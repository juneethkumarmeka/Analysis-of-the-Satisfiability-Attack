module basic_3000_30000_3500_150_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1476,In_1554);
xnor U1 (N_1,In_1488,In_2367);
xnor U2 (N_2,In_1650,In_1443);
and U3 (N_3,In_1292,In_144);
nor U4 (N_4,In_80,In_325);
or U5 (N_5,In_1109,In_2731);
and U6 (N_6,In_2038,In_2173);
xnor U7 (N_7,In_695,In_2845);
or U8 (N_8,In_2234,In_1944);
xnor U9 (N_9,In_2469,In_32);
or U10 (N_10,In_2255,In_419);
nand U11 (N_11,In_408,In_2105);
xor U12 (N_12,In_1841,In_1898);
nor U13 (N_13,In_915,In_2034);
or U14 (N_14,In_2870,In_2466);
nand U15 (N_15,In_158,In_149);
or U16 (N_16,In_612,In_2702);
nor U17 (N_17,In_2370,In_2829);
nand U18 (N_18,In_9,In_2736);
xnor U19 (N_19,In_572,In_916);
nand U20 (N_20,In_1729,In_2347);
xor U21 (N_21,In_2729,In_2429);
and U22 (N_22,In_2265,In_1927);
or U23 (N_23,In_369,In_181);
or U24 (N_24,In_2438,In_660);
nor U25 (N_25,In_2911,In_518);
nand U26 (N_26,In_1696,In_1722);
nand U27 (N_27,In_2812,In_2099);
nand U28 (N_28,In_287,In_1387);
and U29 (N_29,In_364,In_2758);
and U30 (N_30,In_1087,In_634);
nor U31 (N_31,In_1577,In_1874);
xor U32 (N_32,In_1669,In_63);
nor U33 (N_33,In_2409,In_1450);
or U34 (N_34,In_2546,In_1594);
xnor U35 (N_35,In_963,In_1455);
nor U36 (N_36,In_1500,In_753);
xnor U37 (N_37,In_1842,In_2869);
nor U38 (N_38,In_1950,In_2672);
nand U39 (N_39,In_398,In_839);
and U40 (N_40,In_1025,In_681);
nand U41 (N_41,In_2593,In_2396);
or U42 (N_42,In_445,In_1578);
or U43 (N_43,In_969,In_2228);
nor U44 (N_44,In_2144,In_2571);
and U45 (N_45,In_2839,In_1120);
or U46 (N_46,In_44,In_768);
and U47 (N_47,In_866,In_2020);
nand U48 (N_48,In_998,In_2164);
xnor U49 (N_49,In_1561,In_757);
nor U50 (N_50,In_2796,In_35);
nand U51 (N_51,In_1035,In_2909);
xor U52 (N_52,In_2541,In_674);
nor U53 (N_53,In_2956,In_647);
nand U54 (N_54,In_2264,In_377);
nor U55 (N_55,In_1034,In_1308);
or U56 (N_56,In_2786,In_462);
or U57 (N_57,In_250,In_2394);
nand U58 (N_58,In_432,In_262);
nand U59 (N_59,In_781,In_2755);
xor U60 (N_60,In_894,In_2635);
nor U61 (N_61,In_1265,In_1220);
or U62 (N_62,In_1834,In_2237);
nor U63 (N_63,In_1851,In_1987);
or U64 (N_64,In_1521,In_2014);
and U65 (N_65,In_1405,In_2292);
and U66 (N_66,In_2441,In_2420);
xnor U67 (N_67,In_814,In_2591);
or U68 (N_68,In_2055,In_2254);
or U69 (N_69,In_844,In_1546);
or U70 (N_70,In_3,In_2949);
and U71 (N_71,In_2775,In_2566);
xnor U72 (N_72,In_2372,In_2093);
xor U73 (N_73,In_172,In_294);
xnor U74 (N_74,In_954,In_605);
and U75 (N_75,In_116,In_204);
nand U76 (N_76,In_1805,In_88);
and U77 (N_77,In_384,In_360);
and U78 (N_78,In_2457,In_2553);
nand U79 (N_79,In_1690,In_210);
or U80 (N_80,In_1095,In_91);
and U81 (N_81,In_1861,In_1624);
nor U82 (N_82,In_2356,In_2003);
nand U83 (N_83,In_2081,In_1013);
or U84 (N_84,In_2133,In_2686);
nor U85 (N_85,In_1002,In_1936);
and U86 (N_86,In_2768,In_884);
and U87 (N_87,In_2841,In_1829);
or U88 (N_88,In_82,In_1062);
nor U89 (N_89,In_1762,In_1133);
xnor U90 (N_90,In_94,In_593);
xor U91 (N_91,In_2083,In_800);
nor U92 (N_92,In_1963,In_2588);
nor U93 (N_93,In_797,In_2414);
nand U94 (N_94,In_2089,In_2279);
nor U95 (N_95,In_2629,In_1891);
and U96 (N_96,In_2669,In_2652);
xor U97 (N_97,In_1089,In_860);
and U98 (N_98,In_1547,In_1528);
and U99 (N_99,In_2910,In_2456);
xor U100 (N_100,In_983,In_981);
and U101 (N_101,In_2387,In_2223);
nand U102 (N_102,In_673,In_1833);
nor U103 (N_103,In_1417,In_553);
nand U104 (N_104,In_1821,In_2865);
nor U105 (N_105,In_2368,In_1247);
and U106 (N_106,In_2345,In_2194);
xnor U107 (N_107,In_2912,In_1313);
nor U108 (N_108,In_2277,In_1518);
xor U109 (N_109,In_1760,In_2739);
or U110 (N_110,In_1667,In_2026);
or U111 (N_111,In_309,In_1341);
and U112 (N_112,In_1465,In_1770);
or U113 (N_113,In_618,In_2946);
or U114 (N_114,In_1117,In_2310);
nand U115 (N_115,In_698,In_1317);
nand U116 (N_116,In_2085,In_688);
nand U117 (N_117,In_2259,In_1931);
or U118 (N_118,In_549,In_2668);
or U119 (N_119,In_1788,In_2101);
xor U120 (N_120,In_2167,In_591);
nor U121 (N_121,In_2516,In_2680);
or U122 (N_122,In_1966,In_174);
nand U123 (N_123,In_2141,In_1668);
nor U124 (N_124,In_2633,In_2421);
or U125 (N_125,In_1092,In_1586);
and U126 (N_126,In_2106,In_1153);
nand U127 (N_127,In_1145,In_2586);
nand U128 (N_128,In_1381,In_552);
and U129 (N_129,In_1765,In_1370);
or U130 (N_130,In_1176,In_1604);
nand U131 (N_131,In_249,In_978);
or U132 (N_132,In_1552,In_550);
xor U133 (N_133,In_2417,In_14);
xnor U134 (N_134,In_2062,In_2204);
xnor U135 (N_135,In_551,In_1969);
nor U136 (N_136,In_1472,In_1263);
and U137 (N_137,In_1910,In_2432);
nand U138 (N_138,In_2091,In_1406);
xnor U139 (N_139,In_2341,In_476);
xor U140 (N_140,In_2470,In_1451);
xnor U141 (N_141,In_506,In_1671);
nor U142 (N_142,In_999,In_2528);
or U143 (N_143,In_2070,In_2494);
nor U144 (N_144,In_285,In_183);
and U145 (N_145,In_1146,In_1279);
and U146 (N_146,In_1325,In_586);
or U147 (N_147,In_477,In_1132);
nor U148 (N_148,In_465,In_525);
nand U149 (N_149,In_155,In_137);
nor U150 (N_150,In_243,In_1490);
and U151 (N_151,In_81,In_2596);
and U152 (N_152,In_2788,In_2051);
nor U153 (N_153,In_2098,In_1203);
and U154 (N_154,In_1453,In_2705);
or U155 (N_155,In_2561,In_789);
xnor U156 (N_156,In_2479,In_2530);
nor U157 (N_157,In_2894,In_1587);
nand U158 (N_158,In_1394,In_217);
or U159 (N_159,In_2005,In_2882);
nor U160 (N_160,In_376,In_90);
nor U161 (N_161,In_1583,In_2542);
nor U162 (N_162,In_2088,In_1234);
or U163 (N_163,In_2886,In_1198);
or U164 (N_164,In_1674,In_1771);
nor U165 (N_165,In_253,In_561);
and U166 (N_166,In_162,In_2132);
nor U167 (N_167,In_2061,In_1457);
and U168 (N_168,In_463,In_2436);
or U169 (N_169,In_617,In_1517);
nor U170 (N_170,In_441,In_1041);
nand U171 (N_171,In_1032,In_1402);
or U172 (N_172,In_1943,In_1345);
xnor U173 (N_173,In_2451,In_2597);
xor U174 (N_174,In_2278,In_1340);
and U175 (N_175,In_75,In_2868);
or U176 (N_176,In_373,In_139);
and U177 (N_177,In_55,In_1868);
nor U178 (N_178,In_691,In_1536);
or U179 (N_179,In_1735,In_2538);
or U180 (N_180,In_2687,In_132);
nor U181 (N_181,In_1609,In_1459);
xnor U182 (N_182,In_433,In_2554);
xor U183 (N_183,In_1714,In_725);
or U184 (N_184,In_824,In_2326);
or U185 (N_185,In_950,In_2227);
or U186 (N_186,In_1123,In_365);
nand U187 (N_187,In_504,In_1243);
nand U188 (N_188,In_540,In_995);
nor U189 (N_189,In_1887,In_1415);
xor U190 (N_190,In_1090,In_357);
xnor U191 (N_191,In_79,In_1818);
nand U192 (N_192,In_2549,In_668);
nand U193 (N_193,In_2033,In_891);
or U194 (N_194,In_671,In_0);
or U195 (N_195,In_2941,In_1661);
and U196 (N_196,In_2,In_2745);
nand U197 (N_197,In_1201,In_2295);
xnor U198 (N_198,In_1923,In_2484);
xor U199 (N_199,In_1195,In_352);
and U200 (N_200,N_75,In_495);
nand U201 (N_201,In_2382,In_2934);
or U202 (N_202,In_875,In_427);
and U203 (N_203,In_2474,In_2426);
nand U204 (N_204,In_106,N_55);
or U205 (N_205,In_2880,In_404);
nor U206 (N_206,In_96,In_558);
nor U207 (N_207,In_592,In_2428);
or U208 (N_208,In_2049,In_153);
nand U209 (N_209,In_2985,N_50);
and U210 (N_210,In_2856,N_89);
and U211 (N_211,In_1638,In_2532);
and U212 (N_212,In_1892,In_1814);
nand U213 (N_213,In_1316,In_1009);
xor U214 (N_214,In_2166,In_2994);
xnor U215 (N_215,In_1018,In_113);
and U216 (N_216,In_621,In_738);
nand U217 (N_217,In_2373,In_604);
nor U218 (N_218,In_641,In_1189);
nor U219 (N_219,In_2071,In_148);
or U220 (N_220,In_2611,N_138);
or U221 (N_221,In_509,In_1662);
and U222 (N_222,In_1258,In_944);
nand U223 (N_223,In_923,In_2163);
xnor U224 (N_224,In_2662,In_2587);
xnor U225 (N_225,In_1896,In_1764);
nor U226 (N_226,In_2996,In_1965);
and U227 (N_227,In_2364,In_1447);
and U228 (N_228,In_1664,In_693);
xor U229 (N_229,In_1767,In_2826);
and U230 (N_230,In_234,N_110);
nor U231 (N_231,In_1723,In_938);
and U232 (N_232,In_188,In_713);
xor U233 (N_233,N_88,N_60);
xor U234 (N_234,N_118,In_1469);
and U235 (N_235,In_2579,In_415);
or U236 (N_236,In_1571,In_1544);
xnor U237 (N_237,In_2047,In_908);
nor U238 (N_238,In_392,In_1021);
xnor U239 (N_239,In_2517,In_1566);
nand U240 (N_240,In_654,N_156);
xnor U241 (N_241,In_2793,In_1449);
and U242 (N_242,In_1623,In_152);
and U243 (N_243,In_565,In_2460);
or U244 (N_244,In_2908,In_1499);
and U245 (N_245,In_1182,In_92);
and U246 (N_246,In_61,In_156);
or U247 (N_247,In_2626,In_1871);
nor U248 (N_248,In_2261,In_901);
or U249 (N_249,In_2817,In_597);
or U250 (N_250,In_2180,In_101);
xor U251 (N_251,In_951,In_1358);
or U252 (N_252,In_1724,In_692);
and U253 (N_253,In_2746,In_1601);
and U254 (N_254,N_65,In_1286);
or U255 (N_255,In_1565,In_2000);
and U256 (N_256,In_348,In_675);
and U257 (N_257,In_645,In_6);
nand U258 (N_258,In_519,In_286);
xnor U259 (N_259,In_469,In_662);
nor U260 (N_260,In_2154,In_304);
xnor U261 (N_261,In_2651,In_2942);
and U262 (N_262,N_16,In_192);
and U263 (N_263,In_1429,In_2784);
xnor U264 (N_264,In_1085,In_2334);
and U265 (N_265,In_535,In_2375);
or U266 (N_266,In_2217,In_2270);
or U267 (N_267,In_1256,In_133);
and U268 (N_268,In_815,In_1428);
xnor U269 (N_269,In_1970,N_132);
nand U270 (N_270,In_1807,In_1192);
nand U271 (N_271,In_1298,In_929);
or U272 (N_272,In_2594,In_602);
xor U273 (N_273,In_1224,In_1477);
xnor U274 (N_274,In_2518,In_2090);
or U275 (N_275,N_168,In_2770);
nand U276 (N_276,In_2054,In_2772);
nor U277 (N_277,In_1504,In_2735);
xnor U278 (N_278,In_1660,In_1548);
nor U279 (N_279,In_581,In_2883);
nor U280 (N_280,N_101,In_380);
xor U281 (N_281,In_2131,In_1050);
and U282 (N_282,In_2673,In_1217);
xnor U283 (N_283,In_175,In_783);
or U284 (N_284,In_828,In_871);
and U285 (N_285,In_1501,In_744);
and U286 (N_286,In_1337,In_2728);
and U287 (N_287,In_1377,In_2903);
xnor U288 (N_288,In_1678,In_233);
nor U289 (N_289,In_1572,In_1766);
or U290 (N_290,In_2681,In_1218);
xnor U291 (N_291,In_2248,In_2001);
xor U292 (N_292,In_2515,N_186);
nor U293 (N_293,In_1437,In_1769);
nand U294 (N_294,In_120,In_1103);
nor U295 (N_295,In_1017,In_168);
xnor U296 (N_296,In_836,In_1493);
nand U297 (N_297,In_490,In_2342);
and U298 (N_298,In_934,In_2275);
xor U299 (N_299,In_598,In_1404);
xor U300 (N_300,N_10,In_1591);
and U301 (N_301,In_1995,In_2677);
nor U302 (N_302,In_2068,In_2505);
nor U303 (N_303,In_1625,N_127);
nor U304 (N_304,In_105,In_643);
nand U305 (N_305,In_297,N_131);
nor U306 (N_306,In_1626,In_1335);
nand U307 (N_307,In_5,In_1481);
nand U308 (N_308,In_1590,In_129);
nor U309 (N_309,In_2329,In_709);
nand U310 (N_310,In_579,In_2161);
and U311 (N_311,In_312,In_2709);
xor U312 (N_312,In_920,In_1354);
xor U313 (N_313,In_2078,In_2358);
or U314 (N_314,In_885,In_639);
xnor U315 (N_315,In_2979,In_399);
nor U316 (N_316,In_2543,In_717);
or U317 (N_317,In_2143,In_510);
nor U318 (N_318,In_2563,In_627);
or U319 (N_319,In_1101,In_657);
or U320 (N_320,N_169,In_2035);
and U321 (N_321,In_40,In_2762);
and U322 (N_322,In_1811,In_1648);
nand U323 (N_323,In_2365,In_1361);
xnor U324 (N_324,In_39,In_497);
nand U325 (N_325,In_769,In_135);
or U326 (N_326,In_2665,In_2932);
or U327 (N_327,In_1332,N_140);
nor U328 (N_328,In_2535,In_2915);
nand U329 (N_329,In_2117,In_1776);
nand U330 (N_330,In_523,In_1413);
xnor U331 (N_331,In_1968,In_2029);
nor U332 (N_332,In_261,In_288);
nor U333 (N_333,N_69,In_2079);
and U334 (N_334,In_2060,In_326);
or U335 (N_335,In_932,In_486);
nor U336 (N_336,In_2641,In_1219);
nand U337 (N_337,In_240,In_1683);
xor U338 (N_338,In_1142,In_883);
and U339 (N_339,In_2306,In_888);
or U340 (N_340,In_346,In_1057);
and U341 (N_341,In_108,In_1116);
nand U342 (N_342,In_140,In_1467);
or U343 (N_343,In_979,In_2262);
and U344 (N_344,In_1560,In_1114);
nand U345 (N_345,In_661,In_1418);
nor U346 (N_346,In_1301,In_58);
or U347 (N_347,In_2556,N_29);
nor U348 (N_348,In_970,In_2574);
or U349 (N_349,In_1000,In_1508);
and U350 (N_350,In_1732,In_531);
or U351 (N_351,In_242,In_1323);
nand U352 (N_352,In_1695,In_1848);
nor U353 (N_353,In_138,In_1040);
nand U354 (N_354,In_748,In_1126);
nor U355 (N_355,In_21,In_1783);
nand U356 (N_356,In_2952,In_2954);
xnor U357 (N_357,In_2119,In_1704);
and U358 (N_358,In_2599,N_28);
nand U359 (N_359,In_1010,In_2301);
and U360 (N_360,N_153,In_711);
and U361 (N_361,In_1144,In_652);
nor U362 (N_362,N_150,In_1173);
and U363 (N_363,In_19,In_741);
and U364 (N_364,In_2327,In_1971);
and U365 (N_365,In_798,In_2149);
nand U366 (N_366,In_1639,In_2801);
xnor U367 (N_367,In_1734,In_2491);
nor U368 (N_368,In_1348,In_1239);
nor U369 (N_369,In_315,N_98);
nor U370 (N_370,In_1379,In_1775);
nor U371 (N_371,In_1957,In_2854);
and U372 (N_372,In_1366,In_595);
or U373 (N_373,In_2064,In_2723);
nor U374 (N_374,In_1232,In_2448);
or U375 (N_375,In_636,In_2385);
and U376 (N_376,In_2961,In_669);
nand U377 (N_377,In_1640,In_2096);
and U378 (N_378,In_2348,In_2285);
nor U379 (N_379,In_1756,In_2125);
nand U380 (N_380,In_2121,In_374);
xor U381 (N_381,In_2076,In_1593);
or U382 (N_382,In_178,In_2699);
nor U383 (N_383,In_1024,In_564);
xor U384 (N_384,In_2581,In_2468);
nand U385 (N_385,In_2754,In_11);
nor U386 (N_386,In_1642,In_903);
nand U387 (N_387,In_699,N_147);
nand U388 (N_388,In_2339,In_1633);
and U389 (N_389,In_2338,In_1386);
and U390 (N_390,In_2465,In_557);
and U391 (N_391,In_62,In_265);
nor U392 (N_392,In_1634,In_2065);
or U393 (N_393,N_197,In_1044);
nor U394 (N_394,In_864,In_511);
or U395 (N_395,In_2190,In_1152);
nand U396 (N_396,In_1353,In_447);
and U397 (N_397,In_568,In_405);
nor U398 (N_398,In_947,In_791);
nand U399 (N_399,In_2160,In_1495);
and U400 (N_400,In_1259,In_494);
xor U401 (N_401,In_2608,In_2219);
and U402 (N_402,In_2127,In_1863);
and U403 (N_403,In_1761,In_2398);
and U404 (N_404,N_295,In_1549);
xor U405 (N_405,In_2388,In_910);
nor U406 (N_406,In_1885,In_1779);
nor U407 (N_407,In_2239,N_315);
nand U408 (N_408,In_52,In_2963);
nor U409 (N_409,N_319,N_53);
xor U410 (N_410,In_2010,In_2097);
and U411 (N_411,N_196,In_1058);
or U412 (N_412,In_1712,In_1419);
nand U413 (N_413,In_23,In_2455);
nor U414 (N_414,In_1331,In_501);
and U415 (N_415,In_1533,In_1945);
nand U416 (N_416,In_2244,In_913);
and U417 (N_417,In_2811,In_2907);
nor U418 (N_418,In_1797,In_2756);
xnor U419 (N_419,In_1390,In_213);
and U420 (N_420,In_2463,In_865);
nor U421 (N_421,In_1520,In_1906);
nand U422 (N_422,In_56,In_2893);
nand U423 (N_423,In_889,In_2328);
or U424 (N_424,In_2795,In_248);
nor U425 (N_425,In_2011,In_1427);
and U426 (N_426,In_131,In_1351);
and U427 (N_427,In_2782,N_102);
nand U428 (N_428,In_1691,In_608);
or U429 (N_429,In_2998,In_2531);
or U430 (N_430,In_724,In_1854);
nor U431 (N_431,In_1986,In_1038);
nand U432 (N_432,In_1374,N_380);
nand U433 (N_433,N_220,In_206);
or U434 (N_434,In_2130,In_2969);
or U435 (N_435,In_1599,In_629);
nand U436 (N_436,In_2304,In_1793);
and U437 (N_437,In_1154,In_543);
nor U438 (N_438,N_243,In_830);
nand U439 (N_439,In_1180,In_1519);
nor U440 (N_440,In_2986,In_2697);
or U441 (N_441,In_2386,In_232);
nand U442 (N_442,In_1302,N_268);
xnor U443 (N_443,In_776,In_587);
nor U444 (N_444,In_2748,In_1974);
and U445 (N_445,In_2848,In_2140);
and U446 (N_446,In_1107,In_1065);
nand U447 (N_447,In_1082,In_842);
nand U448 (N_448,In_873,In_2073);
nor U449 (N_449,In_1532,N_162);
nor U450 (N_450,In_1605,In_282);
or U451 (N_451,In_255,In_122);
nand U452 (N_452,In_556,In_2926);
nor U453 (N_453,In_2760,In_2240);
and U454 (N_454,In_2437,In_925);
nor U455 (N_455,In_2260,In_2246);
nor U456 (N_456,In_161,In_1270);
and U457 (N_457,In_1365,In_2233);
or U458 (N_458,In_705,In_2767);
nor U459 (N_459,In_1312,In_1226);
nand U460 (N_460,In_560,In_1135);
or U461 (N_461,N_385,In_1251);
and U462 (N_462,In_2852,In_2102);
xnor U463 (N_463,In_87,In_1597);
xor U464 (N_464,In_1272,In_2314);
and U465 (N_465,In_1570,In_60);
xnor U466 (N_466,In_1260,In_2333);
xor U467 (N_467,In_154,In_1478);
and U468 (N_468,In_1815,In_566);
or U469 (N_469,In_704,In_400);
nor U470 (N_470,In_1720,In_1865);
xor U471 (N_471,N_321,In_1952);
or U472 (N_472,In_311,In_505);
and U473 (N_473,In_1649,In_625);
or U474 (N_474,In_291,In_2181);
xor U475 (N_475,In_1847,In_1237);
nor U476 (N_476,In_997,N_182);
and U477 (N_477,In_1707,In_12);
and U478 (N_478,In_1515,In_626);
nand U479 (N_479,In_2846,In_1338);
xnor U480 (N_480,In_750,In_226);
and U481 (N_481,In_994,In_1826);
xnor U482 (N_482,In_1295,N_213);
or U483 (N_483,In_2791,N_37);
and U484 (N_484,In_424,In_1676);
xnor U485 (N_485,In_524,In_194);
nor U486 (N_486,In_1168,In_2427);
and U487 (N_487,In_85,In_1614);
nand U488 (N_488,In_2940,In_457);
or U489 (N_489,In_1894,In_1772);
and U490 (N_490,In_1880,In_2015);
xnor U491 (N_491,In_2012,In_2225);
or U492 (N_492,In_295,In_2918);
xor U493 (N_493,In_235,In_2899);
nand U494 (N_494,In_2006,In_1389);
xor U495 (N_495,In_1229,In_205);
and U496 (N_496,In_193,In_1022);
or U497 (N_497,N_348,In_227);
xor U498 (N_498,In_1327,In_2257);
and U499 (N_499,In_895,In_2603);
or U500 (N_500,In_1291,In_737);
and U501 (N_501,In_931,In_991);
nand U502 (N_502,N_155,In_851);
nor U503 (N_503,In_17,In_2018);
or U504 (N_504,In_1425,In_1080);
and U505 (N_505,In_1271,In_2366);
or U506 (N_506,N_184,In_2445);
xor U507 (N_507,In_1139,In_1737);
nand U508 (N_508,In_54,In_1368);
xnor U509 (N_509,In_258,In_559);
xor U510 (N_510,In_147,In_739);
nor U511 (N_511,In_2743,In_2824);
or U512 (N_512,N_261,In_283);
nor U513 (N_513,In_755,N_250);
nand U514 (N_514,In_846,In_2473);
xor U515 (N_515,In_1104,In_2067);
and U516 (N_516,In_1100,In_2507);
and U517 (N_517,In_2664,In_112);
or U518 (N_518,In_2512,In_1489);
xor U519 (N_519,In_1111,In_1069);
nand U520 (N_520,In_86,In_2488);
xnor U521 (N_521,In_1930,In_2400);
xor U522 (N_522,In_2744,In_343);
or U523 (N_523,In_905,In_2159);
or U524 (N_524,In_1727,In_1924);
or U525 (N_525,In_1812,In_68);
xnor U526 (N_526,In_900,N_208);
nand U527 (N_527,In_2832,In_2769);
xnor U528 (N_528,In_922,In_2609);
nand U529 (N_529,In_2294,N_179);
and U530 (N_530,N_397,In_2241);
nand U531 (N_531,In_2118,In_2890);
or U532 (N_532,In_603,In_2803);
or U533 (N_533,In_2565,In_1787);
xnor U534 (N_534,In_2657,In_2446);
and U535 (N_535,In_1607,N_351);
nor U536 (N_536,In_2268,In_580);
and U537 (N_537,In_631,In_2139);
nor U538 (N_538,In_126,In_906);
and U539 (N_539,In_1199,In_2374);
or U540 (N_540,In_1185,In_431);
and U541 (N_541,In_211,In_1835);
and U542 (N_542,In_2551,In_676);
nor U543 (N_543,In_1458,In_1127);
xnor U544 (N_544,In_1253,In_1531);
nand U545 (N_545,In_2555,N_149);
nand U546 (N_546,In_2742,In_655);
and U547 (N_547,In_2453,In_2108);
and U548 (N_548,In_1267,In_20);
xnor U549 (N_549,In_2972,In_1334);
nand U550 (N_550,In_2607,In_2506);
xor U551 (N_551,In_952,In_416);
and U552 (N_552,N_90,In_123);
xnor U553 (N_553,In_136,In_2562);
or U554 (N_554,In_452,N_368);
nand U555 (N_555,In_1985,N_241);
and U556 (N_556,In_218,In_2525);
nor U557 (N_557,In_2318,In_1978);
and U558 (N_558,In_102,N_383);
nor U559 (N_559,In_1303,In_1551);
and U560 (N_560,N_203,In_2440);
or U561 (N_561,N_276,In_985);
nand U562 (N_562,In_2095,N_267);
nand U563 (N_563,In_1600,N_125);
and U564 (N_564,In_2524,N_157);
and U565 (N_565,In_1837,In_2480);
nand U566 (N_566,N_260,In_1882);
nor U567 (N_567,In_2229,In_458);
and U568 (N_568,In_1073,In_443);
and U569 (N_569,In_2187,In_1221);
xor U570 (N_570,In_199,In_996);
xnor U571 (N_571,In_628,N_165);
and U572 (N_572,In_231,In_2583);
or U573 (N_573,In_853,N_377);
and U574 (N_574,In_1790,In_1984);
and U575 (N_575,In_633,In_401);
or U576 (N_576,In_2849,In_2023);
nand U577 (N_577,N_219,In_664);
nor U578 (N_578,In_2391,In_877);
and U579 (N_579,N_302,In_2416);
nor U580 (N_580,In_2749,N_239);
or U581 (N_581,N_8,N_74);
or U582 (N_582,N_152,In_246);
nand U583 (N_583,In_1193,In_2027);
xnor U584 (N_584,In_2499,In_663);
xor U585 (N_585,In_1392,In_1838);
xor U586 (N_586,In_1610,In_1179);
nor U587 (N_587,In_803,In_177);
or U588 (N_588,In_1036,N_77);
nor U589 (N_589,In_1170,In_1329);
xnor U590 (N_590,In_46,N_214);
or U591 (N_591,In_2497,In_2126);
and U592 (N_592,In_516,In_1911);
or U593 (N_593,In_1928,In_2405);
nand U594 (N_594,N_296,In_2957);
and U595 (N_595,In_2828,In_2544);
nor U596 (N_596,In_182,In_975);
and U597 (N_597,In_324,In_2973);
and U598 (N_598,In_838,In_1194);
nor U599 (N_599,In_1705,In_1976);
xor U600 (N_600,In_1012,In_22);
nor U601 (N_601,In_1914,In_786);
or U602 (N_602,In_807,In_1680);
nand U603 (N_603,In_1763,In_2860);
xor U604 (N_604,In_694,In_254);
nor U605 (N_605,In_646,In_1958);
and U606 (N_606,In_2482,In_833);
nand U607 (N_607,In_2189,N_24);
or U608 (N_608,N_431,In_2874);
nand U609 (N_609,In_735,In_121);
nand U610 (N_610,N_493,N_73);
and U611 (N_611,In_366,In_47);
xnor U612 (N_612,In_902,In_2552);
or U613 (N_613,In_195,In_1191);
or U614 (N_614,In_420,In_1364);
or U615 (N_615,In_1999,In_1411);
xnor U616 (N_616,In_880,N_371);
xnor U617 (N_617,In_2419,In_500);
or U618 (N_618,In_26,In_375);
or U619 (N_619,In_2533,In_973);
and U620 (N_620,In_229,In_1979);
and U621 (N_621,In_1072,In_2293);
xor U622 (N_622,In_1078,N_362);
nand U623 (N_623,In_2175,In_912);
xor U624 (N_624,N_460,In_2124);
xnor U625 (N_625,In_1399,N_137);
xnor U626 (N_626,N_130,N_2);
xor U627 (N_627,In_319,In_1208);
or U628 (N_628,N_562,In_2412);
nand U629 (N_629,In_1227,In_1716);
nand U630 (N_630,In_1689,In_2346);
xor U631 (N_631,In_2842,In_723);
xor U632 (N_632,N_308,In_2211);
or U633 (N_633,In_607,In_1602);
or U634 (N_634,In_1321,In_1921);
or U635 (N_635,N_198,In_2929);
or U636 (N_636,N_297,In_423);
nor U637 (N_637,In_2203,In_1864);
and U638 (N_638,N_223,N_190);
nand U639 (N_639,In_734,N_86);
or U640 (N_640,In_1758,In_1726);
nor U641 (N_641,In_1446,N_404);
nor U642 (N_642,In_749,In_2040);
nand U643 (N_643,In_252,In_1197);
and U644 (N_644,In_2423,In_2514);
and U645 (N_645,In_2286,In_1028);
nor U646 (N_646,In_930,In_2939);
nor U647 (N_647,In_2402,In_2069);
nand U648 (N_648,In_1822,In_808);
nand U649 (N_649,In_2030,In_2776);
nand U650 (N_650,In_1093,In_2443);
nor U651 (N_651,N_393,N_148);
or U652 (N_652,In_2369,In_2316);
nand U653 (N_653,In_329,In_77);
or U654 (N_654,N_201,In_313);
nor U655 (N_655,In_438,In_2464);
xor U656 (N_656,In_2413,In_197);
or U657 (N_657,In_1004,In_2560);
and U658 (N_658,In_1454,In_1975);
xor U659 (N_659,In_2360,In_2726);
xor U660 (N_660,In_498,In_1254);
nor U661 (N_661,In_127,In_539);
or U662 (N_662,In_816,N_440);
and U663 (N_663,In_810,In_2188);
or U664 (N_664,In_1408,N_326);
nor U665 (N_665,In_1524,In_1346);
xor U666 (N_666,N_353,In_2476);
xor U667 (N_667,In_1926,N_463);
or U668 (N_668,In_2982,In_869);
nor U669 (N_669,In_2513,N_579);
nor U670 (N_670,N_506,In_1846);
nor U671 (N_671,In_1456,N_109);
nand U672 (N_672,N_139,N_548);
xnor U673 (N_673,In_70,In_722);
or U674 (N_674,N_30,In_1063);
xor U675 (N_675,In_1148,In_2151);
xnor U676 (N_676,In_1620,In_274);
nor U677 (N_677,N_446,In_2534);
nand U678 (N_678,In_892,N_516);
nor U679 (N_679,In_382,In_341);
and U680 (N_680,In_2733,N_582);
nand U681 (N_681,In_2804,In_1385);
and U682 (N_682,In_1629,In_1768);
or U683 (N_683,In_2297,In_1682);
or U684 (N_684,In_1257,In_2007);
nand U685 (N_685,In_2689,In_601);
nand U686 (N_686,In_1161,N_587);
or U687 (N_687,In_2447,In_1268);
nor U688 (N_688,In_1094,In_2501);
nand U689 (N_689,N_591,In_2224);
nor U690 (N_690,N_501,In_1055);
nand U691 (N_691,In_1037,In_1051);
and U692 (N_692,N_200,In_1523);
or U693 (N_693,N_282,In_2280);
or U694 (N_694,In_2898,In_1980);
nor U695 (N_695,N_426,N_470);
or U696 (N_696,In_124,In_2620);
nor U697 (N_697,In_2287,In_1636);
and U698 (N_698,In_2891,In_858);
xnor U699 (N_699,In_78,In_1129);
nand U700 (N_700,N_305,In_263);
xor U701 (N_701,N_22,In_1574);
and U702 (N_702,In_2645,In_856);
or U703 (N_703,In_1307,In_1096);
or U704 (N_704,In_502,N_500);
nor U705 (N_705,In_1475,N_11);
xor U706 (N_706,In_927,In_436);
or U707 (N_707,In_2621,In_2656);
xor U708 (N_708,In_1698,In_953);
xnor U709 (N_709,In_111,N_369);
or U710 (N_710,In_545,In_1948);
nand U711 (N_711,In_1542,N_154);
xor U712 (N_712,In_1008,In_841);
xor U713 (N_713,In_682,In_1972);
nand U714 (N_714,In_928,In_1172);
nand U715 (N_715,In_1369,In_976);
and U716 (N_716,In_805,In_2357);
or U717 (N_717,In_499,N_85);
or U718 (N_718,In_1916,In_2567);
nand U719 (N_719,In_2258,In_1879);
and U720 (N_720,In_503,In_2250);
or U721 (N_721,In_117,In_809);
or U722 (N_722,In_2232,N_194);
and U723 (N_723,N_61,In_2590);
nand U724 (N_724,In_766,In_2351);
and U725 (N_725,N_427,In_1575);
xor U726 (N_726,In_821,In_95);
nand U727 (N_727,In_703,In_943);
nand U728 (N_728,In_300,In_334);
xor U729 (N_729,In_350,N_329);
or U730 (N_730,In_1448,N_57);
xnor U731 (N_731,In_2660,In_2410);
nor U732 (N_732,In_537,In_1077);
nand U733 (N_733,In_1564,In_2191);
xnor U734 (N_734,In_2251,In_1211);
and U735 (N_735,N_204,In_1907);
xnor U736 (N_736,In_2206,N_474);
xnor U737 (N_737,In_2485,In_2777);
nand U738 (N_738,In_435,In_1494);
nand U739 (N_739,In_1076,In_1982);
nand U740 (N_740,N_346,In_2215);
xor U741 (N_741,In_342,In_1824);
nand U742 (N_742,In_71,In_37);
or U743 (N_743,In_2682,N_122);
nand U744 (N_744,In_1213,In_2344);
nand U745 (N_745,In_2802,In_1171);
xnor U746 (N_746,In_1285,In_1802);
and U747 (N_747,In_848,N_584);
nor U748 (N_748,In_2667,In_2110);
nand U749 (N_749,In_1122,In_770);
and U750 (N_750,In_795,N_453);
and U751 (N_751,In_935,In_2103);
xor U752 (N_752,In_2403,In_2322);
and U753 (N_753,N_465,In_1612);
and U754 (N_754,In_667,In_1395);
and U755 (N_755,In_1214,In_1423);
and U756 (N_756,In_659,In_1383);
and U757 (N_757,In_2462,In_2675);
xor U758 (N_758,In_1960,In_1809);
nor U759 (N_759,In_632,N_211);
and U760 (N_760,In_1615,N_413);
nand U761 (N_761,N_490,In_2177);
xnor U762 (N_762,In_1991,In_2156);
and U763 (N_763,In_2290,In_1266);
nand U764 (N_764,In_1828,In_642);
and U765 (N_765,In_73,In_2866);
or U766 (N_766,In_763,In_2137);
nand U767 (N_767,In_1580,In_1584);
or U768 (N_768,N_62,In_1403);
or U769 (N_769,In_2424,N_327);
or U770 (N_770,In_1973,In_2378);
nor U771 (N_771,In_2631,In_2072);
xor U772 (N_772,In_2162,In_1238);
nor U773 (N_773,In_1954,In_1652);
xor U774 (N_774,In_1487,In_2570);
nand U775 (N_775,In_363,N_256);
and U776 (N_776,In_2013,N_375);
nor U777 (N_777,N_333,N_549);
nor U778 (N_778,In_2335,N_343);
nand U779 (N_779,In_1795,N_66);
xor U780 (N_780,In_2252,In_1844);
and U781 (N_781,In_466,In_1635);
xor U782 (N_782,In_1938,In_2921);
xnor U783 (N_783,In_1042,In_826);
or U784 (N_784,In_610,N_288);
and U785 (N_785,N_189,In_941);
xnor U786 (N_786,In_1981,In_2044);
xor U787 (N_787,In_2605,N_378);
xnor U788 (N_788,N_433,In_989);
nor U789 (N_789,In_245,In_439);
xnor U790 (N_790,In_1915,In_2690);
and U791 (N_791,In_2671,In_1641);
and U792 (N_792,In_269,In_186);
nor U793 (N_793,In_775,N_592);
xnor U794 (N_794,In_609,N_425);
and U795 (N_795,N_278,N_141);
or U796 (N_796,In_620,In_984);
xor U797 (N_797,In_2148,In_1618);
and U798 (N_798,In_412,In_1440);
nor U799 (N_799,N_81,In_2434);
and U800 (N_800,In_1306,In_2897);
nor U801 (N_801,In_679,In_2172);
nand U802 (N_802,In_2389,In_1725);
or U803 (N_803,In_2256,N_357);
and U804 (N_804,N_623,In_1003);
nand U805 (N_805,In_1409,In_1356);
and U806 (N_806,N_104,N_529);
or U807 (N_807,In_759,In_57);
xor U808 (N_808,N_563,In_1901);
or U809 (N_809,In_2838,N_240);
nor U810 (N_810,In_1235,In_2263);
nor U811 (N_811,In_1700,In_471);
xor U812 (N_812,In_1026,N_499);
xnor U813 (N_813,In_1934,In_1988);
xnor U814 (N_814,In_837,In_332);
and U815 (N_815,In_962,N_266);
or U816 (N_816,In_99,In_2582);
nand U817 (N_817,In_1,N_464);
and U818 (N_818,In_2691,In_2509);
or U819 (N_819,In_2114,N_570);
nor U820 (N_820,N_218,In_1595);
and U821 (N_821,In_1831,In_2303);
and U822 (N_822,In_2981,N_534);
nand U823 (N_823,N_777,In_2902);
and U824 (N_824,In_2458,In_1433);
nor U825 (N_825,In_417,In_600);
nor U826 (N_826,In_460,In_247);
nor U827 (N_827,N_310,In_1322);
nor U828 (N_828,In_2041,In_1983);
or U829 (N_829,In_863,In_2235);
and U830 (N_830,In_1410,N_469);
nand U831 (N_831,N_255,In_2325);
xnor U832 (N_832,In_1823,In_2572);
nor U833 (N_833,In_714,In_582);
xnor U834 (N_834,In_2847,In_555);
xor U835 (N_835,N_399,In_1909);
nand U836 (N_836,In_2545,In_1441);
xnor U837 (N_837,N_546,In_710);
nand U838 (N_838,In_792,N_580);
nand U839 (N_839,N_144,In_296);
and U840 (N_840,In_1347,In_2968);
nor U841 (N_841,In_410,In_2100);
and U842 (N_842,In_2823,In_208);
or U843 (N_843,In_2004,In_2877);
nand U844 (N_844,In_496,In_2636);
nor U845 (N_845,In_2578,In_719);
or U846 (N_846,In_806,In_2930);
nor U847 (N_847,N_293,In_353);
or U848 (N_848,In_599,In_1647);
nor U849 (N_849,N_325,N_422);
and U850 (N_850,In_2511,In_2361);
or U851 (N_851,In_1778,In_2613);
nor U852 (N_852,In_1708,In_1016);
nor U853 (N_853,In_1967,In_811);
and U854 (N_854,In_2835,N_669);
nor U855 (N_855,In_1913,In_2618);
and U856 (N_856,In_1684,In_43);
or U857 (N_857,In_2355,In_2688);
xor U858 (N_858,In_986,N_792);
or U859 (N_859,In_2612,In_683);
and U860 (N_860,In_1274,In_179);
nand U861 (N_861,N_773,In_2243);
nand U862 (N_862,In_1052,N_797);
xor U863 (N_863,In_492,In_1514);
nand U864 (N_864,In_649,In_1774);
nand U865 (N_865,N_411,In_2504);
nand U866 (N_866,In_2862,N_417);
nor U867 (N_867,In_146,In_454);
nor U868 (N_868,In_1149,In_1118);
or U869 (N_869,N_778,In_1592);
xnor U870 (N_870,In_2337,N_629);
or U871 (N_871,N_56,In_335);
and U872 (N_872,In_2050,In_1061);
and U873 (N_873,In_1870,In_712);
nand U874 (N_874,In_1319,In_49);
nor U875 (N_875,In_745,In_517);
nand U876 (N_876,N_87,N_586);
xnor U877 (N_877,N_683,In_2780);
xor U878 (N_878,In_730,In_1557);
and U879 (N_879,In_868,In_538);
xor U880 (N_880,In_1442,In_221);
nor U881 (N_881,N_307,In_2273);
nand U882 (N_882,In_1672,In_2025);
nand U883 (N_883,N_347,In_2282);
xnor U884 (N_884,In_2766,In_327);
xor U885 (N_885,In_118,In_2113);
nand U886 (N_886,In_2392,N_694);
xor U887 (N_887,N_555,In_1166);
nor U888 (N_888,In_2500,In_2407);
nand U889 (N_889,In_2135,In_1791);
nor U890 (N_890,In_2821,In_2226);
xnor U891 (N_891,In_1932,In_2195);
or U892 (N_892,In_2152,N_739);
xnor U893 (N_893,In_2266,In_1482);
nor U894 (N_894,N_738,In_1748);
or U895 (N_895,N_568,In_1568);
nand U896 (N_896,In_1773,N_611);
nand U897 (N_897,N_509,In_344);
xor U898 (N_898,In_1352,N_316);
nor U899 (N_899,In_1917,In_2818);
or U900 (N_900,In_1115,In_1020);
or U901 (N_901,In_1873,In_613);
and U902 (N_902,N_389,In_2830);
and U903 (N_903,In_4,N_259);
or U904 (N_904,In_1962,In_2965);
and U905 (N_905,In_1174,In_323);
or U906 (N_906,In_440,In_1471);
xor U907 (N_907,In_1187,In_594);
xor U908 (N_908,In_907,In_1215);
or U909 (N_909,N_13,In_1530);
xnor U910 (N_910,N_655,In_2527);
xor U911 (N_911,In_1786,In_2299);
nand U912 (N_912,In_308,In_189);
xnor U913 (N_913,N_300,N_711);
nand U914 (N_914,In_1740,N_159);
or U915 (N_915,In_1550,N_142);
nand U916 (N_916,In_1645,In_1511);
nor U917 (N_917,N_784,In_2267);
nand U918 (N_918,N_700,N_524);
or U919 (N_919,In_351,N_20);
and U920 (N_920,In_1336,In_1651);
and U921 (N_921,In_716,In_1205);
or U922 (N_922,In_578,N_514);
or U923 (N_923,In_2750,In_1242);
nand U924 (N_924,N_554,In_2785);
and U925 (N_925,N_192,In_2809);
nor U926 (N_926,N_714,In_966);
or U927 (N_927,In_904,N_523);
nand U928 (N_928,In_1382,In_1397);
or U929 (N_929,In_2878,N_191);
nand U930 (N_930,N_108,In_2906);
xor U931 (N_931,In_1430,N_477);
nor U932 (N_932,In_448,In_2142);
xnor U933 (N_933,In_1252,N_269);
nand U934 (N_934,In_115,In_2964);
xnor U935 (N_935,In_758,In_76);
nand U936 (N_936,In_275,N_718);
and U937 (N_937,In_251,In_1105);
nor U938 (N_938,In_2861,In_2487);
nor U939 (N_939,In_955,In_899);
nand U940 (N_940,N_758,N_367);
nand U941 (N_941,In_2340,In_802);
or U942 (N_942,In_1068,In_2642);
nand U943 (N_943,N_445,In_670);
nand U944 (N_944,N_620,In_2418);
nand U945 (N_945,N_473,In_1344);
nor U946 (N_946,In_2057,N_92);
xnor U947 (N_947,In_1250,In_870);
or U948 (N_948,N_666,In_2576);
and U949 (N_949,N_7,In_2028);
nor U950 (N_950,In_2654,In_2425);
or U951 (N_951,N_221,In_2792);
and U952 (N_952,In_2724,In_1169);
nor U953 (N_953,In_2937,In_1752);
and U954 (N_954,In_548,N_522);
xnor U955 (N_955,In_1666,In_1460);
nand U956 (N_956,N_335,N_232);
nand U957 (N_957,In_266,In_371);
nand U958 (N_958,N_598,N_712);
and U959 (N_959,N_113,In_1088);
nand U960 (N_960,In_1810,In_874);
and U961 (N_961,In_230,In_700);
xor U962 (N_962,N_331,In_2837);
nand U963 (N_963,N_656,N_786);
nand U964 (N_964,In_754,In_887);
nand U965 (N_965,In_2205,N_679);
nand U966 (N_966,In_2269,N_719);
xor U967 (N_967,In_2082,N_497);
nor U968 (N_968,In_128,N_116);
or U969 (N_969,N_576,N_704);
nand U970 (N_970,N_419,In_2983);
and U971 (N_971,N_103,In_2676);
nand U972 (N_972,N_699,In_2763);
xnor U973 (N_973,In_2905,N_271);
xnor U974 (N_974,In_241,In_236);
or U975 (N_975,In_512,In_2169);
and U976 (N_976,In_1277,In_854);
xnor U977 (N_977,In_2568,In_2371);
and U978 (N_978,In_574,In_1414);
xnor U979 (N_979,In_1939,In_267);
and U980 (N_980,In_1996,In_1731);
and U981 (N_981,N_4,N_117);
nor U982 (N_982,In_385,In_299);
nor U983 (N_983,In_1432,N_686);
nand U984 (N_984,In_151,In_1742);
xnor U985 (N_985,N_762,In_212);
and U986 (N_986,In_886,N_475);
nand U987 (N_987,N_517,In_696);
xor U988 (N_988,In_130,In_487);
and U989 (N_989,In_1895,N_436);
nor U990 (N_990,N_552,In_1473);
xnor U991 (N_991,N_180,N_143);
xor U992 (N_992,In_1496,N_723);
xnor U993 (N_993,In_157,N_332);
and U994 (N_994,In_544,In_1794);
and U995 (N_995,N_745,In_1850);
xnor U996 (N_996,In_1753,N_312);
and U997 (N_997,N_569,In_2863);
xor U998 (N_998,In_2892,In_1750);
and U999 (N_999,In_1245,In_316);
and U1000 (N_1000,In_18,In_442);
xor U1001 (N_1001,In_1360,N_537);
nor U1002 (N_1002,In_1596,In_395);
nor U1003 (N_1003,N_749,In_1039);
or U1004 (N_1004,In_98,N_258);
or U1005 (N_1005,In_1372,In_402);
and U1006 (N_1006,In_2377,N_476);
nand U1007 (N_1007,In_2978,N_926);
nand U1008 (N_1008,In_2317,In_2363);
xnor U1009 (N_1009,N_481,In_1289);
nand U1010 (N_1010,In_677,In_530);
and U1011 (N_1011,N_951,In_2928);
xor U1012 (N_1012,N_437,N_923);
nor U1013 (N_1013,In_2649,In_1685);
xnor U1014 (N_1014,In_2628,In_1150);
xor U1015 (N_1015,N_969,In_150);
or U1016 (N_1016,In_397,In_2695);
nand U1017 (N_1017,In_2638,N_955);
xor U1018 (N_1018,In_1207,In_2397);
and U1019 (N_1019,N_398,In_69);
or U1020 (N_1020,In_321,In_1576);
xor U1021 (N_1021,N_124,N_817);
nor U1022 (N_1022,In_2519,In_1715);
or U1023 (N_1023,In_2843,N_980);
nor U1024 (N_1024,In_2895,N_967);
and U1025 (N_1025,N_963,In_2332);
nand U1026 (N_1026,N_342,N_750);
and U1027 (N_1027,In_167,N_864);
nor U1028 (N_1028,In_2550,N_919);
or U1029 (N_1029,In_1717,In_388);
nor U1030 (N_1030,In_1659,In_2019);
or U1031 (N_1031,N_942,In_1535);
and U1032 (N_1032,N_870,In_2990);
and U1033 (N_1033,In_1559,N_861);
nand U1034 (N_1034,N_468,N_599);
nor U1035 (N_1035,In_2454,N_622);
nand U1036 (N_1036,N_134,In_2720);
or U1037 (N_1037,In_451,In_508);
and U1038 (N_1038,In_89,In_1287);
nor U1039 (N_1039,In_270,In_968);
and U1040 (N_1040,N_364,In_702);
xnor U1041 (N_1041,In_2401,N_247);
nor U1042 (N_1042,N_225,In_820);
nor U1043 (N_1043,N_107,N_71);
and U1044 (N_1044,N_199,In_2075);
nor U1045 (N_1045,N_237,N_574);
nor U1046 (N_1046,In_303,In_418);
and U1047 (N_1047,In_721,In_2502);
nand U1048 (N_1048,In_614,In_2022);
nand U1049 (N_1049,N_292,In_2887);
or U1050 (N_1050,N_439,In_2478);
nand U1051 (N_1051,In_1165,In_411);
xor U1052 (N_1052,In_2970,N_847);
xnor U1053 (N_1053,In_1658,In_567);
nor U1054 (N_1054,In_937,N_172);
and U1055 (N_1055,N_697,In_992);
xor U1056 (N_1056,In_867,In_2959);
nand U1057 (N_1057,In_238,In_2741);
and U1058 (N_1058,N_234,N_525);
or U1059 (N_1059,In_515,In_1497);
and U1060 (N_1060,In_2045,In_485);
or U1061 (N_1061,N_972,N_573);
xor U1062 (N_1062,In_1516,In_1998);
and U1063 (N_1063,N_930,In_455);
nand U1064 (N_1064,In_2622,N_949);
xor U1065 (N_1065,N_105,In_2624);
and U1066 (N_1066,In_876,In_514);
nand U1067 (N_1067,In_1946,N_698);
nand U1068 (N_1068,In_767,N_688);
and U1069 (N_1069,N_593,In_2221);
and U1070 (N_1070,In_1461,In_1184);
xnor U1071 (N_1071,In_2585,In_1158);
xor U1072 (N_1072,In_2913,N_402);
nand U1073 (N_1073,In_2107,N_806);
nand U1074 (N_1074,N_605,In_665);
or U1075 (N_1075,In_2002,In_430);
nor U1076 (N_1076,N_982,In_100);
xor U1077 (N_1077,In_2569,In_2422);
xnor U1078 (N_1078,In_2122,N_791);
and U1079 (N_1079,N_361,In_2111);
nand U1080 (N_1080,N_280,N_513);
xor U1081 (N_1081,In_2309,In_1859);
nor U1082 (N_1082,N_94,In_2381);
xnor U1083 (N_1083,In_2859,N_63);
or U1084 (N_1084,N_320,In_2925);
or U1085 (N_1085,In_2712,In_1159);
nor U1086 (N_1086,In_1912,In_2059);
nand U1087 (N_1087,In_281,In_2974);
nor U1088 (N_1088,In_1782,In_1759);
or U1089 (N_1089,In_1919,In_1143);
xor U1090 (N_1090,In_1097,In_1628);
xor U1091 (N_1091,In_2222,N_992);
nand U1092 (N_1092,In_1074,N_350);
nor U1093 (N_1093,In_1241,N_810);
and U1094 (N_1094,In_1806,In_2816);
nor U1095 (N_1095,In_2171,In_936);
nand U1096 (N_1096,In_489,In_2698);
xor U1097 (N_1097,In_1177,In_414);
nor U1098 (N_1098,In_526,N_798);
xnor U1099 (N_1099,In_425,In_958);
nand U1100 (N_1100,In_2876,In_2962);
and U1101 (N_1101,In_2799,In_2604);
or U1102 (N_1102,In_1412,In_2230);
nand U1103 (N_1103,In_606,N_510);
nor U1104 (N_1104,In_1738,In_2056);
nor U1105 (N_1105,In_413,In_2717);
and U1106 (N_1106,N_803,In_190);
nor U1107 (N_1107,N_761,In_1739);
nand U1108 (N_1108,In_2885,In_2084);
nand U1109 (N_1109,In_2639,In_1581);
xnor U1110 (N_1110,In_1255,In_1045);
xor U1111 (N_1111,N_167,In_2354);
nand U1112 (N_1112,N_881,In_2300);
nand U1113 (N_1113,In_284,In_1869);
xor U1114 (N_1114,In_653,N_672);
nor U1115 (N_1115,In_2431,In_1933);
nand U1116 (N_1116,N_451,N_627);
and U1117 (N_1117,In_857,In_897);
and U1118 (N_1118,In_2703,In_1777);
nand U1119 (N_1119,In_1693,N_345);
and U1120 (N_1120,In_456,N_421);
and U1121 (N_1121,In_2577,In_2492);
nand U1122 (N_1122,In_678,In_215);
and U1123 (N_1123,N_854,N_814);
nand U1124 (N_1124,In_2610,N_866);
nor U1125 (N_1125,In_1903,In_2298);
or U1126 (N_1126,In_2145,In_638);
or U1127 (N_1127,In_1573,In_1378);
nor U1128 (N_1128,In_2305,In_2548);
or U1129 (N_1129,In_1529,In_1027);
nand U1130 (N_1130,N_678,N_630);
xor U1131 (N_1131,In_879,N_933);
and U1132 (N_1132,In_7,In_2058);
or U1133 (N_1133,In_684,N_748);
nor U1134 (N_1134,N_939,In_1019);
nand U1135 (N_1135,N_747,In_481);
nand U1136 (N_1136,In_391,N_133);
and U1137 (N_1137,In_1479,In_780);
xor U1138 (N_1138,In_2288,N_290);
xnor U1139 (N_1139,N_207,N_226);
and U1140 (N_1140,In_474,In_2123);
nand U1141 (N_1141,In_2520,In_1261);
or U1142 (N_1142,In_2218,In_1262);
nor U1143 (N_1143,In_1875,In_220);
nand U1144 (N_1144,In_1688,N_457);
nand U1145 (N_1145,In_1922,N_311);
nand U1146 (N_1146,In_2201,N_0);
or U1147 (N_1147,In_2917,N_526);
nor U1148 (N_1148,In_2889,In_239);
or U1149 (N_1149,In_2302,N_763);
or U1150 (N_1150,N_43,N_482);
and U1151 (N_1151,In_2798,In_1498);
and U1152 (N_1152,In_2584,In_84);
nand U1153 (N_1153,In_855,N_952);
nand U1154 (N_1154,N_18,In_2376);
or U1155 (N_1155,In_1202,In_2016);
nor U1156 (N_1156,N_663,In_50);
nor U1157 (N_1157,In_114,N_171);
and U1158 (N_1158,In_1110,In_1113);
nor U1159 (N_1159,N_730,In_919);
or U1160 (N_1160,N_878,In_2308);
nand U1161 (N_1161,In_1994,N_853);
nand U1162 (N_1162,In_2663,N_382);
or U1163 (N_1163,In_2158,In_2174);
nand U1164 (N_1164,N_76,In_779);
nor U1165 (N_1165,In_507,In_1853);
nand U1166 (N_1166,N_648,N_272);
nand U1167 (N_1167,N_681,In_651);
and U1168 (N_1168,In_459,N_533);
nand U1169 (N_1169,In_1278,N_740);
nor U1170 (N_1170,In_1491,In_1711);
nand U1171 (N_1171,N_456,In_2120);
xor U1172 (N_1172,In_141,N_863);
nand U1173 (N_1173,N_420,N_640);
nand U1174 (N_1174,N_430,N_129);
nor U1175 (N_1175,N_416,N_231);
xor U1176 (N_1176,In_2537,In_1371);
or U1177 (N_1177,In_1124,In_2200);
nor U1178 (N_1178,In_689,In_832);
nor U1179 (N_1179,N_922,N_929);
xor U1180 (N_1180,N_813,In_765);
nor U1181 (N_1181,N_899,N_759);
nor U1182 (N_1182,In_176,In_1503);
and U1183 (N_1183,N_444,In_2558);
nand U1184 (N_1184,In_1098,N_617);
or U1185 (N_1185,In_1297,N_624);
nand U1186 (N_1186,In_2032,In_1468);
nor U1187 (N_1187,N_571,In_1209);
nor U1188 (N_1188,N_265,In_896);
and U1189 (N_1189,In_2039,In_1632);
and U1190 (N_1190,In_794,N_787);
or U1191 (N_1191,N_423,N_768);
or U1192 (N_1192,In_2738,N_908);
or U1193 (N_1193,In_437,N_917);
nor U1194 (N_1194,N_394,In_1902);
or U1195 (N_1195,N_151,N_956);
and U1196 (N_1196,In_1655,N_64);
xor U1197 (N_1197,In_611,In_2984);
xnor U1198 (N_1198,N_40,N_680);
nand U1199 (N_1199,N_299,In_1400);
xor U1200 (N_1200,N_667,N_491);
and U1201 (N_1201,N_1102,In_909);
or U1202 (N_1202,In_355,In_2716);
or U1203 (N_1203,N_724,In_1947);
nand U1204 (N_1204,N_845,In_1435);
nor U1205 (N_1205,In_829,N_503);
xnor U1206 (N_1206,N_181,N_1072);
xnor U1207 (N_1207,In_30,In_1196);
or U1208 (N_1208,N_435,In_2510);
or U1209 (N_1209,N_274,In_2283);
nand U1210 (N_1210,In_672,In_1883);
nand U1211 (N_1211,N_844,In_2080);
nand U1212 (N_1212,N_210,N_673);
and U1213 (N_1213,N_944,In_822);
and U1214 (N_1214,N_753,In_686);
nor U1215 (N_1215,N_628,N_1130);
and U1216 (N_1216,N_543,N_1061);
or U1217 (N_1217,N_690,N_953);
and U1218 (N_1218,N_164,N_384);
or U1219 (N_1219,N_486,In_222);
and U1220 (N_1220,In_2503,In_2888);
or U1221 (N_1221,In_1866,In_1754);
nor U1222 (N_1222,In_1086,N_54);
and U1223 (N_1223,In_2976,N_772);
nand U1224 (N_1224,In_301,N_508);
or U1225 (N_1225,N_606,In_2707);
nand U1226 (N_1226,N_432,In_1631);
xor U1227 (N_1227,In_2920,N_462);
xor U1228 (N_1228,In_2336,N_1038);
nor U1229 (N_1229,N_400,In_774);
and U1230 (N_1230,N_233,N_957);
and U1231 (N_1231,In_1878,In_2683);
or U1232 (N_1232,In_2430,In_180);
or U1233 (N_1233,N_495,In_2647);
nor U1234 (N_1234,In_354,In_1160);
xnor U1235 (N_1235,N_886,In_1373);
nor U1236 (N_1236,In_1990,In_946);
or U1237 (N_1237,In_728,N_1063);
or U1238 (N_1238,In_1908,N_472);
nor U1239 (N_1239,N_254,In_773);
and U1240 (N_1240,In_2630,N_294);
nand U1241 (N_1241,In_573,In_1318);
nor U1242 (N_1242,N_374,N_691);
or U1243 (N_1243,N_1165,N_1104);
nand U1244 (N_1244,N_1106,In_2722);
and U1245 (N_1245,In_200,In_637);
xor U1246 (N_1246,N_945,In_898);
and U1247 (N_1247,N_187,N_937);
and U1248 (N_1248,In_2168,In_697);
or U1249 (N_1249,N_936,In_2196);
nor U1250 (N_1250,N_406,N_572);
nor U1251 (N_1251,In_1579,N_41);
nand U1252 (N_1252,N_634,In_264);
nor U1253 (N_1253,In_2245,N_641);
nand U1254 (N_1254,N_304,In_1656);
xnor U1255 (N_1255,In_1800,In_166);
or U1256 (N_1256,In_1706,In_125);
nor U1257 (N_1257,In_184,N_682);
nor U1258 (N_1258,N_999,N_868);
nor U1259 (N_1259,In_1054,N_273);
nand U1260 (N_1260,In_338,In_1697);
nor U1261 (N_1261,N_544,N_1111);
xor U1262 (N_1262,In_1162,In_1920);
nand U1263 (N_1263,N_1029,In_104);
nor U1264 (N_1264,In_2209,In_1102);
xnor U1265 (N_1265,N_872,In_2806);
nand U1266 (N_1266,N_706,N_909);
nor U1267 (N_1267,In_2210,N_692);
or U1268 (N_1268,In_2199,In_378);
xnor U1269 (N_1269,N_418,N_1136);
xnor U1270 (N_1270,N_852,N_889);
or U1271 (N_1271,N_1185,In_1675);
and U1272 (N_1272,N_1193,In_2390);
nor U1273 (N_1273,N_484,N_285);
and U1274 (N_1274,N_670,In_732);
xor U1275 (N_1275,In_1643,N_45);
nand U1276 (N_1276,In_302,In_882);
nand U1277 (N_1277,N_1090,N_59);
xor U1278 (N_1278,In_320,In_1803);
nor U1279 (N_1279,N_743,In_1701);
nand U1280 (N_1280,N_877,N_961);
xor U1281 (N_1281,N_334,N_370);
or U1282 (N_1282,N_415,In_2881);
xnor U1283 (N_1283,In_2819,In_1029);
nand U1284 (N_1284,In_2231,In_2564);
nand U1285 (N_1285,In_747,In_119);
xor U1286 (N_1286,In_1188,In_2700);
or U1287 (N_1287,In_2138,N_642);
and U1288 (N_1288,In_845,N_1115);
or U1289 (N_1289,In_918,N_3);
nor U1290 (N_1290,In_28,N_550);
xor U1291 (N_1291,In_1534,N_328);
xnor U1292 (N_1292,In_2493,N_729);
nor U1293 (N_1293,N_1189,In_209);
and U1294 (N_1294,In_1603,N_1062);
or U1295 (N_1295,In_2924,In_1749);
nor U1296 (N_1296,In_1248,N_166);
and U1297 (N_1297,In_2475,N_502);
or U1298 (N_1298,In_1264,N_352);
or U1299 (N_1299,In_1121,N_47);
and U1300 (N_1300,In_1134,N_479);
or U1301 (N_1301,In_1747,In_1567);
or U1302 (N_1302,In_563,N_891);
or U1303 (N_1303,In_2619,In_2950);
or U1304 (N_1304,In_1721,In_2496);
or U1305 (N_1305,N_556,In_2086);
nand U1306 (N_1306,N_496,In_1733);
nand U1307 (N_1307,N_645,N_49);
and U1308 (N_1308,In_2831,In_2192);
nand U1309 (N_1309,In_1622,N_478);
xnor U1310 (N_1310,N_818,In_2975);
nand U1311 (N_1311,In_948,N_839);
or U1312 (N_1312,In_2694,In_322);
or U1313 (N_1313,In_771,N_363);
xor U1314 (N_1314,In_982,In_93);
nand U1315 (N_1315,In_331,N_390);
or U1316 (N_1316,N_1002,N_671);
and U1317 (N_1317,N_1164,In_2008);
nor U1318 (N_1318,N_808,N_983);
or U1319 (N_1319,In_2208,In_2617);
nand U1320 (N_1320,In_1416,In_1718);
xnor U1321 (N_1321,In_965,In_64);
xnor U1322 (N_1322,N_1044,In_2827);
and U1323 (N_1323,N_1127,In_2980);
or U1324 (N_1324,In_2640,N_947);
or U1325 (N_1325,In_993,In_1949);
or U1326 (N_1326,In_31,N_193);
or U1327 (N_1327,N_1131,N_216);
nor U1328 (N_1328,N_635,N_1073);
nand U1329 (N_1329,N_767,In_1611);
xnor U1330 (N_1330,In_2678,In_2477);
nor U1331 (N_1331,N_918,N_687);
xnor U1332 (N_1332,In_1856,In_1466);
xor U1333 (N_1333,N_589,In_8);
nand U1334 (N_1334,In_2794,In_493);
and U1335 (N_1335,In_1483,N_1031);
and U1336 (N_1336,In_2415,In_2053);
and U1337 (N_1337,In_185,In_2960);
nand U1338 (N_1338,In_453,In_191);
or U1339 (N_1339,N_424,N_717);
nand U1340 (N_1340,N_42,In_13);
and U1341 (N_1341,In_2810,In_2547);
or U1342 (N_1342,In_1075,In_1431);
xnor U1343 (N_1343,N_602,In_2176);
and U1344 (N_1344,In_2242,In_1627);
or U1345 (N_1345,N_867,In_1156);
xnor U1346 (N_1346,In_2790,N_1151);
or U1347 (N_1347,N_106,N_217);
and U1348 (N_1348,In_1858,In_2759);
or U1349 (N_1349,N_608,N_317);
and U1350 (N_1350,In_1426,N_1037);
or U1351 (N_1351,In_2704,In_2896);
or U1352 (N_1352,In_1140,In_990);
and U1353 (N_1353,In_2589,In_1081);
nor U1354 (N_1354,In_1210,N_977);
and U1355 (N_1355,N_1191,N_1018);
nor U1356 (N_1356,In_596,In_1872);
nor U1357 (N_1357,N_263,N_931);
nand U1358 (N_1358,In_2879,N_1145);
and U1359 (N_1359,In_1147,N_975);
xnor U1360 (N_1360,In_1525,In_42);
nand U1361 (N_1361,N_809,In_1589);
or U1362 (N_1362,In_2313,N_851);
nor U1363 (N_1363,In_483,N_1050);
or U1364 (N_1364,N_904,N_387);
nand U1365 (N_1365,In_2134,N_684);
nand U1366 (N_1366,In_1309,N_67);
nor U1367 (N_1367,N_974,In_1654);
nor U1368 (N_1368,In_2857,In_450);
nand U1369 (N_1369,In_1918,In_51);
and U1370 (N_1370,In_2526,In_2197);
xnor U1371 (N_1371,In_1311,In_793);
and U1372 (N_1372,In_491,N_707);
or U1373 (N_1373,In_2395,In_1839);
xor U1374 (N_1374,N_920,In_1867);
xnor U1375 (N_1375,N_1118,In_2951);
or U1376 (N_1376,N_1139,N_349);
nand U1377 (N_1377,N_979,In_949);
xnor U1378 (N_1378,N_820,N_1080);
xor U1379 (N_1379,In_2052,N_96);
xor U1380 (N_1380,N_507,N_941);
nand U1381 (N_1381,In_336,In_1225);
or U1382 (N_1382,N_804,N_826);
or U1383 (N_1383,N_647,In_2711);
or U1384 (N_1384,In_1997,N_737);
nand U1385 (N_1385,N_1194,In_1276);
nand U1386 (N_1386,In_2249,N_1074);
nand U1387 (N_1387,In_1886,N_1010);
nor U1388 (N_1388,In_276,In_1730);
and U1389 (N_1389,In_328,N_595);
and U1390 (N_1390,In_1904,In_2557);
xor U1391 (N_1391,N_822,N_693);
and U1392 (N_1392,In_546,In_2320);
nand U1393 (N_1393,In_861,N_236);
or U1394 (N_1394,In_571,In_1687);
nor U1395 (N_1395,In_2807,In_1959);
nand U1396 (N_1396,N_1043,N_821);
xor U1397 (N_1397,N_489,N_906);
nand U1398 (N_1398,N_1171,In_1703);
and U1399 (N_1399,N_79,N_38);
nand U1400 (N_1400,In_528,In_2778);
xor U1401 (N_1401,In_1231,N_907);
or U1402 (N_1402,N_1094,N_1017);
and U1403 (N_1403,N_31,In_2522);
or U1404 (N_1404,In_1007,N_578);
xor U1405 (N_1405,In_1407,N_1);
nor U1406 (N_1406,N_227,N_229);
or U1407 (N_1407,N_1116,In_1941);
xnor U1408 (N_1408,N_841,N_1250);
and U1409 (N_1409,In_1540,In_2155);
or U1410 (N_1410,In_2383,N_1254);
nand U1411 (N_1411,In_640,In_110);
or U1412 (N_1412,In_2214,In_1434);
xnor U1413 (N_1413,N_1394,In_1112);
and U1414 (N_1414,N_405,N_1367);
xor U1415 (N_1415,N_242,In_942);
and U1416 (N_1416,In_2063,In_2404);
xor U1417 (N_1417,N_1290,N_542);
nand U1418 (N_1418,N_539,In_1893);
nand U1419 (N_1419,N_565,In_2271);
nor U1420 (N_1420,In_2943,N_1344);
or U1421 (N_1421,N_776,In_48);
nand U1422 (N_1422,N_480,In_1084);
xnor U1423 (N_1423,N_1221,N_428);
and U1424 (N_1424,N_52,In_2955);
nor U1425 (N_1425,In_1977,N_832);
or U1426 (N_1426,In_2129,N_1121);
nor U1427 (N_1427,In_788,N_1135);
or U1428 (N_1428,N_1051,N_985);
or U1429 (N_1429,N_1361,In_2851);
xnor U1430 (N_1430,N_1095,In_2411);
nor U1431 (N_1431,N_1152,N_1280);
or U1432 (N_1432,In_429,In_778);
and U1433 (N_1433,In_2043,N_1203);
or U1434 (N_1434,N_1310,N_1153);
nand U1435 (N_1435,N_1387,In_1836);
or U1436 (N_1436,N_610,In_2761);
nor U1437 (N_1437,In_1505,N_206);
nor U1438 (N_1438,In_1083,N_1177);
or U1439 (N_1439,In_367,N_441);
and U1440 (N_1440,In_1033,N_795);
nor U1441 (N_1441,N_454,In_547);
xnor U1442 (N_1442,N_1009,N_1020);
and U1443 (N_1443,N_1319,In_1014);
nor U1444 (N_1444,In_940,In_924);
nand U1445 (N_1445,In_2725,In_1305);
nor U1446 (N_1446,N_998,In_1506);
and U1447 (N_1447,In_852,N_959);
nand U1448 (N_1448,N_1187,In_196);
nor U1449 (N_1449,In_862,N_355);
nand U1450 (N_1450,In_1537,In_273);
or U1451 (N_1451,In_1961,N_1205);
or U1452 (N_1452,N_337,N_788);
or U1453 (N_1453,N_449,In_1230);
or U1454 (N_1454,N_264,N_1081);
and U1455 (N_1455,N_1315,N_1068);
xnor U1456 (N_1456,In_1539,In_2685);
nor U1457 (N_1457,N_1124,In_2343);
nand U1458 (N_1458,In_409,In_2147);
nor U1459 (N_1459,In_488,In_1616);
and U1460 (N_1460,N_654,N_800);
and U1461 (N_1461,N_1314,N_705);
and U1462 (N_1462,N_636,In_1136);
xnor U1463 (N_1463,N_403,In_2666);
or U1464 (N_1464,N_948,N_39);
or U1465 (N_1465,N_1091,In_1556);
xor U1466 (N_1466,N_988,N_726);
nor U1467 (N_1467,In_2853,In_2153);
and U1468 (N_1468,N_21,In_289);
xnor U1469 (N_1469,N_676,N_1273);
xnor U1470 (N_1470,N_1230,N_27);
and U1471 (N_1471,In_272,N_257);
nand U1472 (N_1472,In_305,N_1264);
xnor U1473 (N_1473,In_959,N_1379);
xor U1474 (N_1474,In_1375,N_1070);
xor U1475 (N_1475,N_434,N_303);
and U1476 (N_1476,In_964,In_961);
nor U1477 (N_1477,N_1297,N_783);
or U1478 (N_1478,N_1335,N_1272);
nand U1479 (N_1479,N_722,In_1925);
nor U1480 (N_1480,N_1215,N_1030);
or U1481 (N_1481,In_1630,In_554);
xnor U1482 (N_1482,In_2115,In_2247);
xor U1483 (N_1483,N_1128,N_1351);
xor U1484 (N_1484,In_407,N_1064);
xnor U1485 (N_1485,N_1067,N_632);
and U1486 (N_1486,N_1110,N_970);
nand U1487 (N_1487,In_2953,In_2281);
or U1488 (N_1488,N_668,N_36);
nand U1489 (N_1489,N_1155,In_444);
nor U1490 (N_1490,N_161,N_518);
xnor U1491 (N_1491,N_958,In_624);
nand U1492 (N_1492,In_2872,N_782);
nor U1493 (N_1493,In_1884,N_183);
and U1494 (N_1494,In_2993,N_994);
nand U1495 (N_1495,N_1175,In_859);
nand U1496 (N_1496,In_2178,In_1339);
xor U1497 (N_1497,N_577,In_988);
nand U1498 (N_1498,N_1333,In_2238);
nor U1499 (N_1499,N_1036,In_142);
nor U1500 (N_1500,N_322,N_1262);
or U1501 (N_1501,N_1282,In_1290);
nand U1502 (N_1502,In_2916,In_278);
xor U1503 (N_1503,In_630,In_2721);
or U1504 (N_1504,In_347,N_447);
and U1505 (N_1505,N_1035,In_1043);
and U1506 (N_1506,N_323,In_2814);
or U1507 (N_1507,In_850,N_1066);
or U1508 (N_1508,In_1789,N_703);
xnor U1509 (N_1509,N_1241,In_784);
or U1510 (N_1510,N_1206,In_1509);
nand U1511 (N_1511,N_1381,In_1070);
nor U1512 (N_1512,N_858,In_1246);
or U1513 (N_1513,In_1563,N_1093);
nand U1514 (N_1514,N_356,In_1819);
nor U1515 (N_1515,N_551,In_1813);
and U1516 (N_1516,In_389,In_314);
nor U1517 (N_1517,N_927,N_643);
nand U1518 (N_1518,N_890,In_279);
xnor U1519 (N_1519,N_1079,In_2655);
and U1520 (N_1520,N_960,In_225);
nand U1521 (N_1521,In_1047,In_345);
nand U1522 (N_1522,N_467,In_541);
xnor U1523 (N_1523,N_535,In_2185);
xnor U1524 (N_1524,N_1069,In_2362);
nor U1525 (N_1525,In_2945,N_859);
nand U1526 (N_1526,N_1236,N_665);
nor U1527 (N_1527,In_1108,N_224);
nor U1528 (N_1528,In_479,N_120);
and U1529 (N_1529,N_1256,N_1112);
nand U1530 (N_1530,In_1713,N_195);
nor U1531 (N_1531,N_1011,N_78);
nor U1532 (N_1532,N_849,In_2573);
nand U1533 (N_1533,N_631,In_2967);
nor U1534 (N_1534,N_1301,In_2674);
and U1535 (N_1535,In_570,In_207);
and U1536 (N_1536,N_1075,N_536);
xnor U1537 (N_1537,In_823,N_1045);
and U1538 (N_1538,N_1269,N_741);
nand U1539 (N_1539,N_835,In_1845);
nand U1540 (N_1540,In_1608,In_1507);
nor U1541 (N_1541,N_901,In_1011);
xnor U1542 (N_1542,N_318,In_1825);
or U1543 (N_1543,In_1269,N_275);
or U1544 (N_1544,N_869,In_847);
or U1545 (N_1545,In_2834,N_1014);
xnor U1546 (N_1546,N_928,In_2508);
or U1547 (N_1547,In_1452,N_1279);
nor U1548 (N_1548,N_504,In_2779);
xnor U1549 (N_1549,N_897,N_1046);
nor U1550 (N_1550,N_1233,N_1373);
nor U1551 (N_1551,In_1746,N_564);
xnor U1552 (N_1552,In_1855,In_1064);
nor U1553 (N_1553,N_1022,N_984);
nor U1554 (N_1554,In_1030,N_940);
or U1555 (N_1555,N_1204,In_339);
or U1556 (N_1556,In_1798,N_1318);
and U1557 (N_1557,In_1005,In_1282);
and U1558 (N_1558,In_2324,N_1372);
nand U1559 (N_1559,In_1350,In_2104);
xnor U1560 (N_1560,In_1099,N_248);
or U1561 (N_1561,In_2529,N_1281);
nand U1562 (N_1562,N_1329,N_1242);
or U1563 (N_1563,N_685,N_1006);
nand U1564 (N_1564,In_1677,In_470);
nor U1565 (N_1565,In_1006,In_1138);
or U1566 (N_1566,In_2616,N_360);
nor U1567 (N_1567,In_1299,In_219);
nand U1568 (N_1568,N_964,N_366);
nand U1569 (N_1569,N_968,In_1657);
nand U1570 (N_1570,In_1757,In_2989);
nand U1571 (N_1571,N_862,In_1673);
xor U1572 (N_1572,In_1474,In_1899);
nor U1573 (N_1573,In_782,N_856);
xnor U1574 (N_1574,N_1181,In_259);
xnor U1575 (N_1575,In_482,In_2296);
and U1576 (N_1576,N_1209,In_2606);
nand U1577 (N_1577,In_1736,N_1225);
and U1578 (N_1578,In_1860,N_17);
xnor U1579 (N_1579,In_83,In_2991);
or U1580 (N_1580,In_1422,N_1188);
xnor U1581 (N_1581,In_29,N_1259);
xor U1582 (N_1582,N_396,In_687);
xor U1583 (N_1583,N_1192,In_977);
and U1584 (N_1584,In_2997,N_365);
xor U1585 (N_1585,N_429,In_1200);
nand U1586 (N_1586,N_238,In_2315);
or U1587 (N_1587,N_1244,In_2855);
nor U1588 (N_1588,N_987,In_1066);
and U1589 (N_1589,In_1876,N_531);
nor U1590 (N_1590,In_2900,N_1357);
xnor U1591 (N_1591,N_336,N_751);
or U1592 (N_1592,N_771,N_823);
and U1593 (N_1593,N_245,In_1585);
xnor U1594 (N_1594,In_893,N_1196);
or U1595 (N_1595,In_2444,In_1222);
or U1596 (N_1596,In_160,N_1012);
nand U1597 (N_1597,In_1862,N_545);
or U1598 (N_1598,N_209,N_695);
or U1599 (N_1599,N_244,N_1087);
and U1600 (N_1600,In_473,N_291);
or U1601 (N_1601,N_35,In_202);
xor U1602 (N_1602,In_1646,N_893);
and U1603 (N_1603,N_1492,In_223);
and U1604 (N_1604,N_702,N_1154);
xnor U1605 (N_1605,N_251,In_980);
nand U1606 (N_1606,N_1462,In_1512);
or U1607 (N_1607,N_1585,In_1420);
nand U1608 (N_1608,In_2858,N_158);
xor U1609 (N_1609,N_1416,In_65);
nor U1610 (N_1610,N_1120,In_2653);
or U1611 (N_1611,N_793,N_1382);
nand U1612 (N_1612,N_1451,N_1532);
and U1613 (N_1613,N_801,In_914);
nor U1614 (N_1614,In_1206,In_1310);
nor U1615 (N_1615,N_392,N_1513);
nor U1616 (N_1616,In_2627,In_2433);
or U1617 (N_1617,In_987,N_1414);
xnor U1618 (N_1618,N_1252,N_1396);
xor U1619 (N_1619,N_1507,N_1229);
nand U1620 (N_1620,N_802,In_434);
and U1621 (N_1621,In_2116,N_442);
nand U1622 (N_1622,N_1534,N_1564);
nand U1623 (N_1623,N_1566,N_1412);
xnor U1624 (N_1624,N_270,N_1452);
nand U1625 (N_1625,In_1296,N_1041);
nand U1626 (N_1626,In_1053,N_1501);
and U1627 (N_1627,In_2291,N_1573);
and U1628 (N_1628,N_1100,In_2017);
and U1629 (N_1629,N_340,N_1170);
nand U1630 (N_1630,N_176,N_876);
nor U1631 (N_1631,In_2449,In_2495);
xnor U1632 (N_1632,In_34,In_2757);
nand U1633 (N_1633,N_1366,N_309);
and U1634 (N_1634,N_1234,N_842);
nor U1635 (N_1635,In_812,In_2323);
nand U1636 (N_1636,N_136,In_2540);
nand U1637 (N_1637,N_1475,In_2170);
nand U1638 (N_1638,In_972,N_314);
and U1639 (N_1639,N_1535,N_912);
nand U1640 (N_1640,In_650,N_995);
nand U1641 (N_1641,N_774,N_339);
xor U1642 (N_1642,N_932,In_1527);
xnor U1643 (N_1643,N_659,N_660);
and U1644 (N_1644,N_1013,N_1529);
nor U1645 (N_1645,In_945,In_421);
or U1646 (N_1646,N_1419,N_662);
xnor U1647 (N_1647,In_974,N_1293);
nor U1648 (N_1648,N_1352,N_177);
xor U1649 (N_1649,N_888,In_1955);
xnor U1650 (N_1650,N_830,N_6);
xor U1651 (N_1651,N_1509,In_2864);
and U1652 (N_1652,N_1055,N_1527);
nor U1653 (N_1653,In_635,N_612);
or U1654 (N_1654,In_390,N_44);
nand U1655 (N_1655,N_1422,N_619);
xnor U1656 (N_1656,N_675,In_1067);
nand U1657 (N_1657,In_59,In_467);
and U1658 (N_1658,N_775,N_1321);
or U1659 (N_1659,N_14,In_2650);
nand U1660 (N_1660,N_1444,N_1465);
or U1661 (N_1661,N_395,In_449);
or U1662 (N_1662,In_257,N_1132);
xnor U1663 (N_1663,N_1060,In_2311);
or U1664 (N_1664,N_1576,N_1348);
and U1665 (N_1665,In_911,N_1498);
and U1666 (N_1666,N_119,In_340);
nor U1667 (N_1667,N_819,In_1396);
nand U1668 (N_1668,N_1200,In_1137);
nor U1669 (N_1669,N_1168,N_1494);
or U1670 (N_1670,N_834,N_277);
xor U1671 (N_1671,N_1484,In_1644);
nor U1672 (N_1672,In_2710,N_1157);
nor U1673 (N_1673,N_1082,In_381);
nor U1674 (N_1674,In_827,In_1167);
xor U1675 (N_1675,N_414,In_2815);
nand U1676 (N_1676,N_1407,N_80);
or U1677 (N_1677,In_1681,N_174);
nor U1678 (N_1678,N_1593,In_143);
nor U1679 (N_1679,N_1567,N_1485);
xor U1680 (N_1680,N_1184,In_1048);
or U1681 (N_1681,N_756,N_1163);
nand U1682 (N_1682,In_2284,N_1078);
nand U1683 (N_1683,In_1796,In_2274);
or U1684 (N_1684,In_2732,In_804);
xor U1685 (N_1685,In_2467,N_993);
and U1686 (N_1686,N_450,N_1424);
nand U1687 (N_1687,In_2992,N_1320);
nor U1688 (N_1688,N_289,In_228);
or U1689 (N_1689,In_680,N_381);
and U1690 (N_1690,N_1086,In_1744);
nand U1691 (N_1691,In_761,N_1349);
and U1692 (N_1692,N_494,N_1114);
xor U1693 (N_1693,In_733,N_857);
and U1694 (N_1694,N_971,In_171);
nor U1695 (N_1695,N_298,In_2042);
or U1696 (N_1696,N_613,N_696);
and U1697 (N_1697,N_1331,In_1679);
xnor U1698 (N_1698,N_966,In_1304);
nor U1699 (N_1699,N_1584,In_890);
xor U1700 (N_1700,N_1544,In_569);
xnor U1701 (N_1701,N_1467,N_1480);
or U1702 (N_1702,N_638,N_1032);
or U1703 (N_1703,In_1391,N_1561);
xor U1704 (N_1704,N_1228,In_2771);
xor U1705 (N_1705,In_2435,In_1436);
xnor U1706 (N_1706,In_2471,In_464);
nand U1707 (N_1707,N_1240,N_1007);
nand U1708 (N_1708,In_2740,In_2966);
nor U1709 (N_1709,In_1320,N_1308);
nand U1710 (N_1710,N_1496,In_2873);
nor U1711 (N_1711,In_790,In_372);
and U1712 (N_1712,In_2901,N_1528);
nor U1713 (N_1713,N_70,N_1458);
or U1714 (N_1714,N_1393,In_666);
xnor U1715 (N_1715,N_1156,In_74);
nor U1716 (N_1716,N_1299,N_1021);
and U1717 (N_1717,N_900,In_53);
xnor U1718 (N_1718,In_358,N_1506);
and U1719 (N_1719,N_1368,N_1516);
nor U1720 (N_1720,N_1355,N_596);
or U1721 (N_1721,N_976,N_1238);
nand U1722 (N_1722,In_1781,In_2349);
or U1723 (N_1723,N_1300,N_1571);
and U1724 (N_1724,N_1217,In_2461);
nand U1725 (N_1725,N_903,N_990);
nand U1726 (N_1726,N_1085,In_939);
nor U1727 (N_1727,N_1097,N_1138);
nand U1728 (N_1728,N_1176,In_520);
or U1729 (N_1729,N_1572,N_1446);
and U1730 (N_1730,N_558,In_2614);
or U1731 (N_1731,N_1182,N_1531);
nand U1732 (N_1732,In_2066,In_310);
nor U1733 (N_1733,N_1306,N_657);
and U1734 (N_1734,N_1283,N_934);
or U1735 (N_1735,In_2319,N_1391);
or U1736 (N_1736,N_391,N_1580);
xnor U1737 (N_1737,N_746,In_2384);
xnor U1738 (N_1738,N_1302,In_584);
and U1739 (N_1739,N_1574,N_1169);
and U1740 (N_1740,In_1484,In_1249);
and U1741 (N_1741,N_710,N_1243);
or U1742 (N_1742,N_1212,In_198);
or U1743 (N_1743,N_614,In_406);
and U1744 (N_1744,N_1453,N_1015);
nor U1745 (N_1745,In_2836,N_1417);
nor U1746 (N_1746,In_1178,In_562);
and U1747 (N_1747,N_1579,N_896);
nand U1748 (N_1748,In_370,N_170);
and U1749 (N_1749,N_882,N_379);
xor U1750 (N_1750,In_2592,In_1951);
nand U1751 (N_1751,N_581,N_1345);
or U1752 (N_1752,In_2914,N_1161);
or U1753 (N_1753,In_1598,In_2109);
or U1754 (N_1754,In_708,N_1557);
and U1755 (N_1755,In_2797,N_1147);
or U1756 (N_1756,In_2765,In_1522);
or U1757 (N_1757,N_865,In_2999);
or U1758 (N_1758,N_1232,N_286);
nand U1759 (N_1759,N_1546,In_831);
xor U1760 (N_1760,In_1799,In_1294);
and U1761 (N_1761,In_2183,In_2165);
xor U1762 (N_1762,N_1336,In_1485);
and U1763 (N_1763,In_1553,In_271);
or U1764 (N_1764,In_2938,In_1543);
nor U1765 (N_1765,N_1271,In_2399);
nand U1766 (N_1766,In_1281,N_408);
xnor U1767 (N_1767,In_2701,In_2813);
xnor U1768 (N_1768,N_557,N_1477);
nand U1769 (N_1769,In_1463,N_805);
xor U1770 (N_1770,In_2948,N_727);
or U1771 (N_1771,In_306,In_2406);
nand U1772 (N_1772,In_1881,In_393);
and U1773 (N_1773,N_585,N_1303);
nor U1774 (N_1774,N_1178,In_1444);
nor U1775 (N_1775,In_1357,N_1401);
nand U1776 (N_1776,N_1563,In_2359);
nand U1777 (N_1777,N_1195,N_811);
xor U1778 (N_1778,N_128,N_1113);
xnor U1779 (N_1779,N_1219,In_1937);
nor U1780 (N_1780,N_1218,In_2933);
nor U1781 (N_1781,In_10,In_1780);
nand U1782 (N_1782,N_1353,In_1280);
nor U1783 (N_1783,N_1590,N_664);
and U1784 (N_1784,N_1265,N_873);
or U1785 (N_1785,In_2844,N_114);
xor U1786 (N_1786,N_600,In_1929);
or U1787 (N_1787,In_575,N_483);
and U1788 (N_1788,N_1028,N_1479);
or U1789 (N_1789,N_1304,N_528);
or U1790 (N_1790,N_1270,In_1284);
xor U1791 (N_1791,N_1342,In_835);
nor U1792 (N_1792,In_379,In_1362);
xnor U1793 (N_1793,N_1418,N_354);
xor U1794 (N_1794,In_746,In_718);
nand U1795 (N_1795,N_505,N_512);
or U1796 (N_1796,In_726,In_307);
nand U1797 (N_1797,N_650,In_1665);
and U1798 (N_1798,In_170,In_2481);
nand U1799 (N_1799,In_1367,In_762);
nor U1800 (N_1800,N_1325,N_1661);
or U1801 (N_1801,N_1612,In_361);
or U1802 (N_1802,N_991,N_1364);
or U1803 (N_1803,In_825,In_1653);
nand U1804 (N_1804,N_1707,N_1684);
and U1805 (N_1805,In_2995,In_1333);
or U1806 (N_1806,In_1816,N_829);
xnor U1807 (N_1807,N_1720,N_1471);
or U1808 (N_1808,In_2212,In_752);
xnor U1809 (N_1809,N_1675,In_1710);
xnor U1810 (N_1810,N_1713,N_731);
nor U1811 (N_1811,In_840,N_1670);
nor U1812 (N_1812,N_575,In_475);
nand U1813 (N_1813,N_1142,N_1771);
nand U1814 (N_1814,N_827,N_527);
or U1815 (N_1815,N_1278,N_1737);
and U1816 (N_1816,In_533,N_111);
nor U1817 (N_1817,N_58,N_1613);
xor U1818 (N_1818,N_344,N_846);
and U1819 (N_1819,In_1606,N_1326);
and U1820 (N_1820,N_1791,In_2789);
or U1821 (N_1821,N_973,N_1071);
and U1822 (N_1822,N_547,N_1076);
nand U1823 (N_1823,N_1647,In_1792);
xor U1824 (N_1824,In_1421,In_2625);
nand U1825 (N_1825,N_1317,In_2634);
or U1826 (N_1826,In_187,In_1031);
or U1827 (N_1827,N_146,N_1266);
or U1828 (N_1828,N_1739,N_1588);
and U1829 (N_1829,In_1502,N_1753);
or U1830 (N_1830,N_843,N_709);
nor U1831 (N_1831,N_284,N_1350);
or U1832 (N_1832,N_757,N_1313);
nand U1833 (N_1833,N_1552,N_1635);
or U1834 (N_1834,N_1696,N_561);
nor U1835 (N_1835,N_769,In_576);
xor U1836 (N_1836,N_1733,N_1463);
nand U1837 (N_1837,N_1359,N_459);
nand U1838 (N_1838,N_1488,N_1016);
or U1839 (N_1839,N_1665,N_559);
xor U1840 (N_1840,In_787,N_594);
nor U1841 (N_1841,N_1717,N_1277);
nand U1842 (N_1842,N_1117,N_639);
xnor U1843 (N_1843,In_1480,N_1288);
xnor U1844 (N_1844,N_1173,N_1343);
or U1845 (N_1845,N_652,N_1619);
xnor U1846 (N_1846,N_1559,N_1668);
xnor U1847 (N_1847,In_872,N_1482);
and U1848 (N_1848,N_1699,N_51);
and U1849 (N_1849,N_1545,In_2632);
xor U1850 (N_1850,N_649,N_1683);
nor U1851 (N_1851,N_1146,In_97);
nor U1852 (N_1852,N_1049,In_1349);
xnor U1853 (N_1853,In_2787,In_280);
or U1854 (N_1854,In_2489,In_2764);
and U1855 (N_1855,In_2459,N_1540);
nand U1856 (N_1856,In_1992,In_1817);
and U1857 (N_1857,N_916,In_2958);
xor U1858 (N_1858,N_1511,In_2216);
nand U1859 (N_1859,N_1750,N_1503);
and U1860 (N_1860,N_1785,N_1101);
or U1861 (N_1861,In_1380,N_755);
nand U1862 (N_1862,In_1956,N_1211);
and U1863 (N_1863,N_235,In_751);
xnor U1864 (N_1864,N_1466,In_583);
or U1865 (N_1865,In_585,In_1190);
nor U1866 (N_1866,N_1504,N_1766);
nor U1867 (N_1867,In_1993,N_1789);
nor U1868 (N_1868,In_2450,N_874);
xnor U1869 (N_1869,N_633,N_1257);
and U1870 (N_1870,In_2598,N_1674);
xor U1871 (N_1871,In_1857,N_736);
and U1872 (N_1872,In_1273,N_1774);
xor U1873 (N_1873,N_789,N_1727);
xnor U1874 (N_1874,N_1654,In_818);
xor U1875 (N_1875,N_1794,In_521);
nand U1876 (N_1876,N_914,N_1512);
xnor U1877 (N_1877,In_2439,N_1052);
nand U1878 (N_1878,N_376,N_1180);
xnor U1879 (N_1879,N_313,N_1487);
nor U1880 (N_1880,N_540,N_1077);
xor U1881 (N_1881,In_2734,N_1638);
xor U1882 (N_1882,N_1651,N_1415);
and U1883 (N_1883,N_1491,N_1500);
or U1884 (N_1884,N_658,In_878);
nand U1885 (N_1885,In_2330,N_1358);
or U1886 (N_1886,In_1343,In_1613);
xor U1887 (N_1887,N_1762,N_1098);
and U1888 (N_1888,N_1700,N_1123);
nor U1889 (N_1889,N_386,In_318);
nor U1890 (N_1890,N_1449,In_2773);
or U1891 (N_1891,In_2646,In_917);
nor U1892 (N_1892,In_2684,N_1782);
or U1893 (N_1893,In_2236,In_1545);
xor U1894 (N_1894,N_1058,N_1486);
or U1895 (N_1895,N_1772,N_1721);
nand U1896 (N_1896,N_1788,N_1776);
or U1897 (N_1897,In_2714,In_1376);
xor U1898 (N_1898,N_1129,N_742);
xor U1899 (N_1899,N_616,N_1680);
nand U1900 (N_1900,In_616,In_2800);
xnor U1901 (N_1901,N_1723,N_625);
and U1902 (N_1902,N_1213,N_1602);
and U1903 (N_1903,In_1398,N_1311);
or U1904 (N_1904,N_253,N_1143);
or U1905 (N_1905,N_1459,N_1622);
nand U1906 (N_1906,In_1743,N_1141);
nor U1907 (N_1907,N_892,N_287);
and U1908 (N_1908,N_1435,N_653);
xor U1909 (N_1909,In_403,N_1542);
nor U1910 (N_1910,In_72,In_27);
nand U1911 (N_1911,In_2472,N_1538);
xnor U1912 (N_1912,In_2820,N_1653);
xnor U1913 (N_1913,In_277,N_1522);
nand U1914 (N_1914,In_1569,In_777);
nand U1915 (N_1915,N_1553,N_1083);
nor U1916 (N_1916,N_794,N_46);
and U1917 (N_1917,In_173,N_1724);
and U1918 (N_1918,In_2840,N_1442);
nand U1919 (N_1919,N_1202,N_1150);
or U1920 (N_1920,N_1377,In_1001);
and U1921 (N_1921,In_2753,N_1410);
xnor U1922 (N_1922,N_1770,N_1657);
nand U1923 (N_1923,N_1560,N_448);
or U1924 (N_1924,In_1155,N_1740);
nor U1925 (N_1925,In_2833,N_1378);
nand U1926 (N_1926,N_1199,In_292);
nor U1927 (N_1927,In_1621,N_1296);
nand U1928 (N_1928,In_298,In_260);
nor U1929 (N_1929,N_1249,N_1548);
and U1930 (N_1930,N_651,In_834);
nand U1931 (N_1931,N_488,N_1524);
nor U1932 (N_1932,N_840,In_2648);
nor U1933 (N_1933,N_1773,N_1784);
nand U1934 (N_1934,N_1223,N_1757);
and U1935 (N_1935,N_1514,N_1523);
nand U1936 (N_1936,In_203,In_461);
nand U1937 (N_1937,N_590,N_443);
or U1938 (N_1938,In_237,In_2693);
nor U1939 (N_1939,N_1445,N_938);
xor U1940 (N_1940,N_1729,In_1141);
xnor U1941 (N_1941,N_1330,N_1497);
xor U1942 (N_1942,N_721,In_2615);
or U1943 (N_1943,N_1033,N_1054);
and U1944 (N_1944,N_1719,N_1565);
nor U1945 (N_1945,N_1395,In_1877);
or U1946 (N_1946,In_2021,In_2875);
and U1947 (N_1947,N_1339,In_1131);
and U1948 (N_1948,In_2927,N_23);
or U1949 (N_1949,In_956,N_1237);
nor U1950 (N_1950,In_2353,N_796);
or U1951 (N_1951,In_290,In_817);
xor U1952 (N_1952,In_2580,In_1388);
xor U1953 (N_1953,In_577,N_1239);
nor U1954 (N_1954,N_1646,N_1708);
xor U1955 (N_1955,In_1953,In_522);
nand U1956 (N_1956,N_1042,N_1686);
xnor U1957 (N_1957,In_760,N_781);
or U1958 (N_1958,N_1643,N_902);
and U1959 (N_1959,N_1518,In_764);
nor U1960 (N_1960,N_1365,N_1105);
xor U1961 (N_1961,N_1430,N_9);
nand U1962 (N_1962,N_1634,In_658);
or U1963 (N_1963,N_838,In_1244);
and U1964 (N_1964,In_801,In_2321);
and U1965 (N_1965,In_1091,In_333);
and U1966 (N_1966,N_1741,In_2919);
and U1967 (N_1967,In_2307,N_1316);
xor U1968 (N_1968,N_1201,In_1106);
nor U1969 (N_1969,N_1690,N_12);
or U1970 (N_1970,N_306,N_520);
and U1971 (N_1971,N_173,N_1409);
nand U1972 (N_1972,N_1780,N_1263);
and U1973 (N_1973,In_1384,N_1426);
nor U1974 (N_1974,N_1626,In_1617);
or U1975 (N_1975,N_1423,N_1778);
nand U1976 (N_1976,N_1474,In_799);
nor U1977 (N_1977,N_950,N_1607);
nor U1978 (N_1978,N_1639,N_713);
and U1979 (N_1979,N_1652,In_1588);
or U1980 (N_1980,In_2536,In_2092);
or U1981 (N_1981,N_1792,In_2393);
or U1982 (N_1982,In_1300,N_95);
xor U1983 (N_1983,N_1096,N_1667);
and U1984 (N_1984,In_706,N_1411);
xnor U1985 (N_1985,N_135,N_1775);
nand U1986 (N_1986,N_1678,N_674);
or U1987 (N_1987,In_1330,In_656);
nor U1988 (N_1988,N_1630,N_1183);
or U1989 (N_1989,N_766,N_115);
and U1990 (N_1990,N_359,N_452);
nand U1991 (N_1991,N_1658,N_708);
xor U1992 (N_1992,N_1493,N_1758);
and U1993 (N_1993,N_538,N_1671);
nor U1994 (N_1994,N_626,N_790);
and U1995 (N_1995,In_542,N_1227);
nor U1996 (N_1996,N_97,N_1437);
xnor U1997 (N_1997,N_1004,In_1900);
and U1998 (N_1998,N_1371,N_1598);
xor U1999 (N_1999,N_1577,In_513);
and U2000 (N_2000,N_1469,N_1990);
xor U2001 (N_2001,N_1276,In_2805);
or U2002 (N_2002,In_957,N_410);
and U2003 (N_2003,In_1935,N_1831);
xnor U2004 (N_2004,N_1893,N_816);
nand U2005 (N_2005,N_925,N_1998);
and U2006 (N_2006,N_1334,N_1864);
nand U2007 (N_2007,N_1057,N_770);
nor U2008 (N_2008,In_1470,N_1398);
and U2009 (N_2009,N_5,In_1223);
nand U2010 (N_2010,N_1610,N_487);
nor U2011 (N_2011,N_1403,In_2730);
xor U2012 (N_2012,N_1438,N_1508);
and U2013 (N_2013,In_1233,N_1570);
and U2014 (N_2014,N_1900,N_884);
xnor U2015 (N_2015,N_1688,In_2936);
or U2016 (N_2016,N_1827,In_2150);
nor U2017 (N_2017,N_407,N_1003);
and U2018 (N_2018,In_2747,In_1889);
xor U2019 (N_2019,N_1207,N_1460);
nand U2020 (N_2020,In_2198,N_1732);
and U2021 (N_2021,N_1689,N_1380);
xor U2022 (N_2022,In_785,N_962);
nand U2023 (N_2023,N_1669,N_1756);
nor U2024 (N_2024,N_1088,In_2350);
xor U2025 (N_2025,N_93,N_83);
or U2026 (N_2026,N_895,In_2751);
nor U2027 (N_2027,N_1597,N_1374);
or U2028 (N_2028,N_1722,N_1969);
nand U2029 (N_2029,N_1341,N_1384);
or U2030 (N_2030,In_169,In_1637);
nand U2031 (N_2031,N_1938,N_996);
nand U2032 (N_2032,N_1633,In_2692);
nor U2033 (N_2033,N_1167,N_1439);
xor U2034 (N_2034,N_1327,In_1555);
xor U2035 (N_2035,N_1305,N_1231);
nand U2036 (N_2036,N_1197,N_1583);
and U2037 (N_2037,N_1024,In_317);
nand U2038 (N_2038,N_1868,In_1513);
or U2039 (N_2039,N_946,N_1065);
and U2040 (N_2040,N_1681,N_99);
or U2041 (N_2041,N_1604,N_1109);
xor U2042 (N_2042,N_954,N_1805);
and U2043 (N_2043,In_1359,N_1884);
and U2044 (N_2044,N_1470,N_1354);
or U2045 (N_2045,In_2136,In_849);
or U2046 (N_2046,N_1892,N_1850);
and U2047 (N_2047,N_1624,N_1137);
nor U2048 (N_2048,In_742,N_1562);
and U2049 (N_2049,In_2207,N_1994);
xor U2050 (N_2050,In_1820,N_1443);
or U2051 (N_2051,In_394,N_1932);
xnor U2052 (N_2052,N_1911,In_15);
nor U2053 (N_2053,In_268,N_1662);
and U2054 (N_2054,N_1851,In_2193);
nor U2055 (N_2055,N_1873,N_1769);
and U2056 (N_2056,In_163,N_1275);
nand U2057 (N_2057,N_1695,N_1208);
or U2058 (N_2058,N_1744,N_68);
xnor U2059 (N_2059,N_1767,In_1439);
and U2060 (N_2060,N_212,N_1089);
xor U2061 (N_2061,N_760,N_1918);
nor U2062 (N_2062,In_2752,N_1287);
nor U2063 (N_2063,N_860,N_1468);
and U2064 (N_2064,N_1747,In_109);
or U2065 (N_2065,N_338,N_637);
nand U2066 (N_2066,In_1849,N_34);
nand U2067 (N_2067,N_615,N_185);
or U2068 (N_2068,In_720,In_2048);
xnor U2069 (N_2069,In_1510,N_1694);
nand U2070 (N_2070,In_468,N_883);
xnor U2071 (N_2071,N_1925,In_690);
xor U2072 (N_2072,N_924,In_843);
or U2073 (N_2073,N_1582,N_145);
xnor U2074 (N_2074,N_646,N_1781);
xnor U2075 (N_2075,N_1896,In_1315);
and U2076 (N_2076,N_1980,N_1019);
and U2077 (N_2077,N_1510,N_1908);
or U2078 (N_2078,N_716,N_1965);
nand U2079 (N_2079,N_1425,N_1934);
nor U2080 (N_2080,N_1832,N_1428);
and U2081 (N_2081,N_1906,In_33);
xnor U2082 (N_2082,In_2783,N_1697);
xor U2083 (N_2083,In_772,N_732);
and U2084 (N_2084,N_1569,In_1151);
nand U2085 (N_2085,In_1526,N_1408);
and U2086 (N_2086,In_532,N_1605);
nor U2087 (N_2087,N_1235,N_725);
nor U2088 (N_2088,N_1952,In_2670);
nor U2089 (N_2089,N_1447,N_1736);
xor U2090 (N_2090,N_1897,In_1808);
nand U2091 (N_2091,N_1796,N_1144);
and U2092 (N_2092,N_1703,In_2186);
and U2093 (N_2093,N_1790,N_1743);
and U2094 (N_2094,N_1307,N_1846);
nand U2095 (N_2095,In_2718,N_1059);
nand U2096 (N_2096,N_1948,N_1867);
and U2097 (N_2097,N_1706,N_1818);
or U2098 (N_2098,N_1923,N_1951);
and U2099 (N_2099,N_1530,N_1995);
and U2100 (N_2100,In_536,N_583);
xnor U2101 (N_2101,In_921,In_740);
nor U2102 (N_2102,N_1759,In_2825);
xor U2103 (N_2103,N_1611,In_2977);
or U2104 (N_2104,N_1620,N_1478);
nor U2105 (N_2105,N_1617,In_1745);
nand U2106 (N_2106,N_880,In_2600);
xor U2107 (N_2107,In_1288,In_2452);
and U2108 (N_2108,N_1811,N_1537);
or U2109 (N_2109,N_609,N_1457);
xnor U2110 (N_2110,In_588,N_1039);
or U2111 (N_2111,N_1935,N_1258);
nor U2112 (N_2112,N_1970,N_1483);
nor U2113 (N_2113,N_898,N_324);
nand U2114 (N_2114,N_1413,N_701);
xnor U2115 (N_2115,In_589,N_1730);
nor U2116 (N_2116,N_1963,N_879);
nand U2117 (N_2117,N_1833,N_1000);
nor U2118 (N_2118,N_915,N_1210);
and U2119 (N_2119,N_1880,N_1810);
or U2120 (N_2120,N_1536,In_1183);
and U2121 (N_2121,In_1840,In_38);
nand U2122 (N_2122,N_1807,N_1618);
nor U2123 (N_2123,N_15,N_1862);
xnor U2124 (N_2124,N_1476,N_1644);
xnor U2125 (N_2125,N_1974,N_785);
and U2126 (N_2126,N_1985,N_1992);
or U2127 (N_2127,In_2737,N_1879);
xnor U2128 (N_2128,N_1966,In_1890);
nor U2129 (N_2129,In_1164,N_1704);
and U2130 (N_2130,In_480,In_2719);
xor U2131 (N_2131,N_1648,N_981);
or U2132 (N_2132,N_1679,N_1119);
nor U2133 (N_2133,N_887,N_1836);
xor U2134 (N_2134,In_1438,N_560);
nor U2135 (N_2135,N_1979,N_1687);
nor U2136 (N_2136,N_1179,N_1261);
nor U2137 (N_2137,N_1945,In_2774);
nand U2138 (N_2138,N_1843,In_1130);
xnor U2139 (N_2139,N_1190,In_67);
nand U2140 (N_2140,N_1421,In_2644);
xor U2141 (N_2141,In_2922,N_1473);
or U2142 (N_2142,In_971,N_1216);
or U2143 (N_2143,N_1977,In_933);
xor U2144 (N_2144,N_1972,N_850);
xor U2145 (N_2145,In_1719,N_1298);
and U2146 (N_2146,N_485,N_1787);
or U2147 (N_2147,In_2184,In_736);
or U2148 (N_2148,In_1702,N_1863);
or U2149 (N_2149,N_1420,N_1924);
and U2150 (N_2150,In_2521,N_1919);
and U2151 (N_2151,N_1910,N_222);
xnor U2152 (N_2152,N_1253,In_1492);
and U2153 (N_2153,N_1640,N_1885);
xnor U2154 (N_2154,N_855,N_458);
nand U2155 (N_2155,In_2037,N_1958);
or U2156 (N_2156,In_2781,N_1589);
xnor U2157 (N_2157,N_1289,N_1886);
xnor U2158 (N_2158,N_1673,N_1849);
xor U2159 (N_2159,N_779,N_1048);
and U2160 (N_2160,N_1186,In_2379);
xor U2161 (N_2161,N_91,N_1793);
xnor U2162 (N_2162,N_1592,In_2988);
nor U2163 (N_2163,N_1323,In_1046);
and U2164 (N_2164,N_1837,N_1427);
and U2165 (N_2165,N_1858,N_1001);
or U2166 (N_2166,N_828,N_1034);
nand U2167 (N_2167,N_943,In_756);
nand U2168 (N_2168,N_1601,In_529);
nand U2169 (N_2169,N_1549,N_1499);
nand U2170 (N_2170,N_1356,In_1827);
or U2171 (N_2171,In_2483,In_1582);
or U2172 (N_2172,N_875,N_1815);
nand U2173 (N_2173,In_224,In_534);
and U2174 (N_2174,N_1922,N_1107);
nor U2175 (N_2175,In_2602,In_2024);
nand U2176 (N_2176,N_1642,In_796);
and U2177 (N_2177,N_175,In_145);
nand U2178 (N_2178,N_1692,N_764);
or U2179 (N_2179,N_1799,N_744);
and U2180 (N_2180,In_337,N_607);
nor U2181 (N_2181,N_1294,In_1728);
xor U2182 (N_2182,In_1175,In_2331);
nor U2183 (N_2183,N_1159,N_1768);
or U2184 (N_2184,In_2575,N_1763);
or U2185 (N_2185,N_1224,N_72);
and U2186 (N_2186,N_1519,N_1312);
and U2187 (N_2187,N_1716,N_1550);
xor U2188 (N_2188,In_2559,N_1839);
nor U2189 (N_2189,N_1149,N_1978);
or U2190 (N_2190,N_1883,N_1600);
or U2191 (N_2191,N_1655,N_1899);
or U2192 (N_2192,N_1627,N_1222);
and U2193 (N_2193,In_2442,N_1248);
nor U2194 (N_2194,N_461,In_214);
xor U2195 (N_2195,N_1812,N_1148);
xnor U2196 (N_2196,In_731,N_720);
nand U2197 (N_2197,N_1543,N_1973);
and U2198 (N_2198,N_1816,N_1848);
nand U2199 (N_2199,N_1399,N_1292);
or U2200 (N_2200,N_1525,N_1581);
xor U2201 (N_2201,N_2124,N_1650);
or U2202 (N_2202,N_2049,N_1971);
xnor U2203 (N_2203,In_2289,N_1636);
and U2204 (N_2204,N_1976,N_2047);
nand U2205 (N_2205,In_103,In_2661);
or U2206 (N_2206,N_824,N_2086);
and U2207 (N_2207,N_2158,N_2004);
nand U2208 (N_2208,N_279,N_2154);
or U2209 (N_2209,N_2073,N_2114);
or U2210 (N_2210,N_2189,In_1785);
and U2211 (N_2211,N_689,N_2061);
xnor U2212 (N_2212,N_1887,N_2092);
nor U2213 (N_2213,N_2011,N_1539);
nand U2214 (N_2214,In_1562,N_2025);
nand U2215 (N_2215,N_1440,N_2078);
xor U2216 (N_2216,In_2253,In_2947);
and U2217 (N_2217,N_2007,In_743);
or U2218 (N_2218,N_2082,N_1738);
nand U2219 (N_2219,N_1765,N_1578);
nand U2220 (N_2220,N_1702,N_1005);
nand U2221 (N_2221,N_1461,N_1595);
nand U2222 (N_2222,N_2109,N_1889);
xor U2223 (N_2223,In_1741,N_752);
and U2224 (N_2224,N_252,N_2036);
xor U2225 (N_2225,N_2127,N_2182);
or U2226 (N_2226,N_2012,N_2044);
nand U2227 (N_2227,In_2808,N_1558);
or U2228 (N_2228,In_1888,In_926);
or U2229 (N_2229,N_2066,N_1989);
nor U2230 (N_2230,N_2077,N_1804);
nand U2231 (N_2231,N_1441,N_1388);
or U2232 (N_2232,In_2623,N_2001);
and U2233 (N_2233,N_1941,In_2822);
or U2234 (N_2234,N_1606,N_1517);
nand U2235 (N_2235,In_66,N_1246);
or U2236 (N_2236,N_1993,In_2727);
xor U2237 (N_2237,N_1551,N_1751);
nand U2238 (N_2238,N_833,N_1126);
xor U2239 (N_2239,N_1920,N_1625);
nand U2240 (N_2240,N_1734,N_1160);
or U2241 (N_2241,N_1814,N_2172);
and U2242 (N_2242,N_2088,N_2144);
xnor U2243 (N_2243,N_2196,N_1490);
xor U2244 (N_2244,N_1726,N_2023);
or U2245 (N_2245,In_330,N_1434);
nor U2246 (N_2246,In_2923,N_1895);
xor U2247 (N_2247,N_1390,N_2186);
and U2248 (N_2248,N_1260,N_2131);
and U2249 (N_2249,N_1631,N_2098);
or U2250 (N_2250,N_1628,In_2971);
nand U2251 (N_2251,N_2119,N_2106);
xnor U2252 (N_2252,N_1693,N_2176);
and U2253 (N_2253,N_1405,N_1360);
and U2254 (N_2254,N_246,In_1755);
or U2255 (N_2255,In_349,N_1984);
nor U2256 (N_2256,N_1999,N_1346);
and U2257 (N_2257,In_1401,N_553);
or U2258 (N_2258,N_2142,N_1594);
nand U2259 (N_2259,N_1956,N_1134);
and U2260 (N_2260,N_1728,N_2087);
or U2261 (N_2261,N_1711,N_1826);
and U2262 (N_2262,N_2169,In_2213);
and U2263 (N_2263,N_1682,N_2165);
nand U2264 (N_2264,N_1902,N_1866);
xnor U2265 (N_2265,N_733,N_1133);
xor U2266 (N_2266,N_2051,N_1982);
nor U2267 (N_2267,N_1347,N_2108);
and U2268 (N_2268,N_1656,N_2035);
nor U2269 (N_2269,N_1967,In_107);
or U2270 (N_2270,N_2015,N_1285);
nand U2271 (N_2271,N_1855,N_1852);
nor U2272 (N_2272,N_466,N_1842);
nor U2273 (N_2273,In_2408,In_2867);
or U2274 (N_2274,N_1309,N_301);
or U2275 (N_2275,N_2069,N_2139);
nand U2276 (N_2276,N_1928,N_2122);
nor U2277 (N_2277,In_685,In_1692);
and U2278 (N_2278,N_2134,N_2020);
or U2279 (N_2279,N_2096,N_2132);
or U2280 (N_2280,In_2179,In_2486);
and U2281 (N_2281,In_472,N_2046);
nor U2282 (N_2282,N_1672,N_1521);
nand U2283 (N_2283,N_2058,N_1875);
or U2284 (N_2284,In_216,N_1332);
xor U2285 (N_2285,N_2042,N_2079);
nand U2286 (N_2286,N_603,In_2009);
nand U2287 (N_2287,In_159,N_2010);
and U2288 (N_2288,N_1472,N_249);
nand U2289 (N_2289,N_202,N_1914);
and U2290 (N_2290,N_1591,N_1456);
and U2291 (N_2291,In_1538,N_1533);
and U2292 (N_2292,N_1220,N_1056);
and U2293 (N_2293,N_1615,N_2095);
nor U2294 (N_2294,N_1996,N_1844);
or U2295 (N_2295,In_244,N_126);
nand U2296 (N_2296,N_2168,N_1556);
nand U2297 (N_2297,N_2018,In_1445);
and U2298 (N_2298,N_1659,N_754);
nor U2299 (N_2299,N_2040,N_1174);
or U2300 (N_2300,N_2171,N_1541);
nand U2301 (N_2301,N_2183,In_1942);
nor U2302 (N_2302,N_1247,N_2125);
nand U2303 (N_2303,N_1819,N_812);
and U2304 (N_2304,N_2068,N_2166);
or U2305 (N_2305,N_1712,In_2112);
xnor U2306 (N_2306,In_1801,N_1822);
nand U2307 (N_2307,N_1916,N_1869);
or U2308 (N_2308,In_1059,N_2126);
nand U2309 (N_2309,N_1429,N_2039);
nor U2310 (N_2310,N_1854,N_1008);
nor U2311 (N_2311,N_1870,N_1856);
nand U2312 (N_2312,In_293,N_1912);
xnor U2313 (N_2313,N_1385,N_677);
xnor U2314 (N_2314,N_1637,In_2904);
nor U2315 (N_2315,N_1755,In_2036);
xor U2316 (N_2316,N_2057,In_1181);
nand U2317 (N_2317,N_1981,In_24);
nor U2318 (N_2318,N_2157,In_165);
or U2319 (N_2319,In_2935,N_2041);
xnor U2320 (N_2320,In_1216,N_2145);
and U2321 (N_2321,N_2104,In_1784);
and U2322 (N_2322,N_1903,In_1157);
nor U2323 (N_2323,N_1909,N_2199);
xnor U2324 (N_2324,N_2033,In_134);
nor U2325 (N_2325,N_82,N_1779);
or U2326 (N_2326,N_1936,In_1852);
and U2327 (N_2327,N_1226,N_1322);
or U2328 (N_2328,N_2030,N_1432);
or U2329 (N_2329,N_1251,N_341);
nor U2330 (N_2330,N_2151,N_837);
or U2331 (N_2331,N_1663,In_2074);
or U2332 (N_2332,In_1228,N_2152);
xnor U2333 (N_2333,N_1853,N_160);
and U2334 (N_2334,N_2149,N_1122);
or U2335 (N_2335,N_205,N_1800);
and U2336 (N_2336,N_1596,N_2053);
xor U2337 (N_2337,N_2198,In_1023);
xor U2338 (N_2338,N_2136,N_2116);
or U2339 (N_2339,N_935,In_446);
and U2340 (N_2340,In_1283,N_2133);
nand U2341 (N_2341,In_2884,In_1314);
nand U2342 (N_2342,N_2091,N_1783);
or U2343 (N_2343,N_2050,N_2150);
nor U2344 (N_2344,N_100,N_2173);
nor U2345 (N_2345,In_16,N_1907);
nor U2346 (N_2346,N_1701,N_1376);
or U2347 (N_2347,N_2027,In_2202);
and U2348 (N_2348,N_1677,In_1694);
xnor U2349 (N_2349,In_1464,N_885);
xnor U2350 (N_2350,N_1053,In_1060);
xnor U2351 (N_2351,N_1291,N_1502);
nor U2352 (N_2352,In_2352,N_807);
xnor U2353 (N_2353,In_387,N_1214);
xor U2354 (N_2354,In_356,N_1245);
and U2355 (N_2355,N_1954,N_986);
or U2356 (N_2356,N_2019,In_2094);
xnor U2357 (N_2357,N_1166,N_2129);
nand U2358 (N_2358,N_283,N_1450);
or U2359 (N_2359,In_590,N_1198);
nand U2360 (N_2360,In_813,N_1725);
or U2361 (N_2361,N_1991,In_967);
nor U2362 (N_2362,N_2167,N_530);
and U2363 (N_2363,N_1609,N_1975);
nor U2364 (N_2364,N_2185,N_2175);
or U2365 (N_2365,N_1926,In_41);
nand U2366 (N_2366,N_1860,N_2090);
and U2367 (N_2367,N_2111,N_1515);
nor U2368 (N_2368,N_1162,N_1454);
or U2369 (N_2369,N_1942,N_1328);
xor U2370 (N_2370,In_25,N_2121);
nand U2371 (N_2371,In_2696,N_1861);
nor U2372 (N_2372,In_1541,N_2008);
and U2373 (N_2373,N_2177,N_1608);
or U2374 (N_2374,In_2312,N_1337);
or U2375 (N_2375,N_2178,N_1871);
xnor U2376 (N_2376,N_1047,In_1832);
or U2377 (N_2377,N_1505,N_32);
xor U2378 (N_2378,N_2187,N_2017);
xnor U2379 (N_2379,N_601,In_1125);
xnor U2380 (N_2380,N_112,N_1286);
nor U2381 (N_2381,N_1933,N_604);
or U2382 (N_2382,In_2637,N_1859);
nor U2383 (N_2383,In_2987,In_1393);
or U2384 (N_2384,N_2123,N_1632);
nor U2385 (N_2385,N_1950,N_1099);
or U2386 (N_2386,In_2128,N_1324);
and U2387 (N_2387,N_1797,In_2146);
xnor U2388 (N_2388,In_2498,N_1946);
and U2389 (N_2389,N_1026,N_2034);
xor U2390 (N_2390,In_1462,N_2055);
xor U2391 (N_2391,In_1326,N_1338);
and U2392 (N_2392,N_1370,N_388);
and U2393 (N_2393,N_1735,In_426);
or U2394 (N_2394,In_2931,In_2643);
and U2395 (N_2395,In_1071,In_619);
nor U2396 (N_2396,In_1049,N_2024);
xor U2397 (N_2397,N_1786,N_1921);
or U2398 (N_2398,N_1888,In_1709);
nand U2399 (N_2399,N_2014,In_1964);
nand U2400 (N_2400,N_1172,N_2296);
nand U2401 (N_2401,N_1901,In_2046);
nor U2402 (N_2402,N_2056,In_1751);
xor U2403 (N_2403,N_2037,In_1355);
and U2404 (N_2404,N_2278,N_2288);
xor U2405 (N_2405,N_2045,N_2305);
nor U2406 (N_2406,N_2210,N_1691);
and U2407 (N_2407,N_2355,In_362);
nand U2408 (N_2408,N_989,N_2323);
nand U2409 (N_2409,N_1749,N_1997);
or U2410 (N_2410,N_2222,N_2118);
nor U2411 (N_2411,N_2099,N_438);
and U2412 (N_2412,N_2249,N_2128);
xor U2413 (N_2413,In_368,N_2333);
nand U2414 (N_2414,N_1904,N_978);
or U2415 (N_2415,N_2080,In_1663);
xor U2416 (N_2416,In_2380,N_2382);
and U2417 (N_2417,In_2659,N_567);
xnor U2418 (N_2418,In_729,N_2141);
or U2419 (N_2419,In_45,N_2159);
and U2420 (N_2420,N_1929,N_2256);
xor U2421 (N_2421,In_1686,N_1406);
nor U2422 (N_2422,N_2270,In_256);
or U2423 (N_2423,N_2021,N_848);
and U2424 (N_2424,N_2240,N_1748);
and U2425 (N_2425,N_2283,N_2335);
or U2426 (N_2426,In_396,In_201);
or U2427 (N_2427,N_2359,N_1092);
xor U2428 (N_2428,N_871,In_2850);
or U2429 (N_2429,In_1619,N_1960);
xor U2430 (N_2430,N_1761,N_2075);
nor U2431 (N_2431,N_2138,N_2251);
and U2432 (N_2432,N_2137,N_373);
nand U2433 (N_2433,N_1284,N_2101);
xnor U2434 (N_2434,N_2298,N_2361);
and U2435 (N_2435,N_1340,N_1825);
and U2436 (N_2436,In_478,N_1705);
or U2437 (N_2437,N_2234,N_1939);
nand U2438 (N_2438,N_2238,N_2052);
nor U2439 (N_2439,N_2380,N_2362);
and U2440 (N_2440,In_648,N_1709);
and U2441 (N_2441,N_2192,N_178);
nand U2442 (N_2442,N_2016,N_2373);
and U2443 (N_2443,N_2148,N_2225);
nor U2444 (N_2444,N_2337,N_1944);
nand U2445 (N_2445,N_1876,N_2054);
xnor U2446 (N_2446,N_2232,N_1614);
xor U2447 (N_2447,N_566,N_2247);
xor U2448 (N_2448,N_2365,N_2162);
nor U2449 (N_2449,N_1715,N_2241);
nand U2450 (N_2450,N_2297,N_825);
and U2451 (N_2451,N_2327,N_815);
nor U2452 (N_2452,In_527,N_1817);
and U2453 (N_2453,N_19,N_2262);
nor U2454 (N_2454,N_1877,N_2221);
or U2455 (N_2455,In_428,N_1676);
nand U2456 (N_2456,N_2102,N_2164);
xor U2457 (N_2457,N_1431,N_1685);
nor U2458 (N_2458,N_2065,N_48);
nor U2459 (N_2459,N_2006,N_2397);
or U2460 (N_2460,N_1894,N_2315);
nor U2461 (N_2461,N_2339,N_1808);
xor U2462 (N_2462,N_1125,N_1838);
and U2463 (N_2463,N_2100,N_1392);
and U2464 (N_2464,N_230,N_2377);
nand U2465 (N_2465,N_2135,N_1872);
nor U2466 (N_2466,In_2713,N_1714);
or U2467 (N_2467,N_2261,N_2084);
nor U2468 (N_2468,N_2120,N_1881);
xor U2469 (N_2469,In_960,N_2002);
or U2470 (N_2470,N_2268,In_164);
nor U2471 (N_2471,N_1158,N_2153);
nand U2472 (N_2472,N_2230,N_644);
or U2473 (N_2473,N_1947,N_84);
and U2474 (N_2474,N_965,N_2043);
and U2475 (N_2475,N_1362,N_2081);
nand U2476 (N_2476,N_2322,N_1040);
and U2477 (N_2477,N_2223,In_2031);
or U2478 (N_2478,N_1599,In_1204);
xnor U2479 (N_2479,In_615,N_188);
nand U2480 (N_2480,N_372,N_2358);
nand U2481 (N_2481,N_2388,N_2236);
or U2482 (N_2482,N_2293,N_1917);
nor U2483 (N_2483,N_2363,N_1828);
nor U2484 (N_2484,N_2312,In_1163);
nor U2485 (N_2485,N_2105,N_1986);
nand U2486 (N_2486,N_1025,N_1140);
or U2487 (N_2487,In_2272,N_26);
nand U2488 (N_2488,In_1275,N_1464);
xnor U2489 (N_2489,N_799,N_621);
xnor U2490 (N_2490,N_1718,In_1804);
and U2491 (N_2491,In_2490,N_2032);
and U2492 (N_2492,N_910,N_2212);
nor U2493 (N_2493,N_2174,N_1586);
xnor U2494 (N_2494,In_1240,N_1629);
xor U2495 (N_2495,In_1424,In_36);
nand U2496 (N_2496,N_1777,N_2094);
xor U2497 (N_2497,In_1186,In_1293);
and U2498 (N_2498,N_2214,N_123);
and U2499 (N_2499,N_1840,N_1968);
xor U2500 (N_2500,N_2385,N_2246);
xor U2501 (N_2501,N_2194,N_2267);
nor U2502 (N_2502,N_1402,In_2715);
xor U2503 (N_2503,N_2253,N_2258);
nand U2504 (N_2504,N_1027,N_2328);
or U2505 (N_2505,N_2394,N_1813);
or U2506 (N_2506,N_2300,N_1957);
and U2507 (N_2507,N_831,N_2083);
nor U2508 (N_2508,N_836,N_2181);
nand U2509 (N_2509,N_2217,N_1962);
and U2510 (N_2510,N_2260,N_1802);
and U2511 (N_2511,In_2220,N_2204);
nor U2512 (N_2512,N_2378,In_707);
nor U2513 (N_2513,N_2391,N_281);
nand U2514 (N_2514,In_2157,N_2013);
nor U2515 (N_2515,N_1891,In_701);
nand U2516 (N_2516,N_911,N_1448);
and U2517 (N_2517,In_623,N_2218);
or U2518 (N_2518,N_2302,N_2294);
or U2519 (N_2519,N_1953,In_1843);
nor U2520 (N_2520,N_1878,N_1874);
and U2521 (N_2521,N_2250,N_1857);
and U2522 (N_2522,N_1363,N_2389);
nor U2523 (N_2523,In_1079,N_1023);
or U2524 (N_2524,N_1616,N_1760);
nand U2525 (N_2525,N_2399,N_2067);
nand U2526 (N_2526,N_2303,N_2254);
nor U2527 (N_2527,N_1742,N_1821);
or U2528 (N_2528,N_532,N_2320);
and U2529 (N_2529,In_2087,N_2321);
nand U2530 (N_2530,In_2601,In_2182);
nand U2531 (N_2531,N_1829,N_409);
or U2532 (N_2532,N_1400,N_1809);
and U2533 (N_2533,In_2658,N_2226);
or U2534 (N_2534,N_2026,N_2332);
xor U2535 (N_2535,N_1949,In_484);
or U2536 (N_2536,N_2271,N_2370);
xor U2537 (N_2537,N_2304,N_2205);
nor U2538 (N_2538,N_121,N_905);
nor U2539 (N_2539,N_2356,N_1754);
nor U2540 (N_2540,N_2282,N_1547);
nand U2541 (N_2541,N_2264,N_2191);
xnor U2542 (N_2542,N_1295,N_1764);
xor U2543 (N_2543,N_2009,N_2203);
nand U2544 (N_2544,N_1955,N_1526);
nand U2545 (N_2545,N_2330,N_1983);
or U2546 (N_2546,N_1369,N_1623);
xor U2547 (N_2547,In_715,N_1987);
nor U2548 (N_2548,In_1236,N_1731);
and U2549 (N_2549,N_618,In_1328);
xor U2550 (N_2550,In_622,N_2273);
nor U2551 (N_2551,N_2274,N_2000);
or U2552 (N_2552,In_2706,N_2255);
and U2553 (N_2553,N_2383,N_2368);
nor U2554 (N_2554,N_2112,N_1798);
xor U2555 (N_2555,N_1554,N_2197);
xor U2556 (N_2556,N_597,N_515);
and U2557 (N_2557,N_511,N_2350);
and U2558 (N_2558,N_780,N_1375);
nand U2559 (N_2559,N_492,N_2390);
nand U2560 (N_2560,N_1915,N_2289);
nand U2561 (N_2561,In_1989,N_2060);
nor U2562 (N_2562,N_1882,N_2063);
and U2563 (N_2563,N_2295,N_521);
nand U2564 (N_2564,N_1664,In_1558);
xor U2565 (N_2565,N_2245,N_2367);
nor U2566 (N_2566,N_894,N_2265);
nand U2567 (N_2567,N_1898,N_2224);
or U2568 (N_2568,N_2375,In_644);
nand U2569 (N_2569,N_2089,N_2220);
xor U2570 (N_2570,N_2311,N_2338);
and U2571 (N_2571,N_2071,In_1670);
and U2572 (N_2572,N_1841,N_1641);
xnor U2573 (N_2573,N_2343,N_2201);
or U2574 (N_2574,N_2190,In_2679);
and U2575 (N_2575,N_1943,N_1383);
nand U2576 (N_2576,N_2319,N_2028);
or U2577 (N_2577,N_1795,In_1015);
nand U2578 (N_2578,N_2349,In_1830);
xor U2579 (N_2579,N_2147,N_734);
or U2580 (N_2580,N_2263,N_2364);
or U2581 (N_2581,N_1575,N_1386);
nor U2582 (N_2582,N_2398,N_1834);
and U2583 (N_2583,In_1363,N_1905);
and U2584 (N_2584,In_1905,N_228);
or U2585 (N_2585,N_1988,N_1666);
xnor U2586 (N_2586,In_819,N_2279);
nor U2587 (N_2587,N_1436,N_2243);
or U2588 (N_2588,N_2022,In_2944);
nor U2589 (N_2589,In_386,N_1806);
nor U2590 (N_2590,In_2708,N_1801);
xor U2591 (N_2591,N_33,In_1897);
and U2592 (N_2592,N_2379,N_498);
and U2593 (N_2593,N_2345,N_2062);
nor U2594 (N_2594,N_2003,N_2317);
nor U2595 (N_2595,N_1433,N_2366);
or U2596 (N_2596,N_1927,In_881);
xor U2597 (N_2597,N_1108,N_2202);
and U2598 (N_2598,N_471,N_1937);
nand U2599 (N_2599,N_2252,N_2146);
xor U2600 (N_2600,N_2286,N_541);
nand U2601 (N_2601,N_2156,N_2376);
nor U2602 (N_2602,N_2421,N_2170);
xnor U2603 (N_2603,N_2309,N_2576);
xnor U2604 (N_2604,N_358,N_2509);
and U2605 (N_2605,N_2525,N_2405);
xnor U2606 (N_2606,N_2413,N_2275);
xnor U2607 (N_2607,N_2228,N_2541);
or U2608 (N_2608,N_2188,In_2077);
nor U2609 (N_2609,N_2369,N_2479);
xor U2610 (N_2610,N_2248,N_2481);
xor U2611 (N_2611,N_1745,N_2299);
nor U2612 (N_2612,N_1823,N_2209);
and U2613 (N_2613,N_2482,N_2291);
or U2614 (N_2614,N_2466,N_2408);
nor U2615 (N_2615,N_1964,N_2582);
nor U2616 (N_2616,N_2528,N_2184);
or U2617 (N_2617,N_2453,N_2573);
and U2618 (N_2618,N_2517,N_2235);
nor U2619 (N_2619,In_2871,N_2591);
nor U2620 (N_2620,N_2231,N_2499);
nand U2621 (N_2621,N_2371,N_2588);
nand U2622 (N_2622,N_2495,N_2284);
nand U2623 (N_2623,N_2431,N_2005);
and U2624 (N_2624,N_2396,N_2522);
or U2625 (N_2625,N_2354,N_2539);
nand U2626 (N_2626,N_2425,N_2386);
or U2627 (N_2627,N_1803,N_1649);
nor U2628 (N_2628,N_2324,N_2443);
nor U2629 (N_2629,N_2352,N_2244);
nand U2630 (N_2630,N_2587,N_2507);
or U2631 (N_2631,In_422,N_2513);
nand U2632 (N_2632,N_2473,N_1389);
and U2633 (N_2633,N_2546,N_2113);
and U2634 (N_2634,N_1820,N_1865);
nor U2635 (N_2635,N_2393,N_2579);
or U2636 (N_2636,N_2574,N_2277);
xnor U2637 (N_2637,N_2511,N_2492);
xnor U2638 (N_2638,N_2475,N_661);
xnor U2639 (N_2639,N_2357,N_1255);
xnor U2640 (N_2640,N_330,N_1930);
nor U2641 (N_2641,N_2523,N_2329);
and U2642 (N_2642,In_1324,N_2557);
or U2643 (N_2643,N_2360,N_1404);
and U2644 (N_2644,N_2480,N_2444);
and U2645 (N_2645,N_2331,N_2072);
xor U2646 (N_2646,N_1746,N_2059);
xnor U2647 (N_2647,N_2410,N_2287);
and U2648 (N_2648,N_2516,N_1568);
nand U2649 (N_2649,N_2494,N_2430);
and U2650 (N_2650,N_2401,N_2478);
xor U2651 (N_2651,N_2407,N_2403);
nand U2652 (N_2652,N_2458,N_2441);
nor U2653 (N_2653,N_2461,N_2237);
nand U2654 (N_2654,N_2306,N_2486);
nand U2655 (N_2655,N_2347,N_2455);
xor U2656 (N_2656,N_2281,N_2521);
or U2657 (N_2657,N_1752,N_2435);
nand U2658 (N_2658,N_2308,N_2313);
or U2659 (N_2659,N_2484,N_735);
nand U2660 (N_2660,N_2566,N_921);
nand U2661 (N_2661,N_1481,N_2501);
nor U2662 (N_2662,N_2526,N_2213);
nand U2663 (N_2663,N_2549,N_2448);
nor U2664 (N_2664,N_2457,N_2437);
nand U2665 (N_2665,N_2334,N_2316);
xor U2666 (N_2666,N_2551,N_2552);
nor U2667 (N_2667,N_2599,N_2163);
nand U2668 (N_2668,N_2556,N_997);
and U2669 (N_2669,N_2233,N_2227);
and U2670 (N_2670,N_2527,N_2524);
or U2671 (N_2671,N_2342,N_2533);
nor U2672 (N_2672,N_2180,N_2581);
xor U2673 (N_2673,N_2414,N_2519);
or U2674 (N_2674,N_715,N_2586);
and U2675 (N_2675,N_2325,N_2107);
or U2676 (N_2676,N_2422,N_2514);
nand U2677 (N_2677,N_2280,N_2465);
and U2678 (N_2678,N_2314,N_2143);
or U2679 (N_2679,N_2489,N_163);
xor U2680 (N_2680,N_2029,N_2535);
and U2681 (N_2681,In_2595,N_2485);
xor U2682 (N_2682,N_2269,N_2442);
and U2683 (N_2683,N_2471,N_2491);
nor U2684 (N_2684,N_2292,N_2406);
and U2685 (N_2685,N_2215,N_2257);
nand U2686 (N_2686,N_2307,N_2451);
nand U2687 (N_2687,N_2518,N_2577);
and U2688 (N_2688,N_1913,N_1495);
and U2689 (N_2689,N_2548,N_2545);
or U2690 (N_2690,N_2450,N_2229);
and U2691 (N_2691,N_2565,N_2423);
nand U2692 (N_2692,N_2348,N_2572);
and U2693 (N_2693,N_2583,N_2438);
nand U2694 (N_2694,N_2340,N_588);
or U2695 (N_2695,In_1486,N_2070);
nor U2696 (N_2696,N_2567,N_2449);
or U2697 (N_2697,N_2460,N_2140);
nand U2698 (N_2698,N_728,N_2310);
or U2699 (N_2699,N_2477,N_2117);
and U2700 (N_2700,N_2476,N_2464);
and U2701 (N_2701,N_2496,N_2554);
or U2702 (N_2702,N_1931,In_1342);
and U2703 (N_2703,N_2470,N_2239);
xor U2704 (N_2704,N_2543,N_2031);
and U2705 (N_2705,N_2372,N_25);
or U2706 (N_2706,N_2596,N_2439);
nor U2707 (N_2707,N_2540,N_2504);
and U2708 (N_2708,N_2276,N_2207);
nand U2709 (N_2709,N_2416,N_401);
xnor U2710 (N_2710,N_2538,N_2336);
xor U2711 (N_2711,N_2502,N_2193);
nor U2712 (N_2712,In_2539,N_2130);
or U2713 (N_2713,N_2555,N_2436);
nor U2714 (N_2714,N_2593,N_2301);
and U2715 (N_2715,In_1128,N_2427);
nand U2716 (N_2716,N_2590,N_2468);
nor U2717 (N_2717,N_2510,N_2488);
or U2718 (N_2718,In_1940,N_2459);
or U2719 (N_2719,N_2505,N_1890);
or U2720 (N_2720,N_2542,N_2472);
nor U2721 (N_2721,N_2578,N_2076);
and U2722 (N_2722,N_2318,N_2415);
xor U2723 (N_2723,N_2490,N_1103);
or U2724 (N_2724,N_2103,N_412);
xnor U2725 (N_2725,N_2160,N_1698);
nor U2726 (N_2726,N_1824,N_2463);
nor U2727 (N_2727,N_2483,N_2387);
nand U2728 (N_2728,N_2456,N_2446);
and U2729 (N_2729,N_1397,N_2417);
nand U2730 (N_2730,N_2447,N_262);
nor U2731 (N_2731,N_2585,In_1119);
or U2732 (N_2732,N_2272,N_455);
or U2733 (N_2733,N_2412,N_765);
or U2734 (N_2734,N_2155,N_2537);
xnor U2735 (N_2735,N_2553,N_1274);
or U2736 (N_2736,N_1603,N_2558);
xor U2737 (N_2737,N_2474,N_2402);
nand U2738 (N_2738,N_2381,N_2211);
or U2739 (N_2739,N_2048,N_519);
and U2740 (N_2740,N_1455,N_2512);
and U2741 (N_2741,N_2570,N_2400);
nand U2742 (N_2742,N_2419,N_1268);
or U2743 (N_2743,N_2200,N_2085);
nand U2744 (N_2744,N_2550,N_1710);
nand U2745 (N_2745,N_2429,N_2497);
xnor U2746 (N_2746,N_1084,N_1645);
nand U2747 (N_2747,N_2426,N_1940);
or U2748 (N_2748,N_2575,N_2208);
or U2749 (N_2749,N_2392,N_2219);
and U2750 (N_2750,N_1621,N_2597);
nor U2751 (N_2751,N_2487,N_2341);
nand U2752 (N_2752,N_2536,N_2409);
xor U2753 (N_2753,N_1489,N_215);
nand U2754 (N_2754,N_2568,N_2216);
or U2755 (N_2755,N_2285,N_1830);
or U2756 (N_2756,N_2351,N_2547);
nand U2757 (N_2757,N_2266,N_2206);
and U2758 (N_2758,N_2580,N_2592);
and U2759 (N_2759,N_2038,N_1847);
or U2760 (N_2760,N_1267,N_1555);
and U2761 (N_2761,N_2498,In_383);
xor U2762 (N_2762,N_2395,N_2161);
nor U2763 (N_2763,N_2434,In_2276);
nor U2764 (N_2764,N_2326,N_2290);
nor U2765 (N_2765,N_2493,N_2562);
nand U2766 (N_2766,N_2561,N_2259);
and U2767 (N_2767,N_2420,N_2559);
xnor U2768 (N_2768,N_2598,In_727);
xnor U2769 (N_2769,N_2462,N_2531);
nand U2770 (N_2770,N_2508,N_2584);
nand U2771 (N_2771,N_1845,N_2534);
nor U2772 (N_2772,N_2411,In_359);
nor U2773 (N_2773,N_2195,N_2500);
and U2774 (N_2774,N_2344,N_2532);
nand U2775 (N_2775,N_2428,N_2544);
nor U2776 (N_2776,N_2353,N_2074);
or U2777 (N_2777,N_2520,N_2515);
or U2778 (N_2778,N_1660,N_2424);
nand U2779 (N_2779,In_1699,N_1587);
xor U2780 (N_2780,N_2384,N_2560);
nand U2781 (N_2781,N_2569,N_2440);
xor U2782 (N_2782,In_1056,N_2346);
and U2783 (N_2783,N_2452,N_2445);
or U2784 (N_2784,N_2564,N_2097);
xor U2785 (N_2785,N_2467,N_2110);
xnor U2786 (N_2786,N_2469,N_2179);
nor U2787 (N_2787,N_2589,N_2093);
nor U2788 (N_2788,N_1961,N_2506);
or U2789 (N_2789,N_2503,In_2523);
xor U2790 (N_2790,N_2529,N_1835);
or U2791 (N_2791,N_1520,N_2064);
or U2792 (N_2792,N_913,N_2571);
nor U2793 (N_2793,N_2433,In_1212);
xor U2794 (N_2794,N_2242,N_1959);
nor U2795 (N_2795,N_2432,N_2454);
and U2796 (N_2796,N_2594,N_2595);
and U2797 (N_2797,N_2374,N_2115);
nor U2798 (N_2798,N_2530,N_2563);
and U2799 (N_2799,N_2418,N_2404);
or U2800 (N_2800,N_2770,N_2644);
and U2801 (N_2801,N_2682,N_2754);
nand U2802 (N_2802,N_2703,N_2793);
nand U2803 (N_2803,N_2642,N_2621);
nand U2804 (N_2804,N_2677,N_2675);
and U2805 (N_2805,N_2661,N_2766);
nor U2806 (N_2806,N_2776,N_2716);
xor U2807 (N_2807,N_2710,N_2745);
and U2808 (N_2808,N_2764,N_2616);
xnor U2809 (N_2809,N_2797,N_2707);
nand U2810 (N_2810,N_2704,N_2714);
or U2811 (N_2811,N_2645,N_2700);
and U2812 (N_2812,N_2639,N_2780);
nand U2813 (N_2813,N_2692,N_2749);
or U2814 (N_2814,N_2751,N_2606);
xnor U2815 (N_2815,N_2648,N_2734);
nor U2816 (N_2816,N_2673,N_2631);
nor U2817 (N_2817,N_2667,N_2744);
nand U2818 (N_2818,N_2740,N_2701);
nor U2819 (N_2819,N_2638,N_2759);
and U2820 (N_2820,N_2633,N_2671);
nor U2821 (N_2821,N_2722,N_2656);
or U2822 (N_2822,N_2623,N_2630);
xnor U2823 (N_2823,N_2691,N_2628);
nand U2824 (N_2824,N_2627,N_2695);
or U2825 (N_2825,N_2654,N_2634);
xnor U2826 (N_2826,N_2679,N_2785);
nand U2827 (N_2827,N_2624,N_2796);
nor U2828 (N_2828,N_2635,N_2782);
and U2829 (N_2829,N_2659,N_2750);
and U2830 (N_2830,N_2611,N_2657);
nand U2831 (N_2831,N_2632,N_2713);
and U2832 (N_2832,N_2746,N_2727);
and U2833 (N_2833,N_2613,N_2698);
nor U2834 (N_2834,N_2612,N_2795);
nor U2835 (N_2835,N_2672,N_2741);
and U2836 (N_2836,N_2725,N_2689);
or U2837 (N_2837,N_2696,N_2721);
nand U2838 (N_2838,N_2778,N_2752);
nor U2839 (N_2839,N_2678,N_2605);
xor U2840 (N_2840,N_2607,N_2724);
xor U2841 (N_2841,N_2777,N_2761);
and U2842 (N_2842,N_2735,N_2603);
nand U2843 (N_2843,N_2636,N_2646);
nor U2844 (N_2844,N_2769,N_2739);
nor U2845 (N_2845,N_2781,N_2748);
and U2846 (N_2846,N_2681,N_2653);
or U2847 (N_2847,N_2762,N_2765);
or U2848 (N_2848,N_2602,N_2690);
nor U2849 (N_2849,N_2755,N_2614);
and U2850 (N_2850,N_2650,N_2753);
nand U2851 (N_2851,N_2711,N_2660);
or U2852 (N_2852,N_2670,N_2720);
nor U2853 (N_2853,N_2786,N_2723);
nand U2854 (N_2854,N_2699,N_2600);
xnor U2855 (N_2855,N_2747,N_2784);
or U2856 (N_2856,N_2729,N_2774);
nor U2857 (N_2857,N_2773,N_2733);
or U2858 (N_2858,N_2680,N_2662);
and U2859 (N_2859,N_2772,N_2788);
xnor U2860 (N_2860,N_2718,N_2676);
nor U2861 (N_2861,N_2697,N_2640);
and U2862 (N_2862,N_2643,N_2685);
xor U2863 (N_2863,N_2687,N_2688);
nand U2864 (N_2864,N_2647,N_2663);
or U2865 (N_2865,N_2705,N_2649);
nand U2866 (N_2866,N_2775,N_2792);
or U2867 (N_2867,N_2736,N_2622);
xnor U2868 (N_2868,N_2789,N_2655);
xor U2869 (N_2869,N_2668,N_2669);
nand U2870 (N_2870,N_2763,N_2601);
or U2871 (N_2871,N_2768,N_2742);
nor U2872 (N_2872,N_2715,N_2706);
and U2873 (N_2873,N_2717,N_2779);
and U2874 (N_2874,N_2791,N_2767);
nor U2875 (N_2875,N_2625,N_2794);
xnor U2876 (N_2876,N_2608,N_2756);
xnor U2877 (N_2877,N_2629,N_2674);
and U2878 (N_2878,N_2731,N_2738);
and U2879 (N_2879,N_2760,N_2771);
and U2880 (N_2880,N_2743,N_2758);
nor U2881 (N_2881,N_2783,N_2641);
and U2882 (N_2882,N_2651,N_2709);
nand U2883 (N_2883,N_2637,N_2615);
or U2884 (N_2884,N_2652,N_2726);
nand U2885 (N_2885,N_2757,N_2684);
nor U2886 (N_2886,N_2693,N_2618);
and U2887 (N_2887,N_2658,N_2737);
nand U2888 (N_2888,N_2719,N_2610);
nor U2889 (N_2889,N_2617,N_2798);
xor U2890 (N_2890,N_2732,N_2626);
or U2891 (N_2891,N_2683,N_2664);
xnor U2892 (N_2892,N_2790,N_2619);
or U2893 (N_2893,N_2686,N_2604);
xnor U2894 (N_2894,N_2730,N_2799);
nor U2895 (N_2895,N_2787,N_2609);
and U2896 (N_2896,N_2665,N_2620);
and U2897 (N_2897,N_2702,N_2712);
xnor U2898 (N_2898,N_2728,N_2666);
xor U2899 (N_2899,N_2694,N_2708);
nand U2900 (N_2900,N_2667,N_2662);
xor U2901 (N_2901,N_2638,N_2688);
xnor U2902 (N_2902,N_2752,N_2763);
and U2903 (N_2903,N_2765,N_2791);
and U2904 (N_2904,N_2635,N_2642);
or U2905 (N_2905,N_2633,N_2606);
nand U2906 (N_2906,N_2738,N_2733);
nor U2907 (N_2907,N_2748,N_2632);
or U2908 (N_2908,N_2766,N_2616);
nor U2909 (N_2909,N_2761,N_2779);
nor U2910 (N_2910,N_2656,N_2640);
and U2911 (N_2911,N_2672,N_2627);
xnor U2912 (N_2912,N_2647,N_2705);
or U2913 (N_2913,N_2694,N_2636);
and U2914 (N_2914,N_2668,N_2650);
nand U2915 (N_2915,N_2618,N_2783);
or U2916 (N_2916,N_2783,N_2695);
nand U2917 (N_2917,N_2705,N_2675);
nor U2918 (N_2918,N_2627,N_2755);
and U2919 (N_2919,N_2778,N_2609);
xor U2920 (N_2920,N_2658,N_2734);
nand U2921 (N_2921,N_2718,N_2660);
xor U2922 (N_2922,N_2701,N_2652);
and U2923 (N_2923,N_2618,N_2704);
nand U2924 (N_2924,N_2650,N_2648);
xnor U2925 (N_2925,N_2728,N_2674);
and U2926 (N_2926,N_2706,N_2755);
or U2927 (N_2927,N_2788,N_2693);
and U2928 (N_2928,N_2719,N_2757);
or U2929 (N_2929,N_2739,N_2768);
nor U2930 (N_2930,N_2733,N_2741);
nand U2931 (N_2931,N_2721,N_2638);
and U2932 (N_2932,N_2668,N_2734);
and U2933 (N_2933,N_2793,N_2678);
nor U2934 (N_2934,N_2701,N_2771);
and U2935 (N_2935,N_2638,N_2790);
or U2936 (N_2936,N_2666,N_2730);
and U2937 (N_2937,N_2722,N_2688);
or U2938 (N_2938,N_2748,N_2759);
and U2939 (N_2939,N_2647,N_2765);
nand U2940 (N_2940,N_2650,N_2609);
nor U2941 (N_2941,N_2791,N_2774);
or U2942 (N_2942,N_2737,N_2776);
and U2943 (N_2943,N_2615,N_2776);
nor U2944 (N_2944,N_2670,N_2635);
and U2945 (N_2945,N_2702,N_2603);
xor U2946 (N_2946,N_2736,N_2649);
nor U2947 (N_2947,N_2780,N_2783);
nor U2948 (N_2948,N_2651,N_2653);
and U2949 (N_2949,N_2769,N_2705);
or U2950 (N_2950,N_2759,N_2689);
and U2951 (N_2951,N_2660,N_2689);
nor U2952 (N_2952,N_2613,N_2626);
xnor U2953 (N_2953,N_2779,N_2697);
nor U2954 (N_2954,N_2695,N_2628);
nor U2955 (N_2955,N_2724,N_2756);
and U2956 (N_2956,N_2681,N_2667);
or U2957 (N_2957,N_2728,N_2749);
nand U2958 (N_2958,N_2714,N_2769);
xnor U2959 (N_2959,N_2705,N_2657);
nand U2960 (N_2960,N_2714,N_2749);
nand U2961 (N_2961,N_2652,N_2662);
or U2962 (N_2962,N_2698,N_2623);
or U2963 (N_2963,N_2685,N_2648);
and U2964 (N_2964,N_2702,N_2642);
and U2965 (N_2965,N_2670,N_2626);
or U2966 (N_2966,N_2730,N_2739);
and U2967 (N_2967,N_2768,N_2717);
xor U2968 (N_2968,N_2789,N_2784);
xor U2969 (N_2969,N_2693,N_2611);
nand U2970 (N_2970,N_2712,N_2706);
and U2971 (N_2971,N_2677,N_2767);
xnor U2972 (N_2972,N_2630,N_2728);
xor U2973 (N_2973,N_2691,N_2614);
nor U2974 (N_2974,N_2681,N_2759);
nor U2975 (N_2975,N_2783,N_2609);
xor U2976 (N_2976,N_2654,N_2671);
and U2977 (N_2977,N_2716,N_2656);
xor U2978 (N_2978,N_2700,N_2774);
or U2979 (N_2979,N_2638,N_2797);
nand U2980 (N_2980,N_2718,N_2753);
nor U2981 (N_2981,N_2773,N_2746);
nand U2982 (N_2982,N_2614,N_2758);
nor U2983 (N_2983,N_2679,N_2740);
or U2984 (N_2984,N_2729,N_2607);
nand U2985 (N_2985,N_2707,N_2792);
nand U2986 (N_2986,N_2749,N_2779);
nand U2987 (N_2987,N_2795,N_2652);
and U2988 (N_2988,N_2684,N_2741);
or U2989 (N_2989,N_2671,N_2698);
nor U2990 (N_2990,N_2695,N_2608);
xnor U2991 (N_2991,N_2768,N_2689);
xor U2992 (N_2992,N_2703,N_2749);
xor U2993 (N_2993,N_2710,N_2726);
and U2994 (N_2994,N_2663,N_2619);
nor U2995 (N_2995,N_2774,N_2717);
xor U2996 (N_2996,N_2762,N_2712);
or U2997 (N_2997,N_2798,N_2721);
and U2998 (N_2998,N_2655,N_2751);
nor U2999 (N_2999,N_2738,N_2794);
and U3000 (N_3000,N_2974,N_2854);
and U3001 (N_3001,N_2818,N_2907);
nor U3002 (N_3002,N_2834,N_2819);
and U3003 (N_3003,N_2864,N_2979);
nor U3004 (N_3004,N_2845,N_2810);
or U3005 (N_3005,N_2876,N_2860);
xnor U3006 (N_3006,N_2978,N_2981);
nor U3007 (N_3007,N_2921,N_2964);
xor U3008 (N_3008,N_2856,N_2842);
and U3009 (N_3009,N_2820,N_2914);
or U3010 (N_3010,N_2934,N_2982);
or U3011 (N_3011,N_2906,N_2888);
or U3012 (N_3012,N_2983,N_2881);
nand U3013 (N_3013,N_2957,N_2858);
or U3014 (N_3014,N_2877,N_2919);
xnor U3015 (N_3015,N_2951,N_2892);
nand U3016 (N_3016,N_2929,N_2841);
nand U3017 (N_3017,N_2887,N_2867);
xnor U3018 (N_3018,N_2863,N_2931);
and U3019 (N_3019,N_2980,N_2923);
nor U3020 (N_3020,N_2804,N_2975);
or U3021 (N_3021,N_2910,N_2821);
and U3022 (N_3022,N_2893,N_2968);
nor U3023 (N_3023,N_2809,N_2840);
or U3024 (N_3024,N_2855,N_2806);
nor U3025 (N_3025,N_2868,N_2823);
or U3026 (N_3026,N_2882,N_2822);
and U3027 (N_3027,N_2850,N_2994);
or U3028 (N_3028,N_2926,N_2835);
nor U3029 (N_3029,N_2991,N_2947);
xor U3030 (N_3030,N_2862,N_2996);
nand U3031 (N_3031,N_2946,N_2967);
and U3032 (N_3032,N_2824,N_2948);
nand U3033 (N_3033,N_2938,N_2956);
nand U3034 (N_3034,N_2812,N_2857);
nor U3035 (N_3035,N_2993,N_2866);
and U3036 (N_3036,N_2879,N_2941);
or U3037 (N_3037,N_2932,N_2905);
xnor U3038 (N_3038,N_2885,N_2988);
nor U3039 (N_3039,N_2904,N_2992);
or U3040 (N_3040,N_2811,N_2922);
xnor U3041 (N_3041,N_2960,N_2918);
nand U3042 (N_3042,N_2933,N_2954);
nand U3043 (N_3043,N_2817,N_2848);
nor U3044 (N_3044,N_2970,N_2800);
nand U3045 (N_3045,N_2832,N_2838);
and U3046 (N_3046,N_2920,N_2872);
and U3047 (N_3047,N_2895,N_2958);
nor U3048 (N_3048,N_2807,N_2846);
nor U3049 (N_3049,N_2878,N_2942);
nor U3050 (N_3050,N_2903,N_2898);
or U3051 (N_3051,N_2935,N_2897);
nand U3052 (N_3052,N_2963,N_2915);
xor U3053 (N_3053,N_2959,N_2899);
or U3054 (N_3054,N_2976,N_2861);
and U3055 (N_3055,N_2802,N_2816);
nor U3056 (N_3056,N_2873,N_2977);
or U3057 (N_3057,N_2891,N_2869);
and U3058 (N_3058,N_2890,N_2844);
nand U3059 (N_3059,N_2894,N_2883);
or U3060 (N_3060,N_2962,N_2896);
and U3061 (N_3061,N_2971,N_2808);
xor U3062 (N_3062,N_2829,N_2870);
and U3063 (N_3063,N_2949,N_2943);
and U3064 (N_3064,N_2831,N_2825);
nand U3065 (N_3065,N_2999,N_2966);
xnor U3066 (N_3066,N_2853,N_2801);
and U3067 (N_3067,N_2851,N_2839);
nor U3068 (N_3068,N_2952,N_2928);
nand U3069 (N_3069,N_2880,N_2961);
nand U3070 (N_3070,N_2874,N_2987);
xor U3071 (N_3071,N_2813,N_2945);
nor U3072 (N_3072,N_2997,N_2847);
nand U3073 (N_3073,N_2969,N_2805);
or U3074 (N_3074,N_2911,N_2944);
and U3075 (N_3075,N_2927,N_2972);
and U3076 (N_3076,N_2955,N_2875);
or U3077 (N_3077,N_2830,N_2985);
and U3078 (N_3078,N_2900,N_2827);
or U3079 (N_3079,N_2953,N_2828);
and U3080 (N_3080,N_2930,N_2912);
nor U3081 (N_3081,N_2901,N_2836);
nor U3082 (N_3082,N_2995,N_2843);
xnor U3083 (N_3083,N_2998,N_2965);
and U3084 (N_3084,N_2950,N_2939);
nand U3085 (N_3085,N_2865,N_2917);
nor U3086 (N_3086,N_2913,N_2940);
xor U3087 (N_3087,N_2837,N_2871);
xor U3088 (N_3088,N_2826,N_2925);
nor U3089 (N_3089,N_2909,N_2936);
nand U3090 (N_3090,N_2886,N_2889);
and U3091 (N_3091,N_2815,N_2902);
xnor U3092 (N_3092,N_2908,N_2916);
or U3093 (N_3093,N_2924,N_2814);
nor U3094 (N_3094,N_2852,N_2973);
xor U3095 (N_3095,N_2990,N_2989);
or U3096 (N_3096,N_2984,N_2833);
and U3097 (N_3097,N_2937,N_2803);
or U3098 (N_3098,N_2859,N_2986);
and U3099 (N_3099,N_2884,N_2849);
xnor U3100 (N_3100,N_2856,N_2987);
or U3101 (N_3101,N_2986,N_2817);
nor U3102 (N_3102,N_2921,N_2986);
or U3103 (N_3103,N_2847,N_2876);
nor U3104 (N_3104,N_2910,N_2832);
or U3105 (N_3105,N_2942,N_2965);
nor U3106 (N_3106,N_2842,N_2991);
and U3107 (N_3107,N_2958,N_2981);
or U3108 (N_3108,N_2964,N_2947);
nor U3109 (N_3109,N_2824,N_2984);
or U3110 (N_3110,N_2830,N_2953);
and U3111 (N_3111,N_2821,N_2950);
or U3112 (N_3112,N_2819,N_2990);
or U3113 (N_3113,N_2812,N_2874);
xor U3114 (N_3114,N_2975,N_2935);
or U3115 (N_3115,N_2986,N_2953);
or U3116 (N_3116,N_2972,N_2879);
and U3117 (N_3117,N_2941,N_2839);
or U3118 (N_3118,N_2841,N_2871);
or U3119 (N_3119,N_2945,N_2994);
and U3120 (N_3120,N_2839,N_2890);
xor U3121 (N_3121,N_2803,N_2999);
and U3122 (N_3122,N_2869,N_2958);
or U3123 (N_3123,N_2938,N_2864);
and U3124 (N_3124,N_2837,N_2957);
xnor U3125 (N_3125,N_2994,N_2971);
nor U3126 (N_3126,N_2874,N_2864);
nor U3127 (N_3127,N_2816,N_2909);
xnor U3128 (N_3128,N_2929,N_2900);
xor U3129 (N_3129,N_2811,N_2940);
nand U3130 (N_3130,N_2867,N_2916);
nand U3131 (N_3131,N_2824,N_2972);
xnor U3132 (N_3132,N_2811,N_2858);
xor U3133 (N_3133,N_2842,N_2925);
nor U3134 (N_3134,N_2922,N_2931);
nor U3135 (N_3135,N_2968,N_2813);
nor U3136 (N_3136,N_2829,N_2982);
or U3137 (N_3137,N_2848,N_2847);
nor U3138 (N_3138,N_2959,N_2928);
nor U3139 (N_3139,N_2904,N_2807);
xnor U3140 (N_3140,N_2843,N_2888);
or U3141 (N_3141,N_2920,N_2830);
xor U3142 (N_3142,N_2850,N_2903);
or U3143 (N_3143,N_2881,N_2930);
nor U3144 (N_3144,N_2919,N_2856);
nand U3145 (N_3145,N_2812,N_2878);
xnor U3146 (N_3146,N_2929,N_2978);
or U3147 (N_3147,N_2875,N_2904);
and U3148 (N_3148,N_2858,N_2926);
or U3149 (N_3149,N_2939,N_2898);
nand U3150 (N_3150,N_2946,N_2830);
and U3151 (N_3151,N_2887,N_2874);
and U3152 (N_3152,N_2851,N_2880);
or U3153 (N_3153,N_2817,N_2948);
or U3154 (N_3154,N_2800,N_2864);
nor U3155 (N_3155,N_2931,N_2880);
xor U3156 (N_3156,N_2990,N_2800);
or U3157 (N_3157,N_2947,N_2888);
nand U3158 (N_3158,N_2849,N_2994);
xnor U3159 (N_3159,N_2848,N_2919);
xor U3160 (N_3160,N_2884,N_2870);
and U3161 (N_3161,N_2886,N_2815);
and U3162 (N_3162,N_2906,N_2953);
nor U3163 (N_3163,N_2896,N_2948);
nor U3164 (N_3164,N_2931,N_2912);
nor U3165 (N_3165,N_2949,N_2859);
nor U3166 (N_3166,N_2890,N_2903);
nor U3167 (N_3167,N_2884,N_2817);
and U3168 (N_3168,N_2885,N_2970);
nand U3169 (N_3169,N_2856,N_2833);
nor U3170 (N_3170,N_2952,N_2827);
xnor U3171 (N_3171,N_2982,N_2868);
nor U3172 (N_3172,N_2820,N_2989);
nor U3173 (N_3173,N_2876,N_2853);
and U3174 (N_3174,N_2831,N_2916);
xor U3175 (N_3175,N_2824,N_2961);
nand U3176 (N_3176,N_2900,N_2833);
xor U3177 (N_3177,N_2849,N_2996);
xnor U3178 (N_3178,N_2979,N_2824);
nor U3179 (N_3179,N_2828,N_2945);
or U3180 (N_3180,N_2918,N_2872);
xnor U3181 (N_3181,N_2972,N_2850);
xor U3182 (N_3182,N_2852,N_2860);
nor U3183 (N_3183,N_2807,N_2923);
xor U3184 (N_3184,N_2921,N_2888);
and U3185 (N_3185,N_2961,N_2994);
and U3186 (N_3186,N_2872,N_2879);
nor U3187 (N_3187,N_2967,N_2865);
and U3188 (N_3188,N_2962,N_2869);
nand U3189 (N_3189,N_2954,N_2923);
nand U3190 (N_3190,N_2935,N_2995);
xor U3191 (N_3191,N_2803,N_2969);
or U3192 (N_3192,N_2950,N_2812);
nand U3193 (N_3193,N_2939,N_2955);
and U3194 (N_3194,N_2830,N_2822);
xor U3195 (N_3195,N_2949,N_2865);
and U3196 (N_3196,N_2835,N_2854);
and U3197 (N_3197,N_2947,N_2913);
or U3198 (N_3198,N_2934,N_2946);
nand U3199 (N_3199,N_2908,N_2872);
xnor U3200 (N_3200,N_3109,N_3159);
xor U3201 (N_3201,N_3158,N_3069);
and U3202 (N_3202,N_3048,N_3111);
or U3203 (N_3203,N_3171,N_3139);
xnor U3204 (N_3204,N_3065,N_3188);
and U3205 (N_3205,N_3122,N_3006);
nor U3206 (N_3206,N_3191,N_3146);
and U3207 (N_3207,N_3059,N_3103);
nor U3208 (N_3208,N_3027,N_3075);
or U3209 (N_3209,N_3060,N_3101);
or U3210 (N_3210,N_3183,N_3050);
nor U3211 (N_3211,N_3072,N_3024);
or U3212 (N_3212,N_3012,N_3083);
or U3213 (N_3213,N_3091,N_3178);
or U3214 (N_3214,N_3010,N_3029);
and U3215 (N_3215,N_3097,N_3166);
nor U3216 (N_3216,N_3047,N_3123);
or U3217 (N_3217,N_3143,N_3156);
nand U3218 (N_3218,N_3023,N_3070);
xor U3219 (N_3219,N_3022,N_3161);
xor U3220 (N_3220,N_3062,N_3057);
nand U3221 (N_3221,N_3034,N_3112);
xnor U3222 (N_3222,N_3044,N_3189);
nor U3223 (N_3223,N_3100,N_3162);
nor U3224 (N_3224,N_3016,N_3169);
and U3225 (N_3225,N_3179,N_3013);
and U3226 (N_3226,N_3137,N_3011);
xor U3227 (N_3227,N_3092,N_3197);
and U3228 (N_3228,N_3088,N_3190);
xnor U3229 (N_3229,N_3019,N_3008);
or U3230 (N_3230,N_3114,N_3045);
and U3231 (N_3231,N_3110,N_3105);
or U3232 (N_3232,N_3160,N_3026);
and U3233 (N_3233,N_3094,N_3093);
and U3234 (N_3234,N_3030,N_3067);
nand U3235 (N_3235,N_3157,N_3198);
and U3236 (N_3236,N_3118,N_3149);
or U3237 (N_3237,N_3127,N_3079);
or U3238 (N_3238,N_3020,N_3177);
xor U3239 (N_3239,N_3056,N_3098);
nor U3240 (N_3240,N_3038,N_3120);
xnor U3241 (N_3241,N_3192,N_3163);
nand U3242 (N_3242,N_3164,N_3117);
or U3243 (N_3243,N_3170,N_3066);
nand U3244 (N_3244,N_3167,N_3108);
or U3245 (N_3245,N_3174,N_3064);
nor U3246 (N_3246,N_3185,N_3039);
or U3247 (N_3247,N_3193,N_3124);
nor U3248 (N_3248,N_3005,N_3172);
nor U3249 (N_3249,N_3129,N_3053);
xor U3250 (N_3250,N_3154,N_3089);
and U3251 (N_3251,N_3073,N_3141);
or U3252 (N_3252,N_3078,N_3002);
or U3253 (N_3253,N_3014,N_3199);
nor U3254 (N_3254,N_3025,N_3113);
and U3255 (N_3255,N_3090,N_3152);
and U3256 (N_3256,N_3085,N_3133);
xnor U3257 (N_3257,N_3042,N_3130);
xor U3258 (N_3258,N_3142,N_3074);
nand U3259 (N_3259,N_3186,N_3135);
and U3260 (N_3260,N_3028,N_3181);
nand U3261 (N_3261,N_3131,N_3021);
nand U3262 (N_3262,N_3061,N_3081);
or U3263 (N_3263,N_3176,N_3001);
xor U3264 (N_3264,N_3058,N_3151);
nor U3265 (N_3265,N_3033,N_3107);
nand U3266 (N_3266,N_3121,N_3036);
nor U3267 (N_3267,N_3063,N_3187);
and U3268 (N_3268,N_3049,N_3043);
or U3269 (N_3269,N_3068,N_3041);
nor U3270 (N_3270,N_3194,N_3046);
nor U3271 (N_3271,N_3148,N_3147);
xnor U3272 (N_3272,N_3104,N_3145);
or U3273 (N_3273,N_3035,N_3009);
nand U3274 (N_3274,N_3055,N_3150);
and U3275 (N_3275,N_3168,N_3040);
xor U3276 (N_3276,N_3018,N_3102);
xnor U3277 (N_3277,N_3125,N_3000);
or U3278 (N_3278,N_3165,N_3015);
and U3279 (N_3279,N_3132,N_3136);
and U3280 (N_3280,N_3106,N_3128);
nor U3281 (N_3281,N_3180,N_3080);
nor U3282 (N_3282,N_3003,N_3115);
or U3283 (N_3283,N_3138,N_3086);
nand U3284 (N_3284,N_3076,N_3017);
nand U3285 (N_3285,N_3134,N_3031);
xnor U3286 (N_3286,N_3140,N_3195);
nor U3287 (N_3287,N_3082,N_3095);
nand U3288 (N_3288,N_3037,N_3196);
nor U3289 (N_3289,N_3051,N_3077);
or U3290 (N_3290,N_3175,N_3032);
xnor U3291 (N_3291,N_3182,N_3007);
xor U3292 (N_3292,N_3099,N_3155);
or U3293 (N_3293,N_3004,N_3084);
and U3294 (N_3294,N_3184,N_3126);
and U3295 (N_3295,N_3096,N_3116);
and U3296 (N_3296,N_3119,N_3144);
xnor U3297 (N_3297,N_3153,N_3071);
and U3298 (N_3298,N_3052,N_3173);
nand U3299 (N_3299,N_3087,N_3054);
or U3300 (N_3300,N_3147,N_3064);
nor U3301 (N_3301,N_3175,N_3088);
nand U3302 (N_3302,N_3003,N_3016);
nand U3303 (N_3303,N_3051,N_3026);
xnor U3304 (N_3304,N_3012,N_3073);
and U3305 (N_3305,N_3017,N_3014);
or U3306 (N_3306,N_3167,N_3144);
or U3307 (N_3307,N_3092,N_3105);
and U3308 (N_3308,N_3136,N_3104);
and U3309 (N_3309,N_3127,N_3169);
and U3310 (N_3310,N_3054,N_3187);
nand U3311 (N_3311,N_3181,N_3151);
nand U3312 (N_3312,N_3091,N_3089);
and U3313 (N_3313,N_3102,N_3152);
xnor U3314 (N_3314,N_3154,N_3139);
nand U3315 (N_3315,N_3070,N_3051);
or U3316 (N_3316,N_3181,N_3132);
nand U3317 (N_3317,N_3001,N_3003);
nand U3318 (N_3318,N_3068,N_3191);
nand U3319 (N_3319,N_3117,N_3112);
or U3320 (N_3320,N_3008,N_3109);
nor U3321 (N_3321,N_3157,N_3110);
nand U3322 (N_3322,N_3144,N_3198);
nand U3323 (N_3323,N_3144,N_3086);
or U3324 (N_3324,N_3151,N_3043);
and U3325 (N_3325,N_3141,N_3111);
nor U3326 (N_3326,N_3083,N_3193);
nor U3327 (N_3327,N_3175,N_3092);
and U3328 (N_3328,N_3020,N_3139);
xnor U3329 (N_3329,N_3182,N_3143);
or U3330 (N_3330,N_3108,N_3119);
or U3331 (N_3331,N_3083,N_3122);
or U3332 (N_3332,N_3101,N_3181);
or U3333 (N_3333,N_3038,N_3111);
nand U3334 (N_3334,N_3097,N_3135);
xor U3335 (N_3335,N_3032,N_3147);
and U3336 (N_3336,N_3019,N_3027);
and U3337 (N_3337,N_3195,N_3019);
xor U3338 (N_3338,N_3135,N_3125);
or U3339 (N_3339,N_3027,N_3001);
xnor U3340 (N_3340,N_3090,N_3110);
nor U3341 (N_3341,N_3059,N_3126);
and U3342 (N_3342,N_3011,N_3124);
xnor U3343 (N_3343,N_3059,N_3119);
or U3344 (N_3344,N_3108,N_3150);
and U3345 (N_3345,N_3094,N_3135);
and U3346 (N_3346,N_3136,N_3198);
and U3347 (N_3347,N_3062,N_3192);
xnor U3348 (N_3348,N_3141,N_3186);
nand U3349 (N_3349,N_3157,N_3070);
or U3350 (N_3350,N_3188,N_3141);
and U3351 (N_3351,N_3121,N_3192);
or U3352 (N_3352,N_3046,N_3158);
nor U3353 (N_3353,N_3015,N_3008);
nor U3354 (N_3354,N_3145,N_3147);
nand U3355 (N_3355,N_3116,N_3192);
nand U3356 (N_3356,N_3185,N_3149);
or U3357 (N_3357,N_3076,N_3133);
nor U3358 (N_3358,N_3192,N_3093);
and U3359 (N_3359,N_3059,N_3127);
xor U3360 (N_3360,N_3152,N_3198);
nand U3361 (N_3361,N_3146,N_3169);
xor U3362 (N_3362,N_3043,N_3082);
xor U3363 (N_3363,N_3117,N_3181);
xor U3364 (N_3364,N_3104,N_3010);
nand U3365 (N_3365,N_3028,N_3077);
or U3366 (N_3366,N_3188,N_3189);
nand U3367 (N_3367,N_3061,N_3054);
nor U3368 (N_3368,N_3186,N_3179);
nand U3369 (N_3369,N_3101,N_3033);
xor U3370 (N_3370,N_3182,N_3057);
xor U3371 (N_3371,N_3195,N_3122);
or U3372 (N_3372,N_3075,N_3159);
xor U3373 (N_3373,N_3028,N_3008);
nand U3374 (N_3374,N_3005,N_3075);
nor U3375 (N_3375,N_3184,N_3102);
nor U3376 (N_3376,N_3159,N_3060);
and U3377 (N_3377,N_3105,N_3187);
nor U3378 (N_3378,N_3031,N_3058);
nand U3379 (N_3379,N_3163,N_3151);
and U3380 (N_3380,N_3087,N_3150);
or U3381 (N_3381,N_3130,N_3181);
or U3382 (N_3382,N_3141,N_3161);
and U3383 (N_3383,N_3187,N_3185);
xor U3384 (N_3384,N_3052,N_3061);
and U3385 (N_3385,N_3026,N_3151);
xnor U3386 (N_3386,N_3045,N_3100);
nor U3387 (N_3387,N_3132,N_3091);
xnor U3388 (N_3388,N_3133,N_3130);
and U3389 (N_3389,N_3189,N_3184);
and U3390 (N_3390,N_3184,N_3087);
nor U3391 (N_3391,N_3093,N_3143);
nor U3392 (N_3392,N_3167,N_3100);
or U3393 (N_3393,N_3148,N_3181);
and U3394 (N_3394,N_3025,N_3185);
nand U3395 (N_3395,N_3047,N_3049);
or U3396 (N_3396,N_3126,N_3176);
nor U3397 (N_3397,N_3116,N_3011);
nor U3398 (N_3398,N_3161,N_3165);
and U3399 (N_3399,N_3166,N_3153);
or U3400 (N_3400,N_3377,N_3298);
and U3401 (N_3401,N_3273,N_3254);
and U3402 (N_3402,N_3383,N_3336);
xor U3403 (N_3403,N_3361,N_3321);
nor U3404 (N_3404,N_3262,N_3304);
xor U3405 (N_3405,N_3270,N_3268);
and U3406 (N_3406,N_3312,N_3307);
nor U3407 (N_3407,N_3333,N_3286);
xnor U3408 (N_3408,N_3386,N_3330);
and U3409 (N_3409,N_3288,N_3300);
and U3410 (N_3410,N_3311,N_3347);
nor U3411 (N_3411,N_3337,N_3221);
or U3412 (N_3412,N_3399,N_3257);
or U3413 (N_3413,N_3381,N_3244);
nor U3414 (N_3414,N_3385,N_3329);
xnor U3415 (N_3415,N_3351,N_3348);
xor U3416 (N_3416,N_3365,N_3252);
nand U3417 (N_3417,N_3282,N_3261);
and U3418 (N_3418,N_3342,N_3245);
nand U3419 (N_3419,N_3396,N_3322);
xnor U3420 (N_3420,N_3229,N_3379);
and U3421 (N_3421,N_3320,N_3258);
xnor U3422 (N_3422,N_3253,N_3214);
xnor U3423 (N_3423,N_3217,N_3296);
nand U3424 (N_3424,N_3271,N_3269);
and U3425 (N_3425,N_3393,N_3332);
and U3426 (N_3426,N_3309,N_3387);
or U3427 (N_3427,N_3389,N_3220);
or U3428 (N_3428,N_3362,N_3205);
xor U3429 (N_3429,N_3204,N_3283);
and U3430 (N_3430,N_3340,N_3265);
nor U3431 (N_3431,N_3266,N_3302);
and U3432 (N_3432,N_3316,N_3276);
or U3433 (N_3433,N_3228,N_3346);
xnor U3434 (N_3434,N_3289,N_3334);
or U3435 (N_3435,N_3281,N_3236);
and U3436 (N_3436,N_3297,N_3323);
or U3437 (N_3437,N_3219,N_3203);
or U3438 (N_3438,N_3248,N_3212);
nor U3439 (N_3439,N_3339,N_3235);
or U3440 (N_3440,N_3325,N_3284);
or U3441 (N_3441,N_3200,N_3314);
nand U3442 (N_3442,N_3210,N_3263);
xor U3443 (N_3443,N_3274,N_3357);
and U3444 (N_3444,N_3260,N_3301);
xnor U3445 (N_3445,N_3319,N_3291);
and U3446 (N_3446,N_3318,N_3224);
nor U3447 (N_3447,N_3279,N_3369);
nand U3448 (N_3448,N_3264,N_3292);
nor U3449 (N_3449,N_3324,N_3354);
or U3450 (N_3450,N_3384,N_3306);
xor U3451 (N_3451,N_3207,N_3211);
nor U3452 (N_3452,N_3255,N_3237);
or U3453 (N_3453,N_3315,N_3380);
and U3454 (N_3454,N_3226,N_3375);
nor U3455 (N_3455,N_3215,N_3397);
and U3456 (N_3456,N_3326,N_3238);
nor U3457 (N_3457,N_3367,N_3338);
nand U3458 (N_3458,N_3216,N_3349);
or U3459 (N_3459,N_3382,N_3390);
xor U3460 (N_3460,N_3287,N_3294);
nor U3461 (N_3461,N_3267,N_3366);
nand U3462 (N_3462,N_3213,N_3327);
xor U3463 (N_3463,N_3355,N_3372);
nor U3464 (N_3464,N_3232,N_3356);
and U3465 (N_3465,N_3370,N_3395);
or U3466 (N_3466,N_3303,N_3280);
nand U3467 (N_3467,N_3225,N_3305);
nor U3468 (N_3468,N_3368,N_3222);
and U3469 (N_3469,N_3388,N_3308);
nor U3470 (N_3470,N_3239,N_3364);
nor U3471 (N_3471,N_3359,N_3352);
and U3472 (N_3472,N_3247,N_3344);
nand U3473 (N_3473,N_3335,N_3317);
nand U3474 (N_3474,N_3313,N_3394);
nor U3475 (N_3475,N_3230,N_3251);
and U3476 (N_3476,N_3240,N_3241);
xor U3477 (N_3477,N_3360,N_3345);
and U3478 (N_3478,N_3272,N_3206);
nor U3479 (N_3479,N_3285,N_3256);
nand U3480 (N_3480,N_3246,N_3278);
nor U3481 (N_3481,N_3227,N_3392);
and U3482 (N_3482,N_3293,N_3341);
nand U3483 (N_3483,N_3259,N_3231);
nand U3484 (N_3484,N_3331,N_3391);
xnor U3485 (N_3485,N_3234,N_3250);
nand U3486 (N_3486,N_3242,N_3373);
or U3487 (N_3487,N_3218,N_3363);
and U3488 (N_3488,N_3343,N_3202);
nor U3489 (N_3489,N_3295,N_3249);
nor U3490 (N_3490,N_3378,N_3328);
nand U3491 (N_3491,N_3233,N_3376);
nand U3492 (N_3492,N_3299,N_3290);
nand U3493 (N_3493,N_3277,N_3374);
xor U3494 (N_3494,N_3353,N_3223);
nand U3495 (N_3495,N_3201,N_3208);
and U3496 (N_3496,N_3371,N_3350);
nor U3497 (N_3497,N_3275,N_3358);
nand U3498 (N_3498,N_3243,N_3209);
or U3499 (N_3499,N_3398,N_3310);
or U3500 (N_3500,N_3230,N_3342);
nand U3501 (N_3501,N_3312,N_3326);
or U3502 (N_3502,N_3254,N_3228);
xnor U3503 (N_3503,N_3341,N_3218);
and U3504 (N_3504,N_3385,N_3281);
nand U3505 (N_3505,N_3394,N_3276);
nor U3506 (N_3506,N_3387,N_3352);
xnor U3507 (N_3507,N_3250,N_3244);
or U3508 (N_3508,N_3349,N_3385);
xnor U3509 (N_3509,N_3238,N_3237);
xnor U3510 (N_3510,N_3298,N_3312);
or U3511 (N_3511,N_3237,N_3246);
and U3512 (N_3512,N_3202,N_3278);
nand U3513 (N_3513,N_3348,N_3257);
or U3514 (N_3514,N_3385,N_3344);
nand U3515 (N_3515,N_3312,N_3334);
nor U3516 (N_3516,N_3395,N_3238);
xnor U3517 (N_3517,N_3226,N_3240);
and U3518 (N_3518,N_3307,N_3283);
or U3519 (N_3519,N_3279,N_3333);
nor U3520 (N_3520,N_3239,N_3344);
nor U3521 (N_3521,N_3396,N_3204);
nor U3522 (N_3522,N_3313,N_3289);
xnor U3523 (N_3523,N_3256,N_3312);
nor U3524 (N_3524,N_3202,N_3362);
xnor U3525 (N_3525,N_3315,N_3252);
and U3526 (N_3526,N_3345,N_3204);
nand U3527 (N_3527,N_3252,N_3215);
xor U3528 (N_3528,N_3261,N_3254);
and U3529 (N_3529,N_3288,N_3380);
nand U3530 (N_3530,N_3294,N_3296);
and U3531 (N_3531,N_3216,N_3317);
nand U3532 (N_3532,N_3263,N_3365);
and U3533 (N_3533,N_3222,N_3257);
nand U3534 (N_3534,N_3262,N_3333);
nor U3535 (N_3535,N_3374,N_3266);
or U3536 (N_3536,N_3228,N_3378);
or U3537 (N_3537,N_3280,N_3274);
nand U3538 (N_3538,N_3269,N_3376);
or U3539 (N_3539,N_3377,N_3360);
or U3540 (N_3540,N_3204,N_3332);
xor U3541 (N_3541,N_3233,N_3298);
and U3542 (N_3542,N_3264,N_3242);
nor U3543 (N_3543,N_3376,N_3287);
nor U3544 (N_3544,N_3336,N_3386);
or U3545 (N_3545,N_3371,N_3284);
nor U3546 (N_3546,N_3330,N_3259);
nand U3547 (N_3547,N_3274,N_3279);
or U3548 (N_3548,N_3229,N_3393);
and U3549 (N_3549,N_3319,N_3260);
and U3550 (N_3550,N_3310,N_3273);
xnor U3551 (N_3551,N_3210,N_3285);
xor U3552 (N_3552,N_3388,N_3228);
and U3553 (N_3553,N_3349,N_3206);
xnor U3554 (N_3554,N_3229,N_3317);
or U3555 (N_3555,N_3285,N_3320);
and U3556 (N_3556,N_3308,N_3353);
xor U3557 (N_3557,N_3267,N_3316);
or U3558 (N_3558,N_3210,N_3336);
and U3559 (N_3559,N_3289,N_3210);
nor U3560 (N_3560,N_3242,N_3274);
nand U3561 (N_3561,N_3381,N_3252);
nor U3562 (N_3562,N_3278,N_3389);
and U3563 (N_3563,N_3326,N_3217);
nor U3564 (N_3564,N_3362,N_3271);
and U3565 (N_3565,N_3395,N_3206);
or U3566 (N_3566,N_3270,N_3309);
nand U3567 (N_3567,N_3307,N_3270);
xnor U3568 (N_3568,N_3397,N_3378);
and U3569 (N_3569,N_3278,N_3255);
and U3570 (N_3570,N_3229,N_3372);
nor U3571 (N_3571,N_3231,N_3388);
xnor U3572 (N_3572,N_3224,N_3273);
nand U3573 (N_3573,N_3333,N_3223);
or U3574 (N_3574,N_3269,N_3335);
xor U3575 (N_3575,N_3361,N_3269);
nor U3576 (N_3576,N_3254,N_3282);
or U3577 (N_3577,N_3208,N_3319);
xnor U3578 (N_3578,N_3397,N_3365);
nor U3579 (N_3579,N_3333,N_3396);
or U3580 (N_3580,N_3323,N_3210);
xor U3581 (N_3581,N_3346,N_3290);
xor U3582 (N_3582,N_3252,N_3380);
or U3583 (N_3583,N_3399,N_3383);
and U3584 (N_3584,N_3210,N_3311);
nor U3585 (N_3585,N_3302,N_3215);
nand U3586 (N_3586,N_3327,N_3263);
xnor U3587 (N_3587,N_3390,N_3209);
nand U3588 (N_3588,N_3377,N_3220);
or U3589 (N_3589,N_3312,N_3328);
or U3590 (N_3590,N_3232,N_3273);
xnor U3591 (N_3591,N_3204,N_3379);
xnor U3592 (N_3592,N_3347,N_3263);
xnor U3593 (N_3593,N_3280,N_3273);
xor U3594 (N_3594,N_3357,N_3269);
nand U3595 (N_3595,N_3364,N_3291);
or U3596 (N_3596,N_3281,N_3282);
nand U3597 (N_3597,N_3329,N_3259);
and U3598 (N_3598,N_3355,N_3376);
nor U3599 (N_3599,N_3200,N_3315);
and U3600 (N_3600,N_3485,N_3574);
nand U3601 (N_3601,N_3403,N_3593);
or U3602 (N_3602,N_3443,N_3456);
xor U3603 (N_3603,N_3478,N_3514);
and U3604 (N_3604,N_3544,N_3445);
nand U3605 (N_3605,N_3536,N_3554);
and U3606 (N_3606,N_3557,N_3413);
nor U3607 (N_3607,N_3515,N_3429);
nand U3608 (N_3608,N_3532,N_3498);
nand U3609 (N_3609,N_3434,N_3463);
xnor U3610 (N_3610,N_3573,N_3523);
nor U3611 (N_3611,N_3419,N_3596);
and U3612 (N_3612,N_3583,N_3561);
xnor U3613 (N_3613,N_3531,N_3407);
nor U3614 (N_3614,N_3497,N_3422);
nor U3615 (N_3615,N_3464,N_3440);
xnor U3616 (N_3616,N_3468,N_3470);
nand U3617 (N_3617,N_3472,N_3517);
and U3618 (N_3618,N_3474,N_3473);
nor U3619 (N_3619,N_3550,N_3427);
nand U3620 (N_3620,N_3584,N_3476);
nor U3621 (N_3621,N_3452,N_3538);
nand U3622 (N_3622,N_3436,N_3426);
xor U3623 (N_3623,N_3490,N_3585);
xnor U3624 (N_3624,N_3423,N_3562);
nand U3625 (N_3625,N_3457,N_3552);
and U3626 (N_3626,N_3495,N_3526);
or U3627 (N_3627,N_3568,N_3520);
xor U3628 (N_3628,N_3444,N_3535);
nor U3629 (N_3629,N_3494,N_3553);
xnor U3630 (N_3630,N_3459,N_3433);
xor U3631 (N_3631,N_3489,N_3591);
nand U3632 (N_3632,N_3416,N_3549);
nand U3633 (N_3633,N_3481,N_3518);
xnor U3634 (N_3634,N_3402,N_3493);
and U3635 (N_3635,N_3466,N_3516);
nand U3636 (N_3636,N_3559,N_3590);
xnor U3637 (N_3637,N_3558,N_3527);
and U3638 (N_3638,N_3533,N_3406);
or U3639 (N_3639,N_3521,N_3502);
nand U3640 (N_3640,N_3505,N_3408);
or U3641 (N_3641,N_3578,N_3400);
and U3642 (N_3642,N_3556,N_3477);
xnor U3643 (N_3643,N_3441,N_3420);
and U3644 (N_3644,N_3415,N_3582);
or U3645 (N_3645,N_3597,N_3563);
xor U3646 (N_3646,N_3491,N_3525);
nand U3647 (N_3647,N_3453,N_3479);
and U3648 (N_3648,N_3486,N_3522);
nand U3649 (N_3649,N_3487,N_3462);
nand U3650 (N_3650,N_3537,N_3542);
xnor U3651 (N_3651,N_3586,N_3430);
xor U3652 (N_3652,N_3409,N_3460);
xnor U3653 (N_3653,N_3576,N_3581);
xnor U3654 (N_3654,N_3411,N_3572);
xnor U3655 (N_3655,N_3566,N_3543);
and U3656 (N_3656,N_3418,N_3571);
nand U3657 (N_3657,N_3529,N_3555);
nor U3658 (N_3658,N_3579,N_3507);
and U3659 (N_3659,N_3524,N_3528);
and U3660 (N_3660,N_3501,N_3417);
nor U3661 (N_3661,N_3428,N_3570);
nor U3662 (N_3662,N_3421,N_3503);
nor U3663 (N_3663,N_3432,N_3437);
and U3664 (N_3664,N_3480,N_3450);
and U3665 (N_3665,N_3425,N_3404);
nand U3666 (N_3666,N_3500,N_3492);
nor U3667 (N_3667,N_3565,N_3449);
or U3668 (N_3668,N_3469,N_3564);
xnor U3669 (N_3669,N_3438,N_3513);
and U3670 (N_3670,N_3431,N_3599);
xnor U3671 (N_3671,N_3580,N_3448);
nand U3672 (N_3672,N_3465,N_3598);
nor U3673 (N_3673,N_3589,N_3519);
nor U3674 (N_3674,N_3483,N_3512);
and U3675 (N_3675,N_3587,N_3509);
nand U3676 (N_3676,N_3551,N_3410);
nand U3677 (N_3677,N_3592,N_3414);
nand U3678 (N_3678,N_3442,N_3546);
and U3679 (N_3679,N_3504,N_3508);
nor U3680 (N_3680,N_3567,N_3439);
and U3681 (N_3681,N_3412,N_3540);
nand U3682 (N_3682,N_3547,N_3510);
xnor U3683 (N_3683,N_3401,N_3455);
and U3684 (N_3684,N_3545,N_3541);
and U3685 (N_3685,N_3506,N_3446);
xor U3686 (N_3686,N_3467,N_3569);
and U3687 (N_3687,N_3560,N_3451);
or U3688 (N_3688,N_3488,N_3594);
or U3689 (N_3689,N_3471,N_3454);
and U3690 (N_3690,N_3405,N_3511);
xor U3691 (N_3691,N_3499,N_3475);
or U3692 (N_3692,N_3424,N_3595);
or U3693 (N_3693,N_3577,N_3530);
nand U3694 (N_3694,N_3447,N_3496);
and U3695 (N_3695,N_3482,N_3588);
nor U3696 (N_3696,N_3575,N_3461);
xor U3697 (N_3697,N_3539,N_3435);
nor U3698 (N_3698,N_3534,N_3458);
xor U3699 (N_3699,N_3548,N_3484);
nand U3700 (N_3700,N_3432,N_3481);
and U3701 (N_3701,N_3425,N_3570);
nand U3702 (N_3702,N_3513,N_3582);
xor U3703 (N_3703,N_3453,N_3492);
and U3704 (N_3704,N_3546,N_3529);
xnor U3705 (N_3705,N_3424,N_3442);
nand U3706 (N_3706,N_3545,N_3517);
or U3707 (N_3707,N_3485,N_3442);
nand U3708 (N_3708,N_3467,N_3566);
or U3709 (N_3709,N_3536,N_3433);
and U3710 (N_3710,N_3516,N_3508);
nand U3711 (N_3711,N_3551,N_3406);
or U3712 (N_3712,N_3494,N_3546);
nand U3713 (N_3713,N_3439,N_3422);
or U3714 (N_3714,N_3563,N_3539);
and U3715 (N_3715,N_3579,N_3531);
nand U3716 (N_3716,N_3488,N_3420);
nor U3717 (N_3717,N_3525,N_3417);
nand U3718 (N_3718,N_3564,N_3525);
or U3719 (N_3719,N_3501,N_3568);
nand U3720 (N_3720,N_3474,N_3569);
and U3721 (N_3721,N_3493,N_3408);
and U3722 (N_3722,N_3579,N_3528);
xnor U3723 (N_3723,N_3454,N_3537);
xor U3724 (N_3724,N_3433,N_3432);
nor U3725 (N_3725,N_3431,N_3554);
or U3726 (N_3726,N_3548,N_3408);
or U3727 (N_3727,N_3574,N_3481);
nand U3728 (N_3728,N_3578,N_3509);
or U3729 (N_3729,N_3445,N_3556);
nor U3730 (N_3730,N_3593,N_3525);
xnor U3731 (N_3731,N_3473,N_3512);
and U3732 (N_3732,N_3501,N_3531);
xnor U3733 (N_3733,N_3431,N_3586);
nor U3734 (N_3734,N_3528,N_3497);
xor U3735 (N_3735,N_3433,N_3556);
nor U3736 (N_3736,N_3507,N_3483);
nand U3737 (N_3737,N_3563,N_3514);
nand U3738 (N_3738,N_3547,N_3505);
xor U3739 (N_3739,N_3592,N_3537);
nor U3740 (N_3740,N_3550,N_3549);
nor U3741 (N_3741,N_3565,N_3441);
nand U3742 (N_3742,N_3550,N_3422);
nand U3743 (N_3743,N_3476,N_3477);
nand U3744 (N_3744,N_3585,N_3435);
and U3745 (N_3745,N_3586,N_3526);
nor U3746 (N_3746,N_3520,N_3509);
xor U3747 (N_3747,N_3548,N_3425);
and U3748 (N_3748,N_3444,N_3511);
and U3749 (N_3749,N_3570,N_3578);
nor U3750 (N_3750,N_3419,N_3478);
or U3751 (N_3751,N_3565,N_3582);
nand U3752 (N_3752,N_3423,N_3409);
nand U3753 (N_3753,N_3416,N_3561);
xor U3754 (N_3754,N_3542,N_3444);
and U3755 (N_3755,N_3473,N_3437);
nand U3756 (N_3756,N_3478,N_3581);
and U3757 (N_3757,N_3517,N_3577);
or U3758 (N_3758,N_3507,N_3496);
xor U3759 (N_3759,N_3492,N_3445);
nand U3760 (N_3760,N_3531,N_3491);
or U3761 (N_3761,N_3428,N_3496);
xnor U3762 (N_3762,N_3423,N_3526);
xor U3763 (N_3763,N_3412,N_3401);
xor U3764 (N_3764,N_3597,N_3498);
or U3765 (N_3765,N_3504,N_3585);
or U3766 (N_3766,N_3592,N_3570);
nor U3767 (N_3767,N_3470,N_3575);
or U3768 (N_3768,N_3454,N_3473);
or U3769 (N_3769,N_3518,N_3441);
nor U3770 (N_3770,N_3451,N_3453);
nor U3771 (N_3771,N_3422,N_3447);
and U3772 (N_3772,N_3529,N_3549);
or U3773 (N_3773,N_3596,N_3552);
nor U3774 (N_3774,N_3435,N_3486);
xnor U3775 (N_3775,N_3519,N_3547);
xor U3776 (N_3776,N_3510,N_3540);
nand U3777 (N_3777,N_3439,N_3594);
nor U3778 (N_3778,N_3473,N_3560);
xor U3779 (N_3779,N_3506,N_3498);
or U3780 (N_3780,N_3527,N_3478);
xor U3781 (N_3781,N_3516,N_3405);
or U3782 (N_3782,N_3467,N_3558);
xnor U3783 (N_3783,N_3437,N_3558);
xnor U3784 (N_3784,N_3468,N_3578);
xnor U3785 (N_3785,N_3499,N_3486);
nor U3786 (N_3786,N_3469,N_3485);
or U3787 (N_3787,N_3409,N_3451);
or U3788 (N_3788,N_3458,N_3558);
nor U3789 (N_3789,N_3597,N_3565);
nand U3790 (N_3790,N_3525,N_3443);
nand U3791 (N_3791,N_3484,N_3497);
or U3792 (N_3792,N_3463,N_3553);
or U3793 (N_3793,N_3505,N_3581);
xnor U3794 (N_3794,N_3415,N_3544);
or U3795 (N_3795,N_3440,N_3578);
or U3796 (N_3796,N_3440,N_3595);
xor U3797 (N_3797,N_3516,N_3565);
and U3798 (N_3798,N_3418,N_3548);
nor U3799 (N_3799,N_3513,N_3448);
nand U3800 (N_3800,N_3693,N_3669);
and U3801 (N_3801,N_3628,N_3632);
nand U3802 (N_3802,N_3666,N_3723);
and U3803 (N_3803,N_3655,N_3785);
or U3804 (N_3804,N_3694,N_3768);
xnor U3805 (N_3805,N_3659,N_3795);
nand U3806 (N_3806,N_3664,N_3704);
nand U3807 (N_3807,N_3796,N_3620);
xnor U3808 (N_3808,N_3700,N_3654);
nor U3809 (N_3809,N_3610,N_3744);
and U3810 (N_3810,N_3719,N_3641);
xor U3811 (N_3811,N_3626,N_3609);
nand U3812 (N_3812,N_3683,N_3726);
nor U3813 (N_3813,N_3707,N_3789);
nor U3814 (N_3814,N_3710,N_3797);
and U3815 (N_3815,N_3625,N_3601);
and U3816 (N_3816,N_3703,N_3662);
or U3817 (N_3817,N_3712,N_3756);
nor U3818 (N_3818,N_3720,N_3794);
nor U3819 (N_3819,N_3663,N_3758);
nor U3820 (N_3820,N_3631,N_3600);
and U3821 (N_3821,N_3754,N_3698);
xnor U3822 (N_3822,N_3672,N_3781);
nor U3823 (N_3823,N_3671,N_3675);
and U3824 (N_3824,N_3642,N_3779);
and U3825 (N_3825,N_3790,N_3697);
nor U3826 (N_3826,N_3616,N_3660);
or U3827 (N_3827,N_3604,N_3748);
nor U3828 (N_3828,N_3611,N_3668);
nand U3829 (N_3829,N_3645,N_3784);
xnor U3830 (N_3830,N_3711,N_3617);
xor U3831 (N_3831,N_3742,N_3753);
nor U3832 (N_3832,N_3708,N_3636);
nand U3833 (N_3833,N_3691,N_3747);
or U3834 (N_3834,N_3679,N_3650);
nand U3835 (N_3835,N_3637,N_3714);
xor U3836 (N_3836,N_3640,N_3653);
xnor U3837 (N_3837,N_3741,N_3643);
nor U3838 (N_3838,N_3762,N_3721);
or U3839 (N_3839,N_3791,N_3749);
and U3840 (N_3840,N_3624,N_3673);
or U3841 (N_3841,N_3738,N_3761);
xnor U3842 (N_3842,N_3674,N_3798);
nand U3843 (N_3843,N_3792,N_3687);
xor U3844 (N_3844,N_3713,N_3648);
nand U3845 (N_3845,N_3799,N_3770);
or U3846 (N_3846,N_3715,N_3706);
nor U3847 (N_3847,N_3782,N_3705);
nand U3848 (N_3848,N_3733,N_3746);
xor U3849 (N_3849,N_3676,N_3651);
and U3850 (N_3850,N_3670,N_3685);
nor U3851 (N_3851,N_3729,N_3734);
xor U3852 (N_3852,N_3760,N_3725);
nand U3853 (N_3853,N_3627,N_3658);
nand U3854 (N_3854,N_3739,N_3647);
and U3855 (N_3855,N_3765,N_3757);
or U3856 (N_3856,N_3772,N_3764);
and U3857 (N_3857,N_3718,N_3656);
nor U3858 (N_3858,N_3727,N_3716);
xor U3859 (N_3859,N_3633,N_3638);
or U3860 (N_3860,N_3773,N_3689);
xnor U3861 (N_3861,N_3690,N_3682);
or U3862 (N_3862,N_3665,N_3684);
nor U3863 (N_3863,N_3606,N_3692);
xor U3864 (N_3864,N_3759,N_3728);
nor U3865 (N_3865,N_3783,N_3750);
xnor U3866 (N_3866,N_3788,N_3735);
and U3867 (N_3867,N_3639,N_3724);
nand U3868 (N_3868,N_3777,N_3612);
xnor U3869 (N_3869,N_3615,N_3769);
or U3870 (N_3870,N_3786,N_3623);
nor U3871 (N_3871,N_3709,N_3767);
nor U3872 (N_3872,N_3730,N_3635);
nor U3873 (N_3873,N_3774,N_3732);
and U3874 (N_3874,N_3766,N_3644);
or U3875 (N_3875,N_3752,N_3717);
and U3876 (N_3876,N_3613,N_3787);
and U3877 (N_3877,N_3776,N_3618);
nand U3878 (N_3878,N_3661,N_3677);
or U3879 (N_3879,N_3745,N_3680);
and U3880 (N_3880,N_3621,N_3736);
or U3881 (N_3881,N_3619,N_3740);
nand U3882 (N_3882,N_3702,N_3743);
or U3883 (N_3883,N_3649,N_3771);
or U3884 (N_3884,N_3780,N_3630);
nor U3885 (N_3885,N_3763,N_3731);
xnor U3886 (N_3886,N_3614,N_3629);
or U3887 (N_3887,N_3751,N_3605);
nor U3888 (N_3888,N_3608,N_3622);
xnor U3889 (N_3889,N_3699,N_3667);
and U3890 (N_3890,N_3778,N_3607);
xor U3891 (N_3891,N_3634,N_3695);
and U3892 (N_3892,N_3722,N_3652);
nor U3893 (N_3893,N_3775,N_3737);
nor U3894 (N_3894,N_3678,N_3657);
nor U3895 (N_3895,N_3688,N_3696);
or U3896 (N_3896,N_3755,N_3793);
nand U3897 (N_3897,N_3701,N_3646);
nand U3898 (N_3898,N_3681,N_3603);
and U3899 (N_3899,N_3686,N_3602);
and U3900 (N_3900,N_3622,N_3632);
nor U3901 (N_3901,N_3721,N_3704);
or U3902 (N_3902,N_3642,N_3777);
xnor U3903 (N_3903,N_3611,N_3760);
nand U3904 (N_3904,N_3603,N_3634);
nor U3905 (N_3905,N_3648,N_3644);
xor U3906 (N_3906,N_3790,N_3664);
nor U3907 (N_3907,N_3744,N_3730);
xnor U3908 (N_3908,N_3679,N_3633);
and U3909 (N_3909,N_3715,N_3766);
and U3910 (N_3910,N_3707,N_3786);
nand U3911 (N_3911,N_3668,N_3678);
xor U3912 (N_3912,N_3740,N_3798);
nand U3913 (N_3913,N_3654,N_3687);
nand U3914 (N_3914,N_3709,N_3788);
nor U3915 (N_3915,N_3744,N_3663);
xnor U3916 (N_3916,N_3711,N_3722);
and U3917 (N_3917,N_3676,N_3609);
and U3918 (N_3918,N_3769,N_3665);
nor U3919 (N_3919,N_3722,N_3634);
xor U3920 (N_3920,N_3765,N_3660);
or U3921 (N_3921,N_3609,N_3751);
and U3922 (N_3922,N_3691,N_3701);
or U3923 (N_3923,N_3675,N_3736);
nand U3924 (N_3924,N_3601,N_3648);
or U3925 (N_3925,N_3645,N_3753);
and U3926 (N_3926,N_3676,N_3660);
and U3927 (N_3927,N_3662,N_3734);
nor U3928 (N_3928,N_3680,N_3627);
nand U3929 (N_3929,N_3784,N_3685);
xor U3930 (N_3930,N_3668,N_3615);
nor U3931 (N_3931,N_3636,N_3630);
xor U3932 (N_3932,N_3674,N_3789);
or U3933 (N_3933,N_3660,N_3669);
nand U3934 (N_3934,N_3617,N_3770);
nand U3935 (N_3935,N_3708,N_3791);
and U3936 (N_3936,N_3733,N_3634);
and U3937 (N_3937,N_3742,N_3721);
or U3938 (N_3938,N_3660,N_3611);
or U3939 (N_3939,N_3691,N_3787);
and U3940 (N_3940,N_3768,N_3637);
and U3941 (N_3941,N_3636,N_3729);
nor U3942 (N_3942,N_3608,N_3630);
xor U3943 (N_3943,N_3667,N_3676);
or U3944 (N_3944,N_3662,N_3617);
or U3945 (N_3945,N_3661,N_3698);
xnor U3946 (N_3946,N_3709,N_3668);
or U3947 (N_3947,N_3668,N_3692);
nor U3948 (N_3948,N_3797,N_3768);
nand U3949 (N_3949,N_3732,N_3639);
nor U3950 (N_3950,N_3601,N_3771);
or U3951 (N_3951,N_3602,N_3750);
nand U3952 (N_3952,N_3682,N_3684);
or U3953 (N_3953,N_3607,N_3772);
or U3954 (N_3954,N_3729,N_3712);
nor U3955 (N_3955,N_3730,N_3732);
or U3956 (N_3956,N_3654,N_3673);
nand U3957 (N_3957,N_3773,N_3706);
xnor U3958 (N_3958,N_3773,N_3736);
or U3959 (N_3959,N_3610,N_3784);
or U3960 (N_3960,N_3655,N_3671);
xor U3961 (N_3961,N_3745,N_3788);
xnor U3962 (N_3962,N_3772,N_3652);
nand U3963 (N_3963,N_3672,N_3715);
xnor U3964 (N_3964,N_3744,N_3778);
and U3965 (N_3965,N_3724,N_3753);
and U3966 (N_3966,N_3677,N_3795);
nor U3967 (N_3967,N_3747,N_3720);
xor U3968 (N_3968,N_3611,N_3737);
nor U3969 (N_3969,N_3616,N_3753);
or U3970 (N_3970,N_3679,N_3659);
nand U3971 (N_3971,N_3631,N_3768);
nand U3972 (N_3972,N_3716,N_3640);
xnor U3973 (N_3973,N_3717,N_3720);
and U3974 (N_3974,N_3679,N_3704);
and U3975 (N_3975,N_3617,N_3651);
xor U3976 (N_3976,N_3659,N_3639);
nand U3977 (N_3977,N_3728,N_3657);
nor U3978 (N_3978,N_3722,N_3710);
and U3979 (N_3979,N_3640,N_3751);
and U3980 (N_3980,N_3753,N_3780);
or U3981 (N_3981,N_3622,N_3637);
xor U3982 (N_3982,N_3710,N_3644);
nand U3983 (N_3983,N_3730,N_3682);
nor U3984 (N_3984,N_3765,N_3615);
nor U3985 (N_3985,N_3772,N_3670);
xnor U3986 (N_3986,N_3666,N_3774);
and U3987 (N_3987,N_3703,N_3640);
xor U3988 (N_3988,N_3685,N_3699);
nor U3989 (N_3989,N_3799,N_3736);
nor U3990 (N_3990,N_3671,N_3648);
or U3991 (N_3991,N_3600,N_3719);
nand U3992 (N_3992,N_3726,N_3658);
xor U3993 (N_3993,N_3721,N_3734);
xor U3994 (N_3994,N_3605,N_3799);
and U3995 (N_3995,N_3735,N_3790);
nand U3996 (N_3996,N_3768,N_3724);
or U3997 (N_3997,N_3603,N_3767);
xor U3998 (N_3998,N_3612,N_3711);
or U3999 (N_3999,N_3637,N_3725);
or U4000 (N_4000,N_3974,N_3914);
or U4001 (N_4001,N_3975,N_3809);
nand U4002 (N_4002,N_3905,N_3956);
nand U4003 (N_4003,N_3919,N_3811);
xor U4004 (N_4004,N_3904,N_3944);
and U4005 (N_4005,N_3964,N_3885);
and U4006 (N_4006,N_3961,N_3817);
and U4007 (N_4007,N_3854,N_3971);
xor U4008 (N_4008,N_3892,N_3827);
nor U4009 (N_4009,N_3823,N_3832);
xor U4010 (N_4010,N_3824,N_3967);
nand U4011 (N_4011,N_3868,N_3810);
and U4012 (N_4012,N_3951,N_3947);
or U4013 (N_4013,N_3935,N_3912);
nor U4014 (N_4014,N_3926,N_3902);
nand U4015 (N_4015,N_3894,N_3814);
and U4016 (N_4016,N_3922,N_3899);
nand U4017 (N_4017,N_3845,N_3909);
nand U4018 (N_4018,N_3865,N_3920);
xor U4019 (N_4019,N_3883,N_3988);
and U4020 (N_4020,N_3936,N_3999);
nor U4021 (N_4021,N_3896,N_3950);
nor U4022 (N_4022,N_3934,N_3867);
xor U4023 (N_4023,N_3957,N_3958);
nand U4024 (N_4024,N_3910,N_3943);
nand U4025 (N_4025,N_3986,N_3853);
or U4026 (N_4026,N_3913,N_3859);
and U4027 (N_4027,N_3812,N_3887);
nor U4028 (N_4028,N_3939,N_3820);
and U4029 (N_4029,N_3960,N_3816);
xor U4030 (N_4030,N_3856,N_3857);
and U4031 (N_4031,N_3846,N_3860);
nand U4032 (N_4032,N_3869,N_3979);
or U4033 (N_4033,N_3888,N_3933);
nand U4034 (N_4034,N_3841,N_3833);
and U4035 (N_4035,N_3929,N_3901);
nand U4036 (N_4036,N_3927,N_3992);
xor U4037 (N_4037,N_3828,N_3953);
and U4038 (N_4038,N_3965,N_3879);
nor U4039 (N_4039,N_3991,N_3973);
xor U4040 (N_4040,N_3848,N_3923);
and U4041 (N_4041,N_3825,N_3838);
and U4042 (N_4042,N_3878,N_3954);
nor U4043 (N_4043,N_3819,N_3842);
nand U4044 (N_4044,N_3863,N_3995);
nand U4045 (N_4045,N_3998,N_3807);
nor U4046 (N_4046,N_3835,N_3941);
nor U4047 (N_4047,N_3800,N_3925);
nor U4048 (N_4048,N_3806,N_3959);
nand U4049 (N_4049,N_3866,N_3937);
or U4050 (N_4050,N_3963,N_3900);
and U4051 (N_4051,N_3884,N_3803);
nor U4052 (N_4052,N_3906,N_3874);
or U4053 (N_4053,N_3969,N_3968);
xor U4054 (N_4054,N_3924,N_3898);
nor U4055 (N_4055,N_3952,N_3880);
and U4056 (N_4056,N_3847,N_3881);
nor U4057 (N_4057,N_3993,N_3976);
nor U4058 (N_4058,N_3897,N_3921);
nor U4059 (N_4059,N_3984,N_3990);
and U4060 (N_4060,N_3855,N_3882);
nor U4061 (N_4061,N_3858,N_3862);
xor U4062 (N_4062,N_3930,N_3802);
nand U4063 (N_4063,N_3821,N_3918);
nor U4064 (N_4064,N_3851,N_3946);
nand U4065 (N_4065,N_3895,N_3840);
or U4066 (N_4066,N_3945,N_3861);
xor U4067 (N_4067,N_3982,N_3916);
xnor U4068 (N_4068,N_3864,N_3911);
or U4069 (N_4069,N_3889,N_3890);
nand U4070 (N_4070,N_3996,N_3989);
xor U4071 (N_4071,N_3830,N_3938);
or U4072 (N_4072,N_3805,N_3873);
xnor U4073 (N_4073,N_3966,N_3822);
xnor U4074 (N_4074,N_3917,N_3849);
nor U4075 (N_4075,N_3962,N_3970);
or U4076 (N_4076,N_3907,N_3826);
xor U4077 (N_4077,N_3980,N_3829);
nand U4078 (N_4078,N_3804,N_3949);
or U4079 (N_4079,N_3948,N_3839);
nand U4080 (N_4080,N_3987,N_3837);
or U4081 (N_4081,N_3843,N_3985);
xnor U4082 (N_4082,N_3915,N_3836);
nand U4083 (N_4083,N_3981,N_3813);
or U4084 (N_4084,N_3942,N_3875);
nand U4085 (N_4085,N_3972,N_3891);
nand U4086 (N_4086,N_3932,N_3877);
xnor U4087 (N_4087,N_3831,N_3893);
nor U4088 (N_4088,N_3844,N_3834);
nand U4089 (N_4089,N_3928,N_3977);
xor U4090 (N_4090,N_3955,N_3818);
nor U4091 (N_4091,N_3801,N_3872);
or U4092 (N_4092,N_3994,N_3808);
xor U4093 (N_4093,N_3850,N_3931);
nor U4094 (N_4094,N_3876,N_3870);
or U4095 (N_4095,N_3852,N_3978);
and U4096 (N_4096,N_3908,N_3903);
xnor U4097 (N_4097,N_3871,N_3940);
nand U4098 (N_4098,N_3997,N_3983);
nand U4099 (N_4099,N_3815,N_3886);
and U4100 (N_4100,N_3971,N_3881);
nor U4101 (N_4101,N_3802,N_3846);
nor U4102 (N_4102,N_3962,N_3910);
nand U4103 (N_4103,N_3973,N_3945);
nor U4104 (N_4104,N_3842,N_3825);
nand U4105 (N_4105,N_3991,N_3902);
or U4106 (N_4106,N_3917,N_3996);
and U4107 (N_4107,N_3856,N_3918);
nand U4108 (N_4108,N_3877,N_3813);
xor U4109 (N_4109,N_3875,N_3826);
nor U4110 (N_4110,N_3979,N_3807);
or U4111 (N_4111,N_3957,N_3868);
nor U4112 (N_4112,N_3809,N_3903);
and U4113 (N_4113,N_3997,N_3810);
xor U4114 (N_4114,N_3902,N_3972);
and U4115 (N_4115,N_3829,N_3954);
nand U4116 (N_4116,N_3804,N_3901);
and U4117 (N_4117,N_3945,N_3871);
or U4118 (N_4118,N_3977,N_3911);
nand U4119 (N_4119,N_3843,N_3893);
or U4120 (N_4120,N_3982,N_3964);
nor U4121 (N_4121,N_3800,N_3821);
and U4122 (N_4122,N_3817,N_3947);
xnor U4123 (N_4123,N_3963,N_3937);
xor U4124 (N_4124,N_3895,N_3935);
or U4125 (N_4125,N_3818,N_3998);
and U4126 (N_4126,N_3871,N_3949);
nor U4127 (N_4127,N_3940,N_3955);
and U4128 (N_4128,N_3951,N_3840);
nor U4129 (N_4129,N_3890,N_3870);
xnor U4130 (N_4130,N_3953,N_3975);
nor U4131 (N_4131,N_3878,N_3930);
or U4132 (N_4132,N_3825,N_3950);
nand U4133 (N_4133,N_3881,N_3863);
xor U4134 (N_4134,N_3903,N_3829);
or U4135 (N_4135,N_3952,N_3892);
nor U4136 (N_4136,N_3939,N_3889);
nand U4137 (N_4137,N_3868,N_3869);
xor U4138 (N_4138,N_3952,N_3981);
and U4139 (N_4139,N_3834,N_3973);
nor U4140 (N_4140,N_3956,N_3962);
or U4141 (N_4141,N_3811,N_3839);
and U4142 (N_4142,N_3914,N_3989);
nand U4143 (N_4143,N_3975,N_3906);
and U4144 (N_4144,N_3926,N_3840);
nand U4145 (N_4145,N_3836,N_3897);
xnor U4146 (N_4146,N_3972,N_3814);
or U4147 (N_4147,N_3931,N_3882);
nor U4148 (N_4148,N_3958,N_3949);
and U4149 (N_4149,N_3983,N_3825);
nor U4150 (N_4150,N_3939,N_3956);
xor U4151 (N_4151,N_3803,N_3806);
or U4152 (N_4152,N_3828,N_3802);
nand U4153 (N_4153,N_3931,N_3962);
or U4154 (N_4154,N_3926,N_3803);
and U4155 (N_4155,N_3919,N_3852);
and U4156 (N_4156,N_3803,N_3825);
or U4157 (N_4157,N_3919,N_3956);
and U4158 (N_4158,N_3863,N_3938);
xnor U4159 (N_4159,N_3988,N_3851);
xor U4160 (N_4160,N_3911,N_3853);
xor U4161 (N_4161,N_3846,N_3923);
or U4162 (N_4162,N_3864,N_3821);
nor U4163 (N_4163,N_3929,N_3945);
xor U4164 (N_4164,N_3953,N_3928);
nand U4165 (N_4165,N_3878,N_3830);
nand U4166 (N_4166,N_3976,N_3924);
nor U4167 (N_4167,N_3987,N_3925);
or U4168 (N_4168,N_3906,N_3809);
nand U4169 (N_4169,N_3910,N_3834);
or U4170 (N_4170,N_3842,N_3956);
nand U4171 (N_4171,N_3894,N_3949);
nand U4172 (N_4172,N_3912,N_3826);
or U4173 (N_4173,N_3967,N_3875);
and U4174 (N_4174,N_3979,N_3853);
nand U4175 (N_4175,N_3961,N_3831);
or U4176 (N_4176,N_3894,N_3919);
nor U4177 (N_4177,N_3858,N_3873);
nor U4178 (N_4178,N_3966,N_3962);
xor U4179 (N_4179,N_3862,N_3871);
xnor U4180 (N_4180,N_3990,N_3882);
nand U4181 (N_4181,N_3878,N_3923);
and U4182 (N_4182,N_3857,N_3962);
or U4183 (N_4183,N_3917,N_3971);
xnor U4184 (N_4184,N_3889,N_3800);
nor U4185 (N_4185,N_3821,N_3857);
nor U4186 (N_4186,N_3922,N_3896);
nor U4187 (N_4187,N_3889,N_3968);
xor U4188 (N_4188,N_3942,N_3843);
and U4189 (N_4189,N_3903,N_3904);
nand U4190 (N_4190,N_3964,N_3998);
and U4191 (N_4191,N_3990,N_3951);
nor U4192 (N_4192,N_3976,N_3870);
nor U4193 (N_4193,N_3852,N_3805);
xnor U4194 (N_4194,N_3964,N_3842);
and U4195 (N_4195,N_3915,N_3827);
nand U4196 (N_4196,N_3999,N_3882);
and U4197 (N_4197,N_3834,N_3848);
xor U4198 (N_4198,N_3825,N_3877);
and U4199 (N_4199,N_3806,N_3960);
nand U4200 (N_4200,N_4147,N_4053);
xor U4201 (N_4201,N_4127,N_4051);
nand U4202 (N_4202,N_4008,N_4038);
nor U4203 (N_4203,N_4092,N_4026);
nand U4204 (N_4204,N_4137,N_4047);
or U4205 (N_4205,N_4090,N_4198);
nor U4206 (N_4206,N_4037,N_4152);
nor U4207 (N_4207,N_4154,N_4106);
nor U4208 (N_4208,N_4148,N_4141);
or U4209 (N_4209,N_4039,N_4173);
nor U4210 (N_4210,N_4097,N_4195);
and U4211 (N_4211,N_4065,N_4011);
or U4212 (N_4212,N_4183,N_4184);
nor U4213 (N_4213,N_4146,N_4132);
xnor U4214 (N_4214,N_4123,N_4061);
nand U4215 (N_4215,N_4176,N_4186);
xor U4216 (N_4216,N_4188,N_4006);
or U4217 (N_4217,N_4012,N_4165);
and U4218 (N_4218,N_4076,N_4111);
and U4219 (N_4219,N_4005,N_4187);
or U4220 (N_4220,N_4175,N_4018);
nand U4221 (N_4221,N_4072,N_4171);
nand U4222 (N_4222,N_4178,N_4044);
nand U4223 (N_4223,N_4113,N_4073);
and U4224 (N_4224,N_4059,N_4112);
and U4225 (N_4225,N_4172,N_4185);
or U4226 (N_4226,N_4189,N_4055);
nor U4227 (N_4227,N_4030,N_4182);
and U4228 (N_4228,N_4150,N_4046);
xor U4229 (N_4229,N_4194,N_4120);
nor U4230 (N_4230,N_4034,N_4010);
nor U4231 (N_4231,N_4041,N_4169);
or U4232 (N_4232,N_4036,N_4122);
xor U4233 (N_4233,N_4007,N_4089);
and U4234 (N_4234,N_4140,N_4049);
and U4235 (N_4235,N_4013,N_4192);
or U4236 (N_4236,N_4058,N_4079);
nand U4237 (N_4237,N_4048,N_4069);
nand U4238 (N_4238,N_4014,N_4093);
and U4239 (N_4239,N_4094,N_4144);
nand U4240 (N_4240,N_4100,N_4119);
nor U4241 (N_4241,N_4068,N_4096);
xor U4242 (N_4242,N_4027,N_4170);
xnor U4243 (N_4243,N_4168,N_4099);
and U4244 (N_4244,N_4057,N_4062);
and U4245 (N_4245,N_4110,N_4102);
xnor U4246 (N_4246,N_4009,N_4135);
xor U4247 (N_4247,N_4081,N_4043);
nand U4248 (N_4248,N_4136,N_4174);
xor U4249 (N_4249,N_4086,N_4087);
or U4250 (N_4250,N_4196,N_4021);
and U4251 (N_4251,N_4054,N_4035);
xor U4252 (N_4252,N_4180,N_4149);
nor U4253 (N_4253,N_4128,N_4143);
and U4254 (N_4254,N_4134,N_4129);
and U4255 (N_4255,N_4177,N_4131);
nand U4256 (N_4256,N_4060,N_4155);
or U4257 (N_4257,N_4045,N_4084);
xor U4258 (N_4258,N_4016,N_4157);
or U4259 (N_4259,N_4153,N_4190);
and U4260 (N_4260,N_4161,N_4164);
or U4261 (N_4261,N_4114,N_4108);
or U4262 (N_4262,N_4109,N_4004);
nand U4263 (N_4263,N_4124,N_4167);
or U4264 (N_4264,N_4101,N_4017);
xnor U4265 (N_4265,N_4103,N_4029);
nor U4266 (N_4266,N_4071,N_4197);
or U4267 (N_4267,N_4130,N_4085);
and U4268 (N_4268,N_4083,N_4158);
nand U4269 (N_4269,N_4080,N_4052);
or U4270 (N_4270,N_4142,N_4088);
nor U4271 (N_4271,N_4133,N_4078);
or U4272 (N_4272,N_4028,N_4115);
xnor U4273 (N_4273,N_4000,N_4163);
and U4274 (N_4274,N_4020,N_4126);
or U4275 (N_4275,N_4117,N_4077);
nand U4276 (N_4276,N_4179,N_4070);
and U4277 (N_4277,N_4098,N_4095);
or U4278 (N_4278,N_4091,N_4015);
nand U4279 (N_4279,N_4162,N_4042);
xnor U4280 (N_4280,N_4193,N_4022);
nor U4281 (N_4281,N_4138,N_4156);
nor U4282 (N_4282,N_4056,N_4151);
xor U4283 (N_4283,N_4139,N_4159);
xnor U4284 (N_4284,N_4002,N_4066);
nor U4285 (N_4285,N_4074,N_4121);
xor U4286 (N_4286,N_4063,N_4023);
and U4287 (N_4287,N_4075,N_4050);
or U4288 (N_4288,N_4032,N_4019);
or U4289 (N_4289,N_4064,N_4199);
and U4290 (N_4290,N_4107,N_4104);
xor U4291 (N_4291,N_4082,N_4191);
or U4292 (N_4292,N_4166,N_4033);
xor U4293 (N_4293,N_4118,N_4105);
nand U4294 (N_4294,N_4160,N_4001);
and U4295 (N_4295,N_4003,N_4040);
and U4296 (N_4296,N_4031,N_4181);
xnor U4297 (N_4297,N_4067,N_4125);
and U4298 (N_4298,N_4024,N_4025);
or U4299 (N_4299,N_4116,N_4145);
nand U4300 (N_4300,N_4188,N_4022);
and U4301 (N_4301,N_4148,N_4053);
xnor U4302 (N_4302,N_4169,N_4016);
xnor U4303 (N_4303,N_4088,N_4033);
or U4304 (N_4304,N_4139,N_4124);
and U4305 (N_4305,N_4070,N_4193);
and U4306 (N_4306,N_4015,N_4123);
or U4307 (N_4307,N_4086,N_4153);
and U4308 (N_4308,N_4041,N_4174);
and U4309 (N_4309,N_4118,N_4054);
or U4310 (N_4310,N_4143,N_4073);
xnor U4311 (N_4311,N_4077,N_4075);
xnor U4312 (N_4312,N_4079,N_4021);
or U4313 (N_4313,N_4022,N_4162);
nor U4314 (N_4314,N_4005,N_4197);
or U4315 (N_4315,N_4158,N_4174);
and U4316 (N_4316,N_4001,N_4098);
nand U4317 (N_4317,N_4198,N_4039);
or U4318 (N_4318,N_4102,N_4047);
nor U4319 (N_4319,N_4069,N_4112);
and U4320 (N_4320,N_4083,N_4122);
or U4321 (N_4321,N_4161,N_4146);
or U4322 (N_4322,N_4118,N_4057);
and U4323 (N_4323,N_4085,N_4084);
and U4324 (N_4324,N_4045,N_4075);
xor U4325 (N_4325,N_4029,N_4080);
nor U4326 (N_4326,N_4155,N_4185);
or U4327 (N_4327,N_4005,N_4027);
or U4328 (N_4328,N_4064,N_4087);
nor U4329 (N_4329,N_4173,N_4000);
or U4330 (N_4330,N_4070,N_4148);
xnor U4331 (N_4331,N_4086,N_4088);
and U4332 (N_4332,N_4079,N_4114);
or U4333 (N_4333,N_4103,N_4135);
or U4334 (N_4334,N_4028,N_4174);
and U4335 (N_4335,N_4118,N_4142);
or U4336 (N_4336,N_4105,N_4189);
nor U4337 (N_4337,N_4094,N_4102);
or U4338 (N_4338,N_4124,N_4197);
and U4339 (N_4339,N_4189,N_4010);
or U4340 (N_4340,N_4078,N_4096);
xor U4341 (N_4341,N_4165,N_4170);
nand U4342 (N_4342,N_4032,N_4000);
and U4343 (N_4343,N_4067,N_4007);
or U4344 (N_4344,N_4016,N_4066);
nor U4345 (N_4345,N_4024,N_4093);
nor U4346 (N_4346,N_4190,N_4025);
nor U4347 (N_4347,N_4074,N_4067);
and U4348 (N_4348,N_4051,N_4010);
nand U4349 (N_4349,N_4131,N_4081);
nand U4350 (N_4350,N_4054,N_4093);
xor U4351 (N_4351,N_4152,N_4088);
and U4352 (N_4352,N_4187,N_4129);
and U4353 (N_4353,N_4130,N_4009);
and U4354 (N_4354,N_4189,N_4004);
and U4355 (N_4355,N_4042,N_4019);
xnor U4356 (N_4356,N_4185,N_4057);
nand U4357 (N_4357,N_4124,N_4052);
xnor U4358 (N_4358,N_4056,N_4141);
nand U4359 (N_4359,N_4172,N_4012);
or U4360 (N_4360,N_4011,N_4010);
or U4361 (N_4361,N_4133,N_4023);
nor U4362 (N_4362,N_4165,N_4099);
nor U4363 (N_4363,N_4056,N_4135);
nand U4364 (N_4364,N_4157,N_4027);
nand U4365 (N_4365,N_4007,N_4003);
xor U4366 (N_4366,N_4123,N_4192);
xnor U4367 (N_4367,N_4065,N_4067);
nor U4368 (N_4368,N_4085,N_4088);
nand U4369 (N_4369,N_4186,N_4138);
or U4370 (N_4370,N_4112,N_4107);
or U4371 (N_4371,N_4167,N_4044);
xnor U4372 (N_4372,N_4128,N_4070);
xor U4373 (N_4373,N_4130,N_4123);
nand U4374 (N_4374,N_4079,N_4074);
nand U4375 (N_4375,N_4035,N_4021);
nand U4376 (N_4376,N_4136,N_4130);
xor U4377 (N_4377,N_4161,N_4073);
xor U4378 (N_4378,N_4152,N_4195);
nor U4379 (N_4379,N_4009,N_4131);
nor U4380 (N_4380,N_4168,N_4067);
xor U4381 (N_4381,N_4027,N_4181);
nor U4382 (N_4382,N_4075,N_4097);
nor U4383 (N_4383,N_4173,N_4085);
and U4384 (N_4384,N_4049,N_4032);
and U4385 (N_4385,N_4070,N_4037);
xnor U4386 (N_4386,N_4155,N_4174);
nor U4387 (N_4387,N_4160,N_4164);
or U4388 (N_4388,N_4063,N_4052);
or U4389 (N_4389,N_4126,N_4018);
and U4390 (N_4390,N_4183,N_4084);
or U4391 (N_4391,N_4196,N_4093);
or U4392 (N_4392,N_4011,N_4153);
xor U4393 (N_4393,N_4081,N_4154);
and U4394 (N_4394,N_4171,N_4101);
or U4395 (N_4395,N_4036,N_4091);
nand U4396 (N_4396,N_4153,N_4037);
and U4397 (N_4397,N_4095,N_4112);
or U4398 (N_4398,N_4069,N_4026);
nand U4399 (N_4399,N_4014,N_4044);
and U4400 (N_4400,N_4327,N_4319);
xnor U4401 (N_4401,N_4373,N_4372);
nand U4402 (N_4402,N_4320,N_4324);
and U4403 (N_4403,N_4386,N_4216);
xnor U4404 (N_4404,N_4358,N_4314);
nor U4405 (N_4405,N_4300,N_4361);
nor U4406 (N_4406,N_4304,N_4338);
xnor U4407 (N_4407,N_4379,N_4208);
or U4408 (N_4408,N_4253,N_4363);
nor U4409 (N_4409,N_4348,N_4387);
and U4410 (N_4410,N_4290,N_4238);
xnor U4411 (N_4411,N_4384,N_4281);
or U4412 (N_4412,N_4342,N_4241);
nor U4413 (N_4413,N_4318,N_4219);
and U4414 (N_4414,N_4370,N_4233);
and U4415 (N_4415,N_4225,N_4388);
xor U4416 (N_4416,N_4271,N_4261);
or U4417 (N_4417,N_4245,N_4280);
and U4418 (N_4418,N_4336,N_4200);
and U4419 (N_4419,N_4236,N_4207);
nand U4420 (N_4420,N_4391,N_4226);
xor U4421 (N_4421,N_4366,N_4390);
xnor U4422 (N_4422,N_4355,N_4210);
nand U4423 (N_4423,N_4299,N_4275);
or U4424 (N_4424,N_4228,N_4368);
or U4425 (N_4425,N_4301,N_4287);
and U4426 (N_4426,N_4240,N_4311);
and U4427 (N_4427,N_4352,N_4377);
and U4428 (N_4428,N_4214,N_4333);
xnor U4429 (N_4429,N_4360,N_4378);
nand U4430 (N_4430,N_4206,N_4375);
or U4431 (N_4431,N_4298,N_4376);
and U4432 (N_4432,N_4328,N_4211);
and U4433 (N_4433,N_4251,N_4380);
nand U4434 (N_4434,N_4204,N_4274);
xnor U4435 (N_4435,N_4269,N_4242);
nor U4436 (N_4436,N_4349,N_4317);
nand U4437 (N_4437,N_4227,N_4394);
nor U4438 (N_4438,N_4279,N_4247);
and U4439 (N_4439,N_4307,N_4288);
xor U4440 (N_4440,N_4398,N_4237);
or U4441 (N_4441,N_4230,N_4201);
and U4442 (N_4442,N_4213,N_4321);
xnor U4443 (N_4443,N_4256,N_4350);
nor U4444 (N_4444,N_4239,N_4343);
nor U4445 (N_4445,N_4273,N_4202);
nand U4446 (N_4446,N_4277,N_4334);
or U4447 (N_4447,N_4264,N_4395);
xnor U4448 (N_4448,N_4316,N_4203);
or U4449 (N_4449,N_4292,N_4313);
nor U4450 (N_4450,N_4362,N_4255);
or U4451 (N_4451,N_4351,N_4254);
nand U4452 (N_4452,N_4374,N_4340);
and U4453 (N_4453,N_4385,N_4346);
and U4454 (N_4454,N_4283,N_4244);
nand U4455 (N_4455,N_4399,N_4257);
nor U4456 (N_4456,N_4220,N_4235);
or U4457 (N_4457,N_4345,N_4393);
xnor U4458 (N_4458,N_4262,N_4278);
nor U4459 (N_4459,N_4310,N_4323);
or U4460 (N_4460,N_4364,N_4263);
or U4461 (N_4461,N_4260,N_4305);
xnor U4462 (N_4462,N_4356,N_4243);
and U4463 (N_4463,N_4381,N_4250);
and U4464 (N_4464,N_4291,N_4248);
and U4465 (N_4465,N_4282,N_4332);
xnor U4466 (N_4466,N_4331,N_4330);
or U4467 (N_4467,N_4205,N_4383);
nand U4468 (N_4468,N_4382,N_4272);
and U4469 (N_4469,N_4322,N_4258);
or U4470 (N_4470,N_4267,N_4252);
or U4471 (N_4471,N_4222,N_4285);
nor U4472 (N_4472,N_4371,N_4224);
or U4473 (N_4473,N_4265,N_4259);
nor U4474 (N_4474,N_4309,N_4329);
nand U4475 (N_4475,N_4359,N_4339);
xnor U4476 (N_4476,N_4396,N_4326);
nand U4477 (N_4477,N_4212,N_4229);
xor U4478 (N_4478,N_4308,N_4354);
or U4479 (N_4479,N_4303,N_4337);
or U4480 (N_4480,N_4234,N_4232);
and U4481 (N_4481,N_4268,N_4306);
and U4482 (N_4482,N_4286,N_4246);
and U4483 (N_4483,N_4344,N_4341);
and U4484 (N_4484,N_4249,N_4365);
or U4485 (N_4485,N_4335,N_4347);
or U4486 (N_4486,N_4221,N_4289);
or U4487 (N_4487,N_4218,N_4296);
xnor U4488 (N_4488,N_4397,N_4215);
or U4489 (N_4489,N_4270,N_4294);
or U4490 (N_4490,N_4315,N_4353);
xnor U4491 (N_4491,N_4297,N_4266);
nor U4492 (N_4492,N_4223,N_4293);
nor U4493 (N_4493,N_4389,N_4209);
and U4494 (N_4494,N_4367,N_4276);
nor U4495 (N_4495,N_4302,N_4312);
and U4496 (N_4496,N_4325,N_4231);
nor U4497 (N_4497,N_4369,N_4357);
nand U4498 (N_4498,N_4284,N_4392);
and U4499 (N_4499,N_4295,N_4217);
xor U4500 (N_4500,N_4387,N_4371);
nand U4501 (N_4501,N_4302,N_4320);
nand U4502 (N_4502,N_4344,N_4387);
xor U4503 (N_4503,N_4381,N_4232);
nand U4504 (N_4504,N_4353,N_4348);
xnor U4505 (N_4505,N_4347,N_4202);
nor U4506 (N_4506,N_4251,N_4360);
xnor U4507 (N_4507,N_4294,N_4214);
nor U4508 (N_4508,N_4331,N_4328);
or U4509 (N_4509,N_4281,N_4235);
and U4510 (N_4510,N_4392,N_4370);
nand U4511 (N_4511,N_4278,N_4313);
and U4512 (N_4512,N_4387,N_4242);
xor U4513 (N_4513,N_4323,N_4362);
xnor U4514 (N_4514,N_4285,N_4214);
xnor U4515 (N_4515,N_4376,N_4358);
nor U4516 (N_4516,N_4396,N_4358);
xnor U4517 (N_4517,N_4279,N_4317);
xnor U4518 (N_4518,N_4319,N_4328);
nor U4519 (N_4519,N_4377,N_4292);
and U4520 (N_4520,N_4207,N_4204);
nor U4521 (N_4521,N_4364,N_4233);
nand U4522 (N_4522,N_4399,N_4206);
nand U4523 (N_4523,N_4357,N_4307);
nand U4524 (N_4524,N_4337,N_4271);
nor U4525 (N_4525,N_4345,N_4285);
or U4526 (N_4526,N_4274,N_4280);
nor U4527 (N_4527,N_4236,N_4348);
nand U4528 (N_4528,N_4223,N_4388);
and U4529 (N_4529,N_4268,N_4325);
nor U4530 (N_4530,N_4244,N_4344);
or U4531 (N_4531,N_4260,N_4384);
xor U4532 (N_4532,N_4227,N_4383);
and U4533 (N_4533,N_4280,N_4368);
or U4534 (N_4534,N_4391,N_4250);
or U4535 (N_4535,N_4326,N_4342);
nor U4536 (N_4536,N_4276,N_4294);
xor U4537 (N_4537,N_4202,N_4339);
or U4538 (N_4538,N_4331,N_4217);
and U4539 (N_4539,N_4293,N_4338);
nand U4540 (N_4540,N_4306,N_4230);
or U4541 (N_4541,N_4362,N_4213);
xnor U4542 (N_4542,N_4369,N_4354);
xor U4543 (N_4543,N_4290,N_4320);
or U4544 (N_4544,N_4313,N_4231);
nor U4545 (N_4545,N_4384,N_4309);
xnor U4546 (N_4546,N_4224,N_4357);
nand U4547 (N_4547,N_4383,N_4250);
nand U4548 (N_4548,N_4338,N_4350);
nand U4549 (N_4549,N_4224,N_4205);
and U4550 (N_4550,N_4291,N_4202);
and U4551 (N_4551,N_4275,N_4294);
or U4552 (N_4552,N_4394,N_4267);
and U4553 (N_4553,N_4360,N_4223);
xor U4554 (N_4554,N_4293,N_4397);
and U4555 (N_4555,N_4397,N_4315);
or U4556 (N_4556,N_4230,N_4359);
or U4557 (N_4557,N_4337,N_4296);
or U4558 (N_4558,N_4231,N_4349);
and U4559 (N_4559,N_4204,N_4272);
xnor U4560 (N_4560,N_4320,N_4304);
xor U4561 (N_4561,N_4287,N_4312);
and U4562 (N_4562,N_4205,N_4316);
nor U4563 (N_4563,N_4306,N_4293);
or U4564 (N_4564,N_4246,N_4205);
and U4565 (N_4565,N_4347,N_4281);
or U4566 (N_4566,N_4334,N_4308);
xor U4567 (N_4567,N_4200,N_4332);
or U4568 (N_4568,N_4261,N_4311);
and U4569 (N_4569,N_4320,N_4205);
xnor U4570 (N_4570,N_4361,N_4340);
nor U4571 (N_4571,N_4398,N_4233);
and U4572 (N_4572,N_4388,N_4292);
nand U4573 (N_4573,N_4326,N_4329);
and U4574 (N_4574,N_4330,N_4221);
xor U4575 (N_4575,N_4302,N_4366);
and U4576 (N_4576,N_4243,N_4321);
xnor U4577 (N_4577,N_4268,N_4320);
nand U4578 (N_4578,N_4217,N_4385);
nor U4579 (N_4579,N_4299,N_4298);
nor U4580 (N_4580,N_4386,N_4323);
and U4581 (N_4581,N_4272,N_4280);
and U4582 (N_4582,N_4226,N_4296);
nand U4583 (N_4583,N_4242,N_4265);
xor U4584 (N_4584,N_4245,N_4348);
nand U4585 (N_4585,N_4379,N_4253);
nor U4586 (N_4586,N_4388,N_4233);
nor U4587 (N_4587,N_4220,N_4369);
or U4588 (N_4588,N_4218,N_4369);
nand U4589 (N_4589,N_4325,N_4365);
and U4590 (N_4590,N_4258,N_4349);
nor U4591 (N_4591,N_4367,N_4252);
nand U4592 (N_4592,N_4291,N_4236);
nor U4593 (N_4593,N_4244,N_4250);
or U4594 (N_4594,N_4283,N_4356);
and U4595 (N_4595,N_4209,N_4375);
and U4596 (N_4596,N_4249,N_4306);
xnor U4597 (N_4597,N_4378,N_4366);
or U4598 (N_4598,N_4305,N_4399);
or U4599 (N_4599,N_4381,N_4224);
nand U4600 (N_4600,N_4466,N_4491);
and U4601 (N_4601,N_4500,N_4483);
nor U4602 (N_4602,N_4493,N_4574);
or U4603 (N_4603,N_4460,N_4552);
and U4604 (N_4604,N_4584,N_4557);
xnor U4605 (N_4605,N_4496,N_4568);
or U4606 (N_4606,N_4450,N_4418);
or U4607 (N_4607,N_4564,N_4504);
and U4608 (N_4608,N_4407,N_4549);
and U4609 (N_4609,N_4521,N_4404);
xor U4610 (N_4610,N_4461,N_4526);
nand U4611 (N_4611,N_4561,N_4555);
and U4612 (N_4612,N_4513,N_4475);
nand U4613 (N_4613,N_4484,N_4425);
and U4614 (N_4614,N_4575,N_4565);
nand U4615 (N_4615,N_4591,N_4492);
and U4616 (N_4616,N_4485,N_4436);
nand U4617 (N_4617,N_4514,N_4502);
and U4618 (N_4618,N_4452,N_4536);
xor U4619 (N_4619,N_4416,N_4426);
nand U4620 (N_4620,N_4590,N_4563);
nand U4621 (N_4621,N_4402,N_4499);
and U4622 (N_4622,N_4451,N_4419);
xnor U4623 (N_4623,N_4579,N_4535);
nand U4624 (N_4624,N_4468,N_4510);
nor U4625 (N_4625,N_4413,N_4596);
and U4626 (N_4626,N_4415,N_4540);
or U4627 (N_4627,N_4453,N_4562);
and U4628 (N_4628,N_4589,N_4520);
and U4629 (N_4629,N_4403,N_4550);
or U4630 (N_4630,N_4423,N_4541);
nand U4631 (N_4631,N_4581,N_4479);
or U4632 (N_4632,N_4515,N_4480);
nand U4633 (N_4633,N_4446,N_4495);
or U4634 (N_4634,N_4440,N_4482);
nand U4635 (N_4635,N_4434,N_4471);
nand U4636 (N_4636,N_4501,N_4455);
xnor U4637 (N_4637,N_4454,N_4572);
nand U4638 (N_4638,N_4459,N_4544);
and U4639 (N_4639,N_4509,N_4511);
nand U4640 (N_4640,N_4410,N_4437);
nor U4641 (N_4641,N_4585,N_4472);
nand U4642 (N_4642,N_4580,N_4477);
and U4643 (N_4643,N_4538,N_4583);
nor U4644 (N_4644,N_4570,N_4527);
nor U4645 (N_4645,N_4431,N_4530);
nand U4646 (N_4646,N_4448,N_4532);
xnor U4647 (N_4647,N_4476,N_4473);
nand U4648 (N_4648,N_4597,N_4512);
xnor U4649 (N_4649,N_4421,N_4539);
or U4650 (N_4650,N_4588,N_4551);
and U4651 (N_4651,N_4443,N_4505);
nor U4652 (N_4652,N_4592,N_4508);
xor U4653 (N_4653,N_4432,N_4556);
nand U4654 (N_4654,N_4518,N_4409);
or U4655 (N_4655,N_4598,N_4430);
nand U4656 (N_4656,N_4469,N_4488);
or U4657 (N_4657,N_4465,N_4533);
or U4658 (N_4658,N_4490,N_4582);
nand U4659 (N_4659,N_4559,N_4449);
and U4660 (N_4660,N_4467,N_4522);
nand U4661 (N_4661,N_4444,N_4534);
and U4662 (N_4662,N_4558,N_4464);
nor U4663 (N_4663,N_4517,N_4438);
nor U4664 (N_4664,N_4531,N_4422);
xor U4665 (N_4665,N_4401,N_4528);
or U4666 (N_4666,N_4560,N_4458);
and U4667 (N_4667,N_4546,N_4573);
xor U4668 (N_4668,N_4547,N_4577);
and U4669 (N_4669,N_4529,N_4524);
xnor U4670 (N_4670,N_4487,N_4507);
nand U4671 (N_4671,N_4542,N_4506);
or U4672 (N_4672,N_4554,N_4519);
xor U4673 (N_4673,N_4587,N_4481);
xnor U4674 (N_4674,N_4435,N_4489);
nor U4675 (N_4675,N_4523,N_4586);
nor U4676 (N_4676,N_4411,N_4553);
nand U4677 (N_4677,N_4442,N_4408);
xor U4678 (N_4678,N_4445,N_4548);
or U4679 (N_4679,N_4447,N_4594);
or U4680 (N_4680,N_4595,N_4545);
or U4681 (N_4681,N_4433,N_4417);
or U4682 (N_4682,N_4576,N_4566);
and U4683 (N_4683,N_4457,N_4414);
or U4684 (N_4684,N_4486,N_4494);
xor U4685 (N_4685,N_4478,N_4427);
nand U4686 (N_4686,N_4599,N_4516);
or U4687 (N_4687,N_4569,N_4578);
and U4688 (N_4688,N_4429,N_4543);
and U4689 (N_4689,N_4412,N_4405);
and U4690 (N_4690,N_4537,N_4497);
and U4691 (N_4691,N_4593,N_4441);
nor U4692 (N_4692,N_4420,N_4470);
and U4693 (N_4693,N_4424,N_4525);
xnor U4694 (N_4694,N_4463,N_4571);
xor U4695 (N_4695,N_4406,N_4439);
or U4696 (N_4696,N_4474,N_4428);
nor U4697 (N_4697,N_4498,N_4462);
xor U4698 (N_4698,N_4503,N_4456);
nand U4699 (N_4699,N_4567,N_4400);
or U4700 (N_4700,N_4593,N_4428);
nor U4701 (N_4701,N_4423,N_4485);
and U4702 (N_4702,N_4419,N_4454);
or U4703 (N_4703,N_4484,N_4513);
nor U4704 (N_4704,N_4504,N_4496);
xor U4705 (N_4705,N_4581,N_4538);
nand U4706 (N_4706,N_4445,N_4523);
nand U4707 (N_4707,N_4584,N_4435);
nand U4708 (N_4708,N_4457,N_4460);
and U4709 (N_4709,N_4589,N_4532);
or U4710 (N_4710,N_4530,N_4519);
nand U4711 (N_4711,N_4547,N_4514);
and U4712 (N_4712,N_4525,N_4471);
or U4713 (N_4713,N_4456,N_4468);
and U4714 (N_4714,N_4563,N_4581);
or U4715 (N_4715,N_4414,N_4596);
nand U4716 (N_4716,N_4558,N_4415);
or U4717 (N_4717,N_4492,N_4507);
xor U4718 (N_4718,N_4493,N_4478);
nor U4719 (N_4719,N_4425,N_4426);
or U4720 (N_4720,N_4592,N_4511);
and U4721 (N_4721,N_4404,N_4402);
nor U4722 (N_4722,N_4590,N_4513);
and U4723 (N_4723,N_4452,N_4586);
or U4724 (N_4724,N_4538,N_4486);
nor U4725 (N_4725,N_4452,N_4512);
and U4726 (N_4726,N_4408,N_4506);
nand U4727 (N_4727,N_4509,N_4598);
or U4728 (N_4728,N_4481,N_4436);
and U4729 (N_4729,N_4450,N_4540);
and U4730 (N_4730,N_4527,N_4489);
nand U4731 (N_4731,N_4426,N_4541);
nor U4732 (N_4732,N_4527,N_4574);
nand U4733 (N_4733,N_4458,N_4486);
or U4734 (N_4734,N_4522,N_4499);
nand U4735 (N_4735,N_4410,N_4454);
or U4736 (N_4736,N_4497,N_4454);
xor U4737 (N_4737,N_4539,N_4427);
nand U4738 (N_4738,N_4416,N_4440);
or U4739 (N_4739,N_4415,N_4445);
xor U4740 (N_4740,N_4599,N_4505);
nor U4741 (N_4741,N_4455,N_4540);
xnor U4742 (N_4742,N_4518,N_4510);
nor U4743 (N_4743,N_4521,N_4409);
nor U4744 (N_4744,N_4485,N_4448);
nand U4745 (N_4745,N_4580,N_4577);
xor U4746 (N_4746,N_4478,N_4443);
and U4747 (N_4747,N_4551,N_4499);
or U4748 (N_4748,N_4556,N_4439);
and U4749 (N_4749,N_4566,N_4509);
nand U4750 (N_4750,N_4580,N_4403);
or U4751 (N_4751,N_4501,N_4461);
nand U4752 (N_4752,N_4599,N_4423);
nor U4753 (N_4753,N_4485,N_4527);
and U4754 (N_4754,N_4522,N_4454);
or U4755 (N_4755,N_4546,N_4589);
or U4756 (N_4756,N_4568,N_4466);
or U4757 (N_4757,N_4523,N_4561);
nor U4758 (N_4758,N_4521,N_4509);
and U4759 (N_4759,N_4406,N_4461);
nor U4760 (N_4760,N_4484,N_4524);
and U4761 (N_4761,N_4516,N_4464);
xnor U4762 (N_4762,N_4571,N_4586);
nand U4763 (N_4763,N_4591,N_4461);
xnor U4764 (N_4764,N_4542,N_4487);
xor U4765 (N_4765,N_4448,N_4533);
or U4766 (N_4766,N_4475,N_4479);
nand U4767 (N_4767,N_4546,N_4489);
nor U4768 (N_4768,N_4535,N_4470);
xnor U4769 (N_4769,N_4431,N_4430);
nor U4770 (N_4770,N_4511,N_4494);
nor U4771 (N_4771,N_4569,N_4464);
nand U4772 (N_4772,N_4571,N_4563);
xnor U4773 (N_4773,N_4416,N_4531);
or U4774 (N_4774,N_4438,N_4542);
nor U4775 (N_4775,N_4539,N_4473);
and U4776 (N_4776,N_4529,N_4499);
or U4777 (N_4777,N_4464,N_4404);
xor U4778 (N_4778,N_4462,N_4527);
or U4779 (N_4779,N_4570,N_4469);
nor U4780 (N_4780,N_4584,N_4580);
or U4781 (N_4781,N_4594,N_4530);
and U4782 (N_4782,N_4552,N_4535);
or U4783 (N_4783,N_4585,N_4549);
nor U4784 (N_4784,N_4576,N_4431);
or U4785 (N_4785,N_4484,N_4518);
nand U4786 (N_4786,N_4487,N_4552);
and U4787 (N_4787,N_4588,N_4486);
xor U4788 (N_4788,N_4500,N_4436);
and U4789 (N_4789,N_4557,N_4425);
nor U4790 (N_4790,N_4529,N_4541);
nor U4791 (N_4791,N_4507,N_4498);
or U4792 (N_4792,N_4564,N_4422);
and U4793 (N_4793,N_4402,N_4514);
nor U4794 (N_4794,N_4459,N_4565);
nand U4795 (N_4795,N_4551,N_4556);
or U4796 (N_4796,N_4570,N_4420);
and U4797 (N_4797,N_4461,N_4454);
nor U4798 (N_4798,N_4579,N_4518);
or U4799 (N_4799,N_4407,N_4431);
xor U4800 (N_4800,N_4739,N_4689);
nand U4801 (N_4801,N_4737,N_4633);
and U4802 (N_4802,N_4743,N_4614);
nor U4803 (N_4803,N_4666,N_4612);
nand U4804 (N_4804,N_4618,N_4728);
xor U4805 (N_4805,N_4616,N_4690);
nand U4806 (N_4806,N_4695,N_4701);
or U4807 (N_4807,N_4747,N_4613);
or U4808 (N_4808,N_4762,N_4651);
nand U4809 (N_4809,N_4640,N_4604);
xnor U4810 (N_4810,N_4745,N_4776);
and U4811 (N_4811,N_4630,N_4669);
nor U4812 (N_4812,N_4731,N_4746);
xor U4813 (N_4813,N_4719,N_4729);
xnor U4814 (N_4814,N_4702,N_4742);
nor U4815 (N_4815,N_4645,N_4672);
and U4816 (N_4816,N_4647,N_4621);
nand U4817 (N_4817,N_4727,N_4697);
nor U4818 (N_4818,N_4781,N_4664);
or U4819 (N_4819,N_4696,N_4632);
or U4820 (N_4820,N_4755,N_4658);
or U4821 (N_4821,N_4744,N_4656);
or U4822 (N_4822,N_4740,N_4706);
nor U4823 (N_4823,N_4748,N_4665);
nand U4824 (N_4824,N_4767,N_4676);
nor U4825 (N_4825,N_4620,N_4721);
nor U4826 (N_4826,N_4628,N_4793);
or U4827 (N_4827,N_4798,N_4684);
xor U4828 (N_4828,N_4723,N_4714);
nand U4829 (N_4829,N_4769,N_4765);
and U4830 (N_4830,N_4735,N_4787);
or U4831 (N_4831,N_4734,N_4631);
nand U4832 (N_4832,N_4759,N_4786);
nand U4833 (N_4833,N_4603,N_4763);
or U4834 (N_4834,N_4681,N_4653);
xor U4835 (N_4835,N_4758,N_4705);
nand U4836 (N_4836,N_4779,N_4682);
xor U4837 (N_4837,N_4717,N_4650);
nand U4838 (N_4838,N_4615,N_4789);
nand U4839 (N_4839,N_4785,N_4674);
nand U4840 (N_4840,N_4623,N_4625);
and U4841 (N_4841,N_4764,N_4766);
nand U4842 (N_4842,N_4636,N_4677);
nor U4843 (N_4843,N_4709,N_4652);
nand U4844 (N_4844,N_4605,N_4713);
and U4845 (N_4845,N_4638,N_4661);
and U4846 (N_4846,N_4718,N_4752);
nor U4847 (N_4847,N_4768,N_4733);
xor U4848 (N_4848,N_4724,N_4777);
or U4849 (N_4849,N_4760,N_4627);
nand U4850 (N_4850,N_4704,N_4626);
nor U4851 (N_4851,N_4753,N_4601);
nor U4852 (N_4852,N_4700,N_4655);
or U4853 (N_4853,N_4757,N_4639);
and U4854 (N_4854,N_4607,N_4606);
xor U4855 (N_4855,N_4698,N_4751);
nor U4856 (N_4856,N_4750,N_4642);
xor U4857 (N_4857,N_4790,N_4778);
or U4858 (N_4858,N_4610,N_4678);
nand U4859 (N_4859,N_4619,N_4683);
xnor U4860 (N_4860,N_4722,N_4673);
or U4861 (N_4861,N_4761,N_4611);
nand U4862 (N_4862,N_4663,N_4668);
or U4863 (N_4863,N_4791,N_4707);
or U4864 (N_4864,N_4657,N_4715);
nor U4865 (N_4865,N_4725,N_4608);
nor U4866 (N_4866,N_4736,N_4774);
and U4867 (N_4867,N_4726,N_4772);
xnor U4868 (N_4868,N_4662,N_4659);
nor U4869 (N_4869,N_4686,N_4644);
and U4870 (N_4870,N_4679,N_4670);
and U4871 (N_4871,N_4784,N_4716);
nor U4872 (N_4872,N_4691,N_4720);
nand U4873 (N_4873,N_4643,N_4730);
nor U4874 (N_4874,N_4799,N_4741);
or U4875 (N_4875,N_4671,N_4756);
nor U4876 (N_4876,N_4749,N_4710);
nand U4877 (N_4877,N_4667,N_4600);
xor U4878 (N_4878,N_4792,N_4635);
nor U4879 (N_4879,N_4685,N_4629);
and U4880 (N_4880,N_4770,N_4732);
or U4881 (N_4881,N_4637,N_4648);
and U4882 (N_4882,N_4622,N_4675);
and U4883 (N_4883,N_4609,N_4646);
nor U4884 (N_4884,N_4694,N_4680);
xor U4885 (N_4885,N_4738,N_4771);
and U4886 (N_4886,N_4692,N_4624);
nor U4887 (N_4887,N_4688,N_4649);
nand U4888 (N_4888,N_4783,N_4660);
nand U4889 (N_4889,N_4693,N_4711);
or U4890 (N_4890,N_4773,N_4654);
nand U4891 (N_4891,N_4634,N_4602);
xor U4892 (N_4892,N_4703,N_4788);
and U4893 (N_4893,N_4782,N_4797);
xnor U4894 (N_4894,N_4712,N_4699);
or U4895 (N_4895,N_4794,N_4775);
nand U4896 (N_4896,N_4754,N_4796);
xor U4897 (N_4897,N_4687,N_4780);
nand U4898 (N_4898,N_4617,N_4708);
xnor U4899 (N_4899,N_4795,N_4641);
or U4900 (N_4900,N_4695,N_4673);
or U4901 (N_4901,N_4702,N_4754);
xor U4902 (N_4902,N_4636,N_4687);
nand U4903 (N_4903,N_4604,N_4745);
xnor U4904 (N_4904,N_4729,N_4618);
xor U4905 (N_4905,N_4701,N_4768);
nor U4906 (N_4906,N_4621,N_4603);
or U4907 (N_4907,N_4736,N_4669);
nand U4908 (N_4908,N_4676,N_4746);
and U4909 (N_4909,N_4738,N_4765);
nand U4910 (N_4910,N_4643,N_4750);
nand U4911 (N_4911,N_4746,N_4789);
xor U4912 (N_4912,N_4638,N_4622);
nand U4913 (N_4913,N_4746,N_4691);
and U4914 (N_4914,N_4712,N_4697);
nand U4915 (N_4915,N_4764,N_4703);
nor U4916 (N_4916,N_4637,N_4652);
nand U4917 (N_4917,N_4772,N_4771);
or U4918 (N_4918,N_4708,N_4663);
nand U4919 (N_4919,N_4646,N_4739);
nor U4920 (N_4920,N_4662,N_4665);
xor U4921 (N_4921,N_4746,N_4709);
xor U4922 (N_4922,N_4733,N_4648);
nor U4923 (N_4923,N_4774,N_4787);
nor U4924 (N_4924,N_4663,N_4677);
nor U4925 (N_4925,N_4600,N_4773);
xor U4926 (N_4926,N_4602,N_4798);
and U4927 (N_4927,N_4609,N_4614);
nand U4928 (N_4928,N_4707,N_4625);
and U4929 (N_4929,N_4721,N_4683);
and U4930 (N_4930,N_4672,N_4680);
nand U4931 (N_4931,N_4620,N_4739);
xor U4932 (N_4932,N_4613,N_4729);
nor U4933 (N_4933,N_4776,N_4652);
nor U4934 (N_4934,N_4604,N_4775);
nand U4935 (N_4935,N_4798,N_4703);
nor U4936 (N_4936,N_4787,N_4605);
nand U4937 (N_4937,N_4741,N_4714);
nand U4938 (N_4938,N_4684,N_4693);
nand U4939 (N_4939,N_4718,N_4627);
nor U4940 (N_4940,N_4770,N_4665);
and U4941 (N_4941,N_4671,N_4610);
or U4942 (N_4942,N_4688,N_4670);
or U4943 (N_4943,N_4735,N_4607);
nor U4944 (N_4944,N_4783,N_4641);
xor U4945 (N_4945,N_4618,N_4745);
nand U4946 (N_4946,N_4651,N_4771);
or U4947 (N_4947,N_4722,N_4751);
xnor U4948 (N_4948,N_4719,N_4661);
nor U4949 (N_4949,N_4799,N_4657);
or U4950 (N_4950,N_4696,N_4699);
nand U4951 (N_4951,N_4695,N_4697);
and U4952 (N_4952,N_4684,N_4767);
and U4953 (N_4953,N_4669,N_4685);
or U4954 (N_4954,N_4768,N_4647);
nand U4955 (N_4955,N_4623,N_4731);
xor U4956 (N_4956,N_4644,N_4648);
nand U4957 (N_4957,N_4778,N_4758);
or U4958 (N_4958,N_4734,N_4629);
nor U4959 (N_4959,N_4600,N_4767);
or U4960 (N_4960,N_4753,N_4661);
or U4961 (N_4961,N_4702,N_4688);
xor U4962 (N_4962,N_4631,N_4616);
nor U4963 (N_4963,N_4662,N_4748);
or U4964 (N_4964,N_4721,N_4612);
nor U4965 (N_4965,N_4757,N_4610);
xnor U4966 (N_4966,N_4699,N_4759);
nor U4967 (N_4967,N_4611,N_4743);
xor U4968 (N_4968,N_4680,N_4688);
nand U4969 (N_4969,N_4657,N_4679);
nor U4970 (N_4970,N_4626,N_4605);
or U4971 (N_4971,N_4638,N_4635);
and U4972 (N_4972,N_4798,N_4749);
and U4973 (N_4973,N_4742,N_4733);
or U4974 (N_4974,N_4799,N_4766);
nor U4975 (N_4975,N_4726,N_4671);
or U4976 (N_4976,N_4690,N_4753);
nand U4977 (N_4977,N_4668,N_4788);
nand U4978 (N_4978,N_4676,N_4604);
nor U4979 (N_4979,N_4679,N_4691);
xnor U4980 (N_4980,N_4723,N_4765);
and U4981 (N_4981,N_4632,N_4672);
nand U4982 (N_4982,N_4761,N_4740);
or U4983 (N_4983,N_4733,N_4672);
xor U4984 (N_4984,N_4757,N_4713);
nor U4985 (N_4985,N_4762,N_4702);
xor U4986 (N_4986,N_4748,N_4692);
xor U4987 (N_4987,N_4643,N_4646);
nand U4988 (N_4988,N_4669,N_4697);
nand U4989 (N_4989,N_4670,N_4637);
nand U4990 (N_4990,N_4798,N_4645);
nor U4991 (N_4991,N_4620,N_4799);
xnor U4992 (N_4992,N_4777,N_4774);
and U4993 (N_4993,N_4722,N_4689);
nand U4994 (N_4994,N_4722,N_4766);
and U4995 (N_4995,N_4614,N_4764);
or U4996 (N_4996,N_4691,N_4718);
nand U4997 (N_4997,N_4726,N_4633);
nand U4998 (N_4998,N_4737,N_4686);
nor U4999 (N_4999,N_4784,N_4636);
xor U5000 (N_5000,N_4850,N_4803);
nand U5001 (N_5001,N_4848,N_4926);
nor U5002 (N_5002,N_4822,N_4895);
xor U5003 (N_5003,N_4900,N_4819);
nand U5004 (N_5004,N_4947,N_4905);
nand U5005 (N_5005,N_4815,N_4966);
xnor U5006 (N_5006,N_4944,N_4861);
or U5007 (N_5007,N_4888,N_4984);
nor U5008 (N_5008,N_4825,N_4960);
and U5009 (N_5009,N_4835,N_4832);
or U5010 (N_5010,N_4979,N_4989);
and U5011 (N_5011,N_4934,N_4853);
and U5012 (N_5012,N_4912,N_4950);
nand U5013 (N_5013,N_4965,N_4981);
nand U5014 (N_5014,N_4964,N_4869);
or U5015 (N_5015,N_4897,N_4937);
or U5016 (N_5016,N_4930,N_4999);
nor U5017 (N_5017,N_4921,N_4866);
xnor U5018 (N_5018,N_4831,N_4923);
nor U5019 (N_5019,N_4914,N_4892);
or U5020 (N_5020,N_4891,N_4806);
nand U5021 (N_5021,N_4863,N_4844);
nand U5022 (N_5022,N_4980,N_4843);
nand U5023 (N_5023,N_4906,N_4849);
xor U5024 (N_5024,N_4994,N_4973);
nand U5025 (N_5025,N_4882,N_4887);
nor U5026 (N_5026,N_4865,N_4876);
nand U5027 (N_5027,N_4904,N_4935);
xor U5028 (N_5028,N_4933,N_4817);
xor U5029 (N_5029,N_4983,N_4818);
nor U5030 (N_5030,N_4855,N_4948);
nand U5031 (N_5031,N_4873,N_4883);
nand U5032 (N_5032,N_4884,N_4936);
and U5033 (N_5033,N_4801,N_4992);
nor U5034 (N_5034,N_4864,N_4868);
xnor U5035 (N_5035,N_4889,N_4991);
and U5036 (N_5036,N_4945,N_4995);
and U5037 (N_5037,N_4862,N_4978);
or U5038 (N_5038,N_4919,N_4880);
and U5039 (N_5039,N_4929,N_4931);
nor U5040 (N_5040,N_4872,N_4971);
and U5041 (N_5041,N_4968,N_4913);
nor U5042 (N_5042,N_4928,N_4998);
xnor U5043 (N_5043,N_4974,N_4941);
and U5044 (N_5044,N_4939,N_4837);
xor U5045 (N_5045,N_4820,N_4894);
xnor U5046 (N_5046,N_4854,N_4976);
xnor U5047 (N_5047,N_4836,N_4823);
nand U5048 (N_5048,N_4953,N_4970);
nand U5049 (N_5049,N_4902,N_4841);
nor U5050 (N_5050,N_4956,N_4826);
nand U5051 (N_5051,N_4938,N_4969);
and U5052 (N_5052,N_4916,N_4903);
nor U5053 (N_5053,N_4932,N_4918);
xor U5054 (N_5054,N_4893,N_4949);
or U5055 (N_5055,N_4975,N_4952);
xor U5056 (N_5056,N_4990,N_4845);
and U5057 (N_5057,N_4927,N_4804);
or U5058 (N_5058,N_4814,N_4901);
or U5059 (N_5059,N_4986,N_4871);
or U5060 (N_5060,N_4915,N_4886);
xnor U5061 (N_5061,N_4924,N_4957);
and U5062 (N_5062,N_4821,N_4907);
and U5063 (N_5063,N_4811,N_4896);
or U5064 (N_5064,N_4908,N_4852);
nor U5065 (N_5065,N_4961,N_4812);
xnor U5066 (N_5066,N_4885,N_4920);
and U5067 (N_5067,N_4910,N_4824);
nand U5068 (N_5068,N_4959,N_4878);
nand U5069 (N_5069,N_4859,N_4898);
or U5070 (N_5070,N_4899,N_4828);
xnor U5071 (N_5071,N_4972,N_4827);
and U5072 (N_5072,N_4997,N_4958);
nor U5073 (N_5073,N_4911,N_4955);
and U5074 (N_5074,N_4943,N_4881);
nand U5075 (N_5075,N_4963,N_4829);
nand U5076 (N_5076,N_4860,N_4802);
and U5077 (N_5077,N_4890,N_4813);
and U5078 (N_5078,N_4838,N_4816);
xnor U5079 (N_5079,N_4842,N_4851);
or U5080 (N_5080,N_4810,N_4830);
or U5081 (N_5081,N_4856,N_4996);
nor U5082 (N_5082,N_4846,N_4807);
and U5083 (N_5083,N_4839,N_4870);
or U5084 (N_5084,N_4833,N_4909);
nor U5085 (N_5085,N_4993,N_4925);
and U5086 (N_5086,N_4917,N_4942);
or U5087 (N_5087,N_4987,N_4867);
nor U5088 (N_5088,N_4946,N_4847);
nand U5089 (N_5089,N_4922,N_4877);
or U5090 (N_5090,N_4875,N_4834);
nor U5091 (N_5091,N_4954,N_4857);
nand U5092 (N_5092,N_4951,N_4874);
nor U5093 (N_5093,N_4858,N_4879);
or U5094 (N_5094,N_4967,N_4977);
or U5095 (N_5095,N_4805,N_4985);
xnor U5096 (N_5096,N_4808,N_4940);
nand U5097 (N_5097,N_4962,N_4809);
nand U5098 (N_5098,N_4800,N_4840);
xnor U5099 (N_5099,N_4988,N_4982);
nor U5100 (N_5100,N_4800,N_4950);
xnor U5101 (N_5101,N_4806,N_4956);
or U5102 (N_5102,N_4841,N_4982);
and U5103 (N_5103,N_4876,N_4945);
or U5104 (N_5104,N_4964,N_4933);
or U5105 (N_5105,N_4956,N_4822);
nand U5106 (N_5106,N_4996,N_4962);
and U5107 (N_5107,N_4961,N_4932);
nor U5108 (N_5108,N_4886,N_4935);
nor U5109 (N_5109,N_4980,N_4939);
or U5110 (N_5110,N_4900,N_4944);
nor U5111 (N_5111,N_4888,N_4865);
nor U5112 (N_5112,N_4951,N_4868);
xor U5113 (N_5113,N_4908,N_4925);
or U5114 (N_5114,N_4965,N_4984);
or U5115 (N_5115,N_4930,N_4914);
or U5116 (N_5116,N_4977,N_4830);
xnor U5117 (N_5117,N_4824,N_4825);
and U5118 (N_5118,N_4977,N_4864);
xnor U5119 (N_5119,N_4888,N_4843);
nand U5120 (N_5120,N_4805,N_4840);
and U5121 (N_5121,N_4968,N_4859);
nand U5122 (N_5122,N_4922,N_4973);
or U5123 (N_5123,N_4971,N_4926);
nor U5124 (N_5124,N_4854,N_4931);
nor U5125 (N_5125,N_4991,N_4925);
nor U5126 (N_5126,N_4958,N_4846);
and U5127 (N_5127,N_4990,N_4911);
nand U5128 (N_5128,N_4951,N_4883);
nor U5129 (N_5129,N_4870,N_4807);
or U5130 (N_5130,N_4814,N_4982);
and U5131 (N_5131,N_4813,N_4917);
nand U5132 (N_5132,N_4893,N_4975);
nand U5133 (N_5133,N_4862,N_4831);
xnor U5134 (N_5134,N_4937,N_4831);
xnor U5135 (N_5135,N_4870,N_4973);
or U5136 (N_5136,N_4957,N_4969);
nand U5137 (N_5137,N_4990,N_4853);
xor U5138 (N_5138,N_4897,N_4813);
or U5139 (N_5139,N_4909,N_4952);
or U5140 (N_5140,N_4902,N_4931);
and U5141 (N_5141,N_4805,N_4800);
and U5142 (N_5142,N_4935,N_4916);
nand U5143 (N_5143,N_4829,N_4955);
or U5144 (N_5144,N_4873,N_4899);
xnor U5145 (N_5145,N_4860,N_4826);
nand U5146 (N_5146,N_4850,N_4950);
nor U5147 (N_5147,N_4880,N_4955);
xor U5148 (N_5148,N_4872,N_4909);
xor U5149 (N_5149,N_4972,N_4970);
nand U5150 (N_5150,N_4922,N_4930);
or U5151 (N_5151,N_4815,N_4859);
nor U5152 (N_5152,N_4943,N_4986);
nor U5153 (N_5153,N_4925,N_4870);
or U5154 (N_5154,N_4994,N_4990);
nand U5155 (N_5155,N_4970,N_4887);
nor U5156 (N_5156,N_4805,N_4831);
xnor U5157 (N_5157,N_4831,N_4857);
and U5158 (N_5158,N_4934,N_4903);
nand U5159 (N_5159,N_4838,N_4927);
xnor U5160 (N_5160,N_4914,N_4883);
nor U5161 (N_5161,N_4940,N_4970);
or U5162 (N_5162,N_4860,N_4969);
xnor U5163 (N_5163,N_4881,N_4857);
nand U5164 (N_5164,N_4812,N_4837);
nor U5165 (N_5165,N_4945,N_4914);
nand U5166 (N_5166,N_4961,N_4934);
xnor U5167 (N_5167,N_4809,N_4960);
and U5168 (N_5168,N_4978,N_4852);
and U5169 (N_5169,N_4865,N_4808);
or U5170 (N_5170,N_4830,N_4879);
nand U5171 (N_5171,N_4803,N_4857);
and U5172 (N_5172,N_4846,N_4924);
xnor U5173 (N_5173,N_4881,N_4927);
nor U5174 (N_5174,N_4803,N_4913);
or U5175 (N_5175,N_4933,N_4916);
xor U5176 (N_5176,N_4810,N_4819);
nand U5177 (N_5177,N_4828,N_4991);
nor U5178 (N_5178,N_4819,N_4859);
nor U5179 (N_5179,N_4848,N_4802);
nand U5180 (N_5180,N_4924,N_4905);
xnor U5181 (N_5181,N_4873,N_4835);
nand U5182 (N_5182,N_4975,N_4978);
and U5183 (N_5183,N_4813,N_4873);
and U5184 (N_5184,N_4947,N_4807);
nand U5185 (N_5185,N_4920,N_4893);
nand U5186 (N_5186,N_4815,N_4938);
nor U5187 (N_5187,N_4954,N_4816);
nor U5188 (N_5188,N_4987,N_4844);
nor U5189 (N_5189,N_4807,N_4899);
nor U5190 (N_5190,N_4984,N_4838);
nand U5191 (N_5191,N_4889,N_4968);
xnor U5192 (N_5192,N_4824,N_4895);
nand U5193 (N_5193,N_4992,N_4959);
nand U5194 (N_5194,N_4873,N_4962);
xor U5195 (N_5195,N_4902,N_4815);
nand U5196 (N_5196,N_4872,N_4827);
nor U5197 (N_5197,N_4833,N_4859);
and U5198 (N_5198,N_4961,N_4987);
nand U5199 (N_5199,N_4948,N_4938);
nor U5200 (N_5200,N_5162,N_5183);
and U5201 (N_5201,N_5029,N_5111);
nor U5202 (N_5202,N_5186,N_5173);
xnor U5203 (N_5203,N_5081,N_5044);
xnor U5204 (N_5204,N_5161,N_5055);
nand U5205 (N_5205,N_5128,N_5062);
nor U5206 (N_5206,N_5066,N_5061);
or U5207 (N_5207,N_5140,N_5035);
nand U5208 (N_5208,N_5040,N_5042);
nand U5209 (N_5209,N_5129,N_5102);
nand U5210 (N_5210,N_5075,N_5164);
nand U5211 (N_5211,N_5043,N_5086);
xor U5212 (N_5212,N_5108,N_5130);
nand U5213 (N_5213,N_5022,N_5178);
xor U5214 (N_5214,N_5098,N_5009);
xor U5215 (N_5215,N_5182,N_5069);
xor U5216 (N_5216,N_5031,N_5060);
xor U5217 (N_5217,N_5197,N_5045);
and U5218 (N_5218,N_5017,N_5087);
and U5219 (N_5219,N_5125,N_5020);
nand U5220 (N_5220,N_5041,N_5167);
xor U5221 (N_5221,N_5170,N_5100);
nand U5222 (N_5222,N_5056,N_5166);
nor U5223 (N_5223,N_5082,N_5065);
xnor U5224 (N_5224,N_5090,N_5131);
nand U5225 (N_5225,N_5172,N_5033);
nand U5226 (N_5226,N_5169,N_5025);
and U5227 (N_5227,N_5119,N_5126);
nor U5228 (N_5228,N_5059,N_5010);
nor U5229 (N_5229,N_5142,N_5000);
and U5230 (N_5230,N_5146,N_5021);
and U5231 (N_5231,N_5195,N_5192);
or U5232 (N_5232,N_5027,N_5068);
and U5233 (N_5233,N_5063,N_5136);
xnor U5234 (N_5234,N_5004,N_5085);
and U5235 (N_5235,N_5015,N_5171);
xnor U5236 (N_5236,N_5185,N_5077);
or U5237 (N_5237,N_5046,N_5092);
xnor U5238 (N_5238,N_5123,N_5121);
nor U5239 (N_5239,N_5096,N_5093);
xor U5240 (N_5240,N_5156,N_5157);
nand U5241 (N_5241,N_5023,N_5012);
and U5242 (N_5242,N_5113,N_5196);
and U5243 (N_5243,N_5064,N_5104);
or U5244 (N_5244,N_5099,N_5198);
and U5245 (N_5245,N_5188,N_5187);
nand U5246 (N_5246,N_5148,N_5194);
xor U5247 (N_5247,N_5117,N_5003);
xnor U5248 (N_5248,N_5073,N_5080);
xor U5249 (N_5249,N_5165,N_5176);
nand U5250 (N_5250,N_5155,N_5184);
nand U5251 (N_5251,N_5039,N_5071);
nor U5252 (N_5252,N_5137,N_5134);
nor U5253 (N_5253,N_5024,N_5103);
xor U5254 (N_5254,N_5114,N_5118);
and U5255 (N_5255,N_5079,N_5106);
and U5256 (N_5256,N_5135,N_5122);
and U5257 (N_5257,N_5151,N_5149);
nand U5258 (N_5258,N_5175,N_5067);
nand U5259 (N_5259,N_5047,N_5048);
nand U5260 (N_5260,N_5005,N_5091);
nand U5261 (N_5261,N_5002,N_5138);
nand U5262 (N_5262,N_5018,N_5150);
nand U5263 (N_5263,N_5038,N_5174);
xor U5264 (N_5264,N_5132,N_5115);
and U5265 (N_5265,N_5084,N_5070);
nand U5266 (N_5266,N_5034,N_5141);
xnor U5267 (N_5267,N_5158,N_5139);
xnor U5268 (N_5268,N_5057,N_5014);
nand U5269 (N_5269,N_5190,N_5144);
xnor U5270 (N_5270,N_5049,N_5008);
nor U5271 (N_5271,N_5052,N_5036);
xnor U5272 (N_5272,N_5127,N_5006);
and U5273 (N_5273,N_5168,N_5199);
nand U5274 (N_5274,N_5179,N_5112);
and U5275 (N_5275,N_5078,N_5133);
nand U5276 (N_5276,N_5030,N_5097);
nand U5277 (N_5277,N_5189,N_5001);
or U5278 (N_5278,N_5094,N_5083);
nand U5279 (N_5279,N_5153,N_5054);
nor U5280 (N_5280,N_5180,N_5124);
xnor U5281 (N_5281,N_5107,N_5145);
or U5282 (N_5282,N_5028,N_5019);
and U5283 (N_5283,N_5076,N_5058);
nor U5284 (N_5284,N_5051,N_5154);
and U5285 (N_5285,N_5050,N_5072);
xor U5286 (N_5286,N_5026,N_5143);
or U5287 (N_5287,N_5032,N_5074);
and U5288 (N_5288,N_5110,N_5037);
and U5289 (N_5289,N_5016,N_5181);
and U5290 (N_5290,N_5105,N_5011);
xor U5291 (N_5291,N_5159,N_5013);
nand U5292 (N_5292,N_5160,N_5177);
or U5293 (N_5293,N_5088,N_5120);
and U5294 (N_5294,N_5191,N_5095);
nor U5295 (N_5295,N_5152,N_5116);
nand U5296 (N_5296,N_5101,N_5163);
xor U5297 (N_5297,N_5089,N_5147);
or U5298 (N_5298,N_5109,N_5193);
nand U5299 (N_5299,N_5053,N_5007);
xor U5300 (N_5300,N_5089,N_5082);
xnor U5301 (N_5301,N_5154,N_5147);
or U5302 (N_5302,N_5028,N_5078);
nand U5303 (N_5303,N_5134,N_5040);
nor U5304 (N_5304,N_5198,N_5095);
xor U5305 (N_5305,N_5111,N_5181);
xnor U5306 (N_5306,N_5166,N_5180);
nand U5307 (N_5307,N_5169,N_5148);
and U5308 (N_5308,N_5158,N_5138);
xor U5309 (N_5309,N_5066,N_5196);
nand U5310 (N_5310,N_5083,N_5172);
and U5311 (N_5311,N_5077,N_5057);
nor U5312 (N_5312,N_5022,N_5109);
and U5313 (N_5313,N_5005,N_5139);
xor U5314 (N_5314,N_5116,N_5125);
and U5315 (N_5315,N_5136,N_5179);
or U5316 (N_5316,N_5124,N_5145);
nor U5317 (N_5317,N_5042,N_5029);
nand U5318 (N_5318,N_5072,N_5019);
or U5319 (N_5319,N_5083,N_5122);
or U5320 (N_5320,N_5149,N_5183);
nand U5321 (N_5321,N_5145,N_5161);
or U5322 (N_5322,N_5081,N_5187);
and U5323 (N_5323,N_5120,N_5199);
nand U5324 (N_5324,N_5104,N_5088);
or U5325 (N_5325,N_5053,N_5070);
nand U5326 (N_5326,N_5109,N_5106);
or U5327 (N_5327,N_5134,N_5133);
nor U5328 (N_5328,N_5186,N_5059);
nand U5329 (N_5329,N_5061,N_5182);
xnor U5330 (N_5330,N_5177,N_5055);
nand U5331 (N_5331,N_5058,N_5053);
nor U5332 (N_5332,N_5097,N_5187);
or U5333 (N_5333,N_5183,N_5175);
xor U5334 (N_5334,N_5134,N_5001);
and U5335 (N_5335,N_5077,N_5177);
and U5336 (N_5336,N_5018,N_5143);
xor U5337 (N_5337,N_5137,N_5085);
nor U5338 (N_5338,N_5049,N_5119);
xnor U5339 (N_5339,N_5082,N_5199);
nand U5340 (N_5340,N_5118,N_5160);
or U5341 (N_5341,N_5012,N_5103);
or U5342 (N_5342,N_5163,N_5138);
and U5343 (N_5343,N_5081,N_5039);
and U5344 (N_5344,N_5196,N_5131);
xnor U5345 (N_5345,N_5162,N_5091);
nand U5346 (N_5346,N_5166,N_5185);
nand U5347 (N_5347,N_5080,N_5199);
nand U5348 (N_5348,N_5090,N_5197);
nor U5349 (N_5349,N_5070,N_5198);
and U5350 (N_5350,N_5101,N_5084);
nor U5351 (N_5351,N_5144,N_5112);
and U5352 (N_5352,N_5050,N_5156);
xnor U5353 (N_5353,N_5121,N_5165);
xor U5354 (N_5354,N_5124,N_5014);
and U5355 (N_5355,N_5190,N_5025);
and U5356 (N_5356,N_5167,N_5020);
nor U5357 (N_5357,N_5151,N_5059);
nand U5358 (N_5358,N_5189,N_5004);
nor U5359 (N_5359,N_5127,N_5156);
and U5360 (N_5360,N_5036,N_5128);
nor U5361 (N_5361,N_5016,N_5140);
xor U5362 (N_5362,N_5177,N_5137);
and U5363 (N_5363,N_5045,N_5151);
or U5364 (N_5364,N_5063,N_5118);
or U5365 (N_5365,N_5045,N_5006);
nand U5366 (N_5366,N_5171,N_5058);
xor U5367 (N_5367,N_5141,N_5169);
and U5368 (N_5368,N_5102,N_5041);
or U5369 (N_5369,N_5144,N_5165);
xnor U5370 (N_5370,N_5127,N_5182);
nand U5371 (N_5371,N_5115,N_5178);
and U5372 (N_5372,N_5058,N_5018);
nor U5373 (N_5373,N_5003,N_5162);
nor U5374 (N_5374,N_5027,N_5092);
and U5375 (N_5375,N_5031,N_5142);
xor U5376 (N_5376,N_5193,N_5085);
or U5377 (N_5377,N_5121,N_5151);
and U5378 (N_5378,N_5047,N_5175);
nor U5379 (N_5379,N_5036,N_5126);
and U5380 (N_5380,N_5145,N_5027);
xor U5381 (N_5381,N_5117,N_5156);
or U5382 (N_5382,N_5082,N_5134);
or U5383 (N_5383,N_5190,N_5040);
and U5384 (N_5384,N_5134,N_5096);
nand U5385 (N_5385,N_5068,N_5191);
nor U5386 (N_5386,N_5026,N_5101);
and U5387 (N_5387,N_5023,N_5161);
or U5388 (N_5388,N_5085,N_5038);
or U5389 (N_5389,N_5190,N_5009);
or U5390 (N_5390,N_5004,N_5007);
nor U5391 (N_5391,N_5166,N_5107);
xnor U5392 (N_5392,N_5077,N_5058);
nand U5393 (N_5393,N_5006,N_5102);
xnor U5394 (N_5394,N_5150,N_5048);
nand U5395 (N_5395,N_5092,N_5059);
and U5396 (N_5396,N_5087,N_5144);
nor U5397 (N_5397,N_5044,N_5127);
nor U5398 (N_5398,N_5004,N_5042);
and U5399 (N_5399,N_5012,N_5127);
or U5400 (N_5400,N_5264,N_5338);
and U5401 (N_5401,N_5350,N_5301);
and U5402 (N_5402,N_5229,N_5364);
and U5403 (N_5403,N_5304,N_5331);
nand U5404 (N_5404,N_5297,N_5333);
xnor U5405 (N_5405,N_5294,N_5245);
and U5406 (N_5406,N_5319,N_5345);
and U5407 (N_5407,N_5215,N_5390);
or U5408 (N_5408,N_5380,N_5210);
or U5409 (N_5409,N_5286,N_5205);
nor U5410 (N_5410,N_5358,N_5361);
xnor U5411 (N_5411,N_5397,N_5365);
and U5412 (N_5412,N_5256,N_5267);
xnor U5413 (N_5413,N_5370,N_5296);
or U5414 (N_5414,N_5398,N_5399);
xor U5415 (N_5415,N_5271,N_5298);
nor U5416 (N_5416,N_5300,N_5336);
and U5417 (N_5417,N_5248,N_5353);
and U5418 (N_5418,N_5280,N_5208);
xnor U5419 (N_5419,N_5234,N_5363);
or U5420 (N_5420,N_5242,N_5239);
xnor U5421 (N_5421,N_5277,N_5275);
nand U5422 (N_5422,N_5238,N_5213);
nand U5423 (N_5423,N_5263,N_5240);
xnor U5424 (N_5424,N_5295,N_5352);
or U5425 (N_5425,N_5327,N_5261);
xnor U5426 (N_5426,N_5321,N_5232);
xor U5427 (N_5427,N_5235,N_5366);
and U5428 (N_5428,N_5318,N_5257);
nand U5429 (N_5429,N_5285,N_5214);
xor U5430 (N_5430,N_5305,N_5243);
or U5431 (N_5431,N_5332,N_5372);
xnor U5432 (N_5432,N_5273,N_5250);
xor U5433 (N_5433,N_5382,N_5226);
or U5434 (N_5434,N_5346,N_5373);
xor U5435 (N_5435,N_5354,N_5367);
nand U5436 (N_5436,N_5309,N_5322);
nor U5437 (N_5437,N_5231,N_5302);
xor U5438 (N_5438,N_5329,N_5233);
or U5439 (N_5439,N_5282,N_5203);
xnor U5440 (N_5440,N_5375,N_5227);
xor U5441 (N_5441,N_5290,N_5284);
and U5442 (N_5442,N_5216,N_5289);
xnor U5443 (N_5443,N_5310,N_5262);
xor U5444 (N_5444,N_5324,N_5209);
nor U5445 (N_5445,N_5320,N_5357);
and U5446 (N_5446,N_5325,N_5218);
and U5447 (N_5447,N_5288,N_5315);
nand U5448 (N_5448,N_5314,N_5394);
xor U5449 (N_5449,N_5337,N_5342);
and U5450 (N_5450,N_5381,N_5278);
nand U5451 (N_5451,N_5389,N_5312);
and U5452 (N_5452,N_5388,N_5244);
nor U5453 (N_5453,N_5323,N_5204);
nand U5454 (N_5454,N_5279,N_5311);
xnor U5455 (N_5455,N_5307,N_5369);
nor U5456 (N_5456,N_5253,N_5211);
and U5457 (N_5457,N_5384,N_5344);
xor U5458 (N_5458,N_5252,N_5236);
nor U5459 (N_5459,N_5270,N_5317);
and U5460 (N_5460,N_5359,N_5330);
or U5461 (N_5461,N_5228,N_5396);
nand U5462 (N_5462,N_5378,N_5386);
and U5463 (N_5463,N_5392,N_5351);
and U5464 (N_5464,N_5308,N_5376);
nand U5465 (N_5465,N_5268,N_5259);
nand U5466 (N_5466,N_5374,N_5339);
or U5467 (N_5467,N_5241,N_5306);
or U5468 (N_5468,N_5303,N_5276);
nor U5469 (N_5469,N_5393,N_5313);
nand U5470 (N_5470,N_5379,N_5222);
nor U5471 (N_5471,N_5217,N_5219);
and U5472 (N_5472,N_5328,N_5334);
nor U5473 (N_5473,N_5237,N_5343);
nor U5474 (N_5474,N_5377,N_5283);
and U5475 (N_5475,N_5355,N_5395);
nand U5476 (N_5476,N_5347,N_5291);
and U5477 (N_5477,N_5247,N_5212);
xor U5478 (N_5478,N_5200,N_5287);
nand U5479 (N_5479,N_5316,N_5266);
or U5480 (N_5480,N_5362,N_5391);
nor U5481 (N_5481,N_5223,N_5254);
and U5482 (N_5482,N_5207,N_5383);
nand U5483 (N_5483,N_5255,N_5348);
xnor U5484 (N_5484,N_5299,N_5360);
and U5485 (N_5485,N_5292,N_5224);
nand U5486 (N_5486,N_5260,N_5272);
nand U5487 (N_5487,N_5368,N_5387);
nor U5488 (N_5488,N_5293,N_5340);
xor U5489 (N_5489,N_5202,N_5265);
or U5490 (N_5490,N_5326,N_5385);
nor U5491 (N_5491,N_5269,N_5371);
xor U5492 (N_5492,N_5251,N_5246);
xnor U5493 (N_5493,N_5201,N_5356);
nor U5494 (N_5494,N_5335,N_5220);
or U5495 (N_5495,N_5341,N_5349);
and U5496 (N_5496,N_5258,N_5281);
or U5497 (N_5497,N_5249,N_5221);
nor U5498 (N_5498,N_5274,N_5230);
or U5499 (N_5499,N_5225,N_5206);
and U5500 (N_5500,N_5389,N_5301);
and U5501 (N_5501,N_5340,N_5370);
xnor U5502 (N_5502,N_5283,N_5347);
or U5503 (N_5503,N_5399,N_5314);
and U5504 (N_5504,N_5305,N_5281);
xor U5505 (N_5505,N_5314,N_5260);
nor U5506 (N_5506,N_5392,N_5229);
and U5507 (N_5507,N_5278,N_5285);
nand U5508 (N_5508,N_5365,N_5339);
or U5509 (N_5509,N_5382,N_5286);
nor U5510 (N_5510,N_5261,N_5248);
xnor U5511 (N_5511,N_5393,N_5321);
or U5512 (N_5512,N_5285,N_5325);
nor U5513 (N_5513,N_5284,N_5390);
nand U5514 (N_5514,N_5240,N_5228);
nor U5515 (N_5515,N_5399,N_5280);
or U5516 (N_5516,N_5322,N_5237);
and U5517 (N_5517,N_5370,N_5209);
nor U5518 (N_5518,N_5276,N_5257);
xnor U5519 (N_5519,N_5231,N_5366);
nor U5520 (N_5520,N_5260,N_5353);
nor U5521 (N_5521,N_5387,N_5231);
and U5522 (N_5522,N_5339,N_5308);
or U5523 (N_5523,N_5211,N_5390);
nand U5524 (N_5524,N_5267,N_5303);
xor U5525 (N_5525,N_5357,N_5229);
or U5526 (N_5526,N_5302,N_5266);
nor U5527 (N_5527,N_5250,N_5268);
nor U5528 (N_5528,N_5331,N_5371);
and U5529 (N_5529,N_5379,N_5277);
nand U5530 (N_5530,N_5210,N_5246);
and U5531 (N_5531,N_5320,N_5326);
nand U5532 (N_5532,N_5202,N_5293);
or U5533 (N_5533,N_5260,N_5359);
nor U5534 (N_5534,N_5294,N_5240);
nor U5535 (N_5535,N_5285,N_5209);
nand U5536 (N_5536,N_5368,N_5376);
nand U5537 (N_5537,N_5241,N_5244);
or U5538 (N_5538,N_5204,N_5279);
or U5539 (N_5539,N_5298,N_5248);
nor U5540 (N_5540,N_5316,N_5229);
nand U5541 (N_5541,N_5320,N_5377);
nor U5542 (N_5542,N_5347,N_5350);
xor U5543 (N_5543,N_5214,N_5205);
nor U5544 (N_5544,N_5343,N_5285);
nor U5545 (N_5545,N_5272,N_5212);
or U5546 (N_5546,N_5305,N_5303);
nand U5547 (N_5547,N_5378,N_5273);
xnor U5548 (N_5548,N_5320,N_5255);
nand U5549 (N_5549,N_5265,N_5319);
xnor U5550 (N_5550,N_5342,N_5225);
nor U5551 (N_5551,N_5228,N_5248);
nor U5552 (N_5552,N_5263,N_5321);
and U5553 (N_5553,N_5393,N_5210);
or U5554 (N_5554,N_5246,N_5242);
nand U5555 (N_5555,N_5285,N_5247);
and U5556 (N_5556,N_5274,N_5315);
nand U5557 (N_5557,N_5237,N_5394);
xnor U5558 (N_5558,N_5214,N_5222);
and U5559 (N_5559,N_5378,N_5362);
xnor U5560 (N_5560,N_5200,N_5313);
nand U5561 (N_5561,N_5204,N_5360);
or U5562 (N_5562,N_5365,N_5316);
nor U5563 (N_5563,N_5253,N_5355);
xnor U5564 (N_5564,N_5274,N_5237);
and U5565 (N_5565,N_5350,N_5240);
and U5566 (N_5566,N_5241,N_5351);
xnor U5567 (N_5567,N_5284,N_5211);
and U5568 (N_5568,N_5356,N_5242);
nor U5569 (N_5569,N_5378,N_5340);
and U5570 (N_5570,N_5305,N_5344);
nand U5571 (N_5571,N_5240,N_5291);
or U5572 (N_5572,N_5350,N_5273);
nand U5573 (N_5573,N_5253,N_5265);
nor U5574 (N_5574,N_5278,N_5289);
nand U5575 (N_5575,N_5360,N_5283);
nand U5576 (N_5576,N_5361,N_5272);
xor U5577 (N_5577,N_5388,N_5214);
nor U5578 (N_5578,N_5287,N_5236);
nand U5579 (N_5579,N_5205,N_5325);
and U5580 (N_5580,N_5393,N_5346);
and U5581 (N_5581,N_5252,N_5347);
nand U5582 (N_5582,N_5354,N_5373);
or U5583 (N_5583,N_5300,N_5349);
nor U5584 (N_5584,N_5328,N_5351);
or U5585 (N_5585,N_5249,N_5201);
nand U5586 (N_5586,N_5204,N_5361);
xnor U5587 (N_5587,N_5399,N_5307);
nor U5588 (N_5588,N_5226,N_5344);
nand U5589 (N_5589,N_5309,N_5361);
or U5590 (N_5590,N_5221,N_5263);
and U5591 (N_5591,N_5330,N_5342);
xor U5592 (N_5592,N_5360,N_5277);
nor U5593 (N_5593,N_5393,N_5365);
or U5594 (N_5594,N_5352,N_5364);
xor U5595 (N_5595,N_5366,N_5319);
or U5596 (N_5596,N_5222,N_5223);
xnor U5597 (N_5597,N_5391,N_5277);
nand U5598 (N_5598,N_5333,N_5220);
nand U5599 (N_5599,N_5353,N_5376);
nor U5600 (N_5600,N_5497,N_5470);
or U5601 (N_5601,N_5591,N_5402);
and U5602 (N_5602,N_5520,N_5427);
nand U5603 (N_5603,N_5552,N_5474);
and U5604 (N_5604,N_5494,N_5473);
nor U5605 (N_5605,N_5429,N_5525);
and U5606 (N_5606,N_5410,N_5440);
nand U5607 (N_5607,N_5471,N_5422);
and U5608 (N_5608,N_5513,N_5516);
nor U5609 (N_5609,N_5508,N_5523);
and U5610 (N_5610,N_5456,N_5515);
and U5611 (N_5611,N_5448,N_5401);
xor U5612 (N_5612,N_5576,N_5400);
or U5613 (N_5613,N_5495,N_5561);
and U5614 (N_5614,N_5522,N_5578);
xor U5615 (N_5615,N_5535,N_5486);
and U5616 (N_5616,N_5519,N_5594);
xor U5617 (N_5617,N_5595,N_5452);
nor U5618 (N_5618,N_5506,N_5435);
xnor U5619 (N_5619,N_5544,N_5537);
nor U5620 (N_5620,N_5527,N_5458);
nand U5621 (N_5621,N_5479,N_5437);
nor U5622 (N_5622,N_5581,N_5469);
xor U5623 (N_5623,N_5504,N_5500);
and U5624 (N_5624,N_5570,N_5414);
nand U5625 (N_5625,N_5457,N_5450);
xor U5626 (N_5626,N_5404,N_5579);
or U5627 (N_5627,N_5419,N_5518);
and U5628 (N_5628,N_5490,N_5444);
and U5629 (N_5629,N_5511,N_5485);
or U5630 (N_5630,N_5467,N_5549);
or U5631 (N_5631,N_5492,N_5534);
and U5632 (N_5632,N_5586,N_5453);
or U5633 (N_5633,N_5465,N_5558);
or U5634 (N_5634,N_5424,N_5573);
or U5635 (N_5635,N_5460,N_5517);
and U5636 (N_5636,N_5445,N_5464);
or U5637 (N_5637,N_5468,N_5430);
xnor U5638 (N_5638,N_5454,N_5564);
or U5639 (N_5639,N_5597,N_5530);
xor U5640 (N_5640,N_5416,N_5582);
nand U5641 (N_5641,N_5491,N_5569);
xnor U5642 (N_5642,N_5463,N_5590);
or U5643 (N_5643,N_5541,N_5439);
xor U5644 (N_5644,N_5554,N_5426);
nor U5645 (N_5645,N_5560,N_5451);
and U5646 (N_5646,N_5598,N_5483);
or U5647 (N_5647,N_5551,N_5553);
and U5648 (N_5648,N_5428,N_5466);
and U5649 (N_5649,N_5446,N_5487);
or U5650 (N_5650,N_5443,N_5455);
xor U5651 (N_5651,N_5543,N_5447);
nand U5652 (N_5652,N_5555,N_5412);
and U5653 (N_5653,N_5545,N_5559);
nand U5654 (N_5654,N_5565,N_5580);
nand U5655 (N_5655,N_5438,N_5417);
or U5656 (N_5656,N_5584,N_5484);
and U5657 (N_5657,N_5433,N_5538);
xor U5658 (N_5658,N_5481,N_5592);
xnor U5659 (N_5659,N_5585,N_5415);
xnor U5660 (N_5660,N_5524,N_5418);
nor U5661 (N_5661,N_5432,N_5501);
and U5662 (N_5662,N_5461,N_5539);
xor U5663 (N_5663,N_5509,N_5548);
or U5664 (N_5664,N_5434,N_5406);
nand U5665 (N_5665,N_5420,N_5533);
or U5666 (N_5666,N_5512,N_5507);
or U5667 (N_5667,N_5547,N_5557);
xnor U5668 (N_5668,N_5567,N_5472);
nor U5669 (N_5669,N_5587,N_5405);
xnor U5670 (N_5670,N_5514,N_5409);
nand U5671 (N_5671,N_5480,N_5449);
nand U5672 (N_5672,N_5496,N_5599);
xor U5673 (N_5673,N_5566,N_5459);
or U5674 (N_5674,N_5563,N_5413);
xnor U5675 (N_5675,N_5489,N_5482);
nor U5676 (N_5676,N_5540,N_5442);
or U5677 (N_5677,N_5531,N_5403);
and U5678 (N_5678,N_5536,N_5493);
or U5679 (N_5679,N_5577,N_5546);
xnor U5680 (N_5680,N_5571,N_5441);
nand U5681 (N_5681,N_5568,N_5510);
and U5682 (N_5682,N_5550,N_5477);
nand U5683 (N_5683,N_5532,N_5498);
or U5684 (N_5684,N_5476,N_5588);
nand U5685 (N_5685,N_5488,N_5572);
and U5686 (N_5686,N_5436,N_5407);
nand U5687 (N_5687,N_5521,N_5423);
nand U5688 (N_5688,N_5478,N_5583);
nor U5689 (N_5689,N_5502,N_5593);
or U5690 (N_5690,N_5589,N_5505);
nand U5691 (N_5691,N_5556,N_5596);
nor U5692 (N_5692,N_5562,N_5462);
or U5693 (N_5693,N_5499,N_5411);
nand U5694 (N_5694,N_5529,N_5425);
and U5695 (N_5695,N_5431,N_5575);
or U5696 (N_5696,N_5574,N_5421);
and U5697 (N_5697,N_5475,N_5542);
nand U5698 (N_5698,N_5526,N_5528);
nor U5699 (N_5699,N_5408,N_5503);
xor U5700 (N_5700,N_5510,N_5519);
or U5701 (N_5701,N_5413,N_5409);
nor U5702 (N_5702,N_5453,N_5442);
or U5703 (N_5703,N_5507,N_5458);
and U5704 (N_5704,N_5514,N_5463);
and U5705 (N_5705,N_5577,N_5562);
or U5706 (N_5706,N_5467,N_5470);
nor U5707 (N_5707,N_5585,N_5590);
xor U5708 (N_5708,N_5485,N_5571);
xnor U5709 (N_5709,N_5592,N_5451);
nand U5710 (N_5710,N_5584,N_5490);
nand U5711 (N_5711,N_5583,N_5468);
or U5712 (N_5712,N_5549,N_5411);
xnor U5713 (N_5713,N_5466,N_5494);
or U5714 (N_5714,N_5421,N_5496);
xnor U5715 (N_5715,N_5401,N_5414);
or U5716 (N_5716,N_5464,N_5448);
and U5717 (N_5717,N_5510,N_5509);
and U5718 (N_5718,N_5458,N_5547);
nor U5719 (N_5719,N_5501,N_5415);
and U5720 (N_5720,N_5498,N_5453);
xor U5721 (N_5721,N_5438,N_5425);
nand U5722 (N_5722,N_5589,N_5590);
xnor U5723 (N_5723,N_5439,N_5505);
and U5724 (N_5724,N_5579,N_5513);
or U5725 (N_5725,N_5533,N_5531);
nand U5726 (N_5726,N_5516,N_5571);
nand U5727 (N_5727,N_5506,N_5583);
nor U5728 (N_5728,N_5449,N_5411);
nor U5729 (N_5729,N_5452,N_5504);
nor U5730 (N_5730,N_5437,N_5594);
xor U5731 (N_5731,N_5553,N_5416);
and U5732 (N_5732,N_5471,N_5481);
nand U5733 (N_5733,N_5408,N_5453);
and U5734 (N_5734,N_5544,N_5588);
nor U5735 (N_5735,N_5599,N_5436);
xor U5736 (N_5736,N_5479,N_5518);
nand U5737 (N_5737,N_5566,N_5480);
nor U5738 (N_5738,N_5533,N_5583);
nor U5739 (N_5739,N_5419,N_5582);
nor U5740 (N_5740,N_5520,N_5568);
xnor U5741 (N_5741,N_5403,N_5401);
or U5742 (N_5742,N_5491,N_5478);
nand U5743 (N_5743,N_5598,N_5549);
nand U5744 (N_5744,N_5510,N_5497);
or U5745 (N_5745,N_5516,N_5511);
and U5746 (N_5746,N_5480,N_5430);
nand U5747 (N_5747,N_5562,N_5458);
nand U5748 (N_5748,N_5501,N_5523);
or U5749 (N_5749,N_5559,N_5427);
nand U5750 (N_5750,N_5595,N_5406);
xnor U5751 (N_5751,N_5482,N_5475);
or U5752 (N_5752,N_5437,N_5476);
or U5753 (N_5753,N_5562,N_5508);
xor U5754 (N_5754,N_5568,N_5476);
and U5755 (N_5755,N_5469,N_5475);
or U5756 (N_5756,N_5577,N_5541);
and U5757 (N_5757,N_5540,N_5596);
nand U5758 (N_5758,N_5448,N_5533);
or U5759 (N_5759,N_5583,N_5580);
or U5760 (N_5760,N_5565,N_5490);
or U5761 (N_5761,N_5402,N_5568);
or U5762 (N_5762,N_5519,N_5473);
nor U5763 (N_5763,N_5525,N_5515);
and U5764 (N_5764,N_5461,N_5492);
nand U5765 (N_5765,N_5403,N_5500);
or U5766 (N_5766,N_5410,N_5505);
and U5767 (N_5767,N_5484,N_5457);
nor U5768 (N_5768,N_5443,N_5574);
nand U5769 (N_5769,N_5414,N_5550);
xor U5770 (N_5770,N_5512,N_5459);
and U5771 (N_5771,N_5506,N_5590);
nand U5772 (N_5772,N_5599,N_5485);
nor U5773 (N_5773,N_5516,N_5530);
xnor U5774 (N_5774,N_5539,N_5452);
nor U5775 (N_5775,N_5401,N_5564);
nand U5776 (N_5776,N_5505,N_5503);
xor U5777 (N_5777,N_5445,N_5567);
or U5778 (N_5778,N_5535,N_5504);
or U5779 (N_5779,N_5594,N_5517);
and U5780 (N_5780,N_5589,N_5571);
or U5781 (N_5781,N_5575,N_5598);
or U5782 (N_5782,N_5560,N_5447);
nor U5783 (N_5783,N_5541,N_5420);
and U5784 (N_5784,N_5441,N_5471);
xnor U5785 (N_5785,N_5422,N_5535);
nor U5786 (N_5786,N_5545,N_5533);
nor U5787 (N_5787,N_5589,N_5503);
nand U5788 (N_5788,N_5478,N_5451);
nor U5789 (N_5789,N_5569,N_5404);
nor U5790 (N_5790,N_5529,N_5587);
xor U5791 (N_5791,N_5516,N_5558);
xor U5792 (N_5792,N_5534,N_5523);
or U5793 (N_5793,N_5447,N_5454);
or U5794 (N_5794,N_5467,N_5407);
xnor U5795 (N_5795,N_5448,N_5480);
nor U5796 (N_5796,N_5418,N_5594);
xor U5797 (N_5797,N_5566,N_5438);
or U5798 (N_5798,N_5406,N_5402);
xnor U5799 (N_5799,N_5458,N_5535);
or U5800 (N_5800,N_5657,N_5739);
nand U5801 (N_5801,N_5711,N_5617);
and U5802 (N_5802,N_5632,N_5783);
nor U5803 (N_5803,N_5627,N_5729);
and U5804 (N_5804,N_5713,N_5731);
nor U5805 (N_5805,N_5604,N_5695);
and U5806 (N_5806,N_5670,N_5754);
xor U5807 (N_5807,N_5792,N_5672);
and U5808 (N_5808,N_5720,N_5753);
xnor U5809 (N_5809,N_5730,N_5669);
nor U5810 (N_5810,N_5714,N_5796);
and U5811 (N_5811,N_5721,N_5733);
nand U5812 (N_5812,N_5778,N_5775);
xnor U5813 (N_5813,N_5781,N_5660);
or U5814 (N_5814,N_5740,N_5789);
xnor U5815 (N_5815,N_5709,N_5636);
xor U5816 (N_5816,N_5697,N_5654);
nand U5817 (N_5817,N_5759,N_5765);
nor U5818 (N_5818,N_5652,N_5630);
xor U5819 (N_5819,N_5794,N_5722);
xnor U5820 (N_5820,N_5675,N_5743);
xor U5821 (N_5821,N_5648,N_5756);
xnor U5822 (N_5822,N_5708,N_5724);
nand U5823 (N_5823,N_5668,N_5760);
and U5824 (N_5824,N_5767,N_5639);
and U5825 (N_5825,N_5752,N_5622);
or U5826 (N_5826,N_5629,N_5726);
and U5827 (N_5827,N_5791,N_5614);
nand U5828 (N_5828,N_5699,N_5625);
xor U5829 (N_5829,N_5640,N_5600);
nor U5830 (N_5830,N_5725,N_5661);
and U5831 (N_5831,N_5703,N_5676);
nand U5832 (N_5832,N_5601,N_5717);
nand U5833 (N_5833,N_5768,N_5777);
or U5834 (N_5834,N_5665,N_5795);
nor U5835 (N_5835,N_5646,N_5626);
nor U5836 (N_5836,N_5691,N_5749);
or U5837 (N_5837,N_5776,N_5647);
nor U5838 (N_5838,N_5611,N_5613);
and U5839 (N_5839,N_5738,N_5693);
or U5840 (N_5840,N_5719,N_5787);
or U5841 (N_5841,N_5679,N_5698);
nor U5842 (N_5842,N_5710,N_5742);
and U5843 (N_5843,N_5705,N_5655);
xor U5844 (N_5844,N_5761,N_5659);
xnor U5845 (N_5845,N_5690,N_5653);
nand U5846 (N_5846,N_5701,N_5620);
and U5847 (N_5847,N_5638,N_5678);
or U5848 (N_5848,N_5689,N_5658);
xnor U5849 (N_5849,N_5618,N_5764);
and U5850 (N_5850,N_5667,N_5688);
nor U5851 (N_5851,N_5735,N_5737);
and U5852 (N_5852,N_5741,N_5766);
xnor U5853 (N_5853,N_5680,N_5798);
or U5854 (N_5854,N_5758,N_5633);
nor U5855 (N_5855,N_5784,N_5612);
and U5856 (N_5856,N_5694,N_5687);
and U5857 (N_5857,N_5684,N_5619);
or U5858 (N_5858,N_5706,N_5723);
nor U5859 (N_5859,N_5779,N_5769);
nand U5860 (N_5860,N_5797,N_5696);
or U5861 (N_5861,N_5603,N_5606);
nand U5862 (N_5862,N_5677,N_5763);
xor U5863 (N_5863,N_5750,N_5683);
nand U5864 (N_5864,N_5692,N_5650);
or U5865 (N_5865,N_5605,N_5642);
xnor U5866 (N_5866,N_5744,N_5718);
nor U5867 (N_5867,N_5637,N_5727);
xor U5868 (N_5868,N_5634,N_5751);
nand U5869 (N_5869,N_5607,N_5762);
nand U5870 (N_5870,N_5662,N_5685);
and U5871 (N_5871,N_5786,N_5746);
xor U5872 (N_5872,N_5712,N_5773);
nand U5873 (N_5873,N_5715,N_5748);
or U5874 (N_5874,N_5628,N_5608);
nor U5875 (N_5875,N_5610,N_5602);
xor U5876 (N_5876,N_5757,N_5770);
or U5877 (N_5877,N_5674,N_5671);
or U5878 (N_5878,N_5704,N_5774);
nand U5879 (N_5879,N_5621,N_5673);
and U5880 (N_5880,N_5790,N_5651);
xor U5881 (N_5881,N_5780,N_5609);
or U5882 (N_5882,N_5666,N_5641);
or U5883 (N_5883,N_5793,N_5616);
and U5884 (N_5884,N_5799,N_5624);
nand U5885 (N_5885,N_5700,N_5728);
or U5886 (N_5886,N_5707,N_5702);
xor U5887 (N_5887,N_5644,N_5663);
and U5888 (N_5888,N_5747,N_5771);
nor U5889 (N_5889,N_5681,N_5623);
or U5890 (N_5890,N_5772,N_5782);
nor U5891 (N_5891,N_5615,N_5736);
xor U5892 (N_5892,N_5745,N_5645);
and U5893 (N_5893,N_5649,N_5631);
nor U5894 (N_5894,N_5664,N_5755);
xnor U5895 (N_5895,N_5682,N_5635);
or U5896 (N_5896,N_5785,N_5656);
and U5897 (N_5897,N_5732,N_5734);
nand U5898 (N_5898,N_5788,N_5716);
and U5899 (N_5899,N_5686,N_5643);
xnor U5900 (N_5900,N_5767,N_5665);
nand U5901 (N_5901,N_5669,N_5661);
nor U5902 (N_5902,N_5775,N_5755);
or U5903 (N_5903,N_5702,N_5709);
nand U5904 (N_5904,N_5621,N_5785);
nor U5905 (N_5905,N_5640,N_5682);
and U5906 (N_5906,N_5655,N_5632);
xor U5907 (N_5907,N_5613,N_5717);
nor U5908 (N_5908,N_5724,N_5727);
nand U5909 (N_5909,N_5787,N_5684);
and U5910 (N_5910,N_5728,N_5769);
or U5911 (N_5911,N_5783,N_5718);
and U5912 (N_5912,N_5612,N_5724);
and U5913 (N_5913,N_5689,N_5644);
nor U5914 (N_5914,N_5725,N_5784);
or U5915 (N_5915,N_5736,N_5777);
nand U5916 (N_5916,N_5722,N_5628);
nor U5917 (N_5917,N_5699,N_5684);
nor U5918 (N_5918,N_5614,N_5631);
xnor U5919 (N_5919,N_5641,N_5751);
nand U5920 (N_5920,N_5668,N_5612);
and U5921 (N_5921,N_5658,N_5622);
nand U5922 (N_5922,N_5714,N_5636);
nand U5923 (N_5923,N_5756,N_5725);
and U5924 (N_5924,N_5662,N_5734);
nand U5925 (N_5925,N_5717,N_5698);
nand U5926 (N_5926,N_5679,N_5771);
xor U5927 (N_5927,N_5773,N_5767);
nor U5928 (N_5928,N_5729,N_5746);
nor U5929 (N_5929,N_5622,N_5738);
xnor U5930 (N_5930,N_5759,N_5719);
or U5931 (N_5931,N_5691,N_5605);
and U5932 (N_5932,N_5754,N_5679);
nand U5933 (N_5933,N_5675,N_5656);
xnor U5934 (N_5934,N_5749,N_5673);
xnor U5935 (N_5935,N_5787,N_5706);
and U5936 (N_5936,N_5647,N_5778);
nor U5937 (N_5937,N_5708,N_5666);
and U5938 (N_5938,N_5776,N_5728);
nor U5939 (N_5939,N_5643,N_5649);
nand U5940 (N_5940,N_5632,N_5691);
nand U5941 (N_5941,N_5747,N_5756);
and U5942 (N_5942,N_5722,N_5779);
nor U5943 (N_5943,N_5642,N_5610);
nor U5944 (N_5944,N_5754,N_5609);
and U5945 (N_5945,N_5668,N_5741);
nand U5946 (N_5946,N_5798,N_5665);
nand U5947 (N_5947,N_5610,N_5664);
and U5948 (N_5948,N_5608,N_5770);
nor U5949 (N_5949,N_5631,N_5620);
xnor U5950 (N_5950,N_5792,N_5742);
or U5951 (N_5951,N_5651,N_5662);
xor U5952 (N_5952,N_5752,N_5782);
nand U5953 (N_5953,N_5675,N_5650);
and U5954 (N_5954,N_5728,N_5665);
and U5955 (N_5955,N_5678,N_5782);
nand U5956 (N_5956,N_5741,N_5622);
nor U5957 (N_5957,N_5771,N_5769);
or U5958 (N_5958,N_5787,N_5699);
xnor U5959 (N_5959,N_5701,N_5712);
or U5960 (N_5960,N_5798,N_5774);
and U5961 (N_5961,N_5629,N_5670);
nor U5962 (N_5962,N_5731,N_5753);
nand U5963 (N_5963,N_5651,N_5795);
nor U5964 (N_5964,N_5741,N_5702);
and U5965 (N_5965,N_5603,N_5621);
or U5966 (N_5966,N_5777,N_5785);
nand U5967 (N_5967,N_5637,N_5632);
nand U5968 (N_5968,N_5670,N_5605);
or U5969 (N_5969,N_5675,N_5686);
nand U5970 (N_5970,N_5649,N_5779);
nor U5971 (N_5971,N_5680,N_5664);
nor U5972 (N_5972,N_5675,N_5775);
nand U5973 (N_5973,N_5667,N_5789);
nor U5974 (N_5974,N_5733,N_5675);
nand U5975 (N_5975,N_5751,N_5651);
xnor U5976 (N_5976,N_5698,N_5687);
or U5977 (N_5977,N_5628,N_5625);
nor U5978 (N_5978,N_5604,N_5777);
nand U5979 (N_5979,N_5795,N_5768);
xor U5980 (N_5980,N_5781,N_5684);
nor U5981 (N_5981,N_5761,N_5613);
or U5982 (N_5982,N_5727,N_5613);
xor U5983 (N_5983,N_5796,N_5791);
nor U5984 (N_5984,N_5631,N_5732);
nor U5985 (N_5985,N_5659,N_5692);
nand U5986 (N_5986,N_5750,N_5762);
nand U5987 (N_5987,N_5659,N_5661);
and U5988 (N_5988,N_5789,N_5609);
xor U5989 (N_5989,N_5633,N_5699);
or U5990 (N_5990,N_5785,N_5787);
nor U5991 (N_5991,N_5662,N_5655);
nand U5992 (N_5992,N_5682,N_5777);
or U5993 (N_5993,N_5682,N_5697);
nor U5994 (N_5994,N_5682,N_5645);
and U5995 (N_5995,N_5742,N_5757);
or U5996 (N_5996,N_5743,N_5647);
and U5997 (N_5997,N_5688,N_5651);
and U5998 (N_5998,N_5651,N_5608);
nand U5999 (N_5999,N_5775,N_5760);
or U6000 (N_6000,N_5934,N_5814);
and U6001 (N_6001,N_5972,N_5802);
xor U6002 (N_6002,N_5822,N_5821);
and U6003 (N_6003,N_5983,N_5836);
and U6004 (N_6004,N_5908,N_5805);
nor U6005 (N_6005,N_5974,N_5964);
or U6006 (N_6006,N_5896,N_5915);
and U6007 (N_6007,N_5911,N_5900);
or U6008 (N_6008,N_5953,N_5895);
nand U6009 (N_6009,N_5993,N_5941);
or U6010 (N_6010,N_5947,N_5855);
nand U6011 (N_6011,N_5962,N_5882);
nor U6012 (N_6012,N_5827,N_5819);
nand U6013 (N_6013,N_5841,N_5881);
or U6014 (N_6014,N_5879,N_5944);
nand U6015 (N_6015,N_5852,N_5975);
nor U6016 (N_6016,N_5825,N_5919);
nor U6017 (N_6017,N_5935,N_5916);
or U6018 (N_6018,N_5869,N_5999);
nor U6019 (N_6019,N_5865,N_5956);
and U6020 (N_6020,N_5890,N_5998);
and U6021 (N_6021,N_5898,N_5897);
and U6022 (N_6022,N_5812,N_5826);
or U6023 (N_6023,N_5989,N_5988);
nand U6024 (N_6024,N_5970,N_5813);
xor U6025 (N_6025,N_5986,N_5816);
or U6026 (N_6026,N_5857,N_5951);
xor U6027 (N_6027,N_5866,N_5880);
or U6028 (N_6028,N_5884,N_5943);
or U6029 (N_6029,N_5864,N_5845);
or U6030 (N_6030,N_5980,N_5823);
or U6031 (N_6031,N_5914,N_5832);
and U6032 (N_6032,N_5838,N_5818);
and U6033 (N_6033,N_5923,N_5842);
xnor U6034 (N_6034,N_5924,N_5876);
or U6035 (N_6035,N_5967,N_5834);
xor U6036 (N_6036,N_5958,N_5912);
nand U6037 (N_6037,N_5867,N_5885);
or U6038 (N_6038,N_5831,N_5913);
and U6039 (N_6039,N_5917,N_5976);
xor U6040 (N_6040,N_5979,N_5874);
and U6041 (N_6041,N_5850,N_5938);
nand U6042 (N_6042,N_5969,N_5939);
and U6043 (N_6043,N_5846,N_5801);
nand U6044 (N_6044,N_5955,N_5905);
or U6045 (N_6045,N_5977,N_5904);
and U6046 (N_6046,N_5968,N_5839);
xor U6047 (N_6047,N_5806,N_5899);
nand U6048 (N_6048,N_5820,N_5803);
or U6049 (N_6049,N_5982,N_5928);
nor U6050 (N_6050,N_5893,N_5875);
xnor U6051 (N_6051,N_5936,N_5957);
nor U6052 (N_6052,N_5851,N_5978);
xor U6053 (N_6053,N_5960,N_5973);
or U6054 (N_6054,N_5868,N_5872);
or U6055 (N_6055,N_5940,N_5931);
nor U6056 (N_6056,N_5824,N_5918);
nand U6057 (N_6057,N_5861,N_5961);
xnor U6058 (N_6058,N_5995,N_5833);
nor U6059 (N_6059,N_5929,N_5949);
nand U6060 (N_6060,N_5933,N_5844);
or U6061 (N_6061,N_5984,N_5921);
xor U6062 (N_6062,N_5990,N_5849);
and U6063 (N_6063,N_5848,N_5971);
and U6064 (N_6064,N_5992,N_5925);
nand U6065 (N_6065,N_5854,N_5950);
nor U6066 (N_6066,N_5922,N_5829);
or U6067 (N_6067,N_5907,N_5817);
xor U6068 (N_6068,N_5809,N_5870);
nand U6069 (N_6069,N_5952,N_5860);
xor U6070 (N_6070,N_5906,N_5889);
xor U6071 (N_6071,N_5840,N_5996);
xnor U6072 (N_6072,N_5828,N_5966);
nor U6073 (N_6073,N_5891,N_5853);
nor U6074 (N_6074,N_5926,N_5887);
or U6075 (N_6075,N_5862,N_5837);
xor U6076 (N_6076,N_5886,N_5883);
nor U6077 (N_6077,N_5945,N_5811);
nor U6078 (N_6078,N_5808,N_5878);
nor U6079 (N_6079,N_5954,N_5859);
and U6080 (N_6080,N_5835,N_5807);
nor U6081 (N_6081,N_5902,N_5903);
nand U6082 (N_6082,N_5997,N_5920);
and U6083 (N_6083,N_5930,N_5843);
or U6084 (N_6084,N_5847,N_5863);
xnor U6085 (N_6085,N_5858,N_5800);
nand U6086 (N_6086,N_5804,N_5871);
xor U6087 (N_6087,N_5894,N_5810);
and U6088 (N_6088,N_5991,N_5927);
xnor U6089 (N_6089,N_5946,N_5856);
nand U6090 (N_6090,N_5937,N_5888);
nor U6091 (N_6091,N_5942,N_5815);
nor U6092 (N_6092,N_5877,N_5932);
nor U6093 (N_6093,N_5965,N_5959);
or U6094 (N_6094,N_5985,N_5981);
or U6095 (N_6095,N_5948,N_5909);
nor U6096 (N_6096,N_5830,N_5901);
nor U6097 (N_6097,N_5873,N_5987);
xnor U6098 (N_6098,N_5910,N_5963);
nor U6099 (N_6099,N_5994,N_5892);
and U6100 (N_6100,N_5823,N_5875);
nor U6101 (N_6101,N_5877,N_5801);
nand U6102 (N_6102,N_5970,N_5960);
nand U6103 (N_6103,N_5891,N_5930);
and U6104 (N_6104,N_5950,N_5859);
or U6105 (N_6105,N_5847,N_5876);
or U6106 (N_6106,N_5832,N_5926);
or U6107 (N_6107,N_5875,N_5835);
or U6108 (N_6108,N_5958,N_5896);
nor U6109 (N_6109,N_5947,N_5938);
nor U6110 (N_6110,N_5824,N_5831);
and U6111 (N_6111,N_5981,N_5972);
and U6112 (N_6112,N_5951,N_5833);
or U6113 (N_6113,N_5951,N_5865);
and U6114 (N_6114,N_5850,N_5961);
and U6115 (N_6115,N_5886,N_5888);
or U6116 (N_6116,N_5984,N_5884);
and U6117 (N_6117,N_5835,N_5955);
nand U6118 (N_6118,N_5937,N_5914);
xnor U6119 (N_6119,N_5922,N_5950);
nand U6120 (N_6120,N_5967,N_5854);
nor U6121 (N_6121,N_5826,N_5988);
nand U6122 (N_6122,N_5919,N_5912);
nor U6123 (N_6123,N_5951,N_5969);
nand U6124 (N_6124,N_5878,N_5981);
nand U6125 (N_6125,N_5970,N_5901);
xnor U6126 (N_6126,N_5919,N_5911);
nor U6127 (N_6127,N_5888,N_5879);
and U6128 (N_6128,N_5904,N_5938);
nand U6129 (N_6129,N_5900,N_5933);
nand U6130 (N_6130,N_5825,N_5948);
xor U6131 (N_6131,N_5901,N_5921);
xnor U6132 (N_6132,N_5910,N_5915);
nand U6133 (N_6133,N_5812,N_5827);
nand U6134 (N_6134,N_5908,N_5928);
and U6135 (N_6135,N_5982,N_5868);
nor U6136 (N_6136,N_5980,N_5994);
nor U6137 (N_6137,N_5872,N_5869);
xnor U6138 (N_6138,N_5962,N_5870);
or U6139 (N_6139,N_5816,N_5926);
nand U6140 (N_6140,N_5976,N_5870);
or U6141 (N_6141,N_5915,N_5988);
nor U6142 (N_6142,N_5823,N_5872);
and U6143 (N_6143,N_5881,N_5823);
nor U6144 (N_6144,N_5909,N_5885);
xor U6145 (N_6145,N_5836,N_5992);
xnor U6146 (N_6146,N_5894,N_5958);
nor U6147 (N_6147,N_5821,N_5857);
nor U6148 (N_6148,N_5861,N_5955);
and U6149 (N_6149,N_5860,N_5916);
nor U6150 (N_6150,N_5994,N_5929);
or U6151 (N_6151,N_5900,N_5949);
nor U6152 (N_6152,N_5933,N_5943);
xnor U6153 (N_6153,N_5873,N_5957);
or U6154 (N_6154,N_5992,N_5921);
and U6155 (N_6155,N_5857,N_5864);
nor U6156 (N_6156,N_5848,N_5884);
or U6157 (N_6157,N_5947,N_5884);
or U6158 (N_6158,N_5891,N_5916);
nor U6159 (N_6159,N_5960,N_5903);
nand U6160 (N_6160,N_5938,N_5935);
or U6161 (N_6161,N_5924,N_5988);
nor U6162 (N_6162,N_5907,N_5949);
nor U6163 (N_6163,N_5816,N_5938);
xnor U6164 (N_6164,N_5839,N_5960);
and U6165 (N_6165,N_5929,N_5963);
and U6166 (N_6166,N_5815,N_5994);
xor U6167 (N_6167,N_5866,N_5929);
nand U6168 (N_6168,N_5853,N_5885);
or U6169 (N_6169,N_5982,N_5804);
xor U6170 (N_6170,N_5931,N_5843);
and U6171 (N_6171,N_5930,N_5831);
xor U6172 (N_6172,N_5889,N_5900);
xor U6173 (N_6173,N_5872,N_5878);
and U6174 (N_6174,N_5940,N_5908);
nand U6175 (N_6175,N_5921,N_5851);
or U6176 (N_6176,N_5878,N_5852);
xor U6177 (N_6177,N_5986,N_5892);
xnor U6178 (N_6178,N_5912,N_5894);
xnor U6179 (N_6179,N_5854,N_5875);
nand U6180 (N_6180,N_5833,N_5882);
nand U6181 (N_6181,N_5817,N_5924);
and U6182 (N_6182,N_5816,N_5941);
nand U6183 (N_6183,N_5943,N_5870);
xor U6184 (N_6184,N_5946,N_5881);
nor U6185 (N_6185,N_5800,N_5902);
xor U6186 (N_6186,N_5913,N_5916);
or U6187 (N_6187,N_5900,N_5872);
xnor U6188 (N_6188,N_5952,N_5989);
nand U6189 (N_6189,N_5855,N_5996);
nand U6190 (N_6190,N_5962,N_5977);
nand U6191 (N_6191,N_5915,N_5949);
xnor U6192 (N_6192,N_5925,N_5902);
and U6193 (N_6193,N_5923,N_5925);
xnor U6194 (N_6194,N_5886,N_5863);
nand U6195 (N_6195,N_5850,N_5924);
nand U6196 (N_6196,N_5909,N_5854);
nor U6197 (N_6197,N_5906,N_5868);
and U6198 (N_6198,N_5907,N_5803);
nand U6199 (N_6199,N_5883,N_5972);
and U6200 (N_6200,N_6015,N_6142);
xor U6201 (N_6201,N_6057,N_6168);
and U6202 (N_6202,N_6184,N_6053);
nor U6203 (N_6203,N_6122,N_6040);
or U6204 (N_6204,N_6108,N_6069);
nand U6205 (N_6205,N_6066,N_6095);
nand U6206 (N_6206,N_6119,N_6139);
and U6207 (N_6207,N_6141,N_6021);
xor U6208 (N_6208,N_6164,N_6110);
or U6209 (N_6209,N_6172,N_6199);
or U6210 (N_6210,N_6050,N_6170);
and U6211 (N_6211,N_6154,N_6012);
or U6212 (N_6212,N_6183,N_6173);
and U6213 (N_6213,N_6043,N_6077);
and U6214 (N_6214,N_6039,N_6175);
or U6215 (N_6215,N_6135,N_6034);
and U6216 (N_6216,N_6017,N_6149);
xor U6217 (N_6217,N_6174,N_6010);
and U6218 (N_6218,N_6032,N_6071);
and U6219 (N_6219,N_6078,N_6148);
nor U6220 (N_6220,N_6006,N_6145);
xnor U6221 (N_6221,N_6190,N_6136);
or U6222 (N_6222,N_6114,N_6089);
or U6223 (N_6223,N_6099,N_6150);
nand U6224 (N_6224,N_6134,N_6091);
and U6225 (N_6225,N_6002,N_6128);
nand U6226 (N_6226,N_6014,N_6127);
and U6227 (N_6227,N_6079,N_6193);
nor U6228 (N_6228,N_6045,N_6062);
or U6229 (N_6229,N_6093,N_6024);
and U6230 (N_6230,N_6185,N_6027);
nor U6231 (N_6231,N_6033,N_6106);
nand U6232 (N_6232,N_6126,N_6060);
or U6233 (N_6233,N_6038,N_6068);
nand U6234 (N_6234,N_6076,N_6169);
nand U6235 (N_6235,N_6054,N_6125);
xor U6236 (N_6236,N_6132,N_6188);
or U6237 (N_6237,N_6196,N_6044);
or U6238 (N_6238,N_6133,N_6101);
nand U6239 (N_6239,N_6178,N_6022);
or U6240 (N_6240,N_6097,N_6020);
nor U6241 (N_6241,N_6162,N_6109);
nor U6242 (N_6242,N_6023,N_6028);
nor U6243 (N_6243,N_6171,N_6088);
and U6244 (N_6244,N_6105,N_6198);
nand U6245 (N_6245,N_6059,N_6072);
and U6246 (N_6246,N_6195,N_6118);
nor U6247 (N_6247,N_6030,N_6011);
nand U6248 (N_6248,N_6115,N_6009);
and U6249 (N_6249,N_6159,N_6092);
and U6250 (N_6250,N_6081,N_6158);
nor U6251 (N_6251,N_6120,N_6004);
nor U6252 (N_6252,N_6058,N_6049);
and U6253 (N_6253,N_6037,N_6075);
and U6254 (N_6254,N_6177,N_6085);
xnor U6255 (N_6255,N_6182,N_6008);
nor U6256 (N_6256,N_6167,N_6143);
nor U6257 (N_6257,N_6098,N_6035);
nor U6258 (N_6258,N_6137,N_6146);
nor U6259 (N_6259,N_6112,N_6191);
and U6260 (N_6260,N_6123,N_6055);
and U6261 (N_6261,N_6065,N_6061);
xnor U6262 (N_6262,N_6100,N_6003);
xnor U6263 (N_6263,N_6147,N_6155);
xor U6264 (N_6264,N_6111,N_6018);
xnor U6265 (N_6265,N_6063,N_6186);
xnor U6266 (N_6266,N_6082,N_6036);
nand U6267 (N_6267,N_6181,N_6031);
nand U6268 (N_6268,N_6102,N_6090);
nand U6269 (N_6269,N_6073,N_6083);
or U6270 (N_6270,N_6176,N_6192);
or U6271 (N_6271,N_6086,N_6047);
and U6272 (N_6272,N_6187,N_6140);
nor U6273 (N_6273,N_6016,N_6151);
nand U6274 (N_6274,N_6056,N_6052);
nor U6275 (N_6275,N_6084,N_6051);
nand U6276 (N_6276,N_6165,N_6129);
xnor U6277 (N_6277,N_6144,N_6121);
or U6278 (N_6278,N_6029,N_6046);
nor U6279 (N_6279,N_6104,N_6074);
nor U6280 (N_6280,N_6026,N_6042);
nand U6281 (N_6281,N_6107,N_6152);
nor U6282 (N_6282,N_6138,N_6013);
nand U6283 (N_6283,N_6103,N_6130);
and U6284 (N_6284,N_6160,N_6131);
nand U6285 (N_6285,N_6197,N_6001);
xnor U6286 (N_6286,N_6041,N_6000);
nor U6287 (N_6287,N_6080,N_6048);
nand U6288 (N_6288,N_6067,N_6179);
nor U6289 (N_6289,N_6070,N_6157);
xor U6290 (N_6290,N_6116,N_6025);
xnor U6291 (N_6291,N_6189,N_6087);
nand U6292 (N_6292,N_6156,N_6117);
and U6293 (N_6293,N_6166,N_6194);
xor U6294 (N_6294,N_6007,N_6113);
nand U6295 (N_6295,N_6005,N_6096);
xor U6296 (N_6296,N_6094,N_6064);
or U6297 (N_6297,N_6161,N_6019);
and U6298 (N_6298,N_6153,N_6163);
nor U6299 (N_6299,N_6180,N_6124);
and U6300 (N_6300,N_6074,N_6175);
and U6301 (N_6301,N_6051,N_6104);
or U6302 (N_6302,N_6162,N_6187);
and U6303 (N_6303,N_6049,N_6187);
or U6304 (N_6304,N_6168,N_6196);
nor U6305 (N_6305,N_6132,N_6198);
nand U6306 (N_6306,N_6181,N_6068);
xnor U6307 (N_6307,N_6018,N_6105);
nand U6308 (N_6308,N_6162,N_6136);
and U6309 (N_6309,N_6063,N_6048);
and U6310 (N_6310,N_6181,N_6112);
or U6311 (N_6311,N_6187,N_6190);
and U6312 (N_6312,N_6051,N_6002);
and U6313 (N_6313,N_6108,N_6119);
nand U6314 (N_6314,N_6064,N_6046);
xnor U6315 (N_6315,N_6163,N_6082);
and U6316 (N_6316,N_6180,N_6099);
nor U6317 (N_6317,N_6035,N_6142);
and U6318 (N_6318,N_6154,N_6046);
nand U6319 (N_6319,N_6147,N_6041);
nand U6320 (N_6320,N_6129,N_6189);
and U6321 (N_6321,N_6194,N_6145);
and U6322 (N_6322,N_6182,N_6057);
or U6323 (N_6323,N_6022,N_6162);
and U6324 (N_6324,N_6029,N_6122);
nor U6325 (N_6325,N_6098,N_6158);
and U6326 (N_6326,N_6056,N_6091);
and U6327 (N_6327,N_6185,N_6151);
nand U6328 (N_6328,N_6071,N_6146);
nand U6329 (N_6329,N_6065,N_6002);
or U6330 (N_6330,N_6135,N_6150);
or U6331 (N_6331,N_6170,N_6100);
or U6332 (N_6332,N_6064,N_6178);
and U6333 (N_6333,N_6060,N_6033);
xnor U6334 (N_6334,N_6064,N_6056);
xor U6335 (N_6335,N_6119,N_6171);
and U6336 (N_6336,N_6197,N_6075);
nand U6337 (N_6337,N_6029,N_6038);
or U6338 (N_6338,N_6032,N_6183);
and U6339 (N_6339,N_6136,N_6160);
or U6340 (N_6340,N_6121,N_6003);
nand U6341 (N_6341,N_6155,N_6179);
or U6342 (N_6342,N_6183,N_6182);
and U6343 (N_6343,N_6088,N_6070);
and U6344 (N_6344,N_6191,N_6001);
and U6345 (N_6345,N_6049,N_6154);
or U6346 (N_6346,N_6089,N_6036);
nor U6347 (N_6347,N_6163,N_6122);
and U6348 (N_6348,N_6180,N_6021);
and U6349 (N_6349,N_6181,N_6084);
and U6350 (N_6350,N_6120,N_6131);
nor U6351 (N_6351,N_6180,N_6102);
xor U6352 (N_6352,N_6000,N_6144);
xor U6353 (N_6353,N_6192,N_6046);
or U6354 (N_6354,N_6044,N_6099);
nor U6355 (N_6355,N_6035,N_6009);
nor U6356 (N_6356,N_6146,N_6004);
nand U6357 (N_6357,N_6014,N_6129);
nand U6358 (N_6358,N_6194,N_6093);
nand U6359 (N_6359,N_6107,N_6159);
nand U6360 (N_6360,N_6109,N_6163);
and U6361 (N_6361,N_6014,N_6054);
xor U6362 (N_6362,N_6160,N_6106);
xnor U6363 (N_6363,N_6037,N_6052);
xnor U6364 (N_6364,N_6066,N_6026);
and U6365 (N_6365,N_6186,N_6168);
and U6366 (N_6366,N_6068,N_6014);
xnor U6367 (N_6367,N_6109,N_6006);
nand U6368 (N_6368,N_6099,N_6142);
or U6369 (N_6369,N_6095,N_6129);
nor U6370 (N_6370,N_6098,N_6094);
nand U6371 (N_6371,N_6147,N_6169);
nand U6372 (N_6372,N_6051,N_6031);
and U6373 (N_6373,N_6149,N_6155);
nand U6374 (N_6374,N_6111,N_6124);
nand U6375 (N_6375,N_6090,N_6077);
and U6376 (N_6376,N_6058,N_6092);
nand U6377 (N_6377,N_6086,N_6068);
and U6378 (N_6378,N_6156,N_6074);
or U6379 (N_6379,N_6158,N_6150);
and U6380 (N_6380,N_6108,N_6167);
nand U6381 (N_6381,N_6168,N_6106);
xnor U6382 (N_6382,N_6048,N_6011);
xor U6383 (N_6383,N_6169,N_6105);
or U6384 (N_6384,N_6009,N_6195);
nand U6385 (N_6385,N_6142,N_6114);
or U6386 (N_6386,N_6052,N_6196);
or U6387 (N_6387,N_6054,N_6059);
and U6388 (N_6388,N_6048,N_6172);
and U6389 (N_6389,N_6166,N_6118);
nor U6390 (N_6390,N_6085,N_6141);
or U6391 (N_6391,N_6036,N_6047);
nor U6392 (N_6392,N_6110,N_6135);
or U6393 (N_6393,N_6187,N_6194);
nor U6394 (N_6394,N_6125,N_6067);
nor U6395 (N_6395,N_6133,N_6070);
and U6396 (N_6396,N_6056,N_6144);
or U6397 (N_6397,N_6057,N_6093);
nand U6398 (N_6398,N_6113,N_6171);
or U6399 (N_6399,N_6124,N_6161);
and U6400 (N_6400,N_6260,N_6291);
nor U6401 (N_6401,N_6212,N_6205);
nand U6402 (N_6402,N_6374,N_6353);
or U6403 (N_6403,N_6282,N_6362);
or U6404 (N_6404,N_6263,N_6393);
xnor U6405 (N_6405,N_6390,N_6271);
and U6406 (N_6406,N_6342,N_6230);
nor U6407 (N_6407,N_6309,N_6294);
or U6408 (N_6408,N_6376,N_6214);
or U6409 (N_6409,N_6367,N_6299);
nand U6410 (N_6410,N_6217,N_6208);
nand U6411 (N_6411,N_6379,N_6213);
nor U6412 (N_6412,N_6237,N_6224);
or U6413 (N_6413,N_6369,N_6338);
nor U6414 (N_6414,N_6256,N_6312);
xnor U6415 (N_6415,N_6386,N_6301);
nand U6416 (N_6416,N_6226,N_6314);
xnor U6417 (N_6417,N_6281,N_6204);
or U6418 (N_6418,N_6225,N_6356);
or U6419 (N_6419,N_6318,N_6227);
and U6420 (N_6420,N_6372,N_6250);
and U6421 (N_6421,N_6228,N_6262);
nand U6422 (N_6422,N_6245,N_6302);
nand U6423 (N_6423,N_6234,N_6247);
xnor U6424 (N_6424,N_6329,N_6216);
xnor U6425 (N_6425,N_6255,N_6289);
or U6426 (N_6426,N_6220,N_6340);
xor U6427 (N_6427,N_6331,N_6269);
nor U6428 (N_6428,N_6317,N_6239);
and U6429 (N_6429,N_6337,N_6215);
nor U6430 (N_6430,N_6380,N_6360);
nand U6431 (N_6431,N_6257,N_6327);
and U6432 (N_6432,N_6334,N_6378);
and U6433 (N_6433,N_6200,N_6254);
or U6434 (N_6434,N_6259,N_6332);
xnor U6435 (N_6435,N_6206,N_6290);
or U6436 (N_6436,N_6357,N_6298);
nor U6437 (N_6437,N_6354,N_6272);
xor U6438 (N_6438,N_6370,N_6235);
nand U6439 (N_6439,N_6351,N_6313);
and U6440 (N_6440,N_6397,N_6285);
and U6441 (N_6441,N_6373,N_6339);
or U6442 (N_6442,N_6243,N_6365);
and U6443 (N_6443,N_6252,N_6345);
or U6444 (N_6444,N_6201,N_6325);
and U6445 (N_6445,N_6307,N_6296);
nand U6446 (N_6446,N_6276,N_6202);
or U6447 (N_6447,N_6292,N_6388);
or U6448 (N_6448,N_6270,N_6300);
xor U6449 (N_6449,N_6236,N_6371);
and U6450 (N_6450,N_6211,N_6387);
and U6451 (N_6451,N_6203,N_6364);
and U6452 (N_6452,N_6286,N_6368);
or U6453 (N_6453,N_6326,N_6303);
or U6454 (N_6454,N_6207,N_6244);
nor U6455 (N_6455,N_6242,N_6231);
nand U6456 (N_6456,N_6363,N_6383);
and U6457 (N_6457,N_6293,N_6210);
and U6458 (N_6458,N_6350,N_6319);
or U6459 (N_6459,N_6261,N_6359);
or U6460 (N_6460,N_6343,N_6268);
and U6461 (N_6461,N_6229,N_6283);
and U6462 (N_6462,N_6264,N_6391);
xor U6463 (N_6463,N_6223,N_6366);
nand U6464 (N_6464,N_6321,N_6249);
or U6465 (N_6465,N_6241,N_6295);
nand U6466 (N_6466,N_6288,N_6347);
nor U6467 (N_6467,N_6278,N_6346);
nor U6468 (N_6468,N_6248,N_6221);
and U6469 (N_6469,N_6385,N_6381);
or U6470 (N_6470,N_6324,N_6265);
xnor U6471 (N_6471,N_6352,N_6305);
and U6472 (N_6472,N_6219,N_6348);
nand U6473 (N_6473,N_6375,N_6284);
nor U6474 (N_6474,N_6377,N_6209);
xnor U6475 (N_6475,N_6398,N_6389);
nor U6476 (N_6476,N_6341,N_6222);
nand U6477 (N_6477,N_6315,N_6287);
xor U6478 (N_6478,N_6266,N_6258);
nor U6479 (N_6479,N_6280,N_6323);
and U6480 (N_6480,N_6253,N_6399);
and U6481 (N_6481,N_6392,N_6232);
and U6482 (N_6482,N_6218,N_6395);
nand U6483 (N_6483,N_6240,N_6267);
nand U6484 (N_6484,N_6310,N_6306);
nor U6485 (N_6485,N_6335,N_6394);
nor U6486 (N_6486,N_6251,N_6246);
xor U6487 (N_6487,N_6396,N_6328);
and U6488 (N_6488,N_6355,N_6382);
nand U6489 (N_6489,N_6304,N_6279);
and U6490 (N_6490,N_6297,N_6274);
and U6491 (N_6491,N_6275,N_6361);
or U6492 (N_6492,N_6384,N_6316);
and U6493 (N_6493,N_6273,N_6358);
nor U6494 (N_6494,N_6336,N_6277);
and U6495 (N_6495,N_6311,N_6238);
or U6496 (N_6496,N_6344,N_6308);
nor U6497 (N_6497,N_6322,N_6333);
and U6498 (N_6498,N_6320,N_6349);
nand U6499 (N_6499,N_6330,N_6233);
nand U6500 (N_6500,N_6318,N_6200);
or U6501 (N_6501,N_6325,N_6252);
or U6502 (N_6502,N_6378,N_6264);
or U6503 (N_6503,N_6206,N_6215);
or U6504 (N_6504,N_6393,N_6290);
and U6505 (N_6505,N_6397,N_6348);
or U6506 (N_6506,N_6261,N_6357);
nand U6507 (N_6507,N_6305,N_6327);
nand U6508 (N_6508,N_6278,N_6226);
and U6509 (N_6509,N_6290,N_6395);
xnor U6510 (N_6510,N_6265,N_6358);
xor U6511 (N_6511,N_6342,N_6356);
or U6512 (N_6512,N_6361,N_6345);
nand U6513 (N_6513,N_6231,N_6308);
or U6514 (N_6514,N_6361,N_6396);
nor U6515 (N_6515,N_6267,N_6311);
and U6516 (N_6516,N_6223,N_6313);
xnor U6517 (N_6517,N_6278,N_6289);
or U6518 (N_6518,N_6290,N_6242);
nor U6519 (N_6519,N_6352,N_6391);
xnor U6520 (N_6520,N_6312,N_6259);
xnor U6521 (N_6521,N_6272,N_6314);
nor U6522 (N_6522,N_6206,N_6284);
nor U6523 (N_6523,N_6381,N_6220);
xnor U6524 (N_6524,N_6367,N_6326);
nor U6525 (N_6525,N_6299,N_6301);
xnor U6526 (N_6526,N_6246,N_6226);
nor U6527 (N_6527,N_6237,N_6385);
nor U6528 (N_6528,N_6298,N_6296);
xnor U6529 (N_6529,N_6297,N_6232);
nand U6530 (N_6530,N_6251,N_6346);
nor U6531 (N_6531,N_6372,N_6262);
or U6532 (N_6532,N_6324,N_6270);
nor U6533 (N_6533,N_6341,N_6288);
or U6534 (N_6534,N_6277,N_6275);
and U6535 (N_6535,N_6302,N_6293);
nor U6536 (N_6536,N_6228,N_6393);
xor U6537 (N_6537,N_6360,N_6255);
nand U6538 (N_6538,N_6227,N_6361);
nand U6539 (N_6539,N_6379,N_6373);
nor U6540 (N_6540,N_6309,N_6271);
and U6541 (N_6541,N_6229,N_6236);
xnor U6542 (N_6542,N_6267,N_6373);
and U6543 (N_6543,N_6344,N_6362);
xor U6544 (N_6544,N_6397,N_6312);
nand U6545 (N_6545,N_6388,N_6350);
or U6546 (N_6546,N_6312,N_6337);
or U6547 (N_6547,N_6359,N_6230);
nor U6548 (N_6548,N_6224,N_6322);
or U6549 (N_6549,N_6321,N_6377);
or U6550 (N_6550,N_6234,N_6364);
or U6551 (N_6551,N_6326,N_6252);
nor U6552 (N_6552,N_6343,N_6233);
and U6553 (N_6553,N_6253,N_6318);
xor U6554 (N_6554,N_6349,N_6292);
xor U6555 (N_6555,N_6276,N_6277);
xnor U6556 (N_6556,N_6215,N_6311);
and U6557 (N_6557,N_6270,N_6283);
nand U6558 (N_6558,N_6201,N_6334);
and U6559 (N_6559,N_6215,N_6288);
nand U6560 (N_6560,N_6327,N_6330);
and U6561 (N_6561,N_6329,N_6372);
or U6562 (N_6562,N_6220,N_6319);
xnor U6563 (N_6563,N_6323,N_6200);
nand U6564 (N_6564,N_6379,N_6292);
nand U6565 (N_6565,N_6371,N_6394);
nand U6566 (N_6566,N_6293,N_6386);
nand U6567 (N_6567,N_6261,N_6275);
nand U6568 (N_6568,N_6338,N_6210);
nand U6569 (N_6569,N_6215,N_6229);
nand U6570 (N_6570,N_6226,N_6352);
nand U6571 (N_6571,N_6366,N_6302);
nor U6572 (N_6572,N_6265,N_6371);
or U6573 (N_6573,N_6221,N_6258);
or U6574 (N_6574,N_6213,N_6259);
or U6575 (N_6575,N_6383,N_6296);
nor U6576 (N_6576,N_6250,N_6342);
nand U6577 (N_6577,N_6287,N_6212);
and U6578 (N_6578,N_6392,N_6288);
xor U6579 (N_6579,N_6372,N_6278);
nor U6580 (N_6580,N_6206,N_6321);
or U6581 (N_6581,N_6317,N_6251);
nand U6582 (N_6582,N_6272,N_6342);
nand U6583 (N_6583,N_6355,N_6306);
and U6584 (N_6584,N_6337,N_6225);
nor U6585 (N_6585,N_6242,N_6332);
nor U6586 (N_6586,N_6396,N_6300);
or U6587 (N_6587,N_6208,N_6210);
xnor U6588 (N_6588,N_6238,N_6204);
and U6589 (N_6589,N_6336,N_6325);
and U6590 (N_6590,N_6222,N_6396);
nor U6591 (N_6591,N_6303,N_6283);
or U6592 (N_6592,N_6288,N_6251);
or U6593 (N_6593,N_6332,N_6328);
or U6594 (N_6594,N_6392,N_6262);
nor U6595 (N_6595,N_6344,N_6300);
nor U6596 (N_6596,N_6372,N_6214);
and U6597 (N_6597,N_6354,N_6319);
nor U6598 (N_6598,N_6333,N_6291);
nor U6599 (N_6599,N_6300,N_6384);
xnor U6600 (N_6600,N_6445,N_6497);
and U6601 (N_6601,N_6432,N_6558);
xnor U6602 (N_6602,N_6591,N_6502);
nand U6603 (N_6603,N_6403,N_6508);
and U6604 (N_6604,N_6536,N_6420);
or U6605 (N_6605,N_6427,N_6486);
and U6606 (N_6606,N_6480,N_6550);
and U6607 (N_6607,N_6491,N_6423);
xnor U6608 (N_6608,N_6442,N_6462);
nand U6609 (N_6609,N_6541,N_6481);
xor U6610 (N_6610,N_6566,N_6493);
nor U6611 (N_6611,N_6496,N_6531);
nor U6612 (N_6612,N_6511,N_6469);
nand U6613 (N_6613,N_6452,N_6464);
nand U6614 (N_6614,N_6586,N_6440);
nand U6615 (N_6615,N_6507,N_6556);
xnor U6616 (N_6616,N_6447,N_6585);
nand U6617 (N_6617,N_6484,N_6488);
nand U6618 (N_6618,N_6411,N_6574);
nand U6619 (N_6619,N_6404,N_6520);
or U6620 (N_6620,N_6562,N_6425);
or U6621 (N_6621,N_6451,N_6407);
nand U6622 (N_6622,N_6551,N_6519);
nor U6623 (N_6623,N_6448,N_6533);
and U6624 (N_6624,N_6571,N_6514);
nor U6625 (N_6625,N_6592,N_6593);
or U6626 (N_6626,N_6572,N_6466);
and U6627 (N_6627,N_6526,N_6437);
nand U6628 (N_6628,N_6553,N_6573);
and U6629 (N_6629,N_6544,N_6475);
xnor U6630 (N_6630,N_6455,N_6421);
or U6631 (N_6631,N_6577,N_6471);
or U6632 (N_6632,N_6402,N_6564);
nor U6633 (N_6633,N_6428,N_6569);
nor U6634 (N_6634,N_6545,N_6515);
and U6635 (N_6635,N_6501,N_6561);
and U6636 (N_6636,N_6408,N_6542);
nor U6637 (N_6637,N_6430,N_6513);
xnor U6638 (N_6638,N_6560,N_6482);
xnor U6639 (N_6639,N_6559,N_6595);
or U6640 (N_6640,N_6467,N_6458);
or U6641 (N_6641,N_6443,N_6468);
xor U6642 (N_6642,N_6450,N_6419);
or U6643 (N_6643,N_6581,N_6500);
nor U6644 (N_6644,N_6476,N_6439);
and U6645 (N_6645,N_6433,N_6446);
xnor U6646 (N_6646,N_6539,N_6512);
nor U6647 (N_6647,N_6473,N_6552);
xor U6648 (N_6648,N_6495,N_6405);
or U6649 (N_6649,N_6406,N_6540);
or U6650 (N_6650,N_6567,N_6456);
xnor U6651 (N_6651,N_6416,N_6400);
nor U6652 (N_6652,N_6457,N_6530);
nand U6653 (N_6653,N_6584,N_6477);
nand U6654 (N_6654,N_6463,N_6534);
or U6655 (N_6655,N_6459,N_6521);
nor U6656 (N_6656,N_6529,N_6516);
or U6657 (N_6657,N_6576,N_6554);
or U6658 (N_6658,N_6583,N_6532);
or U6659 (N_6659,N_6537,N_6460);
and U6660 (N_6660,N_6453,N_6409);
xor U6661 (N_6661,N_6412,N_6589);
xor U6662 (N_6662,N_6543,N_6429);
nor U6663 (N_6663,N_6506,N_6503);
and U6664 (N_6664,N_6401,N_6413);
or U6665 (N_6665,N_6461,N_6523);
and U6666 (N_6666,N_6546,N_6441);
or U6667 (N_6667,N_6597,N_6575);
xor U6668 (N_6668,N_6528,N_6565);
nand U6669 (N_6669,N_6417,N_6570);
and U6670 (N_6670,N_6489,N_6596);
and U6671 (N_6671,N_6494,N_6548);
nor U6672 (N_6672,N_6431,N_6580);
or U6673 (N_6673,N_6435,N_6599);
nand U6674 (N_6674,N_6434,N_6465);
or U6675 (N_6675,N_6444,N_6479);
nand U6676 (N_6676,N_6522,N_6492);
nor U6677 (N_6677,N_6509,N_6504);
xor U6678 (N_6678,N_6594,N_6418);
and U6679 (N_6679,N_6490,N_6499);
or U6680 (N_6680,N_6414,N_6535);
nor U6681 (N_6681,N_6487,N_6505);
xnor U6682 (N_6682,N_6470,N_6510);
nand U6683 (N_6683,N_6582,N_6587);
and U6684 (N_6684,N_6598,N_6527);
or U6685 (N_6685,N_6525,N_6579);
xnor U6686 (N_6686,N_6563,N_6557);
xnor U6687 (N_6687,N_6588,N_6410);
nor U6688 (N_6688,N_6426,N_6472);
nand U6689 (N_6689,N_6547,N_6498);
or U6690 (N_6690,N_6549,N_6568);
xnor U6691 (N_6691,N_6422,N_6517);
xnor U6692 (N_6692,N_6449,N_6415);
xor U6693 (N_6693,N_6474,N_6578);
xnor U6694 (N_6694,N_6454,N_6538);
nor U6695 (N_6695,N_6436,N_6478);
or U6696 (N_6696,N_6555,N_6524);
or U6697 (N_6697,N_6483,N_6518);
xnor U6698 (N_6698,N_6424,N_6485);
nor U6699 (N_6699,N_6438,N_6590);
nand U6700 (N_6700,N_6571,N_6599);
and U6701 (N_6701,N_6426,N_6489);
or U6702 (N_6702,N_6511,N_6596);
and U6703 (N_6703,N_6547,N_6533);
and U6704 (N_6704,N_6511,N_6493);
and U6705 (N_6705,N_6445,N_6471);
and U6706 (N_6706,N_6596,N_6543);
or U6707 (N_6707,N_6535,N_6476);
or U6708 (N_6708,N_6571,N_6493);
xor U6709 (N_6709,N_6526,N_6454);
or U6710 (N_6710,N_6535,N_6420);
or U6711 (N_6711,N_6598,N_6438);
nand U6712 (N_6712,N_6432,N_6407);
or U6713 (N_6713,N_6506,N_6452);
nand U6714 (N_6714,N_6590,N_6497);
xnor U6715 (N_6715,N_6570,N_6459);
nand U6716 (N_6716,N_6484,N_6523);
nand U6717 (N_6717,N_6418,N_6559);
xor U6718 (N_6718,N_6504,N_6490);
nand U6719 (N_6719,N_6559,N_6503);
xor U6720 (N_6720,N_6419,N_6507);
and U6721 (N_6721,N_6514,N_6540);
xor U6722 (N_6722,N_6406,N_6466);
nand U6723 (N_6723,N_6462,N_6412);
or U6724 (N_6724,N_6561,N_6482);
nand U6725 (N_6725,N_6591,N_6415);
and U6726 (N_6726,N_6595,N_6412);
or U6727 (N_6727,N_6509,N_6572);
or U6728 (N_6728,N_6543,N_6485);
xnor U6729 (N_6729,N_6585,N_6570);
and U6730 (N_6730,N_6520,N_6455);
nand U6731 (N_6731,N_6455,N_6442);
or U6732 (N_6732,N_6477,N_6558);
nor U6733 (N_6733,N_6490,N_6588);
nand U6734 (N_6734,N_6538,N_6483);
nand U6735 (N_6735,N_6564,N_6562);
xnor U6736 (N_6736,N_6538,N_6529);
and U6737 (N_6737,N_6446,N_6486);
nand U6738 (N_6738,N_6470,N_6425);
and U6739 (N_6739,N_6407,N_6463);
xnor U6740 (N_6740,N_6482,N_6430);
nor U6741 (N_6741,N_6580,N_6540);
nor U6742 (N_6742,N_6406,N_6439);
xnor U6743 (N_6743,N_6518,N_6580);
or U6744 (N_6744,N_6580,N_6573);
nor U6745 (N_6745,N_6472,N_6444);
nor U6746 (N_6746,N_6426,N_6474);
or U6747 (N_6747,N_6492,N_6464);
xnor U6748 (N_6748,N_6597,N_6591);
nor U6749 (N_6749,N_6441,N_6511);
nor U6750 (N_6750,N_6431,N_6414);
and U6751 (N_6751,N_6534,N_6510);
nand U6752 (N_6752,N_6495,N_6475);
nand U6753 (N_6753,N_6463,N_6485);
xnor U6754 (N_6754,N_6514,N_6497);
nand U6755 (N_6755,N_6411,N_6521);
nor U6756 (N_6756,N_6530,N_6452);
xor U6757 (N_6757,N_6404,N_6540);
xnor U6758 (N_6758,N_6524,N_6596);
xnor U6759 (N_6759,N_6567,N_6467);
nand U6760 (N_6760,N_6417,N_6562);
and U6761 (N_6761,N_6548,N_6465);
and U6762 (N_6762,N_6416,N_6519);
nand U6763 (N_6763,N_6546,N_6592);
xor U6764 (N_6764,N_6560,N_6509);
nor U6765 (N_6765,N_6459,N_6528);
or U6766 (N_6766,N_6592,N_6568);
or U6767 (N_6767,N_6448,N_6407);
nor U6768 (N_6768,N_6408,N_6456);
nor U6769 (N_6769,N_6457,N_6489);
and U6770 (N_6770,N_6443,N_6499);
nand U6771 (N_6771,N_6548,N_6424);
nand U6772 (N_6772,N_6503,N_6465);
or U6773 (N_6773,N_6410,N_6486);
and U6774 (N_6774,N_6520,N_6427);
and U6775 (N_6775,N_6548,N_6438);
nand U6776 (N_6776,N_6446,N_6414);
xor U6777 (N_6777,N_6442,N_6436);
and U6778 (N_6778,N_6584,N_6570);
or U6779 (N_6779,N_6504,N_6545);
nand U6780 (N_6780,N_6401,N_6538);
nand U6781 (N_6781,N_6562,N_6419);
or U6782 (N_6782,N_6492,N_6513);
nand U6783 (N_6783,N_6573,N_6458);
and U6784 (N_6784,N_6499,N_6471);
nand U6785 (N_6785,N_6574,N_6589);
xnor U6786 (N_6786,N_6568,N_6406);
nor U6787 (N_6787,N_6439,N_6407);
xnor U6788 (N_6788,N_6505,N_6465);
and U6789 (N_6789,N_6588,N_6435);
xnor U6790 (N_6790,N_6511,N_6595);
nor U6791 (N_6791,N_6541,N_6529);
or U6792 (N_6792,N_6483,N_6593);
and U6793 (N_6793,N_6528,N_6560);
and U6794 (N_6794,N_6554,N_6477);
nand U6795 (N_6795,N_6531,N_6440);
nor U6796 (N_6796,N_6525,N_6541);
nor U6797 (N_6797,N_6593,N_6563);
or U6798 (N_6798,N_6412,N_6588);
xor U6799 (N_6799,N_6544,N_6511);
or U6800 (N_6800,N_6728,N_6604);
nor U6801 (N_6801,N_6648,N_6724);
or U6802 (N_6802,N_6759,N_6686);
nor U6803 (N_6803,N_6627,N_6650);
xor U6804 (N_6804,N_6755,N_6729);
or U6805 (N_6805,N_6721,N_6771);
and U6806 (N_6806,N_6754,N_6747);
or U6807 (N_6807,N_6725,N_6688);
nand U6808 (N_6808,N_6766,N_6681);
xor U6809 (N_6809,N_6668,N_6750);
nor U6810 (N_6810,N_6619,N_6740);
nor U6811 (N_6811,N_6675,N_6794);
nand U6812 (N_6812,N_6608,N_6779);
nand U6813 (N_6813,N_6757,N_6611);
nor U6814 (N_6814,N_6605,N_6601);
and U6815 (N_6815,N_6705,N_6761);
xor U6816 (N_6816,N_6723,N_6791);
and U6817 (N_6817,N_6635,N_6719);
or U6818 (N_6818,N_6707,N_6752);
or U6819 (N_6819,N_6777,N_6600);
nor U6820 (N_6820,N_6692,N_6776);
xor U6821 (N_6821,N_6796,N_6620);
or U6822 (N_6822,N_6789,N_6768);
nand U6823 (N_6823,N_6758,N_6733);
nor U6824 (N_6824,N_6615,N_6653);
and U6825 (N_6825,N_6712,N_6775);
xnor U6826 (N_6826,N_6745,N_6661);
or U6827 (N_6827,N_6782,N_6624);
nor U6828 (N_6828,N_6737,N_6645);
xnor U6829 (N_6829,N_6690,N_6603);
or U6830 (N_6830,N_6710,N_6708);
xor U6831 (N_6831,N_6676,N_6765);
or U6832 (N_6832,N_6764,N_6787);
or U6833 (N_6833,N_6660,N_6785);
xor U6834 (N_6834,N_6684,N_6669);
nor U6835 (N_6835,N_6781,N_6727);
nor U6836 (N_6836,N_6683,N_6795);
or U6837 (N_6837,N_6746,N_6762);
and U6838 (N_6838,N_6659,N_6770);
or U6839 (N_6839,N_6632,N_6639);
or U6840 (N_6840,N_6691,N_6689);
and U6841 (N_6841,N_6741,N_6749);
xor U6842 (N_6842,N_6631,N_6714);
nand U6843 (N_6843,N_6778,N_6665);
nor U6844 (N_6844,N_6700,N_6701);
or U6845 (N_6845,N_6732,N_6628);
or U6846 (N_6846,N_6662,N_6621);
xor U6847 (N_6847,N_6695,N_6610);
xor U6848 (N_6848,N_6647,N_6713);
xnor U6849 (N_6849,N_6606,N_6679);
xor U6850 (N_6850,N_6703,N_6636);
or U6851 (N_6851,N_6790,N_6784);
nand U6852 (N_6852,N_6641,N_6706);
nor U6853 (N_6853,N_6715,N_6651);
nand U6854 (N_6854,N_6649,N_6670);
nand U6855 (N_6855,N_6682,N_6613);
and U6856 (N_6856,N_6646,N_6637);
and U6857 (N_6857,N_6704,N_6699);
nand U6858 (N_6858,N_6602,N_6722);
and U6859 (N_6859,N_6638,N_6718);
nor U6860 (N_6860,N_6677,N_6630);
xor U6861 (N_6861,N_6633,N_6634);
or U6862 (N_6862,N_6616,N_6748);
and U6863 (N_6863,N_6663,N_6751);
and U6864 (N_6864,N_6742,N_6717);
nand U6865 (N_6865,N_6618,N_6622);
and U6866 (N_6866,N_6756,N_6797);
nand U6867 (N_6867,N_6774,N_6736);
or U6868 (N_6868,N_6799,N_6786);
or U6869 (N_6869,N_6671,N_6738);
nor U6870 (N_6870,N_6726,N_6617);
xor U6871 (N_6871,N_6698,N_6734);
nor U6872 (N_6872,N_6730,N_6644);
xnor U6873 (N_6873,N_6694,N_6760);
nor U6874 (N_6874,N_6609,N_6793);
nand U6875 (N_6875,N_6652,N_6769);
xor U6876 (N_6876,N_6623,N_6739);
xnor U6877 (N_6877,N_6674,N_6625);
nand U6878 (N_6878,N_6735,N_6685);
xnor U6879 (N_6879,N_6687,N_6607);
and U6880 (N_6880,N_6743,N_6798);
and U6881 (N_6881,N_6763,N_6697);
nand U6882 (N_6882,N_6753,N_6744);
nand U6883 (N_6883,N_6666,N_6664);
nand U6884 (N_6884,N_6678,N_6672);
nand U6885 (N_6885,N_6626,N_6788);
and U6886 (N_6886,N_6640,N_6792);
nand U6887 (N_6887,N_6783,N_6693);
or U6888 (N_6888,N_6673,N_6780);
xnor U6889 (N_6889,N_6656,N_6614);
nand U6890 (N_6890,N_6709,N_6657);
and U6891 (N_6891,N_6767,N_6654);
nor U6892 (N_6892,N_6773,N_6667);
nor U6893 (N_6893,N_6655,N_6612);
or U6894 (N_6894,N_6702,N_6642);
xnor U6895 (N_6895,N_6680,N_6720);
or U6896 (N_6896,N_6772,N_6716);
or U6897 (N_6897,N_6696,N_6711);
nand U6898 (N_6898,N_6643,N_6658);
nor U6899 (N_6899,N_6629,N_6731);
and U6900 (N_6900,N_6717,N_6636);
xnor U6901 (N_6901,N_6772,N_6732);
nor U6902 (N_6902,N_6657,N_6796);
or U6903 (N_6903,N_6776,N_6785);
or U6904 (N_6904,N_6743,N_6759);
nand U6905 (N_6905,N_6762,N_6614);
and U6906 (N_6906,N_6675,N_6761);
and U6907 (N_6907,N_6678,N_6713);
nand U6908 (N_6908,N_6682,N_6678);
xnor U6909 (N_6909,N_6777,N_6694);
and U6910 (N_6910,N_6754,N_6614);
xnor U6911 (N_6911,N_6613,N_6620);
nor U6912 (N_6912,N_6621,N_6677);
nand U6913 (N_6913,N_6720,N_6633);
and U6914 (N_6914,N_6712,N_6707);
or U6915 (N_6915,N_6782,N_6676);
nor U6916 (N_6916,N_6779,N_6759);
xnor U6917 (N_6917,N_6699,N_6642);
and U6918 (N_6918,N_6736,N_6757);
xor U6919 (N_6919,N_6739,N_6610);
xnor U6920 (N_6920,N_6679,N_6708);
and U6921 (N_6921,N_6790,N_6752);
and U6922 (N_6922,N_6770,N_6631);
or U6923 (N_6923,N_6799,N_6728);
and U6924 (N_6924,N_6696,N_6714);
or U6925 (N_6925,N_6688,N_6656);
or U6926 (N_6926,N_6655,N_6634);
xor U6927 (N_6927,N_6795,N_6771);
and U6928 (N_6928,N_6667,N_6723);
and U6929 (N_6929,N_6652,N_6763);
or U6930 (N_6930,N_6649,N_6745);
xor U6931 (N_6931,N_6737,N_6760);
xnor U6932 (N_6932,N_6767,N_6714);
xor U6933 (N_6933,N_6782,N_6621);
nand U6934 (N_6934,N_6693,N_6646);
nor U6935 (N_6935,N_6735,N_6665);
and U6936 (N_6936,N_6780,N_6789);
and U6937 (N_6937,N_6740,N_6689);
nand U6938 (N_6938,N_6727,N_6670);
nor U6939 (N_6939,N_6652,N_6635);
and U6940 (N_6940,N_6777,N_6715);
xnor U6941 (N_6941,N_6751,N_6620);
and U6942 (N_6942,N_6655,N_6789);
nand U6943 (N_6943,N_6649,N_6606);
nand U6944 (N_6944,N_6753,N_6614);
and U6945 (N_6945,N_6785,N_6677);
nand U6946 (N_6946,N_6765,N_6729);
or U6947 (N_6947,N_6620,N_6722);
xnor U6948 (N_6948,N_6697,N_6660);
or U6949 (N_6949,N_6716,N_6770);
xnor U6950 (N_6950,N_6791,N_6693);
xnor U6951 (N_6951,N_6722,N_6713);
nand U6952 (N_6952,N_6722,N_6718);
xor U6953 (N_6953,N_6766,N_6724);
nor U6954 (N_6954,N_6744,N_6661);
or U6955 (N_6955,N_6680,N_6719);
and U6956 (N_6956,N_6624,N_6739);
nor U6957 (N_6957,N_6654,N_6620);
and U6958 (N_6958,N_6709,N_6618);
nand U6959 (N_6959,N_6666,N_6633);
and U6960 (N_6960,N_6669,N_6721);
or U6961 (N_6961,N_6633,N_6704);
nor U6962 (N_6962,N_6791,N_6777);
nor U6963 (N_6963,N_6758,N_6610);
and U6964 (N_6964,N_6728,N_6628);
nand U6965 (N_6965,N_6790,N_6690);
and U6966 (N_6966,N_6605,N_6789);
or U6967 (N_6967,N_6619,N_6629);
nor U6968 (N_6968,N_6632,N_6745);
nor U6969 (N_6969,N_6627,N_6624);
nor U6970 (N_6970,N_6751,N_6742);
nand U6971 (N_6971,N_6724,N_6705);
nand U6972 (N_6972,N_6784,N_6702);
nor U6973 (N_6973,N_6712,N_6764);
nor U6974 (N_6974,N_6726,N_6715);
or U6975 (N_6975,N_6776,N_6749);
and U6976 (N_6976,N_6620,N_6720);
xor U6977 (N_6977,N_6653,N_6646);
or U6978 (N_6978,N_6671,N_6775);
and U6979 (N_6979,N_6700,N_6747);
nand U6980 (N_6980,N_6702,N_6754);
nor U6981 (N_6981,N_6736,N_6765);
or U6982 (N_6982,N_6736,N_6712);
nand U6983 (N_6983,N_6721,N_6711);
and U6984 (N_6984,N_6733,N_6644);
nand U6985 (N_6985,N_6678,N_6714);
nor U6986 (N_6986,N_6780,N_6647);
nand U6987 (N_6987,N_6646,N_6600);
nand U6988 (N_6988,N_6614,N_6636);
nor U6989 (N_6989,N_6609,N_6681);
nor U6990 (N_6990,N_6623,N_6768);
and U6991 (N_6991,N_6665,N_6635);
xor U6992 (N_6992,N_6608,N_6731);
nand U6993 (N_6993,N_6630,N_6717);
and U6994 (N_6994,N_6715,N_6637);
nor U6995 (N_6995,N_6668,N_6687);
nor U6996 (N_6996,N_6782,N_6732);
xor U6997 (N_6997,N_6609,N_6699);
xnor U6998 (N_6998,N_6707,N_6652);
nand U6999 (N_6999,N_6660,N_6747);
nand U7000 (N_7000,N_6813,N_6825);
or U7001 (N_7001,N_6915,N_6856);
or U7002 (N_7002,N_6945,N_6952);
nor U7003 (N_7003,N_6883,N_6843);
xnor U7004 (N_7004,N_6900,N_6949);
or U7005 (N_7005,N_6906,N_6999);
xor U7006 (N_7006,N_6975,N_6817);
xor U7007 (N_7007,N_6888,N_6814);
and U7008 (N_7008,N_6840,N_6966);
nand U7009 (N_7009,N_6917,N_6935);
and U7010 (N_7010,N_6991,N_6996);
nor U7011 (N_7011,N_6943,N_6875);
and U7012 (N_7012,N_6844,N_6861);
and U7013 (N_7013,N_6842,N_6918);
nor U7014 (N_7014,N_6832,N_6908);
or U7015 (N_7015,N_6939,N_6811);
and U7016 (N_7016,N_6971,N_6909);
and U7017 (N_7017,N_6839,N_6870);
nand U7018 (N_7018,N_6893,N_6951);
and U7019 (N_7019,N_6889,N_6863);
xor U7020 (N_7020,N_6987,N_6988);
and U7021 (N_7021,N_6855,N_6852);
nand U7022 (N_7022,N_6983,N_6926);
and U7023 (N_7023,N_6884,N_6807);
nand U7024 (N_7024,N_6824,N_6910);
or U7025 (N_7025,N_6836,N_6891);
and U7026 (N_7026,N_6895,N_6904);
xor U7027 (N_7027,N_6897,N_6853);
or U7028 (N_7028,N_6850,N_6815);
nand U7029 (N_7029,N_6820,N_6858);
nor U7030 (N_7030,N_6961,N_6970);
nor U7031 (N_7031,N_6886,N_6930);
or U7032 (N_7032,N_6955,N_6865);
or U7033 (N_7033,N_6985,N_6879);
nor U7034 (N_7034,N_6907,N_6911);
and U7035 (N_7035,N_6928,N_6986);
or U7036 (N_7036,N_6809,N_6989);
nand U7037 (N_7037,N_6916,N_6838);
or U7038 (N_7038,N_6882,N_6976);
nand U7039 (N_7039,N_6880,N_6803);
nand U7040 (N_7040,N_6956,N_6934);
and U7041 (N_7041,N_6959,N_6936);
xor U7042 (N_7042,N_6835,N_6912);
nand U7043 (N_7043,N_6969,N_6849);
xor U7044 (N_7044,N_6847,N_6854);
nand U7045 (N_7045,N_6867,N_6829);
nor U7046 (N_7046,N_6833,N_6892);
nor U7047 (N_7047,N_6823,N_6885);
xor U7048 (N_7048,N_6804,N_6924);
xnor U7049 (N_7049,N_6837,N_6890);
and U7050 (N_7050,N_6920,N_6972);
or U7051 (N_7051,N_6998,N_6967);
xor U7052 (N_7052,N_6800,N_6913);
nand U7053 (N_7053,N_6876,N_6927);
nor U7054 (N_7054,N_6995,N_6974);
and U7055 (N_7055,N_6905,N_6874);
xor U7056 (N_7056,N_6933,N_6873);
nor U7057 (N_7057,N_6831,N_6957);
or U7058 (N_7058,N_6954,N_6947);
xor U7059 (N_7059,N_6848,N_6931);
or U7060 (N_7060,N_6919,N_6962);
nor U7061 (N_7061,N_6950,N_6818);
xnor U7062 (N_7062,N_6810,N_6960);
nand U7063 (N_7063,N_6846,N_6929);
nand U7064 (N_7064,N_6860,N_6946);
xnor U7065 (N_7065,N_6982,N_6953);
xor U7066 (N_7066,N_6997,N_6802);
and U7067 (N_7067,N_6921,N_6973);
nor U7068 (N_7068,N_6979,N_6830);
or U7069 (N_7069,N_6990,N_6964);
and U7070 (N_7070,N_6941,N_6822);
nor U7071 (N_7071,N_6925,N_6896);
xnor U7072 (N_7072,N_6980,N_6828);
nand U7073 (N_7073,N_6898,N_6805);
or U7074 (N_7074,N_6940,N_6922);
and U7075 (N_7075,N_6887,N_6994);
xor U7076 (N_7076,N_6944,N_6826);
nand U7077 (N_7077,N_6866,N_6821);
and U7078 (N_7078,N_6965,N_6871);
nor U7079 (N_7079,N_6992,N_6978);
and U7080 (N_7080,N_6902,N_6932);
or U7081 (N_7081,N_6948,N_6834);
xor U7082 (N_7082,N_6819,N_6937);
xor U7083 (N_7083,N_6963,N_6993);
and U7084 (N_7084,N_6872,N_6923);
nor U7085 (N_7085,N_6845,N_6808);
nand U7086 (N_7086,N_6806,N_6851);
and U7087 (N_7087,N_6812,N_6857);
nor U7088 (N_7088,N_6899,N_6869);
and U7089 (N_7089,N_6859,N_6914);
xnor U7090 (N_7090,N_6938,N_6958);
nor U7091 (N_7091,N_6968,N_6841);
nand U7092 (N_7092,N_6801,N_6977);
nor U7093 (N_7093,N_6877,N_6878);
and U7094 (N_7094,N_6903,N_6868);
nor U7095 (N_7095,N_6901,N_6981);
or U7096 (N_7096,N_6816,N_6894);
nand U7097 (N_7097,N_6827,N_6984);
nand U7098 (N_7098,N_6864,N_6862);
or U7099 (N_7099,N_6881,N_6942);
nor U7100 (N_7100,N_6851,N_6971);
or U7101 (N_7101,N_6920,N_6863);
xor U7102 (N_7102,N_6942,N_6924);
nor U7103 (N_7103,N_6929,N_6965);
nand U7104 (N_7104,N_6992,N_6812);
nand U7105 (N_7105,N_6940,N_6870);
nand U7106 (N_7106,N_6810,N_6973);
or U7107 (N_7107,N_6801,N_6853);
nand U7108 (N_7108,N_6946,N_6881);
nand U7109 (N_7109,N_6927,N_6904);
and U7110 (N_7110,N_6888,N_6970);
and U7111 (N_7111,N_6893,N_6902);
or U7112 (N_7112,N_6809,N_6914);
xnor U7113 (N_7113,N_6992,N_6875);
or U7114 (N_7114,N_6947,N_6846);
nand U7115 (N_7115,N_6846,N_6942);
or U7116 (N_7116,N_6874,N_6846);
nor U7117 (N_7117,N_6801,N_6866);
or U7118 (N_7118,N_6955,N_6874);
xnor U7119 (N_7119,N_6931,N_6843);
nor U7120 (N_7120,N_6951,N_6997);
and U7121 (N_7121,N_6864,N_6942);
xnor U7122 (N_7122,N_6988,N_6978);
nor U7123 (N_7123,N_6906,N_6991);
and U7124 (N_7124,N_6890,N_6961);
xnor U7125 (N_7125,N_6948,N_6932);
xnor U7126 (N_7126,N_6987,N_6938);
nor U7127 (N_7127,N_6800,N_6834);
or U7128 (N_7128,N_6823,N_6914);
nand U7129 (N_7129,N_6871,N_6843);
and U7130 (N_7130,N_6867,N_6833);
or U7131 (N_7131,N_6900,N_6948);
xor U7132 (N_7132,N_6825,N_6963);
or U7133 (N_7133,N_6843,N_6829);
nand U7134 (N_7134,N_6889,N_6845);
xnor U7135 (N_7135,N_6954,N_6813);
and U7136 (N_7136,N_6932,N_6921);
nor U7137 (N_7137,N_6903,N_6837);
nor U7138 (N_7138,N_6952,N_6946);
nand U7139 (N_7139,N_6926,N_6974);
and U7140 (N_7140,N_6883,N_6818);
nand U7141 (N_7141,N_6911,N_6994);
nand U7142 (N_7142,N_6981,N_6974);
xnor U7143 (N_7143,N_6803,N_6865);
xor U7144 (N_7144,N_6999,N_6994);
xor U7145 (N_7145,N_6939,N_6853);
nor U7146 (N_7146,N_6946,N_6979);
xor U7147 (N_7147,N_6992,N_6826);
or U7148 (N_7148,N_6995,N_6989);
nor U7149 (N_7149,N_6801,N_6858);
or U7150 (N_7150,N_6908,N_6911);
nand U7151 (N_7151,N_6802,N_6929);
and U7152 (N_7152,N_6802,N_6953);
xnor U7153 (N_7153,N_6899,N_6938);
xnor U7154 (N_7154,N_6938,N_6996);
or U7155 (N_7155,N_6878,N_6887);
nand U7156 (N_7156,N_6919,N_6986);
and U7157 (N_7157,N_6847,N_6978);
nand U7158 (N_7158,N_6849,N_6981);
or U7159 (N_7159,N_6919,N_6988);
xor U7160 (N_7160,N_6894,N_6930);
and U7161 (N_7161,N_6865,N_6984);
and U7162 (N_7162,N_6937,N_6836);
xnor U7163 (N_7163,N_6836,N_6815);
and U7164 (N_7164,N_6862,N_6917);
xor U7165 (N_7165,N_6897,N_6869);
xnor U7166 (N_7166,N_6915,N_6962);
nand U7167 (N_7167,N_6870,N_6847);
nand U7168 (N_7168,N_6845,N_6965);
and U7169 (N_7169,N_6983,N_6855);
nor U7170 (N_7170,N_6836,N_6966);
and U7171 (N_7171,N_6855,N_6868);
nor U7172 (N_7172,N_6822,N_6816);
and U7173 (N_7173,N_6980,N_6877);
and U7174 (N_7174,N_6968,N_6813);
and U7175 (N_7175,N_6816,N_6955);
or U7176 (N_7176,N_6897,N_6953);
or U7177 (N_7177,N_6901,N_6998);
or U7178 (N_7178,N_6958,N_6884);
and U7179 (N_7179,N_6834,N_6978);
nand U7180 (N_7180,N_6908,N_6945);
and U7181 (N_7181,N_6872,N_6935);
or U7182 (N_7182,N_6924,N_6829);
or U7183 (N_7183,N_6946,N_6865);
nor U7184 (N_7184,N_6850,N_6842);
or U7185 (N_7185,N_6828,N_6947);
nand U7186 (N_7186,N_6835,N_6991);
or U7187 (N_7187,N_6881,N_6936);
xnor U7188 (N_7188,N_6943,N_6813);
nor U7189 (N_7189,N_6978,N_6854);
or U7190 (N_7190,N_6947,N_6853);
nor U7191 (N_7191,N_6811,N_6917);
nand U7192 (N_7192,N_6882,N_6875);
or U7193 (N_7193,N_6897,N_6849);
or U7194 (N_7194,N_6954,N_6920);
nor U7195 (N_7195,N_6910,N_6984);
nand U7196 (N_7196,N_6896,N_6998);
nor U7197 (N_7197,N_6969,N_6883);
and U7198 (N_7198,N_6946,N_6818);
nand U7199 (N_7199,N_6940,N_6835);
or U7200 (N_7200,N_7109,N_7012);
or U7201 (N_7201,N_7192,N_7016);
nand U7202 (N_7202,N_7163,N_7176);
xor U7203 (N_7203,N_7039,N_7058);
and U7204 (N_7204,N_7088,N_7190);
and U7205 (N_7205,N_7044,N_7020);
or U7206 (N_7206,N_7177,N_7098);
nor U7207 (N_7207,N_7173,N_7031);
or U7208 (N_7208,N_7168,N_7172);
xnor U7209 (N_7209,N_7010,N_7018);
nand U7210 (N_7210,N_7095,N_7151);
nand U7211 (N_7211,N_7140,N_7147);
and U7212 (N_7212,N_7128,N_7053);
xnor U7213 (N_7213,N_7101,N_7111);
nor U7214 (N_7214,N_7171,N_7055);
nor U7215 (N_7215,N_7149,N_7071);
and U7216 (N_7216,N_7129,N_7067);
xnor U7217 (N_7217,N_7092,N_7105);
xnor U7218 (N_7218,N_7054,N_7123);
xnor U7219 (N_7219,N_7076,N_7042);
nor U7220 (N_7220,N_7119,N_7138);
nor U7221 (N_7221,N_7185,N_7112);
and U7222 (N_7222,N_7007,N_7051);
nand U7223 (N_7223,N_7083,N_7079);
and U7224 (N_7224,N_7043,N_7136);
nor U7225 (N_7225,N_7137,N_7028);
nand U7226 (N_7226,N_7046,N_7080);
and U7227 (N_7227,N_7118,N_7022);
or U7228 (N_7228,N_7181,N_7199);
nand U7229 (N_7229,N_7059,N_7170);
and U7230 (N_7230,N_7158,N_7090);
nand U7231 (N_7231,N_7167,N_7062);
nor U7232 (N_7232,N_7078,N_7099);
and U7233 (N_7233,N_7032,N_7120);
xnor U7234 (N_7234,N_7180,N_7125);
and U7235 (N_7235,N_7139,N_7134);
and U7236 (N_7236,N_7144,N_7075);
nand U7237 (N_7237,N_7003,N_7040);
nor U7238 (N_7238,N_7159,N_7184);
nand U7239 (N_7239,N_7198,N_7157);
nand U7240 (N_7240,N_7094,N_7091);
or U7241 (N_7241,N_7093,N_7056);
nand U7242 (N_7242,N_7041,N_7023);
nand U7243 (N_7243,N_7131,N_7179);
nor U7244 (N_7244,N_7126,N_7084);
nor U7245 (N_7245,N_7014,N_7145);
nand U7246 (N_7246,N_7183,N_7188);
nor U7247 (N_7247,N_7006,N_7162);
nand U7248 (N_7248,N_7160,N_7086);
nor U7249 (N_7249,N_7096,N_7100);
and U7250 (N_7250,N_7002,N_7130);
xnor U7251 (N_7251,N_7037,N_7015);
or U7252 (N_7252,N_7035,N_7005);
nand U7253 (N_7253,N_7061,N_7045);
or U7254 (N_7254,N_7009,N_7174);
xor U7255 (N_7255,N_7156,N_7107);
and U7256 (N_7256,N_7036,N_7143);
xnor U7257 (N_7257,N_7030,N_7122);
nor U7258 (N_7258,N_7153,N_7193);
or U7259 (N_7259,N_7034,N_7073);
and U7260 (N_7260,N_7194,N_7197);
nor U7261 (N_7261,N_7102,N_7057);
and U7262 (N_7262,N_7008,N_7148);
nand U7263 (N_7263,N_7178,N_7103);
nand U7264 (N_7264,N_7166,N_7142);
or U7265 (N_7265,N_7038,N_7161);
and U7266 (N_7266,N_7124,N_7026);
nand U7267 (N_7267,N_7050,N_7068);
nor U7268 (N_7268,N_7189,N_7108);
or U7269 (N_7269,N_7047,N_7087);
and U7270 (N_7270,N_7133,N_7175);
or U7271 (N_7271,N_7063,N_7154);
or U7272 (N_7272,N_7074,N_7165);
or U7273 (N_7273,N_7070,N_7127);
xnor U7274 (N_7274,N_7182,N_7132);
and U7275 (N_7275,N_7150,N_7024);
and U7276 (N_7276,N_7013,N_7116);
and U7277 (N_7277,N_7021,N_7017);
and U7278 (N_7278,N_7052,N_7025);
or U7279 (N_7279,N_7164,N_7117);
xnor U7280 (N_7280,N_7104,N_7110);
nor U7281 (N_7281,N_7155,N_7004);
and U7282 (N_7282,N_7066,N_7089);
xor U7283 (N_7283,N_7048,N_7113);
nand U7284 (N_7284,N_7029,N_7064);
or U7285 (N_7285,N_7146,N_7106);
nand U7286 (N_7286,N_7115,N_7019);
nor U7287 (N_7287,N_7114,N_7049);
or U7288 (N_7288,N_7082,N_7033);
and U7289 (N_7289,N_7135,N_7065);
nand U7290 (N_7290,N_7191,N_7081);
or U7291 (N_7291,N_7085,N_7169);
xnor U7292 (N_7292,N_7011,N_7195);
and U7293 (N_7293,N_7000,N_7060);
or U7294 (N_7294,N_7077,N_7097);
nor U7295 (N_7295,N_7186,N_7069);
and U7296 (N_7296,N_7121,N_7072);
nor U7297 (N_7297,N_7001,N_7152);
xor U7298 (N_7298,N_7027,N_7141);
nor U7299 (N_7299,N_7196,N_7187);
or U7300 (N_7300,N_7184,N_7102);
or U7301 (N_7301,N_7152,N_7029);
nor U7302 (N_7302,N_7180,N_7111);
nor U7303 (N_7303,N_7100,N_7002);
nor U7304 (N_7304,N_7143,N_7052);
nor U7305 (N_7305,N_7018,N_7040);
nand U7306 (N_7306,N_7166,N_7199);
nor U7307 (N_7307,N_7017,N_7092);
or U7308 (N_7308,N_7122,N_7181);
or U7309 (N_7309,N_7123,N_7043);
and U7310 (N_7310,N_7125,N_7093);
xnor U7311 (N_7311,N_7068,N_7122);
nor U7312 (N_7312,N_7165,N_7083);
and U7313 (N_7313,N_7046,N_7176);
and U7314 (N_7314,N_7015,N_7111);
or U7315 (N_7315,N_7178,N_7064);
nand U7316 (N_7316,N_7160,N_7044);
nand U7317 (N_7317,N_7118,N_7153);
or U7318 (N_7318,N_7051,N_7197);
or U7319 (N_7319,N_7006,N_7050);
nand U7320 (N_7320,N_7065,N_7053);
nand U7321 (N_7321,N_7058,N_7132);
or U7322 (N_7322,N_7167,N_7192);
nor U7323 (N_7323,N_7005,N_7161);
and U7324 (N_7324,N_7132,N_7198);
and U7325 (N_7325,N_7102,N_7093);
and U7326 (N_7326,N_7018,N_7127);
or U7327 (N_7327,N_7098,N_7058);
nand U7328 (N_7328,N_7119,N_7071);
and U7329 (N_7329,N_7113,N_7169);
nor U7330 (N_7330,N_7058,N_7112);
or U7331 (N_7331,N_7024,N_7159);
xor U7332 (N_7332,N_7093,N_7153);
nor U7333 (N_7333,N_7052,N_7163);
or U7334 (N_7334,N_7095,N_7105);
or U7335 (N_7335,N_7063,N_7103);
nor U7336 (N_7336,N_7137,N_7101);
and U7337 (N_7337,N_7198,N_7094);
and U7338 (N_7338,N_7003,N_7169);
or U7339 (N_7339,N_7079,N_7136);
and U7340 (N_7340,N_7150,N_7029);
nand U7341 (N_7341,N_7078,N_7189);
and U7342 (N_7342,N_7059,N_7197);
xor U7343 (N_7343,N_7189,N_7021);
xnor U7344 (N_7344,N_7174,N_7134);
or U7345 (N_7345,N_7152,N_7042);
nand U7346 (N_7346,N_7141,N_7194);
and U7347 (N_7347,N_7074,N_7142);
or U7348 (N_7348,N_7014,N_7006);
nand U7349 (N_7349,N_7048,N_7107);
nor U7350 (N_7350,N_7103,N_7165);
or U7351 (N_7351,N_7126,N_7115);
and U7352 (N_7352,N_7021,N_7029);
and U7353 (N_7353,N_7181,N_7139);
nand U7354 (N_7354,N_7164,N_7193);
nor U7355 (N_7355,N_7168,N_7022);
xnor U7356 (N_7356,N_7075,N_7159);
or U7357 (N_7357,N_7025,N_7081);
nor U7358 (N_7358,N_7000,N_7126);
or U7359 (N_7359,N_7192,N_7082);
xor U7360 (N_7360,N_7114,N_7154);
xor U7361 (N_7361,N_7175,N_7118);
nand U7362 (N_7362,N_7001,N_7194);
xnor U7363 (N_7363,N_7001,N_7089);
or U7364 (N_7364,N_7162,N_7023);
or U7365 (N_7365,N_7001,N_7018);
nand U7366 (N_7366,N_7182,N_7092);
nand U7367 (N_7367,N_7181,N_7063);
and U7368 (N_7368,N_7064,N_7199);
and U7369 (N_7369,N_7196,N_7147);
nand U7370 (N_7370,N_7120,N_7135);
nand U7371 (N_7371,N_7068,N_7105);
or U7372 (N_7372,N_7038,N_7198);
or U7373 (N_7373,N_7099,N_7164);
xor U7374 (N_7374,N_7034,N_7124);
xor U7375 (N_7375,N_7030,N_7090);
or U7376 (N_7376,N_7032,N_7125);
nor U7377 (N_7377,N_7109,N_7119);
xnor U7378 (N_7378,N_7149,N_7125);
and U7379 (N_7379,N_7096,N_7188);
or U7380 (N_7380,N_7109,N_7168);
or U7381 (N_7381,N_7181,N_7081);
nand U7382 (N_7382,N_7168,N_7151);
and U7383 (N_7383,N_7081,N_7094);
nand U7384 (N_7384,N_7023,N_7051);
nor U7385 (N_7385,N_7136,N_7104);
nor U7386 (N_7386,N_7095,N_7096);
nand U7387 (N_7387,N_7185,N_7158);
or U7388 (N_7388,N_7084,N_7193);
nand U7389 (N_7389,N_7026,N_7164);
xnor U7390 (N_7390,N_7007,N_7008);
and U7391 (N_7391,N_7112,N_7141);
nand U7392 (N_7392,N_7198,N_7099);
xor U7393 (N_7393,N_7002,N_7125);
and U7394 (N_7394,N_7144,N_7038);
or U7395 (N_7395,N_7083,N_7016);
or U7396 (N_7396,N_7138,N_7114);
xor U7397 (N_7397,N_7130,N_7040);
xor U7398 (N_7398,N_7023,N_7187);
nor U7399 (N_7399,N_7181,N_7030);
nand U7400 (N_7400,N_7315,N_7334);
and U7401 (N_7401,N_7336,N_7241);
and U7402 (N_7402,N_7330,N_7240);
xnor U7403 (N_7403,N_7214,N_7351);
nand U7404 (N_7404,N_7231,N_7338);
xor U7405 (N_7405,N_7313,N_7299);
or U7406 (N_7406,N_7305,N_7350);
or U7407 (N_7407,N_7257,N_7337);
nand U7408 (N_7408,N_7347,N_7216);
xnor U7409 (N_7409,N_7385,N_7389);
or U7410 (N_7410,N_7242,N_7223);
xnor U7411 (N_7411,N_7228,N_7275);
xor U7412 (N_7412,N_7369,N_7247);
or U7413 (N_7413,N_7218,N_7279);
xor U7414 (N_7414,N_7249,N_7398);
nor U7415 (N_7415,N_7304,N_7285);
xor U7416 (N_7416,N_7333,N_7264);
or U7417 (N_7417,N_7308,N_7248);
nor U7418 (N_7418,N_7276,N_7206);
nand U7419 (N_7419,N_7290,N_7212);
and U7420 (N_7420,N_7237,N_7387);
xor U7421 (N_7421,N_7380,N_7376);
nand U7422 (N_7422,N_7345,N_7293);
and U7423 (N_7423,N_7256,N_7339);
xor U7424 (N_7424,N_7277,N_7319);
nand U7425 (N_7425,N_7374,N_7349);
nor U7426 (N_7426,N_7233,N_7243);
and U7427 (N_7427,N_7346,N_7245);
xor U7428 (N_7428,N_7384,N_7343);
xnor U7429 (N_7429,N_7399,N_7244);
and U7430 (N_7430,N_7298,N_7282);
nor U7431 (N_7431,N_7395,N_7229);
nand U7432 (N_7432,N_7379,N_7254);
nand U7433 (N_7433,N_7375,N_7225);
and U7434 (N_7434,N_7263,N_7397);
nand U7435 (N_7435,N_7364,N_7221);
and U7436 (N_7436,N_7255,N_7393);
nand U7437 (N_7437,N_7360,N_7222);
and U7438 (N_7438,N_7204,N_7386);
and U7439 (N_7439,N_7213,N_7318);
or U7440 (N_7440,N_7232,N_7252);
nor U7441 (N_7441,N_7265,N_7361);
and U7442 (N_7442,N_7294,N_7238);
xor U7443 (N_7443,N_7224,N_7219);
or U7444 (N_7444,N_7323,N_7365);
nor U7445 (N_7445,N_7239,N_7355);
nand U7446 (N_7446,N_7287,N_7328);
xnor U7447 (N_7447,N_7253,N_7327);
nor U7448 (N_7448,N_7234,N_7390);
and U7449 (N_7449,N_7292,N_7230);
xor U7450 (N_7450,N_7382,N_7217);
nand U7451 (N_7451,N_7363,N_7329);
xor U7452 (N_7452,N_7394,N_7322);
nand U7453 (N_7453,N_7201,N_7280);
and U7454 (N_7454,N_7286,N_7383);
nand U7455 (N_7455,N_7266,N_7296);
xor U7456 (N_7456,N_7340,N_7274);
nor U7457 (N_7457,N_7302,N_7205);
xnor U7458 (N_7458,N_7326,N_7357);
nand U7459 (N_7459,N_7320,N_7200);
xnor U7460 (N_7460,N_7273,N_7203);
nor U7461 (N_7461,N_7353,N_7301);
nor U7462 (N_7462,N_7392,N_7354);
nor U7463 (N_7463,N_7366,N_7291);
and U7464 (N_7464,N_7226,N_7344);
or U7465 (N_7465,N_7295,N_7270);
or U7466 (N_7466,N_7335,N_7283);
nand U7467 (N_7467,N_7310,N_7358);
xnor U7468 (N_7468,N_7381,N_7331);
xor U7469 (N_7469,N_7215,N_7235);
nand U7470 (N_7470,N_7208,N_7314);
and U7471 (N_7471,N_7321,N_7348);
nand U7472 (N_7472,N_7250,N_7260);
nor U7473 (N_7473,N_7377,N_7289);
nand U7474 (N_7474,N_7267,N_7251);
xnor U7475 (N_7475,N_7368,N_7278);
nor U7476 (N_7476,N_7262,N_7281);
or U7477 (N_7477,N_7342,N_7259);
nor U7478 (N_7478,N_7271,N_7268);
xnor U7479 (N_7479,N_7261,N_7325);
and U7480 (N_7480,N_7372,N_7352);
nand U7481 (N_7481,N_7300,N_7202);
xor U7482 (N_7482,N_7311,N_7388);
and U7483 (N_7483,N_7370,N_7258);
nand U7484 (N_7484,N_7316,N_7309);
and U7485 (N_7485,N_7341,N_7312);
xnor U7486 (N_7486,N_7220,N_7378);
or U7487 (N_7487,N_7207,N_7209);
nor U7488 (N_7488,N_7236,N_7324);
nor U7489 (N_7489,N_7246,N_7269);
nor U7490 (N_7490,N_7396,N_7297);
or U7491 (N_7491,N_7272,N_7359);
nand U7492 (N_7492,N_7356,N_7391);
nor U7493 (N_7493,N_7362,N_7210);
nor U7494 (N_7494,N_7284,N_7332);
or U7495 (N_7495,N_7288,N_7306);
nand U7496 (N_7496,N_7211,N_7371);
or U7497 (N_7497,N_7373,N_7367);
nand U7498 (N_7498,N_7303,N_7307);
xor U7499 (N_7499,N_7317,N_7227);
xnor U7500 (N_7500,N_7330,N_7363);
and U7501 (N_7501,N_7245,N_7344);
nand U7502 (N_7502,N_7202,N_7345);
or U7503 (N_7503,N_7319,N_7219);
nand U7504 (N_7504,N_7252,N_7261);
nand U7505 (N_7505,N_7206,N_7330);
or U7506 (N_7506,N_7261,N_7312);
nand U7507 (N_7507,N_7307,N_7222);
or U7508 (N_7508,N_7258,N_7340);
or U7509 (N_7509,N_7277,N_7387);
or U7510 (N_7510,N_7211,N_7385);
xor U7511 (N_7511,N_7290,N_7328);
nor U7512 (N_7512,N_7276,N_7248);
and U7513 (N_7513,N_7396,N_7223);
or U7514 (N_7514,N_7382,N_7313);
nor U7515 (N_7515,N_7236,N_7384);
and U7516 (N_7516,N_7318,N_7355);
or U7517 (N_7517,N_7241,N_7329);
or U7518 (N_7518,N_7398,N_7278);
xnor U7519 (N_7519,N_7234,N_7370);
and U7520 (N_7520,N_7286,N_7377);
xnor U7521 (N_7521,N_7330,N_7304);
or U7522 (N_7522,N_7391,N_7360);
or U7523 (N_7523,N_7232,N_7381);
xnor U7524 (N_7524,N_7366,N_7305);
and U7525 (N_7525,N_7219,N_7240);
and U7526 (N_7526,N_7282,N_7334);
nand U7527 (N_7527,N_7384,N_7217);
nor U7528 (N_7528,N_7322,N_7244);
nor U7529 (N_7529,N_7286,N_7358);
nor U7530 (N_7530,N_7329,N_7246);
and U7531 (N_7531,N_7222,N_7362);
and U7532 (N_7532,N_7391,N_7252);
nand U7533 (N_7533,N_7234,N_7218);
nand U7534 (N_7534,N_7293,N_7371);
nor U7535 (N_7535,N_7380,N_7240);
or U7536 (N_7536,N_7298,N_7250);
nor U7537 (N_7537,N_7266,N_7366);
or U7538 (N_7538,N_7343,N_7233);
or U7539 (N_7539,N_7241,N_7202);
or U7540 (N_7540,N_7270,N_7371);
nor U7541 (N_7541,N_7308,N_7384);
and U7542 (N_7542,N_7219,N_7381);
xor U7543 (N_7543,N_7354,N_7253);
and U7544 (N_7544,N_7340,N_7326);
nor U7545 (N_7545,N_7299,N_7329);
nor U7546 (N_7546,N_7209,N_7336);
and U7547 (N_7547,N_7397,N_7354);
xnor U7548 (N_7548,N_7215,N_7213);
or U7549 (N_7549,N_7347,N_7370);
and U7550 (N_7550,N_7349,N_7288);
nor U7551 (N_7551,N_7362,N_7388);
xor U7552 (N_7552,N_7236,N_7211);
xor U7553 (N_7553,N_7342,N_7275);
nor U7554 (N_7554,N_7339,N_7299);
nor U7555 (N_7555,N_7322,N_7365);
and U7556 (N_7556,N_7361,N_7269);
or U7557 (N_7557,N_7301,N_7246);
nand U7558 (N_7558,N_7287,N_7225);
nand U7559 (N_7559,N_7253,N_7319);
and U7560 (N_7560,N_7354,N_7366);
or U7561 (N_7561,N_7257,N_7382);
and U7562 (N_7562,N_7390,N_7325);
nand U7563 (N_7563,N_7313,N_7239);
xnor U7564 (N_7564,N_7384,N_7213);
nor U7565 (N_7565,N_7250,N_7264);
nand U7566 (N_7566,N_7390,N_7206);
nor U7567 (N_7567,N_7225,N_7285);
nand U7568 (N_7568,N_7388,N_7300);
xor U7569 (N_7569,N_7312,N_7338);
nand U7570 (N_7570,N_7229,N_7223);
and U7571 (N_7571,N_7215,N_7322);
xor U7572 (N_7572,N_7255,N_7296);
or U7573 (N_7573,N_7348,N_7207);
xnor U7574 (N_7574,N_7334,N_7381);
nand U7575 (N_7575,N_7201,N_7373);
nand U7576 (N_7576,N_7389,N_7325);
nand U7577 (N_7577,N_7344,N_7299);
and U7578 (N_7578,N_7323,N_7223);
nand U7579 (N_7579,N_7348,N_7373);
or U7580 (N_7580,N_7228,N_7345);
or U7581 (N_7581,N_7232,N_7334);
nand U7582 (N_7582,N_7285,N_7231);
and U7583 (N_7583,N_7324,N_7328);
nand U7584 (N_7584,N_7211,N_7283);
nor U7585 (N_7585,N_7370,N_7205);
nand U7586 (N_7586,N_7350,N_7290);
nand U7587 (N_7587,N_7395,N_7209);
nor U7588 (N_7588,N_7264,N_7349);
xnor U7589 (N_7589,N_7218,N_7396);
and U7590 (N_7590,N_7219,N_7252);
xnor U7591 (N_7591,N_7236,N_7313);
nand U7592 (N_7592,N_7255,N_7230);
nand U7593 (N_7593,N_7299,N_7260);
and U7594 (N_7594,N_7214,N_7378);
xor U7595 (N_7595,N_7264,N_7392);
or U7596 (N_7596,N_7215,N_7347);
nor U7597 (N_7597,N_7348,N_7307);
and U7598 (N_7598,N_7209,N_7322);
nor U7599 (N_7599,N_7249,N_7337);
or U7600 (N_7600,N_7497,N_7526);
nor U7601 (N_7601,N_7498,N_7449);
or U7602 (N_7602,N_7403,N_7520);
nor U7603 (N_7603,N_7481,N_7470);
or U7604 (N_7604,N_7523,N_7488);
xor U7605 (N_7605,N_7478,N_7530);
and U7606 (N_7606,N_7451,N_7563);
or U7607 (N_7607,N_7516,N_7476);
nor U7608 (N_7608,N_7493,N_7420);
and U7609 (N_7609,N_7594,N_7400);
and U7610 (N_7610,N_7415,N_7557);
or U7611 (N_7611,N_7538,N_7463);
nand U7612 (N_7612,N_7504,N_7568);
nand U7613 (N_7613,N_7510,N_7503);
and U7614 (N_7614,N_7433,N_7529);
nand U7615 (N_7615,N_7465,N_7517);
and U7616 (N_7616,N_7565,N_7522);
nor U7617 (N_7617,N_7427,N_7455);
xor U7618 (N_7618,N_7561,N_7483);
nand U7619 (N_7619,N_7480,N_7460);
or U7620 (N_7620,N_7490,N_7438);
xor U7621 (N_7621,N_7548,N_7461);
or U7622 (N_7622,N_7458,N_7413);
nand U7623 (N_7623,N_7531,N_7596);
and U7624 (N_7624,N_7507,N_7585);
xnor U7625 (N_7625,N_7426,N_7553);
or U7626 (N_7626,N_7508,N_7443);
or U7627 (N_7627,N_7552,N_7527);
nand U7628 (N_7628,N_7467,N_7515);
and U7629 (N_7629,N_7519,N_7569);
nand U7630 (N_7630,N_7572,N_7502);
nand U7631 (N_7631,N_7524,N_7546);
or U7632 (N_7632,N_7414,N_7444);
or U7633 (N_7633,N_7536,N_7584);
and U7634 (N_7634,N_7555,N_7485);
nand U7635 (N_7635,N_7423,N_7582);
and U7636 (N_7636,N_7533,N_7487);
xor U7637 (N_7637,N_7578,N_7580);
nor U7638 (N_7638,N_7469,N_7535);
or U7639 (N_7639,N_7468,N_7597);
and U7640 (N_7640,N_7409,N_7543);
or U7641 (N_7641,N_7491,N_7588);
nand U7642 (N_7642,N_7590,N_7464);
nand U7643 (N_7643,N_7525,N_7573);
nor U7644 (N_7644,N_7450,N_7473);
and U7645 (N_7645,N_7581,N_7571);
or U7646 (N_7646,N_7437,N_7408);
and U7647 (N_7647,N_7435,N_7432);
nor U7648 (N_7648,N_7541,N_7521);
and U7649 (N_7649,N_7591,N_7430);
or U7650 (N_7650,N_7532,N_7537);
xor U7651 (N_7651,N_7466,N_7417);
or U7652 (N_7652,N_7462,N_7482);
or U7653 (N_7653,N_7442,N_7405);
and U7654 (N_7654,N_7471,N_7562);
nand U7655 (N_7655,N_7445,N_7499);
xor U7656 (N_7656,N_7598,N_7419);
or U7657 (N_7657,N_7539,N_7412);
xnor U7658 (N_7658,N_7575,N_7500);
and U7659 (N_7659,N_7439,N_7441);
nand U7660 (N_7660,N_7453,N_7474);
nor U7661 (N_7661,N_7440,N_7501);
nor U7662 (N_7662,N_7551,N_7547);
or U7663 (N_7663,N_7570,N_7406);
nand U7664 (N_7664,N_7472,N_7518);
nor U7665 (N_7665,N_7486,N_7583);
or U7666 (N_7666,N_7505,N_7425);
nand U7667 (N_7667,N_7457,N_7506);
xnor U7668 (N_7668,N_7421,N_7574);
xnor U7669 (N_7669,N_7592,N_7556);
xnor U7670 (N_7670,N_7558,N_7560);
and U7671 (N_7671,N_7511,N_7513);
nand U7672 (N_7672,N_7494,N_7401);
xor U7673 (N_7673,N_7411,N_7495);
nand U7674 (N_7674,N_7484,N_7407);
xor U7675 (N_7675,N_7446,N_7554);
and U7676 (N_7676,N_7595,N_7534);
or U7677 (N_7677,N_7428,N_7528);
nor U7678 (N_7678,N_7512,N_7509);
and U7679 (N_7679,N_7418,N_7577);
xnor U7680 (N_7680,N_7586,N_7410);
nand U7681 (N_7681,N_7540,N_7422);
nand U7682 (N_7682,N_7416,N_7542);
nand U7683 (N_7683,N_7434,N_7479);
or U7684 (N_7684,N_7566,N_7459);
nor U7685 (N_7685,N_7545,N_7550);
nor U7686 (N_7686,N_7447,N_7559);
or U7687 (N_7687,N_7456,N_7579);
or U7688 (N_7688,N_7436,N_7452);
and U7689 (N_7689,N_7402,N_7431);
xor U7690 (N_7690,N_7424,N_7544);
nor U7691 (N_7691,N_7549,N_7599);
or U7692 (N_7692,N_7564,N_7567);
nand U7693 (N_7693,N_7429,N_7496);
nor U7694 (N_7694,N_7489,N_7589);
nand U7695 (N_7695,N_7587,N_7475);
nor U7696 (N_7696,N_7404,N_7448);
and U7697 (N_7697,N_7477,N_7593);
nand U7698 (N_7698,N_7576,N_7514);
or U7699 (N_7699,N_7492,N_7454);
nor U7700 (N_7700,N_7452,N_7477);
xnor U7701 (N_7701,N_7550,N_7517);
nand U7702 (N_7702,N_7573,N_7569);
or U7703 (N_7703,N_7492,N_7513);
and U7704 (N_7704,N_7538,N_7510);
xor U7705 (N_7705,N_7595,N_7551);
nor U7706 (N_7706,N_7599,N_7582);
nor U7707 (N_7707,N_7554,N_7418);
nor U7708 (N_7708,N_7435,N_7415);
and U7709 (N_7709,N_7438,N_7410);
or U7710 (N_7710,N_7582,N_7536);
xor U7711 (N_7711,N_7583,N_7506);
and U7712 (N_7712,N_7581,N_7464);
nand U7713 (N_7713,N_7588,N_7435);
and U7714 (N_7714,N_7498,N_7522);
or U7715 (N_7715,N_7492,N_7549);
nand U7716 (N_7716,N_7531,N_7544);
or U7717 (N_7717,N_7400,N_7447);
or U7718 (N_7718,N_7483,N_7431);
nor U7719 (N_7719,N_7591,N_7417);
and U7720 (N_7720,N_7465,N_7490);
and U7721 (N_7721,N_7538,N_7419);
and U7722 (N_7722,N_7572,N_7556);
or U7723 (N_7723,N_7501,N_7536);
nor U7724 (N_7724,N_7558,N_7457);
xor U7725 (N_7725,N_7422,N_7418);
nand U7726 (N_7726,N_7400,N_7561);
nor U7727 (N_7727,N_7482,N_7555);
nand U7728 (N_7728,N_7561,N_7447);
nor U7729 (N_7729,N_7542,N_7564);
xnor U7730 (N_7730,N_7400,N_7511);
nand U7731 (N_7731,N_7438,N_7504);
nand U7732 (N_7732,N_7454,N_7585);
xnor U7733 (N_7733,N_7451,N_7467);
nor U7734 (N_7734,N_7407,N_7412);
and U7735 (N_7735,N_7421,N_7478);
or U7736 (N_7736,N_7435,N_7409);
xnor U7737 (N_7737,N_7569,N_7454);
nor U7738 (N_7738,N_7407,N_7405);
nand U7739 (N_7739,N_7466,N_7519);
and U7740 (N_7740,N_7492,N_7421);
and U7741 (N_7741,N_7468,N_7449);
and U7742 (N_7742,N_7472,N_7449);
nand U7743 (N_7743,N_7580,N_7522);
or U7744 (N_7744,N_7598,N_7406);
or U7745 (N_7745,N_7498,N_7588);
nand U7746 (N_7746,N_7497,N_7489);
and U7747 (N_7747,N_7435,N_7552);
nor U7748 (N_7748,N_7485,N_7453);
or U7749 (N_7749,N_7535,N_7413);
and U7750 (N_7750,N_7449,N_7421);
and U7751 (N_7751,N_7454,N_7546);
and U7752 (N_7752,N_7566,N_7584);
nor U7753 (N_7753,N_7549,N_7580);
and U7754 (N_7754,N_7405,N_7417);
nor U7755 (N_7755,N_7560,N_7592);
nand U7756 (N_7756,N_7422,N_7472);
nand U7757 (N_7757,N_7591,N_7552);
or U7758 (N_7758,N_7478,N_7532);
or U7759 (N_7759,N_7502,N_7447);
and U7760 (N_7760,N_7562,N_7459);
and U7761 (N_7761,N_7464,N_7421);
and U7762 (N_7762,N_7569,N_7451);
xor U7763 (N_7763,N_7442,N_7527);
or U7764 (N_7764,N_7449,N_7429);
nand U7765 (N_7765,N_7419,N_7408);
nand U7766 (N_7766,N_7573,N_7475);
nor U7767 (N_7767,N_7498,N_7513);
and U7768 (N_7768,N_7455,N_7570);
xor U7769 (N_7769,N_7457,N_7512);
xnor U7770 (N_7770,N_7458,N_7438);
nor U7771 (N_7771,N_7479,N_7519);
or U7772 (N_7772,N_7419,N_7521);
xnor U7773 (N_7773,N_7501,N_7441);
xor U7774 (N_7774,N_7448,N_7465);
nand U7775 (N_7775,N_7554,N_7532);
nand U7776 (N_7776,N_7595,N_7430);
and U7777 (N_7777,N_7459,N_7534);
nor U7778 (N_7778,N_7409,N_7461);
and U7779 (N_7779,N_7475,N_7485);
and U7780 (N_7780,N_7416,N_7551);
nor U7781 (N_7781,N_7428,N_7540);
nand U7782 (N_7782,N_7428,N_7406);
or U7783 (N_7783,N_7507,N_7570);
nand U7784 (N_7784,N_7455,N_7554);
or U7785 (N_7785,N_7518,N_7532);
or U7786 (N_7786,N_7410,N_7418);
nor U7787 (N_7787,N_7558,N_7417);
xnor U7788 (N_7788,N_7594,N_7517);
or U7789 (N_7789,N_7541,N_7510);
nor U7790 (N_7790,N_7487,N_7544);
or U7791 (N_7791,N_7571,N_7481);
nand U7792 (N_7792,N_7401,N_7488);
and U7793 (N_7793,N_7505,N_7431);
xor U7794 (N_7794,N_7456,N_7474);
and U7795 (N_7795,N_7560,N_7543);
and U7796 (N_7796,N_7560,N_7581);
and U7797 (N_7797,N_7440,N_7492);
xor U7798 (N_7798,N_7474,N_7410);
nor U7799 (N_7799,N_7530,N_7507);
nand U7800 (N_7800,N_7770,N_7712);
nor U7801 (N_7801,N_7714,N_7644);
or U7802 (N_7802,N_7761,N_7764);
nand U7803 (N_7803,N_7702,N_7600);
or U7804 (N_7804,N_7662,N_7669);
nand U7805 (N_7805,N_7636,N_7690);
xnor U7806 (N_7806,N_7745,N_7647);
xnor U7807 (N_7807,N_7792,N_7732);
nor U7808 (N_7808,N_7666,N_7789);
or U7809 (N_7809,N_7736,N_7629);
or U7810 (N_7810,N_7760,N_7723);
nand U7811 (N_7811,N_7618,N_7727);
nand U7812 (N_7812,N_7799,N_7706);
nor U7813 (N_7813,N_7741,N_7643);
xnor U7814 (N_7814,N_7729,N_7758);
nor U7815 (N_7815,N_7720,N_7677);
or U7816 (N_7816,N_7766,N_7796);
nor U7817 (N_7817,N_7776,N_7674);
or U7818 (N_7818,N_7721,N_7641);
nor U7819 (N_7819,N_7785,N_7635);
nand U7820 (N_7820,N_7704,N_7794);
nand U7821 (N_7821,N_7718,N_7670);
and U7822 (N_7822,N_7694,N_7784);
nand U7823 (N_7823,N_7683,N_7687);
xnor U7824 (N_7824,N_7747,N_7612);
and U7825 (N_7825,N_7697,N_7752);
nand U7826 (N_7826,N_7744,N_7765);
nand U7827 (N_7827,N_7616,N_7627);
xor U7828 (N_7828,N_7679,N_7711);
or U7829 (N_7829,N_7757,N_7624);
and U7830 (N_7830,N_7671,N_7716);
or U7831 (N_7831,N_7699,N_7790);
xnor U7832 (N_7832,N_7680,N_7622);
and U7833 (N_7833,N_7733,N_7604);
nand U7834 (N_7834,N_7628,N_7780);
nand U7835 (N_7835,N_7638,N_7715);
nor U7836 (N_7836,N_7639,N_7742);
nand U7837 (N_7837,N_7781,N_7611);
nor U7838 (N_7838,N_7713,N_7798);
nor U7839 (N_7839,N_7743,N_7775);
and U7840 (N_7840,N_7667,N_7610);
xor U7841 (N_7841,N_7746,N_7659);
or U7842 (N_7842,N_7652,N_7660);
and U7843 (N_7843,N_7717,N_7709);
xnor U7844 (N_7844,N_7782,N_7707);
and U7845 (N_7845,N_7632,N_7657);
nand U7846 (N_7846,N_7797,N_7726);
xnor U7847 (N_7847,N_7701,N_7719);
and U7848 (N_7848,N_7607,N_7609);
nand U7849 (N_7849,N_7658,N_7602);
xnor U7850 (N_7850,N_7678,N_7751);
nor U7851 (N_7851,N_7735,N_7774);
and U7852 (N_7852,N_7642,N_7793);
nand U7853 (N_7853,N_7705,N_7654);
nand U7854 (N_7854,N_7703,N_7625);
and U7855 (N_7855,N_7739,N_7656);
nor U7856 (N_7856,N_7606,N_7695);
nor U7857 (N_7857,N_7651,N_7672);
and U7858 (N_7858,N_7661,N_7686);
nand U7859 (N_7859,N_7637,N_7768);
and U7860 (N_7860,N_7763,N_7665);
xnor U7861 (N_7861,N_7696,N_7738);
xnor U7862 (N_7862,N_7681,N_7779);
xnor U7863 (N_7863,N_7725,N_7731);
and U7864 (N_7864,N_7689,N_7615);
nand U7865 (N_7865,N_7626,N_7722);
nand U7866 (N_7866,N_7648,N_7688);
nand U7867 (N_7867,N_7676,N_7645);
nor U7868 (N_7868,N_7630,N_7664);
xnor U7869 (N_7869,N_7700,N_7791);
xor U7870 (N_7870,N_7795,N_7750);
and U7871 (N_7871,N_7685,N_7653);
nor U7872 (N_7872,N_7767,N_7693);
xor U7873 (N_7873,N_7777,N_7675);
nor U7874 (N_7874,N_7749,N_7621);
and U7875 (N_7875,N_7769,N_7619);
and U7876 (N_7876,N_7788,N_7754);
nand U7877 (N_7877,N_7620,N_7710);
xor U7878 (N_7878,N_7783,N_7614);
xor U7879 (N_7879,N_7734,N_7663);
nand U7880 (N_7880,N_7759,N_7698);
nand U7881 (N_7881,N_7640,N_7692);
or U7882 (N_7882,N_7755,N_7756);
and U7883 (N_7883,N_7762,N_7601);
nand U7884 (N_7884,N_7608,N_7748);
nor U7885 (N_7885,N_7634,N_7655);
or U7886 (N_7886,N_7649,N_7730);
nand U7887 (N_7887,N_7772,N_7684);
or U7888 (N_7888,N_7682,N_7603);
or U7889 (N_7889,N_7778,N_7650);
xor U7890 (N_7890,N_7605,N_7708);
and U7891 (N_7891,N_7646,N_7668);
nor U7892 (N_7892,N_7737,N_7787);
nor U7893 (N_7893,N_7773,N_7617);
xor U7894 (N_7894,N_7724,N_7771);
or U7895 (N_7895,N_7623,N_7673);
and U7896 (N_7896,N_7613,N_7631);
xor U7897 (N_7897,N_7740,N_7728);
or U7898 (N_7898,N_7691,N_7633);
xnor U7899 (N_7899,N_7753,N_7786);
and U7900 (N_7900,N_7773,N_7714);
xor U7901 (N_7901,N_7618,N_7776);
nand U7902 (N_7902,N_7767,N_7734);
nor U7903 (N_7903,N_7705,N_7667);
and U7904 (N_7904,N_7717,N_7757);
or U7905 (N_7905,N_7707,N_7792);
nand U7906 (N_7906,N_7744,N_7664);
and U7907 (N_7907,N_7775,N_7785);
nor U7908 (N_7908,N_7780,N_7670);
or U7909 (N_7909,N_7668,N_7718);
or U7910 (N_7910,N_7728,N_7664);
xor U7911 (N_7911,N_7681,N_7686);
nor U7912 (N_7912,N_7740,N_7653);
or U7913 (N_7913,N_7662,N_7695);
or U7914 (N_7914,N_7798,N_7785);
or U7915 (N_7915,N_7791,N_7653);
xnor U7916 (N_7916,N_7670,N_7676);
nand U7917 (N_7917,N_7672,N_7711);
and U7918 (N_7918,N_7651,N_7758);
nand U7919 (N_7919,N_7717,N_7652);
nor U7920 (N_7920,N_7733,N_7692);
or U7921 (N_7921,N_7666,N_7765);
or U7922 (N_7922,N_7690,N_7720);
nand U7923 (N_7923,N_7768,N_7767);
and U7924 (N_7924,N_7791,N_7763);
nand U7925 (N_7925,N_7743,N_7741);
xnor U7926 (N_7926,N_7647,N_7703);
nand U7927 (N_7927,N_7731,N_7748);
nand U7928 (N_7928,N_7773,N_7724);
xor U7929 (N_7929,N_7750,N_7619);
or U7930 (N_7930,N_7740,N_7654);
xnor U7931 (N_7931,N_7679,N_7629);
nand U7932 (N_7932,N_7607,N_7781);
nor U7933 (N_7933,N_7629,N_7700);
nor U7934 (N_7934,N_7700,N_7753);
and U7935 (N_7935,N_7785,N_7741);
nand U7936 (N_7936,N_7702,N_7655);
or U7937 (N_7937,N_7628,N_7793);
nand U7938 (N_7938,N_7640,N_7758);
or U7939 (N_7939,N_7732,N_7708);
xnor U7940 (N_7940,N_7689,N_7671);
xnor U7941 (N_7941,N_7651,N_7784);
and U7942 (N_7942,N_7606,N_7749);
xor U7943 (N_7943,N_7648,N_7631);
or U7944 (N_7944,N_7695,N_7736);
nand U7945 (N_7945,N_7749,N_7797);
or U7946 (N_7946,N_7613,N_7642);
and U7947 (N_7947,N_7722,N_7649);
nand U7948 (N_7948,N_7636,N_7716);
and U7949 (N_7949,N_7742,N_7647);
nand U7950 (N_7950,N_7623,N_7795);
and U7951 (N_7951,N_7733,N_7612);
nand U7952 (N_7952,N_7644,N_7660);
nor U7953 (N_7953,N_7604,N_7707);
nor U7954 (N_7954,N_7712,N_7636);
or U7955 (N_7955,N_7640,N_7730);
and U7956 (N_7956,N_7792,N_7720);
nor U7957 (N_7957,N_7793,N_7668);
and U7958 (N_7958,N_7639,N_7752);
and U7959 (N_7959,N_7651,N_7731);
nand U7960 (N_7960,N_7736,N_7763);
nand U7961 (N_7961,N_7792,N_7622);
nor U7962 (N_7962,N_7774,N_7602);
xor U7963 (N_7963,N_7797,N_7663);
and U7964 (N_7964,N_7632,N_7715);
nand U7965 (N_7965,N_7645,N_7644);
or U7966 (N_7966,N_7637,N_7690);
xnor U7967 (N_7967,N_7622,N_7780);
nand U7968 (N_7968,N_7622,N_7608);
nor U7969 (N_7969,N_7773,N_7621);
nand U7970 (N_7970,N_7696,N_7611);
and U7971 (N_7971,N_7699,N_7640);
xor U7972 (N_7972,N_7658,N_7754);
or U7973 (N_7973,N_7613,N_7768);
xor U7974 (N_7974,N_7673,N_7782);
nand U7975 (N_7975,N_7784,N_7791);
nand U7976 (N_7976,N_7750,N_7603);
or U7977 (N_7977,N_7709,N_7705);
nand U7978 (N_7978,N_7631,N_7654);
or U7979 (N_7979,N_7763,N_7742);
xor U7980 (N_7980,N_7762,N_7694);
xnor U7981 (N_7981,N_7736,N_7799);
and U7982 (N_7982,N_7745,N_7799);
xnor U7983 (N_7983,N_7710,N_7674);
and U7984 (N_7984,N_7695,N_7746);
nor U7985 (N_7985,N_7745,N_7785);
nor U7986 (N_7986,N_7724,N_7620);
nor U7987 (N_7987,N_7724,N_7763);
or U7988 (N_7988,N_7734,N_7783);
or U7989 (N_7989,N_7786,N_7705);
nand U7990 (N_7990,N_7749,N_7671);
nand U7991 (N_7991,N_7657,N_7748);
nand U7992 (N_7992,N_7605,N_7759);
nor U7993 (N_7993,N_7712,N_7780);
nand U7994 (N_7994,N_7761,N_7791);
nor U7995 (N_7995,N_7770,N_7634);
xor U7996 (N_7996,N_7749,N_7654);
xnor U7997 (N_7997,N_7741,N_7664);
nand U7998 (N_7998,N_7693,N_7716);
nand U7999 (N_7999,N_7759,N_7613);
nor U8000 (N_8000,N_7867,N_7974);
xor U8001 (N_8001,N_7982,N_7804);
nand U8002 (N_8002,N_7920,N_7874);
xnor U8003 (N_8003,N_7992,N_7859);
nor U8004 (N_8004,N_7943,N_7860);
nand U8005 (N_8005,N_7810,N_7801);
and U8006 (N_8006,N_7897,N_7809);
and U8007 (N_8007,N_7829,N_7939);
or U8008 (N_8008,N_7877,N_7889);
and U8009 (N_8009,N_7987,N_7854);
xor U8010 (N_8010,N_7833,N_7946);
and U8011 (N_8011,N_7928,N_7844);
xnor U8012 (N_8012,N_7983,N_7990);
or U8013 (N_8013,N_7948,N_7848);
nand U8014 (N_8014,N_7816,N_7823);
nand U8015 (N_8015,N_7862,N_7818);
nor U8016 (N_8016,N_7879,N_7807);
nand U8017 (N_8017,N_7985,N_7839);
xor U8018 (N_8018,N_7940,N_7890);
nor U8019 (N_8019,N_7917,N_7808);
and U8020 (N_8020,N_7975,N_7893);
nor U8021 (N_8021,N_7942,N_7956);
nor U8022 (N_8022,N_7955,N_7938);
xor U8023 (N_8023,N_7819,N_7958);
or U8024 (N_8024,N_7842,N_7966);
nand U8025 (N_8025,N_7962,N_7967);
or U8026 (N_8026,N_7909,N_7869);
nor U8027 (N_8027,N_7930,N_7953);
or U8028 (N_8028,N_7872,N_7864);
xnor U8029 (N_8029,N_7994,N_7954);
or U8030 (N_8030,N_7972,N_7927);
and U8031 (N_8031,N_7876,N_7881);
or U8032 (N_8032,N_7904,N_7853);
nand U8033 (N_8033,N_7825,N_7901);
xnor U8034 (N_8034,N_7944,N_7941);
nand U8035 (N_8035,N_7937,N_7849);
nand U8036 (N_8036,N_7878,N_7899);
xor U8037 (N_8037,N_7999,N_7820);
xnor U8038 (N_8038,N_7911,N_7949);
and U8039 (N_8039,N_7986,N_7870);
and U8040 (N_8040,N_7925,N_7906);
nand U8041 (N_8041,N_7905,N_7989);
or U8042 (N_8042,N_7806,N_7970);
and U8043 (N_8043,N_7984,N_7934);
nand U8044 (N_8044,N_7873,N_7815);
and U8045 (N_8045,N_7817,N_7891);
and U8046 (N_8046,N_7981,N_7931);
nor U8047 (N_8047,N_7910,N_7847);
xnor U8048 (N_8048,N_7871,N_7924);
and U8049 (N_8049,N_7821,N_7866);
nand U8050 (N_8050,N_7882,N_7902);
nor U8051 (N_8051,N_7868,N_7834);
and U8052 (N_8052,N_7892,N_7980);
nand U8053 (N_8053,N_7964,N_7945);
nor U8054 (N_8054,N_7957,N_7886);
or U8055 (N_8055,N_7888,N_7908);
xnor U8056 (N_8056,N_7875,N_7998);
xor U8057 (N_8057,N_7926,N_7963);
xnor U8058 (N_8058,N_7968,N_7855);
and U8059 (N_8059,N_7843,N_7947);
xnor U8060 (N_8060,N_7880,N_7827);
xnor U8061 (N_8061,N_7971,N_7973);
and U8062 (N_8062,N_7978,N_7861);
and U8063 (N_8063,N_7933,N_7812);
or U8064 (N_8064,N_7857,N_7929);
nor U8065 (N_8065,N_7831,N_7979);
or U8066 (N_8066,N_7960,N_7997);
xor U8067 (N_8067,N_7916,N_7951);
xnor U8068 (N_8068,N_7977,N_7993);
or U8069 (N_8069,N_7840,N_7838);
nor U8070 (N_8070,N_7835,N_7845);
or U8071 (N_8071,N_7995,N_7894);
xnor U8072 (N_8072,N_7903,N_7907);
and U8073 (N_8073,N_7822,N_7914);
or U8074 (N_8074,N_7863,N_7921);
or U8075 (N_8075,N_7858,N_7885);
and U8076 (N_8076,N_7895,N_7883);
or U8077 (N_8077,N_7802,N_7900);
nor U8078 (N_8078,N_7851,N_7919);
nor U8079 (N_8079,N_7850,N_7837);
and U8080 (N_8080,N_7988,N_7852);
and U8081 (N_8081,N_7803,N_7936);
nor U8082 (N_8082,N_7898,N_7935);
and U8083 (N_8083,N_7826,N_7950);
or U8084 (N_8084,N_7915,N_7811);
nor U8085 (N_8085,N_7913,N_7836);
nor U8086 (N_8086,N_7923,N_7996);
and U8087 (N_8087,N_7828,N_7959);
or U8088 (N_8088,N_7813,N_7965);
xnor U8089 (N_8089,N_7887,N_7856);
or U8090 (N_8090,N_7952,N_7932);
nand U8091 (N_8091,N_7884,N_7824);
or U8092 (N_8092,N_7912,N_7865);
nand U8093 (N_8093,N_7830,N_7805);
or U8094 (N_8094,N_7969,N_7896);
and U8095 (N_8095,N_7841,N_7918);
and U8096 (N_8096,N_7976,N_7800);
xnor U8097 (N_8097,N_7846,N_7961);
and U8098 (N_8098,N_7814,N_7991);
and U8099 (N_8099,N_7832,N_7922);
and U8100 (N_8100,N_7972,N_7911);
nor U8101 (N_8101,N_7815,N_7987);
nand U8102 (N_8102,N_7817,N_7914);
xor U8103 (N_8103,N_7902,N_7962);
nand U8104 (N_8104,N_7905,N_7929);
or U8105 (N_8105,N_7997,N_7822);
nand U8106 (N_8106,N_7883,N_7853);
nand U8107 (N_8107,N_7978,N_7919);
or U8108 (N_8108,N_7906,N_7876);
and U8109 (N_8109,N_7899,N_7952);
nor U8110 (N_8110,N_7901,N_7843);
or U8111 (N_8111,N_7976,N_7941);
and U8112 (N_8112,N_7961,N_7930);
or U8113 (N_8113,N_7949,N_7846);
xnor U8114 (N_8114,N_7983,N_7873);
and U8115 (N_8115,N_7842,N_7902);
or U8116 (N_8116,N_7911,N_7912);
nor U8117 (N_8117,N_7868,N_7850);
or U8118 (N_8118,N_7875,N_7808);
nand U8119 (N_8119,N_7909,N_7844);
nor U8120 (N_8120,N_7801,N_7996);
xor U8121 (N_8121,N_7841,N_7975);
and U8122 (N_8122,N_7992,N_7882);
xor U8123 (N_8123,N_7804,N_7997);
xor U8124 (N_8124,N_7810,N_7918);
xor U8125 (N_8125,N_7974,N_7914);
and U8126 (N_8126,N_7914,N_7868);
nor U8127 (N_8127,N_7844,N_7957);
nand U8128 (N_8128,N_7914,N_7819);
or U8129 (N_8129,N_7866,N_7978);
nand U8130 (N_8130,N_7943,N_7931);
nor U8131 (N_8131,N_7931,N_7970);
or U8132 (N_8132,N_7815,N_7980);
and U8133 (N_8133,N_7823,N_7998);
nor U8134 (N_8134,N_7986,N_7929);
nand U8135 (N_8135,N_7801,N_7886);
or U8136 (N_8136,N_7886,N_7924);
nand U8137 (N_8137,N_7978,N_7838);
nand U8138 (N_8138,N_7878,N_7818);
nor U8139 (N_8139,N_7976,N_7802);
or U8140 (N_8140,N_7883,N_7865);
nand U8141 (N_8141,N_7856,N_7838);
nand U8142 (N_8142,N_7890,N_7869);
and U8143 (N_8143,N_7891,N_7990);
and U8144 (N_8144,N_7920,N_7975);
xnor U8145 (N_8145,N_7955,N_7856);
xor U8146 (N_8146,N_7980,N_7838);
nand U8147 (N_8147,N_7880,N_7866);
or U8148 (N_8148,N_7981,N_7807);
nor U8149 (N_8149,N_7908,N_7862);
nor U8150 (N_8150,N_7800,N_7818);
nand U8151 (N_8151,N_7837,N_7937);
nand U8152 (N_8152,N_7961,N_7904);
xor U8153 (N_8153,N_7827,N_7834);
or U8154 (N_8154,N_7888,N_7979);
and U8155 (N_8155,N_7800,N_7903);
and U8156 (N_8156,N_7928,N_7877);
and U8157 (N_8157,N_7864,N_7874);
nand U8158 (N_8158,N_7999,N_7865);
or U8159 (N_8159,N_7935,N_7950);
nand U8160 (N_8160,N_7952,N_7886);
and U8161 (N_8161,N_7864,N_7961);
nor U8162 (N_8162,N_7890,N_7978);
nor U8163 (N_8163,N_7802,N_7961);
or U8164 (N_8164,N_7887,N_7842);
and U8165 (N_8165,N_7955,N_7887);
or U8166 (N_8166,N_7858,N_7803);
nand U8167 (N_8167,N_7950,N_7878);
and U8168 (N_8168,N_7845,N_7910);
nor U8169 (N_8169,N_7849,N_7844);
and U8170 (N_8170,N_7997,N_7925);
or U8171 (N_8171,N_7917,N_7811);
and U8172 (N_8172,N_7833,N_7943);
or U8173 (N_8173,N_7851,N_7864);
or U8174 (N_8174,N_7863,N_7864);
nand U8175 (N_8175,N_7879,N_7840);
nand U8176 (N_8176,N_7921,N_7868);
xnor U8177 (N_8177,N_7923,N_7928);
and U8178 (N_8178,N_7946,N_7897);
xnor U8179 (N_8179,N_7961,N_7967);
xor U8180 (N_8180,N_7843,N_7863);
and U8181 (N_8181,N_7964,N_7899);
xnor U8182 (N_8182,N_7937,N_7831);
nand U8183 (N_8183,N_7946,N_7846);
xnor U8184 (N_8184,N_7965,N_7885);
nor U8185 (N_8185,N_7851,N_7875);
and U8186 (N_8186,N_7951,N_7920);
and U8187 (N_8187,N_7815,N_7903);
xnor U8188 (N_8188,N_7854,N_7995);
xor U8189 (N_8189,N_7854,N_7835);
xor U8190 (N_8190,N_7820,N_7898);
or U8191 (N_8191,N_7801,N_7939);
xnor U8192 (N_8192,N_7931,N_7883);
nand U8193 (N_8193,N_7848,N_7934);
nand U8194 (N_8194,N_7884,N_7962);
xnor U8195 (N_8195,N_7934,N_7968);
nor U8196 (N_8196,N_7883,N_7862);
and U8197 (N_8197,N_7814,N_7979);
and U8198 (N_8198,N_7881,N_7837);
or U8199 (N_8199,N_7878,N_7881);
nor U8200 (N_8200,N_8028,N_8036);
or U8201 (N_8201,N_8189,N_8124);
nor U8202 (N_8202,N_8080,N_8181);
nand U8203 (N_8203,N_8040,N_8000);
nor U8204 (N_8204,N_8152,N_8017);
and U8205 (N_8205,N_8126,N_8053);
or U8206 (N_8206,N_8161,N_8035);
nor U8207 (N_8207,N_8003,N_8045);
or U8208 (N_8208,N_8113,N_8078);
or U8209 (N_8209,N_8052,N_8039);
nor U8210 (N_8210,N_8073,N_8074);
nand U8211 (N_8211,N_8015,N_8142);
or U8212 (N_8212,N_8058,N_8168);
or U8213 (N_8213,N_8199,N_8021);
nand U8214 (N_8214,N_8062,N_8197);
or U8215 (N_8215,N_8076,N_8125);
or U8216 (N_8216,N_8128,N_8115);
nand U8217 (N_8217,N_8091,N_8041);
nand U8218 (N_8218,N_8098,N_8042);
and U8219 (N_8219,N_8061,N_8109);
nand U8220 (N_8220,N_8046,N_8108);
or U8221 (N_8221,N_8008,N_8079);
nand U8222 (N_8222,N_8116,N_8044);
nor U8223 (N_8223,N_8056,N_8136);
xnor U8224 (N_8224,N_8153,N_8123);
nor U8225 (N_8225,N_8016,N_8112);
nor U8226 (N_8226,N_8166,N_8148);
nand U8227 (N_8227,N_8158,N_8081);
and U8228 (N_8228,N_8169,N_8025);
nor U8229 (N_8229,N_8160,N_8182);
or U8230 (N_8230,N_8100,N_8101);
nand U8231 (N_8231,N_8104,N_8192);
and U8232 (N_8232,N_8032,N_8065);
nor U8233 (N_8233,N_8095,N_8105);
nand U8234 (N_8234,N_8177,N_8193);
nor U8235 (N_8235,N_8180,N_8106);
or U8236 (N_8236,N_8110,N_8029);
xor U8237 (N_8237,N_8114,N_8048);
or U8238 (N_8238,N_8037,N_8075);
or U8239 (N_8239,N_8068,N_8127);
xnor U8240 (N_8240,N_8002,N_8111);
nand U8241 (N_8241,N_8157,N_8084);
xor U8242 (N_8242,N_8151,N_8122);
nand U8243 (N_8243,N_8140,N_8087);
and U8244 (N_8244,N_8130,N_8117);
and U8245 (N_8245,N_8069,N_8131);
nand U8246 (N_8246,N_8059,N_8072);
nor U8247 (N_8247,N_8156,N_8194);
xor U8248 (N_8248,N_8149,N_8171);
xor U8249 (N_8249,N_8012,N_8099);
nor U8250 (N_8250,N_8196,N_8185);
nor U8251 (N_8251,N_8162,N_8159);
nand U8252 (N_8252,N_8082,N_8150);
nand U8253 (N_8253,N_8179,N_8141);
or U8254 (N_8254,N_8018,N_8022);
nor U8255 (N_8255,N_8019,N_8092);
nor U8256 (N_8256,N_8007,N_8057);
and U8257 (N_8257,N_8147,N_8190);
nor U8258 (N_8258,N_8054,N_8013);
or U8259 (N_8259,N_8174,N_8173);
nand U8260 (N_8260,N_8031,N_8184);
or U8261 (N_8261,N_8067,N_8139);
nor U8262 (N_8262,N_8134,N_8055);
xor U8263 (N_8263,N_8186,N_8014);
or U8264 (N_8264,N_8027,N_8175);
xnor U8265 (N_8265,N_8102,N_8144);
and U8266 (N_8266,N_8183,N_8026);
xnor U8267 (N_8267,N_8083,N_8191);
or U8268 (N_8268,N_8088,N_8024);
and U8269 (N_8269,N_8006,N_8178);
and U8270 (N_8270,N_8132,N_8195);
xor U8271 (N_8271,N_8096,N_8135);
and U8272 (N_8272,N_8070,N_8143);
nand U8273 (N_8273,N_8138,N_8043);
and U8274 (N_8274,N_8077,N_8097);
nand U8275 (N_8275,N_8167,N_8085);
xor U8276 (N_8276,N_8063,N_8187);
xnor U8277 (N_8277,N_8107,N_8118);
or U8278 (N_8278,N_8064,N_8034);
nand U8279 (N_8279,N_8020,N_8001);
xor U8280 (N_8280,N_8093,N_8198);
or U8281 (N_8281,N_8155,N_8164);
and U8282 (N_8282,N_8011,N_8172);
or U8283 (N_8283,N_8009,N_8030);
nand U8284 (N_8284,N_8137,N_8121);
nand U8285 (N_8285,N_8010,N_8120);
nor U8286 (N_8286,N_8170,N_8119);
or U8287 (N_8287,N_8023,N_8071);
xnor U8288 (N_8288,N_8129,N_8094);
and U8289 (N_8289,N_8176,N_8050);
nor U8290 (N_8290,N_8154,N_8145);
and U8291 (N_8291,N_8033,N_8163);
nor U8292 (N_8292,N_8089,N_8165);
and U8293 (N_8293,N_8047,N_8049);
or U8294 (N_8294,N_8066,N_8004);
nand U8295 (N_8295,N_8038,N_8103);
nand U8296 (N_8296,N_8005,N_8051);
nor U8297 (N_8297,N_8060,N_8146);
or U8298 (N_8298,N_8086,N_8090);
nor U8299 (N_8299,N_8133,N_8188);
xnor U8300 (N_8300,N_8006,N_8169);
and U8301 (N_8301,N_8010,N_8091);
or U8302 (N_8302,N_8142,N_8084);
and U8303 (N_8303,N_8132,N_8087);
xor U8304 (N_8304,N_8073,N_8143);
nand U8305 (N_8305,N_8099,N_8008);
or U8306 (N_8306,N_8027,N_8192);
or U8307 (N_8307,N_8161,N_8098);
and U8308 (N_8308,N_8006,N_8168);
or U8309 (N_8309,N_8180,N_8174);
nor U8310 (N_8310,N_8041,N_8034);
or U8311 (N_8311,N_8047,N_8113);
nand U8312 (N_8312,N_8075,N_8108);
and U8313 (N_8313,N_8081,N_8172);
or U8314 (N_8314,N_8082,N_8145);
and U8315 (N_8315,N_8137,N_8172);
and U8316 (N_8316,N_8179,N_8053);
or U8317 (N_8317,N_8190,N_8083);
or U8318 (N_8318,N_8102,N_8198);
nand U8319 (N_8319,N_8039,N_8184);
nand U8320 (N_8320,N_8102,N_8087);
or U8321 (N_8321,N_8054,N_8122);
xnor U8322 (N_8322,N_8112,N_8078);
nor U8323 (N_8323,N_8042,N_8092);
or U8324 (N_8324,N_8014,N_8025);
or U8325 (N_8325,N_8001,N_8080);
and U8326 (N_8326,N_8071,N_8027);
and U8327 (N_8327,N_8022,N_8163);
nor U8328 (N_8328,N_8038,N_8069);
nand U8329 (N_8329,N_8017,N_8156);
or U8330 (N_8330,N_8092,N_8020);
nor U8331 (N_8331,N_8129,N_8190);
nand U8332 (N_8332,N_8034,N_8140);
and U8333 (N_8333,N_8126,N_8145);
and U8334 (N_8334,N_8166,N_8091);
xnor U8335 (N_8335,N_8049,N_8137);
nand U8336 (N_8336,N_8128,N_8191);
nand U8337 (N_8337,N_8004,N_8120);
nor U8338 (N_8338,N_8024,N_8015);
nor U8339 (N_8339,N_8006,N_8106);
nand U8340 (N_8340,N_8164,N_8192);
and U8341 (N_8341,N_8103,N_8055);
nand U8342 (N_8342,N_8122,N_8173);
xnor U8343 (N_8343,N_8182,N_8173);
and U8344 (N_8344,N_8076,N_8013);
xor U8345 (N_8345,N_8058,N_8050);
or U8346 (N_8346,N_8000,N_8024);
nor U8347 (N_8347,N_8031,N_8047);
nand U8348 (N_8348,N_8054,N_8021);
and U8349 (N_8349,N_8106,N_8162);
nor U8350 (N_8350,N_8104,N_8181);
xnor U8351 (N_8351,N_8178,N_8068);
nand U8352 (N_8352,N_8108,N_8064);
nand U8353 (N_8353,N_8086,N_8062);
nor U8354 (N_8354,N_8045,N_8110);
and U8355 (N_8355,N_8014,N_8197);
nand U8356 (N_8356,N_8032,N_8028);
nor U8357 (N_8357,N_8163,N_8105);
xnor U8358 (N_8358,N_8042,N_8137);
xnor U8359 (N_8359,N_8056,N_8029);
nor U8360 (N_8360,N_8004,N_8154);
and U8361 (N_8361,N_8109,N_8148);
and U8362 (N_8362,N_8147,N_8020);
or U8363 (N_8363,N_8050,N_8073);
nor U8364 (N_8364,N_8075,N_8089);
nand U8365 (N_8365,N_8077,N_8191);
nor U8366 (N_8366,N_8018,N_8001);
and U8367 (N_8367,N_8064,N_8169);
nand U8368 (N_8368,N_8069,N_8166);
nor U8369 (N_8369,N_8117,N_8082);
and U8370 (N_8370,N_8073,N_8171);
nor U8371 (N_8371,N_8012,N_8002);
and U8372 (N_8372,N_8086,N_8020);
and U8373 (N_8373,N_8186,N_8076);
nand U8374 (N_8374,N_8057,N_8152);
or U8375 (N_8375,N_8179,N_8168);
xnor U8376 (N_8376,N_8019,N_8069);
and U8377 (N_8377,N_8175,N_8038);
xor U8378 (N_8378,N_8112,N_8035);
and U8379 (N_8379,N_8103,N_8147);
or U8380 (N_8380,N_8035,N_8190);
or U8381 (N_8381,N_8150,N_8104);
nor U8382 (N_8382,N_8177,N_8170);
nand U8383 (N_8383,N_8111,N_8051);
and U8384 (N_8384,N_8031,N_8051);
xor U8385 (N_8385,N_8120,N_8083);
or U8386 (N_8386,N_8013,N_8187);
nand U8387 (N_8387,N_8127,N_8076);
nand U8388 (N_8388,N_8189,N_8135);
nand U8389 (N_8389,N_8117,N_8123);
nor U8390 (N_8390,N_8127,N_8049);
nor U8391 (N_8391,N_8167,N_8037);
xor U8392 (N_8392,N_8058,N_8008);
xnor U8393 (N_8393,N_8084,N_8115);
nand U8394 (N_8394,N_8029,N_8021);
nand U8395 (N_8395,N_8064,N_8092);
nor U8396 (N_8396,N_8004,N_8196);
nor U8397 (N_8397,N_8034,N_8167);
and U8398 (N_8398,N_8181,N_8043);
xor U8399 (N_8399,N_8160,N_8163);
xor U8400 (N_8400,N_8392,N_8314);
nor U8401 (N_8401,N_8223,N_8280);
or U8402 (N_8402,N_8332,N_8320);
nor U8403 (N_8403,N_8301,N_8368);
nor U8404 (N_8404,N_8380,N_8328);
nand U8405 (N_8405,N_8394,N_8272);
or U8406 (N_8406,N_8207,N_8202);
nand U8407 (N_8407,N_8307,N_8319);
and U8408 (N_8408,N_8325,N_8287);
and U8409 (N_8409,N_8347,N_8385);
nor U8410 (N_8410,N_8270,N_8267);
or U8411 (N_8411,N_8321,N_8208);
or U8412 (N_8412,N_8260,N_8311);
or U8413 (N_8413,N_8351,N_8342);
xor U8414 (N_8414,N_8290,N_8397);
or U8415 (N_8415,N_8323,N_8356);
xnor U8416 (N_8416,N_8211,N_8308);
nor U8417 (N_8417,N_8337,N_8206);
nand U8418 (N_8418,N_8256,N_8204);
nand U8419 (N_8419,N_8288,N_8292);
and U8420 (N_8420,N_8326,N_8276);
and U8421 (N_8421,N_8262,N_8216);
nand U8422 (N_8422,N_8361,N_8215);
or U8423 (N_8423,N_8239,N_8384);
or U8424 (N_8424,N_8212,N_8263);
or U8425 (N_8425,N_8379,N_8243);
nand U8426 (N_8426,N_8291,N_8362);
or U8427 (N_8427,N_8340,N_8315);
and U8428 (N_8428,N_8218,N_8217);
and U8429 (N_8429,N_8376,N_8274);
and U8430 (N_8430,N_8213,N_8357);
xor U8431 (N_8431,N_8284,N_8331);
xnor U8432 (N_8432,N_8247,N_8258);
nor U8433 (N_8433,N_8203,N_8341);
or U8434 (N_8434,N_8310,N_8309);
nand U8435 (N_8435,N_8220,N_8242);
or U8436 (N_8436,N_8378,N_8339);
or U8437 (N_8437,N_8387,N_8230);
or U8438 (N_8438,N_8396,N_8278);
and U8439 (N_8439,N_8312,N_8381);
or U8440 (N_8440,N_8344,N_8219);
nor U8441 (N_8441,N_8266,N_8214);
nand U8442 (N_8442,N_8329,N_8245);
nand U8443 (N_8443,N_8377,N_8373);
nor U8444 (N_8444,N_8236,N_8375);
nand U8445 (N_8445,N_8201,N_8244);
or U8446 (N_8446,N_8293,N_8285);
and U8447 (N_8447,N_8371,N_8228);
or U8448 (N_8448,N_8359,N_8277);
xor U8449 (N_8449,N_8333,N_8248);
nor U8450 (N_8450,N_8391,N_8393);
xor U8451 (N_8451,N_8388,N_8343);
and U8452 (N_8452,N_8327,N_8268);
or U8453 (N_8453,N_8295,N_8265);
nor U8454 (N_8454,N_8229,N_8350);
xnor U8455 (N_8455,N_8224,N_8313);
nand U8456 (N_8456,N_8364,N_8305);
and U8457 (N_8457,N_8296,N_8241);
and U8458 (N_8458,N_8238,N_8269);
nor U8459 (N_8459,N_8303,N_8281);
xnor U8460 (N_8460,N_8221,N_8358);
nand U8461 (N_8461,N_8317,N_8225);
and U8462 (N_8462,N_8318,N_8289);
nor U8463 (N_8463,N_8349,N_8257);
nand U8464 (N_8464,N_8246,N_8355);
nand U8465 (N_8465,N_8200,N_8226);
xnor U8466 (N_8466,N_8222,N_8300);
and U8467 (N_8467,N_8370,N_8336);
or U8468 (N_8468,N_8227,N_8297);
or U8469 (N_8469,N_8304,N_8275);
xnor U8470 (N_8470,N_8398,N_8240);
nand U8471 (N_8471,N_8210,N_8330);
nand U8472 (N_8472,N_8366,N_8382);
and U8473 (N_8473,N_8302,N_8250);
nand U8474 (N_8474,N_8252,N_8209);
xnor U8475 (N_8475,N_8259,N_8334);
xor U8476 (N_8476,N_8383,N_8205);
and U8477 (N_8477,N_8369,N_8298);
xor U8478 (N_8478,N_8365,N_8389);
nor U8479 (N_8479,N_8322,N_8360);
nor U8480 (N_8480,N_8251,N_8299);
and U8481 (N_8481,N_8237,N_8374);
or U8482 (N_8482,N_8346,N_8279);
or U8483 (N_8483,N_8254,N_8324);
and U8484 (N_8484,N_8372,N_8232);
xnor U8485 (N_8485,N_8255,N_8352);
nor U8486 (N_8486,N_8264,N_8335);
nor U8487 (N_8487,N_8353,N_8363);
nor U8488 (N_8488,N_8235,N_8286);
nand U8489 (N_8489,N_8231,N_8345);
and U8490 (N_8490,N_8261,N_8282);
nor U8491 (N_8491,N_8249,N_8395);
nor U8492 (N_8492,N_8348,N_8273);
nand U8493 (N_8493,N_8253,N_8233);
nand U8494 (N_8494,N_8338,N_8354);
nand U8495 (N_8495,N_8367,N_8294);
or U8496 (N_8496,N_8306,N_8316);
xor U8497 (N_8497,N_8390,N_8283);
nand U8498 (N_8498,N_8271,N_8386);
xor U8499 (N_8499,N_8234,N_8399);
nor U8500 (N_8500,N_8260,N_8316);
or U8501 (N_8501,N_8282,N_8249);
and U8502 (N_8502,N_8267,N_8341);
xor U8503 (N_8503,N_8387,N_8362);
nand U8504 (N_8504,N_8345,N_8240);
and U8505 (N_8505,N_8205,N_8225);
nor U8506 (N_8506,N_8261,N_8229);
nor U8507 (N_8507,N_8205,N_8385);
nand U8508 (N_8508,N_8267,N_8259);
and U8509 (N_8509,N_8272,N_8229);
nor U8510 (N_8510,N_8234,N_8212);
or U8511 (N_8511,N_8371,N_8345);
xnor U8512 (N_8512,N_8397,N_8311);
nand U8513 (N_8513,N_8282,N_8224);
nand U8514 (N_8514,N_8209,N_8297);
and U8515 (N_8515,N_8366,N_8274);
nand U8516 (N_8516,N_8367,N_8377);
nand U8517 (N_8517,N_8203,N_8332);
nor U8518 (N_8518,N_8336,N_8245);
or U8519 (N_8519,N_8321,N_8215);
xor U8520 (N_8520,N_8335,N_8324);
nand U8521 (N_8521,N_8279,N_8309);
nand U8522 (N_8522,N_8308,N_8398);
or U8523 (N_8523,N_8243,N_8370);
xor U8524 (N_8524,N_8301,N_8375);
nor U8525 (N_8525,N_8338,N_8207);
nor U8526 (N_8526,N_8370,N_8205);
nor U8527 (N_8527,N_8303,N_8290);
nor U8528 (N_8528,N_8285,N_8349);
nand U8529 (N_8529,N_8373,N_8298);
nand U8530 (N_8530,N_8327,N_8307);
nor U8531 (N_8531,N_8305,N_8223);
and U8532 (N_8532,N_8383,N_8399);
and U8533 (N_8533,N_8200,N_8264);
xor U8534 (N_8534,N_8282,N_8321);
and U8535 (N_8535,N_8267,N_8398);
nor U8536 (N_8536,N_8340,N_8221);
nor U8537 (N_8537,N_8233,N_8221);
and U8538 (N_8538,N_8261,N_8219);
xor U8539 (N_8539,N_8318,N_8220);
and U8540 (N_8540,N_8304,N_8331);
and U8541 (N_8541,N_8276,N_8318);
or U8542 (N_8542,N_8399,N_8329);
nand U8543 (N_8543,N_8393,N_8208);
nor U8544 (N_8544,N_8316,N_8364);
and U8545 (N_8545,N_8321,N_8357);
or U8546 (N_8546,N_8372,N_8307);
xnor U8547 (N_8547,N_8328,N_8297);
or U8548 (N_8548,N_8345,N_8356);
xor U8549 (N_8549,N_8286,N_8293);
nor U8550 (N_8550,N_8205,N_8333);
nor U8551 (N_8551,N_8244,N_8353);
or U8552 (N_8552,N_8215,N_8233);
xor U8553 (N_8553,N_8235,N_8296);
nand U8554 (N_8554,N_8293,N_8212);
and U8555 (N_8555,N_8205,N_8204);
xnor U8556 (N_8556,N_8337,N_8306);
or U8557 (N_8557,N_8257,N_8268);
and U8558 (N_8558,N_8237,N_8200);
nor U8559 (N_8559,N_8377,N_8368);
and U8560 (N_8560,N_8292,N_8201);
and U8561 (N_8561,N_8207,N_8232);
xor U8562 (N_8562,N_8203,N_8253);
nor U8563 (N_8563,N_8253,N_8284);
nor U8564 (N_8564,N_8312,N_8376);
and U8565 (N_8565,N_8393,N_8374);
or U8566 (N_8566,N_8207,N_8324);
and U8567 (N_8567,N_8218,N_8247);
or U8568 (N_8568,N_8232,N_8274);
or U8569 (N_8569,N_8360,N_8263);
xor U8570 (N_8570,N_8368,N_8254);
and U8571 (N_8571,N_8328,N_8334);
xnor U8572 (N_8572,N_8262,N_8314);
xnor U8573 (N_8573,N_8256,N_8299);
or U8574 (N_8574,N_8267,N_8324);
or U8575 (N_8575,N_8273,N_8266);
xor U8576 (N_8576,N_8269,N_8223);
nand U8577 (N_8577,N_8255,N_8267);
or U8578 (N_8578,N_8322,N_8218);
nand U8579 (N_8579,N_8354,N_8202);
or U8580 (N_8580,N_8261,N_8321);
nand U8581 (N_8581,N_8219,N_8331);
xnor U8582 (N_8582,N_8232,N_8255);
xnor U8583 (N_8583,N_8378,N_8282);
xor U8584 (N_8584,N_8326,N_8338);
and U8585 (N_8585,N_8283,N_8391);
or U8586 (N_8586,N_8302,N_8214);
and U8587 (N_8587,N_8242,N_8328);
xor U8588 (N_8588,N_8371,N_8301);
or U8589 (N_8589,N_8200,N_8262);
nand U8590 (N_8590,N_8325,N_8228);
nand U8591 (N_8591,N_8371,N_8251);
or U8592 (N_8592,N_8351,N_8314);
and U8593 (N_8593,N_8280,N_8367);
nor U8594 (N_8594,N_8307,N_8248);
nand U8595 (N_8595,N_8273,N_8392);
or U8596 (N_8596,N_8253,N_8393);
nor U8597 (N_8597,N_8247,N_8284);
nor U8598 (N_8598,N_8218,N_8314);
nor U8599 (N_8599,N_8337,N_8384);
and U8600 (N_8600,N_8445,N_8577);
nor U8601 (N_8601,N_8460,N_8440);
or U8602 (N_8602,N_8560,N_8478);
nor U8603 (N_8603,N_8527,N_8518);
xnor U8604 (N_8604,N_8463,N_8436);
xor U8605 (N_8605,N_8452,N_8568);
nor U8606 (N_8606,N_8465,N_8493);
or U8607 (N_8607,N_8596,N_8519);
or U8608 (N_8608,N_8488,N_8567);
or U8609 (N_8609,N_8513,N_8491);
and U8610 (N_8610,N_8544,N_8449);
xnor U8611 (N_8611,N_8403,N_8587);
and U8612 (N_8612,N_8459,N_8429);
nand U8613 (N_8613,N_8437,N_8581);
nor U8614 (N_8614,N_8433,N_8575);
or U8615 (N_8615,N_8594,N_8550);
xor U8616 (N_8616,N_8423,N_8599);
and U8617 (N_8617,N_8472,N_8509);
or U8618 (N_8618,N_8534,N_8516);
nand U8619 (N_8619,N_8483,N_8425);
or U8620 (N_8620,N_8554,N_8526);
nand U8621 (N_8621,N_8494,N_8521);
or U8622 (N_8622,N_8411,N_8466);
and U8623 (N_8623,N_8485,N_8502);
xnor U8624 (N_8624,N_8420,N_8572);
and U8625 (N_8625,N_8416,N_8474);
xnor U8626 (N_8626,N_8543,N_8563);
and U8627 (N_8627,N_8454,N_8541);
and U8628 (N_8628,N_8537,N_8515);
nand U8629 (N_8629,N_8582,N_8591);
or U8630 (N_8630,N_8573,N_8532);
nand U8631 (N_8631,N_8428,N_8588);
or U8632 (N_8632,N_8470,N_8487);
nand U8633 (N_8633,N_8476,N_8422);
nor U8634 (N_8634,N_8408,N_8432);
xnor U8635 (N_8635,N_8589,N_8566);
xnor U8636 (N_8636,N_8479,N_8451);
xor U8637 (N_8637,N_8542,N_8419);
or U8638 (N_8638,N_8512,N_8400);
and U8639 (N_8639,N_8435,N_8529);
nor U8640 (N_8640,N_8584,N_8505);
and U8641 (N_8641,N_8475,N_8503);
xor U8642 (N_8642,N_8414,N_8450);
nand U8643 (N_8643,N_8439,N_8536);
or U8644 (N_8644,N_8407,N_8525);
or U8645 (N_8645,N_8413,N_8576);
and U8646 (N_8646,N_8405,N_8480);
nor U8647 (N_8647,N_8421,N_8593);
xnor U8648 (N_8648,N_8524,N_8597);
and U8649 (N_8649,N_8580,N_8464);
or U8650 (N_8650,N_8548,N_8533);
nor U8651 (N_8651,N_8418,N_8511);
and U8652 (N_8652,N_8499,N_8402);
nand U8653 (N_8653,N_8583,N_8434);
xor U8654 (N_8654,N_8569,N_8453);
and U8655 (N_8655,N_8469,N_8562);
and U8656 (N_8656,N_8579,N_8517);
and U8657 (N_8657,N_8506,N_8553);
or U8658 (N_8658,N_8559,N_8424);
nand U8659 (N_8659,N_8508,N_8447);
xor U8660 (N_8660,N_8430,N_8496);
nand U8661 (N_8661,N_8590,N_8522);
nor U8662 (N_8662,N_8561,N_8442);
nand U8663 (N_8663,N_8549,N_8412);
or U8664 (N_8664,N_8482,N_8565);
nand U8665 (N_8665,N_8455,N_8486);
xor U8666 (N_8666,N_8443,N_8535);
nand U8667 (N_8667,N_8458,N_8426);
or U8668 (N_8668,N_8490,N_8586);
nor U8669 (N_8669,N_8415,N_8540);
xnor U8670 (N_8670,N_8547,N_8401);
and U8671 (N_8671,N_8545,N_8462);
or U8672 (N_8672,N_8539,N_8555);
or U8673 (N_8673,N_8523,N_8444);
xnor U8674 (N_8674,N_8551,N_8431);
and U8675 (N_8675,N_8552,N_8510);
and U8676 (N_8676,N_8564,N_8410);
xor U8677 (N_8677,N_8592,N_8473);
xor U8678 (N_8678,N_8484,N_8448);
and U8679 (N_8679,N_8595,N_8514);
nand U8680 (N_8680,N_8489,N_8500);
and U8681 (N_8681,N_8417,N_8504);
or U8682 (N_8682,N_8598,N_8531);
or U8683 (N_8683,N_8404,N_8409);
nand U8684 (N_8684,N_8446,N_8520);
nor U8685 (N_8685,N_8495,N_8477);
xor U8686 (N_8686,N_8481,N_8498);
nand U8687 (N_8687,N_8530,N_8497);
nor U8688 (N_8688,N_8471,N_8585);
nand U8689 (N_8689,N_8538,N_8507);
nand U8690 (N_8690,N_8461,N_8546);
or U8691 (N_8691,N_8406,N_8557);
nand U8692 (N_8692,N_8528,N_8492);
nor U8693 (N_8693,N_8438,N_8574);
or U8694 (N_8694,N_8467,N_8501);
and U8695 (N_8695,N_8570,N_8578);
and U8696 (N_8696,N_8558,N_8556);
or U8697 (N_8697,N_8456,N_8571);
nor U8698 (N_8698,N_8441,N_8427);
nor U8699 (N_8699,N_8468,N_8457);
nand U8700 (N_8700,N_8470,N_8544);
nor U8701 (N_8701,N_8586,N_8504);
nor U8702 (N_8702,N_8498,N_8516);
nor U8703 (N_8703,N_8565,N_8456);
and U8704 (N_8704,N_8542,N_8456);
xnor U8705 (N_8705,N_8467,N_8458);
nand U8706 (N_8706,N_8583,N_8527);
xor U8707 (N_8707,N_8439,N_8554);
nand U8708 (N_8708,N_8442,N_8451);
xnor U8709 (N_8709,N_8508,N_8583);
xor U8710 (N_8710,N_8569,N_8446);
xnor U8711 (N_8711,N_8517,N_8590);
nor U8712 (N_8712,N_8466,N_8437);
or U8713 (N_8713,N_8573,N_8425);
and U8714 (N_8714,N_8555,N_8482);
and U8715 (N_8715,N_8453,N_8497);
nand U8716 (N_8716,N_8586,N_8425);
nor U8717 (N_8717,N_8506,N_8401);
or U8718 (N_8718,N_8491,N_8585);
or U8719 (N_8719,N_8480,N_8568);
and U8720 (N_8720,N_8545,N_8586);
xor U8721 (N_8721,N_8508,N_8585);
and U8722 (N_8722,N_8423,N_8552);
xor U8723 (N_8723,N_8490,N_8540);
xnor U8724 (N_8724,N_8400,N_8509);
or U8725 (N_8725,N_8451,N_8500);
xnor U8726 (N_8726,N_8445,N_8513);
nand U8727 (N_8727,N_8542,N_8513);
xor U8728 (N_8728,N_8503,N_8517);
or U8729 (N_8729,N_8465,N_8529);
xor U8730 (N_8730,N_8421,N_8511);
and U8731 (N_8731,N_8431,N_8473);
or U8732 (N_8732,N_8447,N_8450);
or U8733 (N_8733,N_8584,N_8513);
and U8734 (N_8734,N_8527,N_8568);
and U8735 (N_8735,N_8490,N_8520);
nand U8736 (N_8736,N_8415,N_8471);
xnor U8737 (N_8737,N_8402,N_8421);
xor U8738 (N_8738,N_8569,N_8579);
nand U8739 (N_8739,N_8493,N_8529);
xor U8740 (N_8740,N_8508,N_8434);
nor U8741 (N_8741,N_8565,N_8537);
and U8742 (N_8742,N_8534,N_8544);
nor U8743 (N_8743,N_8545,N_8526);
or U8744 (N_8744,N_8584,N_8436);
nor U8745 (N_8745,N_8561,N_8599);
nor U8746 (N_8746,N_8597,N_8458);
and U8747 (N_8747,N_8518,N_8414);
xor U8748 (N_8748,N_8578,N_8420);
and U8749 (N_8749,N_8403,N_8457);
xnor U8750 (N_8750,N_8540,N_8492);
nor U8751 (N_8751,N_8583,N_8473);
xor U8752 (N_8752,N_8441,N_8518);
nor U8753 (N_8753,N_8563,N_8422);
nand U8754 (N_8754,N_8521,N_8405);
xnor U8755 (N_8755,N_8531,N_8499);
xnor U8756 (N_8756,N_8563,N_8520);
or U8757 (N_8757,N_8441,N_8543);
nor U8758 (N_8758,N_8462,N_8581);
or U8759 (N_8759,N_8493,N_8539);
xnor U8760 (N_8760,N_8450,N_8516);
xor U8761 (N_8761,N_8465,N_8503);
and U8762 (N_8762,N_8432,N_8477);
xnor U8763 (N_8763,N_8461,N_8506);
nor U8764 (N_8764,N_8558,N_8415);
and U8765 (N_8765,N_8533,N_8427);
xnor U8766 (N_8766,N_8581,N_8527);
nand U8767 (N_8767,N_8561,N_8495);
xnor U8768 (N_8768,N_8519,N_8575);
nand U8769 (N_8769,N_8498,N_8443);
nor U8770 (N_8770,N_8512,N_8545);
nand U8771 (N_8771,N_8572,N_8429);
or U8772 (N_8772,N_8559,N_8556);
nor U8773 (N_8773,N_8537,N_8550);
or U8774 (N_8774,N_8412,N_8424);
or U8775 (N_8775,N_8409,N_8412);
and U8776 (N_8776,N_8567,N_8462);
or U8777 (N_8777,N_8455,N_8538);
and U8778 (N_8778,N_8526,N_8556);
nor U8779 (N_8779,N_8491,N_8496);
nand U8780 (N_8780,N_8459,N_8469);
nor U8781 (N_8781,N_8523,N_8522);
nand U8782 (N_8782,N_8404,N_8434);
xor U8783 (N_8783,N_8456,N_8490);
nand U8784 (N_8784,N_8564,N_8519);
and U8785 (N_8785,N_8473,N_8404);
nand U8786 (N_8786,N_8596,N_8416);
nand U8787 (N_8787,N_8512,N_8427);
nor U8788 (N_8788,N_8585,N_8584);
nor U8789 (N_8789,N_8445,N_8414);
or U8790 (N_8790,N_8475,N_8488);
and U8791 (N_8791,N_8487,N_8549);
and U8792 (N_8792,N_8412,N_8464);
nor U8793 (N_8793,N_8581,N_8505);
nand U8794 (N_8794,N_8527,N_8434);
nor U8795 (N_8795,N_8472,N_8510);
or U8796 (N_8796,N_8446,N_8430);
nor U8797 (N_8797,N_8432,N_8526);
and U8798 (N_8798,N_8504,N_8584);
nor U8799 (N_8799,N_8550,N_8557);
nor U8800 (N_8800,N_8790,N_8786);
xnor U8801 (N_8801,N_8646,N_8607);
nand U8802 (N_8802,N_8793,N_8772);
or U8803 (N_8803,N_8675,N_8778);
nand U8804 (N_8804,N_8784,N_8659);
xnor U8805 (N_8805,N_8773,N_8791);
nand U8806 (N_8806,N_8750,N_8644);
nand U8807 (N_8807,N_8738,N_8737);
xnor U8808 (N_8808,N_8782,N_8679);
or U8809 (N_8809,N_8795,N_8765);
nor U8810 (N_8810,N_8726,N_8797);
nand U8811 (N_8811,N_8770,N_8693);
or U8812 (N_8812,N_8733,N_8724);
and U8813 (N_8813,N_8601,N_8688);
nand U8814 (N_8814,N_8613,N_8669);
nor U8815 (N_8815,N_8744,N_8749);
nand U8816 (N_8816,N_8605,N_8643);
xnor U8817 (N_8817,N_8704,N_8645);
xnor U8818 (N_8818,N_8624,N_8678);
nor U8819 (N_8819,N_8687,N_8794);
or U8820 (N_8820,N_8602,N_8742);
nor U8821 (N_8821,N_8676,N_8753);
nor U8822 (N_8822,N_8720,N_8682);
or U8823 (N_8823,N_8713,N_8691);
nor U8824 (N_8824,N_8660,N_8619);
xor U8825 (N_8825,N_8697,N_8756);
nand U8826 (N_8826,N_8684,N_8769);
xnor U8827 (N_8827,N_8783,N_8667);
or U8828 (N_8828,N_8734,N_8799);
or U8829 (N_8829,N_8730,N_8776);
xnor U8830 (N_8830,N_8774,N_8716);
nor U8831 (N_8831,N_8771,N_8775);
xor U8832 (N_8832,N_8761,N_8606);
nor U8833 (N_8833,N_8714,N_8677);
nor U8834 (N_8834,N_8694,N_8642);
nor U8835 (N_8835,N_8628,N_8664);
or U8836 (N_8836,N_8653,N_8681);
xor U8837 (N_8837,N_8666,N_8686);
xor U8838 (N_8838,N_8603,N_8729);
and U8839 (N_8839,N_8674,N_8708);
xnor U8840 (N_8840,N_8768,N_8746);
nor U8841 (N_8841,N_8719,N_8705);
nor U8842 (N_8842,N_8748,N_8710);
nand U8843 (N_8843,N_8661,N_8633);
nand U8844 (N_8844,N_8652,N_8608);
nor U8845 (N_8845,N_8760,N_8777);
nor U8846 (N_8846,N_8656,N_8610);
or U8847 (N_8847,N_8715,N_8609);
and U8848 (N_8848,N_8732,N_8792);
nor U8849 (N_8849,N_8703,N_8739);
xor U8850 (N_8850,N_8764,N_8701);
and U8851 (N_8851,N_8611,N_8709);
or U8852 (N_8852,N_8662,N_8717);
or U8853 (N_8853,N_8604,N_8759);
or U8854 (N_8854,N_8651,N_8630);
or U8855 (N_8855,N_8695,N_8683);
xor U8856 (N_8856,N_8627,N_8745);
nor U8857 (N_8857,N_8655,N_8740);
or U8858 (N_8858,N_8668,N_8623);
nor U8859 (N_8859,N_8672,N_8763);
or U8860 (N_8860,N_8625,N_8796);
and U8861 (N_8861,N_8685,N_8707);
and U8862 (N_8862,N_8781,N_8654);
nand U8863 (N_8863,N_8702,N_8629);
nor U8864 (N_8864,N_8754,N_8712);
or U8865 (N_8865,N_8618,N_8692);
xor U8866 (N_8866,N_8735,N_8725);
or U8867 (N_8867,N_8798,N_8673);
nand U8868 (N_8868,N_8638,N_8657);
xor U8869 (N_8869,N_8711,N_8757);
xnor U8870 (N_8870,N_8612,N_8658);
nand U8871 (N_8871,N_8785,N_8700);
and U8872 (N_8872,N_8640,N_8650);
nand U8873 (N_8873,N_8747,N_8758);
xor U8874 (N_8874,N_8788,N_8647);
nand U8875 (N_8875,N_8743,N_8698);
nor U8876 (N_8876,N_8752,N_8755);
xor U8877 (N_8877,N_8622,N_8649);
xor U8878 (N_8878,N_8637,N_8680);
and U8879 (N_8879,N_8736,N_8718);
and U8880 (N_8880,N_8648,N_8632);
xnor U8881 (N_8881,N_8780,N_8665);
xor U8882 (N_8882,N_8722,N_8614);
nor U8883 (N_8883,N_8689,N_8721);
nand U8884 (N_8884,N_8600,N_8617);
xor U8885 (N_8885,N_8731,N_8728);
nand U8886 (N_8886,N_8690,N_8615);
and U8887 (N_8887,N_8635,N_8766);
xor U8888 (N_8888,N_8620,N_8621);
nor U8889 (N_8889,N_8751,N_8671);
nand U8890 (N_8890,N_8787,N_8723);
and U8891 (N_8891,N_8639,N_8767);
or U8892 (N_8892,N_8616,N_8699);
nor U8893 (N_8893,N_8789,N_8634);
xnor U8894 (N_8894,N_8727,N_8663);
nand U8895 (N_8895,N_8741,N_8641);
nor U8896 (N_8896,N_8631,N_8779);
nor U8897 (N_8897,N_8626,N_8696);
or U8898 (N_8898,N_8762,N_8670);
xor U8899 (N_8899,N_8706,N_8636);
nor U8900 (N_8900,N_8735,N_8617);
nor U8901 (N_8901,N_8797,N_8799);
and U8902 (N_8902,N_8691,N_8637);
nor U8903 (N_8903,N_8675,N_8613);
and U8904 (N_8904,N_8748,N_8650);
nor U8905 (N_8905,N_8689,N_8685);
and U8906 (N_8906,N_8648,N_8732);
or U8907 (N_8907,N_8601,N_8748);
xor U8908 (N_8908,N_8693,N_8646);
and U8909 (N_8909,N_8687,N_8676);
and U8910 (N_8910,N_8650,N_8790);
and U8911 (N_8911,N_8659,N_8733);
nor U8912 (N_8912,N_8743,N_8714);
and U8913 (N_8913,N_8600,N_8798);
xnor U8914 (N_8914,N_8625,N_8684);
nand U8915 (N_8915,N_8756,N_8755);
and U8916 (N_8916,N_8648,N_8643);
nand U8917 (N_8917,N_8637,N_8606);
xnor U8918 (N_8918,N_8666,N_8695);
nand U8919 (N_8919,N_8695,N_8608);
or U8920 (N_8920,N_8708,N_8742);
xnor U8921 (N_8921,N_8699,N_8691);
nor U8922 (N_8922,N_8768,N_8680);
xnor U8923 (N_8923,N_8609,N_8608);
or U8924 (N_8924,N_8748,N_8608);
nand U8925 (N_8925,N_8637,N_8797);
nor U8926 (N_8926,N_8607,N_8704);
nor U8927 (N_8927,N_8703,N_8648);
nor U8928 (N_8928,N_8664,N_8780);
xor U8929 (N_8929,N_8796,N_8682);
and U8930 (N_8930,N_8658,N_8732);
and U8931 (N_8931,N_8678,N_8791);
xor U8932 (N_8932,N_8623,N_8692);
or U8933 (N_8933,N_8761,N_8668);
nand U8934 (N_8934,N_8762,N_8739);
or U8935 (N_8935,N_8729,N_8680);
and U8936 (N_8936,N_8772,N_8739);
or U8937 (N_8937,N_8607,N_8631);
nor U8938 (N_8938,N_8787,N_8781);
nand U8939 (N_8939,N_8636,N_8796);
nand U8940 (N_8940,N_8655,N_8738);
nor U8941 (N_8941,N_8673,N_8606);
nor U8942 (N_8942,N_8781,N_8695);
or U8943 (N_8943,N_8653,N_8749);
and U8944 (N_8944,N_8727,N_8640);
nand U8945 (N_8945,N_8748,N_8653);
or U8946 (N_8946,N_8702,N_8689);
xnor U8947 (N_8947,N_8612,N_8785);
nor U8948 (N_8948,N_8717,N_8785);
and U8949 (N_8949,N_8672,N_8666);
xor U8950 (N_8950,N_8691,N_8756);
or U8951 (N_8951,N_8771,N_8623);
nand U8952 (N_8952,N_8721,N_8755);
nand U8953 (N_8953,N_8625,N_8735);
and U8954 (N_8954,N_8744,N_8773);
nand U8955 (N_8955,N_8602,N_8693);
and U8956 (N_8956,N_8694,N_8726);
or U8957 (N_8957,N_8717,N_8675);
and U8958 (N_8958,N_8635,N_8657);
nor U8959 (N_8959,N_8714,N_8655);
or U8960 (N_8960,N_8711,N_8681);
and U8961 (N_8961,N_8708,N_8795);
and U8962 (N_8962,N_8650,N_8775);
xnor U8963 (N_8963,N_8607,N_8691);
nand U8964 (N_8964,N_8725,N_8729);
xor U8965 (N_8965,N_8677,N_8698);
xor U8966 (N_8966,N_8764,N_8643);
or U8967 (N_8967,N_8658,N_8778);
nand U8968 (N_8968,N_8781,N_8692);
and U8969 (N_8969,N_8734,N_8694);
nor U8970 (N_8970,N_8683,N_8657);
nor U8971 (N_8971,N_8683,N_8765);
xnor U8972 (N_8972,N_8615,N_8786);
xor U8973 (N_8973,N_8673,N_8646);
and U8974 (N_8974,N_8653,N_8739);
nand U8975 (N_8975,N_8721,N_8624);
and U8976 (N_8976,N_8662,N_8653);
or U8977 (N_8977,N_8618,N_8757);
nor U8978 (N_8978,N_8635,N_8628);
xnor U8979 (N_8979,N_8795,N_8633);
nor U8980 (N_8980,N_8638,N_8743);
or U8981 (N_8981,N_8739,N_8727);
and U8982 (N_8982,N_8744,N_8730);
nor U8983 (N_8983,N_8642,N_8727);
or U8984 (N_8984,N_8677,N_8702);
xnor U8985 (N_8985,N_8711,N_8749);
or U8986 (N_8986,N_8773,N_8655);
and U8987 (N_8987,N_8680,N_8635);
nor U8988 (N_8988,N_8625,N_8777);
xor U8989 (N_8989,N_8795,N_8639);
and U8990 (N_8990,N_8662,N_8722);
nor U8991 (N_8991,N_8672,N_8704);
and U8992 (N_8992,N_8781,N_8641);
or U8993 (N_8993,N_8650,N_8660);
xor U8994 (N_8994,N_8634,N_8646);
nand U8995 (N_8995,N_8717,N_8671);
and U8996 (N_8996,N_8763,N_8609);
and U8997 (N_8997,N_8696,N_8732);
nand U8998 (N_8998,N_8715,N_8719);
xor U8999 (N_8999,N_8695,N_8696);
or U9000 (N_9000,N_8979,N_8863);
nor U9001 (N_9001,N_8833,N_8852);
or U9002 (N_9002,N_8871,N_8883);
nor U9003 (N_9003,N_8998,N_8855);
xnor U9004 (N_9004,N_8888,N_8943);
xor U9005 (N_9005,N_8958,N_8927);
and U9006 (N_9006,N_8974,N_8995);
or U9007 (N_9007,N_8886,N_8975);
or U9008 (N_9008,N_8938,N_8894);
xnor U9009 (N_9009,N_8844,N_8820);
nand U9010 (N_9010,N_8857,N_8937);
xnor U9011 (N_9011,N_8895,N_8905);
or U9012 (N_9012,N_8846,N_8824);
nand U9013 (N_9013,N_8869,N_8990);
and U9014 (N_9014,N_8916,N_8813);
and U9015 (N_9015,N_8940,N_8967);
nand U9016 (N_9016,N_8877,N_8887);
nand U9017 (N_9017,N_8901,N_8814);
and U9018 (N_9018,N_8802,N_8851);
and U9019 (N_9019,N_8865,N_8956);
nand U9020 (N_9020,N_8915,N_8910);
nand U9021 (N_9021,N_8931,N_8948);
nand U9022 (N_9022,N_8996,N_8930);
xor U9023 (N_9023,N_8989,N_8929);
nor U9024 (N_9024,N_8973,N_8939);
or U9025 (N_9025,N_8896,N_8983);
xnor U9026 (N_9026,N_8840,N_8897);
and U9027 (N_9027,N_8932,N_8864);
and U9028 (N_9028,N_8841,N_8837);
xor U9029 (N_9029,N_8988,N_8891);
nand U9030 (N_9030,N_8914,N_8853);
xnor U9031 (N_9031,N_8810,N_8811);
nor U9032 (N_9032,N_8859,N_8923);
or U9033 (N_9033,N_8982,N_8807);
nor U9034 (N_9034,N_8893,N_8961);
xor U9035 (N_9035,N_8868,N_8843);
nand U9036 (N_9036,N_8992,N_8816);
xor U9037 (N_9037,N_8968,N_8993);
nand U9038 (N_9038,N_8866,N_8913);
xor U9039 (N_9039,N_8918,N_8952);
xor U9040 (N_9040,N_8953,N_8904);
nor U9041 (N_9041,N_8827,N_8823);
and U9042 (N_9042,N_8994,N_8838);
nand U9043 (N_9043,N_8959,N_8903);
nand U9044 (N_9044,N_8933,N_8858);
nor U9045 (N_9045,N_8861,N_8972);
and U9046 (N_9046,N_8856,N_8954);
or U9047 (N_9047,N_8890,N_8834);
xor U9048 (N_9048,N_8951,N_8819);
nor U9049 (N_9049,N_8808,N_8806);
nand U9050 (N_9050,N_8809,N_8970);
nor U9051 (N_9051,N_8925,N_8980);
and U9052 (N_9052,N_8825,N_8965);
and U9053 (N_9053,N_8949,N_8950);
xor U9054 (N_9054,N_8902,N_8900);
nor U9055 (N_9055,N_8885,N_8804);
or U9056 (N_9056,N_8997,N_8971);
and U9057 (N_9057,N_8935,N_8874);
and U9058 (N_9058,N_8978,N_8981);
nor U9059 (N_9059,N_8803,N_8942);
nor U9060 (N_9060,N_8960,N_8977);
or U9061 (N_9061,N_8907,N_8830);
nand U9062 (N_9062,N_8876,N_8831);
or U9063 (N_9063,N_8991,N_8870);
xnor U9064 (N_9064,N_8862,N_8867);
nand U9065 (N_9065,N_8828,N_8842);
or U9066 (N_9066,N_8800,N_8815);
nor U9067 (N_9067,N_8878,N_8919);
and U9068 (N_9068,N_8926,N_8873);
nand U9069 (N_9069,N_8821,N_8836);
xor U9070 (N_9070,N_8839,N_8964);
and U9071 (N_9071,N_8872,N_8880);
nand U9072 (N_9072,N_8899,N_8969);
xor U9073 (N_9073,N_8922,N_8928);
xor U9074 (N_9074,N_8832,N_8829);
and U9075 (N_9075,N_8879,N_8892);
nand U9076 (N_9076,N_8860,N_8850);
nor U9077 (N_9077,N_8917,N_8884);
nor U9078 (N_9078,N_8962,N_8845);
or U9079 (N_9079,N_8805,N_8875);
xor U9080 (N_9080,N_8906,N_8944);
nor U9081 (N_9081,N_8945,N_8847);
and U9082 (N_9082,N_8882,N_8955);
xor U9083 (N_9083,N_8848,N_8889);
nand U9084 (N_9084,N_8921,N_8911);
xnor U9085 (N_9085,N_8854,N_8812);
nor U9086 (N_9086,N_8924,N_8985);
xnor U9087 (N_9087,N_8966,N_8818);
nand U9088 (N_9088,N_8881,N_8947);
and U9089 (N_9089,N_8912,N_8849);
or U9090 (N_9090,N_8801,N_8941);
or U9091 (N_9091,N_8934,N_8999);
or U9092 (N_9092,N_8817,N_8946);
nor U9093 (N_9093,N_8963,N_8909);
nor U9094 (N_9094,N_8987,N_8976);
nor U9095 (N_9095,N_8822,N_8984);
xor U9096 (N_9096,N_8835,N_8986);
and U9097 (N_9097,N_8920,N_8908);
nor U9098 (N_9098,N_8957,N_8936);
nand U9099 (N_9099,N_8898,N_8826);
nor U9100 (N_9100,N_8900,N_8825);
or U9101 (N_9101,N_8937,N_8992);
xnor U9102 (N_9102,N_8825,N_8845);
nor U9103 (N_9103,N_8871,N_8811);
xnor U9104 (N_9104,N_8932,N_8926);
or U9105 (N_9105,N_8897,N_8969);
xnor U9106 (N_9106,N_8909,N_8890);
nand U9107 (N_9107,N_8866,N_8951);
xnor U9108 (N_9108,N_8873,N_8909);
nand U9109 (N_9109,N_8989,N_8925);
nor U9110 (N_9110,N_8825,N_8820);
nand U9111 (N_9111,N_8878,N_8979);
nor U9112 (N_9112,N_8984,N_8971);
and U9113 (N_9113,N_8938,N_8915);
and U9114 (N_9114,N_8863,N_8847);
xor U9115 (N_9115,N_8855,N_8890);
or U9116 (N_9116,N_8894,N_8812);
and U9117 (N_9117,N_8800,N_8871);
or U9118 (N_9118,N_8958,N_8952);
xor U9119 (N_9119,N_8907,N_8924);
xor U9120 (N_9120,N_8875,N_8857);
and U9121 (N_9121,N_8970,N_8875);
xor U9122 (N_9122,N_8831,N_8843);
or U9123 (N_9123,N_8952,N_8896);
nand U9124 (N_9124,N_8803,N_8801);
xor U9125 (N_9125,N_8915,N_8830);
xnor U9126 (N_9126,N_8841,N_8955);
or U9127 (N_9127,N_8907,N_8958);
xor U9128 (N_9128,N_8872,N_8811);
nor U9129 (N_9129,N_8987,N_8824);
nor U9130 (N_9130,N_8824,N_8898);
nor U9131 (N_9131,N_8996,N_8879);
nand U9132 (N_9132,N_8964,N_8969);
or U9133 (N_9133,N_8914,N_8841);
or U9134 (N_9134,N_8900,N_8953);
nand U9135 (N_9135,N_8959,N_8972);
and U9136 (N_9136,N_8990,N_8804);
nand U9137 (N_9137,N_8931,N_8912);
nand U9138 (N_9138,N_8965,N_8929);
nand U9139 (N_9139,N_8825,N_8864);
and U9140 (N_9140,N_8860,N_8890);
or U9141 (N_9141,N_8844,N_8848);
or U9142 (N_9142,N_8830,N_8839);
nand U9143 (N_9143,N_8998,N_8971);
or U9144 (N_9144,N_8979,N_8987);
xnor U9145 (N_9145,N_8950,N_8882);
xnor U9146 (N_9146,N_8982,N_8827);
nor U9147 (N_9147,N_8833,N_8952);
xnor U9148 (N_9148,N_8806,N_8846);
nor U9149 (N_9149,N_8807,N_8887);
nor U9150 (N_9150,N_8905,N_8844);
nand U9151 (N_9151,N_8888,N_8911);
xnor U9152 (N_9152,N_8802,N_8907);
nor U9153 (N_9153,N_8803,N_8959);
xnor U9154 (N_9154,N_8865,N_8901);
nand U9155 (N_9155,N_8992,N_8952);
or U9156 (N_9156,N_8827,N_8957);
nand U9157 (N_9157,N_8915,N_8927);
xor U9158 (N_9158,N_8949,N_8913);
and U9159 (N_9159,N_8893,N_8932);
or U9160 (N_9160,N_8800,N_8918);
and U9161 (N_9161,N_8844,N_8851);
or U9162 (N_9162,N_8936,N_8843);
or U9163 (N_9163,N_8881,N_8904);
or U9164 (N_9164,N_8977,N_8846);
or U9165 (N_9165,N_8915,N_8991);
nor U9166 (N_9166,N_8993,N_8960);
nand U9167 (N_9167,N_8827,N_8869);
and U9168 (N_9168,N_8877,N_8865);
nand U9169 (N_9169,N_8863,N_8981);
and U9170 (N_9170,N_8842,N_8964);
xor U9171 (N_9171,N_8819,N_8911);
nor U9172 (N_9172,N_8893,N_8971);
and U9173 (N_9173,N_8914,N_8924);
and U9174 (N_9174,N_8996,N_8868);
and U9175 (N_9175,N_8880,N_8955);
xnor U9176 (N_9176,N_8869,N_8823);
and U9177 (N_9177,N_8985,N_8889);
or U9178 (N_9178,N_8858,N_8807);
xnor U9179 (N_9179,N_8835,N_8991);
or U9180 (N_9180,N_8814,N_8957);
and U9181 (N_9181,N_8989,N_8802);
xnor U9182 (N_9182,N_8943,N_8897);
and U9183 (N_9183,N_8883,N_8862);
nor U9184 (N_9184,N_8828,N_8874);
and U9185 (N_9185,N_8967,N_8982);
nand U9186 (N_9186,N_8977,N_8908);
nand U9187 (N_9187,N_8831,N_8812);
xor U9188 (N_9188,N_8880,N_8924);
and U9189 (N_9189,N_8865,N_8894);
nor U9190 (N_9190,N_8821,N_8867);
nor U9191 (N_9191,N_8975,N_8996);
nand U9192 (N_9192,N_8826,N_8933);
or U9193 (N_9193,N_8956,N_8811);
nand U9194 (N_9194,N_8898,N_8916);
nor U9195 (N_9195,N_8857,N_8926);
xor U9196 (N_9196,N_8856,N_8992);
and U9197 (N_9197,N_8855,N_8812);
nor U9198 (N_9198,N_8999,N_8936);
xnor U9199 (N_9199,N_8812,N_8961);
and U9200 (N_9200,N_9109,N_9165);
xor U9201 (N_9201,N_9160,N_9151);
nand U9202 (N_9202,N_9156,N_9054);
nor U9203 (N_9203,N_9002,N_9123);
or U9204 (N_9204,N_9147,N_9001);
nand U9205 (N_9205,N_9133,N_9162);
and U9206 (N_9206,N_9188,N_9115);
and U9207 (N_9207,N_9034,N_9041);
nand U9208 (N_9208,N_9149,N_9171);
and U9209 (N_9209,N_9050,N_9182);
nand U9210 (N_9210,N_9010,N_9022);
and U9211 (N_9211,N_9150,N_9015);
or U9212 (N_9212,N_9076,N_9102);
xnor U9213 (N_9213,N_9166,N_9183);
and U9214 (N_9214,N_9093,N_9044);
xnor U9215 (N_9215,N_9028,N_9191);
and U9216 (N_9216,N_9037,N_9058);
nand U9217 (N_9217,N_9040,N_9027);
or U9218 (N_9218,N_9060,N_9161);
or U9219 (N_9219,N_9023,N_9018);
or U9220 (N_9220,N_9189,N_9116);
or U9221 (N_9221,N_9005,N_9113);
nor U9222 (N_9222,N_9007,N_9118);
nand U9223 (N_9223,N_9091,N_9006);
and U9224 (N_9224,N_9198,N_9132);
or U9225 (N_9225,N_9124,N_9197);
nand U9226 (N_9226,N_9057,N_9142);
nor U9227 (N_9227,N_9143,N_9145);
xor U9228 (N_9228,N_9019,N_9013);
and U9229 (N_9229,N_9032,N_9033);
nand U9230 (N_9230,N_9186,N_9095);
or U9231 (N_9231,N_9167,N_9069);
nor U9232 (N_9232,N_9101,N_9021);
and U9233 (N_9233,N_9117,N_9099);
or U9234 (N_9234,N_9055,N_9114);
and U9235 (N_9235,N_9092,N_9046);
nor U9236 (N_9236,N_9164,N_9187);
nand U9237 (N_9237,N_9084,N_9119);
nor U9238 (N_9238,N_9077,N_9094);
and U9239 (N_9239,N_9081,N_9185);
or U9240 (N_9240,N_9129,N_9126);
or U9241 (N_9241,N_9112,N_9163);
nor U9242 (N_9242,N_9063,N_9088);
and U9243 (N_9243,N_9194,N_9078);
xnor U9244 (N_9244,N_9031,N_9025);
and U9245 (N_9245,N_9174,N_9008);
nor U9246 (N_9246,N_9157,N_9135);
and U9247 (N_9247,N_9098,N_9184);
nor U9248 (N_9248,N_9085,N_9103);
nand U9249 (N_9249,N_9036,N_9053);
xnor U9250 (N_9250,N_9175,N_9065);
and U9251 (N_9251,N_9111,N_9043);
nand U9252 (N_9252,N_9047,N_9072);
nand U9253 (N_9253,N_9169,N_9153);
nand U9254 (N_9254,N_9170,N_9056);
or U9255 (N_9255,N_9154,N_9104);
nor U9256 (N_9256,N_9136,N_9079);
nor U9257 (N_9257,N_9139,N_9075);
xnor U9258 (N_9258,N_9089,N_9176);
xor U9259 (N_9259,N_9090,N_9066);
nand U9260 (N_9260,N_9049,N_9180);
and U9261 (N_9261,N_9140,N_9070);
nand U9262 (N_9262,N_9029,N_9106);
nor U9263 (N_9263,N_9062,N_9148);
nor U9264 (N_9264,N_9181,N_9000);
or U9265 (N_9265,N_9042,N_9038);
nor U9266 (N_9266,N_9128,N_9012);
xor U9267 (N_9267,N_9087,N_9178);
or U9268 (N_9268,N_9100,N_9193);
nor U9269 (N_9269,N_9141,N_9080);
and U9270 (N_9270,N_9120,N_9035);
nor U9271 (N_9271,N_9177,N_9097);
and U9272 (N_9272,N_9026,N_9144);
or U9273 (N_9273,N_9004,N_9039);
and U9274 (N_9274,N_9024,N_9146);
nor U9275 (N_9275,N_9061,N_9196);
xor U9276 (N_9276,N_9125,N_9108);
nand U9277 (N_9277,N_9159,N_9030);
xnor U9278 (N_9278,N_9199,N_9017);
nand U9279 (N_9279,N_9020,N_9195);
nand U9280 (N_9280,N_9122,N_9064);
or U9281 (N_9281,N_9009,N_9011);
nand U9282 (N_9282,N_9045,N_9134);
xor U9283 (N_9283,N_9068,N_9096);
and U9284 (N_9284,N_9168,N_9073);
nand U9285 (N_9285,N_9158,N_9074);
and U9286 (N_9286,N_9105,N_9110);
xor U9287 (N_9287,N_9172,N_9052);
or U9288 (N_9288,N_9016,N_9179);
nor U9289 (N_9289,N_9071,N_9131);
or U9290 (N_9290,N_9086,N_9014);
nand U9291 (N_9291,N_9083,N_9059);
and U9292 (N_9292,N_9190,N_9152);
xor U9293 (N_9293,N_9137,N_9003);
and U9294 (N_9294,N_9082,N_9192);
nand U9295 (N_9295,N_9155,N_9121);
nand U9296 (N_9296,N_9138,N_9051);
and U9297 (N_9297,N_9130,N_9173);
nor U9298 (N_9298,N_9107,N_9127);
nand U9299 (N_9299,N_9048,N_9067);
and U9300 (N_9300,N_9175,N_9070);
or U9301 (N_9301,N_9166,N_9129);
or U9302 (N_9302,N_9074,N_9119);
or U9303 (N_9303,N_9070,N_9049);
or U9304 (N_9304,N_9119,N_9144);
nand U9305 (N_9305,N_9080,N_9108);
and U9306 (N_9306,N_9173,N_9001);
nand U9307 (N_9307,N_9093,N_9005);
xor U9308 (N_9308,N_9177,N_9168);
nand U9309 (N_9309,N_9092,N_9131);
nand U9310 (N_9310,N_9029,N_9003);
nand U9311 (N_9311,N_9007,N_9135);
xor U9312 (N_9312,N_9009,N_9072);
and U9313 (N_9313,N_9162,N_9116);
xnor U9314 (N_9314,N_9037,N_9065);
nor U9315 (N_9315,N_9021,N_9170);
and U9316 (N_9316,N_9093,N_9104);
xnor U9317 (N_9317,N_9044,N_9139);
or U9318 (N_9318,N_9072,N_9198);
xor U9319 (N_9319,N_9098,N_9144);
and U9320 (N_9320,N_9096,N_9082);
and U9321 (N_9321,N_9132,N_9013);
nand U9322 (N_9322,N_9166,N_9132);
and U9323 (N_9323,N_9070,N_9013);
xnor U9324 (N_9324,N_9139,N_9116);
xor U9325 (N_9325,N_9038,N_9003);
xnor U9326 (N_9326,N_9087,N_9113);
xnor U9327 (N_9327,N_9036,N_9160);
nand U9328 (N_9328,N_9156,N_9137);
and U9329 (N_9329,N_9014,N_9137);
nand U9330 (N_9330,N_9097,N_9125);
nor U9331 (N_9331,N_9053,N_9163);
nor U9332 (N_9332,N_9097,N_9020);
xor U9333 (N_9333,N_9098,N_9191);
and U9334 (N_9334,N_9009,N_9153);
nand U9335 (N_9335,N_9191,N_9048);
nand U9336 (N_9336,N_9115,N_9156);
nor U9337 (N_9337,N_9003,N_9076);
or U9338 (N_9338,N_9093,N_9171);
nand U9339 (N_9339,N_9003,N_9167);
xnor U9340 (N_9340,N_9187,N_9094);
nor U9341 (N_9341,N_9112,N_9062);
nor U9342 (N_9342,N_9173,N_9195);
or U9343 (N_9343,N_9148,N_9084);
nand U9344 (N_9344,N_9045,N_9111);
nand U9345 (N_9345,N_9191,N_9125);
xnor U9346 (N_9346,N_9053,N_9002);
xnor U9347 (N_9347,N_9177,N_9092);
nor U9348 (N_9348,N_9049,N_9127);
nor U9349 (N_9349,N_9105,N_9050);
xnor U9350 (N_9350,N_9091,N_9043);
and U9351 (N_9351,N_9134,N_9173);
or U9352 (N_9352,N_9094,N_9121);
nor U9353 (N_9353,N_9183,N_9160);
and U9354 (N_9354,N_9064,N_9137);
and U9355 (N_9355,N_9131,N_9097);
xnor U9356 (N_9356,N_9041,N_9139);
xnor U9357 (N_9357,N_9044,N_9094);
nand U9358 (N_9358,N_9034,N_9035);
and U9359 (N_9359,N_9139,N_9101);
nor U9360 (N_9360,N_9170,N_9086);
nand U9361 (N_9361,N_9051,N_9007);
nor U9362 (N_9362,N_9019,N_9052);
nor U9363 (N_9363,N_9083,N_9155);
nand U9364 (N_9364,N_9060,N_9064);
nor U9365 (N_9365,N_9038,N_9028);
nand U9366 (N_9366,N_9169,N_9180);
xnor U9367 (N_9367,N_9108,N_9156);
or U9368 (N_9368,N_9187,N_9001);
xnor U9369 (N_9369,N_9134,N_9168);
xor U9370 (N_9370,N_9180,N_9117);
nand U9371 (N_9371,N_9169,N_9170);
and U9372 (N_9372,N_9069,N_9004);
nor U9373 (N_9373,N_9158,N_9153);
or U9374 (N_9374,N_9186,N_9125);
and U9375 (N_9375,N_9195,N_9076);
nor U9376 (N_9376,N_9044,N_9095);
and U9377 (N_9377,N_9168,N_9194);
and U9378 (N_9378,N_9095,N_9137);
xnor U9379 (N_9379,N_9149,N_9045);
or U9380 (N_9380,N_9066,N_9010);
nor U9381 (N_9381,N_9024,N_9014);
nor U9382 (N_9382,N_9050,N_9086);
nand U9383 (N_9383,N_9015,N_9062);
xor U9384 (N_9384,N_9003,N_9008);
nand U9385 (N_9385,N_9077,N_9148);
and U9386 (N_9386,N_9156,N_9165);
xnor U9387 (N_9387,N_9082,N_9088);
xor U9388 (N_9388,N_9106,N_9006);
or U9389 (N_9389,N_9052,N_9020);
nor U9390 (N_9390,N_9154,N_9047);
nand U9391 (N_9391,N_9048,N_9070);
and U9392 (N_9392,N_9127,N_9093);
nor U9393 (N_9393,N_9193,N_9049);
xor U9394 (N_9394,N_9131,N_9143);
or U9395 (N_9395,N_9049,N_9196);
nand U9396 (N_9396,N_9131,N_9045);
xor U9397 (N_9397,N_9016,N_9170);
and U9398 (N_9398,N_9147,N_9130);
nor U9399 (N_9399,N_9006,N_9086);
xnor U9400 (N_9400,N_9350,N_9310);
xor U9401 (N_9401,N_9343,N_9263);
xnor U9402 (N_9402,N_9398,N_9209);
nand U9403 (N_9403,N_9237,N_9212);
and U9404 (N_9404,N_9392,N_9359);
and U9405 (N_9405,N_9260,N_9293);
and U9406 (N_9406,N_9201,N_9228);
nor U9407 (N_9407,N_9240,N_9313);
xor U9408 (N_9408,N_9235,N_9262);
xor U9409 (N_9409,N_9290,N_9364);
nand U9410 (N_9410,N_9383,N_9214);
or U9411 (N_9411,N_9251,N_9394);
xor U9412 (N_9412,N_9238,N_9337);
or U9413 (N_9413,N_9381,N_9275);
nand U9414 (N_9414,N_9219,N_9304);
xor U9415 (N_9415,N_9215,N_9236);
xor U9416 (N_9416,N_9301,N_9233);
or U9417 (N_9417,N_9250,N_9306);
and U9418 (N_9418,N_9245,N_9362);
nor U9419 (N_9419,N_9255,N_9295);
nor U9420 (N_9420,N_9248,N_9361);
or U9421 (N_9421,N_9277,N_9208);
and U9422 (N_9422,N_9285,N_9323);
nor U9423 (N_9423,N_9229,N_9391);
xor U9424 (N_9424,N_9396,N_9281);
nor U9425 (N_9425,N_9375,N_9230);
and U9426 (N_9426,N_9355,N_9356);
or U9427 (N_9427,N_9202,N_9234);
xor U9428 (N_9428,N_9397,N_9328);
nor U9429 (N_9429,N_9311,N_9376);
and U9430 (N_9430,N_9268,N_9210);
and U9431 (N_9431,N_9252,N_9284);
xnor U9432 (N_9432,N_9274,N_9385);
and U9433 (N_9433,N_9247,N_9374);
or U9434 (N_9434,N_9388,N_9336);
nor U9435 (N_9435,N_9371,N_9267);
and U9436 (N_9436,N_9324,N_9349);
nand U9437 (N_9437,N_9283,N_9276);
and U9438 (N_9438,N_9205,N_9242);
nor U9439 (N_9439,N_9367,N_9315);
or U9440 (N_9440,N_9372,N_9272);
and U9441 (N_9441,N_9271,N_9317);
nor U9442 (N_9442,N_9329,N_9338);
nor U9443 (N_9443,N_9206,N_9342);
nor U9444 (N_9444,N_9339,N_9207);
nand U9445 (N_9445,N_9270,N_9232);
and U9446 (N_9446,N_9300,N_9340);
or U9447 (N_9447,N_9280,N_9273);
nor U9448 (N_9448,N_9395,N_9389);
nand U9449 (N_9449,N_9223,N_9382);
and U9450 (N_9450,N_9211,N_9370);
xor U9451 (N_9451,N_9312,N_9200);
xnor U9452 (N_9452,N_9261,N_9390);
and U9453 (N_9453,N_9373,N_9341);
nand U9454 (N_9454,N_9241,N_9256);
and U9455 (N_9455,N_9365,N_9298);
nor U9456 (N_9456,N_9353,N_9279);
xnor U9457 (N_9457,N_9243,N_9326);
or U9458 (N_9458,N_9278,N_9331);
or U9459 (N_9459,N_9226,N_9258);
nor U9460 (N_9460,N_9327,N_9282);
or U9461 (N_9461,N_9308,N_9369);
nand U9462 (N_9462,N_9358,N_9354);
xnor U9463 (N_9463,N_9286,N_9289);
or U9464 (N_9464,N_9368,N_9377);
xor U9465 (N_9465,N_9348,N_9239);
or U9466 (N_9466,N_9325,N_9346);
nand U9467 (N_9467,N_9303,N_9321);
and U9468 (N_9468,N_9333,N_9213);
xnor U9469 (N_9469,N_9357,N_9225);
and U9470 (N_9470,N_9291,N_9287);
and U9471 (N_9471,N_9352,N_9314);
xor U9472 (N_9472,N_9302,N_9288);
or U9473 (N_9473,N_9296,N_9387);
xor U9474 (N_9474,N_9379,N_9347);
nand U9475 (N_9475,N_9269,N_9309);
or U9476 (N_9476,N_9292,N_9254);
nand U9477 (N_9477,N_9399,N_9319);
and U9478 (N_9478,N_9217,N_9344);
nand U9479 (N_9479,N_9265,N_9316);
or U9480 (N_9480,N_9244,N_9335);
and U9481 (N_9481,N_9322,N_9257);
xnor U9482 (N_9482,N_9351,N_9294);
nand U9483 (N_9483,N_9384,N_9363);
and U9484 (N_9484,N_9332,N_9204);
and U9485 (N_9485,N_9249,N_9231);
xnor U9486 (N_9486,N_9393,N_9222);
xnor U9487 (N_9487,N_9345,N_9320);
and U9488 (N_9488,N_9227,N_9299);
or U9489 (N_9489,N_9246,N_9360);
and U9490 (N_9490,N_9386,N_9259);
or U9491 (N_9491,N_9264,N_9216);
and U9492 (N_9492,N_9318,N_9297);
and U9493 (N_9493,N_9253,N_9224);
xor U9494 (N_9494,N_9378,N_9380);
or U9495 (N_9495,N_9330,N_9266);
or U9496 (N_9496,N_9220,N_9218);
and U9497 (N_9497,N_9221,N_9203);
xor U9498 (N_9498,N_9334,N_9305);
and U9499 (N_9499,N_9366,N_9307);
nand U9500 (N_9500,N_9356,N_9370);
nand U9501 (N_9501,N_9361,N_9354);
xnor U9502 (N_9502,N_9344,N_9388);
nand U9503 (N_9503,N_9246,N_9206);
and U9504 (N_9504,N_9300,N_9200);
nand U9505 (N_9505,N_9381,N_9339);
nand U9506 (N_9506,N_9353,N_9331);
and U9507 (N_9507,N_9388,N_9261);
and U9508 (N_9508,N_9288,N_9283);
xnor U9509 (N_9509,N_9221,N_9392);
or U9510 (N_9510,N_9218,N_9374);
nand U9511 (N_9511,N_9234,N_9335);
xnor U9512 (N_9512,N_9355,N_9261);
xnor U9513 (N_9513,N_9286,N_9309);
or U9514 (N_9514,N_9294,N_9321);
xor U9515 (N_9515,N_9319,N_9359);
nand U9516 (N_9516,N_9285,N_9361);
nand U9517 (N_9517,N_9312,N_9307);
or U9518 (N_9518,N_9361,N_9215);
nand U9519 (N_9519,N_9390,N_9304);
and U9520 (N_9520,N_9288,N_9242);
and U9521 (N_9521,N_9212,N_9362);
or U9522 (N_9522,N_9377,N_9376);
nand U9523 (N_9523,N_9242,N_9235);
or U9524 (N_9524,N_9398,N_9230);
and U9525 (N_9525,N_9309,N_9302);
nor U9526 (N_9526,N_9230,N_9377);
or U9527 (N_9527,N_9390,N_9215);
or U9528 (N_9528,N_9386,N_9289);
and U9529 (N_9529,N_9247,N_9235);
nor U9530 (N_9530,N_9382,N_9218);
nand U9531 (N_9531,N_9360,N_9363);
or U9532 (N_9532,N_9376,N_9235);
nand U9533 (N_9533,N_9271,N_9399);
and U9534 (N_9534,N_9263,N_9269);
xnor U9535 (N_9535,N_9258,N_9201);
nand U9536 (N_9536,N_9381,N_9207);
xnor U9537 (N_9537,N_9394,N_9376);
xor U9538 (N_9538,N_9248,N_9269);
nor U9539 (N_9539,N_9203,N_9373);
nand U9540 (N_9540,N_9352,N_9287);
xor U9541 (N_9541,N_9236,N_9390);
nor U9542 (N_9542,N_9346,N_9240);
nor U9543 (N_9543,N_9398,N_9326);
xnor U9544 (N_9544,N_9251,N_9344);
or U9545 (N_9545,N_9295,N_9220);
nor U9546 (N_9546,N_9257,N_9360);
or U9547 (N_9547,N_9278,N_9368);
nand U9548 (N_9548,N_9236,N_9203);
xnor U9549 (N_9549,N_9317,N_9368);
and U9550 (N_9550,N_9295,N_9277);
nand U9551 (N_9551,N_9208,N_9331);
nand U9552 (N_9552,N_9369,N_9236);
xor U9553 (N_9553,N_9254,N_9388);
and U9554 (N_9554,N_9244,N_9311);
xor U9555 (N_9555,N_9399,N_9265);
and U9556 (N_9556,N_9372,N_9244);
and U9557 (N_9557,N_9201,N_9235);
and U9558 (N_9558,N_9346,N_9306);
nor U9559 (N_9559,N_9295,N_9268);
nor U9560 (N_9560,N_9322,N_9232);
nor U9561 (N_9561,N_9348,N_9251);
and U9562 (N_9562,N_9364,N_9273);
nand U9563 (N_9563,N_9271,N_9223);
or U9564 (N_9564,N_9297,N_9201);
nor U9565 (N_9565,N_9200,N_9270);
xnor U9566 (N_9566,N_9293,N_9282);
and U9567 (N_9567,N_9326,N_9399);
nor U9568 (N_9568,N_9293,N_9232);
xor U9569 (N_9569,N_9307,N_9348);
xor U9570 (N_9570,N_9276,N_9269);
nand U9571 (N_9571,N_9234,N_9398);
or U9572 (N_9572,N_9241,N_9210);
nor U9573 (N_9573,N_9250,N_9254);
or U9574 (N_9574,N_9395,N_9383);
nand U9575 (N_9575,N_9253,N_9275);
nand U9576 (N_9576,N_9342,N_9263);
nand U9577 (N_9577,N_9237,N_9393);
and U9578 (N_9578,N_9270,N_9214);
nand U9579 (N_9579,N_9327,N_9370);
xnor U9580 (N_9580,N_9316,N_9284);
nand U9581 (N_9581,N_9364,N_9230);
nor U9582 (N_9582,N_9295,N_9256);
nand U9583 (N_9583,N_9240,N_9268);
nor U9584 (N_9584,N_9337,N_9334);
or U9585 (N_9585,N_9351,N_9206);
and U9586 (N_9586,N_9267,N_9341);
or U9587 (N_9587,N_9214,N_9342);
xnor U9588 (N_9588,N_9319,N_9341);
or U9589 (N_9589,N_9284,N_9258);
or U9590 (N_9590,N_9241,N_9227);
and U9591 (N_9591,N_9214,N_9264);
and U9592 (N_9592,N_9320,N_9217);
xnor U9593 (N_9593,N_9299,N_9306);
or U9594 (N_9594,N_9359,N_9240);
xor U9595 (N_9595,N_9242,N_9290);
and U9596 (N_9596,N_9210,N_9229);
xnor U9597 (N_9597,N_9280,N_9229);
xnor U9598 (N_9598,N_9252,N_9324);
xnor U9599 (N_9599,N_9216,N_9368);
nor U9600 (N_9600,N_9514,N_9497);
and U9601 (N_9601,N_9532,N_9446);
nor U9602 (N_9602,N_9495,N_9537);
and U9603 (N_9603,N_9584,N_9513);
xnor U9604 (N_9604,N_9421,N_9587);
nor U9605 (N_9605,N_9466,N_9472);
xor U9606 (N_9606,N_9458,N_9541);
and U9607 (N_9607,N_9451,N_9536);
nand U9608 (N_9608,N_9496,N_9492);
nor U9609 (N_9609,N_9419,N_9564);
xnor U9610 (N_9610,N_9468,N_9475);
nand U9611 (N_9611,N_9510,N_9436);
or U9612 (N_9612,N_9459,N_9546);
xnor U9613 (N_9613,N_9527,N_9518);
xor U9614 (N_9614,N_9453,N_9521);
nor U9615 (N_9615,N_9545,N_9586);
and U9616 (N_9616,N_9413,N_9409);
nand U9617 (N_9617,N_9522,N_9529);
xnor U9618 (N_9618,N_9534,N_9483);
or U9619 (N_9619,N_9535,N_9410);
xnor U9620 (N_9620,N_9543,N_9552);
nand U9621 (N_9621,N_9523,N_9476);
nor U9622 (N_9622,N_9554,N_9542);
and U9623 (N_9623,N_9516,N_9550);
nand U9624 (N_9624,N_9406,N_9593);
nor U9625 (N_9625,N_9427,N_9405);
and U9626 (N_9626,N_9408,N_9504);
and U9627 (N_9627,N_9429,N_9414);
or U9628 (N_9628,N_9460,N_9478);
or U9629 (N_9629,N_9590,N_9547);
nor U9630 (N_9630,N_9508,N_9581);
nand U9631 (N_9631,N_9402,N_9438);
nand U9632 (N_9632,N_9525,N_9563);
nor U9633 (N_9633,N_9592,N_9577);
or U9634 (N_9634,N_9566,N_9580);
nand U9635 (N_9635,N_9403,N_9530);
nand U9636 (N_9636,N_9463,N_9488);
xor U9637 (N_9637,N_9442,N_9417);
or U9638 (N_9638,N_9567,N_9416);
and U9639 (N_9639,N_9556,N_9502);
nand U9640 (N_9640,N_9568,N_9557);
nand U9641 (N_9641,N_9576,N_9553);
xor U9642 (N_9642,N_9520,N_9501);
or U9643 (N_9643,N_9450,N_9594);
nand U9644 (N_9644,N_9435,N_9507);
and U9645 (N_9645,N_9500,N_9505);
nor U9646 (N_9646,N_9517,N_9511);
or U9647 (N_9647,N_9439,N_9582);
nor U9648 (N_9648,N_9578,N_9531);
and U9649 (N_9649,N_9441,N_9509);
nand U9650 (N_9650,N_9434,N_9599);
and U9651 (N_9651,N_9526,N_9482);
or U9652 (N_9652,N_9432,N_9498);
xnor U9653 (N_9653,N_9598,N_9457);
or U9654 (N_9654,N_9512,N_9415);
nor U9655 (N_9655,N_9469,N_9448);
xor U9656 (N_9656,N_9561,N_9503);
nand U9657 (N_9657,N_9575,N_9571);
xnor U9658 (N_9658,N_9430,N_9558);
nand U9659 (N_9659,N_9538,N_9589);
xnor U9660 (N_9660,N_9443,N_9452);
and U9661 (N_9661,N_9551,N_9562);
and U9662 (N_9662,N_9479,N_9515);
xor U9663 (N_9663,N_9440,N_9461);
or U9664 (N_9664,N_9454,N_9528);
nand U9665 (N_9665,N_9539,N_9572);
or U9666 (N_9666,N_9549,N_9473);
or U9667 (N_9667,N_9499,N_9588);
or U9668 (N_9668,N_9560,N_9591);
xor U9669 (N_9669,N_9596,N_9548);
or U9670 (N_9670,N_9565,N_9491);
and U9671 (N_9671,N_9484,N_9540);
xnor U9672 (N_9672,N_9490,N_9445);
xor U9673 (N_9673,N_9407,N_9555);
and U9674 (N_9674,N_9433,N_9506);
nor U9675 (N_9675,N_9533,N_9455);
nand U9676 (N_9676,N_9486,N_9422);
xor U9677 (N_9677,N_9467,N_9579);
or U9678 (N_9678,N_9494,N_9489);
or U9679 (N_9679,N_9493,N_9480);
and U9680 (N_9680,N_9519,N_9595);
xor U9681 (N_9681,N_9424,N_9428);
and U9682 (N_9682,N_9574,N_9559);
nor U9683 (N_9683,N_9400,N_9401);
xor U9684 (N_9684,N_9425,N_9583);
nand U9685 (N_9685,N_9449,N_9471);
xnor U9686 (N_9686,N_9456,N_9426);
nor U9687 (N_9687,N_9481,N_9544);
xnor U9688 (N_9688,N_9437,N_9420);
and U9689 (N_9689,N_9431,N_9570);
nor U9690 (N_9690,N_9423,N_9569);
nor U9691 (N_9691,N_9465,N_9418);
or U9692 (N_9692,N_9524,N_9585);
xnor U9693 (N_9693,N_9487,N_9573);
xnor U9694 (N_9694,N_9470,N_9464);
and U9695 (N_9695,N_9474,N_9444);
nand U9696 (N_9696,N_9411,N_9447);
nand U9697 (N_9697,N_9477,N_9597);
nand U9698 (N_9698,N_9404,N_9462);
xor U9699 (N_9699,N_9412,N_9485);
nor U9700 (N_9700,N_9586,N_9404);
xor U9701 (N_9701,N_9543,N_9422);
xor U9702 (N_9702,N_9518,N_9401);
xor U9703 (N_9703,N_9587,N_9560);
xnor U9704 (N_9704,N_9454,N_9585);
and U9705 (N_9705,N_9525,N_9522);
or U9706 (N_9706,N_9507,N_9414);
xor U9707 (N_9707,N_9414,N_9417);
xor U9708 (N_9708,N_9502,N_9418);
nand U9709 (N_9709,N_9572,N_9421);
xnor U9710 (N_9710,N_9586,N_9421);
and U9711 (N_9711,N_9547,N_9520);
xnor U9712 (N_9712,N_9518,N_9427);
nand U9713 (N_9713,N_9480,N_9591);
nand U9714 (N_9714,N_9460,N_9504);
and U9715 (N_9715,N_9521,N_9488);
or U9716 (N_9716,N_9516,N_9454);
xnor U9717 (N_9717,N_9414,N_9487);
and U9718 (N_9718,N_9441,N_9472);
or U9719 (N_9719,N_9449,N_9440);
and U9720 (N_9720,N_9487,N_9537);
xor U9721 (N_9721,N_9455,N_9441);
xnor U9722 (N_9722,N_9574,N_9567);
xnor U9723 (N_9723,N_9438,N_9578);
or U9724 (N_9724,N_9456,N_9471);
xor U9725 (N_9725,N_9445,N_9598);
or U9726 (N_9726,N_9405,N_9544);
nor U9727 (N_9727,N_9546,N_9470);
xnor U9728 (N_9728,N_9483,N_9517);
nand U9729 (N_9729,N_9444,N_9570);
and U9730 (N_9730,N_9583,N_9416);
and U9731 (N_9731,N_9497,N_9450);
and U9732 (N_9732,N_9514,N_9402);
xor U9733 (N_9733,N_9539,N_9492);
and U9734 (N_9734,N_9454,N_9554);
nand U9735 (N_9735,N_9405,N_9504);
nor U9736 (N_9736,N_9539,N_9429);
nor U9737 (N_9737,N_9571,N_9548);
nor U9738 (N_9738,N_9585,N_9459);
and U9739 (N_9739,N_9479,N_9425);
or U9740 (N_9740,N_9405,N_9534);
nor U9741 (N_9741,N_9482,N_9523);
and U9742 (N_9742,N_9524,N_9512);
nor U9743 (N_9743,N_9412,N_9416);
or U9744 (N_9744,N_9549,N_9410);
xor U9745 (N_9745,N_9476,N_9584);
nor U9746 (N_9746,N_9410,N_9402);
or U9747 (N_9747,N_9456,N_9530);
nand U9748 (N_9748,N_9468,N_9439);
and U9749 (N_9749,N_9490,N_9468);
and U9750 (N_9750,N_9419,N_9503);
nand U9751 (N_9751,N_9499,N_9439);
and U9752 (N_9752,N_9476,N_9597);
or U9753 (N_9753,N_9443,N_9595);
and U9754 (N_9754,N_9555,N_9473);
and U9755 (N_9755,N_9565,N_9496);
nor U9756 (N_9756,N_9532,N_9469);
nor U9757 (N_9757,N_9455,N_9504);
nand U9758 (N_9758,N_9522,N_9475);
and U9759 (N_9759,N_9460,N_9464);
or U9760 (N_9760,N_9534,N_9516);
and U9761 (N_9761,N_9599,N_9433);
nor U9762 (N_9762,N_9588,N_9491);
nor U9763 (N_9763,N_9437,N_9410);
and U9764 (N_9764,N_9410,N_9413);
and U9765 (N_9765,N_9555,N_9580);
xnor U9766 (N_9766,N_9486,N_9451);
xor U9767 (N_9767,N_9577,N_9517);
xnor U9768 (N_9768,N_9572,N_9439);
or U9769 (N_9769,N_9538,N_9586);
nor U9770 (N_9770,N_9534,N_9465);
nor U9771 (N_9771,N_9487,N_9434);
or U9772 (N_9772,N_9417,N_9436);
nand U9773 (N_9773,N_9550,N_9401);
or U9774 (N_9774,N_9494,N_9533);
nor U9775 (N_9775,N_9540,N_9448);
xor U9776 (N_9776,N_9433,N_9545);
nand U9777 (N_9777,N_9497,N_9481);
and U9778 (N_9778,N_9489,N_9406);
or U9779 (N_9779,N_9412,N_9411);
or U9780 (N_9780,N_9556,N_9447);
or U9781 (N_9781,N_9470,N_9456);
or U9782 (N_9782,N_9425,N_9587);
xor U9783 (N_9783,N_9445,N_9504);
or U9784 (N_9784,N_9457,N_9553);
and U9785 (N_9785,N_9416,N_9466);
xor U9786 (N_9786,N_9501,N_9554);
and U9787 (N_9787,N_9476,N_9508);
nor U9788 (N_9788,N_9586,N_9464);
nor U9789 (N_9789,N_9584,N_9535);
or U9790 (N_9790,N_9423,N_9434);
nand U9791 (N_9791,N_9408,N_9503);
nor U9792 (N_9792,N_9470,N_9574);
and U9793 (N_9793,N_9457,N_9472);
xor U9794 (N_9794,N_9408,N_9463);
xor U9795 (N_9795,N_9541,N_9529);
and U9796 (N_9796,N_9497,N_9456);
nand U9797 (N_9797,N_9440,N_9493);
nor U9798 (N_9798,N_9494,N_9577);
nor U9799 (N_9799,N_9429,N_9543);
nor U9800 (N_9800,N_9611,N_9693);
xnor U9801 (N_9801,N_9620,N_9633);
nor U9802 (N_9802,N_9789,N_9761);
xnor U9803 (N_9803,N_9667,N_9795);
nand U9804 (N_9804,N_9624,N_9665);
nor U9805 (N_9805,N_9733,N_9681);
xnor U9806 (N_9806,N_9653,N_9691);
or U9807 (N_9807,N_9771,N_9654);
nor U9808 (N_9808,N_9796,N_9704);
xor U9809 (N_9809,N_9661,N_9788);
and U9810 (N_9810,N_9712,N_9673);
xnor U9811 (N_9811,N_9675,N_9600);
nand U9812 (N_9812,N_9780,N_9669);
xor U9813 (N_9813,N_9629,N_9781);
and U9814 (N_9814,N_9778,N_9775);
nor U9815 (N_9815,N_9762,N_9641);
xnor U9816 (N_9816,N_9790,N_9660);
or U9817 (N_9817,N_9695,N_9649);
nand U9818 (N_9818,N_9770,N_9682);
nor U9819 (N_9819,N_9603,N_9715);
xnor U9820 (N_9820,N_9724,N_9602);
nand U9821 (N_9821,N_9688,N_9619);
nand U9822 (N_9822,N_9754,N_9765);
nand U9823 (N_9823,N_9701,N_9779);
or U9824 (N_9824,N_9747,N_9614);
nand U9825 (N_9825,N_9721,N_9692);
nand U9826 (N_9826,N_9755,N_9612);
nor U9827 (N_9827,N_9737,N_9774);
xor U9828 (N_9828,N_9657,N_9738);
nor U9829 (N_9829,N_9791,N_9750);
nand U9830 (N_9830,N_9698,N_9618);
or U9831 (N_9831,N_9767,N_9787);
nand U9832 (N_9832,N_9783,N_9658);
xor U9833 (N_9833,N_9708,N_9797);
nor U9834 (N_9834,N_9622,N_9792);
and U9835 (N_9835,N_9748,N_9739);
nor U9836 (N_9836,N_9639,N_9606);
nor U9837 (N_9837,N_9719,N_9656);
nor U9838 (N_9838,N_9760,N_9685);
and U9839 (N_9839,N_9670,N_9745);
nor U9840 (N_9840,N_9727,N_9728);
or U9841 (N_9841,N_9758,N_9768);
xor U9842 (N_9842,N_9621,N_9753);
and U9843 (N_9843,N_9652,N_9617);
xor U9844 (N_9844,N_9640,N_9794);
nor U9845 (N_9845,N_9610,N_9752);
nand U9846 (N_9846,N_9632,N_9638);
nand U9847 (N_9847,N_9607,N_9613);
xnor U9848 (N_9848,N_9766,N_9625);
and U9849 (N_9849,N_9683,N_9676);
or U9850 (N_9850,N_9720,N_9679);
xor U9851 (N_9851,N_9655,N_9694);
and U9852 (N_9852,N_9723,N_9671);
nand U9853 (N_9853,N_9687,N_9776);
nand U9854 (N_9854,N_9772,N_9740);
and U9855 (N_9855,N_9734,N_9623);
and U9856 (N_9856,N_9609,N_9648);
nand U9857 (N_9857,N_9746,N_9709);
nor U9858 (N_9858,N_9702,N_9799);
nand U9859 (N_9859,N_9730,N_9785);
xnor U9860 (N_9860,N_9798,N_9793);
nand U9861 (N_9861,N_9616,N_9697);
xnor U9862 (N_9862,N_9615,N_9651);
or U9863 (N_9863,N_9672,N_9725);
or U9864 (N_9864,N_9696,N_9645);
nor U9865 (N_9865,N_9668,N_9703);
nand U9866 (N_9866,N_9732,N_9647);
xor U9867 (N_9867,N_9642,N_9786);
and U9868 (N_9868,N_9678,N_9690);
nor U9869 (N_9869,N_9666,N_9605);
xor U9870 (N_9870,N_9628,N_9711);
nand U9871 (N_9871,N_9777,N_9643);
and U9872 (N_9872,N_9663,N_9636);
xnor U9873 (N_9873,N_9736,N_9700);
nand U9874 (N_9874,N_9751,N_9637);
nand U9875 (N_9875,N_9634,N_9631);
or U9876 (N_9876,N_9757,N_9644);
and U9877 (N_9877,N_9744,N_9749);
and U9878 (N_9878,N_9646,N_9717);
xnor U9879 (N_9879,N_9769,N_9743);
xor U9880 (N_9880,N_9664,N_9773);
nand U9881 (N_9881,N_9650,N_9706);
and U9882 (N_9882,N_9630,N_9726);
nor U9883 (N_9883,N_9782,N_9684);
nor U9884 (N_9884,N_9713,N_9699);
nor U9885 (N_9885,N_9718,N_9722);
nor U9886 (N_9886,N_9604,N_9601);
and U9887 (N_9887,N_9674,N_9735);
nor U9888 (N_9888,N_9705,N_9756);
nor U9889 (N_9889,N_9784,N_9759);
and U9890 (N_9890,N_9710,N_9763);
nor U9891 (N_9891,N_9742,N_9716);
or U9892 (N_9892,N_9714,N_9707);
and U9893 (N_9893,N_9731,N_9608);
nand U9894 (N_9894,N_9729,N_9635);
or U9895 (N_9895,N_9680,N_9689);
xor U9896 (N_9896,N_9659,N_9741);
nand U9897 (N_9897,N_9677,N_9626);
or U9898 (N_9898,N_9662,N_9686);
nand U9899 (N_9899,N_9764,N_9627);
or U9900 (N_9900,N_9723,N_9779);
or U9901 (N_9901,N_9743,N_9600);
xor U9902 (N_9902,N_9758,N_9660);
nor U9903 (N_9903,N_9712,N_9664);
and U9904 (N_9904,N_9655,N_9715);
nor U9905 (N_9905,N_9762,N_9732);
xor U9906 (N_9906,N_9692,N_9710);
or U9907 (N_9907,N_9789,N_9757);
nor U9908 (N_9908,N_9738,N_9689);
and U9909 (N_9909,N_9681,N_9707);
and U9910 (N_9910,N_9767,N_9607);
nand U9911 (N_9911,N_9722,N_9796);
or U9912 (N_9912,N_9694,N_9631);
nor U9913 (N_9913,N_9719,N_9619);
nand U9914 (N_9914,N_9720,N_9600);
and U9915 (N_9915,N_9638,N_9748);
nor U9916 (N_9916,N_9786,N_9659);
xor U9917 (N_9917,N_9637,N_9755);
nand U9918 (N_9918,N_9708,N_9645);
nand U9919 (N_9919,N_9602,N_9650);
or U9920 (N_9920,N_9667,N_9750);
and U9921 (N_9921,N_9698,N_9711);
nand U9922 (N_9922,N_9644,N_9641);
xnor U9923 (N_9923,N_9649,N_9625);
or U9924 (N_9924,N_9625,N_9709);
nand U9925 (N_9925,N_9618,N_9784);
nand U9926 (N_9926,N_9790,N_9719);
or U9927 (N_9927,N_9631,N_9644);
nor U9928 (N_9928,N_9686,N_9671);
xnor U9929 (N_9929,N_9798,N_9676);
nand U9930 (N_9930,N_9659,N_9699);
nand U9931 (N_9931,N_9780,N_9703);
or U9932 (N_9932,N_9619,N_9620);
nand U9933 (N_9933,N_9635,N_9770);
xnor U9934 (N_9934,N_9719,N_9720);
nand U9935 (N_9935,N_9765,N_9625);
and U9936 (N_9936,N_9731,N_9775);
xor U9937 (N_9937,N_9615,N_9728);
and U9938 (N_9938,N_9691,N_9796);
nor U9939 (N_9939,N_9637,N_9649);
nand U9940 (N_9940,N_9703,N_9798);
nor U9941 (N_9941,N_9693,N_9702);
and U9942 (N_9942,N_9756,N_9736);
xor U9943 (N_9943,N_9656,N_9756);
nor U9944 (N_9944,N_9613,N_9756);
nand U9945 (N_9945,N_9717,N_9760);
and U9946 (N_9946,N_9603,N_9622);
nand U9947 (N_9947,N_9613,N_9710);
nand U9948 (N_9948,N_9685,N_9714);
and U9949 (N_9949,N_9734,N_9742);
nand U9950 (N_9950,N_9668,N_9610);
xnor U9951 (N_9951,N_9639,N_9776);
xor U9952 (N_9952,N_9705,N_9788);
and U9953 (N_9953,N_9670,N_9668);
nand U9954 (N_9954,N_9676,N_9705);
and U9955 (N_9955,N_9797,N_9785);
nand U9956 (N_9956,N_9603,N_9655);
nor U9957 (N_9957,N_9707,N_9736);
or U9958 (N_9958,N_9679,N_9770);
nand U9959 (N_9959,N_9671,N_9600);
nor U9960 (N_9960,N_9654,N_9715);
xor U9961 (N_9961,N_9608,N_9654);
nand U9962 (N_9962,N_9609,N_9688);
nor U9963 (N_9963,N_9658,N_9747);
nor U9964 (N_9964,N_9672,N_9784);
and U9965 (N_9965,N_9623,N_9714);
or U9966 (N_9966,N_9783,N_9751);
xnor U9967 (N_9967,N_9769,N_9781);
xor U9968 (N_9968,N_9689,N_9784);
xnor U9969 (N_9969,N_9798,N_9704);
xor U9970 (N_9970,N_9696,N_9735);
and U9971 (N_9971,N_9701,N_9725);
nor U9972 (N_9972,N_9714,N_9671);
or U9973 (N_9973,N_9720,N_9773);
or U9974 (N_9974,N_9720,N_9648);
and U9975 (N_9975,N_9711,N_9638);
and U9976 (N_9976,N_9658,N_9785);
and U9977 (N_9977,N_9709,N_9733);
and U9978 (N_9978,N_9728,N_9788);
or U9979 (N_9979,N_9643,N_9698);
or U9980 (N_9980,N_9632,N_9716);
or U9981 (N_9981,N_9604,N_9602);
nor U9982 (N_9982,N_9740,N_9762);
or U9983 (N_9983,N_9647,N_9655);
nor U9984 (N_9984,N_9770,N_9656);
or U9985 (N_9985,N_9751,N_9761);
nor U9986 (N_9986,N_9798,N_9692);
xnor U9987 (N_9987,N_9641,N_9700);
and U9988 (N_9988,N_9733,N_9700);
xor U9989 (N_9989,N_9689,N_9667);
nor U9990 (N_9990,N_9725,N_9616);
xor U9991 (N_9991,N_9777,N_9653);
nand U9992 (N_9992,N_9735,N_9719);
xnor U9993 (N_9993,N_9653,N_9696);
nor U9994 (N_9994,N_9678,N_9735);
nand U9995 (N_9995,N_9793,N_9766);
nor U9996 (N_9996,N_9775,N_9696);
xnor U9997 (N_9997,N_9628,N_9660);
nor U9998 (N_9998,N_9778,N_9647);
xnor U9999 (N_9999,N_9778,N_9704);
xor U10000 (N_10000,N_9873,N_9884);
or U10001 (N_10001,N_9963,N_9813);
xor U10002 (N_10002,N_9985,N_9941);
or U10003 (N_10003,N_9881,N_9959);
and U10004 (N_10004,N_9912,N_9871);
xor U10005 (N_10005,N_9885,N_9933);
nor U10006 (N_10006,N_9811,N_9927);
nor U10007 (N_10007,N_9895,N_9865);
nand U10008 (N_10008,N_9856,N_9888);
nand U10009 (N_10009,N_9940,N_9847);
or U10010 (N_10010,N_9970,N_9991);
xnor U10011 (N_10011,N_9817,N_9801);
nor U10012 (N_10012,N_9841,N_9976);
nand U10013 (N_10013,N_9859,N_9823);
and U10014 (N_10014,N_9978,N_9848);
nor U10015 (N_10015,N_9879,N_9947);
and U10016 (N_10016,N_9827,N_9808);
and U10017 (N_10017,N_9863,N_9950);
and U10018 (N_10018,N_9953,N_9938);
nor U10019 (N_10019,N_9812,N_9907);
nor U10020 (N_10020,N_9875,N_9843);
or U10021 (N_10021,N_9922,N_9832);
xnor U10022 (N_10022,N_9909,N_9842);
xnor U10023 (N_10023,N_9867,N_9937);
or U10024 (N_10024,N_9840,N_9904);
xnor U10025 (N_10025,N_9844,N_9929);
and U10026 (N_10026,N_9956,N_9911);
xnor U10027 (N_10027,N_9890,N_9854);
nand U10028 (N_10028,N_9852,N_9830);
xnor U10029 (N_10029,N_9908,N_9820);
xor U10030 (N_10030,N_9818,N_9977);
and U10031 (N_10031,N_9825,N_9946);
or U10032 (N_10032,N_9892,N_9920);
or U10033 (N_10033,N_9913,N_9862);
nand U10034 (N_10034,N_9997,N_9928);
or U10035 (N_10035,N_9806,N_9942);
and U10036 (N_10036,N_9845,N_9821);
nand U10037 (N_10037,N_9987,N_9943);
and U10038 (N_10038,N_9849,N_9853);
nand U10039 (N_10039,N_9864,N_9855);
and U10040 (N_10040,N_9926,N_9874);
and U10041 (N_10041,N_9998,N_9819);
xor U10042 (N_10042,N_9981,N_9898);
or U10043 (N_10043,N_9896,N_9994);
or U10044 (N_10044,N_9836,N_9983);
nand U10045 (N_10045,N_9966,N_9804);
nand U10046 (N_10046,N_9858,N_9949);
xnor U10047 (N_10047,N_9971,N_9932);
nand U10048 (N_10048,N_9995,N_9986);
nand U10049 (N_10049,N_9916,N_9989);
nor U10050 (N_10050,N_9883,N_9968);
xor U10051 (N_10051,N_9846,N_9893);
xor U10052 (N_10052,N_9973,N_9872);
nand U10053 (N_10053,N_9954,N_9945);
and U10054 (N_10054,N_9918,N_9955);
and U10055 (N_10055,N_9860,N_9861);
xor U10056 (N_10056,N_9988,N_9967);
or U10057 (N_10057,N_9925,N_9882);
nand U10058 (N_10058,N_9894,N_9900);
nand U10059 (N_10059,N_9980,N_9915);
or U10060 (N_10060,N_9815,N_9880);
nand U10061 (N_10061,N_9901,N_9805);
and U10062 (N_10062,N_9886,N_9951);
and U10063 (N_10063,N_9826,N_9851);
xor U10064 (N_10064,N_9944,N_9975);
xnor U10065 (N_10065,N_9887,N_9877);
and U10066 (N_10066,N_9889,N_9837);
nand U10067 (N_10067,N_9906,N_9809);
or U10068 (N_10068,N_9868,N_9960);
or U10069 (N_10069,N_9993,N_9914);
nor U10070 (N_10070,N_9838,N_9921);
xnor U10071 (N_10071,N_9919,N_9828);
and U10072 (N_10072,N_9972,N_9939);
nor U10073 (N_10073,N_9984,N_9807);
nand U10074 (N_10074,N_9869,N_9810);
xor U10075 (N_10075,N_9948,N_9850);
and U10076 (N_10076,N_9996,N_9917);
and U10077 (N_10077,N_9800,N_9816);
nand U10078 (N_10078,N_9905,N_9924);
nor U10079 (N_10079,N_9990,N_9934);
nor U10080 (N_10080,N_9910,N_9876);
xnor U10081 (N_10081,N_9974,N_9962);
and U10082 (N_10082,N_9935,N_9964);
xor U10083 (N_10083,N_9839,N_9979);
nor U10084 (N_10084,N_9958,N_9822);
nand U10085 (N_10085,N_9961,N_9814);
and U10086 (N_10086,N_9802,N_9969);
nor U10087 (N_10087,N_9891,N_9923);
nor U10088 (N_10088,N_9957,N_9899);
nor U10089 (N_10089,N_9897,N_9834);
nor U10090 (N_10090,N_9878,N_9902);
xnor U10091 (N_10091,N_9992,N_9982);
nor U10092 (N_10092,N_9965,N_9824);
nor U10093 (N_10093,N_9831,N_9870);
xnor U10094 (N_10094,N_9803,N_9829);
nor U10095 (N_10095,N_9857,N_9903);
and U10096 (N_10096,N_9930,N_9936);
xor U10097 (N_10097,N_9866,N_9835);
and U10098 (N_10098,N_9952,N_9931);
nand U10099 (N_10099,N_9833,N_9999);
or U10100 (N_10100,N_9971,N_9819);
nor U10101 (N_10101,N_9865,N_9946);
and U10102 (N_10102,N_9958,N_9832);
or U10103 (N_10103,N_9846,N_9931);
or U10104 (N_10104,N_9902,N_9871);
or U10105 (N_10105,N_9988,N_9937);
nand U10106 (N_10106,N_9967,N_9827);
nor U10107 (N_10107,N_9985,N_9944);
nand U10108 (N_10108,N_9991,N_9911);
nor U10109 (N_10109,N_9947,N_9963);
or U10110 (N_10110,N_9989,N_9867);
or U10111 (N_10111,N_9803,N_9918);
and U10112 (N_10112,N_9893,N_9946);
nor U10113 (N_10113,N_9863,N_9977);
nor U10114 (N_10114,N_9930,N_9887);
and U10115 (N_10115,N_9980,N_9937);
nor U10116 (N_10116,N_9842,N_9988);
or U10117 (N_10117,N_9855,N_9905);
nor U10118 (N_10118,N_9841,N_9835);
nand U10119 (N_10119,N_9975,N_9832);
nand U10120 (N_10120,N_9905,N_9927);
nand U10121 (N_10121,N_9847,N_9926);
and U10122 (N_10122,N_9947,N_9964);
or U10123 (N_10123,N_9969,N_9908);
xnor U10124 (N_10124,N_9873,N_9963);
nand U10125 (N_10125,N_9859,N_9993);
xnor U10126 (N_10126,N_9890,N_9985);
nand U10127 (N_10127,N_9929,N_9860);
xnor U10128 (N_10128,N_9928,N_9853);
nand U10129 (N_10129,N_9858,N_9893);
xor U10130 (N_10130,N_9906,N_9982);
and U10131 (N_10131,N_9977,N_9939);
xor U10132 (N_10132,N_9853,N_9837);
nand U10133 (N_10133,N_9849,N_9937);
or U10134 (N_10134,N_9923,N_9831);
or U10135 (N_10135,N_9986,N_9866);
xor U10136 (N_10136,N_9804,N_9943);
nor U10137 (N_10137,N_9888,N_9883);
or U10138 (N_10138,N_9897,N_9810);
nor U10139 (N_10139,N_9935,N_9838);
or U10140 (N_10140,N_9930,N_9830);
nor U10141 (N_10141,N_9906,N_9933);
and U10142 (N_10142,N_9810,N_9808);
nor U10143 (N_10143,N_9809,N_9863);
nand U10144 (N_10144,N_9884,N_9876);
xnor U10145 (N_10145,N_9855,N_9807);
nor U10146 (N_10146,N_9935,N_9931);
xor U10147 (N_10147,N_9890,N_9915);
or U10148 (N_10148,N_9933,N_9952);
or U10149 (N_10149,N_9828,N_9929);
and U10150 (N_10150,N_9982,N_9926);
and U10151 (N_10151,N_9858,N_9911);
nor U10152 (N_10152,N_9922,N_9877);
nand U10153 (N_10153,N_9973,N_9857);
nor U10154 (N_10154,N_9982,N_9937);
or U10155 (N_10155,N_9876,N_9900);
and U10156 (N_10156,N_9852,N_9935);
xnor U10157 (N_10157,N_9823,N_9829);
and U10158 (N_10158,N_9883,N_9941);
or U10159 (N_10159,N_9914,N_9881);
and U10160 (N_10160,N_9826,N_9923);
or U10161 (N_10161,N_9982,N_9999);
xor U10162 (N_10162,N_9938,N_9970);
and U10163 (N_10163,N_9820,N_9864);
xor U10164 (N_10164,N_9900,N_9873);
nand U10165 (N_10165,N_9893,N_9807);
or U10166 (N_10166,N_9934,N_9860);
nor U10167 (N_10167,N_9801,N_9936);
and U10168 (N_10168,N_9843,N_9932);
or U10169 (N_10169,N_9879,N_9970);
xnor U10170 (N_10170,N_9894,N_9902);
or U10171 (N_10171,N_9963,N_9832);
or U10172 (N_10172,N_9802,N_9952);
or U10173 (N_10173,N_9960,N_9800);
nor U10174 (N_10174,N_9823,N_9875);
xnor U10175 (N_10175,N_9854,N_9801);
xor U10176 (N_10176,N_9938,N_9897);
nand U10177 (N_10177,N_9850,N_9876);
xor U10178 (N_10178,N_9945,N_9933);
nor U10179 (N_10179,N_9981,N_9803);
or U10180 (N_10180,N_9848,N_9898);
nand U10181 (N_10181,N_9943,N_9947);
nand U10182 (N_10182,N_9853,N_9896);
nand U10183 (N_10183,N_9804,N_9973);
xnor U10184 (N_10184,N_9914,N_9938);
or U10185 (N_10185,N_9826,N_9989);
nor U10186 (N_10186,N_9858,N_9894);
nor U10187 (N_10187,N_9849,N_9884);
nand U10188 (N_10188,N_9825,N_9820);
and U10189 (N_10189,N_9960,N_9876);
nor U10190 (N_10190,N_9818,N_9884);
and U10191 (N_10191,N_9942,N_9955);
xor U10192 (N_10192,N_9981,N_9805);
nor U10193 (N_10193,N_9825,N_9894);
and U10194 (N_10194,N_9876,N_9807);
and U10195 (N_10195,N_9950,N_9830);
or U10196 (N_10196,N_9843,N_9854);
nor U10197 (N_10197,N_9803,N_9844);
xnor U10198 (N_10198,N_9987,N_9875);
nand U10199 (N_10199,N_9948,N_9899);
and U10200 (N_10200,N_10179,N_10109);
nor U10201 (N_10201,N_10131,N_10191);
or U10202 (N_10202,N_10065,N_10124);
nand U10203 (N_10203,N_10115,N_10013);
and U10204 (N_10204,N_10097,N_10139);
and U10205 (N_10205,N_10038,N_10057);
or U10206 (N_10206,N_10130,N_10072);
nor U10207 (N_10207,N_10173,N_10146);
or U10208 (N_10208,N_10091,N_10033);
or U10209 (N_10209,N_10068,N_10189);
or U10210 (N_10210,N_10081,N_10090);
or U10211 (N_10211,N_10073,N_10105);
and U10212 (N_10212,N_10087,N_10076);
nor U10213 (N_10213,N_10023,N_10002);
and U10214 (N_10214,N_10066,N_10182);
xnor U10215 (N_10215,N_10082,N_10040);
xor U10216 (N_10216,N_10166,N_10197);
or U10217 (N_10217,N_10047,N_10133);
nand U10218 (N_10218,N_10177,N_10148);
nand U10219 (N_10219,N_10074,N_10093);
nor U10220 (N_10220,N_10046,N_10102);
nor U10221 (N_10221,N_10089,N_10014);
nor U10222 (N_10222,N_10107,N_10017);
nor U10223 (N_10223,N_10001,N_10125);
nor U10224 (N_10224,N_10088,N_10027);
and U10225 (N_10225,N_10180,N_10052);
or U10226 (N_10226,N_10000,N_10170);
and U10227 (N_10227,N_10106,N_10080);
and U10228 (N_10228,N_10021,N_10015);
and U10229 (N_10229,N_10144,N_10003);
and U10230 (N_10230,N_10113,N_10056);
or U10231 (N_10231,N_10099,N_10188);
and U10232 (N_10232,N_10025,N_10181);
or U10233 (N_10233,N_10028,N_10049);
or U10234 (N_10234,N_10054,N_10140);
and U10235 (N_10235,N_10159,N_10194);
nor U10236 (N_10236,N_10085,N_10070);
nand U10237 (N_10237,N_10064,N_10006);
nor U10238 (N_10238,N_10005,N_10042);
xnor U10239 (N_10239,N_10167,N_10030);
nand U10240 (N_10240,N_10032,N_10075);
xor U10241 (N_10241,N_10160,N_10020);
nor U10242 (N_10242,N_10171,N_10035);
and U10243 (N_10243,N_10154,N_10163);
xnor U10244 (N_10244,N_10059,N_10175);
nor U10245 (N_10245,N_10127,N_10184);
xor U10246 (N_10246,N_10039,N_10037);
nand U10247 (N_10247,N_10147,N_10010);
xor U10248 (N_10248,N_10165,N_10162);
or U10249 (N_10249,N_10196,N_10024);
or U10250 (N_10250,N_10004,N_10026);
nand U10251 (N_10251,N_10185,N_10044);
nand U10252 (N_10252,N_10137,N_10009);
or U10253 (N_10253,N_10112,N_10132);
or U10254 (N_10254,N_10161,N_10022);
or U10255 (N_10255,N_10155,N_10098);
nor U10256 (N_10256,N_10018,N_10060);
and U10257 (N_10257,N_10193,N_10101);
nor U10258 (N_10258,N_10183,N_10078);
or U10259 (N_10259,N_10100,N_10008);
and U10260 (N_10260,N_10058,N_10069);
and U10261 (N_10261,N_10152,N_10153);
nand U10262 (N_10262,N_10063,N_10158);
or U10263 (N_10263,N_10129,N_10134);
and U10264 (N_10264,N_10036,N_10117);
nand U10265 (N_10265,N_10053,N_10168);
xnor U10266 (N_10266,N_10103,N_10051);
nor U10267 (N_10267,N_10141,N_10094);
nand U10268 (N_10268,N_10016,N_10142);
and U10269 (N_10269,N_10150,N_10172);
nand U10270 (N_10270,N_10195,N_10029);
nand U10271 (N_10271,N_10138,N_10045);
or U10272 (N_10272,N_10048,N_10192);
nand U10273 (N_10273,N_10186,N_10178);
and U10274 (N_10274,N_10041,N_10120);
or U10275 (N_10275,N_10114,N_10164);
nand U10276 (N_10276,N_10176,N_10067);
nor U10277 (N_10277,N_10104,N_10126);
xnor U10278 (N_10278,N_10092,N_10111);
or U10279 (N_10279,N_10121,N_10157);
and U10280 (N_10280,N_10116,N_10190);
or U10281 (N_10281,N_10135,N_10062);
xor U10282 (N_10282,N_10055,N_10031);
xnor U10283 (N_10283,N_10083,N_10012);
nand U10284 (N_10284,N_10187,N_10169);
nand U10285 (N_10285,N_10086,N_10145);
nor U10286 (N_10286,N_10050,N_10119);
nor U10287 (N_10287,N_10071,N_10019);
nor U10288 (N_10288,N_10151,N_10136);
nor U10289 (N_10289,N_10095,N_10128);
nor U10290 (N_10290,N_10079,N_10122);
or U10291 (N_10291,N_10156,N_10110);
or U10292 (N_10292,N_10007,N_10061);
nor U10293 (N_10293,N_10143,N_10108);
nand U10294 (N_10294,N_10118,N_10011);
nand U10295 (N_10295,N_10199,N_10174);
nand U10296 (N_10296,N_10123,N_10034);
nor U10297 (N_10297,N_10198,N_10084);
or U10298 (N_10298,N_10043,N_10149);
nand U10299 (N_10299,N_10096,N_10077);
nand U10300 (N_10300,N_10188,N_10137);
nor U10301 (N_10301,N_10155,N_10190);
or U10302 (N_10302,N_10187,N_10168);
and U10303 (N_10303,N_10147,N_10016);
and U10304 (N_10304,N_10043,N_10094);
and U10305 (N_10305,N_10040,N_10123);
or U10306 (N_10306,N_10080,N_10014);
and U10307 (N_10307,N_10053,N_10108);
nor U10308 (N_10308,N_10036,N_10123);
xnor U10309 (N_10309,N_10094,N_10191);
and U10310 (N_10310,N_10124,N_10120);
or U10311 (N_10311,N_10019,N_10135);
xor U10312 (N_10312,N_10069,N_10098);
nand U10313 (N_10313,N_10032,N_10185);
or U10314 (N_10314,N_10052,N_10063);
nor U10315 (N_10315,N_10076,N_10180);
nand U10316 (N_10316,N_10025,N_10119);
and U10317 (N_10317,N_10199,N_10197);
nand U10318 (N_10318,N_10081,N_10179);
xnor U10319 (N_10319,N_10136,N_10161);
and U10320 (N_10320,N_10137,N_10049);
nand U10321 (N_10321,N_10192,N_10060);
xor U10322 (N_10322,N_10072,N_10088);
nor U10323 (N_10323,N_10129,N_10088);
nor U10324 (N_10324,N_10188,N_10128);
nand U10325 (N_10325,N_10157,N_10194);
xnor U10326 (N_10326,N_10034,N_10134);
or U10327 (N_10327,N_10061,N_10177);
or U10328 (N_10328,N_10024,N_10007);
nor U10329 (N_10329,N_10137,N_10122);
nor U10330 (N_10330,N_10196,N_10117);
xnor U10331 (N_10331,N_10060,N_10039);
and U10332 (N_10332,N_10198,N_10011);
or U10333 (N_10333,N_10007,N_10012);
and U10334 (N_10334,N_10011,N_10109);
xnor U10335 (N_10335,N_10125,N_10184);
nand U10336 (N_10336,N_10003,N_10057);
nor U10337 (N_10337,N_10105,N_10127);
xnor U10338 (N_10338,N_10149,N_10097);
or U10339 (N_10339,N_10002,N_10125);
xor U10340 (N_10340,N_10152,N_10055);
xor U10341 (N_10341,N_10020,N_10078);
or U10342 (N_10342,N_10124,N_10088);
nand U10343 (N_10343,N_10018,N_10011);
xor U10344 (N_10344,N_10000,N_10082);
nand U10345 (N_10345,N_10071,N_10069);
nor U10346 (N_10346,N_10091,N_10095);
and U10347 (N_10347,N_10061,N_10126);
nor U10348 (N_10348,N_10089,N_10044);
nor U10349 (N_10349,N_10180,N_10027);
nand U10350 (N_10350,N_10050,N_10137);
nand U10351 (N_10351,N_10151,N_10113);
and U10352 (N_10352,N_10143,N_10024);
or U10353 (N_10353,N_10074,N_10162);
and U10354 (N_10354,N_10061,N_10164);
nor U10355 (N_10355,N_10068,N_10197);
nor U10356 (N_10356,N_10040,N_10017);
nand U10357 (N_10357,N_10017,N_10071);
nand U10358 (N_10358,N_10097,N_10047);
nand U10359 (N_10359,N_10117,N_10002);
or U10360 (N_10360,N_10009,N_10025);
nor U10361 (N_10361,N_10038,N_10042);
xor U10362 (N_10362,N_10048,N_10046);
nor U10363 (N_10363,N_10109,N_10149);
and U10364 (N_10364,N_10028,N_10196);
nand U10365 (N_10365,N_10007,N_10086);
nor U10366 (N_10366,N_10116,N_10170);
nand U10367 (N_10367,N_10123,N_10060);
nor U10368 (N_10368,N_10146,N_10182);
or U10369 (N_10369,N_10075,N_10002);
xnor U10370 (N_10370,N_10164,N_10172);
nand U10371 (N_10371,N_10109,N_10020);
nand U10372 (N_10372,N_10167,N_10177);
xor U10373 (N_10373,N_10039,N_10083);
and U10374 (N_10374,N_10191,N_10129);
nor U10375 (N_10375,N_10070,N_10009);
or U10376 (N_10376,N_10135,N_10162);
xnor U10377 (N_10377,N_10049,N_10005);
and U10378 (N_10378,N_10122,N_10061);
or U10379 (N_10379,N_10088,N_10162);
and U10380 (N_10380,N_10189,N_10031);
or U10381 (N_10381,N_10064,N_10039);
xor U10382 (N_10382,N_10029,N_10186);
nand U10383 (N_10383,N_10152,N_10008);
nand U10384 (N_10384,N_10032,N_10033);
and U10385 (N_10385,N_10149,N_10026);
and U10386 (N_10386,N_10096,N_10149);
or U10387 (N_10387,N_10092,N_10113);
nand U10388 (N_10388,N_10027,N_10074);
or U10389 (N_10389,N_10090,N_10070);
nand U10390 (N_10390,N_10167,N_10193);
and U10391 (N_10391,N_10156,N_10168);
and U10392 (N_10392,N_10148,N_10029);
nand U10393 (N_10393,N_10051,N_10090);
nor U10394 (N_10394,N_10174,N_10038);
xnor U10395 (N_10395,N_10127,N_10057);
or U10396 (N_10396,N_10017,N_10136);
xnor U10397 (N_10397,N_10074,N_10160);
and U10398 (N_10398,N_10161,N_10050);
or U10399 (N_10399,N_10094,N_10099);
nor U10400 (N_10400,N_10247,N_10265);
xor U10401 (N_10401,N_10366,N_10271);
nor U10402 (N_10402,N_10278,N_10315);
and U10403 (N_10403,N_10225,N_10252);
or U10404 (N_10404,N_10258,N_10202);
and U10405 (N_10405,N_10390,N_10340);
or U10406 (N_10406,N_10242,N_10356);
and U10407 (N_10407,N_10240,N_10373);
xnor U10408 (N_10408,N_10358,N_10273);
nor U10409 (N_10409,N_10362,N_10305);
xor U10410 (N_10410,N_10359,N_10336);
nor U10411 (N_10411,N_10322,N_10386);
nand U10412 (N_10412,N_10320,N_10351);
nand U10413 (N_10413,N_10397,N_10222);
and U10414 (N_10414,N_10367,N_10343);
and U10415 (N_10415,N_10277,N_10269);
nand U10416 (N_10416,N_10328,N_10243);
nand U10417 (N_10417,N_10207,N_10210);
nor U10418 (N_10418,N_10334,N_10368);
xnor U10419 (N_10419,N_10246,N_10348);
nand U10420 (N_10420,N_10209,N_10268);
or U10421 (N_10421,N_10369,N_10206);
and U10422 (N_10422,N_10357,N_10245);
xor U10423 (N_10423,N_10266,N_10347);
nor U10424 (N_10424,N_10241,N_10352);
nor U10425 (N_10425,N_10337,N_10306);
nand U10426 (N_10426,N_10272,N_10211);
nor U10427 (N_10427,N_10218,N_10360);
nor U10428 (N_10428,N_10301,N_10319);
nor U10429 (N_10429,N_10385,N_10262);
nand U10430 (N_10430,N_10297,N_10208);
nand U10431 (N_10431,N_10214,N_10376);
nor U10432 (N_10432,N_10370,N_10381);
nor U10433 (N_10433,N_10307,N_10205);
xnor U10434 (N_10434,N_10394,N_10313);
nor U10435 (N_10435,N_10310,N_10399);
nand U10436 (N_10436,N_10287,N_10204);
and U10437 (N_10437,N_10325,N_10285);
nor U10438 (N_10438,N_10329,N_10232);
nor U10439 (N_10439,N_10361,N_10349);
and U10440 (N_10440,N_10372,N_10239);
nor U10441 (N_10441,N_10217,N_10371);
nor U10442 (N_10442,N_10282,N_10229);
xor U10443 (N_10443,N_10261,N_10223);
or U10444 (N_10444,N_10383,N_10309);
and U10445 (N_10445,N_10286,N_10248);
or U10446 (N_10446,N_10304,N_10317);
nand U10447 (N_10447,N_10299,N_10374);
xnor U10448 (N_10448,N_10203,N_10251);
or U10449 (N_10449,N_10396,N_10395);
nor U10450 (N_10450,N_10255,N_10378);
nor U10451 (N_10451,N_10249,N_10288);
and U10452 (N_10452,N_10302,N_10219);
and U10453 (N_10453,N_10312,N_10380);
nor U10454 (N_10454,N_10384,N_10281);
or U10455 (N_10455,N_10321,N_10338);
or U10456 (N_10456,N_10226,N_10250);
nor U10457 (N_10457,N_10231,N_10355);
nand U10458 (N_10458,N_10339,N_10311);
nand U10459 (N_10459,N_10379,N_10392);
xnor U10460 (N_10460,N_10341,N_10254);
nor U10461 (N_10461,N_10332,N_10220);
nand U10462 (N_10462,N_10323,N_10387);
and U10463 (N_10463,N_10257,N_10212);
and U10464 (N_10464,N_10267,N_10353);
xor U10465 (N_10465,N_10303,N_10363);
or U10466 (N_10466,N_10234,N_10295);
or U10467 (N_10467,N_10233,N_10327);
xnor U10468 (N_10468,N_10256,N_10235);
or U10469 (N_10469,N_10293,N_10308);
xnor U10470 (N_10470,N_10342,N_10290);
and U10471 (N_10471,N_10259,N_10253);
or U10472 (N_10472,N_10296,N_10200);
nor U10473 (N_10473,N_10314,N_10330);
and U10474 (N_10474,N_10201,N_10375);
nand U10475 (N_10475,N_10275,N_10298);
nand U10476 (N_10476,N_10393,N_10228);
nand U10477 (N_10477,N_10215,N_10280);
or U10478 (N_10478,N_10238,N_10264);
or U10479 (N_10479,N_10354,N_10279);
nor U10480 (N_10480,N_10260,N_10388);
nand U10481 (N_10481,N_10289,N_10291);
and U10482 (N_10482,N_10318,N_10365);
nor U10483 (N_10483,N_10263,N_10230);
nand U10484 (N_10484,N_10294,N_10224);
or U10485 (N_10485,N_10389,N_10364);
or U10486 (N_10486,N_10244,N_10213);
or U10487 (N_10487,N_10324,N_10398);
and U10488 (N_10488,N_10270,N_10326);
or U10489 (N_10489,N_10236,N_10283);
nand U10490 (N_10490,N_10345,N_10284);
nand U10491 (N_10491,N_10221,N_10274);
nand U10492 (N_10492,N_10237,N_10350);
xor U10493 (N_10493,N_10300,N_10333);
or U10494 (N_10494,N_10335,N_10346);
xnor U10495 (N_10495,N_10276,N_10391);
and U10496 (N_10496,N_10292,N_10382);
and U10497 (N_10497,N_10331,N_10377);
nor U10498 (N_10498,N_10344,N_10216);
xor U10499 (N_10499,N_10227,N_10316);
and U10500 (N_10500,N_10235,N_10306);
or U10501 (N_10501,N_10226,N_10219);
and U10502 (N_10502,N_10329,N_10202);
xor U10503 (N_10503,N_10260,N_10272);
nand U10504 (N_10504,N_10355,N_10291);
nand U10505 (N_10505,N_10317,N_10393);
xnor U10506 (N_10506,N_10263,N_10368);
xor U10507 (N_10507,N_10336,N_10244);
or U10508 (N_10508,N_10370,N_10302);
nor U10509 (N_10509,N_10394,N_10300);
and U10510 (N_10510,N_10284,N_10223);
or U10511 (N_10511,N_10378,N_10399);
or U10512 (N_10512,N_10397,N_10326);
or U10513 (N_10513,N_10354,N_10390);
nand U10514 (N_10514,N_10359,N_10259);
xor U10515 (N_10515,N_10293,N_10238);
xor U10516 (N_10516,N_10380,N_10386);
nand U10517 (N_10517,N_10349,N_10304);
xor U10518 (N_10518,N_10292,N_10222);
nor U10519 (N_10519,N_10384,N_10260);
nor U10520 (N_10520,N_10286,N_10201);
nor U10521 (N_10521,N_10306,N_10214);
xnor U10522 (N_10522,N_10385,N_10293);
nor U10523 (N_10523,N_10399,N_10334);
or U10524 (N_10524,N_10258,N_10259);
xnor U10525 (N_10525,N_10211,N_10258);
xor U10526 (N_10526,N_10231,N_10237);
nor U10527 (N_10527,N_10245,N_10285);
or U10528 (N_10528,N_10279,N_10211);
and U10529 (N_10529,N_10254,N_10236);
nand U10530 (N_10530,N_10291,N_10382);
nand U10531 (N_10531,N_10322,N_10327);
or U10532 (N_10532,N_10300,N_10375);
nand U10533 (N_10533,N_10200,N_10349);
and U10534 (N_10534,N_10339,N_10308);
nand U10535 (N_10535,N_10357,N_10301);
nor U10536 (N_10536,N_10257,N_10320);
nor U10537 (N_10537,N_10318,N_10397);
or U10538 (N_10538,N_10362,N_10310);
nand U10539 (N_10539,N_10326,N_10271);
xnor U10540 (N_10540,N_10375,N_10221);
and U10541 (N_10541,N_10375,N_10368);
xnor U10542 (N_10542,N_10324,N_10343);
nor U10543 (N_10543,N_10350,N_10259);
and U10544 (N_10544,N_10293,N_10314);
nor U10545 (N_10545,N_10244,N_10363);
or U10546 (N_10546,N_10206,N_10350);
and U10547 (N_10547,N_10388,N_10330);
or U10548 (N_10548,N_10319,N_10365);
nand U10549 (N_10549,N_10395,N_10236);
and U10550 (N_10550,N_10362,N_10292);
and U10551 (N_10551,N_10367,N_10351);
or U10552 (N_10552,N_10260,N_10348);
nor U10553 (N_10553,N_10360,N_10206);
and U10554 (N_10554,N_10367,N_10276);
xor U10555 (N_10555,N_10368,N_10339);
and U10556 (N_10556,N_10337,N_10394);
nor U10557 (N_10557,N_10229,N_10288);
or U10558 (N_10558,N_10301,N_10247);
nand U10559 (N_10559,N_10373,N_10366);
or U10560 (N_10560,N_10376,N_10323);
nand U10561 (N_10561,N_10297,N_10261);
and U10562 (N_10562,N_10378,N_10307);
nor U10563 (N_10563,N_10391,N_10393);
nand U10564 (N_10564,N_10390,N_10350);
nor U10565 (N_10565,N_10244,N_10203);
xor U10566 (N_10566,N_10310,N_10350);
xor U10567 (N_10567,N_10347,N_10383);
nor U10568 (N_10568,N_10226,N_10207);
nor U10569 (N_10569,N_10299,N_10269);
or U10570 (N_10570,N_10368,N_10320);
nand U10571 (N_10571,N_10349,N_10249);
or U10572 (N_10572,N_10323,N_10277);
nand U10573 (N_10573,N_10344,N_10346);
and U10574 (N_10574,N_10276,N_10258);
or U10575 (N_10575,N_10251,N_10365);
xor U10576 (N_10576,N_10305,N_10204);
nand U10577 (N_10577,N_10284,N_10392);
or U10578 (N_10578,N_10379,N_10364);
nand U10579 (N_10579,N_10211,N_10207);
nand U10580 (N_10580,N_10386,N_10381);
or U10581 (N_10581,N_10221,N_10359);
xnor U10582 (N_10582,N_10244,N_10271);
or U10583 (N_10583,N_10250,N_10249);
or U10584 (N_10584,N_10241,N_10327);
nand U10585 (N_10585,N_10360,N_10385);
xor U10586 (N_10586,N_10212,N_10256);
or U10587 (N_10587,N_10398,N_10224);
and U10588 (N_10588,N_10251,N_10283);
or U10589 (N_10589,N_10216,N_10323);
xnor U10590 (N_10590,N_10339,N_10225);
or U10591 (N_10591,N_10268,N_10394);
nand U10592 (N_10592,N_10287,N_10377);
and U10593 (N_10593,N_10215,N_10223);
and U10594 (N_10594,N_10257,N_10237);
nand U10595 (N_10595,N_10280,N_10359);
or U10596 (N_10596,N_10323,N_10378);
and U10597 (N_10597,N_10386,N_10365);
xor U10598 (N_10598,N_10204,N_10247);
xor U10599 (N_10599,N_10290,N_10221);
nor U10600 (N_10600,N_10544,N_10469);
xnor U10601 (N_10601,N_10414,N_10453);
xnor U10602 (N_10602,N_10562,N_10572);
and U10603 (N_10603,N_10584,N_10542);
xnor U10604 (N_10604,N_10485,N_10431);
nor U10605 (N_10605,N_10459,N_10580);
or U10606 (N_10606,N_10408,N_10458);
nand U10607 (N_10607,N_10593,N_10555);
nand U10608 (N_10608,N_10437,N_10583);
xnor U10609 (N_10609,N_10418,N_10473);
nor U10610 (N_10610,N_10554,N_10409);
or U10611 (N_10611,N_10452,N_10471);
nor U10612 (N_10612,N_10568,N_10441);
nand U10613 (N_10613,N_10543,N_10519);
nor U10614 (N_10614,N_10428,N_10461);
xor U10615 (N_10615,N_10516,N_10528);
or U10616 (N_10616,N_10470,N_10565);
and U10617 (N_10617,N_10468,N_10403);
and U10618 (N_10618,N_10421,N_10521);
or U10619 (N_10619,N_10476,N_10535);
nand U10620 (N_10620,N_10570,N_10429);
nor U10621 (N_10621,N_10569,N_10494);
and U10622 (N_10622,N_10424,N_10430);
xor U10623 (N_10623,N_10456,N_10534);
and U10624 (N_10624,N_10422,N_10435);
nand U10625 (N_10625,N_10412,N_10552);
nor U10626 (N_10626,N_10486,N_10571);
nand U10627 (N_10627,N_10508,N_10513);
xnor U10628 (N_10628,N_10446,N_10488);
nand U10629 (N_10629,N_10523,N_10464);
xnor U10630 (N_10630,N_10445,N_10439);
nand U10631 (N_10631,N_10413,N_10492);
nand U10632 (N_10632,N_10525,N_10481);
and U10633 (N_10633,N_10427,N_10496);
or U10634 (N_10634,N_10587,N_10436);
nand U10635 (N_10635,N_10506,N_10556);
nand U10636 (N_10636,N_10529,N_10498);
and U10637 (N_10637,N_10588,N_10582);
and U10638 (N_10638,N_10457,N_10517);
or U10639 (N_10639,N_10594,N_10530);
and U10640 (N_10640,N_10503,N_10425);
nor U10641 (N_10641,N_10540,N_10433);
nor U10642 (N_10642,N_10567,N_10411);
xor U10643 (N_10643,N_10404,N_10479);
nor U10644 (N_10644,N_10415,N_10559);
xnor U10645 (N_10645,N_10560,N_10491);
nor U10646 (N_10646,N_10475,N_10440);
xnor U10647 (N_10647,N_10472,N_10581);
nand U10648 (N_10648,N_10448,N_10501);
xor U10649 (N_10649,N_10462,N_10443);
or U10650 (N_10650,N_10515,N_10589);
xor U10651 (N_10651,N_10434,N_10507);
and U10652 (N_10652,N_10480,N_10504);
nor U10653 (N_10653,N_10533,N_10487);
xnor U10654 (N_10654,N_10558,N_10574);
nor U10655 (N_10655,N_10591,N_10454);
xnor U10656 (N_10656,N_10531,N_10400);
and U10657 (N_10657,N_10539,N_10463);
and U10658 (N_10658,N_10541,N_10548);
and U10659 (N_10659,N_10490,N_10484);
and U10660 (N_10660,N_10550,N_10465);
nor U10661 (N_10661,N_10520,N_10416);
nor U10662 (N_10662,N_10512,N_10598);
or U10663 (N_10663,N_10546,N_10406);
or U10664 (N_10664,N_10538,N_10522);
and U10665 (N_10665,N_10563,N_10545);
and U10666 (N_10666,N_10438,N_10590);
nor U10667 (N_10667,N_10447,N_10509);
xor U10668 (N_10668,N_10536,N_10505);
and U10669 (N_10669,N_10575,N_10564);
xor U10670 (N_10670,N_10449,N_10502);
or U10671 (N_10671,N_10401,N_10573);
xnor U10672 (N_10672,N_10510,N_10495);
nor U10673 (N_10673,N_10489,N_10578);
and U10674 (N_10674,N_10450,N_10553);
or U10675 (N_10675,N_10474,N_10407);
nand U10676 (N_10676,N_10426,N_10551);
nor U10677 (N_10677,N_10596,N_10402);
nand U10678 (N_10678,N_10592,N_10547);
nand U10679 (N_10679,N_10526,N_10537);
nand U10680 (N_10680,N_10423,N_10419);
or U10681 (N_10681,N_10595,N_10455);
and U10682 (N_10682,N_10460,N_10566);
xnor U10683 (N_10683,N_10579,N_10417);
or U10684 (N_10684,N_10514,N_10442);
nor U10685 (N_10685,N_10518,N_10597);
and U10686 (N_10686,N_10444,N_10483);
nand U10687 (N_10687,N_10576,N_10532);
nor U10688 (N_10688,N_10527,N_10410);
and U10689 (N_10689,N_10432,N_10557);
xor U10690 (N_10690,N_10577,N_10482);
nor U10691 (N_10691,N_10599,N_10477);
xnor U10692 (N_10692,N_10493,N_10585);
or U10693 (N_10693,N_10451,N_10549);
nand U10694 (N_10694,N_10478,N_10497);
and U10695 (N_10695,N_10561,N_10420);
or U10696 (N_10696,N_10499,N_10466);
or U10697 (N_10697,N_10500,N_10405);
or U10698 (N_10698,N_10524,N_10467);
and U10699 (N_10699,N_10586,N_10511);
or U10700 (N_10700,N_10438,N_10423);
nand U10701 (N_10701,N_10496,N_10490);
and U10702 (N_10702,N_10478,N_10561);
xor U10703 (N_10703,N_10458,N_10517);
nor U10704 (N_10704,N_10441,N_10425);
and U10705 (N_10705,N_10432,N_10466);
or U10706 (N_10706,N_10540,N_10439);
nor U10707 (N_10707,N_10589,N_10402);
xor U10708 (N_10708,N_10503,N_10553);
and U10709 (N_10709,N_10490,N_10422);
xnor U10710 (N_10710,N_10544,N_10507);
xnor U10711 (N_10711,N_10557,N_10485);
or U10712 (N_10712,N_10500,N_10486);
nand U10713 (N_10713,N_10432,N_10472);
nor U10714 (N_10714,N_10566,N_10463);
or U10715 (N_10715,N_10429,N_10494);
nor U10716 (N_10716,N_10572,N_10458);
nor U10717 (N_10717,N_10436,N_10534);
or U10718 (N_10718,N_10407,N_10558);
and U10719 (N_10719,N_10484,N_10543);
nand U10720 (N_10720,N_10464,N_10417);
xnor U10721 (N_10721,N_10461,N_10430);
or U10722 (N_10722,N_10560,N_10411);
nand U10723 (N_10723,N_10408,N_10582);
nor U10724 (N_10724,N_10513,N_10463);
and U10725 (N_10725,N_10439,N_10591);
nor U10726 (N_10726,N_10472,N_10564);
nand U10727 (N_10727,N_10492,N_10594);
xor U10728 (N_10728,N_10533,N_10562);
nand U10729 (N_10729,N_10526,N_10494);
nor U10730 (N_10730,N_10471,N_10460);
nor U10731 (N_10731,N_10523,N_10507);
nor U10732 (N_10732,N_10404,N_10530);
or U10733 (N_10733,N_10427,N_10444);
or U10734 (N_10734,N_10412,N_10446);
and U10735 (N_10735,N_10466,N_10490);
nor U10736 (N_10736,N_10557,N_10403);
and U10737 (N_10737,N_10531,N_10530);
and U10738 (N_10738,N_10590,N_10543);
and U10739 (N_10739,N_10559,N_10471);
or U10740 (N_10740,N_10460,N_10549);
and U10741 (N_10741,N_10461,N_10584);
xor U10742 (N_10742,N_10444,N_10574);
or U10743 (N_10743,N_10517,N_10565);
or U10744 (N_10744,N_10566,N_10475);
or U10745 (N_10745,N_10427,N_10469);
nand U10746 (N_10746,N_10455,N_10527);
nand U10747 (N_10747,N_10541,N_10420);
or U10748 (N_10748,N_10561,N_10440);
nor U10749 (N_10749,N_10537,N_10418);
or U10750 (N_10750,N_10501,N_10524);
xor U10751 (N_10751,N_10429,N_10599);
or U10752 (N_10752,N_10561,N_10447);
and U10753 (N_10753,N_10594,N_10523);
nand U10754 (N_10754,N_10596,N_10468);
nor U10755 (N_10755,N_10450,N_10550);
nor U10756 (N_10756,N_10571,N_10595);
nand U10757 (N_10757,N_10421,N_10480);
xor U10758 (N_10758,N_10559,N_10469);
and U10759 (N_10759,N_10421,N_10488);
and U10760 (N_10760,N_10578,N_10434);
nand U10761 (N_10761,N_10565,N_10483);
nor U10762 (N_10762,N_10562,N_10502);
nor U10763 (N_10763,N_10576,N_10567);
xnor U10764 (N_10764,N_10525,N_10529);
nor U10765 (N_10765,N_10431,N_10487);
or U10766 (N_10766,N_10463,N_10410);
nor U10767 (N_10767,N_10550,N_10444);
nor U10768 (N_10768,N_10510,N_10474);
nor U10769 (N_10769,N_10525,N_10482);
or U10770 (N_10770,N_10548,N_10562);
and U10771 (N_10771,N_10455,N_10417);
nand U10772 (N_10772,N_10529,N_10448);
or U10773 (N_10773,N_10499,N_10496);
xor U10774 (N_10774,N_10490,N_10478);
or U10775 (N_10775,N_10463,N_10575);
or U10776 (N_10776,N_10412,N_10573);
xnor U10777 (N_10777,N_10434,N_10584);
nand U10778 (N_10778,N_10448,N_10559);
or U10779 (N_10779,N_10421,N_10559);
and U10780 (N_10780,N_10494,N_10456);
nor U10781 (N_10781,N_10592,N_10515);
nand U10782 (N_10782,N_10468,N_10542);
or U10783 (N_10783,N_10562,N_10440);
xor U10784 (N_10784,N_10522,N_10468);
and U10785 (N_10785,N_10598,N_10515);
or U10786 (N_10786,N_10596,N_10551);
and U10787 (N_10787,N_10525,N_10513);
nor U10788 (N_10788,N_10582,N_10434);
and U10789 (N_10789,N_10470,N_10592);
xnor U10790 (N_10790,N_10452,N_10555);
or U10791 (N_10791,N_10407,N_10471);
or U10792 (N_10792,N_10475,N_10491);
xor U10793 (N_10793,N_10483,N_10515);
xnor U10794 (N_10794,N_10432,N_10568);
xor U10795 (N_10795,N_10556,N_10477);
and U10796 (N_10796,N_10547,N_10562);
xor U10797 (N_10797,N_10586,N_10459);
nand U10798 (N_10798,N_10573,N_10586);
nand U10799 (N_10799,N_10563,N_10539);
or U10800 (N_10800,N_10674,N_10600);
and U10801 (N_10801,N_10772,N_10643);
or U10802 (N_10802,N_10604,N_10633);
xnor U10803 (N_10803,N_10642,N_10777);
and U10804 (N_10804,N_10623,N_10640);
xor U10805 (N_10805,N_10630,N_10690);
nor U10806 (N_10806,N_10771,N_10756);
and U10807 (N_10807,N_10708,N_10779);
nand U10808 (N_10808,N_10785,N_10668);
or U10809 (N_10809,N_10606,N_10629);
nor U10810 (N_10810,N_10795,N_10748);
nor U10811 (N_10811,N_10621,N_10605);
xor U10812 (N_10812,N_10787,N_10758);
xor U10813 (N_10813,N_10740,N_10673);
and U10814 (N_10814,N_10705,N_10653);
nor U10815 (N_10815,N_10737,N_10780);
nor U10816 (N_10816,N_10752,N_10738);
and U10817 (N_10817,N_10683,N_10650);
xor U10818 (N_10818,N_10611,N_10667);
or U10819 (N_10819,N_10691,N_10684);
nor U10820 (N_10820,N_10794,N_10745);
and U10821 (N_10821,N_10680,N_10628);
or U10822 (N_10822,N_10714,N_10725);
xor U10823 (N_10823,N_10636,N_10698);
and U10824 (N_10824,N_10728,N_10688);
or U10825 (N_10825,N_10721,N_10717);
xnor U10826 (N_10826,N_10760,N_10791);
xnor U10827 (N_10827,N_10726,N_10718);
xor U10828 (N_10828,N_10661,N_10746);
nand U10829 (N_10829,N_10655,N_10729);
or U10830 (N_10830,N_10639,N_10602);
xor U10831 (N_10831,N_10652,N_10701);
nand U10832 (N_10832,N_10743,N_10678);
and U10833 (N_10833,N_10637,N_10710);
xor U10834 (N_10834,N_10715,N_10731);
or U10835 (N_10835,N_10751,N_10773);
nor U10836 (N_10836,N_10682,N_10607);
nand U10837 (N_10837,N_10720,N_10749);
xor U10838 (N_10838,N_10736,N_10681);
and U10839 (N_10839,N_10744,N_10687);
nand U10840 (N_10840,N_10796,N_10646);
nand U10841 (N_10841,N_10733,N_10694);
xnor U10842 (N_10842,N_10654,N_10767);
nor U10843 (N_10843,N_10798,N_10739);
and U10844 (N_10844,N_10695,N_10709);
nor U10845 (N_10845,N_10658,N_10665);
and U10846 (N_10846,N_10641,N_10790);
and U10847 (N_10847,N_10625,N_10776);
and U10848 (N_10848,N_10662,N_10723);
nor U10849 (N_10849,N_10699,N_10686);
xnor U10850 (N_10850,N_10703,N_10719);
nand U10851 (N_10851,N_10666,N_10657);
xor U10852 (N_10852,N_10660,N_10693);
and U10853 (N_10853,N_10617,N_10618);
and U10854 (N_10854,N_10775,N_10616);
xor U10855 (N_10855,N_10626,N_10742);
nand U10856 (N_10856,N_10788,N_10645);
nor U10857 (N_10857,N_10781,N_10730);
xor U10858 (N_10858,N_10615,N_10799);
xnor U10859 (N_10859,N_10747,N_10784);
nand U10860 (N_10860,N_10732,N_10706);
or U10861 (N_10861,N_10754,N_10679);
xnor U10862 (N_10862,N_10672,N_10608);
or U10863 (N_10863,N_10757,N_10685);
or U10864 (N_10864,N_10648,N_10631);
nor U10865 (N_10865,N_10632,N_10716);
and U10866 (N_10866,N_10774,N_10638);
nand U10867 (N_10867,N_10764,N_10613);
xor U10868 (N_10868,N_10735,N_10603);
nor U10869 (N_10869,N_10620,N_10670);
or U10870 (N_10870,N_10766,N_10734);
and U10871 (N_10871,N_10769,N_10663);
and U10872 (N_10872,N_10713,N_10761);
xnor U10873 (N_10873,N_10755,N_10647);
nor U10874 (N_10874,N_10612,N_10696);
nand U10875 (N_10875,N_10778,N_10797);
nor U10876 (N_10876,N_10700,N_10677);
and U10877 (N_10877,N_10671,N_10727);
and U10878 (N_10878,N_10644,N_10707);
and U10879 (N_10879,N_10659,N_10627);
or U10880 (N_10880,N_10786,N_10624);
and U10881 (N_10881,N_10762,N_10634);
nor U10882 (N_10882,N_10741,N_10601);
nor U10883 (N_10883,N_10609,N_10704);
or U10884 (N_10884,N_10768,N_10649);
nand U10885 (N_10885,N_10676,N_10619);
or U10886 (N_10886,N_10656,N_10651);
and U10887 (N_10887,N_10692,N_10675);
nand U10888 (N_10888,N_10610,N_10793);
nand U10889 (N_10889,N_10689,N_10614);
or U10890 (N_10890,N_10759,N_10783);
or U10891 (N_10891,N_10792,N_10635);
nor U10892 (N_10892,N_10622,N_10702);
nor U10893 (N_10893,N_10724,N_10697);
nand U10894 (N_10894,N_10765,N_10763);
xnor U10895 (N_10895,N_10669,N_10664);
or U10896 (N_10896,N_10753,N_10782);
xor U10897 (N_10897,N_10789,N_10712);
or U10898 (N_10898,N_10750,N_10722);
and U10899 (N_10899,N_10770,N_10711);
or U10900 (N_10900,N_10729,N_10726);
xor U10901 (N_10901,N_10745,N_10679);
nor U10902 (N_10902,N_10603,N_10771);
nor U10903 (N_10903,N_10602,N_10697);
or U10904 (N_10904,N_10722,N_10700);
nor U10905 (N_10905,N_10603,N_10607);
xor U10906 (N_10906,N_10673,N_10662);
nor U10907 (N_10907,N_10700,N_10656);
or U10908 (N_10908,N_10659,N_10642);
and U10909 (N_10909,N_10738,N_10726);
and U10910 (N_10910,N_10615,N_10680);
or U10911 (N_10911,N_10708,N_10710);
or U10912 (N_10912,N_10704,N_10656);
and U10913 (N_10913,N_10687,N_10644);
nor U10914 (N_10914,N_10680,N_10781);
xor U10915 (N_10915,N_10698,N_10771);
or U10916 (N_10916,N_10622,N_10762);
nor U10917 (N_10917,N_10774,N_10630);
or U10918 (N_10918,N_10653,N_10649);
nor U10919 (N_10919,N_10654,N_10679);
nand U10920 (N_10920,N_10652,N_10646);
nand U10921 (N_10921,N_10600,N_10790);
and U10922 (N_10922,N_10695,N_10745);
or U10923 (N_10923,N_10756,N_10684);
and U10924 (N_10924,N_10648,N_10609);
or U10925 (N_10925,N_10688,N_10664);
and U10926 (N_10926,N_10772,N_10659);
xor U10927 (N_10927,N_10776,N_10690);
xnor U10928 (N_10928,N_10682,N_10779);
nor U10929 (N_10929,N_10740,N_10622);
nand U10930 (N_10930,N_10690,N_10611);
nand U10931 (N_10931,N_10739,N_10722);
nor U10932 (N_10932,N_10671,N_10639);
or U10933 (N_10933,N_10790,N_10603);
xor U10934 (N_10934,N_10650,N_10671);
xnor U10935 (N_10935,N_10744,N_10614);
and U10936 (N_10936,N_10725,N_10607);
xnor U10937 (N_10937,N_10697,N_10604);
nor U10938 (N_10938,N_10712,N_10693);
and U10939 (N_10939,N_10686,N_10687);
nor U10940 (N_10940,N_10608,N_10637);
nor U10941 (N_10941,N_10654,N_10639);
or U10942 (N_10942,N_10721,N_10799);
nor U10943 (N_10943,N_10699,N_10785);
nor U10944 (N_10944,N_10686,N_10713);
xor U10945 (N_10945,N_10732,N_10698);
xnor U10946 (N_10946,N_10634,N_10724);
and U10947 (N_10947,N_10788,N_10698);
and U10948 (N_10948,N_10792,N_10667);
nor U10949 (N_10949,N_10674,N_10788);
and U10950 (N_10950,N_10615,N_10611);
nand U10951 (N_10951,N_10664,N_10682);
nor U10952 (N_10952,N_10619,N_10677);
or U10953 (N_10953,N_10642,N_10734);
nor U10954 (N_10954,N_10789,N_10605);
or U10955 (N_10955,N_10716,N_10633);
xnor U10956 (N_10956,N_10600,N_10679);
and U10957 (N_10957,N_10696,N_10649);
nand U10958 (N_10958,N_10699,N_10645);
nor U10959 (N_10959,N_10666,N_10675);
nand U10960 (N_10960,N_10692,N_10687);
nor U10961 (N_10961,N_10713,N_10771);
nor U10962 (N_10962,N_10695,N_10796);
or U10963 (N_10963,N_10659,N_10791);
and U10964 (N_10964,N_10631,N_10694);
or U10965 (N_10965,N_10680,N_10621);
xnor U10966 (N_10966,N_10631,N_10789);
nand U10967 (N_10967,N_10780,N_10766);
nor U10968 (N_10968,N_10736,N_10615);
and U10969 (N_10969,N_10771,N_10793);
xor U10970 (N_10970,N_10627,N_10732);
or U10971 (N_10971,N_10766,N_10795);
or U10972 (N_10972,N_10624,N_10751);
and U10973 (N_10973,N_10604,N_10669);
or U10974 (N_10974,N_10681,N_10626);
and U10975 (N_10975,N_10609,N_10642);
and U10976 (N_10976,N_10701,N_10694);
or U10977 (N_10977,N_10741,N_10775);
nand U10978 (N_10978,N_10654,N_10603);
and U10979 (N_10979,N_10679,N_10622);
and U10980 (N_10980,N_10699,N_10794);
xnor U10981 (N_10981,N_10700,N_10652);
and U10982 (N_10982,N_10688,N_10727);
xor U10983 (N_10983,N_10728,N_10651);
xor U10984 (N_10984,N_10765,N_10717);
nand U10985 (N_10985,N_10678,N_10721);
nand U10986 (N_10986,N_10628,N_10609);
nor U10987 (N_10987,N_10765,N_10792);
xnor U10988 (N_10988,N_10652,N_10625);
or U10989 (N_10989,N_10792,N_10636);
or U10990 (N_10990,N_10718,N_10767);
xnor U10991 (N_10991,N_10798,N_10771);
nand U10992 (N_10992,N_10732,N_10736);
and U10993 (N_10993,N_10676,N_10783);
or U10994 (N_10994,N_10708,N_10783);
xor U10995 (N_10995,N_10674,N_10722);
or U10996 (N_10996,N_10718,N_10635);
nor U10997 (N_10997,N_10685,N_10734);
nand U10998 (N_10998,N_10641,N_10620);
nand U10999 (N_10999,N_10627,N_10689);
nor U11000 (N_11000,N_10960,N_10973);
xnor U11001 (N_11001,N_10832,N_10807);
xor U11002 (N_11002,N_10908,N_10822);
nand U11003 (N_11003,N_10823,N_10934);
xnor U11004 (N_11004,N_10917,N_10886);
and U11005 (N_11005,N_10880,N_10962);
and U11006 (N_11006,N_10982,N_10829);
and U11007 (N_11007,N_10996,N_10811);
nand U11008 (N_11008,N_10945,N_10994);
xnor U11009 (N_11009,N_10949,N_10935);
and U11010 (N_11010,N_10984,N_10825);
and U11011 (N_11011,N_10853,N_10901);
xnor U11012 (N_11012,N_10841,N_10963);
nand U11013 (N_11013,N_10912,N_10876);
xor U11014 (N_11014,N_10955,N_10992);
and U11015 (N_11015,N_10849,N_10900);
or U11016 (N_11016,N_10855,N_10851);
or U11017 (N_11017,N_10995,N_10896);
and U11018 (N_11018,N_10895,N_10954);
or U11019 (N_11019,N_10815,N_10881);
or U11020 (N_11020,N_10857,N_10980);
and U11021 (N_11021,N_10958,N_10991);
xnor U11022 (N_11022,N_10968,N_10967);
or U11023 (N_11023,N_10861,N_10845);
or U11024 (N_11024,N_10924,N_10905);
and U11025 (N_11025,N_10860,N_10875);
xnor U11026 (N_11026,N_10820,N_10816);
nor U11027 (N_11027,N_10938,N_10877);
or U11028 (N_11028,N_10910,N_10930);
nand U11029 (N_11029,N_10920,N_10902);
nand U11030 (N_11030,N_10810,N_10826);
xor U11031 (N_11031,N_10808,N_10847);
nand U11032 (N_11032,N_10932,N_10862);
nor U11033 (N_11033,N_10941,N_10837);
nand U11034 (N_11034,N_10821,N_10977);
and U11035 (N_11035,N_10830,N_10959);
nor U11036 (N_11036,N_10926,N_10983);
xor U11037 (N_11037,N_10892,N_10843);
or U11038 (N_11038,N_10981,N_10918);
nor U11039 (N_11039,N_10923,N_10819);
xnor U11040 (N_11040,N_10854,N_10871);
nand U11041 (N_11041,N_10928,N_10891);
nand U11042 (N_11042,N_10867,N_10801);
or U11043 (N_11043,N_10887,N_10943);
and U11044 (N_11044,N_10834,N_10971);
or U11045 (N_11045,N_10911,N_10802);
nor U11046 (N_11046,N_10956,N_10974);
nor U11047 (N_11047,N_10869,N_10884);
xnor U11048 (N_11048,N_10868,N_10833);
or U11049 (N_11049,N_10931,N_10953);
xnor U11050 (N_11050,N_10978,N_10872);
and U11051 (N_11051,N_10888,N_10937);
nand U11052 (N_11052,N_10944,N_10865);
and U11053 (N_11053,N_10836,N_10948);
and U11054 (N_11054,N_10870,N_10970);
nand U11055 (N_11055,N_10885,N_10919);
and U11056 (N_11056,N_10961,N_10976);
nor U11057 (N_11057,N_10890,N_10947);
and U11058 (N_11058,N_10927,N_10987);
nand U11059 (N_11059,N_10925,N_10812);
nor U11060 (N_11060,N_10809,N_10979);
nand U11061 (N_11061,N_10824,N_10909);
xor U11062 (N_11062,N_10831,N_10899);
xnor U11063 (N_11063,N_10844,N_10913);
or U11064 (N_11064,N_10990,N_10859);
or U11065 (N_11065,N_10894,N_10950);
and U11066 (N_11066,N_10957,N_10818);
xor U11067 (N_11067,N_10952,N_10827);
or U11068 (N_11068,N_10840,N_10997);
or U11069 (N_11069,N_10889,N_10863);
or U11070 (N_11070,N_10897,N_10904);
nand U11071 (N_11071,N_10874,N_10933);
xor U11072 (N_11072,N_10951,N_10993);
and U11073 (N_11073,N_10929,N_10966);
nand U11074 (N_11074,N_10858,N_10846);
and U11075 (N_11075,N_10848,N_10985);
nor U11076 (N_11076,N_10903,N_10805);
and U11077 (N_11077,N_10965,N_10817);
xor U11078 (N_11078,N_10856,N_10939);
nand U11079 (N_11079,N_10873,N_10882);
nand U11080 (N_11080,N_10828,N_10898);
and U11081 (N_11081,N_10878,N_10989);
or U11082 (N_11082,N_10975,N_10999);
and U11083 (N_11083,N_10883,N_10940);
and U11084 (N_11084,N_10936,N_10988);
nor U11085 (N_11085,N_10813,N_10866);
or U11086 (N_11086,N_10864,N_10921);
and U11087 (N_11087,N_10972,N_10942);
nor U11088 (N_11088,N_10839,N_10922);
or U11089 (N_11089,N_10804,N_10914);
nand U11090 (N_11090,N_10986,N_10842);
nor U11091 (N_11091,N_10946,N_10907);
nand U11092 (N_11092,N_10906,N_10964);
xnor U11093 (N_11093,N_10806,N_10800);
nand U11094 (N_11094,N_10850,N_10915);
nor U11095 (N_11095,N_10998,N_10803);
and U11096 (N_11096,N_10814,N_10916);
nor U11097 (N_11097,N_10835,N_10879);
nand U11098 (N_11098,N_10969,N_10852);
and U11099 (N_11099,N_10893,N_10838);
nand U11100 (N_11100,N_10995,N_10801);
and U11101 (N_11101,N_10860,N_10911);
or U11102 (N_11102,N_10917,N_10823);
nor U11103 (N_11103,N_10951,N_10932);
nand U11104 (N_11104,N_10820,N_10807);
xor U11105 (N_11105,N_10936,N_10912);
xor U11106 (N_11106,N_10989,N_10817);
and U11107 (N_11107,N_10996,N_10879);
xor U11108 (N_11108,N_10835,N_10816);
or U11109 (N_11109,N_10886,N_10980);
or U11110 (N_11110,N_10816,N_10930);
xor U11111 (N_11111,N_10840,N_10895);
or U11112 (N_11112,N_10863,N_10933);
xor U11113 (N_11113,N_10979,N_10978);
nand U11114 (N_11114,N_10997,N_10943);
nand U11115 (N_11115,N_10866,N_10948);
xnor U11116 (N_11116,N_10814,N_10801);
nor U11117 (N_11117,N_10821,N_10926);
xor U11118 (N_11118,N_10857,N_10970);
nand U11119 (N_11119,N_10875,N_10926);
or U11120 (N_11120,N_10801,N_10955);
nor U11121 (N_11121,N_10898,N_10860);
or U11122 (N_11122,N_10957,N_10933);
nand U11123 (N_11123,N_10820,N_10846);
nor U11124 (N_11124,N_10901,N_10813);
nand U11125 (N_11125,N_10863,N_10985);
xor U11126 (N_11126,N_10972,N_10902);
or U11127 (N_11127,N_10822,N_10980);
nand U11128 (N_11128,N_10927,N_10804);
or U11129 (N_11129,N_10840,N_10832);
and U11130 (N_11130,N_10965,N_10923);
xnor U11131 (N_11131,N_10829,N_10980);
nand U11132 (N_11132,N_10998,N_10814);
or U11133 (N_11133,N_10912,N_10969);
nor U11134 (N_11134,N_10871,N_10965);
and U11135 (N_11135,N_10863,N_10875);
nand U11136 (N_11136,N_10808,N_10874);
xnor U11137 (N_11137,N_10855,N_10930);
nor U11138 (N_11138,N_10933,N_10867);
and U11139 (N_11139,N_10805,N_10978);
nand U11140 (N_11140,N_10901,N_10993);
xor U11141 (N_11141,N_10877,N_10887);
and U11142 (N_11142,N_10972,N_10970);
or U11143 (N_11143,N_10995,N_10960);
or U11144 (N_11144,N_10977,N_10972);
or U11145 (N_11145,N_10828,N_10853);
nand U11146 (N_11146,N_10800,N_10815);
nand U11147 (N_11147,N_10982,N_10865);
xnor U11148 (N_11148,N_10882,N_10899);
nor U11149 (N_11149,N_10894,N_10918);
nor U11150 (N_11150,N_10818,N_10950);
or U11151 (N_11151,N_10986,N_10874);
xor U11152 (N_11152,N_10956,N_10997);
nor U11153 (N_11153,N_10848,N_10916);
and U11154 (N_11154,N_10930,N_10951);
and U11155 (N_11155,N_10819,N_10910);
and U11156 (N_11156,N_10838,N_10883);
nor U11157 (N_11157,N_10996,N_10866);
nand U11158 (N_11158,N_10937,N_10972);
nand U11159 (N_11159,N_10808,N_10802);
xor U11160 (N_11160,N_10837,N_10981);
nor U11161 (N_11161,N_10815,N_10834);
xnor U11162 (N_11162,N_10911,N_10924);
or U11163 (N_11163,N_10803,N_10997);
and U11164 (N_11164,N_10947,N_10982);
nor U11165 (N_11165,N_10882,N_10811);
or U11166 (N_11166,N_10807,N_10943);
and U11167 (N_11167,N_10912,N_10996);
nand U11168 (N_11168,N_10830,N_10829);
and U11169 (N_11169,N_10849,N_10899);
nor U11170 (N_11170,N_10920,N_10881);
and U11171 (N_11171,N_10837,N_10992);
xnor U11172 (N_11172,N_10843,N_10817);
or U11173 (N_11173,N_10808,N_10961);
and U11174 (N_11174,N_10996,N_10880);
nor U11175 (N_11175,N_10953,N_10981);
nor U11176 (N_11176,N_10962,N_10985);
nor U11177 (N_11177,N_10911,N_10847);
and U11178 (N_11178,N_10845,N_10872);
or U11179 (N_11179,N_10905,N_10820);
nand U11180 (N_11180,N_10852,N_10923);
nand U11181 (N_11181,N_10960,N_10992);
or U11182 (N_11182,N_10823,N_10833);
or U11183 (N_11183,N_10902,N_10896);
or U11184 (N_11184,N_10895,N_10949);
or U11185 (N_11185,N_10872,N_10861);
and U11186 (N_11186,N_10914,N_10901);
nand U11187 (N_11187,N_10873,N_10834);
xnor U11188 (N_11188,N_10854,N_10878);
or U11189 (N_11189,N_10907,N_10876);
xor U11190 (N_11190,N_10853,N_10943);
nor U11191 (N_11191,N_10882,N_10975);
nor U11192 (N_11192,N_10980,N_10879);
or U11193 (N_11193,N_10922,N_10969);
nand U11194 (N_11194,N_10894,N_10805);
and U11195 (N_11195,N_10889,N_10869);
xnor U11196 (N_11196,N_10966,N_10836);
and U11197 (N_11197,N_10813,N_10918);
nor U11198 (N_11198,N_10854,N_10864);
nand U11199 (N_11199,N_10921,N_10827);
xnor U11200 (N_11200,N_11016,N_11055);
xnor U11201 (N_11201,N_11167,N_11110);
nor U11202 (N_11202,N_11003,N_11047);
nor U11203 (N_11203,N_11041,N_11120);
and U11204 (N_11204,N_11102,N_11159);
and U11205 (N_11205,N_11015,N_11028);
or U11206 (N_11206,N_11031,N_11199);
nand U11207 (N_11207,N_11124,N_11181);
xor U11208 (N_11208,N_11065,N_11054);
nor U11209 (N_11209,N_11088,N_11180);
nand U11210 (N_11210,N_11033,N_11166);
nor U11211 (N_11211,N_11107,N_11068);
nor U11212 (N_11212,N_11182,N_11138);
nand U11213 (N_11213,N_11032,N_11061);
nand U11214 (N_11214,N_11052,N_11184);
nor U11215 (N_11215,N_11073,N_11083);
nand U11216 (N_11216,N_11057,N_11039);
or U11217 (N_11217,N_11070,N_11169);
and U11218 (N_11218,N_11179,N_11013);
nand U11219 (N_11219,N_11037,N_11079);
nor U11220 (N_11220,N_11091,N_11092);
nand U11221 (N_11221,N_11020,N_11171);
nand U11222 (N_11222,N_11130,N_11040);
nor U11223 (N_11223,N_11168,N_11077);
nor U11224 (N_11224,N_11183,N_11150);
or U11225 (N_11225,N_11017,N_11142);
nor U11226 (N_11226,N_11140,N_11178);
xor U11227 (N_11227,N_11008,N_11072);
or U11228 (N_11228,N_11007,N_11044);
nand U11229 (N_11229,N_11074,N_11164);
and U11230 (N_11230,N_11122,N_11121);
and U11231 (N_11231,N_11117,N_11104);
and U11232 (N_11232,N_11030,N_11145);
or U11233 (N_11233,N_11005,N_11112);
nand U11234 (N_11234,N_11177,N_11135);
nor U11235 (N_11235,N_11038,N_11100);
and U11236 (N_11236,N_11006,N_11198);
and U11237 (N_11237,N_11108,N_11196);
nor U11238 (N_11238,N_11018,N_11048);
or U11239 (N_11239,N_11195,N_11134);
or U11240 (N_11240,N_11146,N_11149);
or U11241 (N_11241,N_11123,N_11001);
nor U11242 (N_11242,N_11131,N_11009);
nor U11243 (N_11243,N_11089,N_11049);
and U11244 (N_11244,N_11082,N_11046);
and U11245 (N_11245,N_11059,N_11012);
or U11246 (N_11246,N_11053,N_11187);
nor U11247 (N_11247,N_11098,N_11050);
xor U11248 (N_11248,N_11114,N_11151);
and U11249 (N_11249,N_11034,N_11193);
or U11250 (N_11250,N_11139,N_11078);
nor U11251 (N_11251,N_11148,N_11099);
nand U11252 (N_11252,N_11185,N_11076);
or U11253 (N_11253,N_11192,N_11080);
xor U11254 (N_11254,N_11186,N_11160);
nand U11255 (N_11255,N_11118,N_11105);
nand U11256 (N_11256,N_11188,N_11101);
and U11257 (N_11257,N_11090,N_11109);
nor U11258 (N_11258,N_11060,N_11069);
nand U11259 (N_11259,N_11066,N_11093);
nor U11260 (N_11260,N_11056,N_11154);
and U11261 (N_11261,N_11116,N_11172);
xor U11262 (N_11262,N_11096,N_11143);
nand U11263 (N_11263,N_11111,N_11197);
xnor U11264 (N_11264,N_11141,N_11119);
and U11265 (N_11265,N_11106,N_11024);
or U11266 (N_11266,N_11042,N_11165);
nand U11267 (N_11267,N_11085,N_11062);
nor U11268 (N_11268,N_11132,N_11063);
nor U11269 (N_11269,N_11162,N_11086);
nor U11270 (N_11270,N_11045,N_11155);
or U11271 (N_11271,N_11021,N_11071);
nor U11272 (N_11272,N_11103,N_11027);
nor U11273 (N_11273,N_11084,N_11174);
and U11274 (N_11274,N_11163,N_11097);
nand U11275 (N_11275,N_11023,N_11126);
nor U11276 (N_11276,N_11022,N_11170);
and U11277 (N_11277,N_11025,N_11190);
and U11278 (N_11278,N_11004,N_11036);
nand U11279 (N_11279,N_11029,N_11156);
xnor U11280 (N_11280,N_11035,N_11094);
and U11281 (N_11281,N_11129,N_11136);
xnor U11282 (N_11282,N_11194,N_11189);
and U11283 (N_11283,N_11153,N_11095);
nor U11284 (N_11284,N_11115,N_11158);
or U11285 (N_11285,N_11067,N_11161);
and U11286 (N_11286,N_11051,N_11000);
nor U11287 (N_11287,N_11147,N_11133);
and U11288 (N_11288,N_11026,N_11176);
xor U11289 (N_11289,N_11144,N_11137);
xor U11290 (N_11290,N_11043,N_11128);
and U11291 (N_11291,N_11002,N_11087);
or U11292 (N_11292,N_11019,N_11127);
and U11293 (N_11293,N_11157,N_11058);
and U11294 (N_11294,N_11191,N_11125);
or U11295 (N_11295,N_11011,N_11010);
xor U11296 (N_11296,N_11064,N_11113);
and U11297 (N_11297,N_11173,N_11014);
nand U11298 (N_11298,N_11152,N_11081);
nand U11299 (N_11299,N_11075,N_11175);
nor U11300 (N_11300,N_11032,N_11196);
nor U11301 (N_11301,N_11114,N_11057);
and U11302 (N_11302,N_11006,N_11120);
or U11303 (N_11303,N_11172,N_11080);
nor U11304 (N_11304,N_11014,N_11004);
xnor U11305 (N_11305,N_11199,N_11060);
xnor U11306 (N_11306,N_11112,N_11077);
nand U11307 (N_11307,N_11076,N_11048);
nor U11308 (N_11308,N_11094,N_11136);
and U11309 (N_11309,N_11143,N_11111);
and U11310 (N_11310,N_11190,N_11118);
nand U11311 (N_11311,N_11093,N_11024);
or U11312 (N_11312,N_11024,N_11068);
xor U11313 (N_11313,N_11123,N_11097);
xnor U11314 (N_11314,N_11079,N_11181);
xor U11315 (N_11315,N_11174,N_11170);
xor U11316 (N_11316,N_11005,N_11010);
nand U11317 (N_11317,N_11095,N_11148);
nor U11318 (N_11318,N_11084,N_11007);
nand U11319 (N_11319,N_11175,N_11126);
nand U11320 (N_11320,N_11069,N_11161);
or U11321 (N_11321,N_11107,N_11066);
nand U11322 (N_11322,N_11161,N_11137);
or U11323 (N_11323,N_11138,N_11069);
or U11324 (N_11324,N_11183,N_11178);
or U11325 (N_11325,N_11197,N_11098);
nor U11326 (N_11326,N_11028,N_11163);
nor U11327 (N_11327,N_11059,N_11107);
nand U11328 (N_11328,N_11195,N_11111);
nor U11329 (N_11329,N_11087,N_11182);
nor U11330 (N_11330,N_11180,N_11145);
nand U11331 (N_11331,N_11168,N_11154);
and U11332 (N_11332,N_11159,N_11034);
or U11333 (N_11333,N_11068,N_11074);
nand U11334 (N_11334,N_11051,N_11096);
xor U11335 (N_11335,N_11074,N_11084);
and U11336 (N_11336,N_11190,N_11080);
nor U11337 (N_11337,N_11004,N_11001);
xnor U11338 (N_11338,N_11006,N_11042);
or U11339 (N_11339,N_11148,N_11050);
xor U11340 (N_11340,N_11111,N_11155);
xnor U11341 (N_11341,N_11091,N_11159);
nand U11342 (N_11342,N_11110,N_11095);
or U11343 (N_11343,N_11136,N_11074);
nor U11344 (N_11344,N_11189,N_11174);
nand U11345 (N_11345,N_11178,N_11160);
and U11346 (N_11346,N_11082,N_11054);
or U11347 (N_11347,N_11184,N_11188);
and U11348 (N_11348,N_11032,N_11119);
and U11349 (N_11349,N_11019,N_11119);
and U11350 (N_11350,N_11005,N_11026);
xor U11351 (N_11351,N_11185,N_11058);
nand U11352 (N_11352,N_11072,N_11187);
xor U11353 (N_11353,N_11103,N_11176);
and U11354 (N_11354,N_11023,N_11067);
and U11355 (N_11355,N_11084,N_11176);
or U11356 (N_11356,N_11189,N_11054);
nand U11357 (N_11357,N_11065,N_11135);
nand U11358 (N_11358,N_11000,N_11017);
and U11359 (N_11359,N_11183,N_11016);
or U11360 (N_11360,N_11175,N_11197);
nor U11361 (N_11361,N_11027,N_11074);
and U11362 (N_11362,N_11193,N_11072);
xor U11363 (N_11363,N_11023,N_11137);
nand U11364 (N_11364,N_11080,N_11142);
xnor U11365 (N_11365,N_11147,N_11023);
xor U11366 (N_11366,N_11068,N_11084);
and U11367 (N_11367,N_11042,N_11096);
nor U11368 (N_11368,N_11172,N_11025);
and U11369 (N_11369,N_11042,N_11033);
xnor U11370 (N_11370,N_11199,N_11148);
or U11371 (N_11371,N_11077,N_11004);
xor U11372 (N_11372,N_11004,N_11184);
and U11373 (N_11373,N_11060,N_11093);
xor U11374 (N_11374,N_11150,N_11195);
and U11375 (N_11375,N_11078,N_11156);
and U11376 (N_11376,N_11006,N_11084);
and U11377 (N_11377,N_11183,N_11058);
xor U11378 (N_11378,N_11071,N_11049);
or U11379 (N_11379,N_11024,N_11124);
xor U11380 (N_11380,N_11006,N_11037);
nor U11381 (N_11381,N_11041,N_11074);
nor U11382 (N_11382,N_11044,N_11008);
nor U11383 (N_11383,N_11179,N_11159);
or U11384 (N_11384,N_11012,N_11195);
nand U11385 (N_11385,N_11037,N_11050);
nor U11386 (N_11386,N_11090,N_11134);
and U11387 (N_11387,N_11112,N_11149);
and U11388 (N_11388,N_11101,N_11051);
and U11389 (N_11389,N_11154,N_11083);
nand U11390 (N_11390,N_11194,N_11136);
and U11391 (N_11391,N_11188,N_11071);
xnor U11392 (N_11392,N_11018,N_11108);
nor U11393 (N_11393,N_11136,N_11162);
nand U11394 (N_11394,N_11164,N_11027);
or U11395 (N_11395,N_11060,N_11067);
nand U11396 (N_11396,N_11040,N_11049);
nor U11397 (N_11397,N_11159,N_11152);
xor U11398 (N_11398,N_11182,N_11038);
or U11399 (N_11399,N_11005,N_11036);
xor U11400 (N_11400,N_11266,N_11232);
xnor U11401 (N_11401,N_11240,N_11353);
xor U11402 (N_11402,N_11226,N_11234);
or U11403 (N_11403,N_11205,N_11385);
nor U11404 (N_11404,N_11337,N_11316);
nand U11405 (N_11405,N_11368,N_11397);
or U11406 (N_11406,N_11259,N_11349);
or U11407 (N_11407,N_11283,N_11386);
xnor U11408 (N_11408,N_11229,N_11372);
and U11409 (N_11409,N_11378,N_11258);
nand U11410 (N_11410,N_11328,N_11215);
or U11411 (N_11411,N_11202,N_11216);
or U11412 (N_11412,N_11231,N_11351);
nand U11413 (N_11413,N_11338,N_11246);
nor U11414 (N_11414,N_11369,N_11322);
or U11415 (N_11415,N_11396,N_11302);
nor U11416 (N_11416,N_11294,N_11207);
nor U11417 (N_11417,N_11325,N_11334);
and U11418 (N_11418,N_11279,N_11267);
nand U11419 (N_11419,N_11220,N_11223);
and U11420 (N_11420,N_11305,N_11354);
nor U11421 (N_11421,N_11323,N_11309);
and U11422 (N_11422,N_11212,N_11342);
nor U11423 (N_11423,N_11384,N_11371);
nor U11424 (N_11424,N_11335,N_11208);
nor U11425 (N_11425,N_11376,N_11332);
and U11426 (N_11426,N_11245,N_11331);
xnor U11427 (N_11427,N_11214,N_11343);
xnor U11428 (N_11428,N_11319,N_11224);
and U11429 (N_11429,N_11261,N_11352);
nand U11430 (N_11430,N_11390,N_11284);
nand U11431 (N_11431,N_11285,N_11336);
or U11432 (N_11432,N_11381,N_11228);
or U11433 (N_11433,N_11315,N_11317);
nand U11434 (N_11434,N_11277,N_11255);
nor U11435 (N_11435,N_11311,N_11263);
nor U11436 (N_11436,N_11356,N_11296);
xor U11437 (N_11437,N_11395,N_11257);
nor U11438 (N_11438,N_11290,N_11300);
nand U11439 (N_11439,N_11252,N_11227);
nor U11440 (N_11440,N_11268,N_11236);
or U11441 (N_11441,N_11387,N_11286);
or U11442 (N_11442,N_11270,N_11204);
xor U11443 (N_11443,N_11238,N_11324);
or U11444 (N_11444,N_11295,N_11389);
or U11445 (N_11445,N_11314,N_11373);
nor U11446 (N_11446,N_11347,N_11253);
or U11447 (N_11447,N_11293,N_11248);
xor U11448 (N_11448,N_11289,N_11219);
or U11449 (N_11449,N_11209,N_11312);
and U11450 (N_11450,N_11375,N_11382);
nand U11451 (N_11451,N_11262,N_11237);
and U11452 (N_11452,N_11281,N_11200);
or U11453 (N_11453,N_11221,N_11249);
and U11454 (N_11454,N_11393,N_11276);
nor U11455 (N_11455,N_11287,N_11358);
xor U11456 (N_11456,N_11361,N_11273);
or U11457 (N_11457,N_11307,N_11297);
xnor U11458 (N_11458,N_11201,N_11303);
or U11459 (N_11459,N_11391,N_11340);
or U11460 (N_11460,N_11222,N_11364);
nand U11461 (N_11461,N_11318,N_11239);
and U11462 (N_11462,N_11271,N_11230);
xor U11463 (N_11463,N_11339,N_11394);
xor U11464 (N_11464,N_11365,N_11346);
or U11465 (N_11465,N_11313,N_11244);
nand U11466 (N_11466,N_11374,N_11308);
xor U11467 (N_11467,N_11377,N_11233);
nor U11468 (N_11468,N_11254,N_11392);
nor U11469 (N_11469,N_11304,N_11213);
or U11470 (N_11470,N_11379,N_11366);
xor U11471 (N_11471,N_11383,N_11264);
xnor U11472 (N_11472,N_11211,N_11367);
and U11473 (N_11473,N_11363,N_11345);
xor U11474 (N_11474,N_11329,N_11218);
or U11475 (N_11475,N_11350,N_11243);
xor U11476 (N_11476,N_11370,N_11260);
nor U11477 (N_11477,N_11269,N_11288);
nand U11478 (N_11478,N_11251,N_11320);
nand U11479 (N_11479,N_11241,N_11355);
nor U11480 (N_11480,N_11256,N_11292);
xor U11481 (N_11481,N_11278,N_11282);
and U11482 (N_11482,N_11298,N_11210);
or U11483 (N_11483,N_11301,N_11330);
nor U11484 (N_11484,N_11360,N_11265);
nor U11485 (N_11485,N_11272,N_11206);
and U11486 (N_11486,N_11362,N_11357);
xnor U11487 (N_11487,N_11299,N_11348);
xor U11488 (N_11488,N_11380,N_11359);
xnor U11489 (N_11489,N_11242,N_11388);
xnor U11490 (N_11490,N_11225,N_11333);
xor U11491 (N_11491,N_11341,N_11344);
or U11492 (N_11492,N_11399,N_11203);
nand U11493 (N_11493,N_11280,N_11250);
xnor U11494 (N_11494,N_11274,N_11235);
nor U11495 (N_11495,N_11291,N_11275);
xor U11496 (N_11496,N_11321,N_11217);
and U11497 (N_11497,N_11327,N_11326);
and U11498 (N_11498,N_11247,N_11310);
and U11499 (N_11499,N_11306,N_11398);
nand U11500 (N_11500,N_11284,N_11285);
nand U11501 (N_11501,N_11322,N_11381);
xor U11502 (N_11502,N_11235,N_11224);
or U11503 (N_11503,N_11242,N_11365);
xnor U11504 (N_11504,N_11205,N_11233);
nor U11505 (N_11505,N_11230,N_11318);
and U11506 (N_11506,N_11217,N_11214);
or U11507 (N_11507,N_11222,N_11288);
xor U11508 (N_11508,N_11394,N_11212);
xnor U11509 (N_11509,N_11259,N_11318);
nor U11510 (N_11510,N_11321,N_11387);
nand U11511 (N_11511,N_11243,N_11308);
or U11512 (N_11512,N_11316,N_11264);
nand U11513 (N_11513,N_11285,N_11227);
nor U11514 (N_11514,N_11323,N_11382);
nor U11515 (N_11515,N_11242,N_11390);
nand U11516 (N_11516,N_11331,N_11373);
or U11517 (N_11517,N_11384,N_11397);
nand U11518 (N_11518,N_11381,N_11201);
nor U11519 (N_11519,N_11305,N_11327);
xnor U11520 (N_11520,N_11269,N_11388);
xnor U11521 (N_11521,N_11306,N_11347);
or U11522 (N_11522,N_11338,N_11351);
and U11523 (N_11523,N_11298,N_11251);
and U11524 (N_11524,N_11393,N_11321);
nor U11525 (N_11525,N_11389,N_11232);
and U11526 (N_11526,N_11367,N_11236);
xnor U11527 (N_11527,N_11245,N_11370);
xor U11528 (N_11528,N_11382,N_11357);
xnor U11529 (N_11529,N_11291,N_11260);
and U11530 (N_11530,N_11356,N_11358);
xor U11531 (N_11531,N_11310,N_11284);
nand U11532 (N_11532,N_11369,N_11203);
and U11533 (N_11533,N_11324,N_11377);
or U11534 (N_11534,N_11219,N_11290);
nor U11535 (N_11535,N_11250,N_11219);
and U11536 (N_11536,N_11263,N_11300);
nor U11537 (N_11537,N_11332,N_11247);
xor U11538 (N_11538,N_11334,N_11214);
and U11539 (N_11539,N_11296,N_11376);
and U11540 (N_11540,N_11287,N_11251);
nand U11541 (N_11541,N_11322,N_11221);
nor U11542 (N_11542,N_11389,N_11323);
xor U11543 (N_11543,N_11324,N_11312);
or U11544 (N_11544,N_11322,N_11302);
or U11545 (N_11545,N_11384,N_11325);
nor U11546 (N_11546,N_11210,N_11310);
or U11547 (N_11547,N_11296,N_11395);
nand U11548 (N_11548,N_11395,N_11218);
xor U11549 (N_11549,N_11384,N_11267);
nand U11550 (N_11550,N_11225,N_11396);
nor U11551 (N_11551,N_11259,N_11227);
xnor U11552 (N_11552,N_11359,N_11347);
nor U11553 (N_11553,N_11316,N_11215);
or U11554 (N_11554,N_11374,N_11391);
or U11555 (N_11555,N_11318,N_11348);
and U11556 (N_11556,N_11332,N_11303);
nor U11557 (N_11557,N_11323,N_11267);
xor U11558 (N_11558,N_11361,N_11243);
xnor U11559 (N_11559,N_11348,N_11351);
nand U11560 (N_11560,N_11258,N_11277);
and U11561 (N_11561,N_11262,N_11266);
nand U11562 (N_11562,N_11394,N_11321);
and U11563 (N_11563,N_11355,N_11375);
xnor U11564 (N_11564,N_11395,N_11364);
nor U11565 (N_11565,N_11313,N_11355);
and U11566 (N_11566,N_11227,N_11360);
or U11567 (N_11567,N_11309,N_11397);
or U11568 (N_11568,N_11212,N_11315);
and U11569 (N_11569,N_11339,N_11239);
nor U11570 (N_11570,N_11301,N_11283);
xnor U11571 (N_11571,N_11346,N_11277);
nor U11572 (N_11572,N_11387,N_11398);
nand U11573 (N_11573,N_11265,N_11238);
xor U11574 (N_11574,N_11219,N_11302);
nor U11575 (N_11575,N_11390,N_11355);
nand U11576 (N_11576,N_11248,N_11211);
or U11577 (N_11577,N_11219,N_11296);
and U11578 (N_11578,N_11244,N_11291);
xor U11579 (N_11579,N_11383,N_11203);
xor U11580 (N_11580,N_11348,N_11394);
and U11581 (N_11581,N_11327,N_11243);
nand U11582 (N_11582,N_11214,N_11284);
nand U11583 (N_11583,N_11303,N_11344);
nand U11584 (N_11584,N_11208,N_11266);
and U11585 (N_11585,N_11342,N_11365);
xor U11586 (N_11586,N_11335,N_11342);
nor U11587 (N_11587,N_11278,N_11303);
xor U11588 (N_11588,N_11384,N_11298);
nor U11589 (N_11589,N_11281,N_11291);
nand U11590 (N_11590,N_11340,N_11230);
xor U11591 (N_11591,N_11268,N_11369);
xor U11592 (N_11592,N_11320,N_11301);
xnor U11593 (N_11593,N_11284,N_11327);
and U11594 (N_11594,N_11378,N_11280);
or U11595 (N_11595,N_11347,N_11323);
nand U11596 (N_11596,N_11312,N_11213);
and U11597 (N_11597,N_11226,N_11343);
and U11598 (N_11598,N_11306,N_11268);
or U11599 (N_11599,N_11333,N_11258);
nor U11600 (N_11600,N_11580,N_11453);
nand U11601 (N_11601,N_11534,N_11566);
and U11602 (N_11602,N_11513,N_11537);
and U11603 (N_11603,N_11412,N_11515);
nor U11604 (N_11604,N_11555,N_11583);
and U11605 (N_11605,N_11527,N_11572);
or U11606 (N_11606,N_11519,N_11461);
nor U11607 (N_11607,N_11478,N_11538);
nor U11608 (N_11608,N_11535,N_11496);
nand U11609 (N_11609,N_11545,N_11563);
xor U11610 (N_11610,N_11495,N_11526);
nand U11611 (N_11611,N_11547,N_11469);
nor U11612 (N_11612,N_11414,N_11556);
xor U11613 (N_11613,N_11400,N_11570);
nor U11614 (N_11614,N_11588,N_11521);
xnor U11615 (N_11615,N_11486,N_11559);
xnor U11616 (N_11616,N_11404,N_11574);
nand U11617 (N_11617,N_11464,N_11549);
xnor U11618 (N_11618,N_11592,N_11455);
or U11619 (N_11619,N_11418,N_11440);
or U11620 (N_11620,N_11437,N_11475);
nand U11621 (N_11621,N_11434,N_11500);
nor U11622 (N_11622,N_11462,N_11531);
nor U11623 (N_11623,N_11470,N_11512);
xnor U11624 (N_11624,N_11401,N_11465);
xor U11625 (N_11625,N_11561,N_11503);
xor U11626 (N_11626,N_11528,N_11514);
xor U11627 (N_11627,N_11449,N_11494);
nor U11628 (N_11628,N_11517,N_11571);
nand U11629 (N_11629,N_11430,N_11473);
or U11630 (N_11630,N_11573,N_11459);
xnor U11631 (N_11631,N_11541,N_11553);
nand U11632 (N_11632,N_11522,N_11460);
xnor U11633 (N_11633,N_11581,N_11456);
nand U11634 (N_11634,N_11591,N_11427);
and U11635 (N_11635,N_11468,N_11419);
nor U11636 (N_11636,N_11585,N_11596);
nand U11637 (N_11637,N_11425,N_11407);
xor U11638 (N_11638,N_11524,N_11405);
and U11639 (N_11639,N_11577,N_11586);
xor U11640 (N_11640,N_11540,N_11491);
xnor U11641 (N_11641,N_11584,N_11463);
or U11642 (N_11642,N_11410,N_11450);
xor U11643 (N_11643,N_11428,N_11506);
nand U11644 (N_11644,N_11599,N_11417);
xnor U11645 (N_11645,N_11472,N_11489);
or U11646 (N_11646,N_11546,N_11497);
or U11647 (N_11647,N_11569,N_11516);
and U11648 (N_11648,N_11594,N_11420);
xnor U11649 (N_11649,N_11567,N_11436);
nand U11650 (N_11650,N_11446,N_11415);
nand U11651 (N_11651,N_11426,N_11530);
nand U11652 (N_11652,N_11505,N_11451);
or U11653 (N_11653,N_11507,N_11432);
nor U11654 (N_11654,N_11433,N_11443);
and U11655 (N_11655,N_11467,N_11435);
or U11656 (N_11656,N_11532,N_11422);
nand U11657 (N_11657,N_11552,N_11409);
and U11658 (N_11658,N_11458,N_11402);
and U11659 (N_11659,N_11579,N_11498);
and U11660 (N_11660,N_11424,N_11548);
xnor U11661 (N_11661,N_11593,N_11550);
nor U11662 (N_11662,N_11597,N_11438);
xor U11663 (N_11663,N_11504,N_11476);
xor U11664 (N_11664,N_11565,N_11551);
xor U11665 (N_11665,N_11582,N_11477);
nand U11666 (N_11666,N_11568,N_11501);
or U11667 (N_11667,N_11431,N_11590);
nand U11668 (N_11668,N_11544,N_11490);
xor U11669 (N_11669,N_11487,N_11511);
xnor U11670 (N_11670,N_11510,N_11499);
and U11671 (N_11671,N_11447,N_11480);
xnor U11672 (N_11672,N_11520,N_11576);
nand U11673 (N_11673,N_11423,N_11471);
or U11674 (N_11674,N_11442,N_11482);
nor U11675 (N_11675,N_11558,N_11444);
and U11676 (N_11676,N_11488,N_11587);
nor U11677 (N_11677,N_11598,N_11483);
nor U11678 (N_11678,N_11481,N_11575);
xnor U11679 (N_11679,N_11529,N_11560);
xor U11680 (N_11680,N_11479,N_11474);
nor U11681 (N_11681,N_11493,N_11518);
xnor U11682 (N_11682,N_11454,N_11557);
and U11683 (N_11683,N_11484,N_11445);
nor U11684 (N_11684,N_11421,N_11564);
or U11685 (N_11685,N_11539,N_11408);
or U11686 (N_11686,N_11492,N_11509);
xor U11687 (N_11687,N_11542,N_11429);
or U11688 (N_11688,N_11439,N_11589);
nor U11689 (N_11689,N_11543,N_11448);
and U11690 (N_11690,N_11536,N_11411);
or U11691 (N_11691,N_11595,N_11416);
nor U11692 (N_11692,N_11441,N_11508);
nor U11693 (N_11693,N_11525,N_11466);
and U11694 (N_11694,N_11485,N_11452);
or U11695 (N_11695,N_11502,N_11533);
and U11696 (N_11696,N_11523,N_11554);
xnor U11697 (N_11697,N_11403,N_11457);
nor U11698 (N_11698,N_11578,N_11406);
nand U11699 (N_11699,N_11562,N_11413);
xnor U11700 (N_11700,N_11475,N_11417);
nor U11701 (N_11701,N_11488,N_11538);
xnor U11702 (N_11702,N_11476,N_11584);
nand U11703 (N_11703,N_11554,N_11529);
nor U11704 (N_11704,N_11404,N_11529);
nand U11705 (N_11705,N_11422,N_11478);
xor U11706 (N_11706,N_11407,N_11460);
or U11707 (N_11707,N_11547,N_11551);
nand U11708 (N_11708,N_11506,N_11458);
xor U11709 (N_11709,N_11532,N_11469);
xor U11710 (N_11710,N_11570,N_11589);
xor U11711 (N_11711,N_11576,N_11498);
or U11712 (N_11712,N_11537,N_11409);
nand U11713 (N_11713,N_11418,N_11426);
and U11714 (N_11714,N_11576,N_11596);
nand U11715 (N_11715,N_11510,N_11576);
and U11716 (N_11716,N_11482,N_11542);
nand U11717 (N_11717,N_11473,N_11534);
nor U11718 (N_11718,N_11556,N_11453);
and U11719 (N_11719,N_11477,N_11590);
xor U11720 (N_11720,N_11587,N_11577);
nand U11721 (N_11721,N_11442,N_11522);
nand U11722 (N_11722,N_11562,N_11410);
or U11723 (N_11723,N_11559,N_11497);
nand U11724 (N_11724,N_11591,N_11409);
nand U11725 (N_11725,N_11516,N_11492);
or U11726 (N_11726,N_11413,N_11515);
nor U11727 (N_11727,N_11520,N_11466);
nand U11728 (N_11728,N_11530,N_11555);
or U11729 (N_11729,N_11414,N_11591);
or U11730 (N_11730,N_11512,N_11465);
and U11731 (N_11731,N_11518,N_11434);
and U11732 (N_11732,N_11539,N_11564);
nor U11733 (N_11733,N_11480,N_11482);
nand U11734 (N_11734,N_11551,N_11474);
nand U11735 (N_11735,N_11562,N_11485);
or U11736 (N_11736,N_11524,N_11428);
xor U11737 (N_11737,N_11518,N_11598);
and U11738 (N_11738,N_11449,N_11469);
and U11739 (N_11739,N_11599,N_11430);
or U11740 (N_11740,N_11505,N_11485);
xor U11741 (N_11741,N_11426,N_11427);
xor U11742 (N_11742,N_11403,N_11537);
nor U11743 (N_11743,N_11574,N_11461);
and U11744 (N_11744,N_11456,N_11476);
xor U11745 (N_11745,N_11556,N_11426);
nor U11746 (N_11746,N_11555,N_11552);
xnor U11747 (N_11747,N_11548,N_11583);
or U11748 (N_11748,N_11483,N_11418);
or U11749 (N_11749,N_11581,N_11544);
or U11750 (N_11750,N_11449,N_11510);
nand U11751 (N_11751,N_11528,N_11451);
nand U11752 (N_11752,N_11508,N_11587);
nand U11753 (N_11753,N_11588,N_11458);
or U11754 (N_11754,N_11429,N_11576);
nand U11755 (N_11755,N_11428,N_11514);
nor U11756 (N_11756,N_11494,N_11450);
and U11757 (N_11757,N_11499,N_11477);
nor U11758 (N_11758,N_11452,N_11412);
xnor U11759 (N_11759,N_11458,N_11471);
nor U11760 (N_11760,N_11448,N_11584);
or U11761 (N_11761,N_11457,N_11587);
nand U11762 (N_11762,N_11587,N_11578);
nor U11763 (N_11763,N_11505,N_11466);
and U11764 (N_11764,N_11413,N_11469);
xnor U11765 (N_11765,N_11406,N_11531);
nor U11766 (N_11766,N_11516,N_11475);
and U11767 (N_11767,N_11432,N_11420);
or U11768 (N_11768,N_11476,N_11549);
and U11769 (N_11769,N_11546,N_11566);
nor U11770 (N_11770,N_11516,N_11452);
nor U11771 (N_11771,N_11462,N_11446);
and U11772 (N_11772,N_11438,N_11543);
nor U11773 (N_11773,N_11522,N_11574);
or U11774 (N_11774,N_11474,N_11425);
or U11775 (N_11775,N_11497,N_11504);
nand U11776 (N_11776,N_11476,N_11445);
nor U11777 (N_11777,N_11485,N_11523);
nand U11778 (N_11778,N_11560,N_11524);
nor U11779 (N_11779,N_11487,N_11437);
or U11780 (N_11780,N_11507,N_11556);
or U11781 (N_11781,N_11533,N_11591);
or U11782 (N_11782,N_11481,N_11411);
nand U11783 (N_11783,N_11504,N_11520);
nand U11784 (N_11784,N_11573,N_11454);
nand U11785 (N_11785,N_11574,N_11415);
xnor U11786 (N_11786,N_11511,N_11510);
nand U11787 (N_11787,N_11437,N_11545);
or U11788 (N_11788,N_11572,N_11548);
and U11789 (N_11789,N_11519,N_11564);
nor U11790 (N_11790,N_11410,N_11569);
and U11791 (N_11791,N_11514,N_11530);
or U11792 (N_11792,N_11477,N_11452);
nor U11793 (N_11793,N_11583,N_11449);
or U11794 (N_11794,N_11462,N_11430);
or U11795 (N_11795,N_11432,N_11477);
and U11796 (N_11796,N_11582,N_11507);
xnor U11797 (N_11797,N_11594,N_11513);
xor U11798 (N_11798,N_11510,N_11468);
nand U11799 (N_11799,N_11459,N_11556);
or U11800 (N_11800,N_11646,N_11681);
nand U11801 (N_11801,N_11758,N_11757);
xor U11802 (N_11802,N_11603,N_11718);
xnor U11803 (N_11803,N_11775,N_11694);
and U11804 (N_11804,N_11728,N_11722);
xnor U11805 (N_11805,N_11644,N_11675);
or U11806 (N_11806,N_11659,N_11645);
nor U11807 (N_11807,N_11684,N_11715);
nor U11808 (N_11808,N_11609,N_11739);
and U11809 (N_11809,N_11685,N_11772);
xor U11810 (N_11810,N_11601,N_11726);
or U11811 (N_11811,N_11776,N_11688);
or U11812 (N_11812,N_11752,N_11610);
and U11813 (N_11813,N_11614,N_11611);
or U11814 (N_11814,N_11764,N_11731);
or U11815 (N_11815,N_11689,N_11755);
and U11816 (N_11816,N_11773,N_11662);
nand U11817 (N_11817,N_11736,N_11703);
or U11818 (N_11818,N_11746,N_11637);
or U11819 (N_11819,N_11615,N_11635);
xnor U11820 (N_11820,N_11785,N_11784);
and U11821 (N_11821,N_11788,N_11676);
or U11822 (N_11822,N_11650,N_11799);
nor U11823 (N_11823,N_11741,N_11600);
nor U11824 (N_11824,N_11698,N_11619);
xnor U11825 (N_11825,N_11753,N_11744);
nor U11826 (N_11826,N_11767,N_11648);
and U11827 (N_11827,N_11727,N_11697);
xnor U11828 (N_11828,N_11692,N_11699);
xor U11829 (N_11829,N_11670,N_11702);
or U11830 (N_11830,N_11682,N_11751);
or U11831 (N_11831,N_11626,N_11605);
nor U11832 (N_11832,N_11707,N_11674);
nor U11833 (N_11833,N_11665,N_11745);
and U11834 (N_11834,N_11771,N_11763);
nand U11835 (N_11835,N_11721,N_11725);
nand U11836 (N_11836,N_11616,N_11770);
nand U11837 (N_11837,N_11747,N_11666);
or U11838 (N_11838,N_11663,N_11618);
nor U11839 (N_11839,N_11798,N_11716);
nand U11840 (N_11840,N_11769,N_11696);
nor U11841 (N_11841,N_11677,N_11717);
or U11842 (N_11842,N_11653,N_11733);
xor U11843 (N_11843,N_11797,N_11720);
and U11844 (N_11844,N_11651,N_11606);
or U11845 (N_11845,N_11679,N_11631);
nand U11846 (N_11846,N_11740,N_11749);
or U11847 (N_11847,N_11729,N_11660);
or U11848 (N_11848,N_11734,N_11690);
nor U11849 (N_11849,N_11780,N_11723);
nor U11850 (N_11850,N_11711,N_11641);
and U11851 (N_11851,N_11686,N_11623);
xnor U11852 (N_11852,N_11691,N_11743);
nand U11853 (N_11853,N_11713,N_11652);
nand U11854 (N_11854,N_11777,N_11640);
xnor U11855 (N_11855,N_11786,N_11622);
xor U11856 (N_11856,N_11656,N_11756);
xnor U11857 (N_11857,N_11657,N_11667);
nor U11858 (N_11858,N_11794,N_11709);
nor U11859 (N_11859,N_11658,N_11766);
xnor U11860 (N_11860,N_11649,N_11796);
nor U11861 (N_11861,N_11765,N_11760);
and U11862 (N_11862,N_11624,N_11693);
or U11863 (N_11863,N_11661,N_11732);
or U11864 (N_11864,N_11629,N_11712);
and U11865 (N_11865,N_11617,N_11748);
nor U11866 (N_11866,N_11664,N_11642);
or U11867 (N_11867,N_11672,N_11625);
and U11868 (N_11868,N_11639,N_11669);
xor U11869 (N_11869,N_11774,N_11778);
nand U11870 (N_11870,N_11759,N_11714);
nor U11871 (N_11871,N_11779,N_11654);
nor U11872 (N_11872,N_11792,N_11630);
or U11873 (N_11873,N_11706,N_11750);
and U11874 (N_11874,N_11724,N_11621);
nand U11875 (N_11875,N_11782,N_11613);
nand U11876 (N_11876,N_11655,N_11634);
or U11877 (N_11877,N_11608,N_11704);
xor U11878 (N_11878,N_11737,N_11668);
nand U11879 (N_11879,N_11627,N_11647);
nand U11880 (N_11880,N_11761,N_11793);
and U11881 (N_11881,N_11754,N_11628);
nor U11882 (N_11882,N_11708,N_11638);
xor U11883 (N_11883,N_11643,N_11710);
nand U11884 (N_11884,N_11671,N_11633);
or U11885 (N_11885,N_11673,N_11695);
and U11886 (N_11886,N_11632,N_11680);
xnor U11887 (N_11887,N_11701,N_11700);
xnor U11888 (N_11888,N_11607,N_11735);
or U11889 (N_11889,N_11683,N_11602);
or U11890 (N_11890,N_11738,N_11795);
and U11891 (N_11891,N_11612,N_11705);
or U11892 (N_11892,N_11604,N_11719);
and U11893 (N_11893,N_11620,N_11787);
xor U11894 (N_11894,N_11687,N_11790);
or U11895 (N_11895,N_11762,N_11742);
or U11896 (N_11896,N_11783,N_11678);
nor U11897 (N_11897,N_11730,N_11781);
and U11898 (N_11898,N_11789,N_11791);
or U11899 (N_11899,N_11636,N_11768);
or U11900 (N_11900,N_11604,N_11630);
nand U11901 (N_11901,N_11785,N_11744);
nand U11902 (N_11902,N_11757,N_11657);
xor U11903 (N_11903,N_11693,N_11774);
nand U11904 (N_11904,N_11658,N_11601);
or U11905 (N_11905,N_11604,N_11607);
xor U11906 (N_11906,N_11605,N_11752);
or U11907 (N_11907,N_11645,N_11712);
xor U11908 (N_11908,N_11676,N_11699);
or U11909 (N_11909,N_11735,N_11788);
nor U11910 (N_11910,N_11754,N_11698);
xnor U11911 (N_11911,N_11675,N_11734);
or U11912 (N_11912,N_11621,N_11731);
or U11913 (N_11913,N_11697,N_11748);
and U11914 (N_11914,N_11678,N_11671);
xnor U11915 (N_11915,N_11773,N_11718);
and U11916 (N_11916,N_11640,N_11683);
or U11917 (N_11917,N_11645,N_11713);
or U11918 (N_11918,N_11674,N_11754);
and U11919 (N_11919,N_11657,N_11728);
xnor U11920 (N_11920,N_11670,N_11619);
nor U11921 (N_11921,N_11711,N_11657);
xor U11922 (N_11922,N_11756,N_11637);
or U11923 (N_11923,N_11733,N_11649);
nand U11924 (N_11924,N_11733,N_11701);
nor U11925 (N_11925,N_11613,N_11706);
and U11926 (N_11926,N_11623,N_11708);
or U11927 (N_11927,N_11771,N_11656);
xnor U11928 (N_11928,N_11768,N_11692);
nand U11929 (N_11929,N_11616,N_11618);
nor U11930 (N_11930,N_11664,N_11614);
and U11931 (N_11931,N_11633,N_11751);
and U11932 (N_11932,N_11654,N_11608);
or U11933 (N_11933,N_11634,N_11712);
xor U11934 (N_11934,N_11737,N_11747);
nor U11935 (N_11935,N_11728,N_11772);
nand U11936 (N_11936,N_11615,N_11738);
or U11937 (N_11937,N_11675,N_11639);
or U11938 (N_11938,N_11662,N_11698);
or U11939 (N_11939,N_11756,N_11704);
or U11940 (N_11940,N_11786,N_11760);
xor U11941 (N_11941,N_11791,N_11770);
xor U11942 (N_11942,N_11622,N_11724);
or U11943 (N_11943,N_11706,N_11755);
nand U11944 (N_11944,N_11637,N_11699);
and U11945 (N_11945,N_11669,N_11649);
nand U11946 (N_11946,N_11676,N_11601);
or U11947 (N_11947,N_11627,N_11717);
and U11948 (N_11948,N_11795,N_11720);
or U11949 (N_11949,N_11724,N_11650);
nor U11950 (N_11950,N_11763,N_11698);
and U11951 (N_11951,N_11611,N_11732);
and U11952 (N_11952,N_11770,N_11785);
nor U11953 (N_11953,N_11734,N_11798);
xnor U11954 (N_11954,N_11622,N_11643);
nand U11955 (N_11955,N_11647,N_11628);
and U11956 (N_11956,N_11768,N_11735);
nor U11957 (N_11957,N_11726,N_11682);
xnor U11958 (N_11958,N_11642,N_11654);
or U11959 (N_11959,N_11710,N_11699);
or U11960 (N_11960,N_11720,N_11624);
xor U11961 (N_11961,N_11733,N_11788);
xnor U11962 (N_11962,N_11613,N_11675);
nand U11963 (N_11963,N_11684,N_11692);
nor U11964 (N_11964,N_11674,N_11688);
and U11965 (N_11965,N_11717,N_11794);
nor U11966 (N_11966,N_11780,N_11760);
or U11967 (N_11967,N_11783,N_11658);
and U11968 (N_11968,N_11735,N_11629);
or U11969 (N_11969,N_11741,N_11636);
and U11970 (N_11970,N_11624,N_11727);
nor U11971 (N_11971,N_11751,N_11686);
xnor U11972 (N_11972,N_11601,N_11760);
and U11973 (N_11973,N_11696,N_11641);
nand U11974 (N_11974,N_11650,N_11720);
and U11975 (N_11975,N_11787,N_11685);
nor U11976 (N_11976,N_11731,N_11637);
nor U11977 (N_11977,N_11703,N_11701);
xor U11978 (N_11978,N_11738,N_11709);
or U11979 (N_11979,N_11713,N_11675);
xor U11980 (N_11980,N_11790,N_11704);
or U11981 (N_11981,N_11789,N_11657);
xnor U11982 (N_11982,N_11633,N_11736);
nor U11983 (N_11983,N_11691,N_11687);
and U11984 (N_11984,N_11715,N_11623);
xnor U11985 (N_11985,N_11687,N_11783);
nor U11986 (N_11986,N_11734,N_11622);
or U11987 (N_11987,N_11682,N_11640);
nor U11988 (N_11988,N_11766,N_11613);
and U11989 (N_11989,N_11783,N_11674);
nand U11990 (N_11990,N_11772,N_11698);
or U11991 (N_11991,N_11615,N_11769);
nand U11992 (N_11992,N_11631,N_11605);
nand U11993 (N_11993,N_11736,N_11614);
and U11994 (N_11994,N_11611,N_11762);
nand U11995 (N_11995,N_11635,N_11764);
and U11996 (N_11996,N_11671,N_11714);
and U11997 (N_11997,N_11756,N_11723);
nor U11998 (N_11998,N_11661,N_11706);
nand U11999 (N_11999,N_11770,N_11676);
or U12000 (N_12000,N_11988,N_11871);
nand U12001 (N_12001,N_11893,N_11910);
xnor U12002 (N_12002,N_11925,N_11960);
or U12003 (N_12003,N_11905,N_11916);
or U12004 (N_12004,N_11898,N_11923);
or U12005 (N_12005,N_11825,N_11996);
and U12006 (N_12006,N_11877,N_11803);
nand U12007 (N_12007,N_11858,N_11814);
and U12008 (N_12008,N_11991,N_11878);
nor U12009 (N_12009,N_11849,N_11922);
or U12010 (N_12010,N_11833,N_11896);
nor U12011 (N_12011,N_11894,N_11897);
and U12012 (N_12012,N_11965,N_11911);
or U12013 (N_12013,N_11851,N_11845);
and U12014 (N_12014,N_11956,N_11993);
nand U12015 (N_12015,N_11826,N_11958);
nor U12016 (N_12016,N_11986,N_11946);
nand U12017 (N_12017,N_11954,N_11823);
nor U12018 (N_12018,N_11836,N_11942);
and U12019 (N_12019,N_11868,N_11970);
nor U12020 (N_12020,N_11839,N_11930);
nor U12021 (N_12021,N_11917,N_11907);
nor U12022 (N_12022,N_11857,N_11862);
nor U12023 (N_12023,N_11854,N_11926);
nand U12024 (N_12024,N_11998,N_11844);
nor U12025 (N_12025,N_11966,N_11805);
nand U12026 (N_12026,N_11846,N_11987);
or U12027 (N_12027,N_11948,N_11832);
or U12028 (N_12028,N_11829,N_11884);
xnor U12029 (N_12029,N_11962,N_11856);
nand U12030 (N_12030,N_11999,N_11891);
or U12031 (N_12031,N_11920,N_11974);
nand U12032 (N_12032,N_11850,N_11947);
and U12033 (N_12033,N_11941,N_11932);
nor U12034 (N_12034,N_11913,N_11906);
or U12035 (N_12035,N_11864,N_11853);
nand U12036 (N_12036,N_11837,N_11888);
nand U12037 (N_12037,N_11949,N_11890);
and U12038 (N_12038,N_11934,N_11938);
and U12039 (N_12039,N_11895,N_11872);
or U12040 (N_12040,N_11975,N_11881);
nor U12041 (N_12041,N_11819,N_11800);
xor U12042 (N_12042,N_11951,N_11978);
nand U12043 (N_12043,N_11903,N_11963);
and U12044 (N_12044,N_11852,N_11876);
xnor U12045 (N_12045,N_11924,N_11827);
xor U12046 (N_12046,N_11885,N_11801);
and U12047 (N_12047,N_11859,N_11883);
nor U12048 (N_12048,N_11813,N_11866);
nand U12049 (N_12049,N_11931,N_11967);
and U12050 (N_12050,N_11940,N_11919);
or U12051 (N_12051,N_11870,N_11935);
or U12052 (N_12052,N_11969,N_11972);
xor U12053 (N_12053,N_11808,N_11929);
and U12054 (N_12054,N_11955,N_11806);
nand U12055 (N_12055,N_11810,N_11992);
or U12056 (N_12056,N_11824,N_11882);
nand U12057 (N_12057,N_11889,N_11816);
and U12058 (N_12058,N_11840,N_11860);
nor U12059 (N_12059,N_11982,N_11815);
nor U12060 (N_12060,N_11995,N_11977);
and U12061 (N_12061,N_11964,N_11994);
and U12062 (N_12062,N_11887,N_11933);
nand U12063 (N_12063,N_11950,N_11980);
and U12064 (N_12064,N_11818,N_11820);
or U12065 (N_12065,N_11997,N_11812);
and U12066 (N_12066,N_11869,N_11847);
xnor U12067 (N_12067,N_11886,N_11959);
xor U12068 (N_12068,N_11880,N_11834);
or U12069 (N_12069,N_11953,N_11985);
xor U12070 (N_12070,N_11879,N_11838);
nand U12071 (N_12071,N_11873,N_11957);
or U12072 (N_12072,N_11981,N_11909);
or U12073 (N_12073,N_11900,N_11807);
xor U12074 (N_12074,N_11914,N_11908);
or U12075 (N_12075,N_11841,N_11835);
nand U12076 (N_12076,N_11915,N_11843);
xnor U12077 (N_12077,N_11968,N_11863);
nor U12078 (N_12078,N_11989,N_11848);
xnor U12079 (N_12079,N_11979,N_11984);
nand U12080 (N_12080,N_11927,N_11899);
and U12081 (N_12081,N_11828,N_11817);
nand U12082 (N_12082,N_11875,N_11821);
or U12083 (N_12083,N_11939,N_11961);
xnor U12084 (N_12084,N_11976,N_11830);
nor U12085 (N_12085,N_11944,N_11842);
nor U12086 (N_12086,N_11912,N_11943);
or U12087 (N_12087,N_11901,N_11867);
nand U12088 (N_12088,N_11861,N_11928);
xnor U12089 (N_12089,N_11855,N_11973);
xnor U12090 (N_12090,N_11952,N_11904);
and U12091 (N_12091,N_11921,N_11990);
or U12092 (N_12092,N_11983,N_11809);
xnor U12093 (N_12093,N_11802,N_11902);
nor U12094 (N_12094,N_11865,N_11811);
xor U12095 (N_12095,N_11831,N_11936);
and U12096 (N_12096,N_11892,N_11945);
nor U12097 (N_12097,N_11918,N_11822);
and U12098 (N_12098,N_11874,N_11971);
or U12099 (N_12099,N_11804,N_11937);
or U12100 (N_12100,N_11973,N_11928);
nor U12101 (N_12101,N_11807,N_11855);
or U12102 (N_12102,N_11935,N_11986);
and U12103 (N_12103,N_11829,N_11882);
and U12104 (N_12104,N_11923,N_11962);
or U12105 (N_12105,N_11873,N_11950);
xor U12106 (N_12106,N_11910,N_11935);
and U12107 (N_12107,N_11957,N_11847);
nor U12108 (N_12108,N_11892,N_11913);
or U12109 (N_12109,N_11950,N_11961);
nor U12110 (N_12110,N_11856,N_11910);
nand U12111 (N_12111,N_11809,N_11894);
nor U12112 (N_12112,N_11908,N_11809);
or U12113 (N_12113,N_11949,N_11925);
nand U12114 (N_12114,N_11859,N_11829);
and U12115 (N_12115,N_11893,N_11847);
nor U12116 (N_12116,N_11942,N_11894);
nor U12117 (N_12117,N_11818,N_11992);
or U12118 (N_12118,N_11833,N_11931);
nor U12119 (N_12119,N_11879,N_11857);
or U12120 (N_12120,N_11882,N_11952);
xor U12121 (N_12121,N_11912,N_11867);
nor U12122 (N_12122,N_11981,N_11831);
nand U12123 (N_12123,N_11822,N_11971);
nor U12124 (N_12124,N_11865,N_11905);
xor U12125 (N_12125,N_11925,N_11863);
xor U12126 (N_12126,N_11903,N_11982);
nand U12127 (N_12127,N_11882,N_11808);
nand U12128 (N_12128,N_11865,N_11916);
and U12129 (N_12129,N_11908,N_11880);
and U12130 (N_12130,N_11958,N_11804);
and U12131 (N_12131,N_11875,N_11838);
nand U12132 (N_12132,N_11839,N_11975);
nand U12133 (N_12133,N_11963,N_11977);
nand U12134 (N_12134,N_11957,N_11952);
or U12135 (N_12135,N_11909,N_11805);
nor U12136 (N_12136,N_11920,N_11845);
or U12137 (N_12137,N_11825,N_11939);
nand U12138 (N_12138,N_11851,N_11857);
xor U12139 (N_12139,N_11944,N_11954);
xor U12140 (N_12140,N_11942,N_11864);
xor U12141 (N_12141,N_11871,N_11922);
and U12142 (N_12142,N_11981,N_11976);
nand U12143 (N_12143,N_11837,N_11989);
or U12144 (N_12144,N_11941,N_11845);
nor U12145 (N_12145,N_11889,N_11819);
nor U12146 (N_12146,N_11913,N_11881);
nor U12147 (N_12147,N_11831,N_11963);
and U12148 (N_12148,N_11871,N_11991);
nand U12149 (N_12149,N_11861,N_11814);
or U12150 (N_12150,N_11841,N_11930);
or U12151 (N_12151,N_11965,N_11888);
nand U12152 (N_12152,N_11900,N_11907);
xnor U12153 (N_12153,N_11824,N_11978);
nand U12154 (N_12154,N_11817,N_11864);
and U12155 (N_12155,N_11911,N_11809);
nand U12156 (N_12156,N_11948,N_11926);
xnor U12157 (N_12157,N_11957,N_11811);
and U12158 (N_12158,N_11966,N_11961);
nand U12159 (N_12159,N_11938,N_11959);
or U12160 (N_12160,N_11835,N_11893);
and U12161 (N_12161,N_11952,N_11873);
nand U12162 (N_12162,N_11964,N_11985);
nor U12163 (N_12163,N_11942,N_11934);
and U12164 (N_12164,N_11854,N_11884);
and U12165 (N_12165,N_11892,N_11807);
or U12166 (N_12166,N_11834,N_11840);
nor U12167 (N_12167,N_11947,N_11881);
nor U12168 (N_12168,N_11982,N_11855);
or U12169 (N_12169,N_11979,N_11825);
and U12170 (N_12170,N_11847,N_11826);
and U12171 (N_12171,N_11967,N_11910);
xnor U12172 (N_12172,N_11822,N_11968);
nor U12173 (N_12173,N_11921,N_11950);
nand U12174 (N_12174,N_11873,N_11914);
nor U12175 (N_12175,N_11965,N_11845);
nor U12176 (N_12176,N_11851,N_11822);
nor U12177 (N_12177,N_11977,N_11931);
nor U12178 (N_12178,N_11881,N_11837);
nor U12179 (N_12179,N_11890,N_11818);
nor U12180 (N_12180,N_11982,N_11980);
or U12181 (N_12181,N_11851,N_11936);
xnor U12182 (N_12182,N_11882,N_11975);
nor U12183 (N_12183,N_11968,N_11894);
or U12184 (N_12184,N_11855,N_11899);
nand U12185 (N_12185,N_11981,N_11818);
nand U12186 (N_12186,N_11817,N_11938);
xor U12187 (N_12187,N_11801,N_11943);
and U12188 (N_12188,N_11818,N_11947);
nand U12189 (N_12189,N_11881,N_11826);
xnor U12190 (N_12190,N_11987,N_11913);
nor U12191 (N_12191,N_11851,N_11848);
nor U12192 (N_12192,N_11820,N_11869);
or U12193 (N_12193,N_11916,N_11988);
xor U12194 (N_12194,N_11969,N_11845);
nor U12195 (N_12195,N_11936,N_11803);
nor U12196 (N_12196,N_11866,N_11878);
xor U12197 (N_12197,N_11977,N_11819);
xor U12198 (N_12198,N_11967,N_11882);
nand U12199 (N_12199,N_11913,N_11865);
nand U12200 (N_12200,N_12029,N_12006);
or U12201 (N_12201,N_12026,N_12136);
xor U12202 (N_12202,N_12150,N_12014);
nand U12203 (N_12203,N_12028,N_12170);
nand U12204 (N_12204,N_12063,N_12194);
xnor U12205 (N_12205,N_12101,N_12093);
or U12206 (N_12206,N_12198,N_12178);
nand U12207 (N_12207,N_12095,N_12121);
nand U12208 (N_12208,N_12143,N_12187);
xnor U12209 (N_12209,N_12158,N_12127);
and U12210 (N_12210,N_12070,N_12097);
xor U12211 (N_12211,N_12122,N_12091);
nor U12212 (N_12212,N_12053,N_12061);
and U12213 (N_12213,N_12038,N_12140);
and U12214 (N_12214,N_12126,N_12075);
or U12215 (N_12215,N_12042,N_12106);
nor U12216 (N_12216,N_12002,N_12193);
and U12217 (N_12217,N_12087,N_12155);
or U12218 (N_12218,N_12066,N_12021);
xor U12219 (N_12219,N_12171,N_12147);
nand U12220 (N_12220,N_12092,N_12055);
xnor U12221 (N_12221,N_12031,N_12191);
xnor U12222 (N_12222,N_12088,N_12083);
xor U12223 (N_12223,N_12120,N_12012);
and U12224 (N_12224,N_12128,N_12197);
nand U12225 (N_12225,N_12144,N_12116);
nor U12226 (N_12226,N_12057,N_12084);
xor U12227 (N_12227,N_12033,N_12175);
nor U12228 (N_12228,N_12102,N_12130);
or U12229 (N_12229,N_12161,N_12051);
or U12230 (N_12230,N_12009,N_12184);
nor U12231 (N_12231,N_12050,N_12039);
nor U12232 (N_12232,N_12044,N_12085);
or U12233 (N_12233,N_12145,N_12196);
and U12234 (N_12234,N_12148,N_12164);
nor U12235 (N_12235,N_12156,N_12190);
xnor U12236 (N_12236,N_12181,N_12027);
xor U12237 (N_12237,N_12069,N_12142);
or U12238 (N_12238,N_12081,N_12049);
nor U12239 (N_12239,N_12054,N_12163);
xor U12240 (N_12240,N_12043,N_12005);
and U12241 (N_12241,N_12047,N_12108);
nor U12242 (N_12242,N_12098,N_12001);
or U12243 (N_12243,N_12172,N_12109);
xor U12244 (N_12244,N_12110,N_12169);
and U12245 (N_12245,N_12046,N_12105);
xnor U12246 (N_12246,N_12118,N_12176);
nand U12247 (N_12247,N_12183,N_12146);
nor U12248 (N_12248,N_12134,N_12072);
or U12249 (N_12249,N_12003,N_12064);
or U12250 (N_12250,N_12119,N_12182);
xor U12251 (N_12251,N_12167,N_12131);
nor U12252 (N_12252,N_12125,N_12137);
nand U12253 (N_12253,N_12168,N_12062);
nand U12254 (N_12254,N_12141,N_12112);
nor U12255 (N_12255,N_12133,N_12076);
or U12256 (N_12256,N_12123,N_12185);
nand U12257 (N_12257,N_12004,N_12041);
and U12258 (N_12258,N_12034,N_12199);
xnor U12259 (N_12259,N_12152,N_12025);
or U12260 (N_12260,N_12011,N_12179);
or U12261 (N_12261,N_12030,N_12013);
and U12262 (N_12262,N_12103,N_12099);
xor U12263 (N_12263,N_12078,N_12094);
nor U12264 (N_12264,N_12048,N_12177);
nand U12265 (N_12265,N_12149,N_12114);
and U12266 (N_12266,N_12139,N_12023);
or U12267 (N_12267,N_12086,N_12107);
nor U12268 (N_12268,N_12036,N_12159);
and U12269 (N_12269,N_12074,N_12037);
or U12270 (N_12270,N_12104,N_12067);
or U12271 (N_12271,N_12017,N_12060);
and U12272 (N_12272,N_12089,N_12059);
and U12273 (N_12273,N_12111,N_12068);
and U12274 (N_12274,N_12192,N_12022);
nor U12275 (N_12275,N_12115,N_12166);
xnor U12276 (N_12276,N_12073,N_12000);
nor U12277 (N_12277,N_12056,N_12151);
nand U12278 (N_12278,N_12065,N_12117);
or U12279 (N_12279,N_12165,N_12019);
and U12280 (N_12280,N_12100,N_12035);
nor U12281 (N_12281,N_12188,N_12132);
nand U12282 (N_12282,N_12160,N_12186);
or U12283 (N_12283,N_12154,N_12040);
or U12284 (N_12284,N_12082,N_12008);
and U12285 (N_12285,N_12016,N_12080);
xnor U12286 (N_12286,N_12135,N_12032);
and U12287 (N_12287,N_12157,N_12189);
xnor U12288 (N_12288,N_12058,N_12018);
xnor U12289 (N_12289,N_12153,N_12079);
or U12290 (N_12290,N_12173,N_12129);
and U12291 (N_12291,N_12195,N_12010);
and U12292 (N_12292,N_12174,N_12138);
or U12293 (N_12293,N_12090,N_12162);
xor U12294 (N_12294,N_12096,N_12113);
nand U12295 (N_12295,N_12071,N_12020);
nand U12296 (N_12296,N_12180,N_12052);
and U12297 (N_12297,N_12124,N_12007);
xnor U12298 (N_12298,N_12045,N_12024);
and U12299 (N_12299,N_12077,N_12015);
and U12300 (N_12300,N_12177,N_12127);
nand U12301 (N_12301,N_12113,N_12139);
or U12302 (N_12302,N_12062,N_12190);
xnor U12303 (N_12303,N_12180,N_12167);
nor U12304 (N_12304,N_12048,N_12040);
nor U12305 (N_12305,N_12086,N_12081);
nor U12306 (N_12306,N_12045,N_12008);
nand U12307 (N_12307,N_12036,N_12165);
nand U12308 (N_12308,N_12106,N_12101);
xor U12309 (N_12309,N_12089,N_12074);
xnor U12310 (N_12310,N_12119,N_12014);
nand U12311 (N_12311,N_12048,N_12108);
or U12312 (N_12312,N_12127,N_12055);
and U12313 (N_12313,N_12181,N_12186);
or U12314 (N_12314,N_12071,N_12103);
xor U12315 (N_12315,N_12072,N_12086);
xor U12316 (N_12316,N_12146,N_12048);
xnor U12317 (N_12317,N_12015,N_12126);
xor U12318 (N_12318,N_12136,N_12197);
and U12319 (N_12319,N_12087,N_12113);
xnor U12320 (N_12320,N_12185,N_12075);
or U12321 (N_12321,N_12169,N_12008);
xor U12322 (N_12322,N_12196,N_12126);
nor U12323 (N_12323,N_12183,N_12137);
nand U12324 (N_12324,N_12197,N_12082);
xor U12325 (N_12325,N_12153,N_12183);
or U12326 (N_12326,N_12099,N_12051);
nand U12327 (N_12327,N_12034,N_12141);
nor U12328 (N_12328,N_12079,N_12113);
or U12329 (N_12329,N_12012,N_12061);
xor U12330 (N_12330,N_12198,N_12125);
or U12331 (N_12331,N_12096,N_12160);
and U12332 (N_12332,N_12052,N_12088);
or U12333 (N_12333,N_12003,N_12177);
and U12334 (N_12334,N_12082,N_12032);
or U12335 (N_12335,N_12132,N_12070);
nand U12336 (N_12336,N_12096,N_12068);
xor U12337 (N_12337,N_12150,N_12046);
nor U12338 (N_12338,N_12133,N_12183);
or U12339 (N_12339,N_12002,N_12188);
and U12340 (N_12340,N_12101,N_12169);
or U12341 (N_12341,N_12133,N_12077);
nand U12342 (N_12342,N_12035,N_12199);
xor U12343 (N_12343,N_12167,N_12076);
and U12344 (N_12344,N_12048,N_12046);
or U12345 (N_12345,N_12172,N_12118);
xnor U12346 (N_12346,N_12027,N_12041);
nand U12347 (N_12347,N_12018,N_12057);
nor U12348 (N_12348,N_12115,N_12068);
or U12349 (N_12349,N_12048,N_12122);
xnor U12350 (N_12350,N_12191,N_12028);
nand U12351 (N_12351,N_12066,N_12006);
nor U12352 (N_12352,N_12126,N_12100);
xnor U12353 (N_12353,N_12081,N_12167);
nor U12354 (N_12354,N_12008,N_12121);
nor U12355 (N_12355,N_12063,N_12174);
xnor U12356 (N_12356,N_12184,N_12122);
and U12357 (N_12357,N_12172,N_12187);
nor U12358 (N_12358,N_12143,N_12099);
xnor U12359 (N_12359,N_12053,N_12117);
and U12360 (N_12360,N_12090,N_12059);
and U12361 (N_12361,N_12070,N_12034);
and U12362 (N_12362,N_12001,N_12166);
nand U12363 (N_12363,N_12151,N_12190);
nand U12364 (N_12364,N_12079,N_12020);
or U12365 (N_12365,N_12149,N_12046);
nor U12366 (N_12366,N_12001,N_12044);
or U12367 (N_12367,N_12106,N_12028);
or U12368 (N_12368,N_12138,N_12163);
and U12369 (N_12369,N_12075,N_12000);
nor U12370 (N_12370,N_12077,N_12116);
and U12371 (N_12371,N_12141,N_12074);
nor U12372 (N_12372,N_12126,N_12148);
and U12373 (N_12373,N_12052,N_12166);
or U12374 (N_12374,N_12139,N_12100);
xnor U12375 (N_12375,N_12011,N_12035);
nor U12376 (N_12376,N_12104,N_12040);
and U12377 (N_12377,N_12099,N_12122);
xor U12378 (N_12378,N_12110,N_12147);
nor U12379 (N_12379,N_12111,N_12084);
and U12380 (N_12380,N_12090,N_12030);
or U12381 (N_12381,N_12173,N_12113);
and U12382 (N_12382,N_12035,N_12020);
xor U12383 (N_12383,N_12015,N_12006);
and U12384 (N_12384,N_12134,N_12179);
xnor U12385 (N_12385,N_12115,N_12048);
nand U12386 (N_12386,N_12016,N_12024);
xnor U12387 (N_12387,N_12081,N_12069);
nand U12388 (N_12388,N_12171,N_12037);
xor U12389 (N_12389,N_12098,N_12109);
and U12390 (N_12390,N_12087,N_12166);
nand U12391 (N_12391,N_12171,N_12006);
and U12392 (N_12392,N_12198,N_12164);
nor U12393 (N_12393,N_12043,N_12073);
and U12394 (N_12394,N_12085,N_12139);
xor U12395 (N_12395,N_12111,N_12064);
xnor U12396 (N_12396,N_12198,N_12090);
and U12397 (N_12397,N_12069,N_12099);
or U12398 (N_12398,N_12111,N_12085);
xor U12399 (N_12399,N_12115,N_12054);
or U12400 (N_12400,N_12275,N_12293);
or U12401 (N_12401,N_12226,N_12212);
or U12402 (N_12402,N_12358,N_12354);
and U12403 (N_12403,N_12379,N_12357);
and U12404 (N_12404,N_12238,N_12376);
nor U12405 (N_12405,N_12322,N_12268);
xor U12406 (N_12406,N_12245,N_12292);
or U12407 (N_12407,N_12313,N_12205);
xnor U12408 (N_12408,N_12314,N_12204);
nand U12409 (N_12409,N_12237,N_12398);
nand U12410 (N_12410,N_12290,N_12342);
or U12411 (N_12411,N_12315,N_12251);
or U12412 (N_12412,N_12247,N_12224);
nor U12413 (N_12413,N_12249,N_12317);
xnor U12414 (N_12414,N_12375,N_12360);
and U12415 (N_12415,N_12340,N_12346);
and U12416 (N_12416,N_12272,N_12260);
nor U12417 (N_12417,N_12384,N_12300);
nand U12418 (N_12418,N_12284,N_12378);
nand U12419 (N_12419,N_12296,N_12389);
or U12420 (N_12420,N_12368,N_12264);
nand U12421 (N_12421,N_12230,N_12394);
and U12422 (N_12422,N_12312,N_12280);
nand U12423 (N_12423,N_12201,N_12220);
and U12424 (N_12424,N_12310,N_12203);
nor U12425 (N_12425,N_12323,N_12328);
and U12426 (N_12426,N_12246,N_12253);
nor U12427 (N_12427,N_12285,N_12288);
xor U12428 (N_12428,N_12202,N_12324);
nand U12429 (N_12429,N_12273,N_12343);
and U12430 (N_12430,N_12262,N_12271);
or U12431 (N_12431,N_12371,N_12303);
or U12432 (N_12432,N_12387,N_12355);
nor U12433 (N_12433,N_12261,N_12353);
nor U12434 (N_12434,N_12311,N_12337);
or U12435 (N_12435,N_12279,N_12321);
and U12436 (N_12436,N_12217,N_12373);
and U12437 (N_12437,N_12397,N_12374);
xor U12438 (N_12438,N_12367,N_12307);
xor U12439 (N_12439,N_12298,N_12242);
xnor U12440 (N_12440,N_12327,N_12221);
xnor U12441 (N_12441,N_12319,N_12350);
nand U12442 (N_12442,N_12277,N_12233);
or U12443 (N_12443,N_12255,N_12334);
and U12444 (N_12444,N_12396,N_12281);
nor U12445 (N_12445,N_12291,N_12309);
nor U12446 (N_12446,N_12382,N_12304);
nand U12447 (N_12447,N_12335,N_12339);
or U12448 (N_12448,N_12365,N_12287);
xor U12449 (N_12449,N_12208,N_12211);
nor U12450 (N_12450,N_12227,N_12235);
nand U12451 (N_12451,N_12200,N_12388);
nand U12452 (N_12452,N_12219,N_12370);
nand U12453 (N_12453,N_12206,N_12250);
xor U12454 (N_12454,N_12252,N_12270);
nor U12455 (N_12455,N_12278,N_12348);
nor U12456 (N_12456,N_12383,N_12331);
and U12457 (N_12457,N_12356,N_12305);
xor U12458 (N_12458,N_12257,N_12263);
xnor U12459 (N_12459,N_12240,N_12283);
nand U12460 (N_12460,N_12347,N_12229);
xor U12461 (N_12461,N_12381,N_12266);
or U12462 (N_12462,N_12359,N_12318);
nand U12463 (N_12463,N_12269,N_12294);
and U12464 (N_12464,N_12390,N_12223);
xnor U12465 (N_12465,N_12216,N_12385);
xnor U12466 (N_12466,N_12282,N_12380);
or U12467 (N_12467,N_12333,N_12295);
nor U12468 (N_12468,N_12215,N_12345);
xnor U12469 (N_12469,N_12301,N_12256);
and U12470 (N_12470,N_12344,N_12369);
nand U12471 (N_12471,N_12326,N_12391);
nand U12472 (N_12472,N_12248,N_12332);
nand U12473 (N_12473,N_12349,N_12210);
and U12474 (N_12474,N_12325,N_12393);
nand U12475 (N_12475,N_12209,N_12231);
or U12476 (N_12476,N_12276,N_12259);
and U12477 (N_12477,N_12267,N_12213);
nor U12478 (N_12478,N_12366,N_12218);
and U12479 (N_12479,N_12244,N_12232);
xnor U12480 (N_12480,N_12372,N_12399);
nor U12481 (N_12481,N_12308,N_12297);
nor U12482 (N_12482,N_12286,N_12302);
nor U12483 (N_12483,N_12274,N_12228);
nor U12484 (N_12484,N_12239,N_12364);
or U12485 (N_12485,N_12320,N_12386);
nor U12486 (N_12486,N_12362,N_12265);
and U12487 (N_12487,N_12351,N_12352);
xnor U12488 (N_12488,N_12241,N_12316);
or U12489 (N_12489,N_12330,N_12236);
nand U12490 (N_12490,N_12258,N_12254);
or U12491 (N_12491,N_12363,N_12222);
xor U12492 (N_12492,N_12214,N_12289);
or U12493 (N_12493,N_12336,N_12243);
and U12494 (N_12494,N_12234,N_12341);
and U12495 (N_12495,N_12377,N_12306);
nand U12496 (N_12496,N_12395,N_12207);
nand U12497 (N_12497,N_12361,N_12225);
or U12498 (N_12498,N_12338,N_12299);
nand U12499 (N_12499,N_12329,N_12392);
and U12500 (N_12500,N_12227,N_12388);
xnor U12501 (N_12501,N_12334,N_12327);
and U12502 (N_12502,N_12268,N_12206);
nand U12503 (N_12503,N_12308,N_12271);
nor U12504 (N_12504,N_12384,N_12216);
xnor U12505 (N_12505,N_12370,N_12286);
xnor U12506 (N_12506,N_12376,N_12284);
nor U12507 (N_12507,N_12203,N_12233);
or U12508 (N_12508,N_12359,N_12343);
nand U12509 (N_12509,N_12347,N_12220);
and U12510 (N_12510,N_12376,N_12210);
nand U12511 (N_12511,N_12360,N_12275);
nor U12512 (N_12512,N_12310,N_12214);
or U12513 (N_12513,N_12299,N_12383);
and U12514 (N_12514,N_12201,N_12327);
nor U12515 (N_12515,N_12286,N_12352);
nand U12516 (N_12516,N_12389,N_12263);
xnor U12517 (N_12517,N_12336,N_12277);
or U12518 (N_12518,N_12247,N_12336);
and U12519 (N_12519,N_12332,N_12215);
and U12520 (N_12520,N_12386,N_12372);
or U12521 (N_12521,N_12246,N_12273);
nor U12522 (N_12522,N_12220,N_12331);
and U12523 (N_12523,N_12347,N_12240);
nand U12524 (N_12524,N_12372,N_12390);
nor U12525 (N_12525,N_12263,N_12357);
nand U12526 (N_12526,N_12234,N_12356);
or U12527 (N_12527,N_12322,N_12328);
or U12528 (N_12528,N_12244,N_12308);
xor U12529 (N_12529,N_12217,N_12250);
xnor U12530 (N_12530,N_12345,N_12311);
and U12531 (N_12531,N_12225,N_12277);
nand U12532 (N_12532,N_12368,N_12206);
or U12533 (N_12533,N_12318,N_12297);
xor U12534 (N_12534,N_12338,N_12210);
and U12535 (N_12535,N_12365,N_12324);
nor U12536 (N_12536,N_12246,N_12283);
and U12537 (N_12537,N_12299,N_12337);
nor U12538 (N_12538,N_12365,N_12313);
and U12539 (N_12539,N_12395,N_12292);
nand U12540 (N_12540,N_12293,N_12351);
or U12541 (N_12541,N_12325,N_12355);
xnor U12542 (N_12542,N_12313,N_12210);
nor U12543 (N_12543,N_12235,N_12221);
nor U12544 (N_12544,N_12367,N_12393);
nand U12545 (N_12545,N_12384,N_12280);
or U12546 (N_12546,N_12300,N_12203);
nor U12547 (N_12547,N_12390,N_12200);
xor U12548 (N_12548,N_12266,N_12253);
nor U12549 (N_12549,N_12266,N_12307);
nand U12550 (N_12550,N_12212,N_12311);
xor U12551 (N_12551,N_12345,N_12359);
nor U12552 (N_12552,N_12207,N_12235);
nor U12553 (N_12553,N_12217,N_12265);
nand U12554 (N_12554,N_12216,N_12367);
nand U12555 (N_12555,N_12334,N_12375);
and U12556 (N_12556,N_12327,N_12232);
xnor U12557 (N_12557,N_12251,N_12323);
or U12558 (N_12558,N_12247,N_12380);
and U12559 (N_12559,N_12310,N_12227);
and U12560 (N_12560,N_12302,N_12210);
xnor U12561 (N_12561,N_12222,N_12307);
nand U12562 (N_12562,N_12339,N_12360);
and U12563 (N_12563,N_12345,N_12224);
and U12564 (N_12564,N_12219,N_12232);
xor U12565 (N_12565,N_12204,N_12313);
and U12566 (N_12566,N_12207,N_12242);
and U12567 (N_12567,N_12347,N_12314);
nor U12568 (N_12568,N_12362,N_12268);
or U12569 (N_12569,N_12311,N_12388);
nand U12570 (N_12570,N_12371,N_12360);
nor U12571 (N_12571,N_12245,N_12249);
nand U12572 (N_12572,N_12385,N_12379);
xnor U12573 (N_12573,N_12369,N_12262);
nor U12574 (N_12574,N_12389,N_12210);
xor U12575 (N_12575,N_12212,N_12350);
nor U12576 (N_12576,N_12316,N_12235);
and U12577 (N_12577,N_12317,N_12305);
and U12578 (N_12578,N_12220,N_12319);
or U12579 (N_12579,N_12275,N_12387);
and U12580 (N_12580,N_12276,N_12327);
nor U12581 (N_12581,N_12254,N_12211);
and U12582 (N_12582,N_12381,N_12324);
xnor U12583 (N_12583,N_12334,N_12246);
and U12584 (N_12584,N_12355,N_12385);
and U12585 (N_12585,N_12309,N_12326);
nand U12586 (N_12586,N_12394,N_12318);
and U12587 (N_12587,N_12269,N_12206);
nor U12588 (N_12588,N_12220,N_12324);
nor U12589 (N_12589,N_12257,N_12330);
nand U12590 (N_12590,N_12318,N_12378);
or U12591 (N_12591,N_12319,N_12223);
nand U12592 (N_12592,N_12243,N_12372);
xor U12593 (N_12593,N_12346,N_12274);
nand U12594 (N_12594,N_12370,N_12258);
nand U12595 (N_12595,N_12271,N_12206);
and U12596 (N_12596,N_12325,N_12319);
and U12597 (N_12597,N_12332,N_12390);
nor U12598 (N_12598,N_12348,N_12235);
or U12599 (N_12599,N_12291,N_12214);
or U12600 (N_12600,N_12464,N_12499);
and U12601 (N_12601,N_12527,N_12562);
xnor U12602 (N_12602,N_12439,N_12437);
or U12603 (N_12603,N_12448,N_12554);
nor U12604 (N_12604,N_12461,N_12539);
nand U12605 (N_12605,N_12570,N_12419);
nand U12606 (N_12606,N_12548,N_12444);
nor U12607 (N_12607,N_12434,N_12447);
nand U12608 (N_12608,N_12458,N_12535);
xnor U12609 (N_12609,N_12495,N_12586);
nand U12610 (N_12610,N_12431,N_12463);
nor U12611 (N_12611,N_12582,N_12485);
nand U12612 (N_12612,N_12416,N_12509);
and U12613 (N_12613,N_12438,N_12471);
and U12614 (N_12614,N_12467,N_12454);
or U12615 (N_12615,N_12445,N_12481);
and U12616 (N_12616,N_12493,N_12417);
xnor U12617 (N_12617,N_12522,N_12580);
xor U12618 (N_12618,N_12560,N_12558);
nand U12619 (N_12619,N_12488,N_12414);
or U12620 (N_12620,N_12534,N_12477);
nor U12621 (N_12621,N_12520,N_12588);
xnor U12622 (N_12622,N_12556,N_12486);
xor U12623 (N_12623,N_12430,N_12567);
nor U12624 (N_12624,N_12489,N_12440);
nor U12625 (N_12625,N_12551,N_12446);
nand U12626 (N_12626,N_12421,N_12429);
xor U12627 (N_12627,N_12422,N_12427);
or U12628 (N_12628,N_12571,N_12468);
nand U12629 (N_12629,N_12521,N_12479);
nand U12630 (N_12630,N_12566,N_12546);
and U12631 (N_12631,N_12497,N_12553);
or U12632 (N_12632,N_12518,N_12443);
or U12633 (N_12633,N_12504,N_12523);
and U12634 (N_12634,N_12537,N_12483);
and U12635 (N_12635,N_12524,N_12418);
nor U12636 (N_12636,N_12519,N_12474);
xor U12637 (N_12637,N_12457,N_12424);
and U12638 (N_12638,N_12589,N_12460);
and U12639 (N_12639,N_12576,N_12583);
nor U12640 (N_12640,N_12587,N_12591);
or U12641 (N_12641,N_12478,N_12402);
or U12642 (N_12642,N_12544,N_12406);
nand U12643 (N_12643,N_12572,N_12547);
nand U12644 (N_12644,N_12415,N_12574);
nand U12645 (N_12645,N_12484,N_12436);
xor U12646 (N_12646,N_12473,N_12491);
nor U12647 (N_12647,N_12404,N_12581);
xnor U12648 (N_12648,N_12536,N_12510);
nand U12649 (N_12649,N_12585,N_12578);
nor U12650 (N_12650,N_12528,N_12412);
nand U12651 (N_12651,N_12472,N_12592);
and U12652 (N_12652,N_12595,N_12487);
nand U12653 (N_12653,N_12450,N_12531);
or U12654 (N_12654,N_12449,N_12514);
or U12655 (N_12655,N_12452,N_12530);
or U12656 (N_12656,N_12584,N_12405);
nor U12657 (N_12657,N_12507,N_12563);
xor U12658 (N_12658,N_12469,N_12453);
or U12659 (N_12659,N_12573,N_12515);
nand U12660 (N_12660,N_12423,N_12525);
and U12661 (N_12661,N_12517,N_12596);
xor U12662 (N_12662,N_12492,N_12513);
nor U12663 (N_12663,N_12408,N_12549);
nand U12664 (N_12664,N_12568,N_12409);
nor U12665 (N_12665,N_12425,N_12475);
nand U12666 (N_12666,N_12506,N_12482);
xor U12667 (N_12667,N_12456,N_12532);
or U12668 (N_12668,N_12411,N_12413);
and U12669 (N_12669,N_12503,N_12593);
or U12670 (N_12670,N_12500,N_12401);
xor U12671 (N_12671,N_12579,N_12505);
nand U12672 (N_12672,N_12526,N_12542);
nor U12673 (N_12673,N_12543,N_12462);
and U12674 (N_12674,N_12564,N_12541);
xnor U12675 (N_12675,N_12470,N_12594);
xor U12676 (N_12676,N_12590,N_12433);
xor U12677 (N_12677,N_12565,N_12435);
and U12678 (N_12678,N_12480,N_12529);
and U12679 (N_12679,N_12569,N_12599);
and U12680 (N_12680,N_12575,N_12538);
nor U12681 (N_12681,N_12451,N_12400);
or U12682 (N_12682,N_12459,N_12512);
xnor U12683 (N_12683,N_12597,N_12540);
nand U12684 (N_12684,N_12494,N_12426);
and U12685 (N_12685,N_12559,N_12502);
xnor U12686 (N_12686,N_12441,N_12557);
xnor U12687 (N_12687,N_12516,N_12498);
and U12688 (N_12688,N_12555,N_12432);
nand U12689 (N_12689,N_12407,N_12577);
and U12690 (N_12690,N_12465,N_12496);
and U12691 (N_12691,N_12403,N_12476);
or U12692 (N_12692,N_12466,N_12442);
nand U12693 (N_12693,N_12550,N_12533);
xor U12694 (N_12694,N_12428,N_12598);
nor U12695 (N_12695,N_12545,N_12552);
xor U12696 (N_12696,N_12508,N_12490);
nand U12697 (N_12697,N_12420,N_12561);
or U12698 (N_12698,N_12410,N_12455);
nand U12699 (N_12699,N_12501,N_12511);
nor U12700 (N_12700,N_12526,N_12476);
and U12701 (N_12701,N_12580,N_12458);
nand U12702 (N_12702,N_12522,N_12442);
and U12703 (N_12703,N_12433,N_12400);
and U12704 (N_12704,N_12460,N_12503);
xor U12705 (N_12705,N_12535,N_12541);
xnor U12706 (N_12706,N_12477,N_12435);
and U12707 (N_12707,N_12500,N_12568);
or U12708 (N_12708,N_12516,N_12556);
xor U12709 (N_12709,N_12455,N_12424);
or U12710 (N_12710,N_12451,N_12503);
xnor U12711 (N_12711,N_12466,N_12494);
nand U12712 (N_12712,N_12516,N_12512);
nand U12713 (N_12713,N_12558,N_12457);
nor U12714 (N_12714,N_12474,N_12445);
or U12715 (N_12715,N_12418,N_12478);
nor U12716 (N_12716,N_12594,N_12467);
xor U12717 (N_12717,N_12471,N_12522);
or U12718 (N_12718,N_12561,N_12583);
nand U12719 (N_12719,N_12525,N_12414);
nand U12720 (N_12720,N_12465,N_12590);
or U12721 (N_12721,N_12403,N_12479);
xor U12722 (N_12722,N_12479,N_12574);
or U12723 (N_12723,N_12431,N_12513);
or U12724 (N_12724,N_12467,N_12478);
nor U12725 (N_12725,N_12594,N_12581);
and U12726 (N_12726,N_12517,N_12519);
nand U12727 (N_12727,N_12553,N_12556);
xor U12728 (N_12728,N_12469,N_12448);
and U12729 (N_12729,N_12505,N_12443);
or U12730 (N_12730,N_12563,N_12548);
nand U12731 (N_12731,N_12431,N_12407);
nand U12732 (N_12732,N_12431,N_12543);
nand U12733 (N_12733,N_12537,N_12546);
or U12734 (N_12734,N_12513,N_12595);
or U12735 (N_12735,N_12569,N_12473);
xnor U12736 (N_12736,N_12568,N_12495);
nor U12737 (N_12737,N_12514,N_12407);
or U12738 (N_12738,N_12545,N_12513);
nor U12739 (N_12739,N_12552,N_12591);
nand U12740 (N_12740,N_12570,N_12496);
nand U12741 (N_12741,N_12409,N_12595);
nor U12742 (N_12742,N_12585,N_12506);
nor U12743 (N_12743,N_12411,N_12404);
or U12744 (N_12744,N_12412,N_12489);
nor U12745 (N_12745,N_12438,N_12547);
and U12746 (N_12746,N_12506,N_12492);
xnor U12747 (N_12747,N_12555,N_12582);
nand U12748 (N_12748,N_12562,N_12530);
xnor U12749 (N_12749,N_12469,N_12444);
or U12750 (N_12750,N_12447,N_12558);
or U12751 (N_12751,N_12491,N_12518);
and U12752 (N_12752,N_12431,N_12514);
or U12753 (N_12753,N_12454,N_12459);
and U12754 (N_12754,N_12476,N_12528);
or U12755 (N_12755,N_12555,N_12406);
or U12756 (N_12756,N_12551,N_12495);
nor U12757 (N_12757,N_12468,N_12551);
or U12758 (N_12758,N_12562,N_12445);
nor U12759 (N_12759,N_12560,N_12568);
nand U12760 (N_12760,N_12520,N_12573);
xnor U12761 (N_12761,N_12499,N_12576);
and U12762 (N_12762,N_12429,N_12406);
or U12763 (N_12763,N_12572,N_12504);
or U12764 (N_12764,N_12579,N_12566);
or U12765 (N_12765,N_12474,N_12529);
nor U12766 (N_12766,N_12552,N_12471);
and U12767 (N_12767,N_12466,N_12552);
xor U12768 (N_12768,N_12559,N_12481);
or U12769 (N_12769,N_12426,N_12550);
xor U12770 (N_12770,N_12485,N_12510);
or U12771 (N_12771,N_12500,N_12444);
nand U12772 (N_12772,N_12580,N_12404);
xnor U12773 (N_12773,N_12511,N_12571);
nand U12774 (N_12774,N_12488,N_12557);
nand U12775 (N_12775,N_12484,N_12586);
or U12776 (N_12776,N_12460,N_12411);
or U12777 (N_12777,N_12591,N_12401);
nand U12778 (N_12778,N_12408,N_12588);
nor U12779 (N_12779,N_12560,N_12504);
or U12780 (N_12780,N_12575,N_12470);
nor U12781 (N_12781,N_12482,N_12429);
xor U12782 (N_12782,N_12511,N_12534);
and U12783 (N_12783,N_12534,N_12551);
and U12784 (N_12784,N_12521,N_12504);
nand U12785 (N_12785,N_12415,N_12584);
xor U12786 (N_12786,N_12429,N_12413);
xor U12787 (N_12787,N_12530,N_12509);
or U12788 (N_12788,N_12491,N_12500);
and U12789 (N_12789,N_12489,N_12488);
or U12790 (N_12790,N_12544,N_12501);
nand U12791 (N_12791,N_12589,N_12472);
and U12792 (N_12792,N_12576,N_12504);
and U12793 (N_12793,N_12529,N_12434);
and U12794 (N_12794,N_12415,N_12409);
nand U12795 (N_12795,N_12450,N_12456);
and U12796 (N_12796,N_12445,N_12421);
xor U12797 (N_12797,N_12489,N_12459);
xnor U12798 (N_12798,N_12415,N_12568);
or U12799 (N_12799,N_12447,N_12455);
xnor U12800 (N_12800,N_12604,N_12795);
or U12801 (N_12801,N_12669,N_12602);
and U12802 (N_12802,N_12799,N_12684);
xnor U12803 (N_12803,N_12739,N_12665);
xor U12804 (N_12804,N_12760,N_12693);
and U12805 (N_12805,N_12759,N_12623);
xnor U12806 (N_12806,N_12630,N_12612);
xnor U12807 (N_12807,N_12708,N_12656);
xor U12808 (N_12808,N_12711,N_12709);
or U12809 (N_12809,N_12747,N_12668);
nor U12810 (N_12810,N_12672,N_12779);
nand U12811 (N_12811,N_12676,N_12621);
or U12812 (N_12812,N_12620,N_12784);
xor U12813 (N_12813,N_12696,N_12666);
nor U12814 (N_12814,N_12679,N_12717);
xor U12815 (N_12815,N_12750,N_12689);
nor U12816 (N_12816,N_12682,N_12671);
or U12817 (N_12817,N_12798,N_12628);
xor U12818 (N_12818,N_12748,N_12707);
nand U12819 (N_12819,N_12730,N_12677);
xnor U12820 (N_12820,N_12715,N_12720);
xnor U12821 (N_12821,N_12685,N_12613);
xor U12822 (N_12822,N_12662,N_12757);
nand U12823 (N_12823,N_12751,N_12772);
or U12824 (N_12824,N_12673,N_12758);
nor U12825 (N_12825,N_12789,N_12649);
and U12826 (N_12826,N_12605,N_12729);
or U12827 (N_12827,N_12703,N_12773);
xor U12828 (N_12828,N_12632,N_12695);
xnor U12829 (N_12829,N_12624,N_12634);
nand U12830 (N_12830,N_12701,N_12744);
and U12831 (N_12831,N_12608,N_12713);
and U12832 (N_12832,N_12640,N_12636);
and U12833 (N_12833,N_12650,N_12768);
nand U12834 (N_12834,N_12734,N_12790);
nand U12835 (N_12835,N_12737,N_12704);
or U12836 (N_12836,N_12647,N_12675);
nor U12837 (N_12837,N_12626,N_12687);
or U12838 (N_12838,N_12638,N_12721);
and U12839 (N_12839,N_12637,N_12606);
and U12840 (N_12840,N_12719,N_12654);
and U12841 (N_12841,N_12770,N_12766);
and U12842 (N_12842,N_12791,N_12627);
xnor U12843 (N_12843,N_12635,N_12651);
or U12844 (N_12844,N_12752,N_12670);
or U12845 (N_12845,N_12722,N_12769);
or U12846 (N_12846,N_12680,N_12658);
nor U12847 (N_12847,N_12746,N_12653);
xnor U12848 (N_12848,N_12686,N_12776);
xor U12849 (N_12849,N_12607,N_12774);
xnor U12850 (N_12850,N_12712,N_12629);
nor U12851 (N_12851,N_12780,N_12716);
xor U12852 (N_12852,N_12648,N_12700);
nor U12853 (N_12853,N_12782,N_12681);
xor U12854 (N_12854,N_12783,N_12764);
xnor U12855 (N_12855,N_12688,N_12792);
xor U12856 (N_12856,N_12663,N_12775);
or U12857 (N_12857,N_12692,N_12778);
and U12858 (N_12858,N_12786,N_12618);
xor U12859 (N_12859,N_12615,N_12777);
nor U12860 (N_12860,N_12690,N_12705);
xnor U12861 (N_12861,N_12697,N_12740);
or U12862 (N_12862,N_12762,N_12781);
or U12863 (N_12863,N_12657,N_12702);
and U12864 (N_12864,N_12736,N_12754);
and U12865 (N_12865,N_12753,N_12797);
or U12866 (N_12866,N_12699,N_12787);
xor U12867 (N_12867,N_12742,N_12639);
or U12868 (N_12868,N_12643,N_12725);
and U12869 (N_12869,N_12645,N_12710);
nand U12870 (N_12870,N_12706,N_12714);
xor U12871 (N_12871,N_12659,N_12771);
and U12872 (N_12872,N_12611,N_12794);
xnor U12873 (N_12873,N_12755,N_12732);
and U12874 (N_12874,N_12655,N_12785);
or U12875 (N_12875,N_12633,N_12625);
and U12876 (N_12876,N_12619,N_12661);
nand U12877 (N_12877,N_12761,N_12728);
and U12878 (N_12878,N_12631,N_12641);
nand U12879 (N_12879,N_12745,N_12601);
nor U12880 (N_12880,N_12660,N_12735);
xnor U12881 (N_12881,N_12622,N_12765);
nand U12882 (N_12882,N_12642,N_12616);
nor U12883 (N_12883,N_12756,N_12646);
nand U12884 (N_12884,N_12749,N_12698);
nand U12885 (N_12885,N_12678,N_12683);
nor U12886 (N_12886,N_12600,N_12727);
xor U12887 (N_12887,N_12733,N_12652);
or U12888 (N_12888,N_12788,N_12723);
xor U12889 (N_12889,N_12767,N_12617);
or U12890 (N_12890,N_12603,N_12793);
and U12891 (N_12891,N_12724,N_12796);
and U12892 (N_12892,N_12763,N_12667);
xor U12893 (N_12893,N_12694,N_12743);
xnor U12894 (N_12894,N_12614,N_12609);
nand U12895 (N_12895,N_12610,N_12664);
nor U12896 (N_12896,N_12674,N_12738);
xor U12897 (N_12897,N_12718,N_12741);
and U12898 (N_12898,N_12644,N_12691);
xnor U12899 (N_12899,N_12726,N_12731);
or U12900 (N_12900,N_12636,N_12629);
and U12901 (N_12901,N_12612,N_12786);
xnor U12902 (N_12902,N_12784,N_12655);
and U12903 (N_12903,N_12611,N_12786);
nor U12904 (N_12904,N_12760,N_12646);
nor U12905 (N_12905,N_12688,N_12693);
nor U12906 (N_12906,N_12701,N_12623);
nor U12907 (N_12907,N_12789,N_12707);
and U12908 (N_12908,N_12663,N_12758);
xor U12909 (N_12909,N_12688,N_12774);
or U12910 (N_12910,N_12783,N_12745);
or U12911 (N_12911,N_12647,N_12751);
nor U12912 (N_12912,N_12729,N_12751);
nor U12913 (N_12913,N_12720,N_12747);
nand U12914 (N_12914,N_12730,N_12607);
and U12915 (N_12915,N_12715,N_12696);
or U12916 (N_12916,N_12745,N_12635);
nor U12917 (N_12917,N_12658,N_12626);
or U12918 (N_12918,N_12617,N_12728);
and U12919 (N_12919,N_12748,N_12720);
xnor U12920 (N_12920,N_12633,N_12643);
xnor U12921 (N_12921,N_12646,N_12633);
or U12922 (N_12922,N_12748,N_12614);
or U12923 (N_12923,N_12787,N_12767);
nand U12924 (N_12924,N_12784,N_12678);
or U12925 (N_12925,N_12697,N_12757);
or U12926 (N_12926,N_12747,N_12762);
nor U12927 (N_12927,N_12753,N_12694);
nand U12928 (N_12928,N_12632,N_12764);
and U12929 (N_12929,N_12638,N_12796);
or U12930 (N_12930,N_12705,N_12767);
or U12931 (N_12931,N_12707,N_12644);
nor U12932 (N_12932,N_12794,N_12705);
xnor U12933 (N_12933,N_12656,N_12632);
and U12934 (N_12934,N_12745,N_12625);
xnor U12935 (N_12935,N_12720,N_12633);
and U12936 (N_12936,N_12630,N_12750);
nor U12937 (N_12937,N_12784,N_12731);
and U12938 (N_12938,N_12652,N_12730);
xnor U12939 (N_12939,N_12797,N_12641);
xor U12940 (N_12940,N_12754,N_12772);
xnor U12941 (N_12941,N_12620,N_12654);
or U12942 (N_12942,N_12775,N_12665);
or U12943 (N_12943,N_12647,N_12790);
and U12944 (N_12944,N_12644,N_12717);
nor U12945 (N_12945,N_12767,N_12667);
and U12946 (N_12946,N_12733,N_12724);
and U12947 (N_12947,N_12779,N_12645);
nand U12948 (N_12948,N_12681,N_12724);
or U12949 (N_12949,N_12704,N_12666);
and U12950 (N_12950,N_12706,N_12617);
xor U12951 (N_12951,N_12737,N_12608);
xor U12952 (N_12952,N_12737,N_12741);
nand U12953 (N_12953,N_12654,N_12674);
nor U12954 (N_12954,N_12638,N_12693);
nor U12955 (N_12955,N_12731,N_12663);
nor U12956 (N_12956,N_12695,N_12778);
nor U12957 (N_12957,N_12698,N_12738);
or U12958 (N_12958,N_12727,N_12799);
nand U12959 (N_12959,N_12615,N_12719);
xnor U12960 (N_12960,N_12608,N_12795);
or U12961 (N_12961,N_12687,N_12722);
and U12962 (N_12962,N_12754,N_12624);
nor U12963 (N_12963,N_12774,N_12685);
and U12964 (N_12964,N_12653,N_12777);
nand U12965 (N_12965,N_12679,N_12609);
xor U12966 (N_12966,N_12639,N_12783);
and U12967 (N_12967,N_12679,N_12726);
and U12968 (N_12968,N_12699,N_12666);
and U12969 (N_12969,N_12757,N_12604);
nor U12970 (N_12970,N_12781,N_12603);
nand U12971 (N_12971,N_12787,N_12770);
and U12972 (N_12972,N_12640,N_12733);
nand U12973 (N_12973,N_12702,N_12716);
nand U12974 (N_12974,N_12706,N_12774);
xnor U12975 (N_12975,N_12759,N_12682);
or U12976 (N_12976,N_12682,N_12605);
and U12977 (N_12977,N_12664,N_12604);
nor U12978 (N_12978,N_12644,N_12642);
or U12979 (N_12979,N_12641,N_12698);
or U12980 (N_12980,N_12657,N_12688);
or U12981 (N_12981,N_12725,N_12635);
nor U12982 (N_12982,N_12759,N_12776);
nor U12983 (N_12983,N_12748,N_12787);
nor U12984 (N_12984,N_12784,N_12660);
nor U12985 (N_12985,N_12710,N_12607);
nand U12986 (N_12986,N_12639,N_12752);
and U12987 (N_12987,N_12738,N_12704);
nand U12988 (N_12988,N_12772,N_12709);
or U12989 (N_12989,N_12789,N_12724);
and U12990 (N_12990,N_12734,N_12798);
nand U12991 (N_12991,N_12623,N_12680);
nand U12992 (N_12992,N_12683,N_12659);
and U12993 (N_12993,N_12732,N_12680);
nand U12994 (N_12994,N_12784,N_12600);
and U12995 (N_12995,N_12697,N_12730);
or U12996 (N_12996,N_12705,N_12743);
or U12997 (N_12997,N_12789,N_12741);
or U12998 (N_12998,N_12721,N_12782);
nand U12999 (N_12999,N_12616,N_12671);
nand U13000 (N_13000,N_12869,N_12965);
or U13001 (N_13001,N_12881,N_12818);
nand U13002 (N_13002,N_12887,N_12944);
nand U13003 (N_13003,N_12937,N_12824);
and U13004 (N_13004,N_12963,N_12921);
or U13005 (N_13005,N_12907,N_12968);
nand U13006 (N_13006,N_12977,N_12952);
xor U13007 (N_13007,N_12916,N_12863);
nor U13008 (N_13008,N_12940,N_12846);
and U13009 (N_13009,N_12800,N_12919);
nand U13010 (N_13010,N_12867,N_12872);
nor U13011 (N_13011,N_12813,N_12918);
xnor U13012 (N_13012,N_12949,N_12882);
nand U13013 (N_13013,N_12982,N_12957);
and U13014 (N_13014,N_12900,N_12870);
and U13015 (N_13015,N_12904,N_12898);
nor U13016 (N_13016,N_12874,N_12983);
nand U13017 (N_13017,N_12849,N_12980);
nand U13018 (N_13018,N_12899,N_12978);
or U13019 (N_13019,N_12886,N_12981);
or U13020 (N_13020,N_12804,N_12941);
nor U13021 (N_13021,N_12821,N_12976);
nor U13022 (N_13022,N_12820,N_12806);
nor U13023 (N_13023,N_12987,N_12969);
xnor U13024 (N_13024,N_12997,N_12855);
and U13025 (N_13025,N_12905,N_12845);
xnor U13026 (N_13026,N_12842,N_12923);
or U13027 (N_13027,N_12827,N_12888);
and U13028 (N_13028,N_12920,N_12972);
nand U13029 (N_13029,N_12840,N_12892);
xnor U13030 (N_13030,N_12832,N_12971);
nor U13031 (N_13031,N_12954,N_12803);
or U13032 (N_13032,N_12950,N_12823);
or U13033 (N_13033,N_12808,N_12841);
and U13034 (N_13034,N_12868,N_12939);
or U13035 (N_13035,N_12903,N_12837);
and U13036 (N_13036,N_12848,N_12805);
xor U13037 (N_13037,N_12967,N_12883);
and U13038 (N_13038,N_12909,N_12975);
nor U13039 (N_13039,N_12876,N_12864);
nor U13040 (N_13040,N_12984,N_12853);
nand U13041 (N_13041,N_12973,N_12917);
or U13042 (N_13042,N_12829,N_12850);
nor U13043 (N_13043,N_12955,N_12964);
nand U13044 (N_13044,N_12956,N_12810);
xor U13045 (N_13045,N_12906,N_12947);
nand U13046 (N_13046,N_12946,N_12854);
and U13047 (N_13047,N_12988,N_12930);
nand U13048 (N_13048,N_12807,N_12960);
nand U13049 (N_13049,N_12833,N_12951);
and U13050 (N_13050,N_12902,N_12861);
and U13051 (N_13051,N_12958,N_12885);
or U13052 (N_13052,N_12910,N_12871);
or U13053 (N_13053,N_12927,N_12922);
nand U13054 (N_13054,N_12852,N_12897);
and U13055 (N_13055,N_12817,N_12966);
xor U13056 (N_13056,N_12989,N_12884);
nand U13057 (N_13057,N_12802,N_12986);
nor U13058 (N_13058,N_12873,N_12901);
and U13059 (N_13059,N_12860,N_12908);
and U13060 (N_13060,N_12847,N_12856);
nor U13061 (N_13061,N_12985,N_12894);
and U13062 (N_13062,N_12866,N_12865);
or U13063 (N_13063,N_12844,N_12935);
xor U13064 (N_13064,N_12974,N_12843);
xnor U13065 (N_13065,N_12945,N_12990);
nor U13066 (N_13066,N_12936,N_12809);
nor U13067 (N_13067,N_12914,N_12970);
nor U13068 (N_13068,N_12889,N_12928);
nand U13069 (N_13069,N_12995,N_12831);
nor U13070 (N_13070,N_12924,N_12836);
xnor U13071 (N_13071,N_12979,N_12879);
and U13072 (N_13072,N_12925,N_12830);
or U13073 (N_13073,N_12851,N_12948);
nor U13074 (N_13074,N_12815,N_12993);
or U13075 (N_13075,N_12999,N_12812);
and U13076 (N_13076,N_12878,N_12826);
and U13077 (N_13077,N_12961,N_12998);
nor U13078 (N_13078,N_12825,N_12912);
or U13079 (N_13079,N_12875,N_12880);
nor U13080 (N_13080,N_12877,N_12857);
nand U13081 (N_13081,N_12811,N_12915);
and U13082 (N_13082,N_12835,N_12814);
and U13083 (N_13083,N_12834,N_12911);
xor U13084 (N_13084,N_12893,N_12929);
xor U13085 (N_13085,N_12822,N_12933);
xor U13086 (N_13086,N_12801,N_12996);
and U13087 (N_13087,N_12926,N_12890);
nor U13088 (N_13088,N_12828,N_12943);
or U13089 (N_13089,N_12992,N_12816);
xnor U13090 (N_13090,N_12994,N_12931);
xor U13091 (N_13091,N_12959,N_12938);
nand U13092 (N_13092,N_12932,N_12838);
and U13093 (N_13093,N_12962,N_12839);
nor U13094 (N_13094,N_12891,N_12819);
nand U13095 (N_13095,N_12913,N_12934);
and U13096 (N_13096,N_12895,N_12942);
nor U13097 (N_13097,N_12859,N_12862);
and U13098 (N_13098,N_12858,N_12896);
xnor U13099 (N_13099,N_12953,N_12991);
nor U13100 (N_13100,N_12865,N_12962);
or U13101 (N_13101,N_12870,N_12921);
or U13102 (N_13102,N_12960,N_12941);
nand U13103 (N_13103,N_12958,N_12892);
and U13104 (N_13104,N_12976,N_12926);
nor U13105 (N_13105,N_12899,N_12868);
nor U13106 (N_13106,N_12852,N_12805);
or U13107 (N_13107,N_12973,N_12878);
nor U13108 (N_13108,N_12917,N_12934);
and U13109 (N_13109,N_12817,N_12837);
or U13110 (N_13110,N_12821,N_12989);
and U13111 (N_13111,N_12840,N_12966);
or U13112 (N_13112,N_12994,N_12900);
and U13113 (N_13113,N_12918,N_12883);
or U13114 (N_13114,N_12875,N_12998);
or U13115 (N_13115,N_12958,N_12874);
or U13116 (N_13116,N_12943,N_12867);
xor U13117 (N_13117,N_12820,N_12996);
and U13118 (N_13118,N_12871,N_12858);
xnor U13119 (N_13119,N_12846,N_12867);
and U13120 (N_13120,N_12818,N_12941);
xnor U13121 (N_13121,N_12922,N_12887);
nor U13122 (N_13122,N_12841,N_12972);
nor U13123 (N_13123,N_12879,N_12914);
nand U13124 (N_13124,N_12885,N_12863);
xnor U13125 (N_13125,N_12941,N_12950);
xnor U13126 (N_13126,N_12939,N_12839);
xnor U13127 (N_13127,N_12967,N_12989);
nor U13128 (N_13128,N_12890,N_12857);
nor U13129 (N_13129,N_12998,N_12886);
or U13130 (N_13130,N_12912,N_12861);
xor U13131 (N_13131,N_12858,N_12988);
and U13132 (N_13132,N_12862,N_12923);
nor U13133 (N_13133,N_12957,N_12844);
nand U13134 (N_13134,N_12805,N_12880);
or U13135 (N_13135,N_12930,N_12812);
or U13136 (N_13136,N_12846,N_12995);
or U13137 (N_13137,N_12960,N_12803);
nand U13138 (N_13138,N_12804,N_12998);
nand U13139 (N_13139,N_12989,N_12921);
or U13140 (N_13140,N_12988,N_12868);
nand U13141 (N_13141,N_12934,N_12861);
nand U13142 (N_13142,N_12883,N_12841);
and U13143 (N_13143,N_12971,N_12852);
nor U13144 (N_13144,N_12814,N_12885);
or U13145 (N_13145,N_12909,N_12959);
and U13146 (N_13146,N_12993,N_12899);
or U13147 (N_13147,N_12947,N_12951);
and U13148 (N_13148,N_12811,N_12990);
and U13149 (N_13149,N_12916,N_12883);
or U13150 (N_13150,N_12838,N_12965);
or U13151 (N_13151,N_12973,N_12852);
and U13152 (N_13152,N_12964,N_12935);
xor U13153 (N_13153,N_12881,N_12959);
nor U13154 (N_13154,N_12847,N_12802);
xnor U13155 (N_13155,N_12939,N_12822);
xnor U13156 (N_13156,N_12848,N_12851);
nand U13157 (N_13157,N_12828,N_12825);
nor U13158 (N_13158,N_12923,N_12951);
nand U13159 (N_13159,N_12849,N_12810);
nor U13160 (N_13160,N_12891,N_12909);
or U13161 (N_13161,N_12957,N_12867);
or U13162 (N_13162,N_12946,N_12982);
nor U13163 (N_13163,N_12832,N_12986);
nor U13164 (N_13164,N_12866,N_12827);
nand U13165 (N_13165,N_12959,N_12988);
and U13166 (N_13166,N_12957,N_12945);
or U13167 (N_13167,N_12970,N_12864);
xor U13168 (N_13168,N_12808,N_12834);
nor U13169 (N_13169,N_12931,N_12804);
or U13170 (N_13170,N_12848,N_12970);
xnor U13171 (N_13171,N_12979,N_12949);
nor U13172 (N_13172,N_12852,N_12929);
or U13173 (N_13173,N_12920,N_12831);
nor U13174 (N_13174,N_12906,N_12935);
nand U13175 (N_13175,N_12988,N_12862);
nand U13176 (N_13176,N_12870,N_12844);
nand U13177 (N_13177,N_12999,N_12808);
nor U13178 (N_13178,N_12807,N_12983);
and U13179 (N_13179,N_12994,N_12881);
xnor U13180 (N_13180,N_12820,N_12974);
xnor U13181 (N_13181,N_12893,N_12932);
nand U13182 (N_13182,N_12940,N_12836);
nand U13183 (N_13183,N_12996,N_12946);
or U13184 (N_13184,N_12958,N_12992);
nand U13185 (N_13185,N_12933,N_12816);
nand U13186 (N_13186,N_12811,N_12825);
nand U13187 (N_13187,N_12872,N_12952);
nor U13188 (N_13188,N_12984,N_12822);
and U13189 (N_13189,N_12899,N_12905);
and U13190 (N_13190,N_12839,N_12822);
nand U13191 (N_13191,N_12988,N_12860);
nand U13192 (N_13192,N_12916,N_12843);
nand U13193 (N_13193,N_12860,N_12993);
and U13194 (N_13194,N_12936,N_12992);
nor U13195 (N_13195,N_12911,N_12927);
or U13196 (N_13196,N_12990,N_12978);
xnor U13197 (N_13197,N_12861,N_12807);
xnor U13198 (N_13198,N_12936,N_12822);
xnor U13199 (N_13199,N_12837,N_12957);
and U13200 (N_13200,N_13044,N_13175);
nand U13201 (N_13201,N_13015,N_13006);
nor U13202 (N_13202,N_13143,N_13027);
xnor U13203 (N_13203,N_13181,N_13016);
and U13204 (N_13204,N_13174,N_13045);
xor U13205 (N_13205,N_13099,N_13190);
xor U13206 (N_13206,N_13085,N_13079);
or U13207 (N_13207,N_13157,N_13128);
xnor U13208 (N_13208,N_13165,N_13139);
xnor U13209 (N_13209,N_13168,N_13105);
or U13210 (N_13210,N_13014,N_13194);
and U13211 (N_13211,N_13127,N_13001);
nor U13212 (N_13212,N_13028,N_13057);
or U13213 (N_13213,N_13171,N_13197);
nand U13214 (N_13214,N_13198,N_13107);
nand U13215 (N_13215,N_13152,N_13151);
xnor U13216 (N_13216,N_13004,N_13133);
xor U13217 (N_13217,N_13131,N_13073);
and U13218 (N_13218,N_13034,N_13109);
nand U13219 (N_13219,N_13180,N_13108);
and U13220 (N_13220,N_13160,N_13035);
xnor U13221 (N_13221,N_13040,N_13091);
xnor U13222 (N_13222,N_13162,N_13068);
or U13223 (N_13223,N_13049,N_13067);
xor U13224 (N_13224,N_13191,N_13110);
nor U13225 (N_13225,N_13195,N_13053);
nand U13226 (N_13226,N_13169,N_13173);
xor U13227 (N_13227,N_13059,N_13005);
nor U13228 (N_13228,N_13084,N_13142);
and U13229 (N_13229,N_13043,N_13156);
nand U13230 (N_13230,N_13122,N_13000);
xnor U13231 (N_13231,N_13101,N_13096);
or U13232 (N_13232,N_13126,N_13124);
nor U13233 (N_13233,N_13080,N_13055);
nor U13234 (N_13234,N_13026,N_13095);
or U13235 (N_13235,N_13064,N_13137);
nor U13236 (N_13236,N_13052,N_13003);
and U13237 (N_13237,N_13086,N_13012);
nor U13238 (N_13238,N_13163,N_13187);
nor U13239 (N_13239,N_13058,N_13118);
nand U13240 (N_13240,N_13112,N_13042);
or U13241 (N_13241,N_13141,N_13022);
or U13242 (N_13242,N_13039,N_13177);
or U13243 (N_13243,N_13116,N_13088);
and U13244 (N_13244,N_13150,N_13078);
nor U13245 (N_13245,N_13007,N_13037);
nand U13246 (N_13246,N_13065,N_13036);
xor U13247 (N_13247,N_13129,N_13149);
and U13248 (N_13248,N_13009,N_13071);
nand U13249 (N_13249,N_13054,N_13106);
nor U13250 (N_13250,N_13102,N_13025);
nand U13251 (N_13251,N_13020,N_13094);
nand U13252 (N_13252,N_13083,N_13046);
or U13253 (N_13253,N_13183,N_13061);
xor U13254 (N_13254,N_13038,N_13104);
or U13255 (N_13255,N_13087,N_13048);
nand U13256 (N_13256,N_13184,N_13125);
xor U13257 (N_13257,N_13063,N_13056);
xnor U13258 (N_13258,N_13188,N_13170);
nor U13259 (N_13259,N_13013,N_13135);
or U13260 (N_13260,N_13074,N_13117);
or U13261 (N_13261,N_13111,N_13144);
or U13262 (N_13262,N_13097,N_13070);
or U13263 (N_13263,N_13167,N_13062);
nor U13264 (N_13264,N_13134,N_13178);
xnor U13265 (N_13265,N_13093,N_13089);
nand U13266 (N_13266,N_13164,N_13017);
or U13267 (N_13267,N_13092,N_13132);
nand U13268 (N_13268,N_13008,N_13075);
nand U13269 (N_13269,N_13138,N_13023);
nand U13270 (N_13270,N_13032,N_13147);
xnor U13271 (N_13271,N_13050,N_13186);
xor U13272 (N_13272,N_13161,N_13182);
and U13273 (N_13273,N_13192,N_13030);
nor U13274 (N_13274,N_13098,N_13090);
nor U13275 (N_13275,N_13051,N_13193);
xor U13276 (N_13276,N_13021,N_13154);
nand U13277 (N_13277,N_13189,N_13024);
xor U13278 (N_13278,N_13176,N_13185);
nor U13279 (N_13279,N_13081,N_13120);
nor U13280 (N_13280,N_13100,N_13011);
nor U13281 (N_13281,N_13069,N_13018);
nor U13282 (N_13282,N_13076,N_13010);
nor U13283 (N_13283,N_13130,N_13066);
nor U13284 (N_13284,N_13047,N_13145);
nor U13285 (N_13285,N_13172,N_13029);
or U13286 (N_13286,N_13072,N_13113);
and U13287 (N_13287,N_13123,N_13199);
or U13288 (N_13288,N_13148,N_13019);
nand U13289 (N_13289,N_13119,N_13136);
nor U13290 (N_13290,N_13121,N_13041);
nand U13291 (N_13291,N_13179,N_13146);
or U13292 (N_13292,N_13158,N_13115);
xor U13293 (N_13293,N_13060,N_13155);
and U13294 (N_13294,N_13166,N_13153);
nor U13295 (N_13295,N_13077,N_13031);
nor U13296 (N_13296,N_13159,N_13140);
nor U13297 (N_13297,N_13196,N_13114);
and U13298 (N_13298,N_13033,N_13002);
nor U13299 (N_13299,N_13103,N_13082);
nand U13300 (N_13300,N_13164,N_13140);
xor U13301 (N_13301,N_13025,N_13106);
xor U13302 (N_13302,N_13036,N_13049);
or U13303 (N_13303,N_13152,N_13186);
or U13304 (N_13304,N_13074,N_13098);
and U13305 (N_13305,N_13026,N_13140);
xnor U13306 (N_13306,N_13089,N_13066);
or U13307 (N_13307,N_13070,N_13189);
nand U13308 (N_13308,N_13169,N_13190);
nor U13309 (N_13309,N_13095,N_13031);
nand U13310 (N_13310,N_13196,N_13113);
nor U13311 (N_13311,N_13071,N_13141);
or U13312 (N_13312,N_13080,N_13179);
nor U13313 (N_13313,N_13101,N_13198);
or U13314 (N_13314,N_13008,N_13140);
xnor U13315 (N_13315,N_13193,N_13154);
xor U13316 (N_13316,N_13183,N_13122);
nor U13317 (N_13317,N_13194,N_13153);
and U13318 (N_13318,N_13004,N_13193);
or U13319 (N_13319,N_13198,N_13120);
nor U13320 (N_13320,N_13141,N_13107);
xor U13321 (N_13321,N_13190,N_13171);
or U13322 (N_13322,N_13146,N_13101);
or U13323 (N_13323,N_13029,N_13054);
or U13324 (N_13324,N_13142,N_13090);
or U13325 (N_13325,N_13120,N_13177);
nor U13326 (N_13326,N_13175,N_13186);
or U13327 (N_13327,N_13038,N_13009);
nand U13328 (N_13328,N_13031,N_13191);
xor U13329 (N_13329,N_13160,N_13024);
or U13330 (N_13330,N_13182,N_13196);
and U13331 (N_13331,N_13054,N_13053);
and U13332 (N_13332,N_13015,N_13082);
nor U13333 (N_13333,N_13128,N_13102);
nor U13334 (N_13334,N_13055,N_13074);
or U13335 (N_13335,N_13106,N_13119);
nor U13336 (N_13336,N_13140,N_13141);
nand U13337 (N_13337,N_13133,N_13137);
nand U13338 (N_13338,N_13136,N_13104);
and U13339 (N_13339,N_13059,N_13113);
and U13340 (N_13340,N_13087,N_13186);
nand U13341 (N_13341,N_13170,N_13169);
xor U13342 (N_13342,N_13027,N_13073);
and U13343 (N_13343,N_13195,N_13067);
xor U13344 (N_13344,N_13083,N_13052);
xor U13345 (N_13345,N_13013,N_13046);
nor U13346 (N_13346,N_13006,N_13155);
or U13347 (N_13347,N_13058,N_13055);
or U13348 (N_13348,N_13115,N_13077);
xor U13349 (N_13349,N_13174,N_13081);
xnor U13350 (N_13350,N_13048,N_13185);
nand U13351 (N_13351,N_13127,N_13054);
and U13352 (N_13352,N_13114,N_13110);
and U13353 (N_13353,N_13187,N_13107);
or U13354 (N_13354,N_13079,N_13035);
and U13355 (N_13355,N_13168,N_13162);
nor U13356 (N_13356,N_13107,N_13071);
or U13357 (N_13357,N_13166,N_13184);
or U13358 (N_13358,N_13040,N_13024);
xor U13359 (N_13359,N_13095,N_13007);
nor U13360 (N_13360,N_13147,N_13065);
nand U13361 (N_13361,N_13014,N_13010);
xor U13362 (N_13362,N_13093,N_13162);
and U13363 (N_13363,N_13141,N_13095);
or U13364 (N_13364,N_13162,N_13090);
nand U13365 (N_13365,N_13080,N_13058);
or U13366 (N_13366,N_13124,N_13054);
nor U13367 (N_13367,N_13040,N_13106);
nand U13368 (N_13368,N_13074,N_13163);
nand U13369 (N_13369,N_13151,N_13059);
xnor U13370 (N_13370,N_13072,N_13080);
xnor U13371 (N_13371,N_13044,N_13047);
and U13372 (N_13372,N_13139,N_13019);
nor U13373 (N_13373,N_13098,N_13179);
or U13374 (N_13374,N_13126,N_13011);
and U13375 (N_13375,N_13167,N_13055);
or U13376 (N_13376,N_13029,N_13001);
nand U13377 (N_13377,N_13162,N_13155);
or U13378 (N_13378,N_13033,N_13116);
nand U13379 (N_13379,N_13128,N_13162);
xor U13380 (N_13380,N_13012,N_13024);
and U13381 (N_13381,N_13189,N_13091);
and U13382 (N_13382,N_13091,N_13051);
nand U13383 (N_13383,N_13092,N_13067);
or U13384 (N_13384,N_13087,N_13030);
nand U13385 (N_13385,N_13003,N_13002);
nand U13386 (N_13386,N_13009,N_13172);
nand U13387 (N_13387,N_13043,N_13138);
and U13388 (N_13388,N_13159,N_13188);
or U13389 (N_13389,N_13085,N_13142);
or U13390 (N_13390,N_13157,N_13012);
and U13391 (N_13391,N_13020,N_13140);
xnor U13392 (N_13392,N_13033,N_13134);
and U13393 (N_13393,N_13126,N_13184);
nand U13394 (N_13394,N_13057,N_13156);
and U13395 (N_13395,N_13013,N_13093);
xor U13396 (N_13396,N_13027,N_13176);
nand U13397 (N_13397,N_13070,N_13100);
nor U13398 (N_13398,N_13160,N_13081);
or U13399 (N_13399,N_13131,N_13036);
or U13400 (N_13400,N_13221,N_13324);
nor U13401 (N_13401,N_13271,N_13357);
nand U13402 (N_13402,N_13375,N_13363);
and U13403 (N_13403,N_13372,N_13264);
or U13404 (N_13404,N_13213,N_13371);
and U13405 (N_13405,N_13361,N_13376);
nand U13406 (N_13406,N_13322,N_13308);
xor U13407 (N_13407,N_13380,N_13398);
and U13408 (N_13408,N_13340,N_13311);
nor U13409 (N_13409,N_13339,N_13267);
nand U13410 (N_13410,N_13240,N_13342);
or U13411 (N_13411,N_13210,N_13281);
nor U13412 (N_13412,N_13200,N_13266);
xor U13413 (N_13413,N_13358,N_13208);
or U13414 (N_13414,N_13270,N_13283);
nor U13415 (N_13415,N_13237,N_13291);
nor U13416 (N_13416,N_13222,N_13217);
and U13417 (N_13417,N_13238,N_13223);
or U13418 (N_13418,N_13309,N_13243);
or U13419 (N_13419,N_13337,N_13293);
xor U13420 (N_13420,N_13234,N_13299);
or U13421 (N_13421,N_13352,N_13258);
nor U13422 (N_13422,N_13321,N_13317);
nor U13423 (N_13423,N_13306,N_13335);
xor U13424 (N_13424,N_13360,N_13385);
xor U13425 (N_13425,N_13301,N_13215);
nand U13426 (N_13426,N_13250,N_13367);
nand U13427 (N_13427,N_13316,N_13334);
nor U13428 (N_13428,N_13287,N_13260);
xnor U13429 (N_13429,N_13288,N_13318);
and U13430 (N_13430,N_13297,N_13214);
xor U13431 (N_13431,N_13310,N_13298);
nor U13432 (N_13432,N_13354,N_13303);
nor U13433 (N_13433,N_13265,N_13349);
nor U13434 (N_13434,N_13353,N_13272);
nor U13435 (N_13435,N_13295,N_13290);
xor U13436 (N_13436,N_13255,N_13248);
xor U13437 (N_13437,N_13356,N_13276);
xor U13438 (N_13438,N_13285,N_13379);
nand U13439 (N_13439,N_13278,N_13279);
xnor U13440 (N_13440,N_13331,N_13229);
xnor U13441 (N_13441,N_13241,N_13256);
and U13442 (N_13442,N_13370,N_13239);
and U13443 (N_13443,N_13253,N_13249);
or U13444 (N_13444,N_13254,N_13381);
nand U13445 (N_13445,N_13315,N_13343);
nor U13446 (N_13446,N_13206,N_13368);
xor U13447 (N_13447,N_13232,N_13244);
or U13448 (N_13448,N_13233,N_13228);
or U13449 (N_13449,N_13203,N_13336);
and U13450 (N_13450,N_13323,N_13269);
or U13451 (N_13451,N_13302,N_13224);
or U13452 (N_13452,N_13209,N_13330);
nand U13453 (N_13453,N_13227,N_13319);
xnor U13454 (N_13454,N_13274,N_13390);
nand U13455 (N_13455,N_13235,N_13263);
or U13456 (N_13456,N_13226,N_13350);
nor U13457 (N_13457,N_13219,N_13216);
or U13458 (N_13458,N_13378,N_13369);
and U13459 (N_13459,N_13262,N_13236);
and U13460 (N_13460,N_13383,N_13355);
or U13461 (N_13461,N_13396,N_13364);
or U13462 (N_13462,N_13218,N_13300);
xnor U13463 (N_13463,N_13393,N_13246);
nand U13464 (N_13464,N_13327,N_13391);
and U13465 (N_13465,N_13389,N_13328);
nand U13466 (N_13466,N_13325,N_13280);
nor U13467 (N_13467,N_13252,N_13320);
nor U13468 (N_13468,N_13304,N_13366);
or U13469 (N_13469,N_13201,N_13386);
and U13470 (N_13470,N_13273,N_13387);
nor U13471 (N_13471,N_13332,N_13259);
nand U13472 (N_13472,N_13212,N_13225);
and U13473 (N_13473,N_13351,N_13348);
xnor U13474 (N_13474,N_13314,N_13220);
or U13475 (N_13475,N_13392,N_13268);
or U13476 (N_13476,N_13382,N_13245);
nor U13477 (N_13477,N_13333,N_13230);
and U13478 (N_13478,N_13211,N_13277);
and U13479 (N_13479,N_13261,N_13346);
nand U13480 (N_13480,N_13247,N_13275);
xor U13481 (N_13481,N_13313,N_13202);
and U13482 (N_13482,N_13312,N_13377);
and U13483 (N_13483,N_13344,N_13257);
nand U13484 (N_13484,N_13284,N_13397);
xnor U13485 (N_13485,N_13207,N_13399);
or U13486 (N_13486,N_13286,N_13338);
nand U13487 (N_13487,N_13359,N_13282);
and U13488 (N_13488,N_13345,N_13292);
or U13489 (N_13489,N_13341,N_13374);
nand U13490 (N_13490,N_13307,N_13365);
nand U13491 (N_13491,N_13329,N_13204);
and U13492 (N_13492,N_13388,N_13384);
xor U13493 (N_13493,N_13294,N_13362);
xor U13494 (N_13494,N_13347,N_13305);
nand U13495 (N_13495,N_13373,N_13296);
or U13496 (N_13496,N_13231,N_13395);
nand U13497 (N_13497,N_13326,N_13251);
or U13498 (N_13498,N_13205,N_13242);
or U13499 (N_13499,N_13289,N_13394);
xor U13500 (N_13500,N_13283,N_13386);
nor U13501 (N_13501,N_13345,N_13269);
and U13502 (N_13502,N_13397,N_13249);
and U13503 (N_13503,N_13258,N_13349);
nand U13504 (N_13504,N_13271,N_13395);
xnor U13505 (N_13505,N_13310,N_13271);
and U13506 (N_13506,N_13325,N_13302);
nand U13507 (N_13507,N_13337,N_13280);
xnor U13508 (N_13508,N_13356,N_13283);
nand U13509 (N_13509,N_13323,N_13272);
or U13510 (N_13510,N_13328,N_13278);
nor U13511 (N_13511,N_13297,N_13339);
and U13512 (N_13512,N_13211,N_13312);
and U13513 (N_13513,N_13273,N_13284);
xnor U13514 (N_13514,N_13293,N_13395);
or U13515 (N_13515,N_13362,N_13322);
nor U13516 (N_13516,N_13317,N_13395);
nor U13517 (N_13517,N_13312,N_13246);
and U13518 (N_13518,N_13231,N_13261);
xor U13519 (N_13519,N_13314,N_13328);
nand U13520 (N_13520,N_13386,N_13227);
nand U13521 (N_13521,N_13395,N_13240);
xnor U13522 (N_13522,N_13208,N_13315);
xor U13523 (N_13523,N_13339,N_13238);
and U13524 (N_13524,N_13349,N_13340);
and U13525 (N_13525,N_13382,N_13205);
or U13526 (N_13526,N_13310,N_13305);
nand U13527 (N_13527,N_13371,N_13396);
xor U13528 (N_13528,N_13220,N_13352);
and U13529 (N_13529,N_13226,N_13318);
and U13530 (N_13530,N_13237,N_13331);
nand U13531 (N_13531,N_13210,N_13338);
and U13532 (N_13532,N_13210,N_13202);
nor U13533 (N_13533,N_13353,N_13320);
nand U13534 (N_13534,N_13210,N_13341);
and U13535 (N_13535,N_13244,N_13379);
or U13536 (N_13536,N_13326,N_13369);
or U13537 (N_13537,N_13365,N_13219);
or U13538 (N_13538,N_13337,N_13212);
xnor U13539 (N_13539,N_13236,N_13307);
and U13540 (N_13540,N_13331,N_13396);
or U13541 (N_13541,N_13334,N_13307);
and U13542 (N_13542,N_13317,N_13318);
xnor U13543 (N_13543,N_13344,N_13275);
nor U13544 (N_13544,N_13380,N_13299);
nor U13545 (N_13545,N_13216,N_13265);
nor U13546 (N_13546,N_13305,N_13390);
nand U13547 (N_13547,N_13273,N_13299);
or U13548 (N_13548,N_13314,N_13333);
nor U13549 (N_13549,N_13362,N_13371);
xnor U13550 (N_13550,N_13237,N_13246);
or U13551 (N_13551,N_13299,N_13344);
nor U13552 (N_13552,N_13228,N_13368);
nand U13553 (N_13553,N_13226,N_13369);
nand U13554 (N_13554,N_13212,N_13204);
or U13555 (N_13555,N_13398,N_13235);
nor U13556 (N_13556,N_13350,N_13357);
and U13557 (N_13557,N_13297,N_13232);
and U13558 (N_13558,N_13209,N_13267);
nor U13559 (N_13559,N_13377,N_13211);
nand U13560 (N_13560,N_13313,N_13274);
nand U13561 (N_13561,N_13381,N_13277);
xor U13562 (N_13562,N_13231,N_13217);
and U13563 (N_13563,N_13232,N_13279);
or U13564 (N_13564,N_13244,N_13265);
nor U13565 (N_13565,N_13282,N_13377);
and U13566 (N_13566,N_13315,N_13214);
nand U13567 (N_13567,N_13336,N_13398);
nor U13568 (N_13568,N_13304,N_13298);
and U13569 (N_13569,N_13323,N_13364);
nor U13570 (N_13570,N_13224,N_13380);
nor U13571 (N_13571,N_13362,N_13255);
nor U13572 (N_13572,N_13324,N_13272);
xnor U13573 (N_13573,N_13345,N_13339);
xnor U13574 (N_13574,N_13244,N_13275);
or U13575 (N_13575,N_13320,N_13208);
or U13576 (N_13576,N_13383,N_13352);
nand U13577 (N_13577,N_13280,N_13391);
and U13578 (N_13578,N_13278,N_13236);
nand U13579 (N_13579,N_13224,N_13321);
or U13580 (N_13580,N_13302,N_13300);
nor U13581 (N_13581,N_13257,N_13230);
or U13582 (N_13582,N_13320,N_13373);
nand U13583 (N_13583,N_13305,N_13367);
or U13584 (N_13584,N_13255,N_13321);
nand U13585 (N_13585,N_13286,N_13248);
nand U13586 (N_13586,N_13395,N_13232);
nor U13587 (N_13587,N_13220,N_13334);
nand U13588 (N_13588,N_13282,N_13383);
nor U13589 (N_13589,N_13236,N_13285);
xor U13590 (N_13590,N_13204,N_13243);
xor U13591 (N_13591,N_13393,N_13278);
nor U13592 (N_13592,N_13328,N_13239);
and U13593 (N_13593,N_13397,N_13294);
and U13594 (N_13594,N_13281,N_13249);
nand U13595 (N_13595,N_13223,N_13384);
nand U13596 (N_13596,N_13288,N_13287);
xnor U13597 (N_13597,N_13217,N_13287);
and U13598 (N_13598,N_13307,N_13306);
and U13599 (N_13599,N_13276,N_13259);
xnor U13600 (N_13600,N_13516,N_13507);
xnor U13601 (N_13601,N_13537,N_13591);
or U13602 (N_13602,N_13588,N_13435);
nand U13603 (N_13603,N_13574,N_13590);
nand U13604 (N_13604,N_13517,N_13424);
xor U13605 (N_13605,N_13448,N_13446);
or U13606 (N_13606,N_13442,N_13431);
nand U13607 (N_13607,N_13553,N_13422);
or U13608 (N_13608,N_13562,N_13552);
or U13609 (N_13609,N_13429,N_13572);
xnor U13610 (N_13610,N_13579,N_13593);
or U13611 (N_13611,N_13470,N_13503);
or U13612 (N_13612,N_13462,N_13414);
xnor U13613 (N_13613,N_13556,N_13509);
or U13614 (N_13614,N_13454,N_13559);
and U13615 (N_13615,N_13491,N_13538);
xnor U13616 (N_13616,N_13411,N_13489);
or U13617 (N_13617,N_13499,N_13478);
nor U13618 (N_13618,N_13406,N_13510);
nand U13619 (N_13619,N_13571,N_13599);
or U13620 (N_13620,N_13474,N_13528);
and U13621 (N_13621,N_13465,N_13423);
or U13622 (N_13622,N_13487,N_13594);
nor U13623 (N_13623,N_13535,N_13455);
and U13624 (N_13624,N_13500,N_13586);
or U13625 (N_13625,N_13534,N_13531);
nand U13626 (N_13626,N_13432,N_13473);
and U13627 (N_13627,N_13527,N_13564);
xnor U13628 (N_13628,N_13416,N_13543);
xor U13629 (N_13629,N_13512,N_13549);
xnor U13630 (N_13630,N_13430,N_13480);
nor U13631 (N_13631,N_13496,N_13508);
and U13632 (N_13632,N_13463,N_13519);
or U13633 (N_13633,N_13420,N_13532);
and U13634 (N_13634,N_13436,N_13529);
xor U13635 (N_13635,N_13456,N_13418);
nand U13636 (N_13636,N_13449,N_13567);
nor U13637 (N_13637,N_13505,N_13597);
xor U13638 (N_13638,N_13410,N_13490);
xnor U13639 (N_13639,N_13511,N_13426);
and U13640 (N_13640,N_13539,N_13501);
nand U13641 (N_13641,N_13514,N_13578);
xnor U13642 (N_13642,N_13479,N_13583);
or U13643 (N_13643,N_13485,N_13585);
and U13644 (N_13644,N_13520,N_13550);
and U13645 (N_13645,N_13563,N_13548);
nor U13646 (N_13646,N_13427,N_13450);
nor U13647 (N_13647,N_13544,N_13542);
or U13648 (N_13648,N_13533,N_13481);
xor U13649 (N_13649,N_13400,N_13561);
nand U13650 (N_13650,N_13560,N_13558);
xor U13651 (N_13651,N_13472,N_13407);
and U13652 (N_13652,N_13566,N_13584);
and U13653 (N_13653,N_13513,N_13495);
nand U13654 (N_13654,N_13402,N_13595);
nand U13655 (N_13655,N_13405,N_13545);
and U13656 (N_13656,N_13569,N_13444);
xor U13657 (N_13657,N_13428,N_13441);
or U13658 (N_13658,N_13488,N_13541);
or U13659 (N_13659,N_13547,N_13408);
nand U13660 (N_13660,N_13592,N_13447);
nor U13661 (N_13661,N_13412,N_13482);
and U13662 (N_13662,N_13452,N_13518);
xor U13663 (N_13663,N_13555,N_13522);
or U13664 (N_13664,N_13460,N_13497);
or U13665 (N_13665,N_13443,N_13523);
nand U13666 (N_13666,N_13573,N_13453);
or U13667 (N_13667,N_13475,N_13425);
xor U13668 (N_13668,N_13576,N_13493);
and U13669 (N_13669,N_13434,N_13598);
nor U13670 (N_13670,N_13565,N_13540);
xor U13671 (N_13671,N_13477,N_13467);
xnor U13672 (N_13672,N_13451,N_13587);
xnor U13673 (N_13673,N_13498,N_13580);
xnor U13674 (N_13674,N_13536,N_13471);
or U13675 (N_13675,N_13464,N_13526);
nor U13676 (N_13676,N_13582,N_13417);
and U13677 (N_13677,N_13557,N_13581);
or U13678 (N_13678,N_13524,N_13596);
nor U13679 (N_13679,N_13403,N_13469);
nand U13680 (N_13680,N_13484,N_13437);
nor U13681 (N_13681,N_13445,N_13433);
nor U13682 (N_13682,N_13551,N_13401);
nor U13683 (N_13683,N_13466,N_13515);
xnor U13684 (N_13684,N_13440,N_13413);
or U13685 (N_13685,N_13530,N_13438);
nand U13686 (N_13686,N_13421,N_13483);
nand U13687 (N_13687,N_13459,N_13525);
nand U13688 (N_13688,N_13577,N_13415);
and U13689 (N_13689,N_13492,N_13409);
and U13690 (N_13690,N_13506,N_13521);
and U13691 (N_13691,N_13476,N_13554);
xnor U13692 (N_13692,N_13589,N_13575);
nand U13693 (N_13693,N_13457,N_13546);
and U13694 (N_13694,N_13458,N_13404);
nand U13695 (N_13695,N_13419,N_13494);
and U13696 (N_13696,N_13468,N_13486);
nand U13697 (N_13697,N_13568,N_13461);
nor U13698 (N_13698,N_13570,N_13439);
xor U13699 (N_13699,N_13502,N_13504);
or U13700 (N_13700,N_13557,N_13483);
xor U13701 (N_13701,N_13410,N_13454);
nand U13702 (N_13702,N_13458,N_13529);
and U13703 (N_13703,N_13583,N_13453);
nand U13704 (N_13704,N_13485,N_13524);
nor U13705 (N_13705,N_13445,N_13592);
nor U13706 (N_13706,N_13446,N_13533);
xnor U13707 (N_13707,N_13523,N_13415);
or U13708 (N_13708,N_13407,N_13417);
nor U13709 (N_13709,N_13540,N_13459);
and U13710 (N_13710,N_13447,N_13414);
nand U13711 (N_13711,N_13470,N_13560);
nor U13712 (N_13712,N_13550,N_13443);
nand U13713 (N_13713,N_13562,N_13488);
or U13714 (N_13714,N_13580,N_13566);
and U13715 (N_13715,N_13587,N_13453);
nand U13716 (N_13716,N_13452,N_13564);
nor U13717 (N_13717,N_13596,N_13588);
and U13718 (N_13718,N_13483,N_13417);
xnor U13719 (N_13719,N_13427,N_13471);
xor U13720 (N_13720,N_13502,N_13518);
or U13721 (N_13721,N_13407,N_13466);
nor U13722 (N_13722,N_13509,N_13449);
xnor U13723 (N_13723,N_13528,N_13453);
nand U13724 (N_13724,N_13422,N_13582);
nand U13725 (N_13725,N_13549,N_13557);
nand U13726 (N_13726,N_13482,N_13509);
nand U13727 (N_13727,N_13580,N_13518);
and U13728 (N_13728,N_13522,N_13546);
xor U13729 (N_13729,N_13440,N_13560);
nand U13730 (N_13730,N_13486,N_13560);
nor U13731 (N_13731,N_13585,N_13545);
or U13732 (N_13732,N_13507,N_13466);
nor U13733 (N_13733,N_13423,N_13552);
nor U13734 (N_13734,N_13479,N_13521);
nand U13735 (N_13735,N_13442,N_13550);
nor U13736 (N_13736,N_13418,N_13442);
xnor U13737 (N_13737,N_13404,N_13447);
and U13738 (N_13738,N_13446,N_13514);
nand U13739 (N_13739,N_13530,N_13443);
nand U13740 (N_13740,N_13572,N_13519);
xor U13741 (N_13741,N_13457,N_13535);
xor U13742 (N_13742,N_13427,N_13555);
xnor U13743 (N_13743,N_13473,N_13496);
and U13744 (N_13744,N_13406,N_13430);
xnor U13745 (N_13745,N_13549,N_13441);
nor U13746 (N_13746,N_13524,N_13447);
or U13747 (N_13747,N_13540,N_13525);
xor U13748 (N_13748,N_13444,N_13533);
and U13749 (N_13749,N_13559,N_13501);
nor U13750 (N_13750,N_13535,N_13482);
nor U13751 (N_13751,N_13417,N_13520);
nor U13752 (N_13752,N_13551,N_13495);
nand U13753 (N_13753,N_13480,N_13463);
nand U13754 (N_13754,N_13420,N_13579);
nor U13755 (N_13755,N_13487,N_13520);
xnor U13756 (N_13756,N_13453,N_13497);
and U13757 (N_13757,N_13404,N_13560);
nand U13758 (N_13758,N_13402,N_13429);
and U13759 (N_13759,N_13566,N_13497);
xor U13760 (N_13760,N_13562,N_13483);
nor U13761 (N_13761,N_13504,N_13561);
and U13762 (N_13762,N_13459,N_13561);
nand U13763 (N_13763,N_13506,N_13459);
nor U13764 (N_13764,N_13518,N_13434);
xor U13765 (N_13765,N_13551,N_13474);
and U13766 (N_13766,N_13424,N_13485);
nand U13767 (N_13767,N_13418,N_13574);
nor U13768 (N_13768,N_13429,N_13574);
nand U13769 (N_13769,N_13583,N_13575);
nor U13770 (N_13770,N_13523,N_13460);
nand U13771 (N_13771,N_13420,N_13405);
nand U13772 (N_13772,N_13588,N_13479);
nand U13773 (N_13773,N_13438,N_13488);
nand U13774 (N_13774,N_13595,N_13437);
or U13775 (N_13775,N_13498,N_13564);
xor U13776 (N_13776,N_13571,N_13582);
xnor U13777 (N_13777,N_13564,N_13470);
xnor U13778 (N_13778,N_13503,N_13524);
nand U13779 (N_13779,N_13537,N_13556);
and U13780 (N_13780,N_13577,N_13568);
xnor U13781 (N_13781,N_13474,N_13514);
and U13782 (N_13782,N_13521,N_13495);
nand U13783 (N_13783,N_13543,N_13477);
and U13784 (N_13784,N_13415,N_13552);
xor U13785 (N_13785,N_13589,N_13581);
or U13786 (N_13786,N_13494,N_13410);
nor U13787 (N_13787,N_13506,N_13508);
nand U13788 (N_13788,N_13431,N_13504);
and U13789 (N_13789,N_13564,N_13432);
nand U13790 (N_13790,N_13578,N_13573);
or U13791 (N_13791,N_13575,N_13457);
xnor U13792 (N_13792,N_13486,N_13430);
xnor U13793 (N_13793,N_13478,N_13501);
nor U13794 (N_13794,N_13585,N_13597);
nand U13795 (N_13795,N_13574,N_13416);
xnor U13796 (N_13796,N_13593,N_13464);
nand U13797 (N_13797,N_13415,N_13429);
nor U13798 (N_13798,N_13417,N_13454);
or U13799 (N_13799,N_13422,N_13403);
or U13800 (N_13800,N_13623,N_13744);
xnor U13801 (N_13801,N_13751,N_13765);
or U13802 (N_13802,N_13704,N_13777);
or U13803 (N_13803,N_13637,N_13721);
xnor U13804 (N_13804,N_13643,N_13621);
xor U13805 (N_13805,N_13701,N_13782);
xor U13806 (N_13806,N_13657,N_13702);
nand U13807 (N_13807,N_13709,N_13683);
nor U13808 (N_13808,N_13605,N_13767);
nand U13809 (N_13809,N_13770,N_13611);
nor U13810 (N_13810,N_13668,N_13633);
nor U13811 (N_13811,N_13719,N_13761);
and U13812 (N_13812,N_13635,N_13659);
or U13813 (N_13813,N_13641,N_13732);
and U13814 (N_13814,N_13646,N_13730);
or U13815 (N_13815,N_13707,N_13640);
nor U13816 (N_13816,N_13798,N_13674);
and U13817 (N_13817,N_13792,N_13726);
nand U13818 (N_13818,N_13787,N_13771);
nor U13819 (N_13819,N_13795,N_13727);
or U13820 (N_13820,N_13649,N_13601);
and U13821 (N_13821,N_13741,N_13628);
xnor U13822 (N_13822,N_13630,N_13753);
xor U13823 (N_13823,N_13670,N_13796);
xnor U13824 (N_13824,N_13612,N_13682);
nor U13825 (N_13825,N_13776,N_13626);
nor U13826 (N_13826,N_13661,N_13724);
nor U13827 (N_13827,N_13681,N_13631);
and U13828 (N_13828,N_13642,N_13693);
xnor U13829 (N_13829,N_13757,N_13676);
nor U13830 (N_13830,N_13734,N_13624);
nor U13831 (N_13831,N_13653,N_13699);
nand U13832 (N_13832,N_13691,N_13645);
nand U13833 (N_13833,N_13692,N_13754);
nor U13834 (N_13834,N_13619,N_13662);
xnor U13835 (N_13835,N_13618,N_13717);
and U13836 (N_13836,N_13614,N_13775);
nor U13837 (N_13837,N_13625,N_13783);
xor U13838 (N_13838,N_13784,N_13663);
nor U13839 (N_13839,N_13627,N_13759);
or U13840 (N_13840,N_13684,N_13689);
and U13841 (N_13841,N_13671,N_13742);
or U13842 (N_13842,N_13773,N_13660);
nor U13843 (N_13843,N_13636,N_13698);
xnor U13844 (N_13844,N_13644,N_13603);
nor U13845 (N_13845,N_13779,N_13634);
nor U13846 (N_13846,N_13665,N_13703);
nand U13847 (N_13847,N_13738,N_13685);
xor U13848 (N_13848,N_13791,N_13600);
xnor U13849 (N_13849,N_13788,N_13694);
nor U13850 (N_13850,N_13604,N_13747);
nor U13851 (N_13851,N_13615,N_13655);
nand U13852 (N_13852,N_13743,N_13715);
nor U13853 (N_13853,N_13737,N_13731);
nand U13854 (N_13854,N_13610,N_13652);
or U13855 (N_13855,N_13716,N_13697);
xor U13856 (N_13856,N_13678,N_13772);
or U13857 (N_13857,N_13793,N_13733);
and U13858 (N_13858,N_13718,N_13769);
or U13859 (N_13859,N_13677,N_13735);
or U13860 (N_13860,N_13749,N_13667);
nand U13861 (N_13861,N_13648,N_13745);
xor U13862 (N_13862,N_13764,N_13608);
xor U13863 (N_13863,N_13613,N_13758);
nand U13864 (N_13864,N_13647,N_13755);
and U13865 (N_13865,N_13654,N_13690);
nor U13866 (N_13866,N_13797,N_13713);
or U13867 (N_13867,N_13687,N_13750);
or U13868 (N_13868,N_13658,N_13622);
xnor U13869 (N_13869,N_13760,N_13714);
nor U13870 (N_13870,N_13786,N_13706);
or U13871 (N_13871,N_13638,N_13705);
nand U13872 (N_13872,N_13609,N_13639);
nor U13873 (N_13873,N_13606,N_13680);
or U13874 (N_13874,N_13650,N_13708);
nor U13875 (N_13875,N_13710,N_13728);
nor U13876 (N_13876,N_13763,N_13686);
nand U13877 (N_13877,N_13712,N_13672);
nor U13878 (N_13878,N_13666,N_13790);
or U13879 (N_13879,N_13746,N_13673);
nand U13880 (N_13880,N_13679,N_13656);
nor U13881 (N_13881,N_13688,N_13748);
nor U13882 (N_13882,N_13616,N_13794);
or U13883 (N_13883,N_13740,N_13739);
and U13884 (N_13884,N_13756,N_13711);
or U13885 (N_13885,N_13632,N_13766);
and U13886 (N_13886,N_13785,N_13778);
or U13887 (N_13887,N_13664,N_13729);
nor U13888 (N_13888,N_13736,N_13696);
and U13889 (N_13889,N_13780,N_13725);
and U13890 (N_13890,N_13752,N_13669);
nor U13891 (N_13891,N_13781,N_13695);
xnor U13892 (N_13892,N_13700,N_13620);
xnor U13893 (N_13893,N_13768,N_13651);
nand U13894 (N_13894,N_13762,N_13629);
and U13895 (N_13895,N_13789,N_13799);
and U13896 (N_13896,N_13607,N_13675);
and U13897 (N_13897,N_13720,N_13617);
and U13898 (N_13898,N_13602,N_13774);
xor U13899 (N_13899,N_13723,N_13722);
xor U13900 (N_13900,N_13618,N_13613);
or U13901 (N_13901,N_13766,N_13670);
xnor U13902 (N_13902,N_13649,N_13681);
xnor U13903 (N_13903,N_13669,N_13657);
nor U13904 (N_13904,N_13787,N_13608);
and U13905 (N_13905,N_13735,N_13632);
or U13906 (N_13906,N_13759,N_13739);
xor U13907 (N_13907,N_13718,N_13600);
xnor U13908 (N_13908,N_13638,N_13617);
or U13909 (N_13909,N_13697,N_13634);
nor U13910 (N_13910,N_13651,N_13610);
and U13911 (N_13911,N_13610,N_13769);
and U13912 (N_13912,N_13657,N_13762);
nand U13913 (N_13913,N_13738,N_13611);
or U13914 (N_13914,N_13605,N_13764);
xnor U13915 (N_13915,N_13723,N_13786);
nor U13916 (N_13916,N_13719,N_13747);
or U13917 (N_13917,N_13712,N_13671);
and U13918 (N_13918,N_13660,N_13797);
nand U13919 (N_13919,N_13781,N_13712);
or U13920 (N_13920,N_13657,N_13722);
xnor U13921 (N_13921,N_13673,N_13750);
and U13922 (N_13922,N_13767,N_13753);
nand U13923 (N_13923,N_13621,N_13757);
or U13924 (N_13924,N_13684,N_13659);
and U13925 (N_13925,N_13608,N_13721);
and U13926 (N_13926,N_13690,N_13605);
nand U13927 (N_13927,N_13672,N_13600);
and U13928 (N_13928,N_13757,N_13630);
nand U13929 (N_13929,N_13648,N_13708);
or U13930 (N_13930,N_13691,N_13702);
nand U13931 (N_13931,N_13794,N_13787);
xor U13932 (N_13932,N_13689,N_13743);
nor U13933 (N_13933,N_13614,N_13699);
and U13934 (N_13934,N_13789,N_13671);
nor U13935 (N_13935,N_13694,N_13681);
nand U13936 (N_13936,N_13664,N_13752);
or U13937 (N_13937,N_13762,N_13689);
xor U13938 (N_13938,N_13783,N_13632);
nor U13939 (N_13939,N_13784,N_13716);
xnor U13940 (N_13940,N_13759,N_13726);
xnor U13941 (N_13941,N_13752,N_13774);
xor U13942 (N_13942,N_13605,N_13656);
nand U13943 (N_13943,N_13620,N_13690);
and U13944 (N_13944,N_13712,N_13698);
and U13945 (N_13945,N_13738,N_13784);
or U13946 (N_13946,N_13687,N_13682);
xor U13947 (N_13947,N_13749,N_13709);
nand U13948 (N_13948,N_13780,N_13787);
xor U13949 (N_13949,N_13788,N_13683);
nor U13950 (N_13950,N_13685,N_13725);
or U13951 (N_13951,N_13659,N_13636);
xnor U13952 (N_13952,N_13665,N_13626);
and U13953 (N_13953,N_13605,N_13792);
and U13954 (N_13954,N_13716,N_13710);
nand U13955 (N_13955,N_13733,N_13782);
nand U13956 (N_13956,N_13605,N_13783);
nor U13957 (N_13957,N_13720,N_13630);
nand U13958 (N_13958,N_13658,N_13691);
nand U13959 (N_13959,N_13705,N_13740);
and U13960 (N_13960,N_13630,N_13742);
and U13961 (N_13961,N_13654,N_13605);
xor U13962 (N_13962,N_13717,N_13787);
nand U13963 (N_13963,N_13751,N_13671);
xor U13964 (N_13964,N_13691,N_13674);
or U13965 (N_13965,N_13769,N_13746);
nand U13966 (N_13966,N_13658,N_13696);
or U13967 (N_13967,N_13685,N_13713);
xnor U13968 (N_13968,N_13715,N_13704);
or U13969 (N_13969,N_13659,N_13737);
or U13970 (N_13970,N_13664,N_13731);
or U13971 (N_13971,N_13774,N_13673);
and U13972 (N_13972,N_13640,N_13638);
and U13973 (N_13973,N_13773,N_13605);
or U13974 (N_13974,N_13780,N_13769);
and U13975 (N_13975,N_13736,N_13651);
nand U13976 (N_13976,N_13621,N_13791);
nand U13977 (N_13977,N_13693,N_13672);
xnor U13978 (N_13978,N_13783,N_13759);
nor U13979 (N_13979,N_13693,N_13779);
or U13980 (N_13980,N_13789,N_13653);
or U13981 (N_13981,N_13663,N_13648);
xor U13982 (N_13982,N_13660,N_13631);
xnor U13983 (N_13983,N_13670,N_13644);
or U13984 (N_13984,N_13640,N_13628);
and U13985 (N_13985,N_13643,N_13679);
nor U13986 (N_13986,N_13712,N_13773);
xor U13987 (N_13987,N_13639,N_13737);
nor U13988 (N_13988,N_13713,N_13653);
nor U13989 (N_13989,N_13730,N_13748);
or U13990 (N_13990,N_13662,N_13773);
nand U13991 (N_13991,N_13637,N_13629);
or U13992 (N_13992,N_13655,N_13702);
or U13993 (N_13993,N_13725,N_13665);
xnor U13994 (N_13994,N_13651,N_13717);
nor U13995 (N_13995,N_13723,N_13709);
or U13996 (N_13996,N_13734,N_13694);
and U13997 (N_13997,N_13668,N_13745);
and U13998 (N_13998,N_13725,N_13747);
or U13999 (N_13999,N_13747,N_13640);
or U14000 (N_14000,N_13842,N_13886);
nor U14001 (N_14001,N_13982,N_13864);
xnor U14002 (N_14002,N_13879,N_13805);
xor U14003 (N_14003,N_13899,N_13984);
xnor U14004 (N_14004,N_13845,N_13839);
or U14005 (N_14005,N_13870,N_13862);
and U14006 (N_14006,N_13833,N_13882);
nand U14007 (N_14007,N_13951,N_13876);
nor U14008 (N_14008,N_13841,N_13850);
nor U14009 (N_14009,N_13959,N_13961);
and U14010 (N_14010,N_13902,N_13928);
nor U14011 (N_14011,N_13975,N_13847);
nor U14012 (N_14012,N_13835,N_13884);
nor U14013 (N_14013,N_13904,N_13856);
or U14014 (N_14014,N_13919,N_13848);
and U14015 (N_14015,N_13985,N_13859);
xor U14016 (N_14016,N_13808,N_13943);
nor U14017 (N_14017,N_13916,N_13863);
or U14018 (N_14018,N_13988,N_13939);
nand U14019 (N_14019,N_13986,N_13803);
nor U14020 (N_14020,N_13800,N_13852);
xor U14021 (N_14021,N_13950,N_13924);
or U14022 (N_14022,N_13960,N_13926);
nand U14023 (N_14023,N_13991,N_13962);
and U14024 (N_14024,N_13836,N_13909);
nor U14025 (N_14025,N_13815,N_13963);
nor U14026 (N_14026,N_13958,N_13866);
and U14027 (N_14027,N_13810,N_13898);
xor U14028 (N_14028,N_13905,N_13846);
and U14029 (N_14029,N_13807,N_13925);
nor U14030 (N_14030,N_13908,N_13977);
xor U14031 (N_14031,N_13964,N_13933);
nor U14032 (N_14032,N_13981,N_13947);
nor U14033 (N_14033,N_13930,N_13920);
xnor U14034 (N_14034,N_13997,N_13858);
nor U14035 (N_14035,N_13900,N_13942);
or U14036 (N_14036,N_13914,N_13826);
or U14037 (N_14037,N_13946,N_13891);
nor U14038 (N_14038,N_13918,N_13821);
nand U14039 (N_14039,N_13830,N_13978);
or U14040 (N_14040,N_13813,N_13907);
nand U14041 (N_14041,N_13832,N_13871);
and U14042 (N_14042,N_13910,N_13809);
nor U14043 (N_14043,N_13992,N_13831);
and U14044 (N_14044,N_13817,N_13880);
and U14045 (N_14045,N_13989,N_13921);
or U14046 (N_14046,N_13872,N_13865);
xnor U14047 (N_14047,N_13806,N_13953);
and U14048 (N_14048,N_13893,N_13973);
nand U14049 (N_14049,N_13976,N_13861);
nand U14050 (N_14050,N_13881,N_13811);
or U14051 (N_14051,N_13929,N_13838);
nor U14052 (N_14052,N_13990,N_13972);
nand U14053 (N_14053,N_13954,N_13849);
nor U14054 (N_14054,N_13913,N_13936);
nor U14055 (N_14055,N_13857,N_13874);
xnor U14056 (N_14056,N_13814,N_13843);
xnor U14057 (N_14057,N_13801,N_13935);
or U14058 (N_14058,N_13955,N_13828);
or U14059 (N_14059,N_13877,N_13802);
nor U14060 (N_14060,N_13927,N_13998);
xnor U14061 (N_14061,N_13937,N_13888);
and U14062 (N_14062,N_13906,N_13822);
nand U14063 (N_14063,N_13957,N_13895);
and U14064 (N_14064,N_13940,N_13873);
and U14065 (N_14065,N_13993,N_13867);
xnor U14066 (N_14066,N_13965,N_13853);
xnor U14067 (N_14067,N_13840,N_13854);
nand U14068 (N_14068,N_13892,N_13819);
and U14069 (N_14069,N_13889,N_13970);
nor U14070 (N_14070,N_13878,N_13931);
xnor U14071 (N_14071,N_13829,N_13934);
nor U14072 (N_14072,N_13887,N_13823);
nand U14073 (N_14073,N_13844,N_13868);
nor U14074 (N_14074,N_13952,N_13827);
nor U14075 (N_14075,N_13969,N_13938);
nand U14076 (N_14076,N_13901,N_13818);
nand U14077 (N_14077,N_13804,N_13824);
nor U14078 (N_14078,N_13983,N_13995);
or U14079 (N_14079,N_13979,N_13820);
nor U14080 (N_14080,N_13825,N_13967);
nand U14081 (N_14081,N_13922,N_13855);
xnor U14082 (N_14082,N_13956,N_13834);
nor U14083 (N_14083,N_13885,N_13896);
or U14084 (N_14084,N_13851,N_13915);
nand U14085 (N_14085,N_13897,N_13945);
or U14086 (N_14086,N_13932,N_13812);
or U14087 (N_14087,N_13911,N_13994);
nand U14088 (N_14088,N_13923,N_13974);
nand U14089 (N_14089,N_13883,N_13999);
nand U14090 (N_14090,N_13944,N_13869);
xnor U14091 (N_14091,N_13890,N_13949);
nor U14092 (N_14092,N_13968,N_13875);
nand U14093 (N_14093,N_13816,N_13987);
or U14094 (N_14094,N_13837,N_13966);
or U14095 (N_14095,N_13917,N_13860);
or U14096 (N_14096,N_13980,N_13903);
and U14097 (N_14097,N_13971,N_13941);
nor U14098 (N_14098,N_13912,N_13996);
nor U14099 (N_14099,N_13948,N_13894);
nor U14100 (N_14100,N_13862,N_13873);
or U14101 (N_14101,N_13938,N_13892);
and U14102 (N_14102,N_13800,N_13862);
xnor U14103 (N_14103,N_13888,N_13974);
nor U14104 (N_14104,N_13838,N_13827);
nand U14105 (N_14105,N_13937,N_13966);
and U14106 (N_14106,N_13912,N_13863);
nor U14107 (N_14107,N_13955,N_13925);
and U14108 (N_14108,N_13942,N_13844);
nand U14109 (N_14109,N_13982,N_13801);
or U14110 (N_14110,N_13922,N_13987);
and U14111 (N_14111,N_13923,N_13878);
xor U14112 (N_14112,N_13803,N_13887);
xnor U14113 (N_14113,N_13884,N_13962);
nor U14114 (N_14114,N_13913,N_13958);
nand U14115 (N_14115,N_13997,N_13923);
and U14116 (N_14116,N_13884,N_13973);
or U14117 (N_14117,N_13852,N_13945);
or U14118 (N_14118,N_13824,N_13802);
or U14119 (N_14119,N_13859,N_13819);
xor U14120 (N_14120,N_13941,N_13819);
or U14121 (N_14121,N_13895,N_13882);
xor U14122 (N_14122,N_13857,N_13939);
or U14123 (N_14123,N_13837,N_13950);
xor U14124 (N_14124,N_13970,N_13842);
nand U14125 (N_14125,N_13890,N_13858);
and U14126 (N_14126,N_13921,N_13856);
nand U14127 (N_14127,N_13916,N_13864);
xnor U14128 (N_14128,N_13837,N_13838);
nand U14129 (N_14129,N_13977,N_13879);
and U14130 (N_14130,N_13878,N_13872);
and U14131 (N_14131,N_13845,N_13866);
or U14132 (N_14132,N_13873,N_13842);
or U14133 (N_14133,N_13933,N_13822);
xor U14134 (N_14134,N_13881,N_13918);
and U14135 (N_14135,N_13888,N_13876);
and U14136 (N_14136,N_13941,N_13866);
or U14137 (N_14137,N_13982,N_13981);
nand U14138 (N_14138,N_13980,N_13825);
and U14139 (N_14139,N_13990,N_13944);
nand U14140 (N_14140,N_13914,N_13926);
xor U14141 (N_14141,N_13951,N_13821);
nor U14142 (N_14142,N_13943,N_13856);
or U14143 (N_14143,N_13815,N_13897);
nand U14144 (N_14144,N_13901,N_13989);
and U14145 (N_14145,N_13906,N_13800);
and U14146 (N_14146,N_13883,N_13946);
or U14147 (N_14147,N_13956,N_13962);
nor U14148 (N_14148,N_13922,N_13865);
nor U14149 (N_14149,N_13809,N_13951);
and U14150 (N_14150,N_13969,N_13944);
xor U14151 (N_14151,N_13888,N_13816);
nor U14152 (N_14152,N_13993,N_13953);
nor U14153 (N_14153,N_13840,N_13828);
nor U14154 (N_14154,N_13946,N_13869);
nand U14155 (N_14155,N_13880,N_13871);
nand U14156 (N_14156,N_13986,N_13861);
nand U14157 (N_14157,N_13892,N_13840);
nand U14158 (N_14158,N_13914,N_13843);
xor U14159 (N_14159,N_13953,N_13933);
xnor U14160 (N_14160,N_13921,N_13908);
nand U14161 (N_14161,N_13944,N_13932);
and U14162 (N_14162,N_13994,N_13802);
nor U14163 (N_14163,N_13819,N_13855);
or U14164 (N_14164,N_13813,N_13925);
or U14165 (N_14165,N_13826,N_13802);
and U14166 (N_14166,N_13866,N_13900);
or U14167 (N_14167,N_13907,N_13820);
and U14168 (N_14168,N_13816,N_13957);
nand U14169 (N_14169,N_13874,N_13934);
nor U14170 (N_14170,N_13878,N_13845);
xor U14171 (N_14171,N_13850,N_13810);
nand U14172 (N_14172,N_13941,N_13999);
or U14173 (N_14173,N_13924,N_13892);
nor U14174 (N_14174,N_13976,N_13972);
nand U14175 (N_14175,N_13928,N_13922);
nor U14176 (N_14176,N_13840,N_13803);
xor U14177 (N_14177,N_13976,N_13857);
and U14178 (N_14178,N_13998,N_13905);
or U14179 (N_14179,N_13890,N_13951);
or U14180 (N_14180,N_13845,N_13921);
and U14181 (N_14181,N_13893,N_13921);
xnor U14182 (N_14182,N_13979,N_13830);
xor U14183 (N_14183,N_13901,N_13841);
and U14184 (N_14184,N_13935,N_13845);
nand U14185 (N_14185,N_13934,N_13930);
or U14186 (N_14186,N_13944,N_13827);
and U14187 (N_14187,N_13865,N_13884);
nor U14188 (N_14188,N_13893,N_13830);
and U14189 (N_14189,N_13957,N_13891);
nor U14190 (N_14190,N_13999,N_13820);
and U14191 (N_14191,N_13895,N_13828);
nor U14192 (N_14192,N_13838,N_13834);
nand U14193 (N_14193,N_13987,N_13843);
xor U14194 (N_14194,N_13898,N_13959);
nand U14195 (N_14195,N_13814,N_13866);
or U14196 (N_14196,N_13900,N_13882);
xor U14197 (N_14197,N_13973,N_13945);
and U14198 (N_14198,N_13921,N_13972);
xor U14199 (N_14199,N_13806,N_13917);
nand U14200 (N_14200,N_14192,N_14063);
or U14201 (N_14201,N_14036,N_14178);
and U14202 (N_14202,N_14188,N_14049);
xnor U14203 (N_14203,N_14181,N_14155);
or U14204 (N_14204,N_14170,N_14125);
nand U14205 (N_14205,N_14052,N_14016);
nand U14206 (N_14206,N_14007,N_14120);
and U14207 (N_14207,N_14103,N_14090);
nor U14208 (N_14208,N_14106,N_14080);
xor U14209 (N_14209,N_14145,N_14166);
nor U14210 (N_14210,N_14194,N_14129);
or U14211 (N_14211,N_14061,N_14083);
nor U14212 (N_14212,N_14072,N_14164);
nor U14213 (N_14213,N_14025,N_14035);
and U14214 (N_14214,N_14193,N_14002);
nand U14215 (N_14215,N_14183,N_14086);
nand U14216 (N_14216,N_14173,N_14043);
or U14217 (N_14217,N_14111,N_14009);
nor U14218 (N_14218,N_14059,N_14184);
xor U14219 (N_14219,N_14045,N_14033);
nand U14220 (N_14220,N_14051,N_14134);
nand U14221 (N_14221,N_14130,N_14162);
or U14222 (N_14222,N_14068,N_14180);
and U14223 (N_14223,N_14199,N_14136);
xnor U14224 (N_14224,N_14149,N_14058);
and U14225 (N_14225,N_14095,N_14048);
xnor U14226 (N_14226,N_14022,N_14110);
and U14227 (N_14227,N_14087,N_14138);
and U14228 (N_14228,N_14024,N_14070);
and U14229 (N_14229,N_14042,N_14175);
nor U14230 (N_14230,N_14000,N_14031);
and U14231 (N_14231,N_14137,N_14069);
and U14232 (N_14232,N_14056,N_14084);
nor U14233 (N_14233,N_14053,N_14179);
nor U14234 (N_14234,N_14018,N_14196);
nand U14235 (N_14235,N_14006,N_14112);
xor U14236 (N_14236,N_14122,N_14046);
nand U14237 (N_14237,N_14143,N_14027);
and U14238 (N_14238,N_14158,N_14146);
nand U14239 (N_14239,N_14014,N_14060);
nor U14240 (N_14240,N_14148,N_14077);
nand U14241 (N_14241,N_14156,N_14012);
nand U14242 (N_14242,N_14161,N_14133);
nor U14243 (N_14243,N_14144,N_14139);
nand U14244 (N_14244,N_14029,N_14159);
and U14245 (N_14245,N_14182,N_14115);
or U14246 (N_14246,N_14047,N_14174);
xor U14247 (N_14247,N_14116,N_14050);
nor U14248 (N_14248,N_14123,N_14147);
xnor U14249 (N_14249,N_14001,N_14186);
nor U14250 (N_14250,N_14019,N_14093);
and U14251 (N_14251,N_14150,N_14190);
nand U14252 (N_14252,N_14008,N_14135);
or U14253 (N_14253,N_14023,N_14055);
xor U14254 (N_14254,N_14131,N_14079);
xnor U14255 (N_14255,N_14028,N_14065);
or U14256 (N_14256,N_14064,N_14071);
nor U14257 (N_14257,N_14010,N_14185);
nand U14258 (N_14258,N_14054,N_14141);
nor U14259 (N_14259,N_14039,N_14118);
or U14260 (N_14260,N_14066,N_14020);
or U14261 (N_14261,N_14003,N_14021);
and U14262 (N_14262,N_14100,N_14198);
nand U14263 (N_14263,N_14140,N_14108);
or U14264 (N_14264,N_14096,N_14104);
and U14265 (N_14265,N_14074,N_14169);
nand U14266 (N_14266,N_14126,N_14017);
xor U14267 (N_14267,N_14099,N_14041);
nand U14268 (N_14268,N_14128,N_14105);
xor U14269 (N_14269,N_14189,N_14085);
or U14270 (N_14270,N_14114,N_14073);
xnor U14271 (N_14271,N_14132,N_14153);
nor U14272 (N_14272,N_14078,N_14030);
or U14273 (N_14273,N_14040,N_14152);
nor U14274 (N_14274,N_14088,N_14113);
nor U14275 (N_14275,N_14015,N_14127);
nor U14276 (N_14276,N_14005,N_14195);
nand U14277 (N_14277,N_14076,N_14075);
xor U14278 (N_14278,N_14197,N_14013);
and U14279 (N_14279,N_14176,N_14168);
nand U14280 (N_14280,N_14081,N_14092);
nand U14281 (N_14281,N_14067,N_14163);
xor U14282 (N_14282,N_14160,N_14187);
nor U14283 (N_14283,N_14098,N_14034);
nand U14284 (N_14284,N_14121,N_14057);
and U14285 (N_14285,N_14165,N_14171);
or U14286 (N_14286,N_14037,N_14091);
or U14287 (N_14287,N_14142,N_14004);
nor U14288 (N_14288,N_14167,N_14107);
xor U14289 (N_14289,N_14154,N_14097);
nor U14290 (N_14290,N_14177,N_14032);
and U14291 (N_14291,N_14026,N_14062);
and U14292 (N_14292,N_14102,N_14011);
and U14293 (N_14293,N_14157,N_14109);
and U14294 (N_14294,N_14089,N_14124);
nand U14295 (N_14295,N_14172,N_14038);
or U14296 (N_14296,N_14101,N_14094);
and U14297 (N_14297,N_14082,N_14119);
nand U14298 (N_14298,N_14117,N_14191);
or U14299 (N_14299,N_14044,N_14151);
and U14300 (N_14300,N_14068,N_14191);
or U14301 (N_14301,N_14053,N_14122);
and U14302 (N_14302,N_14149,N_14128);
xnor U14303 (N_14303,N_14034,N_14158);
nor U14304 (N_14304,N_14133,N_14009);
nand U14305 (N_14305,N_14092,N_14058);
xnor U14306 (N_14306,N_14075,N_14017);
or U14307 (N_14307,N_14168,N_14033);
nor U14308 (N_14308,N_14175,N_14074);
xor U14309 (N_14309,N_14054,N_14120);
and U14310 (N_14310,N_14146,N_14180);
nor U14311 (N_14311,N_14090,N_14181);
nand U14312 (N_14312,N_14100,N_14093);
nor U14313 (N_14313,N_14079,N_14127);
or U14314 (N_14314,N_14151,N_14124);
or U14315 (N_14315,N_14057,N_14104);
nor U14316 (N_14316,N_14121,N_14026);
nor U14317 (N_14317,N_14008,N_14088);
xor U14318 (N_14318,N_14071,N_14031);
nand U14319 (N_14319,N_14165,N_14055);
nand U14320 (N_14320,N_14156,N_14034);
nor U14321 (N_14321,N_14060,N_14182);
or U14322 (N_14322,N_14163,N_14117);
nor U14323 (N_14323,N_14016,N_14188);
xnor U14324 (N_14324,N_14178,N_14184);
nor U14325 (N_14325,N_14130,N_14020);
xnor U14326 (N_14326,N_14019,N_14006);
xor U14327 (N_14327,N_14086,N_14079);
nand U14328 (N_14328,N_14097,N_14191);
or U14329 (N_14329,N_14198,N_14090);
and U14330 (N_14330,N_14063,N_14089);
nand U14331 (N_14331,N_14075,N_14157);
nand U14332 (N_14332,N_14104,N_14048);
nor U14333 (N_14333,N_14159,N_14131);
nor U14334 (N_14334,N_14091,N_14032);
nand U14335 (N_14335,N_14051,N_14172);
and U14336 (N_14336,N_14045,N_14136);
nor U14337 (N_14337,N_14141,N_14081);
nor U14338 (N_14338,N_14066,N_14002);
and U14339 (N_14339,N_14041,N_14032);
nand U14340 (N_14340,N_14140,N_14044);
xnor U14341 (N_14341,N_14061,N_14198);
nor U14342 (N_14342,N_14035,N_14049);
xnor U14343 (N_14343,N_14011,N_14041);
or U14344 (N_14344,N_14116,N_14068);
xor U14345 (N_14345,N_14073,N_14120);
and U14346 (N_14346,N_14191,N_14165);
nand U14347 (N_14347,N_14121,N_14053);
nand U14348 (N_14348,N_14172,N_14072);
and U14349 (N_14349,N_14102,N_14045);
or U14350 (N_14350,N_14136,N_14038);
and U14351 (N_14351,N_14145,N_14101);
and U14352 (N_14352,N_14018,N_14015);
nor U14353 (N_14353,N_14042,N_14163);
and U14354 (N_14354,N_14020,N_14072);
and U14355 (N_14355,N_14086,N_14042);
xnor U14356 (N_14356,N_14147,N_14114);
and U14357 (N_14357,N_14037,N_14143);
xnor U14358 (N_14358,N_14183,N_14187);
nor U14359 (N_14359,N_14093,N_14084);
nor U14360 (N_14360,N_14197,N_14007);
xnor U14361 (N_14361,N_14106,N_14023);
and U14362 (N_14362,N_14171,N_14018);
or U14363 (N_14363,N_14012,N_14153);
xor U14364 (N_14364,N_14026,N_14097);
nor U14365 (N_14365,N_14052,N_14018);
and U14366 (N_14366,N_14139,N_14015);
xnor U14367 (N_14367,N_14079,N_14173);
nand U14368 (N_14368,N_14036,N_14129);
nand U14369 (N_14369,N_14095,N_14074);
xor U14370 (N_14370,N_14054,N_14133);
xnor U14371 (N_14371,N_14066,N_14190);
or U14372 (N_14372,N_14088,N_14131);
nand U14373 (N_14373,N_14072,N_14032);
nand U14374 (N_14374,N_14187,N_14066);
or U14375 (N_14375,N_14061,N_14107);
nor U14376 (N_14376,N_14152,N_14184);
nor U14377 (N_14377,N_14162,N_14048);
nand U14378 (N_14378,N_14036,N_14167);
xor U14379 (N_14379,N_14075,N_14025);
xor U14380 (N_14380,N_14159,N_14067);
and U14381 (N_14381,N_14175,N_14022);
nand U14382 (N_14382,N_14079,N_14054);
xor U14383 (N_14383,N_14101,N_14158);
nand U14384 (N_14384,N_14000,N_14061);
nor U14385 (N_14385,N_14007,N_14196);
or U14386 (N_14386,N_14150,N_14144);
nand U14387 (N_14387,N_14115,N_14075);
nor U14388 (N_14388,N_14064,N_14188);
nand U14389 (N_14389,N_14153,N_14188);
nor U14390 (N_14390,N_14080,N_14034);
nor U14391 (N_14391,N_14085,N_14029);
or U14392 (N_14392,N_14062,N_14066);
or U14393 (N_14393,N_14098,N_14104);
nor U14394 (N_14394,N_14100,N_14066);
nand U14395 (N_14395,N_14036,N_14091);
xor U14396 (N_14396,N_14038,N_14039);
or U14397 (N_14397,N_14061,N_14112);
nor U14398 (N_14398,N_14144,N_14019);
xnor U14399 (N_14399,N_14153,N_14187);
xor U14400 (N_14400,N_14391,N_14309);
and U14401 (N_14401,N_14296,N_14351);
nor U14402 (N_14402,N_14273,N_14256);
nor U14403 (N_14403,N_14308,N_14353);
and U14404 (N_14404,N_14320,N_14349);
nand U14405 (N_14405,N_14370,N_14222);
nand U14406 (N_14406,N_14377,N_14281);
or U14407 (N_14407,N_14361,N_14399);
nor U14408 (N_14408,N_14386,N_14364);
nor U14409 (N_14409,N_14328,N_14396);
xor U14410 (N_14410,N_14250,N_14257);
nand U14411 (N_14411,N_14333,N_14231);
nand U14412 (N_14412,N_14219,N_14342);
nor U14413 (N_14413,N_14288,N_14225);
and U14414 (N_14414,N_14265,N_14242);
or U14415 (N_14415,N_14236,N_14372);
xnor U14416 (N_14416,N_14336,N_14346);
nor U14417 (N_14417,N_14326,N_14340);
xnor U14418 (N_14418,N_14247,N_14259);
xnor U14419 (N_14419,N_14356,N_14376);
and U14420 (N_14420,N_14392,N_14316);
or U14421 (N_14421,N_14382,N_14384);
and U14422 (N_14422,N_14365,N_14380);
nor U14423 (N_14423,N_14323,N_14321);
or U14424 (N_14424,N_14211,N_14345);
nor U14425 (N_14425,N_14210,N_14379);
nand U14426 (N_14426,N_14385,N_14358);
and U14427 (N_14427,N_14318,N_14350);
and U14428 (N_14428,N_14233,N_14387);
nor U14429 (N_14429,N_14212,N_14268);
nand U14430 (N_14430,N_14357,N_14334);
and U14431 (N_14431,N_14267,N_14369);
nand U14432 (N_14432,N_14390,N_14279);
nand U14433 (N_14433,N_14398,N_14341);
or U14434 (N_14434,N_14294,N_14374);
xnor U14435 (N_14435,N_14383,N_14324);
xnor U14436 (N_14436,N_14304,N_14389);
and U14437 (N_14437,N_14261,N_14264);
and U14438 (N_14438,N_14395,N_14319);
nand U14439 (N_14439,N_14297,N_14293);
and U14440 (N_14440,N_14315,N_14215);
nor U14441 (N_14441,N_14289,N_14307);
nor U14442 (N_14442,N_14254,N_14394);
xor U14443 (N_14443,N_14317,N_14213);
nor U14444 (N_14444,N_14343,N_14295);
nand U14445 (N_14445,N_14274,N_14246);
and U14446 (N_14446,N_14241,N_14388);
or U14447 (N_14447,N_14339,N_14371);
nand U14448 (N_14448,N_14287,N_14301);
and U14449 (N_14449,N_14255,N_14214);
nand U14450 (N_14450,N_14276,N_14292);
or U14451 (N_14451,N_14206,N_14227);
xor U14452 (N_14452,N_14217,N_14359);
and U14453 (N_14453,N_14205,N_14378);
or U14454 (N_14454,N_14278,N_14362);
xor U14455 (N_14455,N_14305,N_14347);
nand U14456 (N_14456,N_14203,N_14310);
or U14457 (N_14457,N_14332,N_14271);
or U14458 (N_14458,N_14237,N_14303);
xnor U14459 (N_14459,N_14260,N_14245);
xor U14460 (N_14460,N_14313,N_14258);
xor U14461 (N_14461,N_14204,N_14200);
or U14462 (N_14462,N_14327,N_14216);
nor U14463 (N_14463,N_14286,N_14280);
or U14464 (N_14464,N_14285,N_14201);
nand U14465 (N_14465,N_14243,N_14235);
or U14466 (N_14466,N_14290,N_14240);
nor U14467 (N_14467,N_14300,N_14275);
and U14468 (N_14468,N_14311,N_14251);
and U14469 (N_14469,N_14299,N_14352);
and U14470 (N_14470,N_14375,N_14329);
and U14471 (N_14471,N_14253,N_14291);
nor U14472 (N_14472,N_14248,N_14277);
and U14473 (N_14473,N_14244,N_14238);
nand U14474 (N_14474,N_14220,N_14330);
nand U14475 (N_14475,N_14348,N_14335);
and U14476 (N_14476,N_14397,N_14223);
nand U14477 (N_14477,N_14226,N_14354);
or U14478 (N_14478,N_14234,N_14393);
nor U14479 (N_14479,N_14381,N_14331);
nand U14480 (N_14480,N_14366,N_14224);
and U14481 (N_14481,N_14263,N_14252);
nand U14482 (N_14482,N_14269,N_14272);
xnor U14483 (N_14483,N_14282,N_14221);
and U14484 (N_14484,N_14266,N_14228);
nor U14485 (N_14485,N_14283,N_14338);
and U14486 (N_14486,N_14367,N_14208);
xor U14487 (N_14487,N_14306,N_14363);
nor U14488 (N_14488,N_14360,N_14218);
nor U14489 (N_14489,N_14325,N_14262);
xor U14490 (N_14490,N_14202,N_14322);
nor U14491 (N_14491,N_14229,N_14302);
nor U14492 (N_14492,N_14249,N_14344);
or U14493 (N_14493,N_14314,N_14232);
and U14494 (N_14494,N_14312,N_14230);
and U14495 (N_14495,N_14368,N_14284);
xnor U14496 (N_14496,N_14239,N_14270);
nand U14497 (N_14497,N_14355,N_14337);
nor U14498 (N_14498,N_14209,N_14207);
xor U14499 (N_14499,N_14298,N_14373);
and U14500 (N_14500,N_14250,N_14255);
and U14501 (N_14501,N_14383,N_14208);
or U14502 (N_14502,N_14267,N_14341);
nand U14503 (N_14503,N_14391,N_14296);
nand U14504 (N_14504,N_14274,N_14348);
nor U14505 (N_14505,N_14240,N_14344);
nand U14506 (N_14506,N_14374,N_14364);
and U14507 (N_14507,N_14238,N_14253);
nor U14508 (N_14508,N_14227,N_14334);
or U14509 (N_14509,N_14328,N_14399);
or U14510 (N_14510,N_14398,N_14369);
xor U14511 (N_14511,N_14268,N_14373);
nor U14512 (N_14512,N_14347,N_14258);
or U14513 (N_14513,N_14235,N_14257);
or U14514 (N_14514,N_14398,N_14318);
nand U14515 (N_14515,N_14247,N_14280);
nand U14516 (N_14516,N_14260,N_14271);
nor U14517 (N_14517,N_14209,N_14298);
and U14518 (N_14518,N_14324,N_14291);
nand U14519 (N_14519,N_14381,N_14317);
or U14520 (N_14520,N_14279,N_14367);
and U14521 (N_14521,N_14286,N_14257);
and U14522 (N_14522,N_14329,N_14326);
and U14523 (N_14523,N_14229,N_14379);
nand U14524 (N_14524,N_14286,N_14304);
nor U14525 (N_14525,N_14300,N_14315);
nor U14526 (N_14526,N_14264,N_14326);
nor U14527 (N_14527,N_14317,N_14395);
nor U14528 (N_14528,N_14304,N_14339);
or U14529 (N_14529,N_14387,N_14320);
or U14530 (N_14530,N_14393,N_14359);
nand U14531 (N_14531,N_14385,N_14270);
nand U14532 (N_14532,N_14265,N_14355);
or U14533 (N_14533,N_14241,N_14281);
and U14534 (N_14534,N_14240,N_14397);
nand U14535 (N_14535,N_14272,N_14366);
and U14536 (N_14536,N_14201,N_14397);
and U14537 (N_14537,N_14204,N_14270);
xor U14538 (N_14538,N_14376,N_14359);
and U14539 (N_14539,N_14216,N_14294);
nor U14540 (N_14540,N_14224,N_14268);
nand U14541 (N_14541,N_14231,N_14385);
nor U14542 (N_14542,N_14226,N_14328);
nor U14543 (N_14543,N_14245,N_14288);
xor U14544 (N_14544,N_14361,N_14358);
and U14545 (N_14545,N_14378,N_14389);
nor U14546 (N_14546,N_14326,N_14303);
nand U14547 (N_14547,N_14369,N_14246);
and U14548 (N_14548,N_14230,N_14288);
nand U14549 (N_14549,N_14339,N_14378);
xnor U14550 (N_14550,N_14376,N_14393);
and U14551 (N_14551,N_14324,N_14246);
and U14552 (N_14552,N_14338,N_14336);
xnor U14553 (N_14553,N_14225,N_14305);
nand U14554 (N_14554,N_14226,N_14344);
and U14555 (N_14555,N_14362,N_14265);
nor U14556 (N_14556,N_14276,N_14214);
nand U14557 (N_14557,N_14366,N_14319);
nand U14558 (N_14558,N_14313,N_14255);
nand U14559 (N_14559,N_14397,N_14215);
and U14560 (N_14560,N_14238,N_14313);
or U14561 (N_14561,N_14256,N_14355);
nand U14562 (N_14562,N_14295,N_14211);
nor U14563 (N_14563,N_14319,N_14307);
nand U14564 (N_14564,N_14245,N_14213);
and U14565 (N_14565,N_14388,N_14292);
and U14566 (N_14566,N_14335,N_14281);
nand U14567 (N_14567,N_14260,N_14296);
nor U14568 (N_14568,N_14318,N_14385);
xnor U14569 (N_14569,N_14253,N_14337);
xor U14570 (N_14570,N_14217,N_14251);
xnor U14571 (N_14571,N_14305,N_14363);
nor U14572 (N_14572,N_14369,N_14250);
nor U14573 (N_14573,N_14379,N_14237);
xor U14574 (N_14574,N_14320,N_14343);
nor U14575 (N_14575,N_14227,N_14384);
and U14576 (N_14576,N_14235,N_14374);
or U14577 (N_14577,N_14229,N_14324);
xnor U14578 (N_14578,N_14337,N_14321);
and U14579 (N_14579,N_14276,N_14259);
xnor U14580 (N_14580,N_14345,N_14239);
and U14581 (N_14581,N_14262,N_14276);
nand U14582 (N_14582,N_14282,N_14335);
nor U14583 (N_14583,N_14359,N_14333);
or U14584 (N_14584,N_14343,N_14261);
xor U14585 (N_14585,N_14221,N_14335);
and U14586 (N_14586,N_14240,N_14334);
nor U14587 (N_14587,N_14270,N_14272);
or U14588 (N_14588,N_14229,N_14265);
and U14589 (N_14589,N_14333,N_14256);
nor U14590 (N_14590,N_14308,N_14376);
xnor U14591 (N_14591,N_14326,N_14347);
xor U14592 (N_14592,N_14235,N_14393);
nand U14593 (N_14593,N_14278,N_14276);
nor U14594 (N_14594,N_14385,N_14254);
nor U14595 (N_14595,N_14376,N_14378);
and U14596 (N_14596,N_14237,N_14261);
and U14597 (N_14597,N_14222,N_14331);
nand U14598 (N_14598,N_14348,N_14211);
nand U14599 (N_14599,N_14365,N_14358);
or U14600 (N_14600,N_14548,N_14460);
or U14601 (N_14601,N_14493,N_14544);
and U14602 (N_14602,N_14424,N_14547);
xnor U14603 (N_14603,N_14546,N_14496);
and U14604 (N_14604,N_14484,N_14483);
xnor U14605 (N_14605,N_14545,N_14419);
or U14606 (N_14606,N_14442,N_14420);
and U14607 (N_14607,N_14423,N_14551);
or U14608 (N_14608,N_14401,N_14467);
or U14609 (N_14609,N_14566,N_14531);
nor U14610 (N_14610,N_14437,N_14499);
nor U14611 (N_14611,N_14524,N_14425);
xor U14612 (N_14612,N_14511,N_14408);
or U14613 (N_14613,N_14510,N_14446);
and U14614 (N_14614,N_14403,N_14457);
nand U14615 (N_14615,N_14514,N_14575);
xor U14616 (N_14616,N_14404,N_14461);
and U14617 (N_14617,N_14445,N_14549);
xor U14618 (N_14618,N_14422,N_14502);
nor U14619 (N_14619,N_14414,N_14542);
nor U14620 (N_14620,N_14488,N_14491);
xnor U14621 (N_14621,N_14468,N_14498);
or U14622 (N_14622,N_14432,N_14526);
xor U14623 (N_14623,N_14463,N_14417);
nor U14624 (N_14624,N_14582,N_14465);
or U14625 (N_14625,N_14456,N_14504);
nand U14626 (N_14626,N_14589,N_14556);
nor U14627 (N_14627,N_14561,N_14435);
nand U14628 (N_14628,N_14473,N_14434);
or U14629 (N_14629,N_14519,N_14409);
nor U14630 (N_14630,N_14478,N_14454);
nor U14631 (N_14631,N_14477,N_14443);
nor U14632 (N_14632,N_14588,N_14426);
or U14633 (N_14633,N_14453,N_14482);
xor U14634 (N_14634,N_14540,N_14402);
and U14635 (N_14635,N_14428,N_14528);
xor U14636 (N_14636,N_14508,N_14438);
and U14637 (N_14637,N_14449,N_14565);
or U14638 (N_14638,N_14552,N_14523);
nor U14639 (N_14639,N_14427,N_14598);
and U14640 (N_14640,N_14572,N_14543);
xnor U14641 (N_14641,N_14406,N_14571);
or U14642 (N_14642,N_14520,N_14480);
and U14643 (N_14643,N_14574,N_14490);
or U14644 (N_14644,N_14532,N_14489);
or U14645 (N_14645,N_14470,N_14579);
xnor U14646 (N_14646,N_14501,N_14407);
and U14647 (N_14647,N_14464,N_14593);
and U14648 (N_14648,N_14479,N_14517);
xnor U14649 (N_14649,N_14462,N_14440);
and U14650 (N_14650,N_14459,N_14513);
nand U14651 (N_14651,N_14557,N_14573);
nor U14652 (N_14652,N_14530,N_14455);
nor U14653 (N_14653,N_14411,N_14539);
xor U14654 (N_14654,N_14487,N_14469);
nor U14655 (N_14655,N_14592,N_14421);
nand U14656 (N_14656,N_14558,N_14444);
nand U14657 (N_14657,N_14472,N_14591);
xor U14658 (N_14658,N_14481,N_14577);
or U14659 (N_14659,N_14584,N_14509);
and U14660 (N_14660,N_14599,N_14553);
xnor U14661 (N_14661,N_14537,N_14567);
nand U14662 (N_14662,N_14418,N_14535);
nand U14663 (N_14663,N_14431,N_14521);
nor U14664 (N_14664,N_14405,N_14503);
or U14665 (N_14665,N_14564,N_14554);
nand U14666 (N_14666,N_14452,N_14415);
or U14667 (N_14667,N_14585,N_14466);
or U14668 (N_14668,N_14448,N_14534);
nor U14669 (N_14669,N_14512,N_14538);
xor U14670 (N_14670,N_14507,N_14578);
nor U14671 (N_14671,N_14447,N_14580);
xnor U14672 (N_14672,N_14525,N_14590);
and U14673 (N_14673,N_14515,N_14586);
or U14674 (N_14674,N_14476,N_14536);
nand U14675 (N_14675,N_14568,N_14533);
xnor U14676 (N_14676,N_14550,N_14400);
xnor U14677 (N_14677,N_14416,N_14560);
xnor U14678 (N_14678,N_14505,N_14451);
nor U14679 (N_14679,N_14410,N_14569);
xnor U14680 (N_14680,N_14581,N_14595);
nor U14681 (N_14681,N_14475,N_14518);
and U14682 (N_14682,N_14522,N_14506);
nor U14683 (N_14683,N_14494,N_14559);
xnor U14684 (N_14684,N_14563,N_14555);
or U14685 (N_14685,N_14576,N_14497);
and U14686 (N_14686,N_14430,N_14433);
xor U14687 (N_14687,N_14570,N_14474);
xor U14688 (N_14688,N_14429,N_14527);
or U14689 (N_14689,N_14583,N_14597);
or U14690 (N_14690,N_14500,N_14485);
xor U14691 (N_14691,N_14450,N_14516);
nor U14692 (N_14692,N_14412,N_14486);
nand U14693 (N_14693,N_14413,N_14596);
nor U14694 (N_14694,N_14562,N_14541);
nand U14695 (N_14695,N_14439,N_14594);
nand U14696 (N_14696,N_14587,N_14495);
xor U14697 (N_14697,N_14529,N_14441);
and U14698 (N_14698,N_14471,N_14436);
nand U14699 (N_14699,N_14492,N_14458);
and U14700 (N_14700,N_14572,N_14435);
xor U14701 (N_14701,N_14416,N_14540);
nand U14702 (N_14702,N_14564,N_14404);
nor U14703 (N_14703,N_14496,N_14521);
and U14704 (N_14704,N_14556,N_14434);
and U14705 (N_14705,N_14458,N_14549);
nor U14706 (N_14706,N_14536,N_14490);
and U14707 (N_14707,N_14598,N_14534);
and U14708 (N_14708,N_14469,N_14496);
xor U14709 (N_14709,N_14405,N_14514);
or U14710 (N_14710,N_14429,N_14580);
or U14711 (N_14711,N_14453,N_14558);
or U14712 (N_14712,N_14587,N_14411);
and U14713 (N_14713,N_14480,N_14501);
or U14714 (N_14714,N_14528,N_14490);
or U14715 (N_14715,N_14508,N_14568);
xnor U14716 (N_14716,N_14505,N_14538);
nor U14717 (N_14717,N_14596,N_14586);
or U14718 (N_14718,N_14501,N_14599);
nand U14719 (N_14719,N_14422,N_14566);
nand U14720 (N_14720,N_14530,N_14563);
or U14721 (N_14721,N_14528,N_14569);
nand U14722 (N_14722,N_14519,N_14435);
or U14723 (N_14723,N_14555,N_14530);
or U14724 (N_14724,N_14546,N_14563);
xor U14725 (N_14725,N_14596,N_14497);
or U14726 (N_14726,N_14589,N_14499);
nor U14727 (N_14727,N_14582,N_14516);
nor U14728 (N_14728,N_14472,N_14516);
xor U14729 (N_14729,N_14433,N_14530);
or U14730 (N_14730,N_14459,N_14417);
and U14731 (N_14731,N_14522,N_14536);
or U14732 (N_14732,N_14571,N_14430);
nor U14733 (N_14733,N_14468,N_14510);
nor U14734 (N_14734,N_14417,N_14426);
nor U14735 (N_14735,N_14493,N_14480);
and U14736 (N_14736,N_14485,N_14431);
and U14737 (N_14737,N_14512,N_14503);
nand U14738 (N_14738,N_14560,N_14442);
or U14739 (N_14739,N_14576,N_14533);
and U14740 (N_14740,N_14403,N_14564);
nor U14741 (N_14741,N_14533,N_14483);
and U14742 (N_14742,N_14418,N_14482);
and U14743 (N_14743,N_14540,N_14583);
xor U14744 (N_14744,N_14458,N_14461);
nand U14745 (N_14745,N_14509,N_14516);
xnor U14746 (N_14746,N_14434,N_14594);
or U14747 (N_14747,N_14476,N_14498);
and U14748 (N_14748,N_14546,N_14457);
nor U14749 (N_14749,N_14594,N_14555);
nand U14750 (N_14750,N_14500,N_14471);
nand U14751 (N_14751,N_14565,N_14482);
or U14752 (N_14752,N_14467,N_14420);
and U14753 (N_14753,N_14576,N_14557);
nand U14754 (N_14754,N_14531,N_14580);
or U14755 (N_14755,N_14539,N_14501);
or U14756 (N_14756,N_14491,N_14565);
nand U14757 (N_14757,N_14587,N_14577);
nand U14758 (N_14758,N_14559,N_14504);
xor U14759 (N_14759,N_14410,N_14579);
or U14760 (N_14760,N_14411,N_14468);
or U14761 (N_14761,N_14537,N_14461);
nor U14762 (N_14762,N_14571,N_14447);
or U14763 (N_14763,N_14574,N_14529);
nand U14764 (N_14764,N_14558,N_14442);
nand U14765 (N_14765,N_14598,N_14552);
xor U14766 (N_14766,N_14425,N_14484);
nand U14767 (N_14767,N_14586,N_14541);
and U14768 (N_14768,N_14525,N_14541);
or U14769 (N_14769,N_14405,N_14445);
xor U14770 (N_14770,N_14592,N_14532);
or U14771 (N_14771,N_14448,N_14470);
nand U14772 (N_14772,N_14575,N_14587);
or U14773 (N_14773,N_14466,N_14451);
xor U14774 (N_14774,N_14472,N_14491);
or U14775 (N_14775,N_14564,N_14405);
and U14776 (N_14776,N_14435,N_14468);
xor U14777 (N_14777,N_14533,N_14474);
and U14778 (N_14778,N_14537,N_14410);
nand U14779 (N_14779,N_14465,N_14404);
xor U14780 (N_14780,N_14459,N_14440);
nand U14781 (N_14781,N_14451,N_14481);
nor U14782 (N_14782,N_14587,N_14563);
or U14783 (N_14783,N_14448,N_14436);
nand U14784 (N_14784,N_14534,N_14504);
and U14785 (N_14785,N_14499,N_14441);
and U14786 (N_14786,N_14558,N_14433);
nor U14787 (N_14787,N_14458,N_14564);
xor U14788 (N_14788,N_14401,N_14482);
and U14789 (N_14789,N_14565,N_14415);
or U14790 (N_14790,N_14436,N_14555);
and U14791 (N_14791,N_14491,N_14451);
xnor U14792 (N_14792,N_14575,N_14517);
nor U14793 (N_14793,N_14523,N_14415);
xor U14794 (N_14794,N_14440,N_14514);
nor U14795 (N_14795,N_14544,N_14482);
or U14796 (N_14796,N_14483,N_14581);
nor U14797 (N_14797,N_14512,N_14462);
and U14798 (N_14798,N_14566,N_14487);
or U14799 (N_14799,N_14539,N_14569);
and U14800 (N_14800,N_14777,N_14696);
nor U14801 (N_14801,N_14722,N_14609);
nand U14802 (N_14802,N_14607,N_14628);
nor U14803 (N_14803,N_14616,N_14740);
and U14804 (N_14804,N_14752,N_14713);
nor U14805 (N_14805,N_14723,N_14603);
or U14806 (N_14806,N_14701,N_14707);
or U14807 (N_14807,N_14784,N_14756);
xor U14808 (N_14808,N_14738,N_14648);
and U14809 (N_14809,N_14645,N_14759);
nor U14810 (N_14810,N_14695,N_14698);
and U14811 (N_14811,N_14650,N_14733);
and U14812 (N_14812,N_14620,N_14682);
or U14813 (N_14813,N_14769,N_14747);
or U14814 (N_14814,N_14626,N_14797);
and U14815 (N_14815,N_14608,N_14675);
nand U14816 (N_14816,N_14604,N_14680);
and U14817 (N_14817,N_14656,N_14715);
or U14818 (N_14818,N_14765,N_14633);
nor U14819 (N_14819,N_14644,N_14728);
nor U14820 (N_14820,N_14703,N_14766);
or U14821 (N_14821,N_14798,N_14602);
or U14822 (N_14822,N_14767,N_14754);
and U14823 (N_14823,N_14780,N_14643);
nor U14824 (N_14824,N_14658,N_14664);
xnor U14825 (N_14825,N_14711,N_14612);
xnor U14826 (N_14826,N_14625,N_14762);
and U14827 (N_14827,N_14746,N_14716);
nor U14828 (N_14828,N_14743,N_14654);
or U14829 (N_14829,N_14741,N_14727);
nand U14830 (N_14830,N_14630,N_14795);
or U14831 (N_14831,N_14665,N_14773);
and U14832 (N_14832,N_14717,N_14702);
nor U14833 (N_14833,N_14794,N_14788);
and U14834 (N_14834,N_14683,N_14775);
nor U14835 (N_14835,N_14693,N_14779);
and U14836 (N_14836,N_14660,N_14636);
or U14837 (N_14837,N_14774,N_14734);
and U14838 (N_14838,N_14638,N_14708);
nor U14839 (N_14839,N_14611,N_14731);
nand U14840 (N_14840,N_14700,N_14732);
nor U14841 (N_14841,N_14640,N_14686);
or U14842 (N_14842,N_14606,N_14755);
nor U14843 (N_14843,N_14760,N_14748);
nand U14844 (N_14844,N_14689,N_14681);
and U14845 (N_14845,N_14725,N_14624);
or U14846 (N_14846,N_14757,N_14730);
nand U14847 (N_14847,N_14790,N_14618);
xnor U14848 (N_14848,N_14799,N_14676);
nand U14849 (N_14849,N_14623,N_14714);
xor U14850 (N_14850,N_14653,N_14671);
and U14851 (N_14851,N_14615,N_14669);
xnor U14852 (N_14852,N_14685,N_14778);
and U14853 (N_14853,N_14662,N_14646);
nand U14854 (N_14854,N_14786,N_14751);
nor U14855 (N_14855,N_14647,N_14764);
nand U14856 (N_14856,N_14670,N_14758);
or U14857 (N_14857,N_14622,N_14744);
nand U14858 (N_14858,N_14631,N_14635);
xnor U14859 (N_14859,N_14677,N_14694);
nand U14860 (N_14860,N_14627,N_14637);
and U14861 (N_14861,N_14617,N_14783);
and U14862 (N_14862,N_14718,N_14763);
nor U14863 (N_14863,N_14736,N_14642);
nand U14864 (N_14864,N_14737,N_14605);
and U14865 (N_14865,N_14684,N_14668);
or U14866 (N_14866,N_14679,N_14706);
or U14867 (N_14867,N_14651,N_14692);
nor U14868 (N_14868,N_14634,N_14735);
nor U14869 (N_14869,N_14721,N_14657);
xnor U14870 (N_14870,N_14761,N_14771);
nor U14871 (N_14871,N_14782,N_14629);
nor U14872 (N_14872,N_14613,N_14753);
nand U14873 (N_14873,N_14770,N_14705);
and U14874 (N_14874,N_14663,N_14781);
or U14875 (N_14875,N_14719,N_14776);
nand U14876 (N_14876,N_14655,N_14687);
nor U14877 (N_14877,N_14610,N_14619);
nor U14878 (N_14878,N_14712,N_14666);
nand U14879 (N_14879,N_14667,N_14720);
xnor U14880 (N_14880,N_14659,N_14709);
and U14881 (N_14881,N_14699,N_14649);
and U14882 (N_14882,N_14796,N_14785);
or U14883 (N_14883,N_14661,N_14739);
nor U14884 (N_14884,N_14632,N_14639);
nand U14885 (N_14885,N_14729,N_14742);
and U14886 (N_14886,N_14697,N_14793);
or U14887 (N_14887,N_14600,N_14690);
xnor U14888 (N_14888,N_14678,N_14674);
nor U14889 (N_14889,N_14673,N_14745);
or U14890 (N_14890,N_14688,N_14750);
nand U14891 (N_14891,N_14704,N_14726);
xnor U14892 (N_14892,N_14710,N_14768);
and U14893 (N_14893,N_14614,N_14724);
xnor U14894 (N_14894,N_14652,N_14641);
nor U14895 (N_14895,N_14749,N_14621);
or U14896 (N_14896,N_14792,N_14672);
and U14897 (N_14897,N_14791,N_14772);
or U14898 (N_14898,N_14691,N_14601);
or U14899 (N_14899,N_14789,N_14787);
nor U14900 (N_14900,N_14781,N_14686);
nand U14901 (N_14901,N_14600,N_14676);
nor U14902 (N_14902,N_14626,N_14764);
nand U14903 (N_14903,N_14720,N_14628);
or U14904 (N_14904,N_14635,N_14667);
and U14905 (N_14905,N_14651,N_14695);
xor U14906 (N_14906,N_14690,N_14685);
nand U14907 (N_14907,N_14652,N_14729);
nor U14908 (N_14908,N_14763,N_14628);
xor U14909 (N_14909,N_14797,N_14685);
nor U14910 (N_14910,N_14679,N_14610);
xnor U14911 (N_14911,N_14612,N_14690);
xnor U14912 (N_14912,N_14659,N_14681);
nand U14913 (N_14913,N_14612,N_14738);
xor U14914 (N_14914,N_14740,N_14671);
nor U14915 (N_14915,N_14638,N_14644);
and U14916 (N_14916,N_14611,N_14637);
and U14917 (N_14917,N_14734,N_14746);
and U14918 (N_14918,N_14709,N_14762);
nor U14919 (N_14919,N_14775,N_14723);
and U14920 (N_14920,N_14615,N_14752);
and U14921 (N_14921,N_14639,N_14758);
and U14922 (N_14922,N_14645,N_14642);
xor U14923 (N_14923,N_14633,N_14701);
nand U14924 (N_14924,N_14729,N_14678);
nand U14925 (N_14925,N_14631,N_14765);
nand U14926 (N_14926,N_14650,N_14654);
and U14927 (N_14927,N_14780,N_14753);
nor U14928 (N_14928,N_14740,N_14621);
xnor U14929 (N_14929,N_14639,N_14605);
or U14930 (N_14930,N_14661,N_14691);
nand U14931 (N_14931,N_14676,N_14634);
xnor U14932 (N_14932,N_14755,N_14657);
nand U14933 (N_14933,N_14694,N_14683);
or U14934 (N_14934,N_14698,N_14606);
xor U14935 (N_14935,N_14602,N_14603);
and U14936 (N_14936,N_14758,N_14697);
and U14937 (N_14937,N_14618,N_14661);
nor U14938 (N_14938,N_14607,N_14626);
nand U14939 (N_14939,N_14720,N_14691);
nand U14940 (N_14940,N_14633,N_14756);
nand U14941 (N_14941,N_14745,N_14710);
or U14942 (N_14942,N_14787,N_14743);
xor U14943 (N_14943,N_14686,N_14771);
nor U14944 (N_14944,N_14626,N_14782);
nand U14945 (N_14945,N_14724,N_14649);
xor U14946 (N_14946,N_14786,N_14785);
nand U14947 (N_14947,N_14679,N_14787);
nor U14948 (N_14948,N_14752,N_14618);
or U14949 (N_14949,N_14671,N_14667);
or U14950 (N_14950,N_14789,N_14766);
or U14951 (N_14951,N_14781,N_14659);
xor U14952 (N_14952,N_14635,N_14702);
xnor U14953 (N_14953,N_14607,N_14774);
nand U14954 (N_14954,N_14628,N_14666);
nor U14955 (N_14955,N_14769,N_14619);
nor U14956 (N_14956,N_14671,N_14622);
nor U14957 (N_14957,N_14776,N_14705);
nor U14958 (N_14958,N_14643,N_14629);
xor U14959 (N_14959,N_14696,N_14663);
and U14960 (N_14960,N_14749,N_14631);
nand U14961 (N_14961,N_14645,N_14702);
or U14962 (N_14962,N_14785,N_14667);
or U14963 (N_14963,N_14785,N_14648);
nor U14964 (N_14964,N_14659,N_14686);
nor U14965 (N_14965,N_14617,N_14751);
or U14966 (N_14966,N_14743,N_14621);
xnor U14967 (N_14967,N_14689,N_14729);
nor U14968 (N_14968,N_14795,N_14626);
or U14969 (N_14969,N_14621,N_14616);
nand U14970 (N_14970,N_14745,N_14616);
or U14971 (N_14971,N_14652,N_14650);
and U14972 (N_14972,N_14753,N_14664);
or U14973 (N_14973,N_14630,N_14600);
and U14974 (N_14974,N_14763,N_14799);
nor U14975 (N_14975,N_14733,N_14610);
and U14976 (N_14976,N_14636,N_14792);
xor U14977 (N_14977,N_14704,N_14791);
nand U14978 (N_14978,N_14663,N_14798);
xnor U14979 (N_14979,N_14647,N_14782);
or U14980 (N_14980,N_14741,N_14622);
nand U14981 (N_14981,N_14741,N_14701);
and U14982 (N_14982,N_14740,N_14642);
nand U14983 (N_14983,N_14648,N_14622);
or U14984 (N_14984,N_14788,N_14646);
or U14985 (N_14985,N_14713,N_14740);
nand U14986 (N_14986,N_14762,N_14649);
nand U14987 (N_14987,N_14725,N_14784);
nor U14988 (N_14988,N_14741,N_14760);
xnor U14989 (N_14989,N_14613,N_14718);
or U14990 (N_14990,N_14792,N_14623);
xor U14991 (N_14991,N_14690,N_14659);
or U14992 (N_14992,N_14751,N_14672);
xor U14993 (N_14993,N_14632,N_14660);
xnor U14994 (N_14994,N_14682,N_14715);
xnor U14995 (N_14995,N_14604,N_14797);
nor U14996 (N_14996,N_14715,N_14635);
nor U14997 (N_14997,N_14678,N_14701);
nor U14998 (N_14998,N_14796,N_14745);
or U14999 (N_14999,N_14769,N_14622);
or U15000 (N_15000,N_14922,N_14932);
xor U15001 (N_15001,N_14831,N_14857);
or U15002 (N_15002,N_14971,N_14875);
xor U15003 (N_15003,N_14935,N_14841);
xor U15004 (N_15004,N_14833,N_14802);
nand U15005 (N_15005,N_14890,N_14997);
nand U15006 (N_15006,N_14822,N_14901);
or U15007 (N_15007,N_14903,N_14891);
or U15008 (N_15008,N_14917,N_14869);
and U15009 (N_15009,N_14993,N_14871);
or U15010 (N_15010,N_14807,N_14898);
xor U15011 (N_15011,N_14976,N_14945);
or U15012 (N_15012,N_14947,N_14916);
nand U15013 (N_15013,N_14979,N_14940);
nand U15014 (N_15014,N_14938,N_14994);
nor U15015 (N_15015,N_14999,N_14828);
nor U15016 (N_15016,N_14918,N_14937);
nor U15017 (N_15017,N_14970,N_14952);
xor U15018 (N_15018,N_14811,N_14817);
nor U15019 (N_15019,N_14855,N_14928);
xnor U15020 (N_15020,N_14963,N_14850);
and U15021 (N_15021,N_14859,N_14899);
nand U15022 (N_15022,N_14900,N_14824);
xor U15023 (N_15023,N_14830,N_14878);
or U15024 (N_15024,N_14911,N_14853);
nand U15025 (N_15025,N_14998,N_14962);
or U15026 (N_15026,N_14961,N_14924);
nand U15027 (N_15027,N_14879,N_14927);
nor U15028 (N_15028,N_14959,N_14907);
nand U15029 (N_15029,N_14837,N_14810);
nor U15030 (N_15030,N_14861,N_14931);
xor U15031 (N_15031,N_14866,N_14801);
xor U15032 (N_15032,N_14834,N_14863);
xor U15033 (N_15033,N_14967,N_14854);
or U15034 (N_15034,N_14956,N_14930);
xnor U15035 (N_15035,N_14981,N_14934);
nor U15036 (N_15036,N_14887,N_14876);
or U15037 (N_15037,N_14835,N_14896);
nand U15038 (N_15038,N_14953,N_14872);
or U15039 (N_15039,N_14864,N_14987);
and U15040 (N_15040,N_14960,N_14814);
xnor U15041 (N_15041,N_14803,N_14836);
nor U15042 (N_15042,N_14825,N_14882);
and U15043 (N_15043,N_14974,N_14865);
or U15044 (N_15044,N_14925,N_14820);
nor U15045 (N_15045,N_14926,N_14868);
xnor U15046 (N_15046,N_14816,N_14949);
and U15047 (N_15047,N_14951,N_14812);
nor U15048 (N_15048,N_14988,N_14908);
or U15049 (N_15049,N_14968,N_14972);
and U15050 (N_15050,N_14912,N_14893);
nand U15051 (N_15051,N_14941,N_14991);
nor U15052 (N_15052,N_14975,N_14989);
nor U15053 (N_15053,N_14950,N_14889);
and U15054 (N_15054,N_14886,N_14877);
nand U15055 (N_15055,N_14832,N_14884);
or U15056 (N_15056,N_14821,N_14982);
xor U15057 (N_15057,N_14856,N_14885);
xor U15058 (N_15058,N_14929,N_14992);
nand U15059 (N_15059,N_14995,N_14800);
nand U15060 (N_15060,N_14910,N_14915);
xor U15061 (N_15061,N_14874,N_14897);
xor U15062 (N_15062,N_14996,N_14920);
and U15063 (N_15063,N_14838,N_14806);
nand U15064 (N_15064,N_14943,N_14823);
nand U15065 (N_15065,N_14954,N_14902);
and U15066 (N_15066,N_14843,N_14880);
nor U15067 (N_15067,N_14870,N_14809);
or U15068 (N_15068,N_14826,N_14990);
xor U15069 (N_15069,N_14936,N_14986);
xnor U15070 (N_15070,N_14923,N_14819);
or U15071 (N_15071,N_14909,N_14921);
xnor U15072 (N_15072,N_14829,N_14948);
or U15073 (N_15073,N_14860,N_14913);
or U15074 (N_15074,N_14978,N_14946);
nor U15075 (N_15075,N_14905,N_14815);
xnor U15076 (N_15076,N_14858,N_14846);
nor U15077 (N_15077,N_14906,N_14904);
xnor U15078 (N_15078,N_14983,N_14914);
nor U15079 (N_15079,N_14977,N_14958);
and U15080 (N_15080,N_14844,N_14985);
or U15081 (N_15081,N_14805,N_14973);
nand U15082 (N_15082,N_14849,N_14851);
and U15083 (N_15083,N_14881,N_14980);
nor U15084 (N_15084,N_14965,N_14873);
xnor U15085 (N_15085,N_14840,N_14966);
nand U15086 (N_15086,N_14842,N_14888);
nand U15087 (N_15087,N_14894,N_14845);
xor U15088 (N_15088,N_14862,N_14883);
nor U15089 (N_15089,N_14942,N_14919);
nand U15090 (N_15090,N_14933,N_14939);
nand U15091 (N_15091,N_14957,N_14827);
nor U15092 (N_15092,N_14895,N_14867);
or U15093 (N_15093,N_14818,N_14848);
and U15094 (N_15094,N_14847,N_14852);
nor U15095 (N_15095,N_14839,N_14944);
and U15096 (N_15096,N_14964,N_14804);
and U15097 (N_15097,N_14955,N_14892);
and U15098 (N_15098,N_14969,N_14984);
xor U15099 (N_15099,N_14808,N_14813);
xor U15100 (N_15100,N_14842,N_14970);
and U15101 (N_15101,N_14941,N_14852);
xnor U15102 (N_15102,N_14971,N_14815);
nand U15103 (N_15103,N_14885,N_14839);
nor U15104 (N_15104,N_14956,N_14892);
nand U15105 (N_15105,N_14851,N_14983);
nor U15106 (N_15106,N_14817,N_14808);
xor U15107 (N_15107,N_14884,N_14806);
or U15108 (N_15108,N_14987,N_14865);
or U15109 (N_15109,N_14890,N_14977);
or U15110 (N_15110,N_14930,N_14878);
nand U15111 (N_15111,N_14993,N_14870);
and U15112 (N_15112,N_14839,N_14992);
and U15113 (N_15113,N_14838,N_14888);
xnor U15114 (N_15114,N_14903,N_14987);
or U15115 (N_15115,N_14919,N_14988);
nand U15116 (N_15116,N_14837,N_14835);
xnor U15117 (N_15117,N_14885,N_14805);
or U15118 (N_15118,N_14910,N_14877);
nand U15119 (N_15119,N_14835,N_14819);
nor U15120 (N_15120,N_14826,N_14950);
xnor U15121 (N_15121,N_14963,N_14896);
nand U15122 (N_15122,N_14990,N_14838);
and U15123 (N_15123,N_14859,N_14953);
nor U15124 (N_15124,N_14928,N_14917);
xor U15125 (N_15125,N_14860,N_14879);
nand U15126 (N_15126,N_14931,N_14877);
and U15127 (N_15127,N_14860,N_14854);
xor U15128 (N_15128,N_14835,N_14865);
nand U15129 (N_15129,N_14986,N_14998);
nand U15130 (N_15130,N_14998,N_14910);
or U15131 (N_15131,N_14947,N_14826);
or U15132 (N_15132,N_14811,N_14962);
nand U15133 (N_15133,N_14929,N_14832);
nor U15134 (N_15134,N_14955,N_14922);
nand U15135 (N_15135,N_14915,N_14936);
xnor U15136 (N_15136,N_14812,N_14832);
xor U15137 (N_15137,N_14845,N_14988);
nand U15138 (N_15138,N_14844,N_14824);
or U15139 (N_15139,N_14825,N_14819);
nor U15140 (N_15140,N_14904,N_14813);
nor U15141 (N_15141,N_14837,N_14825);
nand U15142 (N_15142,N_14984,N_14854);
nor U15143 (N_15143,N_14834,N_14912);
xor U15144 (N_15144,N_14967,N_14815);
or U15145 (N_15145,N_14811,N_14984);
or U15146 (N_15146,N_14845,N_14985);
or U15147 (N_15147,N_14810,N_14869);
xnor U15148 (N_15148,N_14879,N_14952);
or U15149 (N_15149,N_14909,N_14827);
or U15150 (N_15150,N_14984,N_14951);
and U15151 (N_15151,N_14831,N_14956);
xnor U15152 (N_15152,N_14922,N_14975);
nor U15153 (N_15153,N_14862,N_14985);
nor U15154 (N_15154,N_14805,N_14963);
nand U15155 (N_15155,N_14972,N_14984);
nor U15156 (N_15156,N_14910,N_14996);
xnor U15157 (N_15157,N_14882,N_14904);
xnor U15158 (N_15158,N_14922,N_14808);
or U15159 (N_15159,N_14819,N_14862);
and U15160 (N_15160,N_14905,N_14993);
xor U15161 (N_15161,N_14927,N_14814);
and U15162 (N_15162,N_14952,N_14801);
nand U15163 (N_15163,N_14957,N_14848);
nor U15164 (N_15164,N_14919,N_14853);
xor U15165 (N_15165,N_14948,N_14818);
and U15166 (N_15166,N_14826,N_14939);
nor U15167 (N_15167,N_14968,N_14893);
and U15168 (N_15168,N_14890,N_14827);
and U15169 (N_15169,N_14833,N_14819);
nand U15170 (N_15170,N_14950,N_14809);
nand U15171 (N_15171,N_14902,N_14843);
nor U15172 (N_15172,N_14874,N_14807);
and U15173 (N_15173,N_14970,N_14806);
nand U15174 (N_15174,N_14829,N_14864);
and U15175 (N_15175,N_14992,N_14882);
nor U15176 (N_15176,N_14809,N_14900);
or U15177 (N_15177,N_14864,N_14922);
and U15178 (N_15178,N_14904,N_14949);
nand U15179 (N_15179,N_14823,N_14979);
and U15180 (N_15180,N_14981,N_14956);
xnor U15181 (N_15181,N_14831,N_14862);
or U15182 (N_15182,N_14934,N_14938);
xnor U15183 (N_15183,N_14902,N_14846);
xnor U15184 (N_15184,N_14804,N_14937);
and U15185 (N_15185,N_14845,N_14842);
nand U15186 (N_15186,N_14906,N_14892);
and U15187 (N_15187,N_14937,N_14997);
xor U15188 (N_15188,N_14845,N_14965);
nor U15189 (N_15189,N_14898,N_14921);
nor U15190 (N_15190,N_14827,N_14819);
nor U15191 (N_15191,N_14948,N_14895);
nand U15192 (N_15192,N_14939,N_14889);
xor U15193 (N_15193,N_14963,N_14819);
xnor U15194 (N_15194,N_14816,N_14881);
or U15195 (N_15195,N_14820,N_14845);
nand U15196 (N_15196,N_14816,N_14958);
nand U15197 (N_15197,N_14821,N_14962);
or U15198 (N_15198,N_14911,N_14932);
xor U15199 (N_15199,N_14861,N_14864);
nor U15200 (N_15200,N_15094,N_15183);
and U15201 (N_15201,N_15181,N_15162);
and U15202 (N_15202,N_15103,N_15069);
nor U15203 (N_15203,N_15009,N_15010);
and U15204 (N_15204,N_15168,N_15182);
and U15205 (N_15205,N_15144,N_15122);
nand U15206 (N_15206,N_15025,N_15081);
nor U15207 (N_15207,N_15151,N_15071);
and U15208 (N_15208,N_15119,N_15033);
nor U15209 (N_15209,N_15142,N_15096);
nor U15210 (N_15210,N_15012,N_15185);
or U15211 (N_15211,N_15145,N_15193);
xor U15212 (N_15212,N_15074,N_15179);
nand U15213 (N_15213,N_15005,N_15194);
xor U15214 (N_15214,N_15014,N_15178);
nand U15215 (N_15215,N_15070,N_15196);
and U15216 (N_15216,N_15028,N_15149);
nand U15217 (N_15217,N_15127,N_15006);
and U15218 (N_15218,N_15140,N_15124);
or U15219 (N_15219,N_15163,N_15176);
xor U15220 (N_15220,N_15047,N_15030);
nand U15221 (N_15221,N_15132,N_15035);
nor U15222 (N_15222,N_15195,N_15027);
xnor U15223 (N_15223,N_15092,N_15054);
or U15224 (N_15224,N_15143,N_15101);
or U15225 (N_15225,N_15051,N_15078);
nor U15226 (N_15226,N_15065,N_15186);
nor U15227 (N_15227,N_15073,N_15154);
or U15228 (N_15228,N_15104,N_15164);
nor U15229 (N_15229,N_15088,N_15022);
nor U15230 (N_15230,N_15155,N_15023);
xor U15231 (N_15231,N_15056,N_15068);
and U15232 (N_15232,N_15062,N_15117);
or U15233 (N_15233,N_15123,N_15105);
nor U15234 (N_15234,N_15174,N_15067);
xor U15235 (N_15235,N_15017,N_15130);
and U15236 (N_15236,N_15095,N_15083);
nand U15237 (N_15237,N_15152,N_15192);
nand U15238 (N_15238,N_15125,N_15175);
or U15239 (N_15239,N_15161,N_15001);
nor U15240 (N_15240,N_15066,N_15166);
or U15241 (N_15241,N_15169,N_15141);
xnor U15242 (N_15242,N_15019,N_15053);
xnor U15243 (N_15243,N_15075,N_15102);
nand U15244 (N_15244,N_15058,N_15044);
and U15245 (N_15245,N_15063,N_15126);
xnor U15246 (N_15246,N_15165,N_15170);
nor U15247 (N_15247,N_15000,N_15159);
nand U15248 (N_15248,N_15138,N_15004);
and U15249 (N_15249,N_15049,N_15172);
nor U15250 (N_15250,N_15133,N_15109);
or U15251 (N_15251,N_15055,N_15043);
nand U15252 (N_15252,N_15158,N_15052);
or U15253 (N_15253,N_15120,N_15032);
and U15254 (N_15254,N_15199,N_15050);
xnor U15255 (N_15255,N_15198,N_15137);
nand U15256 (N_15256,N_15110,N_15118);
and U15257 (N_15257,N_15057,N_15189);
xnor U15258 (N_15258,N_15173,N_15188);
and U15259 (N_15259,N_15091,N_15040);
xor U15260 (N_15260,N_15038,N_15018);
or U15261 (N_15261,N_15146,N_15016);
nor U15262 (N_15262,N_15114,N_15041);
or U15263 (N_15263,N_15100,N_15059);
or U15264 (N_15264,N_15082,N_15167);
xor U15265 (N_15265,N_15148,N_15191);
and U15266 (N_15266,N_15157,N_15139);
nand U15267 (N_15267,N_15099,N_15197);
xnor U15268 (N_15268,N_15112,N_15007);
nor U15269 (N_15269,N_15131,N_15128);
xor U15270 (N_15270,N_15037,N_15042);
nand U15271 (N_15271,N_15106,N_15015);
nor U15272 (N_15272,N_15108,N_15011);
or U15273 (N_15273,N_15085,N_15003);
nand U15274 (N_15274,N_15084,N_15029);
xnor U15275 (N_15275,N_15045,N_15190);
or U15276 (N_15276,N_15048,N_15086);
xor U15277 (N_15277,N_15013,N_15026);
xor U15278 (N_15278,N_15171,N_15116);
nand U15279 (N_15279,N_15002,N_15077);
or U15280 (N_15280,N_15111,N_15153);
or U15281 (N_15281,N_15135,N_15031);
and U15282 (N_15282,N_15156,N_15064);
and U15283 (N_15283,N_15129,N_15136);
nand U15284 (N_15284,N_15097,N_15113);
nor U15285 (N_15285,N_15107,N_15021);
nor U15286 (N_15286,N_15061,N_15177);
nand U15287 (N_15287,N_15090,N_15036);
nor U15288 (N_15288,N_15134,N_15187);
xor U15289 (N_15289,N_15046,N_15008);
and U15290 (N_15290,N_15087,N_15115);
or U15291 (N_15291,N_15160,N_15039);
or U15292 (N_15292,N_15079,N_15150);
nor U15293 (N_15293,N_15020,N_15034);
nor U15294 (N_15294,N_15184,N_15024);
xnor U15295 (N_15295,N_15080,N_15121);
and U15296 (N_15296,N_15098,N_15180);
or U15297 (N_15297,N_15076,N_15060);
nor U15298 (N_15298,N_15093,N_15147);
xor U15299 (N_15299,N_15072,N_15089);
and U15300 (N_15300,N_15119,N_15163);
and U15301 (N_15301,N_15175,N_15153);
nor U15302 (N_15302,N_15190,N_15195);
nor U15303 (N_15303,N_15065,N_15090);
or U15304 (N_15304,N_15051,N_15184);
nand U15305 (N_15305,N_15027,N_15066);
nand U15306 (N_15306,N_15196,N_15062);
xor U15307 (N_15307,N_15106,N_15001);
or U15308 (N_15308,N_15166,N_15041);
xnor U15309 (N_15309,N_15165,N_15009);
xor U15310 (N_15310,N_15127,N_15082);
nand U15311 (N_15311,N_15131,N_15129);
nor U15312 (N_15312,N_15100,N_15147);
or U15313 (N_15313,N_15055,N_15086);
xor U15314 (N_15314,N_15183,N_15095);
xor U15315 (N_15315,N_15097,N_15014);
and U15316 (N_15316,N_15142,N_15137);
xnor U15317 (N_15317,N_15125,N_15149);
nor U15318 (N_15318,N_15129,N_15033);
nor U15319 (N_15319,N_15021,N_15000);
nor U15320 (N_15320,N_15013,N_15164);
or U15321 (N_15321,N_15060,N_15070);
nor U15322 (N_15322,N_15199,N_15012);
nor U15323 (N_15323,N_15067,N_15133);
nor U15324 (N_15324,N_15190,N_15184);
or U15325 (N_15325,N_15144,N_15009);
nand U15326 (N_15326,N_15197,N_15181);
xnor U15327 (N_15327,N_15147,N_15141);
xnor U15328 (N_15328,N_15041,N_15085);
or U15329 (N_15329,N_15167,N_15035);
or U15330 (N_15330,N_15023,N_15136);
and U15331 (N_15331,N_15181,N_15155);
xnor U15332 (N_15332,N_15187,N_15111);
nor U15333 (N_15333,N_15054,N_15123);
nand U15334 (N_15334,N_15169,N_15117);
xor U15335 (N_15335,N_15029,N_15156);
nor U15336 (N_15336,N_15197,N_15085);
or U15337 (N_15337,N_15072,N_15023);
and U15338 (N_15338,N_15003,N_15141);
xnor U15339 (N_15339,N_15032,N_15042);
and U15340 (N_15340,N_15109,N_15165);
nor U15341 (N_15341,N_15011,N_15187);
and U15342 (N_15342,N_15134,N_15145);
nand U15343 (N_15343,N_15010,N_15159);
or U15344 (N_15344,N_15090,N_15169);
xor U15345 (N_15345,N_15045,N_15074);
nor U15346 (N_15346,N_15044,N_15132);
and U15347 (N_15347,N_15166,N_15094);
nand U15348 (N_15348,N_15040,N_15148);
xnor U15349 (N_15349,N_15013,N_15143);
and U15350 (N_15350,N_15002,N_15159);
xor U15351 (N_15351,N_15063,N_15102);
nand U15352 (N_15352,N_15037,N_15047);
nor U15353 (N_15353,N_15004,N_15148);
nor U15354 (N_15354,N_15161,N_15044);
and U15355 (N_15355,N_15017,N_15148);
and U15356 (N_15356,N_15039,N_15086);
xor U15357 (N_15357,N_15052,N_15184);
nor U15358 (N_15358,N_15187,N_15097);
and U15359 (N_15359,N_15087,N_15052);
nand U15360 (N_15360,N_15166,N_15180);
xnor U15361 (N_15361,N_15084,N_15023);
nand U15362 (N_15362,N_15133,N_15060);
nand U15363 (N_15363,N_15016,N_15145);
nor U15364 (N_15364,N_15068,N_15169);
nor U15365 (N_15365,N_15104,N_15022);
and U15366 (N_15366,N_15099,N_15150);
xor U15367 (N_15367,N_15045,N_15062);
nand U15368 (N_15368,N_15180,N_15111);
xnor U15369 (N_15369,N_15089,N_15133);
and U15370 (N_15370,N_15005,N_15035);
and U15371 (N_15371,N_15166,N_15186);
xnor U15372 (N_15372,N_15075,N_15120);
and U15373 (N_15373,N_15099,N_15028);
or U15374 (N_15374,N_15006,N_15011);
nor U15375 (N_15375,N_15028,N_15194);
nor U15376 (N_15376,N_15072,N_15010);
nand U15377 (N_15377,N_15083,N_15013);
xnor U15378 (N_15378,N_15160,N_15000);
or U15379 (N_15379,N_15112,N_15012);
and U15380 (N_15380,N_15106,N_15115);
xnor U15381 (N_15381,N_15092,N_15030);
or U15382 (N_15382,N_15076,N_15184);
nor U15383 (N_15383,N_15170,N_15155);
nand U15384 (N_15384,N_15028,N_15011);
and U15385 (N_15385,N_15020,N_15115);
xor U15386 (N_15386,N_15185,N_15036);
nor U15387 (N_15387,N_15076,N_15059);
or U15388 (N_15388,N_15108,N_15167);
xnor U15389 (N_15389,N_15028,N_15190);
nand U15390 (N_15390,N_15055,N_15106);
nor U15391 (N_15391,N_15023,N_15087);
xor U15392 (N_15392,N_15090,N_15138);
nor U15393 (N_15393,N_15138,N_15118);
and U15394 (N_15394,N_15028,N_15066);
nor U15395 (N_15395,N_15019,N_15106);
or U15396 (N_15396,N_15188,N_15171);
or U15397 (N_15397,N_15008,N_15182);
nand U15398 (N_15398,N_15178,N_15033);
nand U15399 (N_15399,N_15062,N_15029);
and U15400 (N_15400,N_15389,N_15255);
nor U15401 (N_15401,N_15357,N_15206);
or U15402 (N_15402,N_15396,N_15254);
or U15403 (N_15403,N_15225,N_15200);
or U15404 (N_15404,N_15323,N_15238);
or U15405 (N_15405,N_15213,N_15372);
nand U15406 (N_15406,N_15349,N_15312);
or U15407 (N_15407,N_15356,N_15368);
nand U15408 (N_15408,N_15335,N_15233);
or U15409 (N_15409,N_15241,N_15310);
or U15410 (N_15410,N_15234,N_15379);
nor U15411 (N_15411,N_15245,N_15275);
or U15412 (N_15412,N_15363,N_15237);
xnor U15413 (N_15413,N_15302,N_15226);
and U15414 (N_15414,N_15290,N_15307);
nor U15415 (N_15415,N_15215,N_15284);
and U15416 (N_15416,N_15220,N_15322);
and U15417 (N_15417,N_15325,N_15311);
nor U15418 (N_15418,N_15384,N_15293);
and U15419 (N_15419,N_15367,N_15385);
nor U15420 (N_15420,N_15364,N_15398);
and U15421 (N_15421,N_15388,N_15395);
nor U15422 (N_15422,N_15279,N_15222);
nand U15423 (N_15423,N_15393,N_15341);
nor U15424 (N_15424,N_15337,N_15281);
and U15425 (N_15425,N_15265,N_15329);
xor U15426 (N_15426,N_15327,N_15294);
nor U15427 (N_15427,N_15274,N_15288);
xnor U15428 (N_15428,N_15257,N_15314);
nor U15429 (N_15429,N_15336,N_15259);
or U15430 (N_15430,N_15375,N_15391);
nand U15431 (N_15431,N_15269,N_15240);
and U15432 (N_15432,N_15242,N_15278);
xor U15433 (N_15433,N_15203,N_15317);
xnor U15434 (N_15434,N_15369,N_15295);
nor U15435 (N_15435,N_15258,N_15286);
nor U15436 (N_15436,N_15320,N_15304);
and U15437 (N_15437,N_15291,N_15287);
or U15438 (N_15438,N_15266,N_15331);
nor U15439 (N_15439,N_15247,N_15271);
xnor U15440 (N_15440,N_15344,N_15352);
and U15441 (N_15441,N_15360,N_15359);
nor U15442 (N_15442,N_15345,N_15253);
nand U15443 (N_15443,N_15216,N_15223);
nor U15444 (N_15444,N_15209,N_15371);
xnor U15445 (N_15445,N_15251,N_15228);
and U15446 (N_15446,N_15208,N_15272);
xor U15447 (N_15447,N_15313,N_15205);
and U15448 (N_15448,N_15218,N_15250);
and U15449 (N_15449,N_15358,N_15297);
nor U15450 (N_15450,N_15256,N_15268);
nand U15451 (N_15451,N_15381,N_15236);
xor U15452 (N_15452,N_15300,N_15227);
nand U15453 (N_15453,N_15267,N_15366);
nand U15454 (N_15454,N_15382,N_15270);
xor U15455 (N_15455,N_15387,N_15229);
or U15456 (N_15456,N_15365,N_15361);
and U15457 (N_15457,N_15210,N_15373);
or U15458 (N_15458,N_15390,N_15342);
or U15459 (N_15459,N_15231,N_15301);
or U15460 (N_15460,N_15232,N_15249);
xnor U15461 (N_15461,N_15333,N_15285);
nor U15462 (N_15462,N_15201,N_15332);
nor U15463 (N_15463,N_15276,N_15211);
nor U15464 (N_15464,N_15383,N_15315);
nand U15465 (N_15465,N_15350,N_15326);
or U15466 (N_15466,N_15212,N_15370);
nor U15467 (N_15467,N_15303,N_15243);
nor U15468 (N_15468,N_15392,N_15282);
and U15469 (N_15469,N_15321,N_15219);
and U15470 (N_15470,N_15207,N_15280);
nand U15471 (N_15471,N_15224,N_15298);
xor U15472 (N_15472,N_15380,N_15362);
or U15473 (N_15473,N_15318,N_15289);
nand U15474 (N_15474,N_15324,N_15204);
xor U15475 (N_15475,N_15394,N_15202);
nor U15476 (N_15476,N_15214,N_15377);
nor U15477 (N_15477,N_15339,N_15221);
and U15478 (N_15478,N_15346,N_15263);
or U15479 (N_15479,N_15283,N_15338);
nand U15480 (N_15480,N_15299,N_15305);
nand U15481 (N_15481,N_15319,N_15347);
and U15482 (N_15482,N_15397,N_15248);
xnor U15483 (N_15483,N_15316,N_15308);
or U15484 (N_15484,N_15348,N_15306);
and U15485 (N_15485,N_15262,N_15386);
or U15486 (N_15486,N_15292,N_15296);
nand U15487 (N_15487,N_15328,N_15376);
and U15488 (N_15488,N_15353,N_15252);
nor U15489 (N_15489,N_15340,N_15351);
or U15490 (N_15490,N_15264,N_15343);
nand U15491 (N_15491,N_15355,N_15239);
nor U15492 (N_15492,N_15378,N_15330);
nand U15493 (N_15493,N_15235,N_15309);
xnor U15494 (N_15494,N_15354,N_15217);
or U15495 (N_15495,N_15334,N_15261);
nor U15496 (N_15496,N_15277,N_15399);
nor U15497 (N_15497,N_15374,N_15230);
nand U15498 (N_15498,N_15246,N_15260);
and U15499 (N_15499,N_15244,N_15273);
nor U15500 (N_15500,N_15300,N_15374);
nand U15501 (N_15501,N_15260,N_15203);
or U15502 (N_15502,N_15254,N_15321);
xnor U15503 (N_15503,N_15388,N_15356);
nor U15504 (N_15504,N_15328,N_15268);
nand U15505 (N_15505,N_15273,N_15238);
nand U15506 (N_15506,N_15373,N_15383);
xnor U15507 (N_15507,N_15369,N_15299);
nand U15508 (N_15508,N_15235,N_15359);
nor U15509 (N_15509,N_15335,N_15220);
nor U15510 (N_15510,N_15394,N_15201);
and U15511 (N_15511,N_15237,N_15231);
nor U15512 (N_15512,N_15316,N_15223);
nand U15513 (N_15513,N_15259,N_15355);
or U15514 (N_15514,N_15229,N_15396);
nand U15515 (N_15515,N_15268,N_15288);
nor U15516 (N_15516,N_15360,N_15324);
nor U15517 (N_15517,N_15294,N_15388);
and U15518 (N_15518,N_15305,N_15312);
xor U15519 (N_15519,N_15368,N_15267);
xnor U15520 (N_15520,N_15330,N_15308);
nor U15521 (N_15521,N_15383,N_15338);
nor U15522 (N_15522,N_15311,N_15396);
nand U15523 (N_15523,N_15319,N_15270);
nand U15524 (N_15524,N_15286,N_15389);
nor U15525 (N_15525,N_15390,N_15228);
and U15526 (N_15526,N_15204,N_15344);
or U15527 (N_15527,N_15291,N_15365);
nand U15528 (N_15528,N_15381,N_15210);
and U15529 (N_15529,N_15257,N_15287);
or U15530 (N_15530,N_15264,N_15272);
nor U15531 (N_15531,N_15258,N_15372);
nor U15532 (N_15532,N_15217,N_15339);
nor U15533 (N_15533,N_15375,N_15241);
nor U15534 (N_15534,N_15251,N_15361);
nor U15535 (N_15535,N_15251,N_15350);
nand U15536 (N_15536,N_15270,N_15373);
nand U15537 (N_15537,N_15256,N_15214);
nor U15538 (N_15538,N_15289,N_15216);
and U15539 (N_15539,N_15220,N_15310);
xor U15540 (N_15540,N_15324,N_15240);
and U15541 (N_15541,N_15224,N_15275);
nor U15542 (N_15542,N_15318,N_15322);
nor U15543 (N_15543,N_15319,N_15294);
or U15544 (N_15544,N_15293,N_15378);
and U15545 (N_15545,N_15231,N_15274);
nor U15546 (N_15546,N_15299,N_15228);
nor U15547 (N_15547,N_15365,N_15316);
xor U15548 (N_15548,N_15346,N_15272);
xor U15549 (N_15549,N_15278,N_15201);
nor U15550 (N_15550,N_15358,N_15274);
xor U15551 (N_15551,N_15263,N_15227);
nand U15552 (N_15552,N_15233,N_15375);
nand U15553 (N_15553,N_15303,N_15398);
or U15554 (N_15554,N_15264,N_15399);
or U15555 (N_15555,N_15381,N_15267);
and U15556 (N_15556,N_15321,N_15236);
nand U15557 (N_15557,N_15237,N_15319);
or U15558 (N_15558,N_15238,N_15267);
or U15559 (N_15559,N_15287,N_15295);
nor U15560 (N_15560,N_15287,N_15385);
nor U15561 (N_15561,N_15289,N_15256);
nand U15562 (N_15562,N_15369,N_15363);
or U15563 (N_15563,N_15268,N_15289);
nor U15564 (N_15564,N_15372,N_15255);
or U15565 (N_15565,N_15325,N_15306);
and U15566 (N_15566,N_15204,N_15254);
nand U15567 (N_15567,N_15349,N_15278);
and U15568 (N_15568,N_15289,N_15355);
nand U15569 (N_15569,N_15223,N_15279);
nand U15570 (N_15570,N_15243,N_15211);
xnor U15571 (N_15571,N_15252,N_15203);
and U15572 (N_15572,N_15380,N_15306);
xor U15573 (N_15573,N_15258,N_15358);
nand U15574 (N_15574,N_15267,N_15338);
and U15575 (N_15575,N_15339,N_15381);
nor U15576 (N_15576,N_15255,N_15300);
and U15577 (N_15577,N_15280,N_15344);
xor U15578 (N_15578,N_15391,N_15341);
nor U15579 (N_15579,N_15365,N_15210);
nor U15580 (N_15580,N_15200,N_15295);
xor U15581 (N_15581,N_15211,N_15240);
or U15582 (N_15582,N_15270,N_15210);
nor U15583 (N_15583,N_15344,N_15250);
and U15584 (N_15584,N_15398,N_15363);
or U15585 (N_15585,N_15220,N_15265);
or U15586 (N_15586,N_15386,N_15305);
xor U15587 (N_15587,N_15269,N_15311);
and U15588 (N_15588,N_15367,N_15215);
or U15589 (N_15589,N_15356,N_15264);
nand U15590 (N_15590,N_15229,N_15250);
nand U15591 (N_15591,N_15223,N_15309);
nand U15592 (N_15592,N_15360,N_15346);
xor U15593 (N_15593,N_15299,N_15372);
and U15594 (N_15594,N_15355,N_15393);
and U15595 (N_15595,N_15354,N_15346);
nand U15596 (N_15596,N_15358,N_15278);
nand U15597 (N_15597,N_15308,N_15249);
nor U15598 (N_15598,N_15326,N_15346);
and U15599 (N_15599,N_15252,N_15399);
nor U15600 (N_15600,N_15517,N_15457);
xor U15601 (N_15601,N_15511,N_15549);
nand U15602 (N_15602,N_15584,N_15513);
or U15603 (N_15603,N_15458,N_15531);
and U15604 (N_15604,N_15523,N_15429);
nand U15605 (N_15605,N_15532,N_15414);
or U15606 (N_15606,N_15569,N_15470);
and U15607 (N_15607,N_15428,N_15502);
xor U15608 (N_15608,N_15504,N_15537);
xnor U15609 (N_15609,N_15555,N_15530);
and U15610 (N_15610,N_15540,N_15560);
or U15611 (N_15611,N_15565,N_15528);
and U15612 (N_15612,N_15475,N_15527);
and U15613 (N_15613,N_15597,N_15587);
nand U15614 (N_15614,N_15455,N_15493);
or U15615 (N_15615,N_15403,N_15407);
and U15616 (N_15616,N_15410,N_15519);
nand U15617 (N_15617,N_15462,N_15417);
nor U15618 (N_15618,N_15592,N_15478);
xnor U15619 (N_15619,N_15481,N_15505);
nor U15620 (N_15620,N_15494,N_15402);
xnor U15621 (N_15621,N_15575,N_15591);
nand U15622 (N_15622,N_15553,N_15415);
xor U15623 (N_15623,N_15421,N_15471);
xor U15624 (N_15624,N_15550,N_15492);
nor U15625 (N_15625,N_15520,N_15413);
nand U15626 (N_15626,N_15525,N_15454);
nand U15627 (N_15627,N_15558,N_15480);
nor U15628 (N_15628,N_15581,N_15408);
nor U15629 (N_15629,N_15518,N_15483);
nand U15630 (N_15630,N_15401,N_15594);
xor U15631 (N_15631,N_15490,N_15541);
xor U15632 (N_15632,N_15524,N_15516);
nand U15633 (N_15633,N_15573,N_15464);
and U15634 (N_15634,N_15445,N_15557);
nor U15635 (N_15635,N_15418,N_15514);
nor U15636 (N_15636,N_15596,N_15497);
xnor U15637 (N_15637,N_15441,N_15499);
nor U15638 (N_15638,N_15500,N_15566);
or U15639 (N_15639,N_15586,N_15585);
nor U15640 (N_15640,N_15437,N_15452);
nor U15641 (N_15641,N_15484,N_15598);
nor U15642 (N_15642,N_15526,N_15595);
or U15643 (N_15643,N_15477,N_15599);
nand U15644 (N_15644,N_15469,N_15577);
nor U15645 (N_15645,N_15488,N_15552);
nand U15646 (N_15646,N_15568,N_15522);
or U15647 (N_15647,N_15486,N_15588);
xnor U15648 (N_15648,N_15442,N_15551);
nand U15649 (N_15649,N_15570,N_15503);
nand U15650 (N_15650,N_15510,N_15456);
xnor U15651 (N_15651,N_15495,N_15479);
nand U15652 (N_15652,N_15539,N_15431);
or U15653 (N_15653,N_15593,N_15554);
nor U15654 (N_15654,N_15512,N_15436);
xor U15655 (N_15655,N_15425,N_15561);
xor U15656 (N_15656,N_15496,N_15461);
nand U15657 (N_15657,N_15485,N_15567);
nor U15658 (N_15658,N_15459,N_15427);
nand U15659 (N_15659,N_15535,N_15571);
nor U15660 (N_15660,N_15433,N_15574);
xor U15661 (N_15661,N_15491,N_15465);
nand U15662 (N_15662,N_15473,N_15444);
nor U15663 (N_15663,N_15533,N_15416);
or U15664 (N_15664,N_15411,N_15424);
and U15665 (N_15665,N_15534,N_15489);
xnor U15666 (N_15666,N_15542,N_15487);
and U15667 (N_15667,N_15590,N_15419);
or U15668 (N_15668,N_15474,N_15468);
and U15669 (N_15669,N_15466,N_15422);
and U15670 (N_15670,N_15546,N_15544);
nor U15671 (N_15671,N_15580,N_15404);
nand U15672 (N_15672,N_15426,N_15547);
nand U15673 (N_15673,N_15508,N_15430);
nor U15674 (N_15674,N_15460,N_15545);
or U15675 (N_15675,N_15451,N_15529);
and U15676 (N_15676,N_15435,N_15423);
xnor U15677 (N_15677,N_15434,N_15507);
or U15678 (N_15678,N_15506,N_15543);
or U15679 (N_15679,N_15521,N_15432);
nor U15680 (N_15680,N_15583,N_15563);
nand U15681 (N_15681,N_15450,N_15440);
xor U15682 (N_15682,N_15405,N_15578);
and U15683 (N_15683,N_15472,N_15446);
nand U15684 (N_15684,N_15572,N_15406);
nor U15685 (N_15685,N_15463,N_15409);
or U15686 (N_15686,N_15559,N_15453);
xnor U15687 (N_15687,N_15443,N_15582);
nor U15688 (N_15688,N_15515,N_15589);
or U15689 (N_15689,N_15562,N_15548);
nand U15690 (N_15690,N_15447,N_15579);
nand U15691 (N_15691,N_15476,N_15536);
or U15692 (N_15692,N_15400,N_15576);
nand U15693 (N_15693,N_15509,N_15448);
nor U15694 (N_15694,N_15556,N_15449);
nand U15695 (N_15695,N_15498,N_15438);
and U15696 (N_15696,N_15467,N_15564);
or U15697 (N_15697,N_15420,N_15482);
and U15698 (N_15698,N_15439,N_15538);
xor U15699 (N_15699,N_15412,N_15501);
nand U15700 (N_15700,N_15426,N_15513);
and U15701 (N_15701,N_15486,N_15466);
or U15702 (N_15702,N_15591,N_15511);
or U15703 (N_15703,N_15435,N_15466);
nand U15704 (N_15704,N_15447,N_15467);
and U15705 (N_15705,N_15407,N_15521);
or U15706 (N_15706,N_15559,N_15555);
and U15707 (N_15707,N_15472,N_15559);
or U15708 (N_15708,N_15597,N_15582);
and U15709 (N_15709,N_15488,N_15529);
or U15710 (N_15710,N_15407,N_15501);
and U15711 (N_15711,N_15569,N_15481);
or U15712 (N_15712,N_15471,N_15595);
or U15713 (N_15713,N_15594,N_15506);
and U15714 (N_15714,N_15442,N_15507);
xnor U15715 (N_15715,N_15542,N_15598);
nor U15716 (N_15716,N_15419,N_15575);
xnor U15717 (N_15717,N_15527,N_15425);
nand U15718 (N_15718,N_15598,N_15526);
and U15719 (N_15719,N_15471,N_15539);
nor U15720 (N_15720,N_15490,N_15496);
xnor U15721 (N_15721,N_15494,N_15412);
and U15722 (N_15722,N_15470,N_15545);
xor U15723 (N_15723,N_15533,N_15562);
or U15724 (N_15724,N_15524,N_15596);
xnor U15725 (N_15725,N_15573,N_15506);
nor U15726 (N_15726,N_15480,N_15486);
or U15727 (N_15727,N_15477,N_15595);
or U15728 (N_15728,N_15472,N_15509);
or U15729 (N_15729,N_15532,N_15558);
nor U15730 (N_15730,N_15443,N_15567);
xnor U15731 (N_15731,N_15524,N_15471);
or U15732 (N_15732,N_15495,N_15478);
or U15733 (N_15733,N_15509,N_15426);
and U15734 (N_15734,N_15558,N_15477);
or U15735 (N_15735,N_15544,N_15577);
nor U15736 (N_15736,N_15502,N_15421);
nor U15737 (N_15737,N_15517,N_15425);
and U15738 (N_15738,N_15532,N_15550);
nor U15739 (N_15739,N_15404,N_15494);
xnor U15740 (N_15740,N_15556,N_15588);
xnor U15741 (N_15741,N_15524,N_15518);
and U15742 (N_15742,N_15410,N_15451);
nor U15743 (N_15743,N_15574,N_15510);
nand U15744 (N_15744,N_15506,N_15576);
nor U15745 (N_15745,N_15571,N_15404);
xor U15746 (N_15746,N_15551,N_15400);
and U15747 (N_15747,N_15466,N_15427);
or U15748 (N_15748,N_15474,N_15426);
or U15749 (N_15749,N_15547,N_15535);
nor U15750 (N_15750,N_15538,N_15416);
and U15751 (N_15751,N_15452,N_15593);
or U15752 (N_15752,N_15479,N_15440);
and U15753 (N_15753,N_15444,N_15424);
and U15754 (N_15754,N_15557,N_15489);
and U15755 (N_15755,N_15577,N_15531);
nor U15756 (N_15756,N_15495,N_15552);
xor U15757 (N_15757,N_15499,N_15502);
nand U15758 (N_15758,N_15514,N_15580);
or U15759 (N_15759,N_15508,N_15518);
xnor U15760 (N_15760,N_15559,N_15468);
and U15761 (N_15761,N_15437,N_15442);
xnor U15762 (N_15762,N_15564,N_15455);
or U15763 (N_15763,N_15580,N_15462);
xor U15764 (N_15764,N_15515,N_15595);
nand U15765 (N_15765,N_15541,N_15567);
xor U15766 (N_15766,N_15563,N_15410);
or U15767 (N_15767,N_15563,N_15559);
xnor U15768 (N_15768,N_15498,N_15419);
xor U15769 (N_15769,N_15565,N_15502);
and U15770 (N_15770,N_15428,N_15527);
nor U15771 (N_15771,N_15416,N_15596);
nand U15772 (N_15772,N_15408,N_15412);
or U15773 (N_15773,N_15575,N_15467);
nor U15774 (N_15774,N_15436,N_15416);
and U15775 (N_15775,N_15457,N_15449);
or U15776 (N_15776,N_15523,N_15573);
nor U15777 (N_15777,N_15439,N_15485);
nand U15778 (N_15778,N_15532,N_15404);
nor U15779 (N_15779,N_15428,N_15412);
and U15780 (N_15780,N_15445,N_15548);
nand U15781 (N_15781,N_15481,N_15513);
xor U15782 (N_15782,N_15430,N_15557);
nand U15783 (N_15783,N_15576,N_15579);
nand U15784 (N_15784,N_15509,N_15444);
or U15785 (N_15785,N_15584,N_15400);
and U15786 (N_15786,N_15554,N_15557);
and U15787 (N_15787,N_15570,N_15578);
nand U15788 (N_15788,N_15508,N_15475);
nand U15789 (N_15789,N_15592,N_15403);
nand U15790 (N_15790,N_15456,N_15552);
or U15791 (N_15791,N_15560,N_15584);
or U15792 (N_15792,N_15576,N_15577);
nand U15793 (N_15793,N_15457,N_15450);
or U15794 (N_15794,N_15594,N_15482);
or U15795 (N_15795,N_15498,N_15425);
or U15796 (N_15796,N_15485,N_15463);
xnor U15797 (N_15797,N_15452,N_15526);
nand U15798 (N_15798,N_15522,N_15524);
and U15799 (N_15799,N_15553,N_15426);
xnor U15800 (N_15800,N_15663,N_15785);
xnor U15801 (N_15801,N_15707,N_15726);
or U15802 (N_15802,N_15610,N_15638);
nand U15803 (N_15803,N_15654,N_15791);
nor U15804 (N_15804,N_15792,N_15781);
xor U15805 (N_15805,N_15754,N_15666);
or U15806 (N_15806,N_15614,N_15772);
nand U15807 (N_15807,N_15661,N_15715);
xor U15808 (N_15808,N_15716,N_15780);
nand U15809 (N_15809,N_15643,N_15681);
nand U15810 (N_15810,N_15758,N_15778);
or U15811 (N_15811,N_15668,N_15602);
and U15812 (N_15812,N_15784,N_15692);
nand U15813 (N_15813,N_15753,N_15672);
and U15814 (N_15814,N_15739,N_15600);
xnor U15815 (N_15815,N_15775,N_15748);
xnor U15816 (N_15816,N_15623,N_15777);
nand U15817 (N_15817,N_15757,N_15679);
nor U15818 (N_15818,N_15616,N_15636);
and U15819 (N_15819,N_15669,N_15608);
nand U15820 (N_15820,N_15655,N_15651);
nand U15821 (N_15821,N_15765,N_15653);
or U15822 (N_15822,N_15646,N_15787);
nor U15823 (N_15823,N_15698,N_15708);
xnor U15824 (N_15824,N_15677,N_15720);
xnor U15825 (N_15825,N_15719,N_15635);
and U15826 (N_15826,N_15745,N_15704);
nor U15827 (N_15827,N_15664,N_15718);
and U15828 (N_15828,N_15671,N_15620);
nor U15829 (N_15829,N_15680,N_15640);
and U15830 (N_15830,N_15710,N_15702);
xor U15831 (N_15831,N_15617,N_15604);
and U15832 (N_15832,N_15737,N_15639);
or U15833 (N_15833,N_15798,N_15774);
nand U15834 (N_15834,N_15606,N_15621);
xor U15835 (N_15835,N_15697,N_15634);
xor U15836 (N_15836,N_15625,N_15794);
nor U15837 (N_15837,N_15797,N_15776);
nor U15838 (N_15838,N_15725,N_15699);
nand U15839 (N_15839,N_15722,N_15603);
xor U15840 (N_15840,N_15733,N_15647);
nor U15841 (N_15841,N_15741,N_15767);
or U15842 (N_15842,N_15632,N_15788);
and U15843 (N_15843,N_15619,N_15690);
nor U15844 (N_15844,N_15644,N_15609);
nand U15845 (N_15845,N_15601,N_15717);
and U15846 (N_15846,N_15631,N_15796);
xor U15847 (N_15847,N_15789,N_15649);
and U15848 (N_15848,N_15626,N_15721);
and U15849 (N_15849,N_15761,N_15607);
nand U15850 (N_15850,N_15770,N_15762);
xnor U15851 (N_15851,N_15645,N_15764);
xnor U15852 (N_15852,N_15740,N_15714);
nand U15853 (N_15853,N_15746,N_15799);
and U15854 (N_15854,N_15633,N_15605);
and U15855 (N_15855,N_15766,N_15695);
or U15856 (N_15856,N_15712,N_15760);
and U15857 (N_15857,N_15612,N_15627);
nand U15858 (N_15858,N_15637,N_15750);
and U15859 (N_15859,N_15658,N_15769);
nand U15860 (N_15860,N_15685,N_15759);
nand U15861 (N_15861,N_15755,N_15657);
xnor U15862 (N_15862,N_15687,N_15738);
and U15863 (N_15863,N_15711,N_15656);
or U15864 (N_15864,N_15706,N_15684);
or U15865 (N_15865,N_15662,N_15630);
nor U15866 (N_15866,N_15786,N_15650);
nand U15867 (N_15867,N_15670,N_15703);
xor U15868 (N_15868,N_15727,N_15756);
nor U15869 (N_15869,N_15743,N_15652);
or U15870 (N_15870,N_15613,N_15729);
and U15871 (N_15871,N_15779,N_15782);
and U15872 (N_15872,N_15783,N_15675);
and U15873 (N_15873,N_15624,N_15660);
nor U15874 (N_15874,N_15676,N_15709);
and U15875 (N_15875,N_15795,N_15689);
and U15876 (N_15876,N_15701,N_15730);
xor U15877 (N_15877,N_15773,N_15629);
or U15878 (N_15878,N_15628,N_15642);
or U15879 (N_15879,N_15744,N_15691);
xnor U15880 (N_15880,N_15688,N_15622);
nand U15881 (N_15881,N_15763,N_15752);
xnor U15882 (N_15882,N_15734,N_15700);
nor U15883 (N_15883,N_15686,N_15705);
nor U15884 (N_15884,N_15731,N_15682);
or U15885 (N_15885,N_15611,N_15641);
or U15886 (N_15886,N_15768,N_15615);
nor U15887 (N_15887,N_15793,N_15667);
or U15888 (N_15888,N_15732,N_15683);
xnor U15889 (N_15889,N_15724,N_15648);
nor U15890 (N_15890,N_15735,N_15674);
or U15891 (N_15891,N_15673,N_15665);
xnor U15892 (N_15892,N_15771,N_15728);
or U15893 (N_15893,N_15747,N_15678);
nand U15894 (N_15894,N_15723,N_15693);
nand U15895 (N_15895,N_15749,N_15742);
or U15896 (N_15896,N_15659,N_15696);
and U15897 (N_15897,N_15694,N_15618);
xnor U15898 (N_15898,N_15790,N_15751);
xnor U15899 (N_15899,N_15736,N_15713);
or U15900 (N_15900,N_15645,N_15733);
xor U15901 (N_15901,N_15650,N_15736);
nand U15902 (N_15902,N_15697,N_15744);
nor U15903 (N_15903,N_15604,N_15600);
xor U15904 (N_15904,N_15676,N_15625);
nand U15905 (N_15905,N_15658,N_15731);
nand U15906 (N_15906,N_15759,N_15761);
xor U15907 (N_15907,N_15693,N_15726);
or U15908 (N_15908,N_15675,N_15786);
or U15909 (N_15909,N_15700,N_15785);
or U15910 (N_15910,N_15716,N_15730);
or U15911 (N_15911,N_15754,N_15605);
nand U15912 (N_15912,N_15713,N_15663);
and U15913 (N_15913,N_15739,N_15702);
and U15914 (N_15914,N_15649,N_15660);
xnor U15915 (N_15915,N_15686,N_15733);
and U15916 (N_15916,N_15655,N_15760);
or U15917 (N_15917,N_15753,N_15768);
nand U15918 (N_15918,N_15656,N_15629);
xnor U15919 (N_15919,N_15667,N_15690);
xor U15920 (N_15920,N_15758,N_15650);
xnor U15921 (N_15921,N_15643,N_15741);
or U15922 (N_15922,N_15682,N_15647);
nor U15923 (N_15923,N_15694,N_15732);
or U15924 (N_15924,N_15632,N_15674);
or U15925 (N_15925,N_15684,N_15712);
xor U15926 (N_15926,N_15737,N_15755);
nand U15927 (N_15927,N_15765,N_15725);
nor U15928 (N_15928,N_15618,N_15624);
xor U15929 (N_15929,N_15789,N_15643);
xnor U15930 (N_15930,N_15750,N_15722);
nand U15931 (N_15931,N_15669,N_15774);
nor U15932 (N_15932,N_15601,N_15659);
and U15933 (N_15933,N_15782,N_15780);
and U15934 (N_15934,N_15716,N_15674);
and U15935 (N_15935,N_15699,N_15762);
xnor U15936 (N_15936,N_15740,N_15626);
xnor U15937 (N_15937,N_15777,N_15751);
nor U15938 (N_15938,N_15639,N_15671);
and U15939 (N_15939,N_15712,N_15783);
and U15940 (N_15940,N_15607,N_15744);
xnor U15941 (N_15941,N_15741,N_15647);
xor U15942 (N_15942,N_15738,N_15618);
or U15943 (N_15943,N_15771,N_15625);
nand U15944 (N_15944,N_15648,N_15686);
xnor U15945 (N_15945,N_15786,N_15719);
nand U15946 (N_15946,N_15642,N_15735);
nand U15947 (N_15947,N_15665,N_15663);
and U15948 (N_15948,N_15604,N_15647);
nand U15949 (N_15949,N_15688,N_15765);
xor U15950 (N_15950,N_15643,N_15653);
and U15951 (N_15951,N_15607,N_15782);
nor U15952 (N_15952,N_15657,N_15610);
nand U15953 (N_15953,N_15658,N_15705);
or U15954 (N_15954,N_15687,N_15723);
xnor U15955 (N_15955,N_15660,N_15712);
or U15956 (N_15956,N_15778,N_15769);
or U15957 (N_15957,N_15756,N_15677);
nand U15958 (N_15958,N_15713,N_15672);
xor U15959 (N_15959,N_15638,N_15763);
xnor U15960 (N_15960,N_15772,N_15699);
and U15961 (N_15961,N_15762,N_15629);
nor U15962 (N_15962,N_15631,N_15774);
xnor U15963 (N_15963,N_15772,N_15602);
or U15964 (N_15964,N_15682,N_15673);
or U15965 (N_15965,N_15775,N_15751);
nor U15966 (N_15966,N_15688,N_15678);
nor U15967 (N_15967,N_15756,N_15683);
xnor U15968 (N_15968,N_15718,N_15713);
xnor U15969 (N_15969,N_15600,N_15744);
and U15970 (N_15970,N_15717,N_15673);
or U15971 (N_15971,N_15613,N_15601);
or U15972 (N_15972,N_15796,N_15687);
nor U15973 (N_15973,N_15656,N_15736);
nor U15974 (N_15974,N_15704,N_15630);
nand U15975 (N_15975,N_15646,N_15672);
nor U15976 (N_15976,N_15741,N_15652);
and U15977 (N_15977,N_15797,N_15796);
nand U15978 (N_15978,N_15635,N_15740);
nor U15979 (N_15979,N_15662,N_15726);
nand U15980 (N_15980,N_15648,N_15612);
and U15981 (N_15981,N_15689,N_15718);
nor U15982 (N_15982,N_15740,N_15769);
and U15983 (N_15983,N_15741,N_15644);
xnor U15984 (N_15984,N_15717,N_15742);
nand U15985 (N_15985,N_15629,N_15611);
xor U15986 (N_15986,N_15605,N_15622);
nor U15987 (N_15987,N_15691,N_15778);
nor U15988 (N_15988,N_15760,N_15603);
nand U15989 (N_15989,N_15634,N_15677);
xnor U15990 (N_15990,N_15684,N_15750);
xnor U15991 (N_15991,N_15776,N_15746);
and U15992 (N_15992,N_15707,N_15681);
nand U15993 (N_15993,N_15629,N_15691);
xor U15994 (N_15994,N_15710,N_15791);
nor U15995 (N_15995,N_15623,N_15667);
xnor U15996 (N_15996,N_15729,N_15618);
nand U15997 (N_15997,N_15666,N_15712);
and U15998 (N_15998,N_15797,N_15788);
nor U15999 (N_15999,N_15676,N_15703);
nor U16000 (N_16000,N_15865,N_15959);
nor U16001 (N_16001,N_15931,N_15935);
and U16002 (N_16002,N_15958,N_15816);
and U16003 (N_16003,N_15966,N_15915);
xnor U16004 (N_16004,N_15900,N_15985);
xnor U16005 (N_16005,N_15812,N_15993);
xnor U16006 (N_16006,N_15882,N_15911);
nor U16007 (N_16007,N_15851,N_15973);
nand U16008 (N_16008,N_15848,N_15908);
nor U16009 (N_16009,N_15877,N_15844);
and U16010 (N_16010,N_15879,N_15946);
and U16011 (N_16011,N_15841,N_15929);
and U16012 (N_16012,N_15912,N_15863);
nand U16013 (N_16013,N_15916,N_15939);
nor U16014 (N_16014,N_15853,N_15962);
xnor U16015 (N_16015,N_15917,N_15855);
nor U16016 (N_16016,N_15803,N_15892);
or U16017 (N_16017,N_15872,N_15899);
xnor U16018 (N_16018,N_15923,N_15997);
and U16019 (N_16019,N_15876,N_15839);
nand U16020 (N_16020,N_15901,N_15984);
and U16021 (N_16021,N_15963,N_15913);
nor U16022 (N_16022,N_15944,N_15989);
and U16023 (N_16023,N_15971,N_15887);
nand U16024 (N_16024,N_15978,N_15981);
nand U16025 (N_16025,N_15858,N_15996);
nand U16026 (N_16026,N_15988,N_15833);
nand U16027 (N_16027,N_15820,N_15895);
nor U16028 (N_16028,N_15807,N_15821);
or U16029 (N_16029,N_15874,N_15834);
and U16030 (N_16030,N_15842,N_15804);
nand U16031 (N_16031,N_15875,N_15802);
and U16032 (N_16032,N_15897,N_15932);
or U16033 (N_16033,N_15925,N_15822);
nand U16034 (N_16034,N_15983,N_15856);
nand U16035 (N_16035,N_15961,N_15881);
xor U16036 (N_16036,N_15960,N_15825);
or U16037 (N_16037,N_15954,N_15835);
nor U16038 (N_16038,N_15927,N_15933);
and U16039 (N_16039,N_15808,N_15850);
nand U16040 (N_16040,N_15937,N_15813);
nor U16041 (N_16041,N_15995,N_15878);
nand U16042 (N_16042,N_15823,N_15871);
xnor U16043 (N_16043,N_15953,N_15936);
and U16044 (N_16044,N_15970,N_15806);
xor U16045 (N_16045,N_15950,N_15969);
nor U16046 (N_16046,N_15906,N_15827);
nor U16047 (N_16047,N_15938,N_15898);
xnor U16048 (N_16048,N_15809,N_15905);
and U16049 (N_16049,N_15964,N_15991);
nor U16050 (N_16050,N_15829,N_15884);
xor U16051 (N_16051,N_15949,N_15818);
xnor U16052 (N_16052,N_15843,N_15928);
xnor U16053 (N_16053,N_15854,N_15845);
or U16054 (N_16054,N_15891,N_15947);
nor U16055 (N_16055,N_15998,N_15860);
and U16056 (N_16056,N_15919,N_15987);
nand U16057 (N_16057,N_15893,N_15999);
nand U16058 (N_16058,N_15904,N_15976);
nor U16059 (N_16059,N_15975,N_15914);
nor U16060 (N_16060,N_15907,N_15942);
nor U16061 (N_16061,N_15889,N_15926);
and U16062 (N_16062,N_15979,N_15885);
and U16063 (N_16063,N_15943,N_15890);
or U16064 (N_16064,N_15852,N_15956);
and U16065 (N_16065,N_15918,N_15861);
and U16066 (N_16066,N_15934,N_15817);
and U16067 (N_16067,N_15952,N_15994);
nor U16068 (N_16068,N_15977,N_15832);
xnor U16069 (N_16069,N_15986,N_15837);
or U16070 (N_16070,N_15849,N_15870);
xor U16071 (N_16071,N_15824,N_15868);
or U16072 (N_16072,N_15800,N_15948);
nor U16073 (N_16073,N_15838,N_15846);
nand U16074 (N_16074,N_15840,N_15862);
or U16075 (N_16075,N_15924,N_15883);
and U16076 (N_16076,N_15992,N_15967);
xnor U16077 (N_16077,N_15888,N_15894);
nand U16078 (N_16078,N_15880,N_15819);
or U16079 (N_16079,N_15869,N_15968);
and U16080 (N_16080,N_15921,N_15940);
or U16081 (N_16081,N_15990,N_15859);
nand U16082 (N_16082,N_15920,N_15836);
xor U16083 (N_16083,N_15815,N_15903);
nor U16084 (N_16084,N_15867,N_15805);
nor U16085 (N_16085,N_15866,N_15982);
nor U16086 (N_16086,N_15873,N_15941);
nor U16087 (N_16087,N_15811,N_15896);
nand U16088 (N_16088,N_15810,N_15831);
nor U16089 (N_16089,N_15910,N_15828);
xnor U16090 (N_16090,N_15857,N_15930);
and U16091 (N_16091,N_15801,N_15826);
and U16092 (N_16092,N_15955,N_15945);
xor U16093 (N_16093,N_15830,N_15974);
nand U16094 (N_16094,N_15951,N_15957);
and U16095 (N_16095,N_15902,N_15922);
and U16096 (N_16096,N_15814,N_15886);
xnor U16097 (N_16097,N_15864,N_15965);
nand U16098 (N_16098,N_15972,N_15980);
nor U16099 (N_16099,N_15909,N_15847);
nand U16100 (N_16100,N_15931,N_15958);
or U16101 (N_16101,N_15957,N_15914);
nor U16102 (N_16102,N_15957,N_15930);
nor U16103 (N_16103,N_15862,N_15981);
or U16104 (N_16104,N_15991,N_15979);
and U16105 (N_16105,N_15956,N_15884);
xor U16106 (N_16106,N_15908,N_15949);
nor U16107 (N_16107,N_15949,N_15803);
nand U16108 (N_16108,N_15983,N_15802);
nand U16109 (N_16109,N_15993,N_15944);
or U16110 (N_16110,N_15995,N_15966);
nor U16111 (N_16111,N_15967,N_15898);
nand U16112 (N_16112,N_15816,N_15993);
nand U16113 (N_16113,N_15921,N_15806);
xor U16114 (N_16114,N_15910,N_15872);
nor U16115 (N_16115,N_15948,N_15819);
xnor U16116 (N_16116,N_15926,N_15803);
nand U16117 (N_16117,N_15914,N_15948);
nor U16118 (N_16118,N_15867,N_15983);
nor U16119 (N_16119,N_15852,N_15906);
nor U16120 (N_16120,N_15934,N_15842);
nand U16121 (N_16121,N_15876,N_15918);
nor U16122 (N_16122,N_15992,N_15979);
and U16123 (N_16123,N_15879,N_15880);
and U16124 (N_16124,N_15957,N_15811);
xnor U16125 (N_16125,N_15980,N_15912);
nand U16126 (N_16126,N_15901,N_15933);
and U16127 (N_16127,N_15809,N_15826);
nor U16128 (N_16128,N_15836,N_15958);
nor U16129 (N_16129,N_15940,N_15970);
nand U16130 (N_16130,N_15944,N_15970);
nor U16131 (N_16131,N_15963,N_15894);
nor U16132 (N_16132,N_15936,N_15805);
xnor U16133 (N_16133,N_15839,N_15912);
nor U16134 (N_16134,N_15836,N_15849);
nand U16135 (N_16135,N_15839,N_15875);
nand U16136 (N_16136,N_15885,N_15963);
xnor U16137 (N_16137,N_15862,N_15982);
nand U16138 (N_16138,N_15847,N_15811);
nand U16139 (N_16139,N_15851,N_15808);
nor U16140 (N_16140,N_15897,N_15814);
or U16141 (N_16141,N_15948,N_15925);
xnor U16142 (N_16142,N_15886,N_15900);
nand U16143 (N_16143,N_15878,N_15961);
and U16144 (N_16144,N_15850,N_15822);
xor U16145 (N_16145,N_15904,N_15847);
nand U16146 (N_16146,N_15923,N_15914);
and U16147 (N_16147,N_15889,N_15913);
nand U16148 (N_16148,N_15970,N_15891);
or U16149 (N_16149,N_15981,N_15865);
and U16150 (N_16150,N_15928,N_15804);
and U16151 (N_16151,N_15958,N_15834);
and U16152 (N_16152,N_15960,N_15993);
or U16153 (N_16153,N_15993,N_15804);
nand U16154 (N_16154,N_15876,N_15813);
or U16155 (N_16155,N_15854,N_15827);
nor U16156 (N_16156,N_15894,N_15847);
nor U16157 (N_16157,N_15841,N_15951);
and U16158 (N_16158,N_15881,N_15815);
nand U16159 (N_16159,N_15926,N_15911);
nor U16160 (N_16160,N_15866,N_15951);
or U16161 (N_16161,N_15963,N_15825);
nand U16162 (N_16162,N_15945,N_15941);
nand U16163 (N_16163,N_15954,N_15836);
nand U16164 (N_16164,N_15885,N_15946);
nand U16165 (N_16165,N_15934,N_15895);
nand U16166 (N_16166,N_15889,N_15834);
and U16167 (N_16167,N_15831,N_15853);
nand U16168 (N_16168,N_15890,N_15884);
and U16169 (N_16169,N_15869,N_15836);
nand U16170 (N_16170,N_15965,N_15916);
nand U16171 (N_16171,N_15843,N_15956);
xnor U16172 (N_16172,N_15860,N_15945);
and U16173 (N_16173,N_15870,N_15987);
nand U16174 (N_16174,N_15954,N_15953);
or U16175 (N_16175,N_15839,N_15928);
and U16176 (N_16176,N_15925,N_15869);
nand U16177 (N_16177,N_15944,N_15997);
and U16178 (N_16178,N_15811,N_15978);
nor U16179 (N_16179,N_15860,N_15949);
and U16180 (N_16180,N_15838,N_15815);
nand U16181 (N_16181,N_15816,N_15995);
or U16182 (N_16182,N_15803,N_15948);
nor U16183 (N_16183,N_15915,N_15811);
nand U16184 (N_16184,N_15918,N_15941);
or U16185 (N_16185,N_15880,N_15914);
and U16186 (N_16186,N_15847,N_15851);
xor U16187 (N_16187,N_15954,N_15895);
nor U16188 (N_16188,N_15856,N_15968);
and U16189 (N_16189,N_15949,N_15964);
xor U16190 (N_16190,N_15833,N_15875);
xnor U16191 (N_16191,N_15937,N_15861);
or U16192 (N_16192,N_15812,N_15816);
and U16193 (N_16193,N_15890,N_15802);
nand U16194 (N_16194,N_15827,N_15810);
nand U16195 (N_16195,N_15942,N_15997);
or U16196 (N_16196,N_15809,N_15948);
and U16197 (N_16197,N_15856,N_15824);
and U16198 (N_16198,N_15946,N_15802);
nand U16199 (N_16199,N_15851,N_15984);
nand U16200 (N_16200,N_16107,N_16019);
xor U16201 (N_16201,N_16101,N_16116);
xnor U16202 (N_16202,N_16035,N_16095);
xor U16203 (N_16203,N_16050,N_16068);
and U16204 (N_16204,N_16181,N_16125);
and U16205 (N_16205,N_16110,N_16184);
and U16206 (N_16206,N_16166,N_16194);
or U16207 (N_16207,N_16142,N_16039);
and U16208 (N_16208,N_16008,N_16165);
nand U16209 (N_16209,N_16078,N_16069);
nand U16210 (N_16210,N_16090,N_16012);
xnor U16211 (N_16211,N_16033,N_16026);
xor U16212 (N_16212,N_16132,N_16042);
xor U16213 (N_16213,N_16156,N_16126);
xnor U16214 (N_16214,N_16017,N_16048);
xor U16215 (N_16215,N_16179,N_16081);
and U16216 (N_16216,N_16106,N_16054);
nor U16217 (N_16217,N_16047,N_16161);
nor U16218 (N_16218,N_16056,N_16046);
or U16219 (N_16219,N_16010,N_16115);
or U16220 (N_16220,N_16134,N_16123);
nand U16221 (N_16221,N_16004,N_16169);
and U16222 (N_16222,N_16024,N_16025);
nor U16223 (N_16223,N_16183,N_16109);
and U16224 (N_16224,N_16067,N_16015);
nor U16225 (N_16225,N_16009,N_16141);
nand U16226 (N_16226,N_16092,N_16160);
or U16227 (N_16227,N_16199,N_16139);
nor U16228 (N_16228,N_16173,N_16167);
or U16229 (N_16229,N_16103,N_16076);
nand U16230 (N_16230,N_16040,N_16182);
xnor U16231 (N_16231,N_16117,N_16195);
xnor U16232 (N_16232,N_16000,N_16120);
xnor U16233 (N_16233,N_16105,N_16062);
nand U16234 (N_16234,N_16197,N_16122);
nand U16235 (N_16235,N_16079,N_16029);
nor U16236 (N_16236,N_16053,N_16178);
nand U16237 (N_16237,N_16086,N_16074);
xor U16238 (N_16238,N_16108,N_16001);
or U16239 (N_16239,N_16177,N_16154);
nor U16240 (N_16240,N_16072,N_16133);
and U16241 (N_16241,N_16070,N_16073);
nor U16242 (N_16242,N_16121,N_16005);
or U16243 (N_16243,N_16096,N_16028);
or U16244 (N_16244,N_16151,N_16027);
and U16245 (N_16245,N_16097,N_16152);
and U16246 (N_16246,N_16051,N_16148);
and U16247 (N_16247,N_16082,N_16087);
nor U16248 (N_16248,N_16061,N_16185);
or U16249 (N_16249,N_16145,N_16146);
and U16250 (N_16250,N_16135,N_16155);
nand U16251 (N_16251,N_16031,N_16071);
nor U16252 (N_16252,N_16118,N_16006);
nand U16253 (N_16253,N_16124,N_16021);
nand U16254 (N_16254,N_16162,N_16180);
nor U16255 (N_16255,N_16198,N_16007);
and U16256 (N_16256,N_16044,N_16144);
and U16257 (N_16257,N_16085,N_16022);
and U16258 (N_16258,N_16127,N_16052);
xor U16259 (N_16259,N_16164,N_16131);
or U16260 (N_16260,N_16196,N_16112);
nor U16261 (N_16261,N_16191,N_16045);
or U16262 (N_16262,N_16037,N_16058);
and U16263 (N_16263,N_16030,N_16114);
nand U16264 (N_16264,N_16088,N_16113);
nor U16265 (N_16265,N_16102,N_16168);
xnor U16266 (N_16266,N_16143,N_16111);
and U16267 (N_16267,N_16077,N_16041);
nor U16268 (N_16268,N_16098,N_16020);
nand U16269 (N_16269,N_16034,N_16055);
xor U16270 (N_16270,N_16036,N_16100);
xnor U16271 (N_16271,N_16170,N_16064);
and U16272 (N_16272,N_16130,N_16032);
and U16273 (N_16273,N_16128,N_16014);
xnor U16274 (N_16274,N_16003,N_16002);
or U16275 (N_16275,N_16150,N_16091);
xnor U16276 (N_16276,N_16171,N_16119);
and U16277 (N_16277,N_16149,N_16172);
and U16278 (N_16278,N_16136,N_16057);
nor U16279 (N_16279,N_16147,N_16129);
and U16280 (N_16280,N_16093,N_16016);
xnor U16281 (N_16281,N_16189,N_16065);
and U16282 (N_16282,N_16080,N_16188);
and U16283 (N_16283,N_16163,N_16138);
nand U16284 (N_16284,N_16193,N_16099);
or U16285 (N_16285,N_16083,N_16190);
and U16286 (N_16286,N_16140,N_16013);
xor U16287 (N_16287,N_16159,N_16187);
xnor U16288 (N_16288,N_16094,N_16104);
and U16289 (N_16289,N_16089,N_16043);
or U16290 (N_16290,N_16075,N_16063);
or U16291 (N_16291,N_16011,N_16192);
or U16292 (N_16292,N_16157,N_16023);
and U16293 (N_16293,N_16084,N_16137);
xor U16294 (N_16294,N_16176,N_16018);
nand U16295 (N_16295,N_16060,N_16049);
xnor U16296 (N_16296,N_16186,N_16066);
or U16297 (N_16297,N_16153,N_16059);
and U16298 (N_16298,N_16175,N_16038);
nor U16299 (N_16299,N_16174,N_16158);
and U16300 (N_16300,N_16164,N_16146);
xnor U16301 (N_16301,N_16050,N_16166);
xnor U16302 (N_16302,N_16032,N_16022);
or U16303 (N_16303,N_16041,N_16121);
nor U16304 (N_16304,N_16189,N_16107);
or U16305 (N_16305,N_16040,N_16039);
and U16306 (N_16306,N_16064,N_16072);
nor U16307 (N_16307,N_16146,N_16049);
nand U16308 (N_16308,N_16195,N_16179);
or U16309 (N_16309,N_16115,N_16192);
nand U16310 (N_16310,N_16175,N_16075);
nor U16311 (N_16311,N_16114,N_16096);
or U16312 (N_16312,N_16178,N_16071);
xor U16313 (N_16313,N_16035,N_16051);
or U16314 (N_16314,N_16149,N_16039);
or U16315 (N_16315,N_16074,N_16131);
xnor U16316 (N_16316,N_16089,N_16153);
xor U16317 (N_16317,N_16179,N_16171);
nor U16318 (N_16318,N_16051,N_16047);
nand U16319 (N_16319,N_16058,N_16109);
xor U16320 (N_16320,N_16050,N_16035);
or U16321 (N_16321,N_16179,N_16042);
or U16322 (N_16322,N_16186,N_16152);
nor U16323 (N_16323,N_16031,N_16053);
xor U16324 (N_16324,N_16103,N_16173);
or U16325 (N_16325,N_16152,N_16174);
nand U16326 (N_16326,N_16017,N_16014);
or U16327 (N_16327,N_16177,N_16173);
nand U16328 (N_16328,N_16157,N_16134);
nor U16329 (N_16329,N_16125,N_16186);
xor U16330 (N_16330,N_16072,N_16008);
nand U16331 (N_16331,N_16104,N_16024);
and U16332 (N_16332,N_16154,N_16132);
and U16333 (N_16333,N_16035,N_16010);
or U16334 (N_16334,N_16187,N_16113);
nor U16335 (N_16335,N_16068,N_16082);
xnor U16336 (N_16336,N_16177,N_16081);
and U16337 (N_16337,N_16187,N_16016);
and U16338 (N_16338,N_16092,N_16076);
xnor U16339 (N_16339,N_16178,N_16028);
xnor U16340 (N_16340,N_16117,N_16141);
or U16341 (N_16341,N_16189,N_16159);
xnor U16342 (N_16342,N_16062,N_16033);
nor U16343 (N_16343,N_16106,N_16124);
nor U16344 (N_16344,N_16049,N_16161);
and U16345 (N_16345,N_16017,N_16167);
nand U16346 (N_16346,N_16029,N_16154);
xor U16347 (N_16347,N_16096,N_16034);
nor U16348 (N_16348,N_16072,N_16134);
nand U16349 (N_16349,N_16139,N_16136);
nor U16350 (N_16350,N_16037,N_16171);
nor U16351 (N_16351,N_16018,N_16118);
nand U16352 (N_16352,N_16158,N_16117);
nand U16353 (N_16353,N_16038,N_16139);
nor U16354 (N_16354,N_16080,N_16079);
and U16355 (N_16355,N_16011,N_16013);
xnor U16356 (N_16356,N_16179,N_16016);
or U16357 (N_16357,N_16110,N_16047);
xor U16358 (N_16358,N_16089,N_16044);
xor U16359 (N_16359,N_16189,N_16171);
nand U16360 (N_16360,N_16076,N_16097);
or U16361 (N_16361,N_16029,N_16174);
or U16362 (N_16362,N_16075,N_16162);
xnor U16363 (N_16363,N_16115,N_16144);
or U16364 (N_16364,N_16014,N_16186);
and U16365 (N_16365,N_16007,N_16071);
and U16366 (N_16366,N_16095,N_16117);
and U16367 (N_16367,N_16038,N_16196);
nand U16368 (N_16368,N_16064,N_16020);
and U16369 (N_16369,N_16023,N_16180);
or U16370 (N_16370,N_16021,N_16123);
or U16371 (N_16371,N_16107,N_16138);
xor U16372 (N_16372,N_16157,N_16173);
and U16373 (N_16373,N_16195,N_16104);
nand U16374 (N_16374,N_16110,N_16192);
nor U16375 (N_16375,N_16069,N_16144);
xor U16376 (N_16376,N_16002,N_16100);
nand U16377 (N_16377,N_16179,N_16029);
or U16378 (N_16378,N_16113,N_16161);
or U16379 (N_16379,N_16002,N_16102);
nand U16380 (N_16380,N_16051,N_16178);
or U16381 (N_16381,N_16165,N_16027);
nor U16382 (N_16382,N_16148,N_16087);
nor U16383 (N_16383,N_16144,N_16105);
and U16384 (N_16384,N_16114,N_16039);
nor U16385 (N_16385,N_16099,N_16168);
and U16386 (N_16386,N_16073,N_16122);
nor U16387 (N_16387,N_16193,N_16055);
or U16388 (N_16388,N_16113,N_16072);
or U16389 (N_16389,N_16119,N_16073);
or U16390 (N_16390,N_16146,N_16149);
xor U16391 (N_16391,N_16061,N_16057);
xnor U16392 (N_16392,N_16012,N_16051);
nor U16393 (N_16393,N_16186,N_16049);
nor U16394 (N_16394,N_16058,N_16069);
nand U16395 (N_16395,N_16178,N_16166);
and U16396 (N_16396,N_16149,N_16092);
nor U16397 (N_16397,N_16099,N_16008);
and U16398 (N_16398,N_16170,N_16182);
and U16399 (N_16399,N_16032,N_16155);
or U16400 (N_16400,N_16385,N_16340);
nor U16401 (N_16401,N_16223,N_16212);
nand U16402 (N_16402,N_16323,N_16315);
xnor U16403 (N_16403,N_16241,N_16394);
nor U16404 (N_16404,N_16344,N_16330);
and U16405 (N_16405,N_16220,N_16318);
and U16406 (N_16406,N_16316,N_16342);
or U16407 (N_16407,N_16262,N_16368);
and U16408 (N_16408,N_16303,N_16313);
and U16409 (N_16409,N_16392,N_16309);
nand U16410 (N_16410,N_16234,N_16387);
nor U16411 (N_16411,N_16213,N_16382);
nand U16412 (N_16412,N_16383,N_16235);
and U16413 (N_16413,N_16364,N_16254);
xnor U16414 (N_16414,N_16244,N_16377);
nor U16415 (N_16415,N_16358,N_16356);
xor U16416 (N_16416,N_16210,N_16232);
or U16417 (N_16417,N_16355,N_16304);
and U16418 (N_16418,N_16273,N_16258);
nand U16419 (N_16419,N_16259,N_16384);
or U16420 (N_16420,N_16204,N_16291);
xor U16421 (N_16421,N_16221,N_16239);
and U16422 (N_16422,N_16278,N_16395);
xnor U16423 (N_16423,N_16374,N_16307);
or U16424 (N_16424,N_16317,N_16231);
nor U16425 (N_16425,N_16396,N_16361);
or U16426 (N_16426,N_16376,N_16202);
nand U16427 (N_16427,N_16351,N_16287);
or U16428 (N_16428,N_16240,N_16299);
or U16429 (N_16429,N_16208,N_16345);
nand U16430 (N_16430,N_16333,N_16267);
or U16431 (N_16431,N_16238,N_16276);
nand U16432 (N_16432,N_16371,N_16296);
and U16433 (N_16433,N_16378,N_16386);
and U16434 (N_16434,N_16380,N_16292);
nand U16435 (N_16435,N_16373,N_16263);
or U16436 (N_16436,N_16247,N_16227);
nor U16437 (N_16437,N_16335,N_16275);
and U16438 (N_16438,N_16334,N_16290);
nand U16439 (N_16439,N_16367,N_16203);
and U16440 (N_16440,N_16269,N_16314);
nand U16441 (N_16441,N_16328,N_16214);
xnor U16442 (N_16442,N_16322,N_16260);
xnor U16443 (N_16443,N_16388,N_16349);
nor U16444 (N_16444,N_16312,N_16390);
xnor U16445 (N_16445,N_16230,N_16346);
nand U16446 (N_16446,N_16353,N_16337);
nand U16447 (N_16447,N_16256,N_16209);
nand U16448 (N_16448,N_16280,N_16372);
nor U16449 (N_16449,N_16215,N_16357);
nor U16450 (N_16450,N_16249,N_16348);
or U16451 (N_16451,N_16237,N_16326);
xnor U16452 (N_16452,N_16257,N_16288);
nor U16453 (N_16453,N_16206,N_16265);
nor U16454 (N_16454,N_16339,N_16228);
or U16455 (N_16455,N_16369,N_16381);
nand U16456 (N_16456,N_16294,N_16293);
nor U16457 (N_16457,N_16266,N_16325);
nand U16458 (N_16458,N_16284,N_16245);
nand U16459 (N_16459,N_16264,N_16305);
and U16460 (N_16460,N_16246,N_16200);
and U16461 (N_16461,N_16252,N_16338);
xnor U16462 (N_16462,N_16310,N_16391);
nand U16463 (N_16463,N_16352,N_16250);
xnor U16464 (N_16464,N_16217,N_16270);
and U16465 (N_16465,N_16242,N_16375);
xnor U16466 (N_16466,N_16393,N_16298);
or U16467 (N_16467,N_16389,N_16222);
nor U16468 (N_16468,N_16274,N_16282);
nand U16469 (N_16469,N_16216,N_16218);
or U16470 (N_16470,N_16201,N_16243);
or U16471 (N_16471,N_16336,N_16233);
or U16472 (N_16472,N_16253,N_16229);
nor U16473 (N_16473,N_16311,N_16224);
or U16474 (N_16474,N_16343,N_16236);
xor U16475 (N_16475,N_16272,N_16277);
xor U16476 (N_16476,N_16286,N_16205);
xnor U16477 (N_16477,N_16359,N_16306);
nand U16478 (N_16478,N_16363,N_16329);
nor U16479 (N_16479,N_16308,N_16324);
and U16480 (N_16480,N_16283,N_16321);
xor U16481 (N_16481,N_16319,N_16301);
nor U16482 (N_16482,N_16397,N_16360);
xor U16483 (N_16483,N_16289,N_16332);
xor U16484 (N_16484,N_16366,N_16248);
and U16485 (N_16485,N_16271,N_16297);
xnor U16486 (N_16486,N_16255,N_16261);
xnor U16487 (N_16487,N_16320,N_16226);
and U16488 (N_16488,N_16350,N_16398);
nor U16489 (N_16489,N_16341,N_16285);
nand U16490 (N_16490,N_16399,N_16362);
nor U16491 (N_16491,N_16370,N_16300);
and U16492 (N_16492,N_16219,N_16331);
or U16493 (N_16493,N_16268,N_16225);
xor U16494 (N_16494,N_16379,N_16347);
or U16495 (N_16495,N_16295,N_16281);
and U16496 (N_16496,N_16207,N_16354);
xor U16497 (N_16497,N_16365,N_16251);
or U16498 (N_16498,N_16279,N_16211);
and U16499 (N_16499,N_16327,N_16302);
xor U16500 (N_16500,N_16360,N_16372);
nand U16501 (N_16501,N_16232,N_16365);
and U16502 (N_16502,N_16372,N_16312);
or U16503 (N_16503,N_16261,N_16324);
and U16504 (N_16504,N_16264,N_16334);
or U16505 (N_16505,N_16287,N_16330);
nand U16506 (N_16506,N_16394,N_16266);
nor U16507 (N_16507,N_16208,N_16232);
nand U16508 (N_16508,N_16235,N_16355);
or U16509 (N_16509,N_16349,N_16226);
or U16510 (N_16510,N_16251,N_16294);
or U16511 (N_16511,N_16243,N_16222);
xnor U16512 (N_16512,N_16377,N_16207);
or U16513 (N_16513,N_16201,N_16240);
nand U16514 (N_16514,N_16352,N_16232);
nand U16515 (N_16515,N_16336,N_16215);
nand U16516 (N_16516,N_16322,N_16256);
nand U16517 (N_16517,N_16268,N_16315);
or U16518 (N_16518,N_16388,N_16367);
xnor U16519 (N_16519,N_16315,N_16361);
and U16520 (N_16520,N_16245,N_16398);
nand U16521 (N_16521,N_16352,N_16342);
or U16522 (N_16522,N_16228,N_16350);
and U16523 (N_16523,N_16314,N_16312);
nand U16524 (N_16524,N_16215,N_16217);
or U16525 (N_16525,N_16244,N_16331);
or U16526 (N_16526,N_16345,N_16232);
xor U16527 (N_16527,N_16397,N_16268);
nand U16528 (N_16528,N_16292,N_16308);
xnor U16529 (N_16529,N_16302,N_16231);
and U16530 (N_16530,N_16312,N_16248);
or U16531 (N_16531,N_16231,N_16344);
nand U16532 (N_16532,N_16389,N_16210);
nor U16533 (N_16533,N_16352,N_16212);
or U16534 (N_16534,N_16246,N_16277);
xor U16535 (N_16535,N_16323,N_16283);
nand U16536 (N_16536,N_16262,N_16253);
xnor U16537 (N_16537,N_16371,N_16301);
xor U16538 (N_16538,N_16344,N_16276);
or U16539 (N_16539,N_16290,N_16311);
xor U16540 (N_16540,N_16201,N_16217);
nor U16541 (N_16541,N_16355,N_16360);
nor U16542 (N_16542,N_16263,N_16300);
nand U16543 (N_16543,N_16212,N_16327);
or U16544 (N_16544,N_16349,N_16322);
or U16545 (N_16545,N_16340,N_16368);
nor U16546 (N_16546,N_16273,N_16279);
xor U16547 (N_16547,N_16346,N_16232);
and U16548 (N_16548,N_16340,N_16389);
nor U16549 (N_16549,N_16214,N_16207);
xor U16550 (N_16550,N_16217,N_16322);
nor U16551 (N_16551,N_16213,N_16340);
nor U16552 (N_16552,N_16394,N_16270);
nand U16553 (N_16553,N_16276,N_16207);
xnor U16554 (N_16554,N_16390,N_16248);
or U16555 (N_16555,N_16364,N_16233);
and U16556 (N_16556,N_16217,N_16210);
or U16557 (N_16557,N_16245,N_16291);
nor U16558 (N_16558,N_16250,N_16217);
or U16559 (N_16559,N_16300,N_16243);
and U16560 (N_16560,N_16268,N_16339);
or U16561 (N_16561,N_16235,N_16337);
nor U16562 (N_16562,N_16219,N_16266);
xnor U16563 (N_16563,N_16320,N_16250);
nand U16564 (N_16564,N_16342,N_16362);
nor U16565 (N_16565,N_16333,N_16389);
and U16566 (N_16566,N_16243,N_16258);
nor U16567 (N_16567,N_16328,N_16297);
or U16568 (N_16568,N_16316,N_16357);
nand U16569 (N_16569,N_16317,N_16222);
nand U16570 (N_16570,N_16232,N_16312);
nor U16571 (N_16571,N_16216,N_16283);
xnor U16572 (N_16572,N_16362,N_16229);
or U16573 (N_16573,N_16328,N_16236);
or U16574 (N_16574,N_16236,N_16304);
or U16575 (N_16575,N_16271,N_16386);
and U16576 (N_16576,N_16395,N_16389);
and U16577 (N_16577,N_16295,N_16244);
nand U16578 (N_16578,N_16385,N_16269);
nor U16579 (N_16579,N_16361,N_16389);
nor U16580 (N_16580,N_16282,N_16243);
or U16581 (N_16581,N_16382,N_16376);
nor U16582 (N_16582,N_16393,N_16207);
xnor U16583 (N_16583,N_16261,N_16246);
nand U16584 (N_16584,N_16325,N_16286);
and U16585 (N_16585,N_16341,N_16355);
xnor U16586 (N_16586,N_16320,N_16283);
and U16587 (N_16587,N_16227,N_16211);
nand U16588 (N_16588,N_16358,N_16216);
nor U16589 (N_16589,N_16227,N_16330);
nor U16590 (N_16590,N_16284,N_16288);
nor U16591 (N_16591,N_16348,N_16344);
nand U16592 (N_16592,N_16349,N_16291);
xnor U16593 (N_16593,N_16319,N_16388);
xor U16594 (N_16594,N_16349,N_16387);
nor U16595 (N_16595,N_16214,N_16259);
nand U16596 (N_16596,N_16318,N_16223);
and U16597 (N_16597,N_16267,N_16273);
or U16598 (N_16598,N_16306,N_16360);
nand U16599 (N_16599,N_16304,N_16249);
and U16600 (N_16600,N_16513,N_16527);
and U16601 (N_16601,N_16533,N_16423);
and U16602 (N_16602,N_16484,N_16406);
and U16603 (N_16603,N_16520,N_16471);
nand U16604 (N_16604,N_16461,N_16591);
xor U16605 (N_16605,N_16452,N_16540);
or U16606 (N_16606,N_16595,N_16511);
nor U16607 (N_16607,N_16524,N_16496);
nor U16608 (N_16608,N_16556,N_16531);
nand U16609 (N_16609,N_16573,N_16514);
or U16610 (N_16610,N_16586,N_16404);
and U16611 (N_16611,N_16434,N_16537);
and U16612 (N_16612,N_16432,N_16580);
nand U16613 (N_16613,N_16592,N_16410);
xnor U16614 (N_16614,N_16541,N_16491);
and U16615 (N_16615,N_16439,N_16467);
xnor U16616 (N_16616,N_16532,N_16530);
nand U16617 (N_16617,N_16510,N_16574);
nor U16618 (N_16618,N_16475,N_16553);
nand U16619 (N_16619,N_16430,N_16518);
and U16620 (N_16620,N_16577,N_16494);
xnor U16621 (N_16621,N_16435,N_16441);
nand U16622 (N_16622,N_16589,N_16488);
or U16623 (N_16623,N_16419,N_16442);
and U16624 (N_16624,N_16490,N_16481);
nand U16625 (N_16625,N_16584,N_16468);
xnor U16626 (N_16626,N_16413,N_16493);
or U16627 (N_16627,N_16550,N_16457);
nand U16628 (N_16628,N_16585,N_16528);
xnor U16629 (N_16629,N_16500,N_16409);
or U16630 (N_16630,N_16499,N_16521);
nand U16631 (N_16631,N_16454,N_16509);
or U16632 (N_16632,N_16558,N_16599);
nor U16633 (N_16633,N_16502,N_16534);
xor U16634 (N_16634,N_16400,N_16578);
or U16635 (N_16635,N_16497,N_16549);
nand U16636 (N_16636,N_16464,N_16562);
nor U16637 (N_16637,N_16449,N_16412);
nand U16638 (N_16638,N_16460,N_16548);
nor U16639 (N_16639,N_16477,N_16448);
or U16640 (N_16640,N_16505,N_16582);
or U16641 (N_16641,N_16424,N_16428);
and U16642 (N_16642,N_16416,N_16450);
nor U16643 (N_16643,N_16529,N_16451);
and U16644 (N_16644,N_16403,N_16411);
nor U16645 (N_16645,N_16455,N_16443);
or U16646 (N_16646,N_16517,N_16405);
xnor U16647 (N_16647,N_16446,N_16485);
or U16648 (N_16648,N_16576,N_16427);
and U16649 (N_16649,N_16483,N_16401);
or U16650 (N_16650,N_16426,N_16551);
xor U16651 (N_16651,N_16503,N_16445);
and U16652 (N_16652,N_16482,N_16526);
or U16653 (N_16653,N_16561,N_16469);
nor U16654 (N_16654,N_16414,N_16437);
nand U16655 (N_16655,N_16564,N_16453);
and U16656 (N_16656,N_16438,N_16570);
and U16657 (N_16657,N_16594,N_16572);
nand U16658 (N_16658,N_16512,N_16458);
or U16659 (N_16659,N_16474,N_16407);
xnor U16660 (N_16660,N_16408,N_16587);
xnor U16661 (N_16661,N_16543,N_16568);
nor U16662 (N_16662,N_16523,N_16590);
xnor U16663 (N_16663,N_16478,N_16486);
and U16664 (N_16664,N_16569,N_16422);
xnor U16665 (N_16665,N_16504,N_16487);
or U16666 (N_16666,N_16421,N_16588);
nand U16667 (N_16667,N_16547,N_16579);
nand U16668 (N_16668,N_16420,N_16470);
nor U16669 (N_16669,N_16473,N_16557);
xnor U16670 (N_16670,N_16535,N_16536);
and U16671 (N_16671,N_16480,N_16417);
xor U16672 (N_16672,N_16593,N_16555);
nand U16673 (N_16673,N_16567,N_16440);
nand U16674 (N_16674,N_16539,N_16542);
nand U16675 (N_16675,N_16566,N_16538);
or U16676 (N_16676,N_16456,N_16465);
xor U16677 (N_16677,N_16516,N_16463);
nand U16678 (N_16678,N_16402,N_16563);
nand U16679 (N_16679,N_16546,N_16476);
nand U16680 (N_16680,N_16519,N_16431);
or U16681 (N_16681,N_16506,N_16522);
or U16682 (N_16682,N_16495,N_16581);
and U16683 (N_16683,N_16525,N_16507);
or U16684 (N_16684,N_16429,N_16508);
or U16685 (N_16685,N_16571,N_16575);
nand U16686 (N_16686,N_16444,N_16425);
xnor U16687 (N_16687,N_16436,N_16565);
nand U16688 (N_16688,N_16559,N_16466);
xor U16689 (N_16689,N_16447,N_16498);
xnor U16690 (N_16690,N_16462,N_16560);
xor U16691 (N_16691,N_16598,N_16492);
xor U16692 (N_16692,N_16597,N_16472);
xnor U16693 (N_16693,N_16552,N_16583);
and U16694 (N_16694,N_16501,N_16459);
nor U16695 (N_16695,N_16489,N_16418);
nor U16696 (N_16696,N_16433,N_16545);
or U16697 (N_16697,N_16544,N_16479);
and U16698 (N_16698,N_16415,N_16554);
or U16699 (N_16699,N_16515,N_16596);
or U16700 (N_16700,N_16450,N_16400);
xnor U16701 (N_16701,N_16410,N_16416);
nand U16702 (N_16702,N_16568,N_16566);
nor U16703 (N_16703,N_16563,N_16595);
nand U16704 (N_16704,N_16439,N_16481);
nor U16705 (N_16705,N_16404,N_16499);
or U16706 (N_16706,N_16524,N_16551);
or U16707 (N_16707,N_16564,N_16401);
or U16708 (N_16708,N_16415,N_16426);
or U16709 (N_16709,N_16403,N_16460);
nand U16710 (N_16710,N_16598,N_16478);
nand U16711 (N_16711,N_16520,N_16405);
nand U16712 (N_16712,N_16514,N_16443);
or U16713 (N_16713,N_16579,N_16450);
nor U16714 (N_16714,N_16460,N_16416);
xnor U16715 (N_16715,N_16526,N_16510);
xor U16716 (N_16716,N_16444,N_16489);
and U16717 (N_16717,N_16553,N_16570);
xor U16718 (N_16718,N_16500,N_16424);
nor U16719 (N_16719,N_16502,N_16420);
or U16720 (N_16720,N_16551,N_16574);
or U16721 (N_16721,N_16472,N_16454);
and U16722 (N_16722,N_16560,N_16484);
xor U16723 (N_16723,N_16528,N_16447);
or U16724 (N_16724,N_16485,N_16566);
or U16725 (N_16725,N_16439,N_16513);
or U16726 (N_16726,N_16532,N_16504);
nand U16727 (N_16727,N_16548,N_16552);
or U16728 (N_16728,N_16424,N_16412);
or U16729 (N_16729,N_16457,N_16488);
nor U16730 (N_16730,N_16482,N_16564);
xor U16731 (N_16731,N_16596,N_16512);
and U16732 (N_16732,N_16442,N_16421);
nor U16733 (N_16733,N_16492,N_16534);
xnor U16734 (N_16734,N_16504,N_16412);
nor U16735 (N_16735,N_16440,N_16501);
nor U16736 (N_16736,N_16538,N_16492);
nand U16737 (N_16737,N_16430,N_16542);
and U16738 (N_16738,N_16403,N_16510);
nand U16739 (N_16739,N_16408,N_16493);
and U16740 (N_16740,N_16431,N_16595);
or U16741 (N_16741,N_16586,N_16595);
or U16742 (N_16742,N_16403,N_16487);
nor U16743 (N_16743,N_16488,N_16422);
and U16744 (N_16744,N_16513,N_16414);
xnor U16745 (N_16745,N_16523,N_16466);
nand U16746 (N_16746,N_16453,N_16442);
nand U16747 (N_16747,N_16433,N_16520);
xnor U16748 (N_16748,N_16542,N_16488);
nand U16749 (N_16749,N_16493,N_16576);
nor U16750 (N_16750,N_16590,N_16447);
or U16751 (N_16751,N_16538,N_16424);
nand U16752 (N_16752,N_16509,N_16568);
nand U16753 (N_16753,N_16597,N_16402);
nor U16754 (N_16754,N_16439,N_16441);
and U16755 (N_16755,N_16503,N_16579);
nand U16756 (N_16756,N_16465,N_16471);
nor U16757 (N_16757,N_16404,N_16508);
and U16758 (N_16758,N_16430,N_16428);
or U16759 (N_16759,N_16582,N_16476);
xnor U16760 (N_16760,N_16578,N_16531);
xor U16761 (N_16761,N_16465,N_16526);
nand U16762 (N_16762,N_16599,N_16455);
or U16763 (N_16763,N_16531,N_16530);
nand U16764 (N_16764,N_16488,N_16576);
or U16765 (N_16765,N_16564,N_16572);
and U16766 (N_16766,N_16413,N_16587);
nand U16767 (N_16767,N_16528,N_16571);
and U16768 (N_16768,N_16597,N_16434);
or U16769 (N_16769,N_16521,N_16462);
or U16770 (N_16770,N_16527,N_16508);
and U16771 (N_16771,N_16472,N_16569);
nand U16772 (N_16772,N_16503,N_16440);
nand U16773 (N_16773,N_16432,N_16467);
nand U16774 (N_16774,N_16505,N_16476);
or U16775 (N_16775,N_16460,N_16573);
or U16776 (N_16776,N_16590,N_16531);
nor U16777 (N_16777,N_16505,N_16532);
xnor U16778 (N_16778,N_16512,N_16555);
nand U16779 (N_16779,N_16488,N_16448);
xor U16780 (N_16780,N_16448,N_16466);
or U16781 (N_16781,N_16420,N_16568);
and U16782 (N_16782,N_16576,N_16405);
or U16783 (N_16783,N_16534,N_16453);
nand U16784 (N_16784,N_16556,N_16553);
and U16785 (N_16785,N_16596,N_16594);
or U16786 (N_16786,N_16531,N_16445);
or U16787 (N_16787,N_16506,N_16491);
xor U16788 (N_16788,N_16443,N_16451);
xnor U16789 (N_16789,N_16551,N_16582);
nand U16790 (N_16790,N_16491,N_16562);
xor U16791 (N_16791,N_16554,N_16491);
xnor U16792 (N_16792,N_16435,N_16514);
nand U16793 (N_16793,N_16577,N_16476);
nor U16794 (N_16794,N_16474,N_16487);
nand U16795 (N_16795,N_16570,N_16492);
nand U16796 (N_16796,N_16436,N_16555);
nand U16797 (N_16797,N_16532,N_16551);
or U16798 (N_16798,N_16537,N_16500);
and U16799 (N_16799,N_16465,N_16583);
xor U16800 (N_16800,N_16624,N_16617);
xor U16801 (N_16801,N_16752,N_16608);
or U16802 (N_16802,N_16674,N_16686);
or U16803 (N_16803,N_16771,N_16706);
and U16804 (N_16804,N_16613,N_16737);
and U16805 (N_16805,N_16754,N_16796);
or U16806 (N_16806,N_16785,N_16725);
and U16807 (N_16807,N_16779,N_16755);
or U16808 (N_16808,N_16703,N_16670);
or U16809 (N_16809,N_16695,N_16681);
nor U16810 (N_16810,N_16627,N_16764);
or U16811 (N_16811,N_16615,N_16741);
and U16812 (N_16812,N_16788,N_16778);
nor U16813 (N_16813,N_16738,N_16787);
xor U16814 (N_16814,N_16731,N_16626);
nor U16815 (N_16815,N_16665,N_16746);
and U16816 (N_16816,N_16740,N_16723);
or U16817 (N_16817,N_16638,N_16628);
nor U16818 (N_16818,N_16791,N_16707);
xnor U16819 (N_16819,N_16636,N_16605);
nor U16820 (N_16820,N_16654,N_16770);
nor U16821 (N_16821,N_16767,N_16679);
or U16822 (N_16822,N_16689,N_16742);
and U16823 (N_16823,N_16783,N_16781);
or U16824 (N_16824,N_16601,N_16727);
nor U16825 (N_16825,N_16696,N_16712);
nor U16826 (N_16826,N_16774,N_16612);
xor U16827 (N_16827,N_16729,N_16691);
and U16828 (N_16828,N_16747,N_16682);
nand U16829 (N_16829,N_16693,N_16713);
nor U16830 (N_16830,N_16611,N_16652);
and U16831 (N_16831,N_16776,N_16694);
nor U16832 (N_16832,N_16784,N_16661);
and U16833 (N_16833,N_16623,N_16633);
or U16834 (N_16834,N_16790,N_16655);
or U16835 (N_16835,N_16692,N_16683);
xnor U16836 (N_16836,N_16688,N_16606);
nand U16837 (N_16837,N_16717,N_16647);
xnor U16838 (N_16838,N_16650,N_16625);
nor U16839 (N_16839,N_16739,N_16634);
and U16840 (N_16840,N_16632,N_16722);
nor U16841 (N_16841,N_16765,N_16672);
or U16842 (N_16842,N_16761,N_16648);
nand U16843 (N_16843,N_16732,N_16645);
nor U16844 (N_16844,N_16667,N_16622);
and U16845 (N_16845,N_16714,N_16753);
or U16846 (N_16846,N_16642,N_16720);
and U16847 (N_16847,N_16794,N_16759);
nand U16848 (N_16848,N_16637,N_16748);
nand U16849 (N_16849,N_16724,N_16671);
xor U16850 (N_16850,N_16676,N_16718);
nand U16851 (N_16851,N_16610,N_16660);
xor U16852 (N_16852,N_16620,N_16616);
and U16853 (N_16853,N_16659,N_16710);
xnor U16854 (N_16854,N_16609,N_16697);
nand U16855 (N_16855,N_16704,N_16711);
and U16856 (N_16856,N_16773,N_16603);
or U16857 (N_16857,N_16777,N_16619);
nor U16858 (N_16858,N_16736,N_16685);
and U16859 (N_16859,N_16658,N_16769);
xnor U16860 (N_16860,N_16621,N_16749);
or U16861 (N_16861,N_16709,N_16675);
and U16862 (N_16862,N_16678,N_16656);
and U16863 (N_16863,N_16630,N_16662);
xor U16864 (N_16864,N_16690,N_16700);
xor U16865 (N_16865,N_16699,N_16677);
nor U16866 (N_16866,N_16701,N_16649);
and U16867 (N_16867,N_16789,N_16756);
nand U16868 (N_16868,N_16726,N_16733);
nand U16869 (N_16869,N_16663,N_16772);
nor U16870 (N_16870,N_16762,N_16716);
xnor U16871 (N_16871,N_16763,N_16728);
nand U16872 (N_16872,N_16640,N_16607);
nor U16873 (N_16873,N_16786,N_16684);
and U16874 (N_16874,N_16639,N_16646);
nand U16875 (N_16875,N_16730,N_16631);
and U16876 (N_16876,N_16687,N_16600);
nor U16877 (N_16877,N_16744,N_16780);
nand U16878 (N_16878,N_16618,N_16664);
nor U16879 (N_16879,N_16766,N_16602);
nand U16880 (N_16880,N_16799,N_16702);
nor U16881 (N_16881,N_16629,N_16768);
nor U16882 (N_16882,N_16669,N_16792);
nor U16883 (N_16883,N_16604,N_16721);
and U16884 (N_16884,N_16719,N_16644);
xnor U16885 (N_16885,N_16651,N_16643);
and U16886 (N_16886,N_16798,N_16680);
xnor U16887 (N_16887,N_16657,N_16797);
nor U16888 (N_16888,N_16734,N_16614);
nor U16889 (N_16889,N_16743,N_16760);
and U16890 (N_16890,N_16795,N_16757);
xnor U16891 (N_16891,N_16751,N_16698);
or U16892 (N_16892,N_16775,N_16673);
or U16893 (N_16893,N_16641,N_16735);
nand U16894 (N_16894,N_16793,N_16758);
or U16895 (N_16895,N_16708,N_16653);
nor U16896 (N_16896,N_16750,N_16715);
xnor U16897 (N_16897,N_16745,N_16705);
nand U16898 (N_16898,N_16668,N_16782);
and U16899 (N_16899,N_16635,N_16666);
nor U16900 (N_16900,N_16622,N_16729);
xnor U16901 (N_16901,N_16632,N_16702);
nor U16902 (N_16902,N_16642,N_16739);
and U16903 (N_16903,N_16679,N_16758);
nand U16904 (N_16904,N_16621,N_16715);
and U16905 (N_16905,N_16727,N_16690);
nor U16906 (N_16906,N_16671,N_16613);
and U16907 (N_16907,N_16793,N_16601);
and U16908 (N_16908,N_16728,N_16700);
nand U16909 (N_16909,N_16607,N_16719);
or U16910 (N_16910,N_16764,N_16671);
nand U16911 (N_16911,N_16762,N_16637);
and U16912 (N_16912,N_16609,N_16699);
nor U16913 (N_16913,N_16763,N_16796);
xnor U16914 (N_16914,N_16755,N_16664);
or U16915 (N_16915,N_16794,N_16782);
nor U16916 (N_16916,N_16626,N_16744);
or U16917 (N_16917,N_16732,N_16733);
xor U16918 (N_16918,N_16688,N_16746);
xnor U16919 (N_16919,N_16760,N_16709);
or U16920 (N_16920,N_16614,N_16735);
or U16921 (N_16921,N_16617,N_16661);
nand U16922 (N_16922,N_16759,N_16797);
and U16923 (N_16923,N_16778,N_16628);
xor U16924 (N_16924,N_16614,N_16791);
nand U16925 (N_16925,N_16760,N_16651);
nor U16926 (N_16926,N_16708,N_16630);
nand U16927 (N_16927,N_16648,N_16673);
or U16928 (N_16928,N_16671,N_16615);
nor U16929 (N_16929,N_16759,N_16677);
xnor U16930 (N_16930,N_16613,N_16604);
or U16931 (N_16931,N_16673,N_16674);
nor U16932 (N_16932,N_16689,N_16782);
nand U16933 (N_16933,N_16782,N_16673);
nor U16934 (N_16934,N_16690,N_16651);
nor U16935 (N_16935,N_16728,N_16786);
or U16936 (N_16936,N_16699,N_16701);
nor U16937 (N_16937,N_16766,N_16786);
xor U16938 (N_16938,N_16752,N_16756);
or U16939 (N_16939,N_16717,N_16691);
nor U16940 (N_16940,N_16639,N_16657);
and U16941 (N_16941,N_16790,N_16601);
and U16942 (N_16942,N_16771,N_16662);
and U16943 (N_16943,N_16749,N_16620);
and U16944 (N_16944,N_16718,N_16648);
and U16945 (N_16945,N_16740,N_16691);
nor U16946 (N_16946,N_16696,N_16676);
xor U16947 (N_16947,N_16725,N_16730);
nand U16948 (N_16948,N_16688,N_16605);
nor U16949 (N_16949,N_16682,N_16660);
nor U16950 (N_16950,N_16758,N_16694);
and U16951 (N_16951,N_16775,N_16658);
and U16952 (N_16952,N_16756,N_16760);
nor U16953 (N_16953,N_16716,N_16697);
nand U16954 (N_16954,N_16652,N_16644);
and U16955 (N_16955,N_16728,N_16790);
and U16956 (N_16956,N_16663,N_16755);
xnor U16957 (N_16957,N_16756,N_16639);
nor U16958 (N_16958,N_16600,N_16638);
nor U16959 (N_16959,N_16660,N_16665);
or U16960 (N_16960,N_16709,N_16716);
or U16961 (N_16961,N_16681,N_16720);
xnor U16962 (N_16962,N_16669,N_16642);
xnor U16963 (N_16963,N_16707,N_16642);
xor U16964 (N_16964,N_16676,N_16615);
xnor U16965 (N_16965,N_16620,N_16768);
nand U16966 (N_16966,N_16792,N_16684);
or U16967 (N_16967,N_16735,N_16682);
xor U16968 (N_16968,N_16680,N_16671);
xnor U16969 (N_16969,N_16616,N_16686);
and U16970 (N_16970,N_16770,N_16641);
and U16971 (N_16971,N_16648,N_16757);
nand U16972 (N_16972,N_16649,N_16641);
xnor U16973 (N_16973,N_16681,N_16791);
xor U16974 (N_16974,N_16733,N_16735);
or U16975 (N_16975,N_16636,N_16731);
or U16976 (N_16976,N_16603,N_16700);
xor U16977 (N_16977,N_16750,N_16720);
xor U16978 (N_16978,N_16722,N_16747);
or U16979 (N_16979,N_16727,N_16703);
xor U16980 (N_16980,N_16713,N_16780);
nor U16981 (N_16981,N_16677,N_16667);
or U16982 (N_16982,N_16626,N_16693);
nand U16983 (N_16983,N_16732,N_16644);
nor U16984 (N_16984,N_16650,N_16657);
xnor U16985 (N_16985,N_16700,N_16715);
xnor U16986 (N_16986,N_16724,N_16755);
or U16987 (N_16987,N_16719,N_16614);
nor U16988 (N_16988,N_16770,N_16622);
nor U16989 (N_16989,N_16652,N_16635);
nor U16990 (N_16990,N_16636,N_16635);
nor U16991 (N_16991,N_16661,N_16603);
nand U16992 (N_16992,N_16653,N_16737);
or U16993 (N_16993,N_16677,N_16727);
and U16994 (N_16994,N_16661,N_16778);
xor U16995 (N_16995,N_16742,N_16638);
or U16996 (N_16996,N_16655,N_16645);
nor U16997 (N_16997,N_16717,N_16779);
xnor U16998 (N_16998,N_16681,N_16723);
or U16999 (N_16999,N_16693,N_16657);
nor U17000 (N_17000,N_16977,N_16946);
nand U17001 (N_17001,N_16989,N_16881);
nand U17002 (N_17002,N_16948,N_16910);
nor U17003 (N_17003,N_16897,N_16916);
and U17004 (N_17004,N_16814,N_16918);
xor U17005 (N_17005,N_16995,N_16834);
xor U17006 (N_17006,N_16923,N_16963);
nor U17007 (N_17007,N_16965,N_16932);
nand U17008 (N_17008,N_16981,N_16927);
nand U17009 (N_17009,N_16872,N_16951);
or U17010 (N_17010,N_16847,N_16828);
nor U17011 (N_17011,N_16898,N_16821);
or U17012 (N_17012,N_16856,N_16836);
nor U17013 (N_17013,N_16956,N_16998);
nand U17014 (N_17014,N_16970,N_16954);
nor U17015 (N_17015,N_16808,N_16961);
nand U17016 (N_17016,N_16876,N_16925);
xor U17017 (N_17017,N_16894,N_16815);
nor U17018 (N_17018,N_16824,N_16907);
or U17019 (N_17019,N_16978,N_16988);
and U17020 (N_17020,N_16950,N_16822);
nor U17021 (N_17021,N_16972,N_16975);
and U17022 (N_17022,N_16813,N_16952);
or U17023 (N_17023,N_16871,N_16841);
xnor U17024 (N_17024,N_16949,N_16940);
nand U17025 (N_17025,N_16987,N_16895);
or U17026 (N_17026,N_16866,N_16921);
and U17027 (N_17027,N_16826,N_16979);
and U17028 (N_17028,N_16830,N_16874);
xor U17029 (N_17029,N_16846,N_16984);
nand U17030 (N_17030,N_16880,N_16862);
xor U17031 (N_17031,N_16868,N_16971);
nand U17032 (N_17032,N_16980,N_16967);
xor U17033 (N_17033,N_16937,N_16805);
nor U17034 (N_17034,N_16867,N_16829);
or U17035 (N_17035,N_16986,N_16827);
or U17036 (N_17036,N_16966,N_16982);
and U17037 (N_17037,N_16877,N_16840);
xor U17038 (N_17038,N_16990,N_16920);
and U17039 (N_17039,N_16800,N_16863);
and U17040 (N_17040,N_16914,N_16983);
nand U17041 (N_17041,N_16930,N_16857);
nand U17042 (N_17042,N_16869,N_16945);
xnor U17043 (N_17043,N_16806,N_16942);
or U17044 (N_17044,N_16964,N_16913);
nand U17045 (N_17045,N_16818,N_16935);
and U17046 (N_17046,N_16973,N_16976);
or U17047 (N_17047,N_16844,N_16999);
nor U17048 (N_17048,N_16802,N_16934);
nand U17049 (N_17049,N_16892,N_16994);
or U17050 (N_17050,N_16947,N_16843);
xnor U17051 (N_17051,N_16996,N_16922);
xor U17052 (N_17052,N_16997,N_16875);
nor U17053 (N_17053,N_16837,N_16931);
nand U17054 (N_17054,N_16850,N_16820);
nor U17055 (N_17055,N_16833,N_16929);
nor U17056 (N_17056,N_16804,N_16953);
or U17057 (N_17057,N_16991,N_16845);
or U17058 (N_17058,N_16878,N_16839);
nand U17059 (N_17059,N_16855,N_16993);
or U17060 (N_17060,N_16882,N_16889);
nand U17061 (N_17061,N_16823,N_16865);
nor U17062 (N_17062,N_16886,N_16899);
nand U17063 (N_17063,N_16807,N_16870);
or U17064 (N_17064,N_16851,N_16810);
xnor U17065 (N_17065,N_16879,N_16884);
and U17066 (N_17066,N_16819,N_16904);
xnor U17067 (N_17067,N_16854,N_16917);
or U17068 (N_17068,N_16803,N_16957);
and U17069 (N_17069,N_16933,N_16812);
or U17070 (N_17070,N_16883,N_16816);
and U17071 (N_17071,N_16974,N_16939);
nand U17072 (N_17072,N_16900,N_16958);
or U17073 (N_17073,N_16873,N_16908);
nand U17074 (N_17074,N_16853,N_16891);
or U17075 (N_17075,N_16938,N_16968);
or U17076 (N_17076,N_16928,N_16825);
and U17077 (N_17077,N_16905,N_16912);
xor U17078 (N_17078,N_16944,N_16861);
nand U17079 (N_17079,N_16848,N_16852);
or U17080 (N_17080,N_16943,N_16864);
and U17081 (N_17081,N_16887,N_16842);
and U17082 (N_17082,N_16962,N_16911);
xor U17083 (N_17083,N_16960,N_16902);
and U17084 (N_17084,N_16924,N_16941);
nand U17085 (N_17085,N_16858,N_16909);
and U17086 (N_17086,N_16896,N_16890);
or U17087 (N_17087,N_16901,N_16969);
xnor U17088 (N_17088,N_16888,N_16801);
xor U17089 (N_17089,N_16832,N_16985);
nand U17090 (N_17090,N_16860,N_16811);
or U17091 (N_17091,N_16926,N_16915);
nand U17092 (N_17092,N_16906,N_16903);
and U17093 (N_17093,N_16936,N_16831);
xnor U17094 (N_17094,N_16885,N_16838);
nor U17095 (N_17095,N_16893,N_16955);
xnor U17096 (N_17096,N_16817,N_16959);
nor U17097 (N_17097,N_16809,N_16919);
and U17098 (N_17098,N_16859,N_16835);
nor U17099 (N_17099,N_16849,N_16992);
and U17100 (N_17100,N_16871,N_16914);
nor U17101 (N_17101,N_16968,N_16900);
or U17102 (N_17102,N_16969,N_16908);
nand U17103 (N_17103,N_16964,N_16977);
or U17104 (N_17104,N_16993,N_16851);
nand U17105 (N_17105,N_16888,N_16944);
or U17106 (N_17106,N_16806,N_16877);
xnor U17107 (N_17107,N_16964,N_16811);
nand U17108 (N_17108,N_16824,N_16963);
or U17109 (N_17109,N_16866,N_16860);
nand U17110 (N_17110,N_16929,N_16838);
nand U17111 (N_17111,N_16928,N_16986);
nor U17112 (N_17112,N_16976,N_16932);
nor U17113 (N_17113,N_16936,N_16854);
nor U17114 (N_17114,N_16805,N_16946);
nand U17115 (N_17115,N_16941,N_16931);
and U17116 (N_17116,N_16839,N_16964);
or U17117 (N_17117,N_16997,N_16969);
nor U17118 (N_17118,N_16997,N_16858);
or U17119 (N_17119,N_16927,N_16921);
or U17120 (N_17120,N_16816,N_16829);
or U17121 (N_17121,N_16954,N_16805);
xor U17122 (N_17122,N_16989,N_16903);
nand U17123 (N_17123,N_16850,N_16925);
nand U17124 (N_17124,N_16884,N_16962);
nor U17125 (N_17125,N_16825,N_16813);
nor U17126 (N_17126,N_16980,N_16837);
xor U17127 (N_17127,N_16978,N_16834);
or U17128 (N_17128,N_16981,N_16906);
nor U17129 (N_17129,N_16868,N_16815);
xor U17130 (N_17130,N_16868,N_16899);
or U17131 (N_17131,N_16914,N_16912);
or U17132 (N_17132,N_16868,N_16923);
or U17133 (N_17133,N_16899,N_16854);
and U17134 (N_17134,N_16962,N_16890);
xor U17135 (N_17135,N_16849,N_16907);
nor U17136 (N_17136,N_16936,N_16988);
nor U17137 (N_17137,N_16986,N_16926);
or U17138 (N_17138,N_16818,N_16841);
nand U17139 (N_17139,N_16998,N_16879);
xnor U17140 (N_17140,N_16832,N_16921);
xnor U17141 (N_17141,N_16947,N_16837);
or U17142 (N_17142,N_16999,N_16882);
and U17143 (N_17143,N_16982,N_16932);
and U17144 (N_17144,N_16814,N_16981);
and U17145 (N_17145,N_16965,N_16949);
and U17146 (N_17146,N_16898,N_16808);
or U17147 (N_17147,N_16996,N_16820);
and U17148 (N_17148,N_16966,N_16962);
nor U17149 (N_17149,N_16936,N_16940);
nand U17150 (N_17150,N_16828,N_16865);
and U17151 (N_17151,N_16949,N_16867);
nand U17152 (N_17152,N_16872,N_16918);
xor U17153 (N_17153,N_16848,N_16808);
nor U17154 (N_17154,N_16803,N_16989);
nor U17155 (N_17155,N_16856,N_16999);
and U17156 (N_17156,N_16868,N_16918);
xor U17157 (N_17157,N_16978,N_16997);
and U17158 (N_17158,N_16857,N_16990);
and U17159 (N_17159,N_16957,N_16980);
xnor U17160 (N_17160,N_16852,N_16975);
nand U17161 (N_17161,N_16835,N_16871);
and U17162 (N_17162,N_16836,N_16845);
and U17163 (N_17163,N_16980,N_16970);
xor U17164 (N_17164,N_16987,N_16904);
xnor U17165 (N_17165,N_16983,N_16944);
and U17166 (N_17166,N_16913,N_16860);
and U17167 (N_17167,N_16900,N_16902);
nor U17168 (N_17168,N_16836,N_16860);
xnor U17169 (N_17169,N_16860,N_16957);
nor U17170 (N_17170,N_16815,N_16883);
nor U17171 (N_17171,N_16953,N_16969);
nand U17172 (N_17172,N_16970,N_16914);
nand U17173 (N_17173,N_16961,N_16874);
nor U17174 (N_17174,N_16868,N_16843);
or U17175 (N_17175,N_16828,N_16971);
nor U17176 (N_17176,N_16879,N_16932);
nand U17177 (N_17177,N_16840,N_16991);
and U17178 (N_17178,N_16916,N_16865);
nand U17179 (N_17179,N_16830,N_16922);
xor U17180 (N_17180,N_16888,N_16925);
nand U17181 (N_17181,N_16920,N_16815);
nor U17182 (N_17182,N_16951,N_16892);
and U17183 (N_17183,N_16832,N_16882);
nor U17184 (N_17184,N_16906,N_16982);
and U17185 (N_17185,N_16848,N_16979);
nand U17186 (N_17186,N_16851,N_16955);
xnor U17187 (N_17187,N_16869,N_16895);
nand U17188 (N_17188,N_16877,N_16815);
xor U17189 (N_17189,N_16814,N_16801);
nand U17190 (N_17190,N_16830,N_16950);
or U17191 (N_17191,N_16989,N_16857);
nor U17192 (N_17192,N_16919,N_16945);
or U17193 (N_17193,N_16875,N_16820);
nand U17194 (N_17194,N_16815,N_16802);
xnor U17195 (N_17195,N_16926,N_16907);
nand U17196 (N_17196,N_16856,N_16899);
and U17197 (N_17197,N_16994,N_16938);
nor U17198 (N_17198,N_16936,N_16968);
or U17199 (N_17199,N_16939,N_16932);
xnor U17200 (N_17200,N_17002,N_17126);
and U17201 (N_17201,N_17017,N_17169);
nor U17202 (N_17202,N_17096,N_17048);
and U17203 (N_17203,N_17092,N_17052);
and U17204 (N_17204,N_17152,N_17187);
or U17205 (N_17205,N_17134,N_17004);
or U17206 (N_17206,N_17069,N_17108);
nand U17207 (N_17207,N_17089,N_17135);
and U17208 (N_17208,N_17129,N_17064);
nand U17209 (N_17209,N_17119,N_17006);
xor U17210 (N_17210,N_17102,N_17094);
nand U17211 (N_17211,N_17074,N_17142);
nor U17212 (N_17212,N_17084,N_17173);
or U17213 (N_17213,N_17055,N_17078);
xnor U17214 (N_17214,N_17071,N_17025);
and U17215 (N_17215,N_17112,N_17062);
and U17216 (N_17216,N_17113,N_17167);
xor U17217 (N_17217,N_17032,N_17028);
and U17218 (N_17218,N_17198,N_17177);
xor U17219 (N_17219,N_17000,N_17082);
or U17220 (N_17220,N_17022,N_17007);
and U17221 (N_17221,N_17088,N_17059);
and U17222 (N_17222,N_17040,N_17015);
and U17223 (N_17223,N_17166,N_17107);
and U17224 (N_17224,N_17189,N_17099);
nor U17225 (N_17225,N_17023,N_17097);
and U17226 (N_17226,N_17011,N_17106);
xnor U17227 (N_17227,N_17033,N_17144);
nand U17228 (N_17228,N_17045,N_17020);
nand U17229 (N_17229,N_17054,N_17125);
and U17230 (N_17230,N_17132,N_17013);
and U17231 (N_17231,N_17061,N_17160);
nor U17232 (N_17232,N_17080,N_17186);
nand U17233 (N_17233,N_17039,N_17188);
or U17234 (N_17234,N_17073,N_17058);
or U17235 (N_17235,N_17197,N_17154);
nand U17236 (N_17236,N_17195,N_17037);
xor U17237 (N_17237,N_17176,N_17036);
and U17238 (N_17238,N_17184,N_17153);
or U17239 (N_17239,N_17170,N_17087);
xnor U17240 (N_17240,N_17041,N_17035);
and U17241 (N_17241,N_17118,N_17063);
nand U17242 (N_17242,N_17042,N_17016);
and U17243 (N_17243,N_17044,N_17149);
or U17244 (N_17244,N_17162,N_17192);
and U17245 (N_17245,N_17180,N_17171);
or U17246 (N_17246,N_17021,N_17026);
nand U17247 (N_17247,N_17090,N_17191);
xnor U17248 (N_17248,N_17070,N_17123);
xnor U17249 (N_17249,N_17141,N_17024);
nor U17250 (N_17250,N_17030,N_17057);
or U17251 (N_17251,N_17196,N_17001);
and U17252 (N_17252,N_17005,N_17120);
or U17253 (N_17253,N_17109,N_17116);
xor U17254 (N_17254,N_17143,N_17105);
or U17255 (N_17255,N_17043,N_17068);
nand U17256 (N_17256,N_17009,N_17185);
nor U17257 (N_17257,N_17179,N_17121);
or U17258 (N_17258,N_17066,N_17072);
nor U17259 (N_17259,N_17174,N_17077);
xnor U17260 (N_17260,N_17095,N_17193);
nand U17261 (N_17261,N_17182,N_17128);
xnor U17262 (N_17262,N_17172,N_17130);
and U17263 (N_17263,N_17161,N_17155);
and U17264 (N_17264,N_17150,N_17098);
or U17265 (N_17265,N_17085,N_17104);
nand U17266 (N_17266,N_17183,N_17147);
and U17267 (N_17267,N_17079,N_17014);
nand U17268 (N_17268,N_17101,N_17083);
nand U17269 (N_17269,N_17164,N_17157);
or U17270 (N_17270,N_17111,N_17060);
nand U17271 (N_17271,N_17081,N_17194);
xnor U17272 (N_17272,N_17133,N_17067);
xnor U17273 (N_17273,N_17034,N_17010);
and U17274 (N_17274,N_17165,N_17139);
xnor U17275 (N_17275,N_17199,N_17031);
and U17276 (N_17276,N_17138,N_17075);
or U17277 (N_17277,N_17124,N_17136);
nand U17278 (N_17278,N_17190,N_17127);
nor U17279 (N_17279,N_17018,N_17140);
xor U17280 (N_17280,N_17110,N_17163);
xnor U17281 (N_17281,N_17156,N_17137);
or U17282 (N_17282,N_17178,N_17065);
xnor U17283 (N_17283,N_17027,N_17093);
nor U17284 (N_17284,N_17103,N_17086);
nor U17285 (N_17285,N_17181,N_17053);
and U17286 (N_17286,N_17008,N_17131);
nand U17287 (N_17287,N_17019,N_17122);
and U17288 (N_17288,N_17175,N_17003);
nand U17289 (N_17289,N_17146,N_17056);
nor U17290 (N_17290,N_17047,N_17158);
or U17291 (N_17291,N_17168,N_17148);
or U17292 (N_17292,N_17076,N_17100);
and U17293 (N_17293,N_17151,N_17038);
nand U17294 (N_17294,N_17159,N_17145);
nand U17295 (N_17295,N_17049,N_17091);
xnor U17296 (N_17296,N_17050,N_17115);
nand U17297 (N_17297,N_17012,N_17051);
or U17298 (N_17298,N_17029,N_17114);
xnor U17299 (N_17299,N_17046,N_17117);
xor U17300 (N_17300,N_17160,N_17044);
nand U17301 (N_17301,N_17167,N_17087);
nor U17302 (N_17302,N_17023,N_17067);
xnor U17303 (N_17303,N_17092,N_17167);
xor U17304 (N_17304,N_17091,N_17116);
or U17305 (N_17305,N_17185,N_17065);
nor U17306 (N_17306,N_17190,N_17135);
or U17307 (N_17307,N_17000,N_17176);
xnor U17308 (N_17308,N_17049,N_17118);
or U17309 (N_17309,N_17065,N_17150);
xnor U17310 (N_17310,N_17139,N_17128);
xnor U17311 (N_17311,N_17185,N_17089);
xor U17312 (N_17312,N_17016,N_17181);
xnor U17313 (N_17313,N_17139,N_17173);
and U17314 (N_17314,N_17154,N_17043);
nand U17315 (N_17315,N_17179,N_17163);
nand U17316 (N_17316,N_17113,N_17075);
nor U17317 (N_17317,N_17132,N_17037);
and U17318 (N_17318,N_17016,N_17053);
xor U17319 (N_17319,N_17059,N_17167);
nand U17320 (N_17320,N_17186,N_17044);
xor U17321 (N_17321,N_17014,N_17139);
or U17322 (N_17322,N_17171,N_17054);
nand U17323 (N_17323,N_17028,N_17110);
nand U17324 (N_17324,N_17155,N_17026);
xnor U17325 (N_17325,N_17059,N_17126);
nand U17326 (N_17326,N_17055,N_17104);
nor U17327 (N_17327,N_17195,N_17147);
xor U17328 (N_17328,N_17091,N_17051);
or U17329 (N_17329,N_17174,N_17157);
or U17330 (N_17330,N_17144,N_17185);
or U17331 (N_17331,N_17005,N_17014);
nor U17332 (N_17332,N_17063,N_17184);
or U17333 (N_17333,N_17004,N_17169);
or U17334 (N_17334,N_17183,N_17128);
nand U17335 (N_17335,N_17007,N_17196);
and U17336 (N_17336,N_17144,N_17145);
xor U17337 (N_17337,N_17125,N_17143);
xnor U17338 (N_17338,N_17005,N_17092);
nand U17339 (N_17339,N_17032,N_17040);
and U17340 (N_17340,N_17126,N_17122);
nand U17341 (N_17341,N_17160,N_17028);
or U17342 (N_17342,N_17102,N_17040);
nand U17343 (N_17343,N_17164,N_17079);
or U17344 (N_17344,N_17145,N_17164);
and U17345 (N_17345,N_17170,N_17088);
nor U17346 (N_17346,N_17097,N_17119);
xnor U17347 (N_17347,N_17148,N_17173);
nor U17348 (N_17348,N_17068,N_17050);
xnor U17349 (N_17349,N_17044,N_17169);
and U17350 (N_17350,N_17083,N_17002);
nor U17351 (N_17351,N_17002,N_17171);
nor U17352 (N_17352,N_17038,N_17060);
and U17353 (N_17353,N_17118,N_17164);
or U17354 (N_17354,N_17146,N_17121);
or U17355 (N_17355,N_17138,N_17046);
nor U17356 (N_17356,N_17037,N_17107);
or U17357 (N_17357,N_17173,N_17057);
nand U17358 (N_17358,N_17179,N_17100);
or U17359 (N_17359,N_17192,N_17095);
or U17360 (N_17360,N_17027,N_17194);
and U17361 (N_17361,N_17000,N_17133);
xnor U17362 (N_17362,N_17121,N_17112);
nand U17363 (N_17363,N_17060,N_17152);
nor U17364 (N_17364,N_17125,N_17145);
or U17365 (N_17365,N_17036,N_17062);
or U17366 (N_17366,N_17134,N_17058);
nand U17367 (N_17367,N_17066,N_17109);
nor U17368 (N_17368,N_17058,N_17189);
or U17369 (N_17369,N_17087,N_17162);
or U17370 (N_17370,N_17141,N_17010);
or U17371 (N_17371,N_17073,N_17085);
or U17372 (N_17372,N_17071,N_17032);
nand U17373 (N_17373,N_17044,N_17089);
nand U17374 (N_17374,N_17078,N_17003);
and U17375 (N_17375,N_17148,N_17070);
nand U17376 (N_17376,N_17071,N_17116);
nor U17377 (N_17377,N_17083,N_17125);
or U17378 (N_17378,N_17021,N_17082);
and U17379 (N_17379,N_17069,N_17142);
and U17380 (N_17380,N_17103,N_17132);
xor U17381 (N_17381,N_17054,N_17199);
nor U17382 (N_17382,N_17070,N_17004);
xor U17383 (N_17383,N_17056,N_17162);
and U17384 (N_17384,N_17147,N_17122);
xnor U17385 (N_17385,N_17135,N_17157);
or U17386 (N_17386,N_17045,N_17124);
xor U17387 (N_17387,N_17025,N_17003);
xnor U17388 (N_17388,N_17047,N_17060);
nand U17389 (N_17389,N_17024,N_17130);
xnor U17390 (N_17390,N_17017,N_17141);
nor U17391 (N_17391,N_17160,N_17114);
xor U17392 (N_17392,N_17106,N_17042);
and U17393 (N_17393,N_17128,N_17113);
or U17394 (N_17394,N_17136,N_17110);
nor U17395 (N_17395,N_17190,N_17156);
and U17396 (N_17396,N_17167,N_17116);
nor U17397 (N_17397,N_17047,N_17049);
nor U17398 (N_17398,N_17177,N_17071);
nor U17399 (N_17399,N_17191,N_17157);
or U17400 (N_17400,N_17289,N_17265);
or U17401 (N_17401,N_17261,N_17361);
and U17402 (N_17402,N_17344,N_17272);
or U17403 (N_17403,N_17293,N_17247);
nor U17404 (N_17404,N_17214,N_17352);
xnor U17405 (N_17405,N_17300,N_17309);
and U17406 (N_17406,N_17369,N_17365);
or U17407 (N_17407,N_17224,N_17276);
nand U17408 (N_17408,N_17207,N_17371);
or U17409 (N_17409,N_17345,N_17304);
and U17410 (N_17410,N_17322,N_17288);
or U17411 (N_17411,N_17241,N_17318);
nor U17412 (N_17412,N_17399,N_17251);
xor U17413 (N_17413,N_17294,N_17372);
nand U17414 (N_17414,N_17366,N_17301);
xor U17415 (N_17415,N_17228,N_17308);
nor U17416 (N_17416,N_17230,N_17200);
nand U17417 (N_17417,N_17271,N_17392);
and U17418 (N_17418,N_17397,N_17394);
or U17419 (N_17419,N_17331,N_17270);
or U17420 (N_17420,N_17215,N_17296);
xor U17421 (N_17421,N_17235,N_17395);
xor U17422 (N_17422,N_17226,N_17256);
nand U17423 (N_17423,N_17375,N_17238);
or U17424 (N_17424,N_17209,N_17391);
nor U17425 (N_17425,N_17257,N_17274);
or U17426 (N_17426,N_17273,N_17396);
or U17427 (N_17427,N_17355,N_17266);
nand U17428 (N_17428,N_17259,N_17347);
nand U17429 (N_17429,N_17232,N_17383);
nand U17430 (N_17430,N_17389,N_17337);
nand U17431 (N_17431,N_17370,N_17386);
nand U17432 (N_17432,N_17341,N_17313);
xnor U17433 (N_17433,N_17326,N_17217);
nor U17434 (N_17434,N_17282,N_17306);
nand U17435 (N_17435,N_17390,N_17393);
nor U17436 (N_17436,N_17373,N_17292);
xor U17437 (N_17437,N_17220,N_17385);
or U17438 (N_17438,N_17280,N_17245);
and U17439 (N_17439,N_17335,N_17284);
or U17440 (N_17440,N_17240,N_17277);
and U17441 (N_17441,N_17219,N_17317);
or U17442 (N_17442,N_17242,N_17367);
xor U17443 (N_17443,N_17260,N_17298);
nor U17444 (N_17444,N_17269,N_17229);
xnor U17445 (N_17445,N_17210,N_17204);
and U17446 (N_17446,N_17312,N_17233);
nor U17447 (N_17447,N_17384,N_17286);
xnor U17448 (N_17448,N_17246,N_17223);
xor U17449 (N_17449,N_17380,N_17249);
or U17450 (N_17450,N_17354,N_17332);
xor U17451 (N_17451,N_17205,N_17333);
or U17452 (N_17452,N_17303,N_17348);
nor U17453 (N_17453,N_17221,N_17325);
and U17454 (N_17454,N_17315,N_17360);
and U17455 (N_17455,N_17218,N_17324);
xor U17456 (N_17456,N_17263,N_17329);
and U17457 (N_17457,N_17237,N_17234);
nor U17458 (N_17458,N_17202,N_17239);
and U17459 (N_17459,N_17227,N_17358);
and U17460 (N_17460,N_17314,N_17213);
or U17461 (N_17461,N_17252,N_17350);
nand U17462 (N_17462,N_17336,N_17378);
and U17463 (N_17463,N_17216,N_17248);
nor U17464 (N_17464,N_17334,N_17291);
or U17465 (N_17465,N_17363,N_17244);
xor U17466 (N_17466,N_17340,N_17330);
or U17467 (N_17467,N_17243,N_17305);
and U17468 (N_17468,N_17287,N_17381);
xnor U17469 (N_17469,N_17342,N_17253);
xor U17470 (N_17470,N_17353,N_17338);
or U17471 (N_17471,N_17250,N_17320);
or U17472 (N_17472,N_17255,N_17225);
nand U17473 (N_17473,N_17254,N_17379);
or U17474 (N_17474,N_17349,N_17374);
nand U17475 (N_17475,N_17368,N_17307);
xnor U17476 (N_17476,N_17264,N_17281);
nor U17477 (N_17477,N_17290,N_17327);
or U17478 (N_17478,N_17203,N_17268);
nand U17479 (N_17479,N_17357,N_17302);
xnor U17480 (N_17480,N_17211,N_17323);
xnor U17481 (N_17481,N_17316,N_17319);
or U17482 (N_17482,N_17206,N_17295);
nand U17483 (N_17483,N_17258,N_17359);
nand U17484 (N_17484,N_17278,N_17364);
and U17485 (N_17485,N_17362,N_17339);
xor U17486 (N_17486,N_17377,N_17387);
or U17487 (N_17487,N_17285,N_17328);
and U17488 (N_17488,N_17275,N_17346);
xnor U17489 (N_17489,N_17311,N_17388);
nand U17490 (N_17490,N_17351,N_17231);
or U17491 (N_17491,N_17222,N_17398);
nand U17492 (N_17492,N_17201,N_17283);
nand U17493 (N_17493,N_17382,N_17267);
nor U17494 (N_17494,N_17356,N_17262);
nor U17495 (N_17495,N_17321,N_17212);
and U17496 (N_17496,N_17208,N_17343);
or U17497 (N_17497,N_17299,N_17376);
and U17498 (N_17498,N_17236,N_17279);
and U17499 (N_17499,N_17297,N_17310);
nor U17500 (N_17500,N_17301,N_17353);
and U17501 (N_17501,N_17330,N_17395);
and U17502 (N_17502,N_17207,N_17316);
nand U17503 (N_17503,N_17385,N_17323);
xnor U17504 (N_17504,N_17323,N_17265);
or U17505 (N_17505,N_17342,N_17258);
or U17506 (N_17506,N_17240,N_17207);
or U17507 (N_17507,N_17205,N_17321);
or U17508 (N_17508,N_17280,N_17337);
and U17509 (N_17509,N_17304,N_17207);
xnor U17510 (N_17510,N_17283,N_17234);
and U17511 (N_17511,N_17293,N_17287);
nand U17512 (N_17512,N_17283,N_17223);
nor U17513 (N_17513,N_17271,N_17274);
and U17514 (N_17514,N_17339,N_17347);
and U17515 (N_17515,N_17224,N_17306);
and U17516 (N_17516,N_17226,N_17260);
or U17517 (N_17517,N_17377,N_17310);
and U17518 (N_17518,N_17312,N_17305);
or U17519 (N_17519,N_17358,N_17326);
or U17520 (N_17520,N_17369,N_17233);
xor U17521 (N_17521,N_17329,N_17211);
or U17522 (N_17522,N_17390,N_17225);
and U17523 (N_17523,N_17261,N_17291);
and U17524 (N_17524,N_17380,N_17220);
nor U17525 (N_17525,N_17258,N_17214);
nand U17526 (N_17526,N_17342,N_17372);
xnor U17527 (N_17527,N_17318,N_17399);
nor U17528 (N_17528,N_17394,N_17375);
nor U17529 (N_17529,N_17353,N_17357);
nand U17530 (N_17530,N_17392,N_17349);
nor U17531 (N_17531,N_17374,N_17384);
and U17532 (N_17532,N_17388,N_17239);
or U17533 (N_17533,N_17257,N_17382);
nor U17534 (N_17534,N_17365,N_17212);
nor U17535 (N_17535,N_17381,N_17377);
and U17536 (N_17536,N_17236,N_17310);
xor U17537 (N_17537,N_17374,N_17318);
nor U17538 (N_17538,N_17317,N_17385);
nand U17539 (N_17539,N_17210,N_17353);
xor U17540 (N_17540,N_17391,N_17282);
nand U17541 (N_17541,N_17376,N_17317);
xor U17542 (N_17542,N_17374,N_17311);
xor U17543 (N_17543,N_17304,N_17296);
nand U17544 (N_17544,N_17306,N_17278);
and U17545 (N_17545,N_17377,N_17314);
nor U17546 (N_17546,N_17230,N_17316);
nand U17547 (N_17547,N_17325,N_17316);
nor U17548 (N_17548,N_17228,N_17248);
nor U17549 (N_17549,N_17237,N_17209);
and U17550 (N_17550,N_17384,N_17298);
xnor U17551 (N_17551,N_17290,N_17339);
nand U17552 (N_17552,N_17278,N_17370);
nor U17553 (N_17553,N_17276,N_17294);
nor U17554 (N_17554,N_17241,N_17302);
nand U17555 (N_17555,N_17251,N_17373);
and U17556 (N_17556,N_17396,N_17378);
nor U17557 (N_17557,N_17222,N_17347);
xnor U17558 (N_17558,N_17245,N_17210);
xnor U17559 (N_17559,N_17336,N_17386);
and U17560 (N_17560,N_17319,N_17248);
and U17561 (N_17561,N_17314,N_17237);
or U17562 (N_17562,N_17389,N_17233);
or U17563 (N_17563,N_17211,N_17366);
and U17564 (N_17564,N_17366,N_17236);
nand U17565 (N_17565,N_17214,N_17346);
and U17566 (N_17566,N_17220,N_17201);
nand U17567 (N_17567,N_17243,N_17399);
xor U17568 (N_17568,N_17270,N_17353);
nand U17569 (N_17569,N_17234,N_17365);
and U17570 (N_17570,N_17252,N_17390);
nand U17571 (N_17571,N_17268,N_17262);
nand U17572 (N_17572,N_17389,N_17390);
and U17573 (N_17573,N_17322,N_17202);
xor U17574 (N_17574,N_17226,N_17399);
xnor U17575 (N_17575,N_17361,N_17288);
nor U17576 (N_17576,N_17319,N_17268);
and U17577 (N_17577,N_17285,N_17213);
and U17578 (N_17578,N_17210,N_17344);
or U17579 (N_17579,N_17206,N_17277);
xor U17580 (N_17580,N_17306,N_17221);
xor U17581 (N_17581,N_17203,N_17339);
nand U17582 (N_17582,N_17363,N_17230);
xnor U17583 (N_17583,N_17310,N_17238);
xor U17584 (N_17584,N_17226,N_17259);
xnor U17585 (N_17585,N_17284,N_17268);
and U17586 (N_17586,N_17377,N_17318);
or U17587 (N_17587,N_17215,N_17272);
nor U17588 (N_17588,N_17380,N_17229);
nor U17589 (N_17589,N_17289,N_17232);
xnor U17590 (N_17590,N_17271,N_17390);
or U17591 (N_17591,N_17362,N_17306);
or U17592 (N_17592,N_17313,N_17294);
nand U17593 (N_17593,N_17201,N_17365);
xor U17594 (N_17594,N_17329,N_17356);
and U17595 (N_17595,N_17222,N_17283);
nor U17596 (N_17596,N_17342,N_17210);
nor U17597 (N_17597,N_17285,N_17248);
or U17598 (N_17598,N_17357,N_17212);
or U17599 (N_17599,N_17304,N_17328);
or U17600 (N_17600,N_17526,N_17401);
nor U17601 (N_17601,N_17423,N_17472);
nor U17602 (N_17602,N_17504,N_17407);
nor U17603 (N_17603,N_17537,N_17413);
and U17604 (N_17604,N_17575,N_17490);
nor U17605 (N_17605,N_17498,N_17559);
and U17606 (N_17606,N_17597,N_17454);
nand U17607 (N_17607,N_17469,N_17480);
and U17608 (N_17608,N_17534,N_17539);
nand U17609 (N_17609,N_17594,N_17515);
nor U17610 (N_17610,N_17556,N_17543);
xor U17611 (N_17611,N_17506,N_17592);
xor U17612 (N_17612,N_17493,N_17536);
and U17613 (N_17613,N_17446,N_17478);
nand U17614 (N_17614,N_17570,N_17557);
nand U17615 (N_17615,N_17421,N_17591);
nand U17616 (N_17616,N_17548,N_17488);
xor U17617 (N_17617,N_17447,N_17513);
xnor U17618 (N_17618,N_17462,N_17468);
nand U17619 (N_17619,N_17538,N_17475);
nand U17620 (N_17620,N_17520,N_17517);
nor U17621 (N_17621,N_17579,N_17562);
nand U17622 (N_17622,N_17400,N_17542);
and U17623 (N_17623,N_17551,N_17561);
or U17624 (N_17624,N_17435,N_17598);
nor U17625 (N_17625,N_17408,N_17463);
or U17626 (N_17626,N_17477,N_17524);
and U17627 (N_17627,N_17405,N_17596);
nor U17628 (N_17628,N_17574,N_17521);
nand U17629 (N_17629,N_17495,N_17431);
or U17630 (N_17630,N_17494,N_17585);
and U17631 (N_17631,N_17569,N_17560);
and U17632 (N_17632,N_17587,N_17403);
or U17633 (N_17633,N_17424,N_17530);
nand U17634 (N_17634,N_17415,N_17476);
and U17635 (N_17635,N_17540,N_17568);
and U17636 (N_17636,N_17426,N_17471);
and U17637 (N_17637,N_17558,N_17564);
nor U17638 (N_17638,N_17547,N_17550);
nand U17639 (N_17639,N_17440,N_17467);
or U17640 (N_17640,N_17406,N_17442);
nand U17641 (N_17641,N_17450,N_17546);
or U17642 (N_17642,N_17503,N_17554);
xor U17643 (N_17643,N_17438,N_17528);
nor U17644 (N_17644,N_17582,N_17418);
nand U17645 (N_17645,N_17437,N_17419);
nor U17646 (N_17646,N_17500,N_17483);
or U17647 (N_17647,N_17492,N_17588);
nor U17648 (N_17648,N_17573,N_17518);
or U17649 (N_17649,N_17531,N_17441);
or U17650 (N_17650,N_17527,N_17566);
nand U17651 (N_17651,N_17460,N_17402);
nand U17652 (N_17652,N_17510,N_17416);
nand U17653 (N_17653,N_17535,N_17571);
xor U17654 (N_17654,N_17464,N_17482);
nand U17655 (N_17655,N_17411,N_17599);
nand U17656 (N_17656,N_17507,N_17481);
nand U17657 (N_17657,N_17514,N_17451);
nand U17658 (N_17658,N_17410,N_17457);
xnor U17659 (N_17659,N_17448,N_17443);
and U17660 (N_17660,N_17544,N_17436);
or U17661 (N_17661,N_17412,N_17455);
xnor U17662 (N_17662,N_17549,N_17496);
nor U17663 (N_17663,N_17529,N_17577);
xnor U17664 (N_17664,N_17502,N_17473);
or U17665 (N_17665,N_17470,N_17586);
xor U17666 (N_17666,N_17453,N_17555);
xor U17667 (N_17667,N_17512,N_17525);
and U17668 (N_17668,N_17580,N_17439);
xor U17669 (N_17669,N_17414,N_17474);
nor U17670 (N_17670,N_17428,N_17461);
or U17671 (N_17671,N_17523,N_17466);
and U17672 (N_17672,N_17430,N_17589);
xor U17673 (N_17673,N_17417,N_17583);
and U17674 (N_17674,N_17489,N_17445);
xor U17675 (N_17675,N_17516,N_17459);
and U17676 (N_17676,N_17563,N_17509);
nand U17677 (N_17677,N_17576,N_17572);
nor U17678 (N_17678,N_17422,N_17499);
xor U17679 (N_17679,N_17501,N_17541);
nor U17680 (N_17680,N_17545,N_17409);
xor U17681 (N_17681,N_17567,N_17456);
nor U17682 (N_17682,N_17420,N_17434);
and U17683 (N_17683,N_17565,N_17491);
xor U17684 (N_17684,N_17427,N_17595);
or U17685 (N_17685,N_17511,N_17465);
and U17686 (N_17686,N_17487,N_17404);
nand U17687 (N_17687,N_17479,N_17486);
nand U17688 (N_17688,N_17533,N_17458);
nor U17689 (N_17689,N_17584,N_17449);
and U17690 (N_17690,N_17578,N_17505);
and U17691 (N_17691,N_17581,N_17552);
or U17692 (N_17692,N_17425,N_17485);
and U17693 (N_17693,N_17432,N_17444);
nor U17694 (N_17694,N_17532,N_17497);
nor U17695 (N_17695,N_17590,N_17593);
nand U17696 (N_17696,N_17429,N_17519);
xor U17697 (N_17697,N_17433,N_17452);
or U17698 (N_17698,N_17508,N_17522);
and U17699 (N_17699,N_17484,N_17553);
or U17700 (N_17700,N_17513,N_17433);
or U17701 (N_17701,N_17587,N_17406);
xnor U17702 (N_17702,N_17475,N_17424);
nand U17703 (N_17703,N_17416,N_17474);
nor U17704 (N_17704,N_17569,N_17545);
xnor U17705 (N_17705,N_17408,N_17484);
or U17706 (N_17706,N_17403,N_17422);
or U17707 (N_17707,N_17517,N_17531);
nand U17708 (N_17708,N_17587,N_17599);
xnor U17709 (N_17709,N_17403,N_17590);
nor U17710 (N_17710,N_17485,N_17412);
xor U17711 (N_17711,N_17406,N_17496);
nand U17712 (N_17712,N_17570,N_17441);
and U17713 (N_17713,N_17529,N_17471);
nand U17714 (N_17714,N_17527,N_17470);
or U17715 (N_17715,N_17416,N_17531);
and U17716 (N_17716,N_17452,N_17453);
or U17717 (N_17717,N_17583,N_17594);
or U17718 (N_17718,N_17587,N_17467);
and U17719 (N_17719,N_17500,N_17442);
nor U17720 (N_17720,N_17407,N_17525);
xor U17721 (N_17721,N_17400,N_17567);
nand U17722 (N_17722,N_17503,N_17469);
nor U17723 (N_17723,N_17594,N_17559);
xnor U17724 (N_17724,N_17497,N_17400);
or U17725 (N_17725,N_17443,N_17510);
xnor U17726 (N_17726,N_17524,N_17579);
and U17727 (N_17727,N_17580,N_17488);
nand U17728 (N_17728,N_17570,N_17438);
and U17729 (N_17729,N_17487,N_17575);
xor U17730 (N_17730,N_17599,N_17524);
and U17731 (N_17731,N_17595,N_17459);
and U17732 (N_17732,N_17582,N_17546);
xnor U17733 (N_17733,N_17538,N_17554);
and U17734 (N_17734,N_17459,N_17590);
xor U17735 (N_17735,N_17432,N_17544);
and U17736 (N_17736,N_17582,N_17495);
xor U17737 (N_17737,N_17503,N_17526);
or U17738 (N_17738,N_17559,N_17556);
nand U17739 (N_17739,N_17440,N_17405);
xnor U17740 (N_17740,N_17597,N_17496);
and U17741 (N_17741,N_17400,N_17595);
and U17742 (N_17742,N_17577,N_17567);
nand U17743 (N_17743,N_17426,N_17593);
or U17744 (N_17744,N_17464,N_17409);
nor U17745 (N_17745,N_17426,N_17468);
xnor U17746 (N_17746,N_17433,N_17424);
nor U17747 (N_17747,N_17596,N_17566);
xnor U17748 (N_17748,N_17415,N_17547);
nand U17749 (N_17749,N_17400,N_17587);
or U17750 (N_17750,N_17567,N_17489);
nor U17751 (N_17751,N_17495,N_17538);
nor U17752 (N_17752,N_17549,N_17543);
nor U17753 (N_17753,N_17526,N_17488);
xor U17754 (N_17754,N_17568,N_17498);
nand U17755 (N_17755,N_17471,N_17593);
nor U17756 (N_17756,N_17415,N_17493);
nand U17757 (N_17757,N_17505,N_17529);
nand U17758 (N_17758,N_17490,N_17478);
and U17759 (N_17759,N_17481,N_17502);
nand U17760 (N_17760,N_17481,N_17460);
and U17761 (N_17761,N_17571,N_17479);
nor U17762 (N_17762,N_17550,N_17544);
nand U17763 (N_17763,N_17429,N_17527);
and U17764 (N_17764,N_17443,N_17540);
nand U17765 (N_17765,N_17588,N_17505);
nor U17766 (N_17766,N_17509,N_17456);
xor U17767 (N_17767,N_17486,N_17503);
nor U17768 (N_17768,N_17452,N_17438);
and U17769 (N_17769,N_17513,N_17558);
and U17770 (N_17770,N_17478,N_17495);
or U17771 (N_17771,N_17547,N_17554);
nor U17772 (N_17772,N_17571,N_17423);
and U17773 (N_17773,N_17509,N_17529);
xnor U17774 (N_17774,N_17565,N_17451);
and U17775 (N_17775,N_17520,N_17444);
and U17776 (N_17776,N_17545,N_17568);
and U17777 (N_17777,N_17489,N_17493);
and U17778 (N_17778,N_17446,N_17475);
and U17779 (N_17779,N_17451,N_17462);
xnor U17780 (N_17780,N_17526,N_17500);
nand U17781 (N_17781,N_17574,N_17542);
xor U17782 (N_17782,N_17418,N_17461);
or U17783 (N_17783,N_17457,N_17517);
nor U17784 (N_17784,N_17540,N_17509);
and U17785 (N_17785,N_17470,N_17431);
and U17786 (N_17786,N_17438,N_17493);
or U17787 (N_17787,N_17497,N_17486);
xor U17788 (N_17788,N_17550,N_17404);
nand U17789 (N_17789,N_17491,N_17410);
nand U17790 (N_17790,N_17573,N_17482);
nand U17791 (N_17791,N_17454,N_17462);
xnor U17792 (N_17792,N_17549,N_17536);
or U17793 (N_17793,N_17455,N_17503);
xor U17794 (N_17794,N_17468,N_17470);
nor U17795 (N_17795,N_17476,N_17478);
xor U17796 (N_17796,N_17433,N_17483);
and U17797 (N_17797,N_17444,N_17515);
and U17798 (N_17798,N_17480,N_17507);
or U17799 (N_17799,N_17424,N_17460);
and U17800 (N_17800,N_17789,N_17683);
nand U17801 (N_17801,N_17739,N_17622);
nand U17802 (N_17802,N_17704,N_17730);
nor U17803 (N_17803,N_17763,N_17773);
or U17804 (N_17804,N_17641,N_17639);
nor U17805 (N_17805,N_17708,N_17626);
and U17806 (N_17806,N_17729,N_17666);
and U17807 (N_17807,N_17621,N_17676);
xor U17808 (N_17808,N_17712,N_17681);
and U17809 (N_17809,N_17718,N_17726);
and U17810 (N_17810,N_17790,N_17647);
and U17811 (N_17811,N_17757,N_17689);
and U17812 (N_17812,N_17664,N_17637);
nand U17813 (N_17813,N_17736,N_17693);
xnor U17814 (N_17814,N_17652,N_17651);
or U17815 (N_17815,N_17768,N_17677);
xor U17816 (N_17816,N_17684,N_17728);
xnor U17817 (N_17817,N_17662,N_17692);
or U17818 (N_17818,N_17737,N_17770);
nand U17819 (N_17819,N_17719,N_17654);
xor U17820 (N_17820,N_17752,N_17608);
nand U17821 (N_17821,N_17786,N_17782);
xor U17822 (N_17822,N_17743,N_17754);
and U17823 (N_17823,N_17611,N_17791);
and U17824 (N_17824,N_17795,N_17706);
and U17825 (N_17825,N_17631,N_17648);
or U17826 (N_17826,N_17784,N_17727);
and U17827 (N_17827,N_17705,N_17682);
xnor U17828 (N_17828,N_17643,N_17673);
xor U17829 (N_17829,N_17620,N_17694);
and U17830 (N_17830,N_17794,N_17649);
or U17831 (N_17831,N_17640,N_17615);
nor U17832 (N_17832,N_17765,N_17613);
or U17833 (N_17833,N_17783,N_17630);
xnor U17834 (N_17834,N_17634,N_17685);
xor U17835 (N_17835,N_17711,N_17655);
nor U17836 (N_17836,N_17687,N_17690);
and U17837 (N_17837,N_17760,N_17788);
and U17838 (N_17838,N_17638,N_17761);
and U17839 (N_17839,N_17781,N_17632);
nor U17840 (N_17840,N_17793,N_17753);
xor U17841 (N_17841,N_17715,N_17751);
and U17842 (N_17842,N_17619,N_17656);
nand U17843 (N_17843,N_17635,N_17735);
xor U17844 (N_17844,N_17720,N_17721);
and U17845 (N_17845,N_17710,N_17755);
nand U17846 (N_17846,N_17688,N_17742);
xnor U17847 (N_17847,N_17623,N_17778);
nand U17848 (N_17848,N_17600,N_17602);
or U17849 (N_17849,N_17799,N_17725);
nor U17850 (N_17850,N_17767,N_17766);
and U17851 (N_17851,N_17776,N_17741);
xnor U17852 (N_17852,N_17624,N_17775);
nand U17853 (N_17853,N_17700,N_17695);
nor U17854 (N_17854,N_17774,N_17732);
and U17855 (N_17855,N_17716,N_17644);
and U17856 (N_17856,N_17702,N_17738);
xor U17857 (N_17857,N_17747,N_17612);
or U17858 (N_17858,N_17653,N_17678);
nand U17859 (N_17859,N_17750,N_17714);
nor U17860 (N_17860,N_17625,N_17764);
and U17861 (N_17861,N_17731,N_17713);
or U17862 (N_17862,N_17796,N_17792);
nor U17863 (N_17863,N_17675,N_17745);
nor U17864 (N_17864,N_17628,N_17646);
nor U17865 (N_17865,N_17603,N_17645);
nor U17866 (N_17866,N_17629,N_17609);
xor U17867 (N_17867,N_17663,N_17618);
or U17868 (N_17868,N_17642,N_17733);
nand U17869 (N_17869,N_17659,N_17698);
or U17870 (N_17870,N_17748,N_17616);
or U17871 (N_17871,N_17758,N_17779);
xnor U17872 (N_17872,N_17769,N_17671);
and U17873 (N_17873,N_17756,N_17746);
and U17874 (N_17874,N_17749,N_17691);
xor U17875 (N_17875,N_17787,N_17772);
and U17876 (N_17876,N_17606,N_17670);
nor U17877 (N_17877,N_17798,N_17762);
nand U17878 (N_17878,N_17701,N_17657);
nor U17879 (N_17879,N_17679,N_17601);
xnor U17880 (N_17880,N_17680,N_17744);
xnor U17881 (N_17881,N_17667,N_17607);
xnor U17882 (N_17882,N_17717,N_17660);
xor U17883 (N_17883,N_17780,N_17658);
nor U17884 (N_17884,N_17636,N_17771);
and U17885 (N_17885,N_17604,N_17650);
nand U17886 (N_17886,N_17759,N_17665);
nand U17887 (N_17887,N_17740,N_17703);
xnor U17888 (N_17888,N_17724,N_17777);
and U17889 (N_17889,N_17699,N_17674);
xnor U17890 (N_17890,N_17686,N_17723);
nor U17891 (N_17891,N_17697,N_17627);
nand U17892 (N_17892,N_17785,N_17614);
or U17893 (N_17893,N_17668,N_17610);
xor U17894 (N_17894,N_17672,N_17707);
and U17895 (N_17895,N_17661,N_17734);
nor U17896 (N_17896,N_17633,N_17617);
xor U17897 (N_17897,N_17709,N_17797);
xor U17898 (N_17898,N_17605,N_17696);
or U17899 (N_17899,N_17669,N_17722);
nand U17900 (N_17900,N_17707,N_17787);
nor U17901 (N_17901,N_17781,N_17651);
xor U17902 (N_17902,N_17746,N_17682);
nor U17903 (N_17903,N_17689,N_17710);
and U17904 (N_17904,N_17606,N_17723);
or U17905 (N_17905,N_17609,N_17745);
xnor U17906 (N_17906,N_17765,N_17628);
nand U17907 (N_17907,N_17621,N_17760);
xor U17908 (N_17908,N_17662,N_17793);
and U17909 (N_17909,N_17637,N_17750);
xor U17910 (N_17910,N_17698,N_17667);
and U17911 (N_17911,N_17622,N_17697);
and U17912 (N_17912,N_17770,N_17773);
xnor U17913 (N_17913,N_17778,N_17767);
or U17914 (N_17914,N_17642,N_17675);
xnor U17915 (N_17915,N_17770,N_17649);
and U17916 (N_17916,N_17797,N_17750);
nor U17917 (N_17917,N_17675,N_17794);
or U17918 (N_17918,N_17628,N_17741);
nand U17919 (N_17919,N_17763,N_17680);
xnor U17920 (N_17920,N_17701,N_17779);
nand U17921 (N_17921,N_17634,N_17682);
nand U17922 (N_17922,N_17678,N_17665);
nor U17923 (N_17923,N_17747,N_17727);
and U17924 (N_17924,N_17692,N_17794);
xnor U17925 (N_17925,N_17700,N_17620);
xor U17926 (N_17926,N_17616,N_17689);
nor U17927 (N_17927,N_17632,N_17643);
nand U17928 (N_17928,N_17603,N_17724);
or U17929 (N_17929,N_17673,N_17782);
nand U17930 (N_17930,N_17666,N_17681);
xnor U17931 (N_17931,N_17629,N_17716);
and U17932 (N_17932,N_17753,N_17766);
nor U17933 (N_17933,N_17779,N_17659);
nand U17934 (N_17934,N_17668,N_17685);
and U17935 (N_17935,N_17771,N_17775);
or U17936 (N_17936,N_17611,N_17767);
nor U17937 (N_17937,N_17776,N_17707);
and U17938 (N_17938,N_17641,N_17774);
or U17939 (N_17939,N_17712,N_17618);
nand U17940 (N_17940,N_17697,N_17703);
nor U17941 (N_17941,N_17770,N_17762);
nand U17942 (N_17942,N_17686,N_17680);
nand U17943 (N_17943,N_17646,N_17638);
or U17944 (N_17944,N_17661,N_17738);
xnor U17945 (N_17945,N_17686,N_17773);
nor U17946 (N_17946,N_17634,N_17623);
and U17947 (N_17947,N_17688,N_17616);
nand U17948 (N_17948,N_17658,N_17642);
or U17949 (N_17949,N_17689,N_17778);
xnor U17950 (N_17950,N_17620,N_17768);
and U17951 (N_17951,N_17678,N_17622);
xnor U17952 (N_17952,N_17623,N_17735);
and U17953 (N_17953,N_17778,N_17659);
and U17954 (N_17954,N_17652,N_17716);
or U17955 (N_17955,N_17703,N_17747);
nand U17956 (N_17956,N_17711,N_17667);
xnor U17957 (N_17957,N_17789,N_17721);
and U17958 (N_17958,N_17791,N_17751);
and U17959 (N_17959,N_17747,N_17744);
xor U17960 (N_17960,N_17788,N_17676);
nand U17961 (N_17961,N_17735,N_17753);
xnor U17962 (N_17962,N_17711,N_17653);
and U17963 (N_17963,N_17752,N_17612);
or U17964 (N_17964,N_17646,N_17716);
and U17965 (N_17965,N_17626,N_17767);
nor U17966 (N_17966,N_17726,N_17715);
nand U17967 (N_17967,N_17784,N_17789);
and U17968 (N_17968,N_17637,N_17672);
nand U17969 (N_17969,N_17666,N_17708);
nor U17970 (N_17970,N_17640,N_17741);
nor U17971 (N_17971,N_17648,N_17695);
nor U17972 (N_17972,N_17605,N_17673);
nor U17973 (N_17973,N_17675,N_17760);
nor U17974 (N_17974,N_17723,N_17738);
xor U17975 (N_17975,N_17732,N_17794);
or U17976 (N_17976,N_17662,N_17656);
and U17977 (N_17977,N_17635,N_17774);
and U17978 (N_17978,N_17647,N_17793);
nor U17979 (N_17979,N_17752,N_17688);
xnor U17980 (N_17980,N_17761,N_17660);
nor U17981 (N_17981,N_17616,N_17782);
xnor U17982 (N_17982,N_17694,N_17753);
and U17983 (N_17983,N_17763,N_17724);
nor U17984 (N_17984,N_17725,N_17633);
and U17985 (N_17985,N_17696,N_17738);
nor U17986 (N_17986,N_17743,N_17735);
or U17987 (N_17987,N_17744,N_17696);
nor U17988 (N_17988,N_17794,N_17756);
nor U17989 (N_17989,N_17608,N_17751);
or U17990 (N_17990,N_17633,N_17761);
or U17991 (N_17991,N_17651,N_17799);
xor U17992 (N_17992,N_17696,N_17656);
nand U17993 (N_17993,N_17686,N_17646);
nor U17994 (N_17994,N_17654,N_17689);
and U17995 (N_17995,N_17704,N_17789);
nor U17996 (N_17996,N_17789,N_17794);
nand U17997 (N_17997,N_17796,N_17716);
nand U17998 (N_17998,N_17766,N_17725);
and U17999 (N_17999,N_17779,N_17610);
nor U18000 (N_18000,N_17963,N_17835);
or U18001 (N_18001,N_17980,N_17820);
xnor U18002 (N_18002,N_17983,N_17882);
nand U18003 (N_18003,N_17833,N_17848);
xor U18004 (N_18004,N_17839,N_17809);
and U18005 (N_18005,N_17818,N_17807);
nor U18006 (N_18006,N_17940,N_17805);
nor U18007 (N_18007,N_17808,N_17878);
nor U18008 (N_18008,N_17959,N_17895);
nand U18009 (N_18009,N_17975,N_17933);
nand U18010 (N_18010,N_17854,N_17864);
or U18011 (N_18011,N_17969,N_17894);
nor U18012 (N_18012,N_17921,N_17948);
nor U18013 (N_18013,N_17986,N_17887);
or U18014 (N_18014,N_17923,N_17967);
nor U18015 (N_18015,N_17919,N_17852);
and U18016 (N_18016,N_17806,N_17982);
nor U18017 (N_18017,N_17996,N_17965);
and U18018 (N_18018,N_17821,N_17896);
nor U18019 (N_18019,N_17960,N_17961);
or U18020 (N_18020,N_17814,N_17883);
or U18021 (N_18021,N_17881,N_17911);
nand U18022 (N_18022,N_17897,N_17800);
or U18023 (N_18023,N_17968,N_17999);
nand U18024 (N_18024,N_17804,N_17870);
nand U18025 (N_18025,N_17927,N_17861);
and U18026 (N_18026,N_17838,N_17908);
or U18027 (N_18027,N_17802,N_17928);
nor U18028 (N_18028,N_17836,N_17992);
nand U18029 (N_18029,N_17958,N_17872);
nor U18030 (N_18030,N_17931,N_17850);
nor U18031 (N_18031,N_17834,N_17981);
and U18032 (N_18032,N_17966,N_17823);
nor U18033 (N_18033,N_17817,N_17873);
and U18034 (N_18034,N_17916,N_17841);
nor U18035 (N_18035,N_17830,N_17810);
nor U18036 (N_18036,N_17903,N_17946);
or U18037 (N_18037,N_17890,N_17867);
or U18038 (N_18038,N_17912,N_17939);
xnor U18039 (N_18039,N_17902,N_17970);
xor U18040 (N_18040,N_17950,N_17846);
nand U18041 (N_18041,N_17913,N_17879);
and U18042 (N_18042,N_17816,N_17888);
and U18043 (N_18043,N_17801,N_17899);
nor U18044 (N_18044,N_17866,N_17917);
nor U18045 (N_18045,N_17853,N_17952);
nor U18046 (N_18046,N_17974,N_17844);
xnor U18047 (N_18047,N_17877,N_17837);
xnor U18048 (N_18048,N_17865,N_17856);
xor U18049 (N_18049,N_17932,N_17987);
nand U18050 (N_18050,N_17842,N_17825);
xnor U18051 (N_18051,N_17910,N_17937);
xnor U18052 (N_18052,N_17860,N_17874);
and U18053 (N_18053,N_17924,N_17811);
and U18054 (N_18054,N_17957,N_17824);
nor U18055 (N_18055,N_17972,N_17956);
or U18056 (N_18056,N_17847,N_17951);
or U18057 (N_18057,N_17925,N_17871);
or U18058 (N_18058,N_17934,N_17914);
nor U18059 (N_18059,N_17953,N_17828);
nand U18060 (N_18060,N_17898,N_17971);
nor U18061 (N_18061,N_17857,N_17995);
xnor U18062 (N_18062,N_17851,N_17858);
nor U18063 (N_18063,N_17979,N_17826);
and U18064 (N_18064,N_17984,N_17884);
or U18065 (N_18065,N_17892,N_17901);
and U18066 (N_18066,N_17926,N_17930);
nand U18067 (N_18067,N_17922,N_17949);
nand U18068 (N_18068,N_17822,N_17920);
nand U18069 (N_18069,N_17812,N_17875);
and U18070 (N_18070,N_17889,N_17863);
and U18071 (N_18071,N_17880,N_17954);
nand U18072 (N_18072,N_17915,N_17905);
nor U18073 (N_18073,N_17827,N_17904);
nor U18074 (N_18074,N_17997,N_17843);
nor U18075 (N_18075,N_17989,N_17815);
xor U18076 (N_18076,N_17985,N_17998);
xnor U18077 (N_18077,N_17977,N_17849);
nand U18078 (N_18078,N_17876,N_17907);
nand U18079 (N_18079,N_17973,N_17900);
xnor U18080 (N_18080,N_17993,N_17909);
or U18081 (N_18081,N_17906,N_17893);
nor U18082 (N_18082,N_17976,N_17938);
nor U18083 (N_18083,N_17991,N_17941);
nor U18084 (N_18084,N_17845,N_17813);
xor U18085 (N_18085,N_17942,N_17929);
and U18086 (N_18086,N_17947,N_17955);
xnor U18087 (N_18087,N_17819,N_17832);
nand U18088 (N_18088,N_17945,N_17885);
and U18089 (N_18089,N_17829,N_17840);
xor U18090 (N_18090,N_17990,N_17964);
or U18091 (N_18091,N_17855,N_17862);
xor U18092 (N_18092,N_17988,N_17831);
and U18093 (N_18093,N_17935,N_17869);
and U18094 (N_18094,N_17803,N_17868);
xnor U18095 (N_18095,N_17886,N_17891);
and U18096 (N_18096,N_17994,N_17859);
or U18097 (N_18097,N_17962,N_17978);
xor U18098 (N_18098,N_17918,N_17944);
nand U18099 (N_18099,N_17943,N_17936);
nand U18100 (N_18100,N_17866,N_17807);
nand U18101 (N_18101,N_17983,N_17853);
nand U18102 (N_18102,N_17934,N_17944);
nand U18103 (N_18103,N_17915,N_17844);
or U18104 (N_18104,N_17851,N_17978);
nand U18105 (N_18105,N_17987,N_17813);
nand U18106 (N_18106,N_17973,N_17849);
and U18107 (N_18107,N_17804,N_17855);
and U18108 (N_18108,N_17871,N_17982);
xor U18109 (N_18109,N_17915,N_17950);
and U18110 (N_18110,N_17926,N_17834);
xor U18111 (N_18111,N_17936,N_17859);
and U18112 (N_18112,N_17983,N_17921);
nand U18113 (N_18113,N_17863,N_17941);
xor U18114 (N_18114,N_17988,N_17953);
or U18115 (N_18115,N_17805,N_17910);
xnor U18116 (N_18116,N_17902,N_17955);
or U18117 (N_18117,N_17916,N_17801);
and U18118 (N_18118,N_17975,N_17885);
nand U18119 (N_18119,N_17956,N_17917);
nor U18120 (N_18120,N_17924,N_17831);
and U18121 (N_18121,N_17832,N_17985);
and U18122 (N_18122,N_17892,N_17978);
and U18123 (N_18123,N_17914,N_17892);
nor U18124 (N_18124,N_17858,N_17995);
or U18125 (N_18125,N_17801,N_17965);
xor U18126 (N_18126,N_17986,N_17815);
and U18127 (N_18127,N_17888,N_17916);
nand U18128 (N_18128,N_17901,N_17903);
or U18129 (N_18129,N_17934,N_17920);
xor U18130 (N_18130,N_17873,N_17900);
or U18131 (N_18131,N_17812,N_17877);
xor U18132 (N_18132,N_17991,N_17892);
nor U18133 (N_18133,N_17837,N_17858);
xor U18134 (N_18134,N_17899,N_17944);
and U18135 (N_18135,N_17817,N_17810);
and U18136 (N_18136,N_17965,N_17980);
and U18137 (N_18137,N_17954,N_17853);
xor U18138 (N_18138,N_17872,N_17920);
nor U18139 (N_18139,N_17828,N_17860);
and U18140 (N_18140,N_17931,N_17924);
xor U18141 (N_18141,N_17815,N_17964);
xor U18142 (N_18142,N_17945,N_17980);
and U18143 (N_18143,N_17889,N_17841);
nand U18144 (N_18144,N_17815,N_17821);
and U18145 (N_18145,N_17879,N_17919);
nor U18146 (N_18146,N_17882,N_17963);
xnor U18147 (N_18147,N_17904,N_17938);
nor U18148 (N_18148,N_17962,N_17990);
and U18149 (N_18149,N_17978,N_17959);
and U18150 (N_18150,N_17931,N_17922);
nor U18151 (N_18151,N_17912,N_17977);
and U18152 (N_18152,N_17817,N_17845);
nor U18153 (N_18153,N_17889,N_17972);
or U18154 (N_18154,N_17883,N_17900);
and U18155 (N_18155,N_17978,N_17953);
nor U18156 (N_18156,N_17989,N_17829);
nor U18157 (N_18157,N_17902,N_17929);
or U18158 (N_18158,N_17929,N_17925);
and U18159 (N_18159,N_17838,N_17888);
or U18160 (N_18160,N_17953,N_17863);
nor U18161 (N_18161,N_17979,N_17987);
and U18162 (N_18162,N_17941,N_17885);
or U18163 (N_18163,N_17823,N_17906);
nand U18164 (N_18164,N_17872,N_17964);
xor U18165 (N_18165,N_17904,N_17921);
or U18166 (N_18166,N_17838,N_17999);
or U18167 (N_18167,N_17869,N_17823);
nor U18168 (N_18168,N_17982,N_17863);
nor U18169 (N_18169,N_17976,N_17887);
nand U18170 (N_18170,N_17865,N_17838);
nor U18171 (N_18171,N_17975,N_17893);
or U18172 (N_18172,N_17836,N_17993);
nand U18173 (N_18173,N_17960,N_17944);
and U18174 (N_18174,N_17938,N_17885);
xnor U18175 (N_18175,N_17963,N_17863);
nor U18176 (N_18176,N_17968,N_17867);
or U18177 (N_18177,N_17899,N_17921);
nor U18178 (N_18178,N_17834,N_17921);
or U18179 (N_18179,N_17929,N_17828);
and U18180 (N_18180,N_17800,N_17801);
nor U18181 (N_18181,N_17826,N_17932);
or U18182 (N_18182,N_17894,N_17919);
and U18183 (N_18183,N_17850,N_17824);
nor U18184 (N_18184,N_17867,N_17813);
and U18185 (N_18185,N_17810,N_17818);
and U18186 (N_18186,N_17807,N_17831);
xor U18187 (N_18187,N_17993,N_17824);
nor U18188 (N_18188,N_17992,N_17945);
nor U18189 (N_18189,N_17953,N_17982);
nand U18190 (N_18190,N_17924,N_17953);
xnor U18191 (N_18191,N_17986,N_17833);
and U18192 (N_18192,N_17877,N_17960);
xor U18193 (N_18193,N_17992,N_17875);
nand U18194 (N_18194,N_17826,N_17977);
nor U18195 (N_18195,N_17950,N_17975);
nand U18196 (N_18196,N_17830,N_17959);
nand U18197 (N_18197,N_17965,N_17991);
nor U18198 (N_18198,N_17901,N_17921);
and U18199 (N_18199,N_17888,N_17955);
or U18200 (N_18200,N_18173,N_18051);
xnor U18201 (N_18201,N_18171,N_18089);
nor U18202 (N_18202,N_18197,N_18053);
or U18203 (N_18203,N_18008,N_18014);
xor U18204 (N_18204,N_18195,N_18085);
or U18205 (N_18205,N_18184,N_18021);
nand U18206 (N_18206,N_18097,N_18078);
xor U18207 (N_18207,N_18086,N_18146);
nand U18208 (N_18208,N_18028,N_18136);
and U18209 (N_18209,N_18161,N_18090);
or U18210 (N_18210,N_18133,N_18128);
nand U18211 (N_18211,N_18149,N_18134);
nand U18212 (N_18212,N_18026,N_18072);
or U18213 (N_18213,N_18169,N_18162);
nor U18214 (N_18214,N_18007,N_18054);
and U18215 (N_18215,N_18144,N_18187);
nand U18216 (N_18216,N_18125,N_18073);
and U18217 (N_18217,N_18063,N_18045);
or U18218 (N_18218,N_18104,N_18101);
xnor U18219 (N_18219,N_18003,N_18015);
nand U18220 (N_18220,N_18009,N_18175);
nor U18221 (N_18221,N_18194,N_18127);
xnor U18222 (N_18222,N_18040,N_18132);
or U18223 (N_18223,N_18177,N_18099);
xnor U18224 (N_18224,N_18172,N_18034);
or U18225 (N_18225,N_18141,N_18048);
nor U18226 (N_18226,N_18036,N_18105);
xnor U18227 (N_18227,N_18140,N_18057);
or U18228 (N_18228,N_18055,N_18186);
xnor U18229 (N_18229,N_18166,N_18093);
and U18230 (N_18230,N_18096,N_18150);
nor U18231 (N_18231,N_18060,N_18157);
nand U18232 (N_18232,N_18155,N_18153);
and U18233 (N_18233,N_18147,N_18022);
nand U18234 (N_18234,N_18091,N_18016);
xor U18235 (N_18235,N_18081,N_18083);
nand U18236 (N_18236,N_18118,N_18043);
nand U18237 (N_18237,N_18154,N_18182);
nand U18238 (N_18238,N_18124,N_18044);
nor U18239 (N_18239,N_18075,N_18106);
xor U18240 (N_18240,N_18029,N_18095);
nand U18241 (N_18241,N_18061,N_18148);
and U18242 (N_18242,N_18114,N_18019);
nand U18243 (N_18243,N_18084,N_18199);
and U18244 (N_18244,N_18145,N_18117);
nor U18245 (N_18245,N_18087,N_18137);
xnor U18246 (N_18246,N_18102,N_18005);
or U18247 (N_18247,N_18107,N_18004);
and U18248 (N_18248,N_18024,N_18049);
xor U18249 (N_18249,N_18039,N_18030);
xor U18250 (N_18250,N_18143,N_18192);
xnor U18251 (N_18251,N_18109,N_18188);
nor U18252 (N_18252,N_18158,N_18066);
or U18253 (N_18253,N_18038,N_18065);
nor U18254 (N_18254,N_18165,N_18151);
xnor U18255 (N_18255,N_18198,N_18047);
nand U18256 (N_18256,N_18167,N_18018);
nand U18257 (N_18257,N_18135,N_18006);
xnor U18258 (N_18258,N_18176,N_18010);
nor U18259 (N_18259,N_18120,N_18079);
nor U18260 (N_18260,N_18142,N_18160);
xor U18261 (N_18261,N_18023,N_18002);
xor U18262 (N_18262,N_18011,N_18183);
xnor U18263 (N_18263,N_18068,N_18103);
or U18264 (N_18264,N_18112,N_18031);
nand U18265 (N_18265,N_18138,N_18163);
nand U18266 (N_18266,N_18070,N_18001);
nor U18267 (N_18267,N_18092,N_18035);
nand U18268 (N_18268,N_18115,N_18174);
xor U18269 (N_18269,N_18111,N_18168);
nand U18270 (N_18270,N_18067,N_18178);
nor U18271 (N_18271,N_18121,N_18046);
and U18272 (N_18272,N_18041,N_18069);
or U18273 (N_18273,N_18185,N_18159);
or U18274 (N_18274,N_18110,N_18170);
and U18275 (N_18275,N_18179,N_18020);
nor U18276 (N_18276,N_18094,N_18122);
and U18277 (N_18277,N_18130,N_18033);
nand U18278 (N_18278,N_18074,N_18077);
nand U18279 (N_18279,N_18050,N_18116);
nand U18280 (N_18280,N_18058,N_18156);
xnor U18281 (N_18281,N_18100,N_18000);
or U18282 (N_18282,N_18052,N_18013);
and U18283 (N_18283,N_18080,N_18126);
xnor U18284 (N_18284,N_18076,N_18098);
nor U18285 (N_18285,N_18071,N_18012);
xnor U18286 (N_18286,N_18181,N_18113);
nor U18287 (N_18287,N_18189,N_18088);
xnor U18288 (N_18288,N_18082,N_18062);
xor U18289 (N_18289,N_18017,N_18064);
xor U18290 (N_18290,N_18123,N_18193);
xnor U18291 (N_18291,N_18190,N_18042);
and U18292 (N_18292,N_18059,N_18129);
nand U18293 (N_18293,N_18056,N_18196);
or U18294 (N_18294,N_18139,N_18131);
and U18295 (N_18295,N_18180,N_18032);
nor U18296 (N_18296,N_18025,N_18027);
or U18297 (N_18297,N_18037,N_18108);
and U18298 (N_18298,N_18119,N_18152);
or U18299 (N_18299,N_18164,N_18191);
nand U18300 (N_18300,N_18195,N_18104);
xnor U18301 (N_18301,N_18032,N_18174);
and U18302 (N_18302,N_18049,N_18127);
nor U18303 (N_18303,N_18065,N_18033);
or U18304 (N_18304,N_18017,N_18180);
nor U18305 (N_18305,N_18107,N_18034);
nand U18306 (N_18306,N_18155,N_18006);
or U18307 (N_18307,N_18086,N_18069);
or U18308 (N_18308,N_18125,N_18011);
and U18309 (N_18309,N_18110,N_18191);
or U18310 (N_18310,N_18095,N_18190);
xor U18311 (N_18311,N_18106,N_18051);
nand U18312 (N_18312,N_18109,N_18152);
nand U18313 (N_18313,N_18096,N_18149);
and U18314 (N_18314,N_18118,N_18194);
or U18315 (N_18315,N_18044,N_18195);
xnor U18316 (N_18316,N_18168,N_18189);
nor U18317 (N_18317,N_18020,N_18150);
xnor U18318 (N_18318,N_18106,N_18030);
nor U18319 (N_18319,N_18048,N_18098);
nor U18320 (N_18320,N_18067,N_18043);
xnor U18321 (N_18321,N_18065,N_18192);
and U18322 (N_18322,N_18040,N_18171);
or U18323 (N_18323,N_18054,N_18099);
nor U18324 (N_18324,N_18074,N_18174);
nand U18325 (N_18325,N_18017,N_18113);
nand U18326 (N_18326,N_18185,N_18122);
nand U18327 (N_18327,N_18120,N_18105);
nor U18328 (N_18328,N_18056,N_18177);
nor U18329 (N_18329,N_18000,N_18184);
xor U18330 (N_18330,N_18120,N_18181);
or U18331 (N_18331,N_18011,N_18151);
nor U18332 (N_18332,N_18013,N_18123);
nand U18333 (N_18333,N_18137,N_18053);
xor U18334 (N_18334,N_18170,N_18195);
xor U18335 (N_18335,N_18065,N_18159);
xnor U18336 (N_18336,N_18024,N_18084);
and U18337 (N_18337,N_18011,N_18143);
and U18338 (N_18338,N_18120,N_18062);
nand U18339 (N_18339,N_18129,N_18198);
nor U18340 (N_18340,N_18172,N_18052);
and U18341 (N_18341,N_18125,N_18057);
xor U18342 (N_18342,N_18048,N_18050);
or U18343 (N_18343,N_18061,N_18035);
and U18344 (N_18344,N_18135,N_18003);
or U18345 (N_18345,N_18034,N_18122);
nor U18346 (N_18346,N_18019,N_18194);
xnor U18347 (N_18347,N_18046,N_18103);
nand U18348 (N_18348,N_18034,N_18016);
or U18349 (N_18349,N_18181,N_18079);
and U18350 (N_18350,N_18172,N_18183);
xnor U18351 (N_18351,N_18136,N_18067);
nand U18352 (N_18352,N_18011,N_18177);
nor U18353 (N_18353,N_18151,N_18189);
nand U18354 (N_18354,N_18052,N_18050);
and U18355 (N_18355,N_18183,N_18131);
and U18356 (N_18356,N_18164,N_18142);
and U18357 (N_18357,N_18089,N_18197);
nor U18358 (N_18358,N_18071,N_18198);
or U18359 (N_18359,N_18122,N_18003);
and U18360 (N_18360,N_18064,N_18085);
nor U18361 (N_18361,N_18000,N_18067);
or U18362 (N_18362,N_18067,N_18110);
or U18363 (N_18363,N_18121,N_18150);
xnor U18364 (N_18364,N_18093,N_18149);
xor U18365 (N_18365,N_18058,N_18003);
nand U18366 (N_18366,N_18066,N_18017);
nor U18367 (N_18367,N_18091,N_18035);
or U18368 (N_18368,N_18112,N_18197);
xor U18369 (N_18369,N_18059,N_18096);
nor U18370 (N_18370,N_18077,N_18006);
xor U18371 (N_18371,N_18152,N_18193);
or U18372 (N_18372,N_18139,N_18134);
or U18373 (N_18373,N_18132,N_18118);
nand U18374 (N_18374,N_18052,N_18133);
or U18375 (N_18375,N_18017,N_18174);
or U18376 (N_18376,N_18019,N_18146);
nand U18377 (N_18377,N_18174,N_18055);
or U18378 (N_18378,N_18104,N_18156);
or U18379 (N_18379,N_18092,N_18136);
or U18380 (N_18380,N_18015,N_18155);
and U18381 (N_18381,N_18124,N_18001);
xor U18382 (N_18382,N_18089,N_18182);
or U18383 (N_18383,N_18000,N_18120);
and U18384 (N_18384,N_18058,N_18108);
xor U18385 (N_18385,N_18165,N_18109);
and U18386 (N_18386,N_18116,N_18031);
and U18387 (N_18387,N_18117,N_18050);
nand U18388 (N_18388,N_18060,N_18075);
nor U18389 (N_18389,N_18058,N_18124);
nor U18390 (N_18390,N_18035,N_18018);
or U18391 (N_18391,N_18152,N_18173);
xnor U18392 (N_18392,N_18003,N_18179);
and U18393 (N_18393,N_18128,N_18058);
or U18394 (N_18394,N_18070,N_18188);
xnor U18395 (N_18395,N_18018,N_18147);
nand U18396 (N_18396,N_18016,N_18139);
or U18397 (N_18397,N_18173,N_18070);
xnor U18398 (N_18398,N_18098,N_18040);
or U18399 (N_18399,N_18186,N_18121);
or U18400 (N_18400,N_18321,N_18218);
or U18401 (N_18401,N_18287,N_18225);
and U18402 (N_18402,N_18342,N_18290);
xnor U18403 (N_18403,N_18212,N_18214);
xor U18404 (N_18404,N_18327,N_18242);
nor U18405 (N_18405,N_18394,N_18313);
and U18406 (N_18406,N_18357,N_18215);
nor U18407 (N_18407,N_18333,N_18314);
nand U18408 (N_18408,N_18339,N_18228);
xnor U18409 (N_18409,N_18326,N_18344);
xor U18410 (N_18410,N_18237,N_18234);
and U18411 (N_18411,N_18292,N_18373);
and U18412 (N_18412,N_18389,N_18244);
and U18413 (N_18413,N_18289,N_18251);
nand U18414 (N_18414,N_18220,N_18209);
xnor U18415 (N_18415,N_18345,N_18227);
or U18416 (N_18416,N_18391,N_18278);
nand U18417 (N_18417,N_18248,N_18211);
and U18418 (N_18418,N_18388,N_18294);
or U18419 (N_18419,N_18386,N_18265);
or U18420 (N_18420,N_18281,N_18208);
or U18421 (N_18421,N_18332,N_18359);
xnor U18422 (N_18422,N_18396,N_18243);
nor U18423 (N_18423,N_18207,N_18328);
nand U18424 (N_18424,N_18239,N_18219);
nand U18425 (N_18425,N_18360,N_18379);
nand U18426 (N_18426,N_18368,N_18270);
nor U18427 (N_18427,N_18329,N_18201);
nand U18428 (N_18428,N_18341,N_18323);
nor U18429 (N_18429,N_18267,N_18399);
nand U18430 (N_18430,N_18262,N_18249);
nand U18431 (N_18431,N_18306,N_18307);
xor U18432 (N_18432,N_18320,N_18277);
and U18433 (N_18433,N_18305,N_18376);
xor U18434 (N_18434,N_18318,N_18216);
nand U18435 (N_18435,N_18362,N_18253);
or U18436 (N_18436,N_18238,N_18334);
or U18437 (N_18437,N_18392,N_18246);
and U18438 (N_18438,N_18365,N_18263);
nand U18439 (N_18439,N_18247,N_18347);
nor U18440 (N_18440,N_18202,N_18203);
xnor U18441 (N_18441,N_18271,N_18351);
xnor U18442 (N_18442,N_18395,N_18297);
and U18443 (N_18443,N_18390,N_18268);
or U18444 (N_18444,N_18380,N_18325);
and U18445 (N_18445,N_18363,N_18322);
xor U18446 (N_18446,N_18222,N_18298);
or U18447 (N_18447,N_18301,N_18282);
nor U18448 (N_18448,N_18276,N_18335);
xnor U18449 (N_18449,N_18261,N_18346);
and U18450 (N_18450,N_18358,N_18230);
nor U18451 (N_18451,N_18378,N_18293);
nand U18452 (N_18452,N_18284,N_18235);
or U18453 (N_18453,N_18217,N_18223);
xor U18454 (N_18454,N_18309,N_18349);
and U18455 (N_18455,N_18353,N_18348);
nand U18456 (N_18456,N_18303,N_18264);
or U18457 (N_18457,N_18317,N_18393);
and U18458 (N_18458,N_18210,N_18331);
and U18459 (N_18459,N_18383,N_18308);
xnor U18460 (N_18460,N_18352,N_18260);
nor U18461 (N_18461,N_18275,N_18355);
xor U18462 (N_18462,N_18224,N_18385);
nand U18463 (N_18463,N_18254,N_18371);
or U18464 (N_18464,N_18377,N_18205);
and U18465 (N_18465,N_18319,N_18374);
nor U18466 (N_18466,N_18255,N_18231);
and U18467 (N_18467,N_18367,N_18382);
xor U18468 (N_18468,N_18397,N_18233);
and U18469 (N_18469,N_18279,N_18310);
xnor U18470 (N_18470,N_18296,N_18300);
xor U18471 (N_18471,N_18245,N_18384);
nor U18472 (N_18472,N_18252,N_18288);
and U18473 (N_18473,N_18213,N_18398);
xnor U18474 (N_18474,N_18259,N_18299);
xnor U18475 (N_18475,N_18302,N_18257);
or U18476 (N_18476,N_18272,N_18258);
or U18477 (N_18477,N_18356,N_18250);
or U18478 (N_18478,N_18283,N_18204);
and U18479 (N_18479,N_18240,N_18266);
nand U18480 (N_18480,N_18269,N_18336);
nor U18481 (N_18481,N_18316,N_18295);
nor U18482 (N_18482,N_18387,N_18350);
and U18483 (N_18483,N_18337,N_18256);
nor U18484 (N_18484,N_18311,N_18241);
and U18485 (N_18485,N_18324,N_18343);
or U18486 (N_18486,N_18274,N_18372);
or U18487 (N_18487,N_18200,N_18232);
xnor U18488 (N_18488,N_18338,N_18330);
and U18489 (N_18489,N_18221,N_18369);
xor U18490 (N_18490,N_18236,N_18361);
nor U18491 (N_18491,N_18291,N_18229);
or U18492 (N_18492,N_18226,N_18354);
or U18493 (N_18493,N_18381,N_18286);
and U18494 (N_18494,N_18315,N_18206);
nor U18495 (N_18495,N_18273,N_18370);
and U18496 (N_18496,N_18280,N_18340);
and U18497 (N_18497,N_18285,N_18366);
nor U18498 (N_18498,N_18312,N_18364);
and U18499 (N_18499,N_18304,N_18375);
xnor U18500 (N_18500,N_18383,N_18281);
and U18501 (N_18501,N_18259,N_18334);
xor U18502 (N_18502,N_18393,N_18321);
and U18503 (N_18503,N_18325,N_18387);
nand U18504 (N_18504,N_18289,N_18236);
xor U18505 (N_18505,N_18204,N_18377);
xnor U18506 (N_18506,N_18247,N_18217);
and U18507 (N_18507,N_18244,N_18367);
and U18508 (N_18508,N_18230,N_18282);
or U18509 (N_18509,N_18396,N_18350);
nand U18510 (N_18510,N_18229,N_18324);
nor U18511 (N_18511,N_18295,N_18379);
and U18512 (N_18512,N_18293,N_18398);
and U18513 (N_18513,N_18391,N_18289);
nand U18514 (N_18514,N_18306,N_18351);
xnor U18515 (N_18515,N_18351,N_18291);
and U18516 (N_18516,N_18372,N_18233);
or U18517 (N_18517,N_18298,N_18363);
nor U18518 (N_18518,N_18311,N_18235);
xnor U18519 (N_18519,N_18362,N_18236);
nand U18520 (N_18520,N_18366,N_18221);
and U18521 (N_18521,N_18371,N_18279);
nand U18522 (N_18522,N_18350,N_18291);
xnor U18523 (N_18523,N_18232,N_18231);
and U18524 (N_18524,N_18351,N_18374);
and U18525 (N_18525,N_18345,N_18209);
and U18526 (N_18526,N_18391,N_18310);
or U18527 (N_18527,N_18201,N_18275);
or U18528 (N_18528,N_18283,N_18308);
or U18529 (N_18529,N_18258,N_18346);
or U18530 (N_18530,N_18356,N_18282);
and U18531 (N_18531,N_18231,N_18332);
or U18532 (N_18532,N_18303,N_18286);
or U18533 (N_18533,N_18216,N_18341);
or U18534 (N_18534,N_18283,N_18216);
nor U18535 (N_18535,N_18231,N_18337);
xnor U18536 (N_18536,N_18385,N_18371);
or U18537 (N_18537,N_18348,N_18235);
nand U18538 (N_18538,N_18255,N_18270);
or U18539 (N_18539,N_18265,N_18304);
xor U18540 (N_18540,N_18224,N_18375);
nand U18541 (N_18541,N_18300,N_18264);
nand U18542 (N_18542,N_18219,N_18252);
nand U18543 (N_18543,N_18297,N_18241);
or U18544 (N_18544,N_18253,N_18279);
or U18545 (N_18545,N_18218,N_18394);
or U18546 (N_18546,N_18203,N_18379);
nand U18547 (N_18547,N_18311,N_18267);
or U18548 (N_18548,N_18218,N_18236);
or U18549 (N_18549,N_18296,N_18382);
and U18550 (N_18550,N_18219,N_18369);
xor U18551 (N_18551,N_18203,N_18256);
xor U18552 (N_18552,N_18214,N_18294);
nor U18553 (N_18553,N_18314,N_18376);
or U18554 (N_18554,N_18235,N_18283);
nor U18555 (N_18555,N_18334,N_18233);
nand U18556 (N_18556,N_18287,N_18273);
and U18557 (N_18557,N_18216,N_18311);
nor U18558 (N_18558,N_18351,N_18303);
nand U18559 (N_18559,N_18227,N_18365);
or U18560 (N_18560,N_18233,N_18235);
nand U18561 (N_18561,N_18330,N_18258);
nor U18562 (N_18562,N_18239,N_18275);
nand U18563 (N_18563,N_18367,N_18245);
xnor U18564 (N_18564,N_18392,N_18283);
and U18565 (N_18565,N_18339,N_18250);
nand U18566 (N_18566,N_18392,N_18217);
nor U18567 (N_18567,N_18314,N_18353);
nand U18568 (N_18568,N_18258,N_18390);
xnor U18569 (N_18569,N_18392,N_18216);
nand U18570 (N_18570,N_18299,N_18200);
or U18571 (N_18571,N_18397,N_18257);
xnor U18572 (N_18572,N_18219,N_18245);
or U18573 (N_18573,N_18339,N_18291);
or U18574 (N_18574,N_18289,N_18223);
or U18575 (N_18575,N_18362,N_18206);
nor U18576 (N_18576,N_18339,N_18377);
nand U18577 (N_18577,N_18353,N_18264);
or U18578 (N_18578,N_18301,N_18242);
and U18579 (N_18579,N_18383,N_18224);
nand U18580 (N_18580,N_18275,N_18335);
xor U18581 (N_18581,N_18362,N_18311);
or U18582 (N_18582,N_18201,N_18392);
and U18583 (N_18583,N_18326,N_18284);
nand U18584 (N_18584,N_18315,N_18385);
nor U18585 (N_18585,N_18306,N_18340);
nand U18586 (N_18586,N_18312,N_18205);
or U18587 (N_18587,N_18351,N_18242);
and U18588 (N_18588,N_18263,N_18344);
and U18589 (N_18589,N_18285,N_18290);
and U18590 (N_18590,N_18370,N_18294);
and U18591 (N_18591,N_18207,N_18372);
nor U18592 (N_18592,N_18259,N_18210);
or U18593 (N_18593,N_18268,N_18272);
xnor U18594 (N_18594,N_18370,N_18224);
or U18595 (N_18595,N_18333,N_18283);
xor U18596 (N_18596,N_18247,N_18239);
xnor U18597 (N_18597,N_18393,N_18397);
or U18598 (N_18598,N_18255,N_18315);
and U18599 (N_18599,N_18392,N_18331);
xnor U18600 (N_18600,N_18479,N_18570);
or U18601 (N_18601,N_18580,N_18409);
xnor U18602 (N_18602,N_18463,N_18469);
nor U18603 (N_18603,N_18538,N_18517);
xnor U18604 (N_18604,N_18443,N_18497);
and U18605 (N_18605,N_18412,N_18429);
xor U18606 (N_18606,N_18598,N_18427);
xor U18607 (N_18607,N_18460,N_18439);
xor U18608 (N_18608,N_18430,N_18449);
or U18609 (N_18609,N_18406,N_18554);
or U18610 (N_18610,N_18544,N_18504);
xor U18611 (N_18611,N_18458,N_18532);
nor U18612 (N_18612,N_18572,N_18541);
or U18613 (N_18613,N_18501,N_18540);
and U18614 (N_18614,N_18481,N_18564);
and U18615 (N_18615,N_18550,N_18563);
xnor U18616 (N_18616,N_18405,N_18576);
xnor U18617 (N_18617,N_18592,N_18494);
and U18618 (N_18618,N_18492,N_18596);
or U18619 (N_18619,N_18491,N_18448);
nor U18620 (N_18620,N_18461,N_18431);
and U18621 (N_18621,N_18545,N_18578);
and U18622 (N_18622,N_18509,N_18503);
or U18623 (N_18623,N_18444,N_18586);
xor U18624 (N_18624,N_18599,N_18573);
nor U18625 (N_18625,N_18456,N_18520);
nand U18626 (N_18626,N_18528,N_18574);
and U18627 (N_18627,N_18476,N_18556);
nor U18628 (N_18628,N_18529,N_18459);
and U18629 (N_18629,N_18425,N_18447);
nor U18630 (N_18630,N_18511,N_18557);
and U18631 (N_18631,N_18519,N_18414);
or U18632 (N_18632,N_18416,N_18499);
and U18633 (N_18633,N_18507,N_18558);
nand U18634 (N_18634,N_18483,N_18513);
nand U18635 (N_18635,N_18400,N_18546);
xnor U18636 (N_18636,N_18583,N_18446);
nand U18637 (N_18637,N_18410,N_18506);
and U18638 (N_18638,N_18473,N_18423);
and U18639 (N_18639,N_18471,N_18589);
or U18640 (N_18640,N_18549,N_18522);
nor U18641 (N_18641,N_18445,N_18585);
or U18642 (N_18642,N_18435,N_18560);
xnor U18643 (N_18643,N_18488,N_18486);
and U18644 (N_18644,N_18593,N_18542);
xor U18645 (N_18645,N_18581,N_18547);
nand U18646 (N_18646,N_18407,N_18464);
and U18647 (N_18647,N_18437,N_18417);
or U18648 (N_18648,N_18568,N_18401);
or U18649 (N_18649,N_18434,N_18531);
or U18650 (N_18650,N_18515,N_18595);
and U18651 (N_18651,N_18582,N_18478);
nor U18652 (N_18652,N_18579,N_18575);
or U18653 (N_18653,N_18487,N_18510);
nand U18654 (N_18654,N_18432,N_18590);
nand U18655 (N_18655,N_18455,N_18418);
nand U18656 (N_18656,N_18477,N_18421);
nor U18657 (N_18657,N_18569,N_18553);
nor U18658 (N_18658,N_18404,N_18584);
and U18659 (N_18659,N_18426,N_18587);
nand U18660 (N_18660,N_18440,N_18567);
xnor U18661 (N_18661,N_18502,N_18535);
nand U18662 (N_18662,N_18408,N_18490);
xnor U18663 (N_18663,N_18571,N_18411);
nand U18664 (N_18664,N_18561,N_18548);
nand U18665 (N_18665,N_18462,N_18505);
or U18666 (N_18666,N_18419,N_18493);
xor U18667 (N_18667,N_18527,N_18465);
or U18668 (N_18668,N_18536,N_18597);
and U18669 (N_18669,N_18534,N_18524);
or U18670 (N_18670,N_18450,N_18516);
nor U18671 (N_18671,N_18433,N_18480);
nand U18672 (N_18672,N_18565,N_18415);
xor U18673 (N_18673,N_18424,N_18518);
and U18674 (N_18674,N_18453,N_18514);
nand U18675 (N_18675,N_18533,N_18539);
and U18676 (N_18676,N_18472,N_18403);
and U18677 (N_18677,N_18537,N_18482);
or U18678 (N_18678,N_18438,N_18428);
xnor U18679 (N_18679,N_18454,N_18451);
xnor U18680 (N_18680,N_18489,N_18468);
nand U18681 (N_18681,N_18562,N_18441);
or U18682 (N_18682,N_18594,N_18498);
or U18683 (N_18683,N_18508,N_18466);
nand U18684 (N_18684,N_18484,N_18474);
nand U18685 (N_18685,N_18566,N_18475);
nor U18686 (N_18686,N_18555,N_18577);
nor U18687 (N_18687,N_18467,N_18470);
or U18688 (N_18688,N_18485,N_18496);
and U18689 (N_18689,N_18420,N_18500);
and U18690 (N_18690,N_18551,N_18457);
nor U18691 (N_18691,N_18543,N_18552);
xor U18692 (N_18692,N_18413,N_18422);
or U18693 (N_18693,N_18512,N_18526);
and U18694 (N_18694,N_18591,N_18559);
and U18695 (N_18695,N_18525,N_18521);
nand U18696 (N_18696,N_18402,N_18442);
xnor U18697 (N_18697,N_18523,N_18495);
and U18698 (N_18698,N_18588,N_18452);
xor U18699 (N_18699,N_18436,N_18530);
xnor U18700 (N_18700,N_18527,N_18531);
nand U18701 (N_18701,N_18437,N_18413);
and U18702 (N_18702,N_18449,N_18508);
nand U18703 (N_18703,N_18534,N_18423);
xor U18704 (N_18704,N_18469,N_18475);
or U18705 (N_18705,N_18558,N_18555);
xor U18706 (N_18706,N_18541,N_18575);
nor U18707 (N_18707,N_18439,N_18551);
nand U18708 (N_18708,N_18489,N_18412);
nor U18709 (N_18709,N_18526,N_18597);
nor U18710 (N_18710,N_18445,N_18580);
and U18711 (N_18711,N_18462,N_18578);
and U18712 (N_18712,N_18527,N_18494);
xnor U18713 (N_18713,N_18570,N_18498);
xnor U18714 (N_18714,N_18597,N_18537);
or U18715 (N_18715,N_18504,N_18560);
or U18716 (N_18716,N_18487,N_18489);
or U18717 (N_18717,N_18401,N_18472);
and U18718 (N_18718,N_18463,N_18565);
or U18719 (N_18719,N_18447,N_18533);
nor U18720 (N_18720,N_18582,N_18474);
or U18721 (N_18721,N_18496,N_18498);
xor U18722 (N_18722,N_18598,N_18484);
xnor U18723 (N_18723,N_18509,N_18492);
nor U18724 (N_18724,N_18413,N_18448);
nor U18725 (N_18725,N_18570,N_18458);
nand U18726 (N_18726,N_18538,N_18575);
nand U18727 (N_18727,N_18517,N_18407);
xnor U18728 (N_18728,N_18436,N_18429);
nor U18729 (N_18729,N_18432,N_18525);
and U18730 (N_18730,N_18416,N_18524);
and U18731 (N_18731,N_18480,N_18461);
and U18732 (N_18732,N_18491,N_18407);
or U18733 (N_18733,N_18403,N_18544);
and U18734 (N_18734,N_18486,N_18409);
xnor U18735 (N_18735,N_18445,N_18406);
nor U18736 (N_18736,N_18409,N_18560);
and U18737 (N_18737,N_18483,N_18492);
nand U18738 (N_18738,N_18509,N_18516);
and U18739 (N_18739,N_18434,N_18442);
and U18740 (N_18740,N_18476,N_18429);
nand U18741 (N_18741,N_18549,N_18488);
xor U18742 (N_18742,N_18516,N_18403);
nor U18743 (N_18743,N_18453,N_18523);
nor U18744 (N_18744,N_18457,N_18506);
and U18745 (N_18745,N_18493,N_18510);
xor U18746 (N_18746,N_18528,N_18578);
and U18747 (N_18747,N_18445,N_18541);
nor U18748 (N_18748,N_18572,N_18507);
nor U18749 (N_18749,N_18444,N_18493);
or U18750 (N_18750,N_18552,N_18432);
and U18751 (N_18751,N_18588,N_18585);
xor U18752 (N_18752,N_18410,N_18580);
and U18753 (N_18753,N_18516,N_18423);
or U18754 (N_18754,N_18476,N_18597);
and U18755 (N_18755,N_18546,N_18511);
xnor U18756 (N_18756,N_18523,N_18489);
nand U18757 (N_18757,N_18403,N_18495);
nor U18758 (N_18758,N_18421,N_18587);
nor U18759 (N_18759,N_18559,N_18488);
nor U18760 (N_18760,N_18528,N_18475);
or U18761 (N_18761,N_18401,N_18549);
nand U18762 (N_18762,N_18524,N_18550);
or U18763 (N_18763,N_18532,N_18503);
and U18764 (N_18764,N_18478,N_18469);
xor U18765 (N_18765,N_18552,N_18536);
or U18766 (N_18766,N_18496,N_18413);
nor U18767 (N_18767,N_18525,N_18541);
nand U18768 (N_18768,N_18456,N_18524);
nand U18769 (N_18769,N_18444,N_18448);
and U18770 (N_18770,N_18491,N_18571);
and U18771 (N_18771,N_18442,N_18461);
and U18772 (N_18772,N_18591,N_18497);
nor U18773 (N_18773,N_18410,N_18420);
nor U18774 (N_18774,N_18404,N_18501);
and U18775 (N_18775,N_18528,N_18576);
or U18776 (N_18776,N_18593,N_18572);
or U18777 (N_18777,N_18479,N_18566);
nand U18778 (N_18778,N_18462,N_18546);
xor U18779 (N_18779,N_18484,N_18546);
nand U18780 (N_18780,N_18573,N_18449);
nor U18781 (N_18781,N_18535,N_18461);
nand U18782 (N_18782,N_18506,N_18552);
nor U18783 (N_18783,N_18414,N_18520);
and U18784 (N_18784,N_18400,N_18584);
xnor U18785 (N_18785,N_18446,N_18419);
nor U18786 (N_18786,N_18542,N_18440);
or U18787 (N_18787,N_18552,N_18487);
nor U18788 (N_18788,N_18497,N_18488);
nor U18789 (N_18789,N_18531,N_18439);
and U18790 (N_18790,N_18566,N_18493);
nand U18791 (N_18791,N_18539,N_18549);
xor U18792 (N_18792,N_18416,N_18439);
and U18793 (N_18793,N_18484,N_18446);
nor U18794 (N_18794,N_18537,N_18542);
or U18795 (N_18795,N_18496,N_18591);
and U18796 (N_18796,N_18470,N_18569);
xnor U18797 (N_18797,N_18581,N_18560);
nand U18798 (N_18798,N_18481,N_18488);
nor U18799 (N_18799,N_18453,N_18510);
xor U18800 (N_18800,N_18694,N_18714);
and U18801 (N_18801,N_18666,N_18735);
and U18802 (N_18802,N_18721,N_18682);
xnor U18803 (N_18803,N_18741,N_18753);
nor U18804 (N_18804,N_18709,N_18797);
or U18805 (N_18805,N_18712,N_18609);
and U18806 (N_18806,N_18762,N_18707);
or U18807 (N_18807,N_18605,N_18780);
and U18808 (N_18808,N_18646,N_18670);
or U18809 (N_18809,N_18621,N_18787);
nor U18810 (N_18810,N_18748,N_18789);
or U18811 (N_18811,N_18662,N_18677);
nand U18812 (N_18812,N_18659,N_18760);
or U18813 (N_18813,N_18740,N_18600);
nor U18814 (N_18814,N_18743,N_18726);
or U18815 (N_18815,N_18676,N_18658);
or U18816 (N_18816,N_18624,N_18643);
and U18817 (N_18817,N_18706,N_18655);
or U18818 (N_18818,N_18717,N_18784);
or U18819 (N_18819,N_18631,N_18625);
xnor U18820 (N_18820,N_18751,N_18685);
xor U18821 (N_18821,N_18680,N_18733);
or U18822 (N_18822,N_18757,N_18672);
nor U18823 (N_18823,N_18703,N_18622);
xor U18824 (N_18824,N_18749,N_18696);
nor U18825 (N_18825,N_18610,N_18619);
or U18826 (N_18826,N_18665,N_18771);
nor U18827 (N_18827,N_18661,N_18752);
xor U18828 (N_18828,N_18701,N_18615);
nor U18829 (N_18829,N_18683,N_18794);
or U18830 (N_18830,N_18634,N_18747);
or U18831 (N_18831,N_18776,N_18681);
xnor U18832 (N_18832,N_18795,N_18614);
or U18833 (N_18833,N_18766,N_18732);
or U18834 (N_18834,N_18688,N_18637);
or U18835 (N_18835,N_18710,N_18671);
and U18836 (N_18836,N_18628,N_18723);
xnor U18837 (N_18837,N_18773,N_18768);
and U18838 (N_18838,N_18664,N_18692);
or U18839 (N_18839,N_18746,N_18686);
nor U18840 (N_18840,N_18675,N_18704);
xor U18841 (N_18841,N_18604,N_18779);
nand U18842 (N_18842,N_18744,N_18790);
xnor U18843 (N_18843,N_18636,N_18742);
nand U18844 (N_18844,N_18611,N_18711);
nand U18845 (N_18845,N_18715,N_18679);
nand U18846 (N_18846,N_18695,N_18654);
or U18847 (N_18847,N_18772,N_18651);
xnor U18848 (N_18848,N_18728,N_18668);
xor U18849 (N_18849,N_18754,N_18687);
nor U18850 (N_18850,N_18777,N_18758);
nand U18851 (N_18851,N_18786,N_18775);
nand U18852 (N_18852,N_18799,N_18700);
nor U18853 (N_18853,N_18620,N_18623);
nor U18854 (N_18854,N_18781,N_18645);
xnor U18855 (N_18855,N_18727,N_18761);
nand U18856 (N_18856,N_18647,N_18630);
nand U18857 (N_18857,N_18739,N_18793);
and U18858 (N_18858,N_18756,N_18783);
xnor U18859 (N_18859,N_18719,N_18767);
and U18860 (N_18860,N_18725,N_18638);
xnor U18861 (N_18861,N_18641,N_18750);
and U18862 (N_18862,N_18626,N_18674);
and U18863 (N_18863,N_18649,N_18755);
nor U18864 (N_18864,N_18633,N_18693);
nand U18865 (N_18865,N_18632,N_18653);
nor U18866 (N_18866,N_18607,N_18734);
xnor U18867 (N_18867,N_18603,N_18782);
xor U18868 (N_18868,N_18763,N_18644);
or U18869 (N_18869,N_18698,N_18718);
nor U18870 (N_18870,N_18639,N_18669);
nand U18871 (N_18871,N_18765,N_18730);
and U18872 (N_18872,N_18656,N_18796);
and U18873 (N_18873,N_18764,N_18705);
xnor U18874 (N_18874,N_18697,N_18617);
and U18875 (N_18875,N_18678,N_18660);
nor U18876 (N_18876,N_18788,N_18627);
and U18877 (N_18877,N_18613,N_18720);
or U18878 (N_18878,N_18759,N_18736);
xor U18879 (N_18879,N_18769,N_18798);
or U18880 (N_18880,N_18785,N_18642);
nor U18881 (N_18881,N_18648,N_18663);
and U18882 (N_18882,N_18792,N_18699);
nand U18883 (N_18883,N_18724,N_18778);
or U18884 (N_18884,N_18729,N_18708);
xor U18885 (N_18885,N_18612,N_18657);
nand U18886 (N_18886,N_18629,N_18738);
nand U18887 (N_18887,N_18606,N_18691);
and U18888 (N_18888,N_18608,N_18731);
and U18889 (N_18889,N_18602,N_18722);
and U18890 (N_18890,N_18713,N_18770);
nor U18891 (N_18891,N_18650,N_18635);
xor U18892 (N_18892,N_18601,N_18640);
nand U18893 (N_18893,N_18616,N_18667);
or U18894 (N_18894,N_18745,N_18737);
and U18895 (N_18895,N_18673,N_18684);
xnor U18896 (N_18896,N_18791,N_18689);
or U18897 (N_18897,N_18652,N_18716);
or U18898 (N_18898,N_18690,N_18774);
or U18899 (N_18899,N_18618,N_18702);
nor U18900 (N_18900,N_18689,N_18709);
and U18901 (N_18901,N_18663,N_18694);
or U18902 (N_18902,N_18615,N_18713);
xnor U18903 (N_18903,N_18699,N_18783);
nor U18904 (N_18904,N_18721,N_18625);
nor U18905 (N_18905,N_18690,N_18601);
and U18906 (N_18906,N_18703,N_18794);
xnor U18907 (N_18907,N_18680,N_18634);
nand U18908 (N_18908,N_18679,N_18756);
xnor U18909 (N_18909,N_18755,N_18763);
nor U18910 (N_18910,N_18743,N_18612);
nand U18911 (N_18911,N_18688,N_18765);
or U18912 (N_18912,N_18711,N_18608);
or U18913 (N_18913,N_18678,N_18738);
nand U18914 (N_18914,N_18606,N_18761);
xor U18915 (N_18915,N_18743,N_18635);
xor U18916 (N_18916,N_18651,N_18752);
and U18917 (N_18917,N_18715,N_18739);
nand U18918 (N_18918,N_18719,N_18639);
nor U18919 (N_18919,N_18677,N_18780);
xnor U18920 (N_18920,N_18661,N_18685);
or U18921 (N_18921,N_18670,N_18722);
nand U18922 (N_18922,N_18653,N_18606);
or U18923 (N_18923,N_18791,N_18729);
and U18924 (N_18924,N_18682,N_18713);
nor U18925 (N_18925,N_18754,N_18685);
and U18926 (N_18926,N_18737,N_18629);
xnor U18927 (N_18927,N_18617,N_18619);
or U18928 (N_18928,N_18749,N_18688);
and U18929 (N_18929,N_18715,N_18716);
or U18930 (N_18930,N_18660,N_18625);
or U18931 (N_18931,N_18614,N_18672);
xor U18932 (N_18932,N_18684,N_18781);
xor U18933 (N_18933,N_18710,N_18787);
nor U18934 (N_18934,N_18736,N_18772);
and U18935 (N_18935,N_18693,N_18621);
and U18936 (N_18936,N_18640,N_18622);
and U18937 (N_18937,N_18703,N_18691);
xnor U18938 (N_18938,N_18777,N_18755);
nor U18939 (N_18939,N_18745,N_18603);
nor U18940 (N_18940,N_18778,N_18705);
and U18941 (N_18941,N_18641,N_18734);
nand U18942 (N_18942,N_18757,N_18698);
nor U18943 (N_18943,N_18727,N_18783);
or U18944 (N_18944,N_18776,N_18796);
nand U18945 (N_18945,N_18612,N_18628);
and U18946 (N_18946,N_18767,N_18753);
xor U18947 (N_18947,N_18738,N_18671);
and U18948 (N_18948,N_18629,N_18688);
nand U18949 (N_18949,N_18703,N_18712);
nor U18950 (N_18950,N_18759,N_18614);
xnor U18951 (N_18951,N_18673,N_18669);
xor U18952 (N_18952,N_18682,N_18693);
xor U18953 (N_18953,N_18601,N_18631);
nor U18954 (N_18954,N_18783,N_18618);
xor U18955 (N_18955,N_18713,N_18660);
nand U18956 (N_18956,N_18666,N_18799);
nor U18957 (N_18957,N_18690,N_18612);
or U18958 (N_18958,N_18761,N_18645);
nand U18959 (N_18959,N_18658,N_18643);
or U18960 (N_18960,N_18637,N_18679);
and U18961 (N_18961,N_18737,N_18648);
or U18962 (N_18962,N_18778,N_18670);
or U18963 (N_18963,N_18678,N_18662);
nor U18964 (N_18964,N_18662,N_18688);
and U18965 (N_18965,N_18727,N_18652);
and U18966 (N_18966,N_18797,N_18682);
or U18967 (N_18967,N_18726,N_18738);
or U18968 (N_18968,N_18770,N_18787);
and U18969 (N_18969,N_18600,N_18617);
or U18970 (N_18970,N_18646,N_18787);
xnor U18971 (N_18971,N_18760,N_18684);
nor U18972 (N_18972,N_18791,N_18787);
or U18973 (N_18973,N_18748,N_18675);
and U18974 (N_18974,N_18788,N_18766);
nor U18975 (N_18975,N_18684,N_18697);
nor U18976 (N_18976,N_18613,N_18605);
nand U18977 (N_18977,N_18794,N_18753);
nor U18978 (N_18978,N_18621,N_18663);
and U18979 (N_18979,N_18666,N_18692);
nor U18980 (N_18980,N_18661,N_18722);
xor U18981 (N_18981,N_18703,N_18765);
xnor U18982 (N_18982,N_18778,N_18654);
and U18983 (N_18983,N_18725,N_18667);
xnor U18984 (N_18984,N_18666,N_18685);
or U18985 (N_18985,N_18631,N_18654);
or U18986 (N_18986,N_18732,N_18632);
or U18987 (N_18987,N_18793,N_18624);
nand U18988 (N_18988,N_18687,N_18703);
nand U18989 (N_18989,N_18652,N_18656);
and U18990 (N_18990,N_18618,N_18661);
nor U18991 (N_18991,N_18799,N_18767);
and U18992 (N_18992,N_18686,N_18715);
and U18993 (N_18993,N_18607,N_18671);
or U18994 (N_18994,N_18615,N_18793);
or U18995 (N_18995,N_18633,N_18707);
or U18996 (N_18996,N_18760,N_18761);
or U18997 (N_18997,N_18787,N_18657);
nand U18998 (N_18998,N_18789,N_18655);
xor U18999 (N_18999,N_18692,N_18706);
nand U19000 (N_19000,N_18916,N_18888);
and U19001 (N_19001,N_18945,N_18880);
nor U19002 (N_19002,N_18805,N_18915);
and U19003 (N_19003,N_18820,N_18956);
and U19004 (N_19004,N_18854,N_18839);
nor U19005 (N_19005,N_18816,N_18871);
and U19006 (N_19006,N_18996,N_18911);
nand U19007 (N_19007,N_18931,N_18971);
or U19008 (N_19008,N_18873,N_18906);
and U19009 (N_19009,N_18851,N_18860);
and U19010 (N_19010,N_18987,N_18837);
nand U19011 (N_19011,N_18947,N_18949);
and U19012 (N_19012,N_18998,N_18882);
and U19013 (N_19013,N_18954,N_18898);
nand U19014 (N_19014,N_18813,N_18967);
nand U19015 (N_19015,N_18923,N_18867);
xnor U19016 (N_19016,N_18870,N_18921);
and U19017 (N_19017,N_18908,N_18913);
or U19018 (N_19018,N_18874,N_18876);
xnor U19019 (N_19019,N_18917,N_18830);
nand U19020 (N_19020,N_18843,N_18952);
xnor U19021 (N_19021,N_18853,N_18803);
nor U19022 (N_19022,N_18819,N_18896);
or U19023 (N_19023,N_18920,N_18928);
nand U19024 (N_19024,N_18907,N_18978);
nand U19025 (N_19025,N_18862,N_18857);
xnor U19026 (N_19026,N_18895,N_18881);
and U19027 (N_19027,N_18955,N_18926);
and U19028 (N_19028,N_18840,N_18884);
and U19029 (N_19029,N_18941,N_18994);
nor U19030 (N_19030,N_18958,N_18897);
xor U19031 (N_19031,N_18891,N_18903);
xor U19032 (N_19032,N_18957,N_18815);
nor U19033 (N_19033,N_18997,N_18868);
nor U19034 (N_19034,N_18912,N_18909);
xnor U19035 (N_19035,N_18800,N_18914);
xnor U19036 (N_19036,N_18883,N_18865);
or U19037 (N_19037,N_18834,N_18889);
nand U19038 (N_19038,N_18810,N_18885);
and U19039 (N_19039,N_18801,N_18919);
xnor U19040 (N_19040,N_18948,N_18993);
and U19041 (N_19041,N_18877,N_18864);
nand U19042 (N_19042,N_18965,N_18981);
nor U19043 (N_19043,N_18972,N_18899);
or U19044 (N_19044,N_18910,N_18963);
nor U19045 (N_19045,N_18863,N_18844);
or U19046 (N_19046,N_18959,N_18973);
and U19047 (N_19047,N_18809,N_18950);
and U19048 (N_19048,N_18875,N_18841);
nand U19049 (N_19049,N_18814,N_18934);
xor U19050 (N_19050,N_18939,N_18852);
nor U19051 (N_19051,N_18850,N_18825);
or U19052 (N_19052,N_18964,N_18823);
nand U19053 (N_19053,N_18869,N_18848);
or U19054 (N_19054,N_18835,N_18836);
xor U19055 (N_19055,N_18827,N_18845);
nor U19056 (N_19056,N_18804,N_18861);
nor U19057 (N_19057,N_18927,N_18886);
and U19058 (N_19058,N_18808,N_18822);
or U19059 (N_19059,N_18930,N_18961);
nor U19060 (N_19060,N_18849,N_18890);
nand U19061 (N_19061,N_18918,N_18829);
nor U19062 (N_19062,N_18855,N_18935);
nor U19063 (N_19063,N_18859,N_18932);
xor U19064 (N_19064,N_18892,N_18944);
and U19065 (N_19065,N_18976,N_18938);
xor U19066 (N_19066,N_18806,N_18905);
xnor U19067 (N_19067,N_18924,N_18975);
and U19068 (N_19068,N_18966,N_18977);
nand U19069 (N_19069,N_18879,N_18847);
nor U19070 (N_19070,N_18802,N_18925);
xor U19071 (N_19071,N_18807,N_18982);
and U19072 (N_19072,N_18902,N_18828);
xnor U19073 (N_19073,N_18818,N_18811);
nor U19074 (N_19074,N_18980,N_18821);
nand U19075 (N_19075,N_18969,N_18922);
nand U19076 (N_19076,N_18824,N_18940);
xor U19077 (N_19077,N_18929,N_18974);
or U19078 (N_19078,N_18894,N_18838);
nand U19079 (N_19079,N_18831,N_18832);
nor U19080 (N_19080,N_18936,N_18933);
xor U19081 (N_19081,N_18900,N_18887);
xnor U19082 (N_19082,N_18962,N_18992);
nand U19083 (N_19083,N_18985,N_18937);
xor U19084 (N_19084,N_18951,N_18856);
and U19085 (N_19085,N_18904,N_18943);
xnor U19086 (N_19086,N_18968,N_18991);
or U19087 (N_19087,N_18999,N_18893);
xnor U19088 (N_19088,N_18953,N_18858);
or U19089 (N_19089,N_18960,N_18817);
and U19090 (N_19090,N_18990,N_18901);
nor U19091 (N_19091,N_18988,N_18812);
xor U19092 (N_19092,N_18866,N_18946);
nor U19093 (N_19093,N_18986,N_18984);
xnor U19094 (N_19094,N_18846,N_18878);
or U19095 (N_19095,N_18872,N_18983);
or U19096 (N_19096,N_18826,N_18942);
xor U19097 (N_19097,N_18979,N_18833);
nor U19098 (N_19098,N_18970,N_18842);
or U19099 (N_19099,N_18995,N_18989);
nand U19100 (N_19100,N_18918,N_18820);
nand U19101 (N_19101,N_18865,N_18995);
nand U19102 (N_19102,N_18969,N_18837);
xor U19103 (N_19103,N_18934,N_18905);
xnor U19104 (N_19104,N_18852,N_18945);
or U19105 (N_19105,N_18888,N_18844);
xnor U19106 (N_19106,N_18812,N_18973);
nor U19107 (N_19107,N_18847,N_18937);
or U19108 (N_19108,N_18951,N_18998);
nand U19109 (N_19109,N_18927,N_18983);
nand U19110 (N_19110,N_18969,N_18903);
or U19111 (N_19111,N_18908,N_18907);
xnor U19112 (N_19112,N_18816,N_18830);
xnor U19113 (N_19113,N_18834,N_18959);
and U19114 (N_19114,N_18815,N_18878);
and U19115 (N_19115,N_18822,N_18850);
and U19116 (N_19116,N_18920,N_18861);
and U19117 (N_19117,N_18834,N_18849);
or U19118 (N_19118,N_18825,N_18938);
nand U19119 (N_19119,N_18989,N_18893);
xor U19120 (N_19120,N_18953,N_18826);
and U19121 (N_19121,N_18929,N_18813);
or U19122 (N_19122,N_18988,N_18887);
xor U19123 (N_19123,N_18905,N_18920);
or U19124 (N_19124,N_18897,N_18844);
and U19125 (N_19125,N_18867,N_18881);
or U19126 (N_19126,N_18818,N_18925);
or U19127 (N_19127,N_18810,N_18959);
nor U19128 (N_19128,N_18835,N_18898);
or U19129 (N_19129,N_18991,N_18940);
nor U19130 (N_19130,N_18924,N_18879);
or U19131 (N_19131,N_18916,N_18935);
xnor U19132 (N_19132,N_18838,N_18978);
xnor U19133 (N_19133,N_18875,N_18868);
or U19134 (N_19134,N_18998,N_18824);
xor U19135 (N_19135,N_18908,N_18986);
and U19136 (N_19136,N_18813,N_18905);
and U19137 (N_19137,N_18871,N_18987);
xor U19138 (N_19138,N_18878,N_18924);
or U19139 (N_19139,N_18810,N_18868);
xor U19140 (N_19140,N_18977,N_18814);
nor U19141 (N_19141,N_18861,N_18896);
nand U19142 (N_19142,N_18940,N_18875);
nand U19143 (N_19143,N_18942,N_18959);
xor U19144 (N_19144,N_18958,N_18836);
xor U19145 (N_19145,N_18955,N_18804);
nor U19146 (N_19146,N_18884,N_18870);
and U19147 (N_19147,N_18970,N_18962);
nand U19148 (N_19148,N_18817,N_18928);
and U19149 (N_19149,N_18910,N_18970);
xnor U19150 (N_19150,N_18907,N_18874);
nand U19151 (N_19151,N_18823,N_18897);
xnor U19152 (N_19152,N_18946,N_18956);
and U19153 (N_19153,N_18949,N_18822);
nand U19154 (N_19154,N_18865,N_18981);
xnor U19155 (N_19155,N_18834,N_18967);
nor U19156 (N_19156,N_18922,N_18847);
nor U19157 (N_19157,N_18875,N_18995);
xnor U19158 (N_19158,N_18824,N_18890);
xor U19159 (N_19159,N_18902,N_18955);
nor U19160 (N_19160,N_18853,N_18953);
or U19161 (N_19161,N_18949,N_18873);
nor U19162 (N_19162,N_18973,N_18928);
nand U19163 (N_19163,N_18860,N_18863);
nand U19164 (N_19164,N_18950,N_18982);
nand U19165 (N_19165,N_18993,N_18926);
nand U19166 (N_19166,N_18800,N_18834);
nand U19167 (N_19167,N_18880,N_18861);
and U19168 (N_19168,N_18880,N_18830);
xor U19169 (N_19169,N_18999,N_18906);
xor U19170 (N_19170,N_18887,N_18984);
nand U19171 (N_19171,N_18874,N_18993);
xnor U19172 (N_19172,N_18873,N_18897);
xnor U19173 (N_19173,N_18839,N_18919);
or U19174 (N_19174,N_18850,N_18900);
and U19175 (N_19175,N_18900,N_18868);
and U19176 (N_19176,N_18964,N_18981);
nor U19177 (N_19177,N_18928,N_18840);
nor U19178 (N_19178,N_18982,N_18812);
nor U19179 (N_19179,N_18893,N_18994);
or U19180 (N_19180,N_18826,N_18938);
and U19181 (N_19181,N_18991,N_18999);
nor U19182 (N_19182,N_18985,N_18892);
nor U19183 (N_19183,N_18977,N_18815);
and U19184 (N_19184,N_18871,N_18826);
xnor U19185 (N_19185,N_18818,N_18861);
or U19186 (N_19186,N_18923,N_18808);
nor U19187 (N_19187,N_18829,N_18908);
xor U19188 (N_19188,N_18885,N_18820);
nor U19189 (N_19189,N_18935,N_18842);
nand U19190 (N_19190,N_18980,N_18951);
and U19191 (N_19191,N_18953,N_18902);
or U19192 (N_19192,N_18908,N_18861);
nor U19193 (N_19193,N_18812,N_18837);
and U19194 (N_19194,N_18940,N_18988);
or U19195 (N_19195,N_18824,N_18974);
nor U19196 (N_19196,N_18814,N_18822);
and U19197 (N_19197,N_18950,N_18900);
nor U19198 (N_19198,N_18872,N_18875);
or U19199 (N_19199,N_18818,N_18942);
or U19200 (N_19200,N_19083,N_19047);
and U19201 (N_19201,N_19077,N_19171);
and U19202 (N_19202,N_19089,N_19036);
nand U19203 (N_19203,N_19199,N_19010);
nor U19204 (N_19204,N_19151,N_19000);
xor U19205 (N_19205,N_19141,N_19155);
nor U19206 (N_19206,N_19197,N_19068);
or U19207 (N_19207,N_19052,N_19118);
nor U19208 (N_19208,N_19086,N_19099);
nand U19209 (N_19209,N_19008,N_19034);
or U19210 (N_19210,N_19075,N_19098);
and U19211 (N_19211,N_19006,N_19056);
and U19212 (N_19212,N_19003,N_19159);
and U19213 (N_19213,N_19101,N_19031);
or U19214 (N_19214,N_19029,N_19169);
and U19215 (N_19215,N_19027,N_19001);
nor U19216 (N_19216,N_19102,N_19125);
nor U19217 (N_19217,N_19119,N_19080);
xor U19218 (N_19218,N_19175,N_19126);
and U19219 (N_19219,N_19134,N_19011);
or U19220 (N_19220,N_19127,N_19040);
or U19221 (N_19221,N_19137,N_19084);
and U19222 (N_19222,N_19092,N_19009);
nand U19223 (N_19223,N_19053,N_19121);
or U19224 (N_19224,N_19024,N_19196);
nor U19225 (N_19225,N_19046,N_19018);
xnor U19226 (N_19226,N_19090,N_19161);
or U19227 (N_19227,N_19050,N_19166);
nor U19228 (N_19228,N_19026,N_19167);
xor U19229 (N_19229,N_19117,N_19035);
or U19230 (N_19230,N_19045,N_19019);
xor U19231 (N_19231,N_19016,N_19174);
nand U19232 (N_19232,N_19022,N_19023);
xnor U19233 (N_19233,N_19032,N_19181);
and U19234 (N_19234,N_19051,N_19191);
xnor U19235 (N_19235,N_19108,N_19184);
or U19236 (N_19236,N_19073,N_19147);
nor U19237 (N_19237,N_19061,N_19177);
nand U19238 (N_19238,N_19195,N_19055);
or U19239 (N_19239,N_19145,N_19064);
and U19240 (N_19240,N_19135,N_19168);
or U19241 (N_19241,N_19105,N_19180);
nand U19242 (N_19242,N_19091,N_19063);
nand U19243 (N_19243,N_19115,N_19002);
and U19244 (N_19244,N_19087,N_19148);
or U19245 (N_19245,N_19107,N_19185);
or U19246 (N_19246,N_19085,N_19094);
nand U19247 (N_19247,N_19097,N_19067);
and U19248 (N_19248,N_19041,N_19049);
xor U19249 (N_19249,N_19198,N_19071);
and U19250 (N_19250,N_19078,N_19178);
or U19251 (N_19251,N_19189,N_19060);
or U19252 (N_19252,N_19039,N_19179);
xnor U19253 (N_19253,N_19143,N_19070);
nor U19254 (N_19254,N_19069,N_19072);
nand U19255 (N_19255,N_19033,N_19110);
and U19256 (N_19256,N_19150,N_19096);
or U19257 (N_19257,N_19088,N_19100);
xnor U19258 (N_19258,N_19025,N_19095);
xor U19259 (N_19259,N_19131,N_19173);
and U19260 (N_19260,N_19038,N_19176);
nor U19261 (N_19261,N_19021,N_19193);
nand U19262 (N_19262,N_19013,N_19048);
and U19263 (N_19263,N_19065,N_19042);
and U19264 (N_19264,N_19183,N_19163);
nand U19265 (N_19265,N_19111,N_19076);
or U19266 (N_19266,N_19170,N_19109);
nand U19267 (N_19267,N_19140,N_19012);
nor U19268 (N_19268,N_19142,N_19136);
and U19269 (N_19269,N_19152,N_19059);
and U19270 (N_19270,N_19160,N_19156);
xnor U19271 (N_19271,N_19112,N_19128);
or U19272 (N_19272,N_19133,N_19165);
xnor U19273 (N_19273,N_19172,N_19004);
xor U19274 (N_19274,N_19062,N_19153);
or U19275 (N_19275,N_19164,N_19120);
or U19276 (N_19276,N_19192,N_19116);
or U19277 (N_19277,N_19058,N_19149);
nand U19278 (N_19278,N_19028,N_19186);
xor U19279 (N_19279,N_19182,N_19030);
nor U19280 (N_19280,N_19015,N_19138);
xnor U19281 (N_19281,N_19093,N_19114);
xor U19282 (N_19282,N_19081,N_19054);
and U19283 (N_19283,N_19158,N_19130);
or U19284 (N_19284,N_19074,N_19113);
and U19285 (N_19285,N_19157,N_19146);
nor U19286 (N_19286,N_19014,N_19017);
xnor U19287 (N_19287,N_19124,N_19154);
or U19288 (N_19288,N_19082,N_19104);
and U19289 (N_19289,N_19187,N_19122);
and U19290 (N_19290,N_19132,N_19194);
and U19291 (N_19291,N_19057,N_19043);
nor U19292 (N_19292,N_19123,N_19188);
nand U19293 (N_19293,N_19037,N_19106);
xnor U19294 (N_19294,N_19162,N_19005);
nand U19295 (N_19295,N_19103,N_19129);
and U19296 (N_19296,N_19139,N_19144);
or U19297 (N_19297,N_19079,N_19190);
or U19298 (N_19298,N_19020,N_19066);
or U19299 (N_19299,N_19044,N_19007);
nand U19300 (N_19300,N_19138,N_19069);
xor U19301 (N_19301,N_19194,N_19010);
xnor U19302 (N_19302,N_19132,N_19037);
and U19303 (N_19303,N_19093,N_19174);
nand U19304 (N_19304,N_19076,N_19087);
nor U19305 (N_19305,N_19006,N_19183);
nand U19306 (N_19306,N_19016,N_19123);
or U19307 (N_19307,N_19093,N_19046);
nor U19308 (N_19308,N_19168,N_19194);
xor U19309 (N_19309,N_19180,N_19070);
and U19310 (N_19310,N_19163,N_19141);
and U19311 (N_19311,N_19147,N_19029);
xnor U19312 (N_19312,N_19065,N_19045);
xnor U19313 (N_19313,N_19130,N_19135);
nor U19314 (N_19314,N_19098,N_19061);
nor U19315 (N_19315,N_19011,N_19185);
and U19316 (N_19316,N_19163,N_19102);
nor U19317 (N_19317,N_19076,N_19133);
nand U19318 (N_19318,N_19071,N_19157);
or U19319 (N_19319,N_19025,N_19188);
nand U19320 (N_19320,N_19119,N_19039);
or U19321 (N_19321,N_19020,N_19179);
and U19322 (N_19322,N_19192,N_19113);
nand U19323 (N_19323,N_19185,N_19127);
nand U19324 (N_19324,N_19035,N_19094);
or U19325 (N_19325,N_19005,N_19076);
or U19326 (N_19326,N_19118,N_19088);
nor U19327 (N_19327,N_19122,N_19088);
xnor U19328 (N_19328,N_19146,N_19138);
nor U19329 (N_19329,N_19197,N_19151);
nand U19330 (N_19330,N_19196,N_19164);
or U19331 (N_19331,N_19170,N_19112);
nor U19332 (N_19332,N_19157,N_19065);
and U19333 (N_19333,N_19020,N_19128);
nand U19334 (N_19334,N_19123,N_19038);
xnor U19335 (N_19335,N_19089,N_19130);
nand U19336 (N_19336,N_19016,N_19012);
or U19337 (N_19337,N_19082,N_19070);
xnor U19338 (N_19338,N_19183,N_19047);
and U19339 (N_19339,N_19047,N_19033);
xor U19340 (N_19340,N_19013,N_19172);
or U19341 (N_19341,N_19189,N_19050);
or U19342 (N_19342,N_19027,N_19117);
nand U19343 (N_19343,N_19176,N_19193);
or U19344 (N_19344,N_19053,N_19168);
nand U19345 (N_19345,N_19145,N_19123);
or U19346 (N_19346,N_19185,N_19027);
and U19347 (N_19347,N_19186,N_19169);
nor U19348 (N_19348,N_19153,N_19139);
xor U19349 (N_19349,N_19036,N_19187);
and U19350 (N_19350,N_19029,N_19033);
xnor U19351 (N_19351,N_19145,N_19172);
nor U19352 (N_19352,N_19122,N_19023);
xnor U19353 (N_19353,N_19105,N_19126);
and U19354 (N_19354,N_19179,N_19038);
nor U19355 (N_19355,N_19189,N_19008);
or U19356 (N_19356,N_19094,N_19083);
nor U19357 (N_19357,N_19186,N_19007);
xor U19358 (N_19358,N_19156,N_19190);
nand U19359 (N_19359,N_19001,N_19148);
or U19360 (N_19360,N_19135,N_19033);
and U19361 (N_19361,N_19123,N_19195);
nor U19362 (N_19362,N_19010,N_19070);
nor U19363 (N_19363,N_19111,N_19100);
or U19364 (N_19364,N_19072,N_19110);
xor U19365 (N_19365,N_19097,N_19021);
nor U19366 (N_19366,N_19128,N_19100);
nor U19367 (N_19367,N_19119,N_19012);
nand U19368 (N_19368,N_19172,N_19132);
xor U19369 (N_19369,N_19148,N_19099);
xnor U19370 (N_19370,N_19123,N_19023);
or U19371 (N_19371,N_19078,N_19087);
nand U19372 (N_19372,N_19137,N_19197);
and U19373 (N_19373,N_19163,N_19085);
nand U19374 (N_19374,N_19158,N_19019);
nand U19375 (N_19375,N_19080,N_19142);
nor U19376 (N_19376,N_19089,N_19066);
or U19377 (N_19377,N_19119,N_19045);
xnor U19378 (N_19378,N_19003,N_19018);
or U19379 (N_19379,N_19174,N_19054);
nor U19380 (N_19380,N_19142,N_19088);
and U19381 (N_19381,N_19112,N_19034);
nor U19382 (N_19382,N_19064,N_19089);
nor U19383 (N_19383,N_19135,N_19026);
and U19384 (N_19384,N_19069,N_19167);
nand U19385 (N_19385,N_19051,N_19049);
or U19386 (N_19386,N_19013,N_19001);
nor U19387 (N_19387,N_19195,N_19115);
and U19388 (N_19388,N_19004,N_19157);
nor U19389 (N_19389,N_19003,N_19188);
and U19390 (N_19390,N_19175,N_19122);
xnor U19391 (N_19391,N_19137,N_19187);
nand U19392 (N_19392,N_19022,N_19141);
nor U19393 (N_19393,N_19168,N_19141);
xor U19394 (N_19394,N_19105,N_19198);
and U19395 (N_19395,N_19152,N_19093);
nand U19396 (N_19396,N_19101,N_19159);
or U19397 (N_19397,N_19025,N_19164);
nand U19398 (N_19398,N_19165,N_19163);
or U19399 (N_19399,N_19002,N_19070);
nand U19400 (N_19400,N_19249,N_19369);
nor U19401 (N_19401,N_19301,N_19384);
nor U19402 (N_19402,N_19397,N_19353);
xnor U19403 (N_19403,N_19268,N_19212);
or U19404 (N_19404,N_19234,N_19213);
or U19405 (N_19405,N_19326,N_19344);
or U19406 (N_19406,N_19224,N_19377);
nand U19407 (N_19407,N_19280,N_19365);
nand U19408 (N_19408,N_19254,N_19395);
or U19409 (N_19409,N_19287,N_19363);
or U19410 (N_19410,N_19229,N_19310);
and U19411 (N_19411,N_19276,N_19385);
nand U19412 (N_19412,N_19255,N_19330);
nor U19413 (N_19413,N_19362,N_19207);
nand U19414 (N_19414,N_19299,N_19282);
xor U19415 (N_19415,N_19317,N_19230);
or U19416 (N_19416,N_19240,N_19336);
nor U19417 (N_19417,N_19259,N_19246);
nor U19418 (N_19418,N_19323,N_19354);
and U19419 (N_19419,N_19297,N_19235);
and U19420 (N_19420,N_19380,N_19352);
nor U19421 (N_19421,N_19300,N_19327);
nor U19422 (N_19422,N_19347,N_19201);
nand U19423 (N_19423,N_19263,N_19269);
or U19424 (N_19424,N_19225,N_19227);
nor U19425 (N_19425,N_19203,N_19298);
or U19426 (N_19426,N_19370,N_19375);
and U19427 (N_19427,N_19284,N_19209);
or U19428 (N_19428,N_19244,N_19231);
xnor U19429 (N_19429,N_19256,N_19245);
nor U19430 (N_19430,N_19305,N_19315);
xor U19431 (N_19431,N_19223,N_19381);
xor U19432 (N_19432,N_19309,N_19366);
xor U19433 (N_19433,N_19260,N_19202);
xnor U19434 (N_19434,N_19343,N_19364);
xnor U19435 (N_19435,N_19393,N_19359);
xor U19436 (N_19436,N_19341,N_19200);
nor U19437 (N_19437,N_19316,N_19220);
or U19438 (N_19438,N_19290,N_19355);
nand U19439 (N_19439,N_19281,N_19337);
xor U19440 (N_19440,N_19348,N_19239);
nand U19441 (N_19441,N_19342,N_19289);
nor U19442 (N_19442,N_19358,N_19295);
nor U19443 (N_19443,N_19304,N_19217);
and U19444 (N_19444,N_19376,N_19206);
nor U19445 (N_19445,N_19367,N_19215);
nand U19446 (N_19446,N_19286,N_19398);
nand U19447 (N_19447,N_19250,N_19332);
and U19448 (N_19448,N_19262,N_19350);
and U19449 (N_19449,N_19266,N_19346);
nand U19450 (N_19450,N_19288,N_19325);
nand U19451 (N_19451,N_19216,N_19324);
nand U19452 (N_19452,N_19253,N_19389);
nor U19453 (N_19453,N_19228,N_19318);
nor U19454 (N_19454,N_19320,N_19351);
and U19455 (N_19455,N_19372,N_19356);
and U19456 (N_19456,N_19222,N_19291);
and U19457 (N_19457,N_19232,N_19241);
or U19458 (N_19458,N_19270,N_19285);
or U19459 (N_19459,N_19329,N_19219);
or U19460 (N_19460,N_19373,N_19283);
nor U19461 (N_19461,N_19391,N_19236);
nor U19462 (N_19462,N_19390,N_19382);
nand U19463 (N_19463,N_19258,N_19328);
and U19464 (N_19464,N_19221,N_19392);
and U19465 (N_19465,N_19378,N_19394);
nor U19466 (N_19466,N_19360,N_19273);
nor U19467 (N_19467,N_19383,N_19248);
and U19468 (N_19468,N_19349,N_19296);
and U19469 (N_19469,N_19226,N_19307);
xor U19470 (N_19470,N_19275,N_19312);
xnor U19471 (N_19471,N_19303,N_19357);
nand U19472 (N_19472,N_19267,N_19274);
or U19473 (N_19473,N_19210,N_19243);
and U19474 (N_19474,N_19321,N_19339);
or U19475 (N_19475,N_19242,N_19251);
and U19476 (N_19476,N_19361,N_19388);
and U19477 (N_19477,N_19264,N_19233);
xor U19478 (N_19478,N_19308,N_19265);
and U19479 (N_19479,N_19257,N_19338);
nand U19480 (N_19480,N_19311,N_19371);
and U19481 (N_19481,N_19319,N_19247);
or U19482 (N_19482,N_19218,N_19334);
nor U19483 (N_19483,N_19374,N_19399);
or U19484 (N_19484,N_19261,N_19306);
and U19485 (N_19485,N_19204,N_19322);
nand U19486 (N_19486,N_19278,N_19293);
and U19487 (N_19487,N_19272,N_19386);
or U19488 (N_19488,N_19279,N_19333);
and U19489 (N_19489,N_19340,N_19292);
nor U19490 (N_19490,N_19335,N_19271);
or U19491 (N_19491,N_19313,N_19205);
nor U19492 (N_19492,N_19294,N_19252);
or U19493 (N_19493,N_19387,N_19277);
or U19494 (N_19494,N_19214,N_19331);
xnor U19495 (N_19495,N_19208,N_19379);
or U19496 (N_19496,N_19314,N_19211);
or U19497 (N_19497,N_19396,N_19345);
and U19498 (N_19498,N_19302,N_19237);
nor U19499 (N_19499,N_19368,N_19238);
or U19500 (N_19500,N_19211,N_19238);
or U19501 (N_19501,N_19282,N_19254);
nand U19502 (N_19502,N_19321,N_19211);
xnor U19503 (N_19503,N_19373,N_19268);
nor U19504 (N_19504,N_19260,N_19220);
and U19505 (N_19505,N_19388,N_19309);
and U19506 (N_19506,N_19269,N_19239);
nor U19507 (N_19507,N_19352,N_19309);
xnor U19508 (N_19508,N_19270,N_19399);
xnor U19509 (N_19509,N_19270,N_19351);
and U19510 (N_19510,N_19366,N_19268);
nand U19511 (N_19511,N_19295,N_19325);
nor U19512 (N_19512,N_19390,N_19263);
nor U19513 (N_19513,N_19363,N_19253);
and U19514 (N_19514,N_19270,N_19274);
nand U19515 (N_19515,N_19269,N_19350);
nand U19516 (N_19516,N_19234,N_19253);
nand U19517 (N_19517,N_19217,N_19250);
or U19518 (N_19518,N_19230,N_19327);
and U19519 (N_19519,N_19312,N_19371);
nor U19520 (N_19520,N_19222,N_19234);
xnor U19521 (N_19521,N_19250,N_19251);
nand U19522 (N_19522,N_19247,N_19236);
or U19523 (N_19523,N_19201,N_19260);
nor U19524 (N_19524,N_19203,N_19283);
xor U19525 (N_19525,N_19326,N_19223);
or U19526 (N_19526,N_19351,N_19357);
or U19527 (N_19527,N_19366,N_19290);
nor U19528 (N_19528,N_19280,N_19200);
xnor U19529 (N_19529,N_19345,N_19312);
and U19530 (N_19530,N_19349,N_19293);
or U19531 (N_19531,N_19386,N_19267);
and U19532 (N_19532,N_19224,N_19353);
or U19533 (N_19533,N_19382,N_19228);
or U19534 (N_19534,N_19299,N_19228);
or U19535 (N_19535,N_19342,N_19224);
nor U19536 (N_19536,N_19333,N_19270);
and U19537 (N_19537,N_19307,N_19250);
nand U19538 (N_19538,N_19241,N_19357);
xor U19539 (N_19539,N_19356,N_19362);
nor U19540 (N_19540,N_19228,N_19317);
and U19541 (N_19541,N_19277,N_19389);
nor U19542 (N_19542,N_19289,N_19311);
and U19543 (N_19543,N_19325,N_19347);
nand U19544 (N_19544,N_19372,N_19328);
xor U19545 (N_19545,N_19349,N_19287);
and U19546 (N_19546,N_19373,N_19232);
nor U19547 (N_19547,N_19285,N_19259);
xnor U19548 (N_19548,N_19336,N_19365);
nor U19549 (N_19549,N_19320,N_19212);
xnor U19550 (N_19550,N_19235,N_19264);
nor U19551 (N_19551,N_19296,N_19283);
or U19552 (N_19552,N_19327,N_19252);
or U19553 (N_19553,N_19214,N_19249);
nor U19554 (N_19554,N_19271,N_19303);
nor U19555 (N_19555,N_19252,N_19395);
nor U19556 (N_19556,N_19318,N_19348);
nor U19557 (N_19557,N_19296,N_19294);
nand U19558 (N_19558,N_19304,N_19201);
xnor U19559 (N_19559,N_19368,N_19366);
xnor U19560 (N_19560,N_19204,N_19309);
xnor U19561 (N_19561,N_19261,N_19273);
nor U19562 (N_19562,N_19239,N_19267);
nand U19563 (N_19563,N_19208,N_19299);
and U19564 (N_19564,N_19354,N_19383);
nand U19565 (N_19565,N_19321,N_19316);
xor U19566 (N_19566,N_19331,N_19221);
nand U19567 (N_19567,N_19346,N_19242);
xnor U19568 (N_19568,N_19258,N_19299);
or U19569 (N_19569,N_19351,N_19300);
and U19570 (N_19570,N_19311,N_19343);
xor U19571 (N_19571,N_19280,N_19390);
and U19572 (N_19572,N_19291,N_19299);
xnor U19573 (N_19573,N_19362,N_19244);
or U19574 (N_19574,N_19244,N_19230);
and U19575 (N_19575,N_19380,N_19360);
xor U19576 (N_19576,N_19347,N_19279);
xor U19577 (N_19577,N_19312,N_19204);
nand U19578 (N_19578,N_19268,N_19271);
nor U19579 (N_19579,N_19354,N_19238);
nor U19580 (N_19580,N_19246,N_19266);
or U19581 (N_19581,N_19397,N_19240);
or U19582 (N_19582,N_19298,N_19333);
nand U19583 (N_19583,N_19338,N_19334);
or U19584 (N_19584,N_19217,N_19393);
nand U19585 (N_19585,N_19390,N_19314);
or U19586 (N_19586,N_19365,N_19369);
nand U19587 (N_19587,N_19308,N_19225);
or U19588 (N_19588,N_19397,N_19248);
and U19589 (N_19589,N_19379,N_19282);
nor U19590 (N_19590,N_19347,N_19348);
and U19591 (N_19591,N_19321,N_19369);
nor U19592 (N_19592,N_19378,N_19290);
xor U19593 (N_19593,N_19336,N_19233);
nand U19594 (N_19594,N_19217,N_19342);
nor U19595 (N_19595,N_19215,N_19293);
nor U19596 (N_19596,N_19384,N_19258);
or U19597 (N_19597,N_19378,N_19240);
or U19598 (N_19598,N_19350,N_19377);
and U19599 (N_19599,N_19304,N_19281);
nand U19600 (N_19600,N_19482,N_19543);
and U19601 (N_19601,N_19437,N_19472);
and U19602 (N_19602,N_19423,N_19486);
and U19603 (N_19603,N_19502,N_19500);
and U19604 (N_19604,N_19456,N_19462);
nand U19605 (N_19605,N_19537,N_19592);
nor U19606 (N_19606,N_19448,N_19480);
and U19607 (N_19607,N_19407,N_19416);
or U19608 (N_19608,N_19470,N_19505);
nor U19609 (N_19609,N_19409,N_19524);
and U19610 (N_19610,N_19517,N_19564);
xor U19611 (N_19611,N_19549,N_19597);
nand U19612 (N_19612,N_19526,N_19501);
and U19613 (N_19613,N_19532,N_19488);
and U19614 (N_19614,N_19552,N_19405);
and U19615 (N_19615,N_19506,N_19417);
nor U19616 (N_19616,N_19463,N_19520);
nor U19617 (N_19617,N_19507,N_19584);
nor U19618 (N_19618,N_19446,N_19447);
or U19619 (N_19619,N_19554,N_19535);
or U19620 (N_19620,N_19550,N_19579);
and U19621 (N_19621,N_19563,N_19578);
or U19622 (N_19622,N_19491,N_19594);
xnor U19623 (N_19623,N_19411,N_19547);
and U19624 (N_19624,N_19586,N_19542);
nand U19625 (N_19625,N_19402,N_19516);
xor U19626 (N_19626,N_19531,N_19565);
xor U19627 (N_19627,N_19573,N_19561);
and U19628 (N_19628,N_19414,N_19460);
and U19629 (N_19629,N_19459,N_19533);
and U19630 (N_19630,N_19498,N_19449);
or U19631 (N_19631,N_19475,N_19465);
xor U19632 (N_19632,N_19540,N_19559);
or U19633 (N_19633,N_19404,N_19548);
and U19634 (N_19634,N_19461,N_19483);
xnor U19635 (N_19635,N_19551,N_19509);
nand U19636 (N_19636,N_19539,N_19494);
and U19637 (N_19637,N_19599,N_19485);
and U19638 (N_19638,N_19588,N_19495);
nand U19639 (N_19639,N_19490,N_19515);
nand U19640 (N_19640,N_19585,N_19435);
xor U19641 (N_19641,N_19439,N_19431);
and U19642 (N_19642,N_19410,N_19541);
and U19643 (N_19643,N_19581,N_19438);
nand U19644 (N_19644,N_19430,N_19511);
and U19645 (N_19645,N_19413,N_19527);
nor U19646 (N_19646,N_19427,N_19534);
nor U19647 (N_19647,N_19576,N_19504);
nand U19648 (N_19648,N_19451,N_19477);
or U19649 (N_19649,N_19412,N_19545);
nand U19650 (N_19650,N_19426,N_19421);
and U19651 (N_19651,N_19583,N_19590);
nor U19652 (N_19652,N_19525,N_19476);
nor U19653 (N_19653,N_19441,N_19445);
nand U19654 (N_19654,N_19418,N_19508);
nor U19655 (N_19655,N_19493,N_19489);
xor U19656 (N_19656,N_19454,N_19466);
xor U19657 (N_19657,N_19521,N_19598);
nand U19658 (N_19658,N_19464,N_19419);
nor U19659 (N_19659,N_19514,N_19450);
xnor U19660 (N_19660,N_19593,N_19513);
or U19661 (N_19661,N_19452,N_19510);
nand U19662 (N_19662,N_19406,N_19569);
nor U19663 (N_19663,N_19503,N_19468);
or U19664 (N_19664,N_19432,N_19492);
nand U19665 (N_19665,N_19415,N_19560);
nand U19666 (N_19666,N_19469,N_19474);
or U19667 (N_19667,N_19487,N_19496);
and U19668 (N_19668,N_19444,N_19455);
xor U19669 (N_19669,N_19436,N_19570);
or U19670 (N_19670,N_19420,N_19555);
nand U19671 (N_19671,N_19473,N_19467);
or U19672 (N_19672,N_19479,N_19442);
nand U19673 (N_19673,N_19589,N_19497);
nand U19674 (N_19674,N_19422,N_19434);
xor U19675 (N_19675,N_19562,N_19566);
or U19676 (N_19676,N_19453,N_19575);
nand U19677 (N_19677,N_19536,N_19425);
nand U19678 (N_19678,N_19458,N_19522);
nand U19679 (N_19679,N_19401,N_19567);
or U19680 (N_19680,N_19553,N_19546);
nand U19681 (N_19681,N_19400,N_19481);
or U19682 (N_19682,N_19528,N_19499);
xnor U19683 (N_19683,N_19557,N_19484);
or U19684 (N_19684,N_19471,N_19478);
xor U19685 (N_19685,N_19424,N_19572);
and U19686 (N_19686,N_19558,N_19591);
or U19687 (N_19687,N_19443,N_19538);
nand U19688 (N_19688,N_19568,N_19433);
xor U19689 (N_19689,N_19582,N_19512);
or U19690 (N_19690,N_19530,N_19518);
xor U19691 (N_19691,N_19596,N_19529);
nand U19692 (N_19692,N_19587,N_19556);
and U19693 (N_19693,N_19544,N_19523);
nand U19694 (N_19694,N_19428,N_19440);
and U19695 (N_19695,N_19457,N_19429);
nor U19696 (N_19696,N_19595,N_19577);
or U19697 (N_19697,N_19574,N_19408);
and U19698 (N_19698,N_19403,N_19571);
nand U19699 (N_19699,N_19580,N_19519);
and U19700 (N_19700,N_19483,N_19505);
and U19701 (N_19701,N_19576,N_19484);
nand U19702 (N_19702,N_19546,N_19403);
xor U19703 (N_19703,N_19523,N_19525);
nand U19704 (N_19704,N_19489,N_19572);
nand U19705 (N_19705,N_19447,N_19592);
nor U19706 (N_19706,N_19548,N_19577);
nand U19707 (N_19707,N_19421,N_19437);
or U19708 (N_19708,N_19412,N_19575);
nor U19709 (N_19709,N_19558,N_19447);
nor U19710 (N_19710,N_19542,N_19529);
or U19711 (N_19711,N_19545,N_19483);
xnor U19712 (N_19712,N_19577,N_19509);
nand U19713 (N_19713,N_19583,N_19481);
or U19714 (N_19714,N_19474,N_19414);
and U19715 (N_19715,N_19508,N_19510);
or U19716 (N_19716,N_19482,N_19484);
nand U19717 (N_19717,N_19594,N_19448);
nor U19718 (N_19718,N_19434,N_19481);
xor U19719 (N_19719,N_19533,N_19401);
nor U19720 (N_19720,N_19408,N_19576);
nor U19721 (N_19721,N_19426,N_19454);
nand U19722 (N_19722,N_19507,N_19423);
and U19723 (N_19723,N_19416,N_19429);
xor U19724 (N_19724,N_19525,N_19457);
nor U19725 (N_19725,N_19445,N_19414);
nor U19726 (N_19726,N_19502,N_19471);
or U19727 (N_19727,N_19596,N_19530);
and U19728 (N_19728,N_19459,N_19549);
nor U19729 (N_19729,N_19422,N_19479);
nand U19730 (N_19730,N_19442,N_19524);
nor U19731 (N_19731,N_19543,N_19584);
or U19732 (N_19732,N_19470,N_19582);
nor U19733 (N_19733,N_19420,N_19529);
or U19734 (N_19734,N_19473,N_19408);
or U19735 (N_19735,N_19561,N_19563);
or U19736 (N_19736,N_19431,N_19539);
or U19737 (N_19737,N_19555,N_19413);
nor U19738 (N_19738,N_19529,N_19481);
or U19739 (N_19739,N_19447,N_19512);
nand U19740 (N_19740,N_19472,N_19447);
nand U19741 (N_19741,N_19584,N_19570);
nand U19742 (N_19742,N_19464,N_19416);
nand U19743 (N_19743,N_19415,N_19516);
nand U19744 (N_19744,N_19556,N_19530);
nand U19745 (N_19745,N_19522,N_19400);
xnor U19746 (N_19746,N_19465,N_19579);
nand U19747 (N_19747,N_19468,N_19480);
nand U19748 (N_19748,N_19445,N_19514);
xor U19749 (N_19749,N_19527,N_19567);
nor U19750 (N_19750,N_19536,N_19573);
xnor U19751 (N_19751,N_19585,N_19541);
nand U19752 (N_19752,N_19482,N_19426);
xor U19753 (N_19753,N_19407,N_19414);
xnor U19754 (N_19754,N_19526,N_19574);
or U19755 (N_19755,N_19464,N_19459);
nor U19756 (N_19756,N_19437,N_19467);
nand U19757 (N_19757,N_19515,N_19465);
nand U19758 (N_19758,N_19467,N_19440);
or U19759 (N_19759,N_19502,N_19533);
or U19760 (N_19760,N_19428,N_19496);
nor U19761 (N_19761,N_19552,N_19445);
nor U19762 (N_19762,N_19426,N_19504);
xnor U19763 (N_19763,N_19407,N_19499);
and U19764 (N_19764,N_19499,N_19491);
and U19765 (N_19765,N_19424,N_19524);
nand U19766 (N_19766,N_19502,N_19413);
xnor U19767 (N_19767,N_19538,N_19581);
or U19768 (N_19768,N_19469,N_19433);
xnor U19769 (N_19769,N_19585,N_19554);
nand U19770 (N_19770,N_19516,N_19419);
nor U19771 (N_19771,N_19421,N_19528);
or U19772 (N_19772,N_19599,N_19426);
nor U19773 (N_19773,N_19460,N_19573);
or U19774 (N_19774,N_19525,N_19417);
nand U19775 (N_19775,N_19407,N_19430);
nand U19776 (N_19776,N_19438,N_19463);
nor U19777 (N_19777,N_19518,N_19480);
xnor U19778 (N_19778,N_19403,N_19428);
nor U19779 (N_19779,N_19532,N_19519);
and U19780 (N_19780,N_19495,N_19570);
nand U19781 (N_19781,N_19539,N_19433);
nand U19782 (N_19782,N_19536,N_19584);
and U19783 (N_19783,N_19468,N_19490);
nor U19784 (N_19784,N_19586,N_19485);
and U19785 (N_19785,N_19465,N_19552);
and U19786 (N_19786,N_19468,N_19564);
and U19787 (N_19787,N_19514,N_19598);
xor U19788 (N_19788,N_19441,N_19571);
xor U19789 (N_19789,N_19513,N_19425);
nand U19790 (N_19790,N_19547,N_19563);
xor U19791 (N_19791,N_19497,N_19556);
or U19792 (N_19792,N_19527,N_19428);
and U19793 (N_19793,N_19462,N_19476);
xnor U19794 (N_19794,N_19452,N_19523);
and U19795 (N_19795,N_19545,N_19498);
nor U19796 (N_19796,N_19470,N_19426);
xnor U19797 (N_19797,N_19477,N_19522);
or U19798 (N_19798,N_19483,N_19531);
nand U19799 (N_19799,N_19476,N_19530);
or U19800 (N_19800,N_19763,N_19748);
or U19801 (N_19801,N_19712,N_19725);
or U19802 (N_19802,N_19630,N_19628);
nand U19803 (N_19803,N_19680,N_19679);
or U19804 (N_19804,N_19684,N_19785);
xnor U19805 (N_19805,N_19726,N_19638);
nand U19806 (N_19806,N_19757,N_19784);
nor U19807 (N_19807,N_19646,N_19603);
and U19808 (N_19808,N_19790,N_19621);
nand U19809 (N_19809,N_19606,N_19731);
and U19810 (N_19810,N_19741,N_19791);
or U19811 (N_19811,N_19775,N_19718);
and U19812 (N_19812,N_19685,N_19764);
and U19813 (N_19813,N_19616,N_19737);
and U19814 (N_19814,N_19602,N_19634);
or U19815 (N_19815,N_19734,N_19736);
or U19816 (N_19816,N_19774,N_19600);
nor U19817 (N_19817,N_19674,N_19691);
xnor U19818 (N_19818,N_19798,N_19742);
xor U19819 (N_19819,N_19717,N_19622);
nor U19820 (N_19820,N_19677,N_19779);
and U19821 (N_19821,N_19673,N_19765);
xnor U19822 (N_19822,N_19728,N_19651);
and U19823 (N_19823,N_19781,N_19727);
or U19824 (N_19824,N_19759,N_19658);
and U19825 (N_19825,N_19796,N_19740);
or U19826 (N_19826,N_19730,N_19705);
and U19827 (N_19827,N_19665,N_19642);
and U19828 (N_19828,N_19693,N_19789);
nor U19829 (N_19829,N_19795,N_19635);
nor U19830 (N_19830,N_19656,N_19702);
xor U19831 (N_19831,N_19743,N_19671);
and U19832 (N_19832,N_19607,N_19697);
or U19833 (N_19833,N_19722,N_19608);
and U19834 (N_19834,N_19624,N_19661);
and U19835 (N_19835,N_19636,N_19681);
xnor U19836 (N_19836,N_19766,N_19675);
xnor U19837 (N_19837,N_19704,N_19772);
or U19838 (N_19838,N_19794,N_19639);
or U19839 (N_19839,N_19601,N_19672);
xnor U19840 (N_19840,N_19650,N_19771);
xor U19841 (N_19841,N_19776,N_19687);
and U19842 (N_19842,N_19778,N_19696);
or U19843 (N_19843,N_19641,N_19719);
nor U19844 (N_19844,N_19611,N_19746);
or U19845 (N_19845,N_19749,N_19793);
or U19846 (N_19846,N_19604,N_19744);
nor U19847 (N_19847,N_19760,N_19733);
or U19848 (N_19848,N_19662,N_19620);
or U19849 (N_19849,N_19762,N_19657);
xnor U19850 (N_19850,N_19666,N_19683);
xor U19851 (N_19851,N_19700,N_19773);
xnor U19852 (N_19852,N_19709,N_19655);
xnor U19853 (N_19853,N_19738,N_19723);
nand U19854 (N_19854,N_19788,N_19669);
xnor U19855 (N_19855,N_19632,N_19627);
or U19856 (N_19856,N_19782,N_19724);
or U19857 (N_19857,N_19714,N_19735);
nand U19858 (N_19858,N_19711,N_19786);
nand U19859 (N_19859,N_19644,N_19755);
nand U19860 (N_19860,N_19613,N_19750);
and U19861 (N_19861,N_19756,N_19645);
or U19862 (N_19862,N_19631,N_19707);
or U19863 (N_19863,N_19694,N_19663);
xor U19864 (N_19864,N_19640,N_19710);
xor U19865 (N_19865,N_19637,N_19626);
nor U19866 (N_19866,N_19695,N_19783);
or U19867 (N_19867,N_19643,N_19769);
nand U19868 (N_19868,N_19689,N_19767);
and U19869 (N_19869,N_19690,N_19761);
or U19870 (N_19870,N_19614,N_19720);
and U19871 (N_19871,N_19701,N_19618);
or U19872 (N_19872,N_19647,N_19653);
nor U19873 (N_19873,N_19660,N_19747);
and U19874 (N_19874,N_19633,N_19792);
xnor U19875 (N_19875,N_19649,N_19623);
nand U19876 (N_19876,N_19768,N_19751);
nor U19877 (N_19877,N_19667,N_19799);
or U19878 (N_19878,N_19698,N_19752);
or U19879 (N_19879,N_19780,N_19617);
and U19880 (N_19880,N_19670,N_19787);
nand U19881 (N_19881,N_19664,N_19703);
nand U19882 (N_19882,N_19699,N_19619);
or U19883 (N_19883,N_19688,N_19654);
xnor U19884 (N_19884,N_19732,N_19713);
or U19885 (N_19885,N_19678,N_19753);
or U19886 (N_19886,N_19629,N_19715);
xnor U19887 (N_19887,N_19605,N_19729);
nand U19888 (N_19888,N_19739,N_19609);
xor U19889 (N_19889,N_19754,N_19615);
xnor U19890 (N_19890,N_19659,N_19758);
nand U19891 (N_19891,N_19610,N_19797);
nand U19892 (N_19892,N_19682,N_19770);
nor U19893 (N_19893,N_19625,N_19706);
and U19894 (N_19894,N_19652,N_19721);
nor U19895 (N_19895,N_19745,N_19668);
nand U19896 (N_19896,N_19648,N_19686);
and U19897 (N_19897,N_19777,N_19612);
nor U19898 (N_19898,N_19692,N_19676);
or U19899 (N_19899,N_19716,N_19708);
xnor U19900 (N_19900,N_19646,N_19692);
nor U19901 (N_19901,N_19685,N_19672);
xnor U19902 (N_19902,N_19714,N_19778);
or U19903 (N_19903,N_19646,N_19627);
nand U19904 (N_19904,N_19602,N_19645);
and U19905 (N_19905,N_19625,N_19634);
nor U19906 (N_19906,N_19670,N_19689);
xor U19907 (N_19907,N_19618,N_19716);
nand U19908 (N_19908,N_19629,N_19649);
or U19909 (N_19909,N_19649,N_19764);
nand U19910 (N_19910,N_19757,N_19683);
nand U19911 (N_19911,N_19790,N_19767);
and U19912 (N_19912,N_19729,N_19742);
and U19913 (N_19913,N_19798,N_19628);
and U19914 (N_19914,N_19732,N_19692);
xnor U19915 (N_19915,N_19737,N_19645);
and U19916 (N_19916,N_19723,N_19654);
nor U19917 (N_19917,N_19709,N_19764);
or U19918 (N_19918,N_19775,N_19607);
and U19919 (N_19919,N_19716,N_19600);
nor U19920 (N_19920,N_19760,N_19670);
or U19921 (N_19921,N_19688,N_19684);
and U19922 (N_19922,N_19785,N_19644);
nor U19923 (N_19923,N_19648,N_19629);
nor U19924 (N_19924,N_19622,N_19691);
xnor U19925 (N_19925,N_19650,N_19764);
nor U19926 (N_19926,N_19701,N_19631);
or U19927 (N_19927,N_19621,N_19669);
nand U19928 (N_19928,N_19733,N_19708);
nand U19929 (N_19929,N_19613,N_19759);
or U19930 (N_19930,N_19796,N_19771);
and U19931 (N_19931,N_19760,N_19618);
or U19932 (N_19932,N_19627,N_19716);
xnor U19933 (N_19933,N_19768,N_19697);
nand U19934 (N_19934,N_19680,N_19714);
and U19935 (N_19935,N_19754,N_19622);
nand U19936 (N_19936,N_19615,N_19717);
and U19937 (N_19937,N_19659,N_19662);
nand U19938 (N_19938,N_19654,N_19731);
and U19939 (N_19939,N_19677,N_19792);
and U19940 (N_19940,N_19699,N_19622);
and U19941 (N_19941,N_19646,N_19656);
nand U19942 (N_19942,N_19735,N_19727);
or U19943 (N_19943,N_19731,N_19701);
nor U19944 (N_19944,N_19725,N_19636);
and U19945 (N_19945,N_19746,N_19629);
and U19946 (N_19946,N_19725,N_19610);
nand U19947 (N_19947,N_19673,N_19777);
xnor U19948 (N_19948,N_19747,N_19686);
xor U19949 (N_19949,N_19798,N_19632);
xor U19950 (N_19950,N_19761,N_19769);
and U19951 (N_19951,N_19783,N_19626);
nand U19952 (N_19952,N_19684,N_19770);
and U19953 (N_19953,N_19688,N_19695);
or U19954 (N_19954,N_19638,N_19640);
or U19955 (N_19955,N_19686,N_19637);
and U19956 (N_19956,N_19608,N_19623);
xor U19957 (N_19957,N_19604,N_19637);
or U19958 (N_19958,N_19680,N_19662);
nand U19959 (N_19959,N_19709,N_19742);
xor U19960 (N_19960,N_19605,N_19685);
and U19961 (N_19961,N_19750,N_19746);
or U19962 (N_19962,N_19768,N_19661);
nor U19963 (N_19963,N_19769,N_19733);
or U19964 (N_19964,N_19780,N_19704);
or U19965 (N_19965,N_19794,N_19795);
and U19966 (N_19966,N_19747,N_19650);
and U19967 (N_19967,N_19673,N_19619);
or U19968 (N_19968,N_19725,N_19608);
xnor U19969 (N_19969,N_19634,N_19682);
xnor U19970 (N_19970,N_19761,N_19619);
nand U19971 (N_19971,N_19734,N_19712);
nand U19972 (N_19972,N_19753,N_19673);
and U19973 (N_19973,N_19656,N_19721);
and U19974 (N_19974,N_19747,N_19685);
nand U19975 (N_19975,N_19699,N_19798);
or U19976 (N_19976,N_19767,N_19647);
nand U19977 (N_19977,N_19717,N_19616);
xnor U19978 (N_19978,N_19671,N_19672);
nand U19979 (N_19979,N_19727,N_19670);
nor U19980 (N_19980,N_19619,N_19781);
nand U19981 (N_19981,N_19725,N_19650);
xor U19982 (N_19982,N_19799,N_19776);
xnor U19983 (N_19983,N_19629,N_19668);
xor U19984 (N_19984,N_19747,N_19600);
and U19985 (N_19985,N_19682,N_19620);
and U19986 (N_19986,N_19684,N_19759);
nor U19987 (N_19987,N_19794,N_19666);
nor U19988 (N_19988,N_19617,N_19651);
and U19989 (N_19989,N_19696,N_19773);
nand U19990 (N_19990,N_19618,N_19666);
nand U19991 (N_19991,N_19644,N_19611);
and U19992 (N_19992,N_19679,N_19619);
or U19993 (N_19993,N_19621,N_19674);
nor U19994 (N_19994,N_19715,N_19740);
xnor U19995 (N_19995,N_19701,N_19660);
and U19996 (N_19996,N_19610,N_19781);
or U19997 (N_19997,N_19724,N_19658);
nor U19998 (N_19998,N_19697,N_19749);
xor U19999 (N_19999,N_19678,N_19659);
nor U20000 (N_20000,N_19901,N_19869);
nor U20001 (N_20001,N_19935,N_19946);
xor U20002 (N_20002,N_19954,N_19964);
nor U20003 (N_20003,N_19864,N_19876);
and U20004 (N_20004,N_19833,N_19915);
nand U20005 (N_20005,N_19846,N_19938);
nor U20006 (N_20006,N_19868,N_19897);
and U20007 (N_20007,N_19815,N_19867);
and U20008 (N_20008,N_19953,N_19894);
nor U20009 (N_20009,N_19863,N_19908);
nand U20010 (N_20010,N_19810,N_19822);
and U20011 (N_20011,N_19959,N_19976);
xnor U20012 (N_20012,N_19984,N_19978);
nand U20013 (N_20013,N_19805,N_19813);
and U20014 (N_20014,N_19830,N_19851);
nand U20015 (N_20015,N_19880,N_19877);
or U20016 (N_20016,N_19930,N_19801);
nor U20017 (N_20017,N_19970,N_19860);
and U20018 (N_20018,N_19961,N_19809);
nand U20019 (N_20019,N_19855,N_19923);
xnor U20020 (N_20020,N_19804,N_19972);
nor U20021 (N_20021,N_19862,N_19837);
or U20022 (N_20022,N_19811,N_19802);
or U20023 (N_20023,N_19937,N_19999);
nand U20024 (N_20024,N_19940,N_19861);
and U20025 (N_20025,N_19920,N_19950);
and U20026 (N_20026,N_19882,N_19866);
nand U20027 (N_20027,N_19878,N_19956);
and U20028 (N_20028,N_19887,N_19952);
nand U20029 (N_20029,N_19884,N_19841);
nor U20030 (N_20030,N_19821,N_19857);
nor U20031 (N_20031,N_19906,N_19893);
or U20032 (N_20032,N_19928,N_19800);
nand U20033 (N_20033,N_19945,N_19913);
nand U20034 (N_20034,N_19816,N_19896);
nor U20035 (N_20035,N_19820,N_19829);
or U20036 (N_20036,N_19844,N_19947);
and U20037 (N_20037,N_19831,N_19995);
nand U20038 (N_20038,N_19842,N_19951);
nand U20039 (N_20039,N_19997,N_19912);
nor U20040 (N_20040,N_19989,N_19990);
and U20041 (N_20041,N_19962,N_19942);
or U20042 (N_20042,N_19807,N_19900);
or U20043 (N_20043,N_19826,N_19949);
or U20044 (N_20044,N_19870,N_19828);
nand U20045 (N_20045,N_19839,N_19981);
xnor U20046 (N_20046,N_19886,N_19873);
or U20047 (N_20047,N_19958,N_19922);
and U20048 (N_20048,N_19819,N_19827);
nand U20049 (N_20049,N_19838,N_19987);
and U20050 (N_20050,N_19992,N_19803);
xor U20051 (N_20051,N_19933,N_19824);
or U20052 (N_20052,N_19968,N_19914);
or U20053 (N_20053,N_19973,N_19926);
and U20054 (N_20054,N_19890,N_19966);
and U20055 (N_20055,N_19874,N_19998);
or U20056 (N_20056,N_19888,N_19818);
or U20057 (N_20057,N_19852,N_19872);
or U20058 (N_20058,N_19932,N_19927);
nand U20059 (N_20059,N_19994,N_19965);
or U20060 (N_20060,N_19895,N_19865);
xor U20061 (N_20061,N_19967,N_19918);
or U20062 (N_20062,N_19911,N_19924);
nor U20063 (N_20063,N_19921,N_19835);
and U20064 (N_20064,N_19849,N_19969);
nand U20065 (N_20065,N_19977,N_19948);
and U20066 (N_20066,N_19892,N_19903);
nand U20067 (N_20067,N_19936,N_19960);
or U20068 (N_20068,N_19891,N_19982);
nor U20069 (N_20069,N_19904,N_19883);
nor U20070 (N_20070,N_19993,N_19850);
nand U20071 (N_20071,N_19910,N_19856);
nand U20072 (N_20072,N_19941,N_19817);
and U20073 (N_20073,N_19843,N_19917);
or U20074 (N_20074,N_19898,N_19929);
and U20075 (N_20075,N_19983,N_19823);
and U20076 (N_20076,N_19979,N_19902);
xnor U20077 (N_20077,N_19985,N_19907);
or U20078 (N_20078,N_19944,N_19939);
or U20079 (N_20079,N_19854,N_19848);
nand U20080 (N_20080,N_19840,N_19834);
or U20081 (N_20081,N_19899,N_19879);
nand U20082 (N_20082,N_19980,N_19875);
nor U20083 (N_20083,N_19847,N_19916);
and U20084 (N_20084,N_19934,N_19957);
and U20085 (N_20085,N_19812,N_19986);
nand U20086 (N_20086,N_19988,N_19974);
and U20087 (N_20087,N_19905,N_19925);
or U20088 (N_20088,N_19808,N_19991);
nand U20089 (N_20089,N_19955,N_19814);
xnor U20090 (N_20090,N_19836,N_19963);
nand U20091 (N_20091,N_19919,N_19885);
xnor U20092 (N_20092,N_19859,N_19871);
xnor U20093 (N_20093,N_19943,N_19996);
and U20094 (N_20094,N_19971,N_19931);
and U20095 (N_20095,N_19858,N_19845);
or U20096 (N_20096,N_19853,N_19975);
or U20097 (N_20097,N_19806,N_19889);
or U20098 (N_20098,N_19832,N_19825);
and U20099 (N_20099,N_19909,N_19881);
or U20100 (N_20100,N_19969,N_19845);
or U20101 (N_20101,N_19951,N_19999);
nand U20102 (N_20102,N_19847,N_19934);
nor U20103 (N_20103,N_19965,N_19887);
nand U20104 (N_20104,N_19992,N_19857);
nand U20105 (N_20105,N_19855,N_19871);
nor U20106 (N_20106,N_19841,N_19839);
nand U20107 (N_20107,N_19804,N_19896);
nand U20108 (N_20108,N_19879,N_19921);
nor U20109 (N_20109,N_19999,N_19952);
nor U20110 (N_20110,N_19981,N_19950);
nor U20111 (N_20111,N_19839,N_19932);
and U20112 (N_20112,N_19912,N_19898);
and U20113 (N_20113,N_19947,N_19915);
nor U20114 (N_20114,N_19929,N_19879);
xnor U20115 (N_20115,N_19983,N_19964);
xnor U20116 (N_20116,N_19953,N_19959);
nand U20117 (N_20117,N_19877,N_19909);
xnor U20118 (N_20118,N_19936,N_19993);
or U20119 (N_20119,N_19914,N_19817);
or U20120 (N_20120,N_19803,N_19826);
nor U20121 (N_20121,N_19854,N_19917);
nor U20122 (N_20122,N_19936,N_19897);
nand U20123 (N_20123,N_19831,N_19936);
nand U20124 (N_20124,N_19819,N_19927);
nand U20125 (N_20125,N_19808,N_19830);
and U20126 (N_20126,N_19860,N_19997);
and U20127 (N_20127,N_19999,N_19867);
or U20128 (N_20128,N_19903,N_19882);
nor U20129 (N_20129,N_19953,N_19835);
nand U20130 (N_20130,N_19848,N_19874);
nand U20131 (N_20131,N_19843,N_19969);
nand U20132 (N_20132,N_19959,N_19956);
nand U20133 (N_20133,N_19866,N_19910);
xnor U20134 (N_20134,N_19879,N_19993);
nor U20135 (N_20135,N_19977,N_19980);
and U20136 (N_20136,N_19988,N_19901);
nor U20137 (N_20137,N_19855,N_19941);
nor U20138 (N_20138,N_19980,N_19931);
and U20139 (N_20139,N_19826,N_19869);
or U20140 (N_20140,N_19920,N_19808);
nor U20141 (N_20141,N_19887,N_19982);
xor U20142 (N_20142,N_19832,N_19952);
and U20143 (N_20143,N_19959,N_19828);
nor U20144 (N_20144,N_19829,N_19987);
and U20145 (N_20145,N_19879,N_19954);
xor U20146 (N_20146,N_19940,N_19871);
or U20147 (N_20147,N_19958,N_19847);
and U20148 (N_20148,N_19935,N_19874);
nand U20149 (N_20149,N_19981,N_19962);
nand U20150 (N_20150,N_19838,N_19823);
nor U20151 (N_20151,N_19942,N_19887);
or U20152 (N_20152,N_19985,N_19820);
nand U20153 (N_20153,N_19941,N_19802);
or U20154 (N_20154,N_19838,N_19898);
nor U20155 (N_20155,N_19927,N_19880);
xor U20156 (N_20156,N_19866,N_19999);
and U20157 (N_20157,N_19865,N_19911);
or U20158 (N_20158,N_19890,N_19881);
and U20159 (N_20159,N_19898,N_19844);
xor U20160 (N_20160,N_19955,N_19938);
nor U20161 (N_20161,N_19917,N_19874);
and U20162 (N_20162,N_19824,N_19954);
nor U20163 (N_20163,N_19917,N_19802);
and U20164 (N_20164,N_19976,N_19971);
nand U20165 (N_20165,N_19877,N_19818);
xnor U20166 (N_20166,N_19946,N_19960);
xor U20167 (N_20167,N_19940,N_19959);
nor U20168 (N_20168,N_19843,N_19982);
or U20169 (N_20169,N_19964,N_19953);
xnor U20170 (N_20170,N_19865,N_19953);
nor U20171 (N_20171,N_19876,N_19814);
xnor U20172 (N_20172,N_19930,N_19926);
nor U20173 (N_20173,N_19973,N_19885);
and U20174 (N_20174,N_19892,N_19834);
or U20175 (N_20175,N_19800,N_19954);
nand U20176 (N_20176,N_19986,N_19834);
nor U20177 (N_20177,N_19915,N_19970);
xnor U20178 (N_20178,N_19924,N_19804);
or U20179 (N_20179,N_19947,N_19964);
nor U20180 (N_20180,N_19877,N_19964);
nor U20181 (N_20181,N_19850,N_19802);
or U20182 (N_20182,N_19804,N_19999);
and U20183 (N_20183,N_19871,N_19901);
nor U20184 (N_20184,N_19862,N_19966);
or U20185 (N_20185,N_19888,N_19977);
xnor U20186 (N_20186,N_19817,N_19901);
and U20187 (N_20187,N_19801,N_19816);
nor U20188 (N_20188,N_19839,N_19984);
nand U20189 (N_20189,N_19868,N_19926);
nand U20190 (N_20190,N_19954,N_19992);
xor U20191 (N_20191,N_19971,N_19986);
nand U20192 (N_20192,N_19847,N_19985);
or U20193 (N_20193,N_19851,N_19964);
or U20194 (N_20194,N_19934,N_19968);
and U20195 (N_20195,N_19890,N_19956);
nor U20196 (N_20196,N_19818,N_19960);
or U20197 (N_20197,N_19801,N_19807);
or U20198 (N_20198,N_19814,N_19806);
nor U20199 (N_20199,N_19889,N_19938);
or U20200 (N_20200,N_20128,N_20048);
nor U20201 (N_20201,N_20065,N_20151);
and U20202 (N_20202,N_20060,N_20080);
and U20203 (N_20203,N_20056,N_20019);
or U20204 (N_20204,N_20091,N_20161);
xor U20205 (N_20205,N_20153,N_20068);
or U20206 (N_20206,N_20147,N_20028);
nor U20207 (N_20207,N_20087,N_20045);
and U20208 (N_20208,N_20088,N_20038);
or U20209 (N_20209,N_20130,N_20111);
or U20210 (N_20210,N_20067,N_20044);
nor U20211 (N_20211,N_20018,N_20109);
nand U20212 (N_20212,N_20084,N_20174);
and U20213 (N_20213,N_20073,N_20057);
and U20214 (N_20214,N_20159,N_20096);
nand U20215 (N_20215,N_20197,N_20094);
nor U20216 (N_20216,N_20034,N_20086);
nand U20217 (N_20217,N_20050,N_20122);
and U20218 (N_20218,N_20104,N_20141);
and U20219 (N_20219,N_20132,N_20119);
and U20220 (N_20220,N_20121,N_20191);
nand U20221 (N_20221,N_20015,N_20185);
nand U20222 (N_20222,N_20009,N_20131);
nor U20223 (N_20223,N_20032,N_20106);
or U20224 (N_20224,N_20033,N_20012);
nand U20225 (N_20225,N_20199,N_20144);
nor U20226 (N_20226,N_20116,N_20102);
nor U20227 (N_20227,N_20095,N_20188);
xor U20228 (N_20228,N_20142,N_20155);
or U20229 (N_20229,N_20016,N_20179);
or U20230 (N_20230,N_20108,N_20154);
nor U20231 (N_20231,N_20007,N_20198);
xor U20232 (N_20232,N_20140,N_20114);
or U20233 (N_20233,N_20182,N_20129);
xor U20234 (N_20234,N_20165,N_20162);
nor U20235 (N_20235,N_20186,N_20052);
and U20236 (N_20236,N_20047,N_20105);
nand U20237 (N_20237,N_20089,N_20011);
and U20238 (N_20238,N_20002,N_20171);
xor U20239 (N_20239,N_20103,N_20049);
xnor U20240 (N_20240,N_20143,N_20134);
nand U20241 (N_20241,N_20146,N_20187);
or U20242 (N_20242,N_20101,N_20027);
and U20243 (N_20243,N_20125,N_20136);
and U20244 (N_20244,N_20195,N_20118);
nor U20245 (N_20245,N_20075,N_20036);
nand U20246 (N_20246,N_20093,N_20078);
nor U20247 (N_20247,N_20099,N_20040);
or U20248 (N_20248,N_20112,N_20123);
nor U20249 (N_20249,N_20006,N_20115);
xnor U20250 (N_20250,N_20022,N_20030);
xnor U20251 (N_20251,N_20062,N_20066);
xor U20252 (N_20252,N_20037,N_20069);
and U20253 (N_20253,N_20063,N_20156);
nand U20254 (N_20254,N_20043,N_20029);
nor U20255 (N_20255,N_20149,N_20074);
xnor U20256 (N_20256,N_20059,N_20085);
or U20257 (N_20257,N_20177,N_20178);
nand U20258 (N_20258,N_20024,N_20124);
xor U20259 (N_20259,N_20127,N_20020);
or U20260 (N_20260,N_20092,N_20023);
nor U20261 (N_20261,N_20003,N_20041);
xor U20262 (N_20262,N_20113,N_20166);
or U20263 (N_20263,N_20017,N_20051);
nor U20264 (N_20264,N_20005,N_20170);
and U20265 (N_20265,N_20175,N_20137);
nand U20266 (N_20266,N_20193,N_20070);
nor U20267 (N_20267,N_20077,N_20039);
xor U20268 (N_20268,N_20054,N_20097);
nand U20269 (N_20269,N_20139,N_20181);
nor U20270 (N_20270,N_20164,N_20035);
or U20271 (N_20271,N_20172,N_20169);
xnor U20272 (N_20272,N_20180,N_20120);
nor U20273 (N_20273,N_20072,N_20163);
nand U20274 (N_20274,N_20173,N_20192);
nor U20275 (N_20275,N_20183,N_20194);
nand U20276 (N_20276,N_20001,N_20190);
nor U20277 (N_20277,N_20098,N_20107);
and U20278 (N_20278,N_20083,N_20079);
or U20279 (N_20279,N_20176,N_20110);
nor U20280 (N_20280,N_20031,N_20013);
and U20281 (N_20281,N_20025,N_20076);
xnor U20282 (N_20282,N_20152,N_20053);
and U20283 (N_20283,N_20010,N_20055);
and U20284 (N_20284,N_20046,N_20081);
and U20285 (N_20285,N_20090,N_20184);
xnor U20286 (N_20286,N_20145,N_20135);
nand U20287 (N_20287,N_20004,N_20138);
nand U20288 (N_20288,N_20014,N_20160);
or U20289 (N_20289,N_20133,N_20117);
nor U20290 (N_20290,N_20071,N_20126);
nand U20291 (N_20291,N_20008,N_20042);
xor U20292 (N_20292,N_20061,N_20021);
nor U20293 (N_20293,N_20158,N_20167);
or U20294 (N_20294,N_20000,N_20100);
nand U20295 (N_20295,N_20157,N_20026);
or U20296 (N_20296,N_20064,N_20196);
or U20297 (N_20297,N_20082,N_20058);
nand U20298 (N_20298,N_20168,N_20189);
and U20299 (N_20299,N_20150,N_20148);
and U20300 (N_20300,N_20167,N_20039);
xor U20301 (N_20301,N_20016,N_20013);
nand U20302 (N_20302,N_20173,N_20001);
nand U20303 (N_20303,N_20038,N_20115);
xor U20304 (N_20304,N_20150,N_20041);
or U20305 (N_20305,N_20074,N_20155);
or U20306 (N_20306,N_20045,N_20033);
xnor U20307 (N_20307,N_20138,N_20055);
nand U20308 (N_20308,N_20030,N_20194);
xnor U20309 (N_20309,N_20025,N_20169);
or U20310 (N_20310,N_20105,N_20146);
and U20311 (N_20311,N_20101,N_20050);
nand U20312 (N_20312,N_20175,N_20006);
and U20313 (N_20313,N_20102,N_20178);
or U20314 (N_20314,N_20140,N_20004);
or U20315 (N_20315,N_20086,N_20159);
nor U20316 (N_20316,N_20043,N_20002);
nand U20317 (N_20317,N_20153,N_20167);
nor U20318 (N_20318,N_20116,N_20032);
nor U20319 (N_20319,N_20032,N_20139);
nand U20320 (N_20320,N_20173,N_20157);
xor U20321 (N_20321,N_20027,N_20059);
nand U20322 (N_20322,N_20103,N_20034);
nor U20323 (N_20323,N_20005,N_20095);
xnor U20324 (N_20324,N_20165,N_20098);
xnor U20325 (N_20325,N_20042,N_20080);
nand U20326 (N_20326,N_20059,N_20129);
nand U20327 (N_20327,N_20002,N_20020);
or U20328 (N_20328,N_20046,N_20047);
xnor U20329 (N_20329,N_20054,N_20189);
nand U20330 (N_20330,N_20030,N_20117);
xnor U20331 (N_20331,N_20170,N_20195);
nand U20332 (N_20332,N_20188,N_20044);
nand U20333 (N_20333,N_20134,N_20071);
nand U20334 (N_20334,N_20114,N_20082);
nand U20335 (N_20335,N_20008,N_20076);
nand U20336 (N_20336,N_20095,N_20148);
or U20337 (N_20337,N_20181,N_20132);
and U20338 (N_20338,N_20105,N_20191);
nor U20339 (N_20339,N_20179,N_20102);
nor U20340 (N_20340,N_20082,N_20052);
nor U20341 (N_20341,N_20110,N_20038);
nor U20342 (N_20342,N_20116,N_20189);
nor U20343 (N_20343,N_20118,N_20184);
nand U20344 (N_20344,N_20108,N_20181);
nor U20345 (N_20345,N_20114,N_20083);
xor U20346 (N_20346,N_20019,N_20017);
nor U20347 (N_20347,N_20183,N_20128);
nand U20348 (N_20348,N_20113,N_20068);
and U20349 (N_20349,N_20107,N_20196);
nand U20350 (N_20350,N_20030,N_20172);
nand U20351 (N_20351,N_20088,N_20108);
nand U20352 (N_20352,N_20132,N_20156);
or U20353 (N_20353,N_20098,N_20144);
nor U20354 (N_20354,N_20066,N_20073);
and U20355 (N_20355,N_20110,N_20167);
nor U20356 (N_20356,N_20060,N_20152);
and U20357 (N_20357,N_20154,N_20181);
or U20358 (N_20358,N_20112,N_20193);
xor U20359 (N_20359,N_20023,N_20136);
nor U20360 (N_20360,N_20025,N_20160);
nor U20361 (N_20361,N_20161,N_20131);
nor U20362 (N_20362,N_20015,N_20122);
nand U20363 (N_20363,N_20050,N_20152);
xnor U20364 (N_20364,N_20191,N_20093);
nor U20365 (N_20365,N_20169,N_20009);
or U20366 (N_20366,N_20083,N_20059);
xor U20367 (N_20367,N_20036,N_20117);
nor U20368 (N_20368,N_20156,N_20076);
nand U20369 (N_20369,N_20113,N_20182);
nand U20370 (N_20370,N_20178,N_20190);
xor U20371 (N_20371,N_20105,N_20167);
nand U20372 (N_20372,N_20010,N_20093);
xnor U20373 (N_20373,N_20008,N_20086);
or U20374 (N_20374,N_20189,N_20132);
or U20375 (N_20375,N_20087,N_20140);
nand U20376 (N_20376,N_20150,N_20053);
nand U20377 (N_20377,N_20158,N_20108);
xnor U20378 (N_20378,N_20041,N_20083);
and U20379 (N_20379,N_20069,N_20012);
xor U20380 (N_20380,N_20053,N_20186);
nor U20381 (N_20381,N_20140,N_20010);
or U20382 (N_20382,N_20014,N_20075);
nor U20383 (N_20383,N_20060,N_20107);
and U20384 (N_20384,N_20072,N_20196);
nand U20385 (N_20385,N_20157,N_20091);
or U20386 (N_20386,N_20161,N_20198);
nand U20387 (N_20387,N_20190,N_20118);
nor U20388 (N_20388,N_20186,N_20090);
xor U20389 (N_20389,N_20134,N_20037);
nor U20390 (N_20390,N_20006,N_20039);
and U20391 (N_20391,N_20091,N_20009);
or U20392 (N_20392,N_20109,N_20144);
xor U20393 (N_20393,N_20045,N_20102);
nand U20394 (N_20394,N_20183,N_20100);
nand U20395 (N_20395,N_20111,N_20025);
nor U20396 (N_20396,N_20000,N_20127);
or U20397 (N_20397,N_20036,N_20141);
nand U20398 (N_20398,N_20082,N_20174);
or U20399 (N_20399,N_20115,N_20194);
xor U20400 (N_20400,N_20209,N_20284);
nand U20401 (N_20401,N_20305,N_20279);
or U20402 (N_20402,N_20310,N_20268);
or U20403 (N_20403,N_20215,N_20345);
or U20404 (N_20404,N_20346,N_20368);
nand U20405 (N_20405,N_20271,N_20285);
nor U20406 (N_20406,N_20396,N_20201);
nand U20407 (N_20407,N_20302,N_20385);
or U20408 (N_20408,N_20233,N_20333);
and U20409 (N_20409,N_20200,N_20249);
nand U20410 (N_20410,N_20252,N_20384);
nand U20411 (N_20411,N_20280,N_20243);
and U20412 (N_20412,N_20321,N_20246);
nand U20413 (N_20413,N_20223,N_20218);
nor U20414 (N_20414,N_20307,N_20267);
nor U20415 (N_20415,N_20324,N_20269);
or U20416 (N_20416,N_20358,N_20287);
or U20417 (N_20417,N_20213,N_20281);
xor U20418 (N_20418,N_20372,N_20343);
and U20419 (N_20419,N_20361,N_20236);
or U20420 (N_20420,N_20290,N_20381);
xor U20421 (N_20421,N_20389,N_20262);
nor U20422 (N_20422,N_20313,N_20292);
nor U20423 (N_20423,N_20210,N_20322);
or U20424 (N_20424,N_20335,N_20317);
nor U20425 (N_20425,N_20234,N_20383);
or U20426 (N_20426,N_20296,N_20391);
nor U20427 (N_20427,N_20352,N_20206);
and U20428 (N_20428,N_20222,N_20349);
nor U20429 (N_20429,N_20247,N_20394);
and U20430 (N_20430,N_20388,N_20202);
nand U20431 (N_20431,N_20339,N_20278);
and U20432 (N_20432,N_20261,N_20363);
nand U20433 (N_20433,N_20379,N_20238);
nand U20434 (N_20434,N_20330,N_20242);
nor U20435 (N_20435,N_20295,N_20211);
or U20436 (N_20436,N_20320,N_20229);
or U20437 (N_20437,N_20277,N_20283);
or U20438 (N_20438,N_20297,N_20289);
or U20439 (N_20439,N_20275,N_20338);
and U20440 (N_20440,N_20364,N_20318);
xnor U20441 (N_20441,N_20212,N_20353);
or U20442 (N_20442,N_20397,N_20378);
nand U20443 (N_20443,N_20235,N_20257);
and U20444 (N_20444,N_20336,N_20365);
or U20445 (N_20445,N_20327,N_20203);
or U20446 (N_20446,N_20393,N_20299);
and U20447 (N_20447,N_20311,N_20226);
and U20448 (N_20448,N_20342,N_20208);
nand U20449 (N_20449,N_20273,N_20354);
nor U20450 (N_20450,N_20237,N_20390);
xor U20451 (N_20451,N_20264,N_20253);
nor U20452 (N_20452,N_20265,N_20293);
xnor U20453 (N_20453,N_20227,N_20228);
or U20454 (N_20454,N_20387,N_20366);
nand U20455 (N_20455,N_20351,N_20348);
nand U20456 (N_20456,N_20308,N_20350);
or U20457 (N_20457,N_20224,N_20325);
or U20458 (N_20458,N_20312,N_20386);
xnor U20459 (N_20459,N_20254,N_20282);
and U20460 (N_20460,N_20377,N_20214);
or U20461 (N_20461,N_20248,N_20326);
nor U20462 (N_20462,N_20306,N_20266);
nand U20463 (N_20463,N_20255,N_20270);
and U20464 (N_20464,N_20276,N_20207);
and U20465 (N_20465,N_20375,N_20300);
nor U20466 (N_20466,N_20328,N_20298);
or U20467 (N_20467,N_20376,N_20360);
nand U20468 (N_20468,N_20225,N_20357);
or U20469 (N_20469,N_20369,N_20316);
or U20470 (N_20470,N_20244,N_20240);
nor U20471 (N_20471,N_20309,N_20371);
or U20472 (N_20472,N_20239,N_20232);
and U20473 (N_20473,N_20251,N_20219);
or U20474 (N_20474,N_20220,N_20221);
xnor U20475 (N_20475,N_20286,N_20245);
nor U20476 (N_20476,N_20337,N_20373);
and U20477 (N_20477,N_20399,N_20341);
and U20478 (N_20478,N_20340,N_20301);
nor U20479 (N_20479,N_20250,N_20260);
and U20480 (N_20480,N_20204,N_20231);
nor U20481 (N_20481,N_20217,N_20334);
nor U20482 (N_20482,N_20374,N_20205);
xnor U20483 (N_20483,N_20329,N_20303);
or U20484 (N_20484,N_20395,N_20323);
nand U20485 (N_20485,N_20332,N_20319);
xor U20486 (N_20486,N_20314,N_20398);
and U20487 (N_20487,N_20382,N_20362);
or U20488 (N_20488,N_20272,N_20291);
nand U20489 (N_20489,N_20230,N_20274);
and U20490 (N_20490,N_20216,N_20347);
nand U20491 (N_20491,N_20356,N_20344);
or U20492 (N_20492,N_20258,N_20331);
nand U20493 (N_20493,N_20294,N_20370);
or U20494 (N_20494,N_20304,N_20256);
and U20495 (N_20495,N_20259,N_20392);
nand U20496 (N_20496,N_20380,N_20315);
xor U20497 (N_20497,N_20241,N_20288);
nor U20498 (N_20498,N_20355,N_20367);
and U20499 (N_20499,N_20263,N_20359);
and U20500 (N_20500,N_20354,N_20234);
and U20501 (N_20501,N_20328,N_20390);
xnor U20502 (N_20502,N_20359,N_20208);
xor U20503 (N_20503,N_20294,N_20313);
xnor U20504 (N_20504,N_20234,N_20254);
and U20505 (N_20505,N_20328,N_20349);
or U20506 (N_20506,N_20356,N_20271);
nand U20507 (N_20507,N_20373,N_20288);
and U20508 (N_20508,N_20283,N_20321);
and U20509 (N_20509,N_20291,N_20233);
and U20510 (N_20510,N_20293,N_20285);
xor U20511 (N_20511,N_20260,N_20259);
nor U20512 (N_20512,N_20324,N_20343);
or U20513 (N_20513,N_20280,N_20300);
nand U20514 (N_20514,N_20213,N_20274);
and U20515 (N_20515,N_20310,N_20326);
nor U20516 (N_20516,N_20368,N_20306);
nand U20517 (N_20517,N_20259,N_20239);
nand U20518 (N_20518,N_20242,N_20296);
and U20519 (N_20519,N_20245,N_20235);
xnor U20520 (N_20520,N_20327,N_20240);
nor U20521 (N_20521,N_20308,N_20312);
nand U20522 (N_20522,N_20238,N_20279);
xor U20523 (N_20523,N_20228,N_20221);
or U20524 (N_20524,N_20332,N_20388);
nor U20525 (N_20525,N_20322,N_20384);
and U20526 (N_20526,N_20393,N_20268);
xnor U20527 (N_20527,N_20392,N_20283);
and U20528 (N_20528,N_20225,N_20267);
nor U20529 (N_20529,N_20276,N_20307);
or U20530 (N_20530,N_20258,N_20234);
and U20531 (N_20531,N_20294,N_20350);
nor U20532 (N_20532,N_20358,N_20370);
xor U20533 (N_20533,N_20377,N_20282);
nor U20534 (N_20534,N_20359,N_20306);
or U20535 (N_20535,N_20337,N_20227);
xnor U20536 (N_20536,N_20292,N_20305);
nand U20537 (N_20537,N_20277,N_20338);
nor U20538 (N_20538,N_20326,N_20330);
nor U20539 (N_20539,N_20312,N_20259);
xor U20540 (N_20540,N_20201,N_20226);
nor U20541 (N_20541,N_20270,N_20338);
xnor U20542 (N_20542,N_20243,N_20389);
nor U20543 (N_20543,N_20320,N_20283);
or U20544 (N_20544,N_20261,N_20337);
nand U20545 (N_20545,N_20201,N_20242);
or U20546 (N_20546,N_20228,N_20256);
and U20547 (N_20547,N_20289,N_20242);
and U20548 (N_20548,N_20332,N_20308);
xnor U20549 (N_20549,N_20359,N_20343);
nor U20550 (N_20550,N_20294,N_20298);
nand U20551 (N_20551,N_20247,N_20234);
xor U20552 (N_20552,N_20239,N_20207);
xor U20553 (N_20553,N_20321,N_20380);
and U20554 (N_20554,N_20280,N_20232);
and U20555 (N_20555,N_20216,N_20286);
or U20556 (N_20556,N_20220,N_20375);
nor U20557 (N_20557,N_20276,N_20340);
or U20558 (N_20558,N_20264,N_20250);
nand U20559 (N_20559,N_20320,N_20215);
nor U20560 (N_20560,N_20319,N_20214);
nor U20561 (N_20561,N_20360,N_20398);
and U20562 (N_20562,N_20363,N_20373);
and U20563 (N_20563,N_20352,N_20309);
and U20564 (N_20564,N_20352,N_20339);
xnor U20565 (N_20565,N_20220,N_20307);
and U20566 (N_20566,N_20221,N_20330);
xnor U20567 (N_20567,N_20312,N_20352);
xor U20568 (N_20568,N_20212,N_20232);
or U20569 (N_20569,N_20307,N_20384);
nand U20570 (N_20570,N_20219,N_20217);
nor U20571 (N_20571,N_20296,N_20270);
and U20572 (N_20572,N_20243,N_20360);
or U20573 (N_20573,N_20240,N_20227);
nor U20574 (N_20574,N_20343,N_20351);
or U20575 (N_20575,N_20301,N_20288);
xnor U20576 (N_20576,N_20203,N_20202);
xnor U20577 (N_20577,N_20385,N_20263);
nand U20578 (N_20578,N_20310,N_20232);
nor U20579 (N_20579,N_20245,N_20239);
or U20580 (N_20580,N_20234,N_20355);
nor U20581 (N_20581,N_20216,N_20240);
or U20582 (N_20582,N_20235,N_20260);
nor U20583 (N_20583,N_20204,N_20322);
nor U20584 (N_20584,N_20314,N_20252);
nand U20585 (N_20585,N_20269,N_20259);
xnor U20586 (N_20586,N_20289,N_20374);
nor U20587 (N_20587,N_20211,N_20398);
and U20588 (N_20588,N_20278,N_20219);
and U20589 (N_20589,N_20228,N_20359);
xnor U20590 (N_20590,N_20352,N_20307);
and U20591 (N_20591,N_20360,N_20346);
xnor U20592 (N_20592,N_20245,N_20277);
nand U20593 (N_20593,N_20373,N_20296);
nor U20594 (N_20594,N_20329,N_20308);
and U20595 (N_20595,N_20216,N_20362);
and U20596 (N_20596,N_20296,N_20210);
nor U20597 (N_20597,N_20250,N_20386);
nor U20598 (N_20598,N_20320,N_20328);
xnor U20599 (N_20599,N_20223,N_20266);
xnor U20600 (N_20600,N_20544,N_20527);
or U20601 (N_20601,N_20449,N_20417);
and U20602 (N_20602,N_20463,N_20507);
and U20603 (N_20603,N_20530,N_20457);
or U20604 (N_20604,N_20427,N_20518);
and U20605 (N_20605,N_20466,N_20418);
nor U20606 (N_20606,N_20487,N_20574);
and U20607 (N_20607,N_20520,N_20425);
and U20608 (N_20608,N_20585,N_20592);
or U20609 (N_20609,N_20563,N_20435);
xnor U20610 (N_20610,N_20571,N_20562);
and U20611 (N_20611,N_20515,N_20479);
and U20612 (N_20612,N_20411,N_20483);
and U20613 (N_20613,N_20413,N_20416);
nand U20614 (N_20614,N_20490,N_20473);
xnor U20615 (N_20615,N_20454,N_20565);
nor U20616 (N_20616,N_20485,N_20489);
or U20617 (N_20617,N_20525,N_20501);
and U20618 (N_20618,N_20465,N_20524);
and U20619 (N_20619,N_20421,N_20533);
nor U20620 (N_20620,N_20475,N_20514);
xor U20621 (N_20621,N_20517,N_20458);
nor U20622 (N_20622,N_20597,N_20498);
or U20623 (N_20623,N_20503,N_20464);
xnor U20624 (N_20624,N_20477,N_20513);
and U20625 (N_20625,N_20570,N_20439);
xnor U20626 (N_20626,N_20596,N_20561);
xnor U20627 (N_20627,N_20535,N_20552);
and U20628 (N_20628,N_20512,N_20493);
and U20629 (N_20629,N_20505,N_20408);
nor U20630 (N_20630,N_20492,N_20547);
xnor U20631 (N_20631,N_20460,N_20419);
nand U20632 (N_20632,N_20495,N_20557);
or U20633 (N_20633,N_20587,N_20566);
or U20634 (N_20634,N_20409,N_20494);
xor U20635 (N_20635,N_20567,N_20484);
nand U20636 (N_20636,N_20516,N_20526);
nand U20637 (N_20637,N_20538,N_20588);
nor U20638 (N_20638,N_20443,N_20590);
nor U20639 (N_20639,N_20448,N_20450);
or U20640 (N_20640,N_20441,N_20482);
and U20641 (N_20641,N_20433,N_20474);
xnor U20642 (N_20642,N_20559,N_20540);
xor U20643 (N_20643,N_20414,N_20444);
and U20644 (N_20644,N_20436,N_20442);
or U20645 (N_20645,N_20400,N_20437);
and U20646 (N_20646,N_20415,N_20446);
or U20647 (N_20647,N_20541,N_20575);
xor U20648 (N_20648,N_20556,N_20598);
xor U20649 (N_20649,N_20583,N_20470);
nor U20650 (N_20650,N_20510,N_20462);
or U20651 (N_20651,N_20573,N_20546);
nor U20652 (N_20652,N_20511,N_20542);
and U20653 (N_20653,N_20496,N_20553);
nand U20654 (N_20654,N_20543,N_20521);
nand U20655 (N_20655,N_20586,N_20432);
nor U20656 (N_20656,N_20407,N_20549);
or U20657 (N_20657,N_20480,N_20534);
and U20658 (N_20658,N_20591,N_20456);
or U20659 (N_20659,N_20429,N_20476);
xnor U20660 (N_20660,N_20582,N_20523);
xnor U20661 (N_20661,N_20595,N_20469);
xor U20662 (N_20662,N_20545,N_20584);
or U20663 (N_20663,N_20434,N_20551);
xor U20664 (N_20664,N_20519,N_20569);
and U20665 (N_20665,N_20593,N_20451);
xor U20666 (N_20666,N_20426,N_20580);
xnor U20667 (N_20667,N_20445,N_20431);
nand U20668 (N_20668,N_20423,N_20478);
and U20669 (N_20669,N_20529,N_20430);
nor U20670 (N_20670,N_20504,N_20481);
xor U20671 (N_20671,N_20536,N_20472);
xnor U20672 (N_20672,N_20412,N_20459);
nand U20673 (N_20673,N_20522,N_20539);
and U20674 (N_20674,N_20420,N_20453);
and U20675 (N_20675,N_20568,N_20554);
xnor U20676 (N_20676,N_20532,N_20558);
nor U20677 (N_20677,N_20405,N_20438);
xnor U20678 (N_20678,N_20447,N_20468);
and U20679 (N_20679,N_20467,N_20422);
nand U20680 (N_20680,N_20572,N_20528);
nor U20681 (N_20681,N_20531,N_20440);
and U20682 (N_20682,N_20577,N_20502);
nor U20683 (N_20683,N_20488,N_20491);
nand U20684 (N_20684,N_20576,N_20508);
nand U20685 (N_20685,N_20424,N_20461);
or U20686 (N_20686,N_20579,N_20410);
or U20687 (N_20687,N_20555,N_20537);
and U20688 (N_20688,N_20499,N_20560);
nor U20689 (N_20689,N_20506,N_20455);
nor U20690 (N_20690,N_20594,N_20403);
and U20691 (N_20691,N_20599,N_20509);
and U20692 (N_20692,N_20548,N_20497);
nor U20693 (N_20693,N_20578,N_20404);
xor U20694 (N_20694,N_20402,N_20500);
nand U20695 (N_20695,N_20406,N_20589);
and U20696 (N_20696,N_20564,N_20471);
and U20697 (N_20697,N_20428,N_20581);
and U20698 (N_20698,N_20401,N_20550);
and U20699 (N_20699,N_20452,N_20486);
and U20700 (N_20700,N_20504,N_20581);
and U20701 (N_20701,N_20417,N_20475);
nand U20702 (N_20702,N_20412,N_20548);
nor U20703 (N_20703,N_20518,N_20524);
xnor U20704 (N_20704,N_20585,N_20406);
nand U20705 (N_20705,N_20523,N_20443);
and U20706 (N_20706,N_20559,N_20447);
and U20707 (N_20707,N_20523,N_20429);
nand U20708 (N_20708,N_20535,N_20442);
or U20709 (N_20709,N_20460,N_20472);
nand U20710 (N_20710,N_20460,N_20440);
xor U20711 (N_20711,N_20427,N_20548);
or U20712 (N_20712,N_20596,N_20420);
nand U20713 (N_20713,N_20440,N_20581);
and U20714 (N_20714,N_20598,N_20480);
nor U20715 (N_20715,N_20440,N_20579);
nand U20716 (N_20716,N_20446,N_20570);
nor U20717 (N_20717,N_20594,N_20413);
and U20718 (N_20718,N_20541,N_20455);
and U20719 (N_20719,N_20540,N_20518);
nor U20720 (N_20720,N_20548,N_20429);
and U20721 (N_20721,N_20583,N_20475);
xor U20722 (N_20722,N_20448,N_20475);
or U20723 (N_20723,N_20598,N_20422);
and U20724 (N_20724,N_20486,N_20408);
or U20725 (N_20725,N_20456,N_20464);
xor U20726 (N_20726,N_20419,N_20414);
or U20727 (N_20727,N_20529,N_20514);
and U20728 (N_20728,N_20465,N_20411);
xor U20729 (N_20729,N_20456,N_20519);
nand U20730 (N_20730,N_20538,N_20542);
and U20731 (N_20731,N_20483,N_20534);
nand U20732 (N_20732,N_20415,N_20577);
nand U20733 (N_20733,N_20447,N_20515);
nand U20734 (N_20734,N_20528,N_20402);
nor U20735 (N_20735,N_20521,N_20414);
nand U20736 (N_20736,N_20463,N_20581);
xnor U20737 (N_20737,N_20580,N_20590);
or U20738 (N_20738,N_20498,N_20453);
or U20739 (N_20739,N_20579,N_20508);
nor U20740 (N_20740,N_20427,N_20496);
or U20741 (N_20741,N_20477,N_20425);
nand U20742 (N_20742,N_20565,N_20486);
xor U20743 (N_20743,N_20591,N_20593);
xor U20744 (N_20744,N_20566,N_20545);
and U20745 (N_20745,N_20598,N_20459);
xor U20746 (N_20746,N_20511,N_20578);
or U20747 (N_20747,N_20509,N_20441);
nand U20748 (N_20748,N_20478,N_20467);
nor U20749 (N_20749,N_20428,N_20540);
xor U20750 (N_20750,N_20510,N_20553);
and U20751 (N_20751,N_20407,N_20541);
nand U20752 (N_20752,N_20443,N_20407);
nand U20753 (N_20753,N_20540,N_20427);
or U20754 (N_20754,N_20405,N_20430);
or U20755 (N_20755,N_20508,N_20433);
or U20756 (N_20756,N_20415,N_20468);
and U20757 (N_20757,N_20569,N_20471);
nor U20758 (N_20758,N_20479,N_20572);
nor U20759 (N_20759,N_20481,N_20499);
nor U20760 (N_20760,N_20503,N_20572);
and U20761 (N_20761,N_20534,N_20407);
xnor U20762 (N_20762,N_20503,N_20437);
or U20763 (N_20763,N_20473,N_20430);
nand U20764 (N_20764,N_20587,N_20538);
and U20765 (N_20765,N_20561,N_20473);
xor U20766 (N_20766,N_20528,N_20563);
nand U20767 (N_20767,N_20457,N_20449);
or U20768 (N_20768,N_20437,N_20424);
and U20769 (N_20769,N_20473,N_20581);
nand U20770 (N_20770,N_20434,N_20504);
nand U20771 (N_20771,N_20479,N_20489);
and U20772 (N_20772,N_20568,N_20523);
nand U20773 (N_20773,N_20571,N_20536);
or U20774 (N_20774,N_20544,N_20487);
xor U20775 (N_20775,N_20439,N_20484);
or U20776 (N_20776,N_20420,N_20586);
xnor U20777 (N_20777,N_20478,N_20598);
and U20778 (N_20778,N_20517,N_20547);
nand U20779 (N_20779,N_20539,N_20537);
or U20780 (N_20780,N_20427,N_20400);
or U20781 (N_20781,N_20428,N_20458);
nand U20782 (N_20782,N_20576,N_20581);
or U20783 (N_20783,N_20535,N_20549);
xnor U20784 (N_20784,N_20426,N_20449);
xor U20785 (N_20785,N_20599,N_20430);
and U20786 (N_20786,N_20508,N_20525);
or U20787 (N_20787,N_20414,N_20464);
nor U20788 (N_20788,N_20595,N_20409);
xnor U20789 (N_20789,N_20500,N_20555);
or U20790 (N_20790,N_20479,N_20503);
or U20791 (N_20791,N_20573,N_20464);
xnor U20792 (N_20792,N_20581,N_20590);
nor U20793 (N_20793,N_20598,N_20574);
and U20794 (N_20794,N_20458,N_20451);
nor U20795 (N_20795,N_20504,N_20402);
nor U20796 (N_20796,N_20523,N_20434);
nor U20797 (N_20797,N_20458,N_20447);
nand U20798 (N_20798,N_20401,N_20442);
nor U20799 (N_20799,N_20444,N_20579);
nand U20800 (N_20800,N_20790,N_20615);
and U20801 (N_20801,N_20784,N_20728);
xor U20802 (N_20802,N_20672,N_20717);
or U20803 (N_20803,N_20750,N_20791);
or U20804 (N_20804,N_20629,N_20666);
and U20805 (N_20805,N_20754,N_20739);
xnor U20806 (N_20806,N_20619,N_20676);
and U20807 (N_20807,N_20718,N_20731);
or U20808 (N_20808,N_20742,N_20639);
or U20809 (N_20809,N_20767,N_20755);
or U20810 (N_20810,N_20668,N_20797);
and U20811 (N_20811,N_20609,N_20626);
or U20812 (N_20812,N_20643,N_20765);
and U20813 (N_20813,N_20727,N_20770);
or U20814 (N_20814,N_20627,N_20617);
and U20815 (N_20815,N_20624,N_20723);
or U20816 (N_20816,N_20748,N_20611);
nand U20817 (N_20817,N_20692,N_20669);
and U20818 (N_20818,N_20777,N_20735);
or U20819 (N_20819,N_20684,N_20712);
or U20820 (N_20820,N_20786,N_20794);
nor U20821 (N_20821,N_20635,N_20788);
and U20822 (N_20822,N_20760,N_20690);
nand U20823 (N_20823,N_20715,N_20657);
nand U20824 (N_20824,N_20787,N_20764);
or U20825 (N_20825,N_20673,N_20753);
xnor U20826 (N_20826,N_20688,N_20710);
xnor U20827 (N_20827,N_20707,N_20689);
nand U20828 (N_20828,N_20756,N_20714);
xor U20829 (N_20829,N_20693,N_20785);
xor U20830 (N_20830,N_20660,N_20655);
or U20831 (N_20831,N_20651,N_20771);
and U20832 (N_20832,N_20780,N_20618);
or U20833 (N_20833,N_20706,N_20621);
or U20834 (N_20834,N_20730,N_20773);
nand U20835 (N_20835,N_20661,N_20766);
xor U20836 (N_20836,N_20695,N_20628);
or U20837 (N_20837,N_20600,N_20604);
xnor U20838 (N_20838,N_20736,N_20782);
nor U20839 (N_20839,N_20696,N_20740);
nand U20840 (N_20840,N_20682,N_20607);
nand U20841 (N_20841,N_20670,N_20758);
or U20842 (N_20842,N_20795,N_20783);
or U20843 (N_20843,N_20711,N_20603);
nand U20844 (N_20844,N_20798,N_20649);
or U20845 (N_20845,N_20648,N_20664);
nor U20846 (N_20846,N_20637,N_20776);
nand U20847 (N_20847,N_20665,N_20700);
or U20848 (N_20848,N_20761,N_20671);
nor U20849 (N_20849,N_20719,N_20614);
nor U20850 (N_20850,N_20602,N_20779);
xnor U20851 (N_20851,N_20792,N_20733);
and U20852 (N_20852,N_20633,N_20701);
nand U20853 (N_20853,N_20658,N_20720);
nor U20854 (N_20854,N_20738,N_20694);
nor U20855 (N_20855,N_20737,N_20702);
nand U20856 (N_20856,N_20726,N_20622);
or U20857 (N_20857,N_20679,N_20747);
nand U20858 (N_20858,N_20732,N_20749);
or U20859 (N_20859,N_20653,N_20613);
nand U20860 (N_20860,N_20608,N_20685);
and U20861 (N_20861,N_20646,N_20691);
nand U20862 (N_20862,N_20631,N_20751);
and U20863 (N_20863,N_20610,N_20743);
xnor U20864 (N_20864,N_20687,N_20667);
nand U20865 (N_20865,N_20699,N_20636);
or U20866 (N_20866,N_20678,N_20762);
nor U20867 (N_20867,N_20708,N_20725);
nor U20868 (N_20868,N_20796,N_20674);
or U20869 (N_20869,N_20663,N_20675);
nor U20870 (N_20870,N_20680,N_20704);
or U20871 (N_20871,N_20752,N_20721);
xnor U20872 (N_20872,N_20645,N_20641);
xnor U20873 (N_20873,N_20775,N_20642);
or U20874 (N_20874,N_20763,N_20662);
nand U20875 (N_20875,N_20774,N_20757);
and U20876 (N_20876,N_20625,N_20605);
nand U20877 (N_20877,N_20656,N_20746);
xor U20878 (N_20878,N_20620,N_20745);
nand U20879 (N_20879,N_20713,N_20647);
and U20880 (N_20880,N_20778,N_20799);
nor U20881 (N_20881,N_20781,N_20722);
nand U20882 (N_20882,N_20640,N_20729);
nand U20883 (N_20883,N_20634,N_20734);
or U20884 (N_20884,N_20654,N_20741);
and U20885 (N_20885,N_20652,N_20759);
nor U20886 (N_20886,N_20697,N_20724);
and U20887 (N_20887,N_20716,N_20703);
and U20888 (N_20888,N_20612,N_20644);
and U20889 (N_20889,N_20630,N_20769);
or U20890 (N_20890,N_20686,N_20681);
nor U20891 (N_20891,N_20650,N_20632);
nor U20892 (N_20892,N_20793,N_20638);
nor U20893 (N_20893,N_20772,N_20601);
nand U20894 (N_20894,N_20683,N_20606);
nor U20895 (N_20895,N_20677,N_20789);
nand U20896 (N_20896,N_20744,N_20659);
nor U20897 (N_20897,N_20709,N_20616);
nor U20898 (N_20898,N_20768,N_20623);
xor U20899 (N_20899,N_20698,N_20705);
or U20900 (N_20900,N_20762,N_20679);
xor U20901 (N_20901,N_20764,N_20782);
or U20902 (N_20902,N_20630,N_20779);
nand U20903 (N_20903,N_20627,N_20659);
xnor U20904 (N_20904,N_20768,N_20639);
xnor U20905 (N_20905,N_20683,N_20739);
or U20906 (N_20906,N_20766,N_20640);
or U20907 (N_20907,N_20766,N_20659);
and U20908 (N_20908,N_20772,N_20666);
nor U20909 (N_20909,N_20627,N_20691);
nand U20910 (N_20910,N_20692,N_20758);
or U20911 (N_20911,N_20639,N_20687);
and U20912 (N_20912,N_20663,N_20790);
and U20913 (N_20913,N_20691,N_20668);
and U20914 (N_20914,N_20770,N_20719);
and U20915 (N_20915,N_20720,N_20637);
nand U20916 (N_20916,N_20749,N_20629);
xor U20917 (N_20917,N_20788,N_20726);
nand U20918 (N_20918,N_20653,N_20618);
or U20919 (N_20919,N_20714,N_20672);
nor U20920 (N_20920,N_20762,N_20690);
nor U20921 (N_20921,N_20612,N_20708);
and U20922 (N_20922,N_20618,N_20654);
nor U20923 (N_20923,N_20792,N_20672);
nor U20924 (N_20924,N_20649,N_20797);
nor U20925 (N_20925,N_20781,N_20634);
nor U20926 (N_20926,N_20673,N_20617);
nand U20927 (N_20927,N_20784,N_20766);
xnor U20928 (N_20928,N_20620,N_20621);
xnor U20929 (N_20929,N_20763,N_20731);
and U20930 (N_20930,N_20625,N_20720);
nor U20931 (N_20931,N_20646,N_20676);
xnor U20932 (N_20932,N_20603,N_20714);
xor U20933 (N_20933,N_20741,N_20653);
xnor U20934 (N_20934,N_20799,N_20789);
nor U20935 (N_20935,N_20674,N_20777);
nand U20936 (N_20936,N_20612,N_20762);
and U20937 (N_20937,N_20777,N_20718);
nand U20938 (N_20938,N_20625,N_20614);
nand U20939 (N_20939,N_20661,N_20782);
and U20940 (N_20940,N_20705,N_20709);
xnor U20941 (N_20941,N_20796,N_20777);
and U20942 (N_20942,N_20681,N_20710);
xor U20943 (N_20943,N_20601,N_20623);
and U20944 (N_20944,N_20694,N_20672);
xnor U20945 (N_20945,N_20791,N_20620);
xnor U20946 (N_20946,N_20722,N_20732);
xnor U20947 (N_20947,N_20761,N_20632);
and U20948 (N_20948,N_20733,N_20662);
xor U20949 (N_20949,N_20684,N_20659);
or U20950 (N_20950,N_20642,N_20610);
or U20951 (N_20951,N_20758,N_20744);
nand U20952 (N_20952,N_20700,N_20612);
or U20953 (N_20953,N_20784,N_20714);
nand U20954 (N_20954,N_20707,N_20624);
nand U20955 (N_20955,N_20619,N_20783);
xor U20956 (N_20956,N_20663,N_20635);
xnor U20957 (N_20957,N_20602,N_20730);
or U20958 (N_20958,N_20677,N_20738);
xnor U20959 (N_20959,N_20646,N_20689);
nor U20960 (N_20960,N_20687,N_20701);
and U20961 (N_20961,N_20635,N_20763);
or U20962 (N_20962,N_20717,N_20766);
or U20963 (N_20963,N_20747,N_20741);
or U20964 (N_20964,N_20734,N_20674);
nand U20965 (N_20965,N_20790,N_20709);
nand U20966 (N_20966,N_20724,N_20763);
nor U20967 (N_20967,N_20737,N_20704);
xnor U20968 (N_20968,N_20668,N_20603);
xnor U20969 (N_20969,N_20739,N_20603);
nor U20970 (N_20970,N_20662,N_20794);
nand U20971 (N_20971,N_20704,N_20688);
xor U20972 (N_20972,N_20603,N_20637);
nand U20973 (N_20973,N_20605,N_20724);
nand U20974 (N_20974,N_20653,N_20754);
xnor U20975 (N_20975,N_20787,N_20645);
nor U20976 (N_20976,N_20752,N_20716);
and U20977 (N_20977,N_20796,N_20665);
or U20978 (N_20978,N_20771,N_20752);
or U20979 (N_20979,N_20723,N_20716);
or U20980 (N_20980,N_20727,N_20746);
nor U20981 (N_20981,N_20608,N_20734);
nor U20982 (N_20982,N_20615,N_20656);
and U20983 (N_20983,N_20793,N_20786);
nand U20984 (N_20984,N_20754,N_20688);
or U20985 (N_20985,N_20710,N_20620);
and U20986 (N_20986,N_20743,N_20785);
or U20987 (N_20987,N_20694,N_20755);
nand U20988 (N_20988,N_20781,N_20791);
or U20989 (N_20989,N_20721,N_20628);
and U20990 (N_20990,N_20675,N_20727);
xnor U20991 (N_20991,N_20690,N_20651);
and U20992 (N_20992,N_20716,N_20666);
or U20993 (N_20993,N_20764,N_20664);
or U20994 (N_20994,N_20670,N_20608);
nand U20995 (N_20995,N_20635,N_20784);
nor U20996 (N_20996,N_20635,N_20733);
nand U20997 (N_20997,N_20799,N_20755);
xor U20998 (N_20998,N_20671,N_20603);
and U20999 (N_20999,N_20699,N_20655);
or U21000 (N_21000,N_20976,N_20924);
nand U21001 (N_21001,N_20847,N_20809);
or U21002 (N_21002,N_20882,N_20985);
nand U21003 (N_21003,N_20867,N_20932);
nor U21004 (N_21004,N_20906,N_20897);
or U21005 (N_21005,N_20835,N_20859);
nor U21006 (N_21006,N_20977,N_20903);
and U21007 (N_21007,N_20834,N_20826);
nand U21008 (N_21008,N_20990,N_20822);
nor U21009 (N_21009,N_20804,N_20857);
nand U21010 (N_21010,N_20896,N_20808);
nand U21011 (N_21011,N_20872,N_20862);
nand U21012 (N_21012,N_20814,N_20930);
or U21013 (N_21013,N_20860,N_20806);
or U21014 (N_21014,N_20838,N_20979);
nor U21015 (N_21015,N_20908,N_20858);
nor U21016 (N_21016,N_20950,N_20933);
nor U21017 (N_21017,N_20855,N_20900);
and U21018 (N_21018,N_20807,N_20892);
and U21019 (N_21019,N_20907,N_20958);
nor U21020 (N_21020,N_20815,N_20854);
or U21021 (N_21021,N_20851,N_20883);
and U21022 (N_21022,N_20888,N_20849);
xor U21023 (N_21023,N_20839,N_20841);
or U21024 (N_21024,N_20966,N_20880);
and U21025 (N_21025,N_20845,N_20821);
or U21026 (N_21026,N_20902,N_20866);
nor U21027 (N_21027,N_20819,N_20960);
nor U21028 (N_21028,N_20813,N_20800);
nor U21029 (N_21029,N_20968,N_20949);
nor U21030 (N_21030,N_20864,N_20991);
and U21031 (N_21031,N_20853,N_20827);
and U21032 (N_21032,N_20962,N_20861);
nand U21033 (N_21033,N_20925,N_20947);
xnor U21034 (N_21034,N_20890,N_20928);
xnor U21035 (N_21035,N_20891,N_20901);
nor U21036 (N_21036,N_20831,N_20940);
xnor U21037 (N_21037,N_20915,N_20944);
nor U21038 (N_21038,N_20879,N_20911);
and U21039 (N_21039,N_20934,N_20913);
or U21040 (N_21040,N_20869,N_20811);
nand U21041 (N_21041,N_20801,N_20810);
xnor U21042 (N_21042,N_20941,N_20923);
xnor U21043 (N_21043,N_20812,N_20983);
and U21044 (N_21044,N_20887,N_20978);
nor U21045 (N_21045,N_20886,N_20836);
and U21046 (N_21046,N_20863,N_20927);
and U21047 (N_21047,N_20936,N_20984);
or U21048 (N_21048,N_20829,N_20889);
and U21049 (N_21049,N_20999,N_20969);
xnor U21050 (N_21050,N_20994,N_20917);
and U21051 (N_21051,N_20973,N_20850);
nor U21052 (N_21052,N_20955,N_20824);
nor U21053 (N_21053,N_20848,N_20895);
nor U21054 (N_21054,N_20825,N_20942);
or U21055 (N_21055,N_20884,N_20993);
xor U21056 (N_21056,N_20982,N_20894);
or U21057 (N_21057,N_20943,N_20856);
nand U21058 (N_21058,N_20989,N_20997);
nand U21059 (N_21059,N_20840,N_20914);
xor U21060 (N_21060,N_20877,N_20967);
and U21061 (N_21061,N_20921,N_20878);
and U21062 (N_21062,N_20904,N_20951);
xor U21063 (N_21063,N_20975,N_20843);
xnor U21064 (N_21064,N_20885,N_20912);
xnor U21065 (N_21065,N_20893,N_20931);
or U21066 (N_21066,N_20956,N_20980);
nand U21067 (N_21067,N_20935,N_20981);
xnor U21068 (N_21068,N_20948,N_20963);
xor U21069 (N_21069,N_20874,N_20996);
nand U21070 (N_21070,N_20922,N_20803);
and U21071 (N_21071,N_20916,N_20972);
nand U21072 (N_21072,N_20986,N_20920);
and U21073 (N_21073,N_20926,N_20817);
nand U21074 (N_21074,N_20871,N_20876);
or U21075 (N_21075,N_20909,N_20828);
xnor U21076 (N_21076,N_20961,N_20953);
nor U21077 (N_21077,N_20905,N_20959);
nand U21078 (N_21078,N_20820,N_20974);
nor U21079 (N_21079,N_20918,N_20805);
nor U21080 (N_21080,N_20873,N_20898);
nor U21081 (N_21081,N_20833,N_20998);
or U21082 (N_21082,N_20992,N_20939);
and U21083 (N_21083,N_20945,N_20837);
nor U21084 (N_21084,N_20881,N_20946);
nand U21085 (N_21085,N_20842,N_20995);
or U21086 (N_21086,N_20964,N_20987);
xnor U21087 (N_21087,N_20988,N_20938);
or U21088 (N_21088,N_20830,N_20954);
nand U21089 (N_21089,N_20957,N_20899);
or U21090 (N_21090,N_20919,N_20823);
xor U21091 (N_21091,N_20852,N_20816);
and U21092 (N_21092,N_20965,N_20870);
nor U21093 (N_21093,N_20929,N_20868);
and U21094 (N_21094,N_20865,N_20844);
or U21095 (N_21095,N_20818,N_20832);
nand U21096 (N_21096,N_20875,N_20910);
and U21097 (N_21097,N_20970,N_20952);
xor U21098 (N_21098,N_20802,N_20971);
or U21099 (N_21099,N_20846,N_20937);
or U21100 (N_21100,N_20940,N_20934);
nand U21101 (N_21101,N_20981,N_20941);
nor U21102 (N_21102,N_20949,N_20940);
nor U21103 (N_21103,N_20954,N_20803);
nand U21104 (N_21104,N_20850,N_20805);
nor U21105 (N_21105,N_20887,N_20815);
nand U21106 (N_21106,N_20836,N_20970);
nand U21107 (N_21107,N_20952,N_20871);
xnor U21108 (N_21108,N_20877,N_20894);
or U21109 (N_21109,N_20819,N_20840);
nand U21110 (N_21110,N_20883,N_20903);
and U21111 (N_21111,N_20962,N_20991);
xnor U21112 (N_21112,N_20974,N_20986);
xnor U21113 (N_21113,N_20827,N_20890);
nand U21114 (N_21114,N_20967,N_20911);
or U21115 (N_21115,N_20889,N_20932);
nor U21116 (N_21116,N_20920,N_20973);
or U21117 (N_21117,N_20920,N_20911);
xnor U21118 (N_21118,N_20857,N_20993);
nand U21119 (N_21119,N_20943,N_20892);
or U21120 (N_21120,N_20894,N_20804);
nand U21121 (N_21121,N_20891,N_20897);
xnor U21122 (N_21122,N_20815,N_20940);
and U21123 (N_21123,N_20864,N_20895);
or U21124 (N_21124,N_20894,N_20913);
nor U21125 (N_21125,N_20954,N_20891);
or U21126 (N_21126,N_20989,N_20880);
nor U21127 (N_21127,N_20918,N_20838);
and U21128 (N_21128,N_20820,N_20905);
and U21129 (N_21129,N_20848,N_20925);
or U21130 (N_21130,N_20954,N_20883);
nand U21131 (N_21131,N_20815,N_20802);
and U21132 (N_21132,N_20936,N_20983);
xor U21133 (N_21133,N_20938,N_20839);
nor U21134 (N_21134,N_20958,N_20838);
xnor U21135 (N_21135,N_20891,N_20889);
nor U21136 (N_21136,N_20831,N_20913);
nand U21137 (N_21137,N_20948,N_20801);
nor U21138 (N_21138,N_20888,N_20880);
or U21139 (N_21139,N_20811,N_20961);
or U21140 (N_21140,N_20995,N_20893);
xnor U21141 (N_21141,N_20957,N_20997);
nand U21142 (N_21142,N_20919,N_20829);
nand U21143 (N_21143,N_20963,N_20830);
xnor U21144 (N_21144,N_20922,N_20875);
and U21145 (N_21145,N_20825,N_20800);
nor U21146 (N_21146,N_20896,N_20853);
xor U21147 (N_21147,N_20820,N_20977);
xnor U21148 (N_21148,N_20856,N_20854);
and U21149 (N_21149,N_20915,N_20927);
or U21150 (N_21150,N_20814,N_20903);
nand U21151 (N_21151,N_20894,N_20814);
nand U21152 (N_21152,N_20836,N_20863);
and U21153 (N_21153,N_20817,N_20935);
nor U21154 (N_21154,N_20835,N_20949);
or U21155 (N_21155,N_20999,N_20907);
nand U21156 (N_21156,N_20882,N_20858);
xor U21157 (N_21157,N_20846,N_20815);
nand U21158 (N_21158,N_20900,N_20965);
or U21159 (N_21159,N_20995,N_20908);
or U21160 (N_21160,N_20954,N_20852);
or U21161 (N_21161,N_20856,N_20953);
and U21162 (N_21162,N_20923,N_20966);
and U21163 (N_21163,N_20862,N_20937);
and U21164 (N_21164,N_20880,N_20907);
or U21165 (N_21165,N_20948,N_20864);
or U21166 (N_21166,N_20850,N_20833);
nand U21167 (N_21167,N_20847,N_20880);
xnor U21168 (N_21168,N_20916,N_20800);
nand U21169 (N_21169,N_20902,N_20868);
xor U21170 (N_21170,N_20952,N_20879);
nand U21171 (N_21171,N_20890,N_20957);
nand U21172 (N_21172,N_20988,N_20939);
or U21173 (N_21173,N_20989,N_20969);
or U21174 (N_21174,N_20962,N_20891);
and U21175 (N_21175,N_20965,N_20850);
xor U21176 (N_21176,N_20810,N_20925);
nor U21177 (N_21177,N_20811,N_20989);
nor U21178 (N_21178,N_20966,N_20982);
nor U21179 (N_21179,N_20905,N_20876);
xnor U21180 (N_21180,N_20837,N_20950);
xnor U21181 (N_21181,N_20951,N_20898);
and U21182 (N_21182,N_20817,N_20979);
or U21183 (N_21183,N_20895,N_20906);
and U21184 (N_21184,N_20832,N_20897);
or U21185 (N_21185,N_20982,N_20944);
nor U21186 (N_21186,N_20909,N_20905);
xor U21187 (N_21187,N_20839,N_20871);
and U21188 (N_21188,N_20861,N_20833);
nand U21189 (N_21189,N_20959,N_20886);
xnor U21190 (N_21190,N_20992,N_20867);
and U21191 (N_21191,N_20895,N_20999);
nand U21192 (N_21192,N_20919,N_20915);
nor U21193 (N_21193,N_20822,N_20866);
nor U21194 (N_21194,N_20950,N_20971);
xor U21195 (N_21195,N_20861,N_20913);
nand U21196 (N_21196,N_20904,N_20988);
and U21197 (N_21197,N_20814,N_20851);
xnor U21198 (N_21198,N_20948,N_20953);
nor U21199 (N_21199,N_20958,N_20865);
or U21200 (N_21200,N_21194,N_21185);
and U21201 (N_21201,N_21047,N_21161);
nor U21202 (N_21202,N_21158,N_21028);
and U21203 (N_21203,N_21086,N_21004);
xor U21204 (N_21204,N_21180,N_21038);
nor U21205 (N_21205,N_21034,N_21113);
nor U21206 (N_21206,N_21046,N_21131);
or U21207 (N_21207,N_21159,N_21017);
xor U21208 (N_21208,N_21021,N_21013);
and U21209 (N_21209,N_21056,N_21177);
nand U21210 (N_21210,N_21150,N_21167);
nor U21211 (N_21211,N_21139,N_21045);
nand U21212 (N_21212,N_21066,N_21190);
xnor U21213 (N_21213,N_21101,N_21140);
and U21214 (N_21214,N_21076,N_21174);
or U21215 (N_21215,N_21157,N_21042);
nor U21216 (N_21216,N_21057,N_21077);
and U21217 (N_21217,N_21039,N_21054);
nor U21218 (N_21218,N_21058,N_21033);
nand U21219 (N_21219,N_21070,N_21093);
or U21220 (N_21220,N_21043,N_21097);
nor U21221 (N_21221,N_21120,N_21079);
nor U21222 (N_21222,N_21108,N_21105);
and U21223 (N_21223,N_21016,N_21106);
or U21224 (N_21224,N_21130,N_21169);
xor U21225 (N_21225,N_21145,N_21136);
or U21226 (N_21226,N_21068,N_21026);
or U21227 (N_21227,N_21142,N_21188);
nand U21228 (N_21228,N_21084,N_21110);
nor U21229 (N_21229,N_21029,N_21125);
nor U21230 (N_21230,N_21064,N_21162);
nand U21231 (N_21231,N_21176,N_21193);
xnor U21232 (N_21232,N_21137,N_21005);
nand U21233 (N_21233,N_21001,N_21144);
xnor U21234 (N_21234,N_21119,N_21006);
or U21235 (N_21235,N_21025,N_21148);
nor U21236 (N_21236,N_21087,N_21023);
xor U21237 (N_21237,N_21126,N_21069);
xnor U21238 (N_21238,N_21189,N_21133);
nand U21239 (N_21239,N_21184,N_21081);
xnor U21240 (N_21240,N_21165,N_21063);
nor U21241 (N_21241,N_21051,N_21114);
nand U21242 (N_21242,N_21109,N_21096);
nor U21243 (N_21243,N_21031,N_21022);
or U21244 (N_21244,N_21037,N_21098);
nor U21245 (N_21245,N_21020,N_21135);
nor U21246 (N_21246,N_21143,N_21155);
nor U21247 (N_21247,N_21099,N_21012);
and U21248 (N_21248,N_21062,N_21082);
xor U21249 (N_21249,N_21186,N_21112);
nand U21250 (N_21250,N_21027,N_21091);
nor U21251 (N_21251,N_21015,N_21030);
nand U21252 (N_21252,N_21040,N_21024);
nor U21253 (N_21253,N_21198,N_21192);
xnor U21254 (N_21254,N_21124,N_21168);
xnor U21255 (N_21255,N_21089,N_21094);
nand U21256 (N_21256,N_21059,N_21014);
nor U21257 (N_21257,N_21141,N_21151);
and U21258 (N_21258,N_21052,N_21060);
and U21259 (N_21259,N_21011,N_21072);
and U21260 (N_21260,N_21129,N_21127);
or U21261 (N_21261,N_21122,N_21041);
and U21262 (N_21262,N_21116,N_21050);
or U21263 (N_21263,N_21118,N_21195);
and U21264 (N_21264,N_21191,N_21163);
xor U21265 (N_21265,N_21035,N_21196);
and U21266 (N_21266,N_21010,N_21055);
nand U21267 (N_21267,N_21197,N_21103);
and U21268 (N_21268,N_21156,N_21173);
or U21269 (N_21269,N_21074,N_21147);
nor U21270 (N_21270,N_21009,N_21067);
xnor U21271 (N_21271,N_21134,N_21053);
xor U21272 (N_21272,N_21049,N_21061);
xnor U21273 (N_21273,N_21036,N_21115);
and U21274 (N_21274,N_21154,N_21111);
nor U21275 (N_21275,N_21175,N_21090);
and U21276 (N_21276,N_21171,N_21071);
nor U21277 (N_21277,N_21065,N_21019);
nand U21278 (N_21278,N_21138,N_21000);
or U21279 (N_21279,N_21080,N_21172);
nand U21280 (N_21280,N_21032,N_21107);
xor U21281 (N_21281,N_21100,N_21146);
nor U21282 (N_21282,N_21102,N_21073);
nand U21283 (N_21283,N_21092,N_21178);
or U21284 (N_21284,N_21187,N_21182);
and U21285 (N_21285,N_21104,N_21007);
nand U21286 (N_21286,N_21083,N_21170);
xor U21287 (N_21287,N_21085,N_21117);
nor U21288 (N_21288,N_21149,N_21078);
xor U21289 (N_21289,N_21160,N_21132);
xor U21290 (N_21290,N_21048,N_21088);
nor U21291 (N_21291,N_21003,N_21008);
xor U21292 (N_21292,N_21181,N_21199);
nor U21293 (N_21293,N_21179,N_21075);
nor U21294 (N_21294,N_21002,N_21123);
nand U21295 (N_21295,N_21153,N_21166);
xnor U21296 (N_21296,N_21095,N_21018);
xnor U21297 (N_21297,N_21164,N_21152);
and U21298 (N_21298,N_21183,N_21044);
and U21299 (N_21299,N_21128,N_21121);
and U21300 (N_21300,N_21180,N_21077);
xnor U21301 (N_21301,N_21003,N_21038);
and U21302 (N_21302,N_21143,N_21074);
nor U21303 (N_21303,N_21074,N_21177);
xor U21304 (N_21304,N_21086,N_21130);
nor U21305 (N_21305,N_21126,N_21015);
xor U21306 (N_21306,N_21183,N_21123);
or U21307 (N_21307,N_21092,N_21090);
nand U21308 (N_21308,N_21162,N_21136);
xor U21309 (N_21309,N_21059,N_21187);
nor U21310 (N_21310,N_21141,N_21126);
nor U21311 (N_21311,N_21033,N_21075);
nor U21312 (N_21312,N_21072,N_21139);
nand U21313 (N_21313,N_21057,N_21070);
nor U21314 (N_21314,N_21040,N_21128);
or U21315 (N_21315,N_21102,N_21163);
or U21316 (N_21316,N_21007,N_21182);
or U21317 (N_21317,N_21008,N_21020);
or U21318 (N_21318,N_21026,N_21004);
or U21319 (N_21319,N_21038,N_21041);
or U21320 (N_21320,N_21072,N_21119);
or U21321 (N_21321,N_21145,N_21032);
or U21322 (N_21322,N_21130,N_21017);
nor U21323 (N_21323,N_21112,N_21076);
nor U21324 (N_21324,N_21097,N_21050);
nand U21325 (N_21325,N_21003,N_21134);
nand U21326 (N_21326,N_21137,N_21020);
nand U21327 (N_21327,N_21103,N_21180);
nor U21328 (N_21328,N_21073,N_21173);
xor U21329 (N_21329,N_21050,N_21047);
or U21330 (N_21330,N_21098,N_21123);
nor U21331 (N_21331,N_21111,N_21063);
nor U21332 (N_21332,N_21192,N_21100);
nor U21333 (N_21333,N_21168,N_21006);
xnor U21334 (N_21334,N_21055,N_21104);
nor U21335 (N_21335,N_21043,N_21002);
nand U21336 (N_21336,N_21110,N_21129);
nor U21337 (N_21337,N_21076,N_21193);
and U21338 (N_21338,N_21093,N_21030);
and U21339 (N_21339,N_21091,N_21193);
nor U21340 (N_21340,N_21004,N_21145);
or U21341 (N_21341,N_21032,N_21116);
xor U21342 (N_21342,N_21076,N_21139);
and U21343 (N_21343,N_21117,N_21156);
nand U21344 (N_21344,N_21006,N_21135);
nor U21345 (N_21345,N_21172,N_21135);
xor U21346 (N_21346,N_21078,N_21009);
nand U21347 (N_21347,N_21121,N_21175);
xor U21348 (N_21348,N_21106,N_21183);
and U21349 (N_21349,N_21181,N_21008);
nor U21350 (N_21350,N_21033,N_21035);
nor U21351 (N_21351,N_21160,N_21108);
nand U21352 (N_21352,N_21063,N_21038);
nand U21353 (N_21353,N_21116,N_21158);
or U21354 (N_21354,N_21108,N_21100);
or U21355 (N_21355,N_21157,N_21095);
xnor U21356 (N_21356,N_21138,N_21002);
xnor U21357 (N_21357,N_21010,N_21091);
nand U21358 (N_21358,N_21011,N_21064);
or U21359 (N_21359,N_21196,N_21136);
xnor U21360 (N_21360,N_21029,N_21173);
and U21361 (N_21361,N_21002,N_21189);
nand U21362 (N_21362,N_21094,N_21076);
and U21363 (N_21363,N_21002,N_21046);
xor U21364 (N_21364,N_21151,N_21091);
nor U21365 (N_21365,N_21075,N_21110);
xnor U21366 (N_21366,N_21051,N_21040);
and U21367 (N_21367,N_21026,N_21041);
nand U21368 (N_21368,N_21031,N_21093);
nand U21369 (N_21369,N_21078,N_21151);
or U21370 (N_21370,N_21040,N_21033);
nor U21371 (N_21371,N_21169,N_21006);
xor U21372 (N_21372,N_21164,N_21010);
nand U21373 (N_21373,N_21027,N_21143);
or U21374 (N_21374,N_21031,N_21069);
xnor U21375 (N_21375,N_21037,N_21169);
xnor U21376 (N_21376,N_21009,N_21143);
or U21377 (N_21377,N_21057,N_21042);
nor U21378 (N_21378,N_21173,N_21196);
xor U21379 (N_21379,N_21143,N_21067);
and U21380 (N_21380,N_21030,N_21173);
nand U21381 (N_21381,N_21077,N_21053);
nor U21382 (N_21382,N_21078,N_21133);
and U21383 (N_21383,N_21042,N_21131);
and U21384 (N_21384,N_21088,N_21056);
nor U21385 (N_21385,N_21138,N_21053);
nand U21386 (N_21386,N_21017,N_21139);
xnor U21387 (N_21387,N_21058,N_21145);
or U21388 (N_21388,N_21097,N_21129);
xnor U21389 (N_21389,N_21151,N_21073);
nor U21390 (N_21390,N_21088,N_21188);
or U21391 (N_21391,N_21087,N_21092);
or U21392 (N_21392,N_21166,N_21124);
and U21393 (N_21393,N_21047,N_21180);
or U21394 (N_21394,N_21022,N_21091);
xor U21395 (N_21395,N_21189,N_21048);
nand U21396 (N_21396,N_21013,N_21023);
xnor U21397 (N_21397,N_21113,N_21100);
xnor U21398 (N_21398,N_21021,N_21117);
nand U21399 (N_21399,N_21115,N_21044);
xnor U21400 (N_21400,N_21381,N_21339);
nor U21401 (N_21401,N_21348,N_21261);
nand U21402 (N_21402,N_21320,N_21385);
nand U21403 (N_21403,N_21291,N_21301);
and U21404 (N_21404,N_21352,N_21215);
and U21405 (N_21405,N_21296,N_21266);
nor U21406 (N_21406,N_21246,N_21303);
nor U21407 (N_21407,N_21250,N_21248);
or U21408 (N_21408,N_21325,N_21384);
xor U21409 (N_21409,N_21207,N_21363);
or U21410 (N_21410,N_21213,N_21298);
or U21411 (N_21411,N_21333,N_21226);
and U21412 (N_21412,N_21257,N_21390);
xnor U21413 (N_21413,N_21350,N_21393);
and U21414 (N_21414,N_21377,N_21369);
or U21415 (N_21415,N_21287,N_21368);
nor U21416 (N_21416,N_21208,N_21217);
or U21417 (N_21417,N_21313,N_21254);
nand U21418 (N_21418,N_21346,N_21372);
or U21419 (N_21419,N_21335,N_21206);
or U21420 (N_21420,N_21280,N_21211);
or U21421 (N_21421,N_21290,N_21326);
nor U21422 (N_21422,N_21227,N_21225);
nor U21423 (N_21423,N_21391,N_21302);
nand U21424 (N_21424,N_21252,N_21315);
nand U21425 (N_21425,N_21281,N_21224);
xor U21426 (N_21426,N_21260,N_21338);
nand U21427 (N_21427,N_21233,N_21263);
and U21428 (N_21428,N_21230,N_21396);
xnor U21429 (N_21429,N_21240,N_21262);
xor U21430 (N_21430,N_21265,N_21221);
or U21431 (N_21431,N_21316,N_21319);
xnor U21432 (N_21432,N_21375,N_21355);
xnor U21433 (N_21433,N_21395,N_21289);
nand U21434 (N_21434,N_21276,N_21256);
or U21435 (N_21435,N_21274,N_21336);
nand U21436 (N_21436,N_21330,N_21380);
xor U21437 (N_21437,N_21202,N_21389);
nand U21438 (N_21438,N_21209,N_21249);
nand U21439 (N_21439,N_21340,N_21358);
nand U21440 (N_21440,N_21297,N_21397);
nor U21441 (N_21441,N_21272,N_21307);
xor U21442 (N_21442,N_21271,N_21200);
nor U21443 (N_21443,N_21270,N_21317);
and U21444 (N_21444,N_21223,N_21318);
nor U21445 (N_21445,N_21267,N_21360);
and U21446 (N_21446,N_21361,N_21204);
or U21447 (N_21447,N_21399,N_21214);
and U21448 (N_21448,N_21294,N_21388);
or U21449 (N_21449,N_21321,N_21324);
and U21450 (N_21450,N_21387,N_21218);
nor U21451 (N_21451,N_21362,N_21253);
nand U21452 (N_21452,N_21332,N_21382);
nand U21453 (N_21453,N_21285,N_21283);
xor U21454 (N_21454,N_21394,N_21251);
nand U21455 (N_21455,N_21354,N_21323);
xnor U21456 (N_21456,N_21231,N_21305);
and U21457 (N_21457,N_21247,N_21284);
and U21458 (N_21458,N_21311,N_21229);
nor U21459 (N_21459,N_21299,N_21349);
xnor U21460 (N_21460,N_21232,N_21365);
nor U21461 (N_21461,N_21376,N_21308);
or U21462 (N_21462,N_21259,N_21269);
nand U21463 (N_21463,N_21237,N_21242);
and U21464 (N_21464,N_21220,N_21378);
xnor U21465 (N_21465,N_21241,N_21342);
and U21466 (N_21466,N_21243,N_21245);
or U21467 (N_21467,N_21334,N_21373);
and U21468 (N_21468,N_21312,N_21219);
nor U21469 (N_21469,N_21364,N_21383);
nand U21470 (N_21470,N_21345,N_21392);
or U21471 (N_21471,N_21351,N_21304);
and U21472 (N_21472,N_21337,N_21329);
xnor U21473 (N_21473,N_21353,N_21344);
or U21474 (N_21474,N_21322,N_21292);
xnor U21475 (N_21475,N_21343,N_21386);
xor U21476 (N_21476,N_21216,N_21244);
nand U21477 (N_21477,N_21286,N_21306);
or U21478 (N_21478,N_21293,N_21228);
xor U21479 (N_21479,N_21279,N_21278);
nand U21480 (N_21480,N_21212,N_21359);
nor U21481 (N_21481,N_21277,N_21255);
xor U21482 (N_21482,N_21379,N_21203);
xor U21483 (N_21483,N_21357,N_21201);
and U21484 (N_21484,N_21258,N_21239);
nand U21485 (N_21485,N_21295,N_21236);
or U21486 (N_21486,N_21356,N_21328);
xnor U21487 (N_21487,N_21398,N_21341);
nor U21488 (N_21488,N_21275,N_21374);
nand U21489 (N_21489,N_21300,N_21234);
xor U21490 (N_21490,N_21282,N_21327);
and U21491 (N_21491,N_21288,N_21314);
xnor U21492 (N_21492,N_21264,N_21205);
xnor U21493 (N_21493,N_21366,N_21367);
nand U21494 (N_21494,N_21370,N_21210);
xnor U21495 (N_21495,N_21309,N_21310);
xor U21496 (N_21496,N_21371,N_21331);
and U21497 (N_21497,N_21273,N_21347);
or U21498 (N_21498,N_21222,N_21238);
nand U21499 (N_21499,N_21235,N_21268);
and U21500 (N_21500,N_21391,N_21394);
and U21501 (N_21501,N_21201,N_21277);
or U21502 (N_21502,N_21319,N_21203);
nand U21503 (N_21503,N_21305,N_21208);
nand U21504 (N_21504,N_21311,N_21254);
nor U21505 (N_21505,N_21304,N_21335);
or U21506 (N_21506,N_21304,N_21224);
nor U21507 (N_21507,N_21265,N_21305);
or U21508 (N_21508,N_21341,N_21209);
xor U21509 (N_21509,N_21314,N_21305);
and U21510 (N_21510,N_21273,N_21362);
xnor U21511 (N_21511,N_21242,N_21318);
and U21512 (N_21512,N_21283,N_21276);
and U21513 (N_21513,N_21283,N_21229);
xor U21514 (N_21514,N_21324,N_21308);
nand U21515 (N_21515,N_21246,N_21333);
or U21516 (N_21516,N_21213,N_21375);
and U21517 (N_21517,N_21338,N_21247);
nor U21518 (N_21518,N_21208,N_21207);
nor U21519 (N_21519,N_21356,N_21292);
nand U21520 (N_21520,N_21359,N_21232);
or U21521 (N_21521,N_21277,N_21252);
nor U21522 (N_21522,N_21223,N_21348);
xnor U21523 (N_21523,N_21204,N_21287);
nand U21524 (N_21524,N_21216,N_21209);
or U21525 (N_21525,N_21239,N_21271);
nor U21526 (N_21526,N_21338,N_21281);
nor U21527 (N_21527,N_21359,N_21254);
nor U21528 (N_21528,N_21318,N_21336);
xnor U21529 (N_21529,N_21204,N_21233);
or U21530 (N_21530,N_21312,N_21361);
nand U21531 (N_21531,N_21360,N_21309);
nor U21532 (N_21532,N_21212,N_21332);
nor U21533 (N_21533,N_21201,N_21230);
nand U21534 (N_21534,N_21281,N_21388);
nor U21535 (N_21535,N_21391,N_21333);
nor U21536 (N_21536,N_21385,N_21209);
and U21537 (N_21537,N_21327,N_21242);
or U21538 (N_21538,N_21226,N_21256);
nor U21539 (N_21539,N_21380,N_21349);
nand U21540 (N_21540,N_21262,N_21387);
nor U21541 (N_21541,N_21381,N_21235);
or U21542 (N_21542,N_21364,N_21389);
xor U21543 (N_21543,N_21316,N_21330);
nand U21544 (N_21544,N_21212,N_21277);
xor U21545 (N_21545,N_21264,N_21334);
nor U21546 (N_21546,N_21375,N_21382);
nor U21547 (N_21547,N_21325,N_21210);
and U21548 (N_21548,N_21248,N_21231);
nand U21549 (N_21549,N_21301,N_21358);
and U21550 (N_21550,N_21382,N_21312);
xor U21551 (N_21551,N_21219,N_21272);
or U21552 (N_21552,N_21338,N_21301);
and U21553 (N_21553,N_21345,N_21214);
and U21554 (N_21554,N_21395,N_21371);
nor U21555 (N_21555,N_21372,N_21359);
nand U21556 (N_21556,N_21243,N_21326);
xnor U21557 (N_21557,N_21339,N_21273);
nand U21558 (N_21558,N_21280,N_21332);
xnor U21559 (N_21559,N_21327,N_21336);
xor U21560 (N_21560,N_21282,N_21279);
or U21561 (N_21561,N_21236,N_21315);
nor U21562 (N_21562,N_21241,N_21258);
and U21563 (N_21563,N_21261,N_21321);
or U21564 (N_21564,N_21347,N_21243);
and U21565 (N_21565,N_21398,N_21364);
nand U21566 (N_21566,N_21212,N_21391);
nor U21567 (N_21567,N_21254,N_21273);
nor U21568 (N_21568,N_21391,N_21255);
xor U21569 (N_21569,N_21311,N_21325);
nand U21570 (N_21570,N_21339,N_21398);
and U21571 (N_21571,N_21253,N_21361);
or U21572 (N_21572,N_21313,N_21270);
nor U21573 (N_21573,N_21360,N_21315);
xor U21574 (N_21574,N_21349,N_21284);
xor U21575 (N_21575,N_21253,N_21262);
or U21576 (N_21576,N_21321,N_21365);
xor U21577 (N_21577,N_21220,N_21380);
xnor U21578 (N_21578,N_21339,N_21201);
or U21579 (N_21579,N_21303,N_21287);
nor U21580 (N_21580,N_21316,N_21374);
xnor U21581 (N_21581,N_21341,N_21314);
nand U21582 (N_21582,N_21358,N_21399);
or U21583 (N_21583,N_21385,N_21257);
nand U21584 (N_21584,N_21229,N_21236);
nor U21585 (N_21585,N_21353,N_21360);
nor U21586 (N_21586,N_21303,N_21272);
nor U21587 (N_21587,N_21307,N_21321);
nor U21588 (N_21588,N_21286,N_21225);
nor U21589 (N_21589,N_21284,N_21396);
or U21590 (N_21590,N_21270,N_21242);
nor U21591 (N_21591,N_21339,N_21223);
xnor U21592 (N_21592,N_21333,N_21377);
nand U21593 (N_21593,N_21364,N_21336);
nand U21594 (N_21594,N_21305,N_21350);
xor U21595 (N_21595,N_21313,N_21223);
nor U21596 (N_21596,N_21315,N_21226);
or U21597 (N_21597,N_21371,N_21222);
nor U21598 (N_21598,N_21230,N_21342);
or U21599 (N_21599,N_21393,N_21320);
and U21600 (N_21600,N_21589,N_21462);
or U21601 (N_21601,N_21440,N_21506);
nor U21602 (N_21602,N_21590,N_21432);
nand U21603 (N_21603,N_21470,N_21403);
or U21604 (N_21604,N_21425,N_21499);
and U21605 (N_21605,N_21463,N_21428);
nor U21606 (N_21606,N_21578,N_21493);
nand U21607 (N_21607,N_21515,N_21526);
or U21608 (N_21608,N_21449,N_21594);
and U21609 (N_21609,N_21460,N_21430);
and U21610 (N_21610,N_21560,N_21489);
and U21611 (N_21611,N_21473,N_21441);
xnor U21612 (N_21612,N_21537,N_21431);
xnor U21613 (N_21613,N_21471,N_21402);
nand U21614 (N_21614,N_21404,N_21567);
nor U21615 (N_21615,N_21447,N_21445);
and U21616 (N_21616,N_21521,N_21446);
nand U21617 (N_21617,N_21583,N_21479);
nor U21618 (N_21618,N_21465,N_21407);
or U21619 (N_21619,N_21448,N_21454);
and U21620 (N_21620,N_21482,N_21474);
xnor U21621 (N_21621,N_21557,N_21480);
nand U21622 (N_21622,N_21536,N_21467);
nand U21623 (N_21623,N_21481,N_21426);
and U21624 (N_21624,N_21512,N_21565);
or U21625 (N_21625,N_21504,N_21412);
xor U21626 (N_21626,N_21591,N_21555);
xor U21627 (N_21627,N_21476,N_21523);
and U21628 (N_21628,N_21478,N_21429);
or U21629 (N_21629,N_21486,N_21542);
nand U21630 (N_21630,N_21524,N_21417);
xnor U21631 (N_21631,N_21528,N_21502);
and U21632 (N_21632,N_21421,N_21541);
or U21633 (N_21633,N_21546,N_21527);
xor U21634 (N_21634,N_21405,N_21522);
and U21635 (N_21635,N_21571,N_21595);
or U21636 (N_21636,N_21458,N_21517);
nand U21637 (N_21637,N_21510,N_21501);
xor U21638 (N_21638,N_21436,N_21490);
nand U21639 (N_21639,N_21409,N_21566);
and U21640 (N_21640,N_21495,N_21535);
and U21641 (N_21641,N_21576,N_21586);
nand U21642 (N_21642,N_21497,N_21545);
nand U21643 (N_21643,N_21433,N_21410);
and U21644 (N_21644,N_21456,N_21599);
xor U21645 (N_21645,N_21573,N_21487);
xnor U21646 (N_21646,N_21548,N_21503);
nand U21647 (N_21647,N_21558,N_21435);
xnor U21648 (N_21648,N_21400,N_21437);
nor U21649 (N_21649,N_21508,N_21559);
nand U21650 (N_21650,N_21550,N_21549);
xnor U21651 (N_21651,N_21511,N_21563);
or U21652 (N_21652,N_21513,N_21498);
xor U21653 (N_21653,N_21581,N_21547);
nor U21654 (N_21654,N_21416,N_21569);
and U21655 (N_21655,N_21453,N_21485);
and U21656 (N_21656,N_21516,N_21411);
xor U21657 (N_21657,N_21418,N_21444);
and U21658 (N_21658,N_21584,N_21488);
nand U21659 (N_21659,N_21424,N_21450);
or U21660 (N_21660,N_21544,N_21543);
or U21661 (N_21661,N_21530,N_21423);
nand U21662 (N_21662,N_21455,N_21457);
or U21663 (N_21663,N_21492,N_21593);
nand U21664 (N_21664,N_21468,N_21434);
and U21665 (N_21665,N_21509,N_21451);
nor U21666 (N_21666,N_21551,N_21494);
or U21667 (N_21667,N_21529,N_21596);
and U21668 (N_21668,N_21408,N_21464);
and U21669 (N_21669,N_21556,N_21531);
and U21670 (N_21670,N_21427,N_21597);
and U21671 (N_21671,N_21598,N_21588);
nand U21672 (N_21672,N_21572,N_21419);
xor U21673 (N_21673,N_21401,N_21466);
or U21674 (N_21674,N_21592,N_21525);
or U21675 (N_21675,N_21459,N_21484);
or U21676 (N_21676,N_21422,N_21534);
xor U21677 (N_21677,N_21472,N_21538);
xnor U21678 (N_21678,N_21483,N_21577);
nor U21679 (N_21679,N_21539,N_21461);
nor U21680 (N_21680,N_21570,N_21475);
nor U21681 (N_21681,N_21518,N_21532);
nor U21682 (N_21682,N_21442,N_21415);
and U21683 (N_21683,N_21564,N_21469);
nand U21684 (N_21684,N_21520,N_21561);
nor U21685 (N_21685,N_21420,N_21443);
nor U21686 (N_21686,N_21552,N_21452);
or U21687 (N_21687,N_21438,N_21582);
nand U21688 (N_21688,N_21579,N_21568);
and U21689 (N_21689,N_21414,N_21580);
xnor U21690 (N_21690,N_21439,N_21507);
nor U21691 (N_21691,N_21533,N_21574);
xor U21692 (N_21692,N_21491,N_21587);
nand U21693 (N_21693,N_21505,N_21406);
and U21694 (N_21694,N_21585,N_21519);
and U21695 (N_21695,N_21500,N_21554);
nand U21696 (N_21696,N_21413,N_21575);
or U21697 (N_21697,N_21514,N_21496);
and U21698 (N_21698,N_21553,N_21540);
and U21699 (N_21699,N_21477,N_21562);
or U21700 (N_21700,N_21577,N_21576);
nor U21701 (N_21701,N_21550,N_21478);
nand U21702 (N_21702,N_21540,N_21518);
nand U21703 (N_21703,N_21530,N_21441);
xor U21704 (N_21704,N_21571,N_21587);
xor U21705 (N_21705,N_21451,N_21596);
nand U21706 (N_21706,N_21476,N_21474);
nand U21707 (N_21707,N_21565,N_21532);
nor U21708 (N_21708,N_21451,N_21469);
or U21709 (N_21709,N_21500,N_21424);
or U21710 (N_21710,N_21411,N_21582);
xor U21711 (N_21711,N_21426,N_21530);
and U21712 (N_21712,N_21526,N_21513);
xor U21713 (N_21713,N_21420,N_21452);
xor U21714 (N_21714,N_21584,N_21524);
and U21715 (N_21715,N_21499,N_21537);
nand U21716 (N_21716,N_21426,N_21550);
and U21717 (N_21717,N_21466,N_21531);
xor U21718 (N_21718,N_21433,N_21435);
nand U21719 (N_21719,N_21428,N_21430);
xor U21720 (N_21720,N_21471,N_21483);
or U21721 (N_21721,N_21498,N_21589);
and U21722 (N_21722,N_21583,N_21458);
or U21723 (N_21723,N_21571,N_21479);
xnor U21724 (N_21724,N_21566,N_21586);
xor U21725 (N_21725,N_21422,N_21486);
and U21726 (N_21726,N_21514,N_21459);
and U21727 (N_21727,N_21511,N_21478);
nand U21728 (N_21728,N_21454,N_21584);
or U21729 (N_21729,N_21419,N_21524);
nor U21730 (N_21730,N_21483,N_21556);
or U21731 (N_21731,N_21583,N_21427);
or U21732 (N_21732,N_21429,N_21470);
xnor U21733 (N_21733,N_21493,N_21536);
xnor U21734 (N_21734,N_21589,N_21417);
nand U21735 (N_21735,N_21402,N_21421);
nor U21736 (N_21736,N_21594,N_21572);
and U21737 (N_21737,N_21420,N_21570);
xnor U21738 (N_21738,N_21565,N_21527);
nand U21739 (N_21739,N_21415,N_21488);
nor U21740 (N_21740,N_21445,N_21461);
xnor U21741 (N_21741,N_21593,N_21431);
and U21742 (N_21742,N_21453,N_21412);
and U21743 (N_21743,N_21525,N_21540);
and U21744 (N_21744,N_21411,N_21548);
nand U21745 (N_21745,N_21575,N_21443);
nor U21746 (N_21746,N_21477,N_21598);
or U21747 (N_21747,N_21559,N_21424);
and U21748 (N_21748,N_21429,N_21575);
xnor U21749 (N_21749,N_21481,N_21552);
and U21750 (N_21750,N_21496,N_21488);
nor U21751 (N_21751,N_21565,N_21523);
or U21752 (N_21752,N_21573,N_21586);
or U21753 (N_21753,N_21515,N_21452);
xor U21754 (N_21754,N_21518,N_21429);
nor U21755 (N_21755,N_21419,N_21426);
and U21756 (N_21756,N_21547,N_21544);
nand U21757 (N_21757,N_21547,N_21522);
nand U21758 (N_21758,N_21459,N_21571);
nor U21759 (N_21759,N_21434,N_21589);
or U21760 (N_21760,N_21514,N_21442);
nand U21761 (N_21761,N_21475,N_21450);
xnor U21762 (N_21762,N_21417,N_21577);
nor U21763 (N_21763,N_21427,N_21591);
nor U21764 (N_21764,N_21467,N_21497);
nand U21765 (N_21765,N_21502,N_21431);
xor U21766 (N_21766,N_21571,N_21425);
nand U21767 (N_21767,N_21591,N_21533);
nor U21768 (N_21768,N_21480,N_21505);
or U21769 (N_21769,N_21538,N_21430);
and U21770 (N_21770,N_21569,N_21558);
or U21771 (N_21771,N_21576,N_21557);
xnor U21772 (N_21772,N_21468,N_21492);
xor U21773 (N_21773,N_21511,N_21489);
nor U21774 (N_21774,N_21488,N_21526);
and U21775 (N_21775,N_21557,N_21597);
nor U21776 (N_21776,N_21588,N_21494);
nor U21777 (N_21777,N_21530,N_21440);
nand U21778 (N_21778,N_21540,N_21503);
or U21779 (N_21779,N_21491,N_21561);
xnor U21780 (N_21780,N_21465,N_21400);
or U21781 (N_21781,N_21529,N_21440);
xnor U21782 (N_21782,N_21597,N_21542);
and U21783 (N_21783,N_21476,N_21597);
xnor U21784 (N_21784,N_21423,N_21417);
nand U21785 (N_21785,N_21470,N_21595);
and U21786 (N_21786,N_21414,N_21460);
and U21787 (N_21787,N_21424,N_21445);
nor U21788 (N_21788,N_21531,N_21452);
nand U21789 (N_21789,N_21564,N_21541);
or U21790 (N_21790,N_21586,N_21568);
or U21791 (N_21791,N_21463,N_21511);
nor U21792 (N_21792,N_21461,N_21426);
xor U21793 (N_21793,N_21544,N_21555);
xnor U21794 (N_21794,N_21487,N_21562);
nor U21795 (N_21795,N_21418,N_21495);
or U21796 (N_21796,N_21411,N_21578);
nand U21797 (N_21797,N_21555,N_21571);
nor U21798 (N_21798,N_21582,N_21498);
nor U21799 (N_21799,N_21590,N_21561);
or U21800 (N_21800,N_21651,N_21675);
or U21801 (N_21801,N_21607,N_21656);
and U21802 (N_21802,N_21682,N_21646);
or U21803 (N_21803,N_21748,N_21691);
and U21804 (N_21804,N_21718,N_21662);
and U21805 (N_21805,N_21739,N_21780);
and U21806 (N_21806,N_21647,N_21772);
and U21807 (N_21807,N_21658,N_21620);
xor U21808 (N_21808,N_21705,N_21613);
xnor U21809 (N_21809,N_21737,N_21758);
xor U21810 (N_21810,N_21615,N_21761);
nor U21811 (N_21811,N_21688,N_21717);
and U21812 (N_21812,N_21765,N_21794);
nor U21813 (N_21813,N_21669,N_21619);
nor U21814 (N_21814,N_21792,N_21751);
or U21815 (N_21815,N_21775,N_21707);
and U21816 (N_21816,N_21660,N_21612);
nand U21817 (N_21817,N_21655,N_21695);
nand U21818 (N_21818,N_21611,N_21652);
nand U21819 (N_21819,N_21648,N_21782);
or U21820 (N_21820,N_21668,N_21636);
nand U21821 (N_21821,N_21769,N_21664);
and U21822 (N_21822,N_21689,N_21784);
nor U21823 (N_21823,N_21706,N_21630);
nor U21824 (N_21824,N_21754,N_21745);
xor U21825 (N_21825,N_21633,N_21730);
nand U21826 (N_21826,N_21632,N_21679);
xor U21827 (N_21827,N_21733,N_21603);
nor U21828 (N_21828,N_21755,N_21740);
and U21829 (N_21829,N_21614,N_21616);
and U21830 (N_21830,N_21610,N_21684);
and U21831 (N_21831,N_21635,N_21697);
or U21832 (N_21832,N_21624,N_21771);
nor U21833 (N_21833,N_21791,N_21713);
nor U21834 (N_21834,N_21638,N_21731);
nand U21835 (N_21835,N_21628,N_21665);
nor U21836 (N_21836,N_21673,N_21753);
or U21837 (N_21837,N_21642,N_21768);
and U21838 (N_21838,N_21685,N_21732);
and U21839 (N_21839,N_21694,N_21721);
nor U21840 (N_21840,N_21779,N_21618);
nand U21841 (N_21841,N_21726,N_21634);
nor U21842 (N_21842,N_21774,N_21760);
and U21843 (N_21843,N_21738,N_21617);
xor U21844 (N_21844,N_21671,N_21702);
and U21845 (N_21845,N_21708,N_21698);
and U21846 (N_21846,N_21750,N_21604);
and U21847 (N_21847,N_21683,N_21622);
xnor U21848 (N_21848,N_21605,N_21757);
and U21849 (N_21849,N_21729,N_21746);
nor U21850 (N_21850,N_21667,N_21627);
or U21851 (N_21851,N_21722,N_21744);
and U21852 (N_21852,N_21720,N_21654);
nor U21853 (N_21853,N_21621,N_21709);
xnor U21854 (N_21854,N_21777,N_21600);
xor U21855 (N_21855,N_21645,N_21797);
nand U21856 (N_21856,N_21747,N_21723);
nor U21857 (N_21857,N_21734,N_21700);
or U21858 (N_21858,N_21736,N_21699);
xor U21859 (N_21859,N_21742,N_21696);
nor U21860 (N_21860,N_21785,N_21743);
nor U21861 (N_21861,N_21767,N_21631);
nor U21862 (N_21862,N_21653,N_21678);
or U21863 (N_21863,N_21650,N_21677);
or U21864 (N_21864,N_21639,N_21623);
and U21865 (N_21865,N_21762,N_21770);
and U21866 (N_21866,N_21672,N_21778);
nor U21867 (N_21867,N_21609,N_21786);
xnor U21868 (N_21868,N_21759,N_21712);
and U21869 (N_21869,N_21763,N_21663);
and U21870 (N_21870,N_21741,N_21626);
and U21871 (N_21871,N_21783,N_21661);
nand U21872 (N_21872,N_21681,N_21716);
and U21873 (N_21873,N_21703,N_21724);
nor U21874 (N_21874,N_21756,N_21796);
or U21875 (N_21875,N_21781,N_21629);
xor U21876 (N_21876,N_21788,N_21659);
nand U21877 (N_21877,N_21798,N_21725);
and U21878 (N_21878,N_21787,N_21752);
nand U21879 (N_21879,N_21674,N_21711);
or U21880 (N_21880,N_21649,N_21690);
or U21881 (N_21881,N_21773,N_21749);
xnor U21882 (N_21882,N_21657,N_21790);
nand U21883 (N_21883,N_21625,N_21701);
nand U21884 (N_21884,N_21641,N_21692);
nor U21885 (N_21885,N_21608,N_21766);
nor U21886 (N_21886,N_21687,N_21704);
nand U21887 (N_21887,N_21637,N_21735);
nor U21888 (N_21888,N_21666,N_21793);
xnor U21889 (N_21889,N_21764,N_21686);
xor U21890 (N_21890,N_21714,N_21640);
and U21891 (N_21891,N_21799,N_21680);
or U21892 (N_21892,N_21776,N_21710);
nor U21893 (N_21893,N_21795,N_21644);
xnor U21894 (N_21894,N_21727,N_21789);
nand U21895 (N_21895,N_21676,N_21643);
xnor U21896 (N_21896,N_21693,N_21728);
or U21897 (N_21897,N_21602,N_21670);
nand U21898 (N_21898,N_21601,N_21715);
or U21899 (N_21899,N_21606,N_21719);
or U21900 (N_21900,N_21761,N_21702);
and U21901 (N_21901,N_21695,N_21633);
xor U21902 (N_21902,N_21690,N_21747);
or U21903 (N_21903,N_21709,N_21744);
xnor U21904 (N_21904,N_21668,N_21631);
and U21905 (N_21905,N_21788,N_21774);
and U21906 (N_21906,N_21660,N_21658);
nor U21907 (N_21907,N_21796,N_21785);
nand U21908 (N_21908,N_21610,N_21780);
nand U21909 (N_21909,N_21710,N_21697);
or U21910 (N_21910,N_21781,N_21787);
nor U21911 (N_21911,N_21610,N_21669);
nand U21912 (N_21912,N_21798,N_21652);
or U21913 (N_21913,N_21657,N_21723);
nand U21914 (N_21914,N_21682,N_21799);
nor U21915 (N_21915,N_21731,N_21686);
or U21916 (N_21916,N_21659,N_21646);
nand U21917 (N_21917,N_21671,N_21788);
nand U21918 (N_21918,N_21611,N_21621);
xnor U21919 (N_21919,N_21694,N_21731);
nand U21920 (N_21920,N_21740,N_21718);
nand U21921 (N_21921,N_21796,N_21698);
nand U21922 (N_21922,N_21749,N_21644);
nand U21923 (N_21923,N_21665,N_21721);
nand U21924 (N_21924,N_21779,N_21707);
nand U21925 (N_21925,N_21772,N_21681);
nor U21926 (N_21926,N_21666,N_21620);
nand U21927 (N_21927,N_21733,N_21688);
nand U21928 (N_21928,N_21714,N_21633);
nor U21929 (N_21929,N_21759,N_21643);
nand U21930 (N_21930,N_21769,N_21644);
nor U21931 (N_21931,N_21656,N_21715);
or U21932 (N_21932,N_21790,N_21653);
nand U21933 (N_21933,N_21744,N_21661);
nor U21934 (N_21934,N_21620,N_21643);
xor U21935 (N_21935,N_21704,N_21645);
nand U21936 (N_21936,N_21740,N_21733);
or U21937 (N_21937,N_21732,N_21748);
nor U21938 (N_21938,N_21607,N_21768);
and U21939 (N_21939,N_21762,N_21767);
nor U21940 (N_21940,N_21626,N_21692);
nand U21941 (N_21941,N_21637,N_21687);
nor U21942 (N_21942,N_21607,N_21788);
xor U21943 (N_21943,N_21634,N_21742);
nor U21944 (N_21944,N_21688,N_21755);
and U21945 (N_21945,N_21778,N_21711);
and U21946 (N_21946,N_21788,N_21783);
nand U21947 (N_21947,N_21638,N_21726);
nor U21948 (N_21948,N_21798,N_21632);
xor U21949 (N_21949,N_21787,N_21796);
xor U21950 (N_21950,N_21715,N_21639);
nand U21951 (N_21951,N_21631,N_21724);
nor U21952 (N_21952,N_21774,N_21633);
nor U21953 (N_21953,N_21606,N_21790);
nor U21954 (N_21954,N_21625,N_21602);
nand U21955 (N_21955,N_21700,N_21725);
xnor U21956 (N_21956,N_21714,N_21776);
nand U21957 (N_21957,N_21753,N_21725);
nand U21958 (N_21958,N_21706,N_21633);
xor U21959 (N_21959,N_21687,N_21720);
or U21960 (N_21960,N_21686,N_21653);
xor U21961 (N_21961,N_21697,N_21625);
or U21962 (N_21962,N_21704,N_21629);
xnor U21963 (N_21963,N_21795,N_21767);
nor U21964 (N_21964,N_21602,N_21629);
nand U21965 (N_21965,N_21757,N_21726);
and U21966 (N_21966,N_21662,N_21602);
nor U21967 (N_21967,N_21798,N_21643);
xnor U21968 (N_21968,N_21625,N_21773);
xnor U21969 (N_21969,N_21756,N_21621);
nor U21970 (N_21970,N_21719,N_21623);
nand U21971 (N_21971,N_21772,N_21786);
nor U21972 (N_21972,N_21748,N_21714);
nand U21973 (N_21973,N_21760,N_21730);
xnor U21974 (N_21974,N_21768,N_21645);
xnor U21975 (N_21975,N_21723,N_21750);
and U21976 (N_21976,N_21674,N_21666);
nor U21977 (N_21977,N_21619,N_21624);
or U21978 (N_21978,N_21761,N_21651);
and U21979 (N_21979,N_21678,N_21638);
nand U21980 (N_21980,N_21778,N_21666);
nand U21981 (N_21981,N_21631,N_21654);
nand U21982 (N_21982,N_21796,N_21696);
nand U21983 (N_21983,N_21736,N_21777);
xnor U21984 (N_21984,N_21664,N_21783);
and U21985 (N_21985,N_21696,N_21763);
or U21986 (N_21986,N_21759,N_21645);
and U21987 (N_21987,N_21624,N_21782);
or U21988 (N_21988,N_21782,N_21632);
xor U21989 (N_21989,N_21745,N_21781);
and U21990 (N_21990,N_21766,N_21763);
nand U21991 (N_21991,N_21734,N_21797);
or U21992 (N_21992,N_21624,N_21726);
and U21993 (N_21993,N_21750,N_21678);
nor U21994 (N_21994,N_21774,N_21641);
nand U21995 (N_21995,N_21634,N_21737);
nor U21996 (N_21996,N_21738,N_21675);
nor U21997 (N_21997,N_21658,N_21636);
xor U21998 (N_21998,N_21662,N_21737);
xnor U21999 (N_21999,N_21786,N_21610);
xor U22000 (N_22000,N_21965,N_21801);
nand U22001 (N_22001,N_21853,N_21932);
or U22002 (N_22002,N_21950,N_21958);
xnor U22003 (N_22003,N_21944,N_21945);
nand U22004 (N_22004,N_21880,N_21829);
or U22005 (N_22005,N_21802,N_21828);
nor U22006 (N_22006,N_21873,N_21878);
or U22007 (N_22007,N_21896,N_21888);
xor U22008 (N_22008,N_21941,N_21893);
and U22009 (N_22009,N_21961,N_21832);
nor U22010 (N_22010,N_21972,N_21843);
and U22011 (N_22011,N_21835,N_21844);
nor U22012 (N_22012,N_21865,N_21846);
nor U22013 (N_22013,N_21892,N_21823);
and U22014 (N_22014,N_21962,N_21871);
or U22015 (N_22015,N_21909,N_21803);
nor U22016 (N_22016,N_21904,N_21948);
xnor U22017 (N_22017,N_21947,N_21842);
nand U22018 (N_22018,N_21805,N_21991);
nand U22019 (N_22019,N_21920,N_21915);
nand U22020 (N_22020,N_21862,N_21860);
and U22021 (N_22021,N_21851,N_21960);
nand U22022 (N_22022,N_21913,N_21907);
nor U22023 (N_22023,N_21867,N_21983);
nand U22024 (N_22024,N_21859,N_21976);
nor U22025 (N_22025,N_21968,N_21822);
nand U22026 (N_22026,N_21815,N_21898);
or U22027 (N_22027,N_21930,N_21837);
nor U22028 (N_22028,N_21916,N_21981);
or U22029 (N_22029,N_21877,N_21914);
nor U22030 (N_22030,N_21998,N_21818);
xnor U22031 (N_22031,N_21955,N_21923);
xor U22032 (N_22032,N_21970,N_21912);
and U22033 (N_22033,N_21813,N_21831);
and U22034 (N_22034,N_21868,N_21845);
xor U22035 (N_22035,N_21886,N_21870);
xor U22036 (N_22036,N_21926,N_21850);
or U22037 (N_22037,N_21977,N_21937);
xor U22038 (N_22038,N_21999,N_21890);
xnor U22039 (N_22039,N_21839,N_21942);
xor U22040 (N_22040,N_21804,N_21833);
or U22041 (N_22041,N_21939,N_21899);
or U22042 (N_22042,N_21966,N_21992);
xor U22043 (N_22043,N_21973,N_21919);
xnor U22044 (N_22044,N_21943,N_21967);
and U22045 (N_22045,N_21817,N_21901);
nand U22046 (N_22046,N_21935,N_21993);
nand U22047 (N_22047,N_21986,N_21875);
or U22048 (N_22048,N_21979,N_21849);
nand U22049 (N_22049,N_21994,N_21820);
xor U22050 (N_22050,N_21963,N_21940);
nor U22051 (N_22051,N_21985,N_21808);
xor U22052 (N_22052,N_21969,N_21934);
nor U22053 (N_22053,N_21897,N_21929);
xnor U22054 (N_22054,N_21952,N_21964);
xor U22055 (N_22055,N_21995,N_21905);
nor U22056 (N_22056,N_21956,N_21874);
nand U22057 (N_22057,N_21816,N_21987);
xnor U22058 (N_22058,N_21910,N_21924);
nor U22059 (N_22059,N_21869,N_21911);
nand U22060 (N_22060,N_21827,N_21996);
or U22061 (N_22061,N_21882,N_21903);
or U22062 (N_22062,N_21938,N_21811);
or U22063 (N_22063,N_21980,N_21821);
nand U22064 (N_22064,N_21847,N_21885);
and U22065 (N_22065,N_21806,N_21982);
nor U22066 (N_22066,N_21978,N_21819);
xnor U22067 (N_22067,N_21864,N_21984);
xnor U22068 (N_22068,N_21830,N_21848);
nand U22069 (N_22069,N_21936,N_21918);
nor U22070 (N_22070,N_21989,N_21836);
and U22071 (N_22071,N_21834,N_21951);
nand U22072 (N_22072,N_21933,N_21990);
or U22073 (N_22073,N_21974,N_21809);
or U22074 (N_22074,N_21906,N_21810);
or U22075 (N_22075,N_21887,N_21946);
xor U22076 (N_22076,N_21953,N_21858);
or U22077 (N_22077,N_21800,N_21866);
xnor U22078 (N_22078,N_21957,N_21876);
or U22079 (N_22079,N_21838,N_21883);
or U22080 (N_22080,N_21959,N_21863);
nand U22081 (N_22081,N_21807,N_21988);
or U22082 (N_22082,N_21856,N_21971);
xor U22083 (N_22083,N_21889,N_21921);
nor U22084 (N_22084,N_21922,N_21884);
nand U22085 (N_22085,N_21902,N_21881);
nor U22086 (N_22086,N_21928,N_21894);
or U22087 (N_22087,N_21852,N_21825);
or U22088 (N_22088,N_21997,N_21931);
and U22089 (N_22089,N_21841,N_21855);
and U22090 (N_22090,N_21925,N_21954);
nand U22091 (N_22091,N_21872,N_21975);
nor U22092 (N_22092,N_21895,N_21857);
or U22093 (N_22093,N_21900,N_21854);
and U22094 (N_22094,N_21879,N_21814);
nand U22095 (N_22095,N_21824,N_21840);
nor U22096 (N_22096,N_21908,N_21861);
or U22097 (N_22097,N_21949,N_21891);
and U22098 (N_22098,N_21826,N_21812);
xor U22099 (N_22099,N_21917,N_21927);
xnor U22100 (N_22100,N_21851,N_21968);
and U22101 (N_22101,N_21924,N_21864);
or U22102 (N_22102,N_21862,N_21889);
and U22103 (N_22103,N_21955,N_21802);
xnor U22104 (N_22104,N_21898,N_21983);
and U22105 (N_22105,N_21859,N_21885);
and U22106 (N_22106,N_21857,N_21994);
nor U22107 (N_22107,N_21850,N_21833);
and U22108 (N_22108,N_21912,N_21903);
xnor U22109 (N_22109,N_21868,N_21849);
or U22110 (N_22110,N_21840,N_21915);
or U22111 (N_22111,N_21820,N_21976);
nand U22112 (N_22112,N_21926,N_21887);
or U22113 (N_22113,N_21860,N_21898);
nand U22114 (N_22114,N_21939,N_21903);
xor U22115 (N_22115,N_21961,N_21991);
xnor U22116 (N_22116,N_21872,N_21997);
xor U22117 (N_22117,N_21959,N_21812);
xor U22118 (N_22118,N_21886,N_21881);
nand U22119 (N_22119,N_21961,N_21815);
or U22120 (N_22120,N_21899,N_21839);
or U22121 (N_22121,N_21950,N_21817);
xor U22122 (N_22122,N_21903,N_21850);
or U22123 (N_22123,N_21981,N_21914);
xnor U22124 (N_22124,N_21899,N_21934);
xnor U22125 (N_22125,N_21954,N_21958);
or U22126 (N_22126,N_21879,N_21928);
nor U22127 (N_22127,N_21802,N_21826);
xor U22128 (N_22128,N_21975,N_21846);
and U22129 (N_22129,N_21959,N_21893);
xor U22130 (N_22130,N_21925,N_21910);
and U22131 (N_22131,N_21804,N_21969);
and U22132 (N_22132,N_21925,N_21946);
nor U22133 (N_22133,N_21924,N_21898);
xnor U22134 (N_22134,N_21802,N_21839);
nand U22135 (N_22135,N_21965,N_21803);
or U22136 (N_22136,N_21861,N_21950);
and U22137 (N_22137,N_21844,N_21979);
nor U22138 (N_22138,N_21835,N_21847);
nand U22139 (N_22139,N_21974,N_21921);
nor U22140 (N_22140,N_21801,N_21976);
or U22141 (N_22141,N_21828,N_21870);
or U22142 (N_22142,N_21854,N_21871);
xor U22143 (N_22143,N_21877,N_21903);
or U22144 (N_22144,N_21952,N_21847);
and U22145 (N_22145,N_21959,N_21895);
nand U22146 (N_22146,N_21970,N_21879);
xnor U22147 (N_22147,N_21864,N_21958);
and U22148 (N_22148,N_21872,N_21915);
nor U22149 (N_22149,N_21941,N_21864);
xnor U22150 (N_22150,N_21977,N_21818);
nor U22151 (N_22151,N_21965,N_21858);
nor U22152 (N_22152,N_21894,N_21830);
and U22153 (N_22153,N_21809,N_21802);
xnor U22154 (N_22154,N_21861,N_21943);
nand U22155 (N_22155,N_21881,N_21944);
and U22156 (N_22156,N_21847,N_21903);
nand U22157 (N_22157,N_21818,N_21949);
xnor U22158 (N_22158,N_21840,N_21942);
nor U22159 (N_22159,N_21800,N_21966);
and U22160 (N_22160,N_21952,N_21867);
or U22161 (N_22161,N_21964,N_21907);
or U22162 (N_22162,N_21827,N_21983);
xnor U22163 (N_22163,N_21947,N_21888);
xnor U22164 (N_22164,N_21820,N_21990);
xnor U22165 (N_22165,N_21907,N_21909);
xor U22166 (N_22166,N_21825,N_21916);
nand U22167 (N_22167,N_21813,N_21871);
xor U22168 (N_22168,N_21989,N_21921);
and U22169 (N_22169,N_21958,N_21868);
xor U22170 (N_22170,N_21996,N_21989);
or U22171 (N_22171,N_21940,N_21811);
and U22172 (N_22172,N_21821,N_21885);
nor U22173 (N_22173,N_21958,N_21999);
or U22174 (N_22174,N_21904,N_21811);
or U22175 (N_22175,N_21852,N_21847);
nor U22176 (N_22176,N_21814,N_21928);
and U22177 (N_22177,N_21865,N_21968);
or U22178 (N_22178,N_21884,N_21915);
xor U22179 (N_22179,N_21923,N_21861);
xnor U22180 (N_22180,N_21813,N_21845);
and U22181 (N_22181,N_21906,N_21909);
nor U22182 (N_22182,N_21908,N_21821);
nor U22183 (N_22183,N_21994,N_21876);
and U22184 (N_22184,N_21928,N_21934);
xnor U22185 (N_22185,N_21811,N_21888);
and U22186 (N_22186,N_21881,N_21873);
nand U22187 (N_22187,N_21833,N_21908);
nor U22188 (N_22188,N_21951,N_21805);
and U22189 (N_22189,N_21854,N_21923);
or U22190 (N_22190,N_21827,N_21949);
nor U22191 (N_22191,N_21999,N_21957);
nor U22192 (N_22192,N_21888,N_21921);
nand U22193 (N_22193,N_21914,N_21978);
and U22194 (N_22194,N_21893,N_21956);
or U22195 (N_22195,N_21865,N_21824);
or U22196 (N_22196,N_21934,N_21945);
and U22197 (N_22197,N_21814,N_21816);
nand U22198 (N_22198,N_21827,N_21938);
nand U22199 (N_22199,N_21840,N_21933);
or U22200 (N_22200,N_22025,N_22182);
nor U22201 (N_22201,N_22089,N_22164);
and U22202 (N_22202,N_22049,N_22058);
or U22203 (N_22203,N_22096,N_22119);
nor U22204 (N_22204,N_22002,N_22067);
and U22205 (N_22205,N_22151,N_22059);
xor U22206 (N_22206,N_22028,N_22142);
xor U22207 (N_22207,N_22101,N_22020);
or U22208 (N_22208,N_22161,N_22055);
nor U22209 (N_22209,N_22043,N_22186);
or U22210 (N_22210,N_22039,N_22197);
nand U22211 (N_22211,N_22183,N_22083);
nor U22212 (N_22212,N_22162,N_22037);
or U22213 (N_22213,N_22149,N_22194);
xnor U22214 (N_22214,N_22184,N_22031);
xnor U22215 (N_22215,N_22065,N_22198);
and U22216 (N_22216,N_22073,N_22195);
nand U22217 (N_22217,N_22085,N_22010);
nand U22218 (N_22218,N_22106,N_22179);
and U22219 (N_22219,N_22047,N_22018);
xor U22220 (N_22220,N_22094,N_22013);
and U22221 (N_22221,N_22045,N_22076);
and U22222 (N_22222,N_22092,N_22057);
and U22223 (N_22223,N_22030,N_22160);
nand U22224 (N_22224,N_22177,N_22107);
and U22225 (N_22225,N_22087,N_22185);
or U22226 (N_22226,N_22064,N_22146);
nor U22227 (N_22227,N_22122,N_22144);
xnor U22228 (N_22228,N_22128,N_22000);
nor U22229 (N_22229,N_22109,N_22044);
nor U22230 (N_22230,N_22034,N_22007);
nor U22231 (N_22231,N_22021,N_22040);
nand U22232 (N_22232,N_22170,N_22052);
nor U22233 (N_22233,N_22078,N_22102);
xor U22234 (N_22234,N_22100,N_22036);
nor U22235 (N_22235,N_22108,N_22066);
or U22236 (N_22236,N_22086,N_22095);
xnor U22237 (N_22237,N_22143,N_22019);
nand U22238 (N_22238,N_22169,N_22014);
nand U22239 (N_22239,N_22113,N_22104);
or U22240 (N_22240,N_22015,N_22115);
nand U22241 (N_22241,N_22081,N_22153);
nor U22242 (N_22242,N_22071,N_22112);
or U22243 (N_22243,N_22121,N_22068);
xnor U22244 (N_22244,N_22004,N_22165);
or U22245 (N_22245,N_22105,N_22080);
and U22246 (N_22246,N_22134,N_22125);
nor U22247 (N_22247,N_22166,N_22070);
xor U22248 (N_22248,N_22190,N_22074);
and U22249 (N_22249,N_22154,N_22003);
xnor U22250 (N_22250,N_22079,N_22111);
nand U22251 (N_22251,N_22022,N_22145);
xor U22252 (N_22252,N_22054,N_22168);
nand U22253 (N_22253,N_22163,N_22041);
xnor U22254 (N_22254,N_22118,N_22050);
xnor U22255 (N_22255,N_22131,N_22141);
or U22256 (N_22256,N_22140,N_22192);
xnor U22257 (N_22257,N_22093,N_22061);
or U22258 (N_22258,N_22199,N_22187);
or U22259 (N_22259,N_22193,N_22167);
xnor U22260 (N_22260,N_22088,N_22042);
xnor U22261 (N_22261,N_22126,N_22117);
nand U22262 (N_22262,N_22129,N_22172);
and U22263 (N_22263,N_22016,N_22051);
or U22264 (N_22264,N_22176,N_22060);
or U22265 (N_22265,N_22048,N_22124);
xor U22266 (N_22266,N_22120,N_22046);
and U22267 (N_22267,N_22178,N_22099);
xnor U22268 (N_22268,N_22011,N_22006);
or U22269 (N_22269,N_22038,N_22147);
xor U22270 (N_22270,N_22158,N_22132);
nor U22271 (N_22271,N_22171,N_22084);
nand U22272 (N_22272,N_22024,N_22114);
nor U22273 (N_22273,N_22133,N_22138);
xor U22274 (N_22274,N_22150,N_22116);
and U22275 (N_22275,N_22180,N_22026);
nand U22276 (N_22276,N_22191,N_22137);
nor U22277 (N_22277,N_22157,N_22152);
nand U22278 (N_22278,N_22072,N_22097);
and U22279 (N_22279,N_22127,N_22027);
nor U22280 (N_22280,N_22005,N_22181);
nor U22281 (N_22281,N_22156,N_22130);
nor U22282 (N_22282,N_22056,N_22090);
or U22283 (N_22283,N_22035,N_22091);
xor U22284 (N_22284,N_22196,N_22159);
or U22285 (N_22285,N_22053,N_22062);
and U22286 (N_22286,N_22082,N_22033);
or U22287 (N_22287,N_22175,N_22001);
or U22288 (N_22288,N_22098,N_22063);
xnor U22289 (N_22289,N_22110,N_22174);
and U22290 (N_22290,N_22188,N_22135);
nor U22291 (N_22291,N_22155,N_22069);
nand U22292 (N_22292,N_22023,N_22173);
nor U22293 (N_22293,N_22075,N_22148);
and U22294 (N_22294,N_22009,N_22077);
nor U22295 (N_22295,N_22123,N_22136);
nor U22296 (N_22296,N_22189,N_22017);
nand U22297 (N_22297,N_22012,N_22008);
and U22298 (N_22298,N_22139,N_22032);
xor U22299 (N_22299,N_22103,N_22029);
and U22300 (N_22300,N_22103,N_22120);
nor U22301 (N_22301,N_22157,N_22025);
nor U22302 (N_22302,N_22075,N_22166);
nand U22303 (N_22303,N_22102,N_22149);
and U22304 (N_22304,N_22155,N_22087);
and U22305 (N_22305,N_22196,N_22184);
nand U22306 (N_22306,N_22178,N_22029);
or U22307 (N_22307,N_22070,N_22103);
and U22308 (N_22308,N_22084,N_22196);
nor U22309 (N_22309,N_22075,N_22090);
and U22310 (N_22310,N_22106,N_22183);
nand U22311 (N_22311,N_22127,N_22103);
or U22312 (N_22312,N_22028,N_22043);
xor U22313 (N_22313,N_22154,N_22086);
and U22314 (N_22314,N_22132,N_22061);
or U22315 (N_22315,N_22097,N_22046);
nand U22316 (N_22316,N_22017,N_22091);
or U22317 (N_22317,N_22160,N_22025);
nand U22318 (N_22318,N_22100,N_22094);
and U22319 (N_22319,N_22092,N_22165);
xnor U22320 (N_22320,N_22152,N_22150);
xnor U22321 (N_22321,N_22167,N_22153);
or U22322 (N_22322,N_22052,N_22190);
or U22323 (N_22323,N_22179,N_22174);
nand U22324 (N_22324,N_22120,N_22189);
or U22325 (N_22325,N_22067,N_22070);
xnor U22326 (N_22326,N_22145,N_22095);
or U22327 (N_22327,N_22057,N_22124);
and U22328 (N_22328,N_22179,N_22093);
and U22329 (N_22329,N_22038,N_22099);
nand U22330 (N_22330,N_22180,N_22039);
nor U22331 (N_22331,N_22020,N_22081);
xor U22332 (N_22332,N_22139,N_22159);
and U22333 (N_22333,N_22123,N_22143);
and U22334 (N_22334,N_22127,N_22165);
nor U22335 (N_22335,N_22197,N_22185);
and U22336 (N_22336,N_22158,N_22136);
nor U22337 (N_22337,N_22102,N_22130);
nor U22338 (N_22338,N_22120,N_22010);
nor U22339 (N_22339,N_22109,N_22100);
and U22340 (N_22340,N_22123,N_22174);
and U22341 (N_22341,N_22131,N_22027);
or U22342 (N_22342,N_22014,N_22195);
nor U22343 (N_22343,N_22126,N_22082);
nand U22344 (N_22344,N_22149,N_22091);
nor U22345 (N_22345,N_22024,N_22150);
xnor U22346 (N_22346,N_22130,N_22170);
nor U22347 (N_22347,N_22050,N_22054);
and U22348 (N_22348,N_22052,N_22199);
nand U22349 (N_22349,N_22068,N_22123);
nor U22350 (N_22350,N_22092,N_22051);
nand U22351 (N_22351,N_22084,N_22001);
nor U22352 (N_22352,N_22107,N_22108);
and U22353 (N_22353,N_22139,N_22121);
nand U22354 (N_22354,N_22037,N_22168);
nor U22355 (N_22355,N_22109,N_22139);
or U22356 (N_22356,N_22144,N_22063);
and U22357 (N_22357,N_22005,N_22133);
nor U22358 (N_22358,N_22079,N_22153);
or U22359 (N_22359,N_22040,N_22176);
xor U22360 (N_22360,N_22149,N_22195);
and U22361 (N_22361,N_22129,N_22101);
xnor U22362 (N_22362,N_22085,N_22082);
and U22363 (N_22363,N_22011,N_22136);
and U22364 (N_22364,N_22184,N_22083);
xnor U22365 (N_22365,N_22042,N_22026);
and U22366 (N_22366,N_22137,N_22143);
nand U22367 (N_22367,N_22068,N_22141);
nor U22368 (N_22368,N_22069,N_22192);
xor U22369 (N_22369,N_22005,N_22007);
and U22370 (N_22370,N_22025,N_22149);
or U22371 (N_22371,N_22182,N_22139);
and U22372 (N_22372,N_22102,N_22172);
xnor U22373 (N_22373,N_22090,N_22043);
or U22374 (N_22374,N_22113,N_22047);
and U22375 (N_22375,N_22189,N_22171);
or U22376 (N_22376,N_22096,N_22039);
nand U22377 (N_22377,N_22197,N_22084);
nor U22378 (N_22378,N_22066,N_22107);
xor U22379 (N_22379,N_22121,N_22164);
nand U22380 (N_22380,N_22007,N_22110);
xnor U22381 (N_22381,N_22036,N_22027);
or U22382 (N_22382,N_22057,N_22094);
and U22383 (N_22383,N_22151,N_22135);
nor U22384 (N_22384,N_22054,N_22137);
nor U22385 (N_22385,N_22147,N_22077);
nand U22386 (N_22386,N_22139,N_22144);
and U22387 (N_22387,N_22159,N_22136);
and U22388 (N_22388,N_22194,N_22183);
nand U22389 (N_22389,N_22016,N_22183);
and U22390 (N_22390,N_22076,N_22062);
xnor U22391 (N_22391,N_22140,N_22095);
and U22392 (N_22392,N_22061,N_22041);
or U22393 (N_22393,N_22061,N_22053);
or U22394 (N_22394,N_22197,N_22055);
nand U22395 (N_22395,N_22030,N_22185);
and U22396 (N_22396,N_22174,N_22199);
xnor U22397 (N_22397,N_22060,N_22145);
xor U22398 (N_22398,N_22130,N_22083);
nor U22399 (N_22399,N_22056,N_22181);
and U22400 (N_22400,N_22397,N_22266);
nor U22401 (N_22401,N_22261,N_22207);
or U22402 (N_22402,N_22217,N_22253);
xor U22403 (N_22403,N_22359,N_22386);
and U22404 (N_22404,N_22333,N_22241);
xnor U22405 (N_22405,N_22204,N_22220);
xnor U22406 (N_22406,N_22358,N_22340);
or U22407 (N_22407,N_22210,N_22327);
nand U22408 (N_22408,N_22395,N_22249);
nand U22409 (N_22409,N_22259,N_22376);
and U22410 (N_22410,N_22320,N_22339);
xor U22411 (N_22411,N_22342,N_22301);
xor U22412 (N_22412,N_22276,N_22390);
xnor U22413 (N_22413,N_22265,N_22236);
or U22414 (N_22414,N_22350,N_22307);
or U22415 (N_22415,N_22293,N_22300);
or U22416 (N_22416,N_22349,N_22393);
and U22417 (N_22417,N_22343,N_22371);
nand U22418 (N_22418,N_22351,N_22360);
xor U22419 (N_22419,N_22332,N_22235);
or U22420 (N_22420,N_22305,N_22285);
xor U22421 (N_22421,N_22385,N_22312);
xnor U22422 (N_22422,N_22231,N_22304);
xor U22423 (N_22423,N_22200,N_22341);
or U22424 (N_22424,N_22330,N_22257);
nand U22425 (N_22425,N_22337,N_22211);
nand U22426 (N_22426,N_22348,N_22223);
or U22427 (N_22427,N_22338,N_22316);
and U22428 (N_22428,N_22357,N_22203);
and U22429 (N_22429,N_22329,N_22234);
nor U22430 (N_22430,N_22399,N_22388);
xnor U22431 (N_22431,N_22296,N_22324);
and U22432 (N_22432,N_22273,N_22391);
or U22433 (N_22433,N_22284,N_22379);
nand U22434 (N_22434,N_22290,N_22322);
nor U22435 (N_22435,N_22201,N_22226);
nor U22436 (N_22436,N_22370,N_22228);
nor U22437 (N_22437,N_22238,N_22209);
or U22438 (N_22438,N_22323,N_22274);
nand U22439 (N_22439,N_22287,N_22394);
or U22440 (N_22440,N_22381,N_22263);
or U22441 (N_22441,N_22354,N_22278);
nand U22442 (N_22442,N_22315,N_22355);
xor U22443 (N_22443,N_22294,N_22272);
nor U22444 (N_22444,N_22310,N_22346);
nor U22445 (N_22445,N_22214,N_22363);
nor U22446 (N_22446,N_22365,N_22206);
xnor U22447 (N_22447,N_22202,N_22280);
and U22448 (N_22448,N_22392,N_22335);
nor U22449 (N_22449,N_22283,N_22375);
nand U22450 (N_22450,N_22242,N_22245);
xor U22451 (N_22451,N_22275,N_22254);
xnor U22452 (N_22452,N_22225,N_22309);
xnor U22453 (N_22453,N_22252,N_22318);
nand U22454 (N_22454,N_22213,N_22319);
and U22455 (N_22455,N_22384,N_22295);
and U22456 (N_22456,N_22291,N_22255);
nor U22457 (N_22457,N_22344,N_22215);
and U22458 (N_22458,N_22240,N_22328);
nand U22459 (N_22459,N_22270,N_22308);
and U22460 (N_22460,N_22297,N_22369);
or U22461 (N_22461,N_22282,N_22247);
and U22462 (N_22462,N_22380,N_22281);
xor U22463 (N_22463,N_22248,N_22377);
and U22464 (N_22464,N_22227,N_22233);
nand U22465 (N_22465,N_22298,N_22239);
nand U22466 (N_22466,N_22260,N_22230);
xnor U22467 (N_22467,N_22387,N_22237);
nor U22468 (N_22468,N_22258,N_22378);
nand U22469 (N_22469,N_22398,N_22311);
or U22470 (N_22470,N_22262,N_22222);
nor U22471 (N_22471,N_22372,N_22205);
or U22472 (N_22472,N_22219,N_22269);
and U22473 (N_22473,N_22251,N_22208);
or U22474 (N_22474,N_22336,N_22221);
nand U22475 (N_22475,N_22292,N_22317);
or U22476 (N_22476,N_22347,N_22383);
nand U22477 (N_22477,N_22216,N_22288);
nor U22478 (N_22478,N_22345,N_22353);
nand U22479 (N_22479,N_22389,N_22250);
and U22480 (N_22480,N_22362,N_22368);
or U22481 (N_22481,N_22218,N_22279);
xnor U22482 (N_22482,N_22321,N_22373);
and U22483 (N_22483,N_22303,N_22246);
and U22484 (N_22484,N_22314,N_22229);
or U22485 (N_22485,N_22244,N_22352);
nor U22486 (N_22486,N_22364,N_22326);
xnor U22487 (N_22487,N_22382,N_22267);
or U22488 (N_22488,N_22232,N_22313);
xnor U22489 (N_22489,N_22367,N_22243);
and U22490 (N_22490,N_22331,N_22264);
nor U22491 (N_22491,N_22212,N_22299);
and U22492 (N_22492,N_22374,N_22286);
and U22493 (N_22493,N_22361,N_22334);
or U22494 (N_22494,N_22256,N_22268);
and U22495 (N_22495,N_22271,N_22366);
nor U22496 (N_22496,N_22325,N_22277);
nor U22497 (N_22497,N_22224,N_22302);
xnor U22498 (N_22498,N_22356,N_22306);
or U22499 (N_22499,N_22396,N_22289);
xor U22500 (N_22500,N_22234,N_22300);
or U22501 (N_22501,N_22369,N_22319);
xor U22502 (N_22502,N_22391,N_22251);
xor U22503 (N_22503,N_22210,N_22239);
nand U22504 (N_22504,N_22278,N_22221);
or U22505 (N_22505,N_22293,N_22315);
nand U22506 (N_22506,N_22213,N_22292);
xor U22507 (N_22507,N_22283,N_22350);
nor U22508 (N_22508,N_22397,N_22348);
nand U22509 (N_22509,N_22273,N_22314);
nand U22510 (N_22510,N_22323,N_22269);
nor U22511 (N_22511,N_22329,N_22291);
nand U22512 (N_22512,N_22352,N_22390);
xor U22513 (N_22513,N_22245,N_22258);
and U22514 (N_22514,N_22292,N_22268);
nor U22515 (N_22515,N_22322,N_22269);
nand U22516 (N_22516,N_22274,N_22263);
xnor U22517 (N_22517,N_22386,N_22255);
nand U22518 (N_22518,N_22252,N_22209);
nor U22519 (N_22519,N_22389,N_22280);
xnor U22520 (N_22520,N_22378,N_22248);
and U22521 (N_22521,N_22392,N_22214);
and U22522 (N_22522,N_22344,N_22285);
nand U22523 (N_22523,N_22254,N_22206);
or U22524 (N_22524,N_22221,N_22327);
nand U22525 (N_22525,N_22255,N_22202);
and U22526 (N_22526,N_22218,N_22243);
nor U22527 (N_22527,N_22335,N_22212);
xor U22528 (N_22528,N_22358,N_22284);
and U22529 (N_22529,N_22323,N_22392);
nand U22530 (N_22530,N_22329,N_22350);
nand U22531 (N_22531,N_22211,N_22352);
nand U22532 (N_22532,N_22229,N_22399);
and U22533 (N_22533,N_22322,N_22284);
nand U22534 (N_22534,N_22208,N_22392);
nand U22535 (N_22535,N_22367,N_22285);
nor U22536 (N_22536,N_22259,N_22295);
nand U22537 (N_22537,N_22218,N_22355);
nor U22538 (N_22538,N_22381,N_22367);
nand U22539 (N_22539,N_22370,N_22289);
and U22540 (N_22540,N_22227,N_22257);
nand U22541 (N_22541,N_22316,N_22279);
nand U22542 (N_22542,N_22313,N_22345);
nor U22543 (N_22543,N_22363,N_22306);
xor U22544 (N_22544,N_22382,N_22291);
xor U22545 (N_22545,N_22361,N_22220);
nor U22546 (N_22546,N_22209,N_22215);
or U22547 (N_22547,N_22315,N_22269);
or U22548 (N_22548,N_22333,N_22252);
nor U22549 (N_22549,N_22367,N_22234);
or U22550 (N_22550,N_22360,N_22251);
xnor U22551 (N_22551,N_22272,N_22298);
nand U22552 (N_22552,N_22392,N_22330);
xnor U22553 (N_22553,N_22344,N_22338);
or U22554 (N_22554,N_22341,N_22285);
nand U22555 (N_22555,N_22256,N_22381);
nor U22556 (N_22556,N_22361,N_22321);
xnor U22557 (N_22557,N_22373,N_22316);
nand U22558 (N_22558,N_22382,N_22289);
xor U22559 (N_22559,N_22303,N_22266);
nand U22560 (N_22560,N_22354,N_22350);
nand U22561 (N_22561,N_22204,N_22371);
nor U22562 (N_22562,N_22367,N_22284);
or U22563 (N_22563,N_22215,N_22361);
xnor U22564 (N_22564,N_22261,N_22349);
or U22565 (N_22565,N_22268,N_22329);
and U22566 (N_22566,N_22350,N_22252);
xor U22567 (N_22567,N_22395,N_22292);
nand U22568 (N_22568,N_22327,N_22204);
nand U22569 (N_22569,N_22266,N_22342);
nor U22570 (N_22570,N_22302,N_22375);
and U22571 (N_22571,N_22340,N_22250);
nor U22572 (N_22572,N_22323,N_22344);
nand U22573 (N_22573,N_22330,N_22361);
xnor U22574 (N_22574,N_22233,N_22232);
or U22575 (N_22575,N_22299,N_22309);
and U22576 (N_22576,N_22381,N_22328);
xor U22577 (N_22577,N_22239,N_22332);
nor U22578 (N_22578,N_22253,N_22329);
and U22579 (N_22579,N_22346,N_22366);
or U22580 (N_22580,N_22301,N_22389);
or U22581 (N_22581,N_22300,N_22373);
and U22582 (N_22582,N_22322,N_22326);
xnor U22583 (N_22583,N_22207,N_22300);
or U22584 (N_22584,N_22392,N_22331);
xnor U22585 (N_22585,N_22316,N_22342);
and U22586 (N_22586,N_22278,N_22290);
nand U22587 (N_22587,N_22363,N_22253);
nand U22588 (N_22588,N_22271,N_22215);
nand U22589 (N_22589,N_22309,N_22265);
nand U22590 (N_22590,N_22291,N_22289);
or U22591 (N_22591,N_22227,N_22258);
xnor U22592 (N_22592,N_22207,N_22294);
nand U22593 (N_22593,N_22247,N_22304);
or U22594 (N_22594,N_22321,N_22216);
nand U22595 (N_22595,N_22209,N_22376);
or U22596 (N_22596,N_22206,N_22244);
nor U22597 (N_22597,N_22244,N_22346);
xor U22598 (N_22598,N_22229,N_22204);
nand U22599 (N_22599,N_22317,N_22214);
xor U22600 (N_22600,N_22529,N_22447);
and U22601 (N_22601,N_22593,N_22523);
or U22602 (N_22602,N_22406,N_22528);
xor U22603 (N_22603,N_22589,N_22525);
or U22604 (N_22604,N_22400,N_22401);
xor U22605 (N_22605,N_22557,N_22452);
xor U22606 (N_22606,N_22503,N_22496);
nor U22607 (N_22607,N_22542,N_22515);
xor U22608 (N_22608,N_22538,N_22508);
and U22609 (N_22609,N_22552,N_22489);
or U22610 (N_22610,N_22514,N_22502);
or U22611 (N_22611,N_22449,N_22428);
nor U22612 (N_22612,N_22486,N_22591);
nand U22613 (N_22613,N_22582,N_22472);
and U22614 (N_22614,N_22580,N_22469);
nand U22615 (N_22615,N_22459,N_22468);
xnor U22616 (N_22616,N_22439,N_22554);
nor U22617 (N_22617,N_22539,N_22461);
nand U22618 (N_22618,N_22563,N_22540);
and U22619 (N_22619,N_22555,N_22446);
nand U22620 (N_22620,N_22596,N_22430);
xor U22621 (N_22621,N_22408,N_22403);
nor U22622 (N_22622,N_22465,N_22471);
and U22623 (N_22623,N_22498,N_22432);
and U22624 (N_22624,N_22442,N_22577);
nor U22625 (N_22625,N_22492,N_22588);
and U22626 (N_22626,N_22512,N_22586);
or U22627 (N_22627,N_22473,N_22445);
or U22628 (N_22628,N_22463,N_22526);
or U22629 (N_22629,N_22494,N_22487);
xnor U22630 (N_22630,N_22417,N_22553);
or U22631 (N_22631,N_22477,N_22569);
and U22632 (N_22632,N_22533,N_22575);
nand U22633 (N_22633,N_22592,N_22579);
xor U22634 (N_22634,N_22490,N_22506);
and U22635 (N_22635,N_22546,N_22545);
and U22636 (N_22636,N_22541,N_22427);
nand U22637 (N_22637,N_22424,N_22572);
and U22638 (N_22638,N_22462,N_22423);
or U22639 (N_22639,N_22455,N_22466);
xnor U22640 (N_22640,N_22426,N_22482);
or U22641 (N_22641,N_22532,N_22556);
xor U22642 (N_22642,N_22583,N_22561);
nor U22643 (N_22643,N_22510,N_22527);
nor U22644 (N_22644,N_22507,N_22504);
and U22645 (N_22645,N_22484,N_22571);
nor U22646 (N_22646,N_22500,N_22522);
and U22647 (N_22647,N_22438,N_22543);
xor U22648 (N_22648,N_22479,N_22505);
or U22649 (N_22649,N_22495,N_22414);
nor U22650 (N_22650,N_22488,N_22590);
or U22651 (N_22651,N_22568,N_22413);
and U22652 (N_22652,N_22458,N_22530);
and U22653 (N_22653,N_22535,N_22402);
xor U22654 (N_22654,N_22436,N_22520);
nor U22655 (N_22655,N_22464,N_22407);
and U22656 (N_22656,N_22470,N_22581);
nor U22657 (N_22657,N_22574,N_22444);
nand U22658 (N_22658,N_22480,N_22431);
xnor U22659 (N_22659,N_22567,N_22598);
and U22660 (N_22660,N_22564,N_22565);
nor U22661 (N_22661,N_22599,N_22421);
or U22662 (N_22662,N_22422,N_22474);
and U22663 (N_22663,N_22544,N_22405);
xor U22664 (N_22664,N_22493,N_22485);
xnor U22665 (N_22665,N_22476,N_22437);
or U22666 (N_22666,N_22456,N_22410);
nand U22667 (N_22667,N_22518,N_22429);
and U22668 (N_22668,N_22576,N_22451);
xnor U22669 (N_22669,N_22453,N_22570);
nand U22670 (N_22670,N_22549,N_22481);
xor U22671 (N_22671,N_22566,N_22483);
nand U22672 (N_22672,N_22560,N_22416);
and U22673 (N_22673,N_22516,N_22467);
xnor U22674 (N_22674,N_22578,N_22517);
xnor U22675 (N_22675,N_22534,N_22562);
or U22676 (N_22676,N_22411,N_22412);
nor U22677 (N_22677,N_22587,N_22450);
xnor U22678 (N_22678,N_22454,N_22478);
nor U22679 (N_22679,N_22448,N_22501);
or U22680 (N_22680,N_22597,N_22499);
or U22681 (N_22681,N_22460,N_22548);
or U22682 (N_22682,N_22475,N_22585);
xnor U22683 (N_22683,N_22511,N_22491);
nor U22684 (N_22684,N_22558,N_22584);
nand U22685 (N_22685,N_22441,N_22433);
nor U22686 (N_22686,N_22547,N_22415);
nand U22687 (N_22687,N_22443,N_22509);
nand U22688 (N_22688,N_22531,N_22513);
nor U22689 (N_22689,N_22409,N_22420);
nand U22690 (N_22690,N_22425,N_22497);
nor U22691 (N_22691,N_22550,N_22595);
xor U22692 (N_22692,N_22519,N_22524);
and U22693 (N_22693,N_22559,N_22594);
and U22694 (N_22694,N_22404,N_22536);
and U22695 (N_22695,N_22435,N_22434);
or U22696 (N_22696,N_22537,N_22521);
and U22697 (N_22697,N_22418,N_22440);
nand U22698 (N_22698,N_22419,N_22457);
or U22699 (N_22699,N_22573,N_22551);
xor U22700 (N_22700,N_22533,N_22545);
xor U22701 (N_22701,N_22424,N_22422);
nor U22702 (N_22702,N_22418,N_22495);
nor U22703 (N_22703,N_22507,N_22454);
or U22704 (N_22704,N_22417,N_22412);
nand U22705 (N_22705,N_22477,N_22558);
xnor U22706 (N_22706,N_22441,N_22406);
nor U22707 (N_22707,N_22502,N_22558);
and U22708 (N_22708,N_22411,N_22566);
xnor U22709 (N_22709,N_22417,N_22481);
and U22710 (N_22710,N_22535,N_22561);
xnor U22711 (N_22711,N_22579,N_22587);
xnor U22712 (N_22712,N_22536,N_22457);
nand U22713 (N_22713,N_22590,N_22408);
nor U22714 (N_22714,N_22522,N_22593);
and U22715 (N_22715,N_22419,N_22594);
xnor U22716 (N_22716,N_22576,N_22442);
and U22717 (N_22717,N_22426,N_22445);
and U22718 (N_22718,N_22497,N_22547);
and U22719 (N_22719,N_22464,N_22412);
nor U22720 (N_22720,N_22491,N_22408);
xnor U22721 (N_22721,N_22453,N_22510);
xnor U22722 (N_22722,N_22403,N_22404);
nor U22723 (N_22723,N_22442,N_22453);
and U22724 (N_22724,N_22471,N_22474);
or U22725 (N_22725,N_22462,N_22485);
nor U22726 (N_22726,N_22415,N_22491);
or U22727 (N_22727,N_22509,N_22506);
nand U22728 (N_22728,N_22464,N_22506);
or U22729 (N_22729,N_22412,N_22408);
or U22730 (N_22730,N_22440,N_22564);
and U22731 (N_22731,N_22514,N_22580);
and U22732 (N_22732,N_22439,N_22450);
xnor U22733 (N_22733,N_22422,N_22457);
xor U22734 (N_22734,N_22541,N_22417);
and U22735 (N_22735,N_22434,N_22451);
xor U22736 (N_22736,N_22538,N_22468);
xnor U22737 (N_22737,N_22509,N_22407);
xnor U22738 (N_22738,N_22552,N_22426);
or U22739 (N_22739,N_22480,N_22425);
nor U22740 (N_22740,N_22469,N_22576);
nand U22741 (N_22741,N_22569,N_22451);
nor U22742 (N_22742,N_22455,N_22547);
and U22743 (N_22743,N_22488,N_22594);
and U22744 (N_22744,N_22485,N_22463);
and U22745 (N_22745,N_22500,N_22489);
nor U22746 (N_22746,N_22508,N_22522);
nand U22747 (N_22747,N_22497,N_22455);
nor U22748 (N_22748,N_22470,N_22418);
xor U22749 (N_22749,N_22524,N_22569);
nand U22750 (N_22750,N_22566,N_22451);
nand U22751 (N_22751,N_22450,N_22536);
nor U22752 (N_22752,N_22512,N_22455);
nor U22753 (N_22753,N_22487,N_22593);
nor U22754 (N_22754,N_22450,N_22472);
or U22755 (N_22755,N_22461,N_22523);
or U22756 (N_22756,N_22544,N_22425);
nor U22757 (N_22757,N_22586,N_22593);
and U22758 (N_22758,N_22553,N_22419);
and U22759 (N_22759,N_22528,N_22484);
or U22760 (N_22760,N_22520,N_22426);
xor U22761 (N_22761,N_22594,N_22574);
or U22762 (N_22762,N_22491,N_22595);
xor U22763 (N_22763,N_22576,N_22564);
or U22764 (N_22764,N_22494,N_22404);
xnor U22765 (N_22765,N_22496,N_22458);
xor U22766 (N_22766,N_22453,N_22446);
nand U22767 (N_22767,N_22549,N_22512);
nor U22768 (N_22768,N_22567,N_22413);
and U22769 (N_22769,N_22501,N_22462);
xnor U22770 (N_22770,N_22412,N_22586);
nand U22771 (N_22771,N_22559,N_22497);
nand U22772 (N_22772,N_22564,N_22446);
and U22773 (N_22773,N_22465,N_22409);
and U22774 (N_22774,N_22593,N_22434);
xnor U22775 (N_22775,N_22549,N_22592);
or U22776 (N_22776,N_22484,N_22550);
xnor U22777 (N_22777,N_22520,N_22526);
nand U22778 (N_22778,N_22558,N_22461);
or U22779 (N_22779,N_22439,N_22505);
nor U22780 (N_22780,N_22588,N_22528);
and U22781 (N_22781,N_22540,N_22586);
nor U22782 (N_22782,N_22581,N_22483);
xnor U22783 (N_22783,N_22563,N_22537);
nand U22784 (N_22784,N_22495,N_22569);
nor U22785 (N_22785,N_22405,N_22582);
nand U22786 (N_22786,N_22423,N_22526);
nand U22787 (N_22787,N_22494,N_22470);
or U22788 (N_22788,N_22585,N_22442);
or U22789 (N_22789,N_22550,N_22483);
nor U22790 (N_22790,N_22548,N_22511);
xnor U22791 (N_22791,N_22509,N_22530);
or U22792 (N_22792,N_22560,N_22577);
or U22793 (N_22793,N_22536,N_22420);
xnor U22794 (N_22794,N_22582,N_22525);
nand U22795 (N_22795,N_22468,N_22522);
xor U22796 (N_22796,N_22549,N_22566);
xor U22797 (N_22797,N_22553,N_22577);
and U22798 (N_22798,N_22534,N_22479);
xor U22799 (N_22799,N_22573,N_22450);
nor U22800 (N_22800,N_22764,N_22777);
and U22801 (N_22801,N_22791,N_22720);
or U22802 (N_22802,N_22774,N_22625);
or U22803 (N_22803,N_22716,N_22704);
xnor U22804 (N_22804,N_22645,N_22708);
nor U22805 (N_22805,N_22613,N_22780);
nand U22806 (N_22806,N_22799,N_22741);
nand U22807 (N_22807,N_22680,N_22734);
xnor U22808 (N_22808,N_22711,N_22695);
nor U22809 (N_22809,N_22767,N_22631);
and U22810 (N_22810,N_22601,N_22758);
or U22811 (N_22811,N_22713,N_22697);
nand U22812 (N_22812,N_22615,N_22635);
xor U22813 (N_22813,N_22640,N_22740);
xor U22814 (N_22814,N_22678,N_22687);
xnor U22815 (N_22815,N_22779,N_22626);
nand U22816 (N_22816,N_22651,N_22657);
and U22817 (N_22817,N_22775,N_22796);
xnor U22818 (N_22818,N_22795,N_22628);
nor U22819 (N_22819,N_22658,N_22709);
and U22820 (N_22820,N_22637,N_22676);
nand U22821 (N_22821,N_22743,N_22660);
or U22822 (N_22822,N_22632,N_22792);
and U22823 (N_22823,N_22689,N_22798);
and U22824 (N_22824,N_22617,N_22702);
xnor U22825 (N_22825,N_22733,N_22683);
nor U22826 (N_22826,N_22725,N_22655);
nand U22827 (N_22827,N_22784,N_22608);
nor U22828 (N_22828,N_22662,N_22664);
or U22829 (N_22829,N_22648,N_22751);
nand U22830 (N_22830,N_22790,N_22673);
xnor U22831 (N_22831,N_22794,N_22686);
and U22832 (N_22832,N_22739,N_22762);
nand U22833 (N_22833,N_22752,N_22726);
nand U22834 (N_22834,N_22723,N_22641);
or U22835 (N_22835,N_22624,N_22787);
xnor U22836 (N_22836,N_22778,N_22724);
nand U22837 (N_22837,N_22756,N_22736);
and U22838 (N_22838,N_22682,N_22776);
and U22839 (N_22839,N_22769,N_22643);
nor U22840 (N_22840,N_22620,N_22692);
or U22841 (N_22841,N_22735,N_22715);
or U22842 (N_22842,N_22714,N_22621);
nor U22843 (N_22843,N_22750,N_22732);
or U22844 (N_22844,N_22604,N_22674);
or U22845 (N_22845,N_22647,N_22694);
xor U22846 (N_22846,N_22610,N_22696);
and U22847 (N_22847,N_22705,N_22727);
and U22848 (N_22848,N_22654,N_22688);
nand U22849 (N_22849,N_22761,N_22738);
and U22850 (N_22850,N_22669,N_22785);
and U22851 (N_22851,N_22656,N_22719);
xor U22852 (N_22852,N_22759,N_22611);
and U22853 (N_22853,N_22786,N_22665);
nand U22854 (N_22854,N_22731,N_22685);
and U22855 (N_22855,N_22793,N_22693);
nor U22856 (N_22856,N_22710,N_22772);
nor U22857 (N_22857,N_22707,N_22609);
or U22858 (N_22858,N_22712,N_22753);
xnor U22859 (N_22859,N_22700,N_22630);
xor U22860 (N_22860,N_22763,N_22638);
or U22861 (N_22861,N_22745,N_22627);
nand U22862 (N_22862,N_22771,N_22757);
nand U22863 (N_22863,N_22639,N_22633);
nand U22864 (N_22864,N_22766,N_22679);
nor U22865 (N_22865,N_22797,N_22703);
or U22866 (N_22866,N_22644,N_22607);
and U22867 (N_22867,N_22622,N_22783);
nand U22868 (N_22868,N_22650,N_22698);
nor U22869 (N_22869,N_22649,N_22749);
xor U22870 (N_22870,N_22642,N_22754);
and U22871 (N_22871,N_22614,N_22619);
xnor U22872 (N_22872,N_22652,N_22768);
xnor U22873 (N_22873,N_22653,N_22742);
or U22874 (N_22874,N_22606,N_22663);
and U22875 (N_22875,N_22646,N_22717);
nor U22876 (N_22876,N_22721,N_22684);
nor U22877 (N_22877,N_22661,N_22765);
nand U22878 (N_22878,N_22782,N_22618);
and U22879 (N_22879,N_22755,N_22773);
xnor U22880 (N_22880,N_22629,N_22701);
xor U22881 (N_22881,N_22722,N_22681);
nor U22882 (N_22882,N_22677,N_22728);
nand U22883 (N_22883,N_22760,N_22675);
and U22884 (N_22884,N_22788,N_22666);
and U22885 (N_22885,N_22667,N_22668);
nor U22886 (N_22886,N_22671,N_22706);
or U22887 (N_22887,N_22690,N_22602);
or U22888 (N_22888,N_22672,N_22748);
xnor U22889 (N_22889,N_22612,N_22781);
nand U22890 (N_22890,N_22603,N_22770);
nor U22891 (N_22891,N_22737,N_22746);
xor U22892 (N_22892,N_22699,N_22729);
xor U22893 (N_22893,N_22691,N_22605);
nand U22894 (N_22894,N_22747,N_22634);
xor U22895 (N_22895,N_22600,N_22659);
nor U22896 (N_22896,N_22789,N_22636);
nor U22897 (N_22897,N_22744,N_22616);
or U22898 (N_22898,N_22623,N_22670);
or U22899 (N_22899,N_22718,N_22730);
nor U22900 (N_22900,N_22793,N_22704);
nor U22901 (N_22901,N_22756,N_22658);
nor U22902 (N_22902,N_22670,N_22619);
and U22903 (N_22903,N_22640,N_22763);
or U22904 (N_22904,N_22779,N_22770);
or U22905 (N_22905,N_22606,N_22797);
xor U22906 (N_22906,N_22637,N_22631);
and U22907 (N_22907,N_22764,N_22667);
nand U22908 (N_22908,N_22797,N_22682);
or U22909 (N_22909,N_22738,N_22684);
nand U22910 (N_22910,N_22711,N_22686);
nor U22911 (N_22911,N_22673,N_22727);
xor U22912 (N_22912,N_22793,N_22629);
nor U22913 (N_22913,N_22651,N_22724);
nor U22914 (N_22914,N_22758,N_22642);
and U22915 (N_22915,N_22636,N_22610);
and U22916 (N_22916,N_22622,N_22718);
xor U22917 (N_22917,N_22743,N_22618);
nor U22918 (N_22918,N_22746,N_22638);
and U22919 (N_22919,N_22665,N_22791);
nor U22920 (N_22920,N_22728,N_22647);
nand U22921 (N_22921,N_22738,N_22653);
or U22922 (N_22922,N_22747,N_22688);
nand U22923 (N_22923,N_22772,N_22630);
or U22924 (N_22924,N_22694,N_22601);
and U22925 (N_22925,N_22653,N_22753);
and U22926 (N_22926,N_22640,N_22758);
and U22927 (N_22927,N_22769,N_22792);
nor U22928 (N_22928,N_22732,N_22698);
xnor U22929 (N_22929,N_22743,N_22669);
xnor U22930 (N_22930,N_22778,N_22712);
xnor U22931 (N_22931,N_22625,N_22756);
nor U22932 (N_22932,N_22662,N_22749);
or U22933 (N_22933,N_22702,N_22715);
nor U22934 (N_22934,N_22710,N_22762);
nor U22935 (N_22935,N_22798,N_22765);
nor U22936 (N_22936,N_22691,N_22724);
xnor U22937 (N_22937,N_22733,N_22773);
and U22938 (N_22938,N_22770,N_22726);
and U22939 (N_22939,N_22726,N_22795);
xor U22940 (N_22940,N_22679,N_22648);
or U22941 (N_22941,N_22610,N_22776);
nand U22942 (N_22942,N_22796,N_22687);
or U22943 (N_22943,N_22754,N_22669);
nor U22944 (N_22944,N_22745,N_22747);
nand U22945 (N_22945,N_22684,N_22604);
xnor U22946 (N_22946,N_22669,N_22748);
or U22947 (N_22947,N_22651,N_22632);
nand U22948 (N_22948,N_22644,N_22751);
or U22949 (N_22949,N_22634,N_22629);
xnor U22950 (N_22950,N_22760,N_22791);
xor U22951 (N_22951,N_22732,N_22668);
nor U22952 (N_22952,N_22639,N_22647);
and U22953 (N_22953,N_22697,N_22668);
nand U22954 (N_22954,N_22727,N_22742);
and U22955 (N_22955,N_22727,N_22717);
nor U22956 (N_22956,N_22614,N_22662);
and U22957 (N_22957,N_22634,N_22669);
or U22958 (N_22958,N_22704,N_22675);
nand U22959 (N_22959,N_22704,N_22739);
nor U22960 (N_22960,N_22749,N_22708);
or U22961 (N_22961,N_22680,N_22673);
or U22962 (N_22962,N_22774,N_22758);
and U22963 (N_22963,N_22728,N_22655);
xnor U22964 (N_22964,N_22700,N_22715);
nand U22965 (N_22965,N_22698,N_22701);
or U22966 (N_22966,N_22724,N_22736);
or U22967 (N_22967,N_22629,N_22685);
nor U22968 (N_22968,N_22764,N_22746);
and U22969 (N_22969,N_22757,N_22684);
and U22970 (N_22970,N_22650,N_22651);
and U22971 (N_22971,N_22770,N_22784);
nor U22972 (N_22972,N_22675,N_22668);
or U22973 (N_22973,N_22780,N_22668);
nor U22974 (N_22974,N_22650,N_22677);
nor U22975 (N_22975,N_22630,N_22774);
and U22976 (N_22976,N_22773,N_22797);
xor U22977 (N_22977,N_22785,N_22624);
xor U22978 (N_22978,N_22799,N_22743);
nand U22979 (N_22979,N_22737,N_22660);
nand U22980 (N_22980,N_22700,N_22791);
and U22981 (N_22981,N_22774,N_22714);
nor U22982 (N_22982,N_22705,N_22614);
and U22983 (N_22983,N_22728,N_22752);
or U22984 (N_22984,N_22604,N_22754);
or U22985 (N_22985,N_22780,N_22734);
or U22986 (N_22986,N_22719,N_22686);
or U22987 (N_22987,N_22750,N_22656);
xor U22988 (N_22988,N_22715,N_22658);
and U22989 (N_22989,N_22788,N_22736);
and U22990 (N_22990,N_22677,N_22611);
and U22991 (N_22991,N_22697,N_22638);
or U22992 (N_22992,N_22704,N_22760);
or U22993 (N_22993,N_22709,N_22713);
nand U22994 (N_22994,N_22642,N_22738);
nand U22995 (N_22995,N_22737,N_22717);
and U22996 (N_22996,N_22707,N_22783);
nor U22997 (N_22997,N_22632,N_22708);
nand U22998 (N_22998,N_22641,N_22660);
nor U22999 (N_22999,N_22641,N_22733);
xor U23000 (N_23000,N_22823,N_22964);
and U23001 (N_23001,N_22839,N_22932);
or U23002 (N_23002,N_22901,N_22885);
nor U23003 (N_23003,N_22939,N_22894);
or U23004 (N_23004,N_22959,N_22911);
nand U23005 (N_23005,N_22877,N_22899);
or U23006 (N_23006,N_22814,N_22929);
or U23007 (N_23007,N_22968,N_22847);
nand U23008 (N_23008,N_22937,N_22888);
nor U23009 (N_23009,N_22897,N_22851);
or U23010 (N_23010,N_22913,N_22846);
or U23011 (N_23011,N_22994,N_22955);
nand U23012 (N_23012,N_22902,N_22821);
nor U23013 (N_23013,N_22996,N_22870);
xor U23014 (N_23014,N_22872,N_22834);
nor U23015 (N_23015,N_22944,N_22855);
nand U23016 (N_23016,N_22815,N_22950);
nand U23017 (N_23017,N_22984,N_22988);
or U23018 (N_23018,N_22809,N_22912);
nor U23019 (N_23019,N_22827,N_22945);
and U23020 (N_23020,N_22975,N_22930);
nor U23021 (N_23021,N_22942,N_22801);
or U23022 (N_23022,N_22933,N_22845);
xnor U23023 (N_23023,N_22841,N_22893);
nand U23024 (N_23024,N_22992,N_22892);
xnor U23025 (N_23025,N_22931,N_22832);
nor U23026 (N_23026,N_22824,N_22878);
nor U23027 (N_23027,N_22866,N_22938);
xor U23028 (N_23028,N_22915,N_22914);
xor U23029 (N_23029,N_22922,N_22977);
nor U23030 (N_23030,N_22907,N_22880);
xor U23031 (N_23031,N_22807,N_22919);
and U23032 (N_23032,N_22863,N_22825);
or U23033 (N_23033,N_22802,N_22963);
nand U23034 (N_23034,N_22848,N_22812);
and U23035 (N_23035,N_22829,N_22856);
and U23036 (N_23036,N_22983,N_22859);
nand U23037 (N_23037,N_22862,N_22917);
or U23038 (N_23038,N_22954,N_22895);
or U23039 (N_23039,N_22987,N_22966);
nand U23040 (N_23040,N_22886,N_22943);
nand U23041 (N_23041,N_22905,N_22949);
nand U23042 (N_23042,N_22813,N_22879);
or U23043 (N_23043,N_22948,N_22806);
or U23044 (N_23044,N_22852,N_22820);
and U23045 (N_23045,N_22810,N_22920);
and U23046 (N_23046,N_22916,N_22926);
nand U23047 (N_23047,N_22969,N_22836);
nand U23048 (N_23048,N_22860,N_22858);
or U23049 (N_23049,N_22921,N_22874);
or U23050 (N_23050,N_22924,N_22993);
nor U23051 (N_23051,N_22881,N_22904);
and U23052 (N_23052,N_22854,N_22818);
or U23053 (N_23053,N_22960,N_22837);
or U23054 (N_23054,N_22971,N_22889);
xnor U23055 (N_23055,N_22972,N_22869);
or U23056 (N_23056,N_22936,N_22967);
nor U23057 (N_23057,N_22838,N_22828);
and U23058 (N_23058,N_22898,N_22927);
xor U23059 (N_23059,N_22840,N_22952);
nor U23060 (N_23060,N_22982,N_22816);
nand U23061 (N_23061,N_22962,N_22961);
nor U23062 (N_23062,N_22998,N_22946);
xnor U23063 (N_23063,N_22951,N_22953);
and U23064 (N_23064,N_22999,N_22903);
xnor U23065 (N_23065,N_22803,N_22910);
xnor U23066 (N_23066,N_22857,N_22986);
or U23067 (N_23067,N_22864,N_22918);
nor U23068 (N_23068,N_22883,N_22844);
or U23069 (N_23069,N_22978,N_22976);
xnor U23070 (N_23070,N_22991,N_22835);
nand U23071 (N_23071,N_22884,N_22842);
nand U23072 (N_23072,N_22887,N_22867);
and U23073 (N_23073,N_22906,N_22853);
xnor U23074 (N_23074,N_22980,N_22850);
and U23075 (N_23075,N_22882,N_22896);
or U23076 (N_23076,N_22811,N_22979);
nand U23077 (N_23077,N_22956,N_22941);
and U23078 (N_23078,N_22805,N_22958);
and U23079 (N_23079,N_22819,N_22876);
or U23080 (N_23080,N_22990,N_22833);
nand U23081 (N_23081,N_22947,N_22830);
or U23082 (N_23082,N_22973,N_22974);
nor U23083 (N_23083,N_22826,N_22940);
and U23084 (N_23084,N_22923,N_22865);
nor U23085 (N_23085,N_22800,N_22985);
or U23086 (N_23086,N_22970,N_22934);
nor U23087 (N_23087,N_22843,N_22935);
nand U23088 (N_23088,N_22831,N_22995);
xor U23089 (N_23089,N_22891,N_22900);
xor U23090 (N_23090,N_22981,N_22817);
nor U23091 (N_23091,N_22804,N_22909);
nor U23092 (N_23092,N_22808,N_22849);
nor U23093 (N_23093,N_22868,N_22925);
xnor U23094 (N_23094,N_22871,N_22822);
nor U23095 (N_23095,N_22908,N_22875);
nor U23096 (N_23096,N_22861,N_22957);
nor U23097 (N_23097,N_22873,N_22965);
xor U23098 (N_23098,N_22997,N_22890);
and U23099 (N_23099,N_22928,N_22989);
or U23100 (N_23100,N_22803,N_22903);
and U23101 (N_23101,N_22822,N_22924);
nand U23102 (N_23102,N_22868,N_22811);
nand U23103 (N_23103,N_22896,N_22930);
nor U23104 (N_23104,N_22826,N_22978);
or U23105 (N_23105,N_22910,N_22930);
nand U23106 (N_23106,N_22989,N_22889);
nor U23107 (N_23107,N_22821,N_22940);
xor U23108 (N_23108,N_22930,N_22949);
and U23109 (N_23109,N_22866,N_22990);
xnor U23110 (N_23110,N_22878,N_22924);
and U23111 (N_23111,N_22943,N_22856);
nand U23112 (N_23112,N_22846,N_22883);
nand U23113 (N_23113,N_22835,N_22997);
and U23114 (N_23114,N_22925,N_22949);
and U23115 (N_23115,N_22996,N_22983);
or U23116 (N_23116,N_22936,N_22812);
or U23117 (N_23117,N_22868,N_22901);
nand U23118 (N_23118,N_22925,N_22887);
or U23119 (N_23119,N_22962,N_22846);
nand U23120 (N_23120,N_22957,N_22981);
or U23121 (N_23121,N_22903,N_22830);
or U23122 (N_23122,N_22911,N_22832);
or U23123 (N_23123,N_22975,N_22934);
and U23124 (N_23124,N_22929,N_22917);
or U23125 (N_23125,N_22818,N_22943);
nor U23126 (N_23126,N_22818,N_22835);
and U23127 (N_23127,N_22868,N_22977);
or U23128 (N_23128,N_22875,N_22963);
nand U23129 (N_23129,N_22966,N_22841);
or U23130 (N_23130,N_22908,N_22895);
nand U23131 (N_23131,N_22966,N_22852);
and U23132 (N_23132,N_22889,N_22895);
nand U23133 (N_23133,N_22804,N_22939);
nor U23134 (N_23134,N_22859,N_22867);
and U23135 (N_23135,N_22866,N_22818);
or U23136 (N_23136,N_22956,N_22804);
nand U23137 (N_23137,N_22832,N_22880);
and U23138 (N_23138,N_22820,N_22808);
nor U23139 (N_23139,N_22957,N_22970);
xor U23140 (N_23140,N_22916,N_22830);
or U23141 (N_23141,N_22892,N_22901);
nand U23142 (N_23142,N_22978,N_22809);
nor U23143 (N_23143,N_22861,N_22923);
and U23144 (N_23144,N_22867,N_22943);
and U23145 (N_23145,N_22856,N_22818);
nor U23146 (N_23146,N_22876,N_22899);
xnor U23147 (N_23147,N_22921,N_22858);
nand U23148 (N_23148,N_22896,N_22999);
nor U23149 (N_23149,N_22887,N_22929);
and U23150 (N_23150,N_22911,N_22920);
nand U23151 (N_23151,N_22950,N_22958);
nor U23152 (N_23152,N_22994,N_22878);
or U23153 (N_23153,N_22848,N_22860);
xnor U23154 (N_23154,N_22802,N_22876);
and U23155 (N_23155,N_22875,N_22867);
xor U23156 (N_23156,N_22956,N_22859);
and U23157 (N_23157,N_22963,N_22987);
xor U23158 (N_23158,N_22812,N_22915);
nor U23159 (N_23159,N_22848,N_22855);
or U23160 (N_23160,N_22836,N_22952);
nor U23161 (N_23161,N_22894,N_22827);
or U23162 (N_23162,N_22951,N_22993);
xor U23163 (N_23163,N_22976,N_22942);
and U23164 (N_23164,N_22975,N_22827);
nor U23165 (N_23165,N_22893,N_22909);
xnor U23166 (N_23166,N_22838,N_22898);
and U23167 (N_23167,N_22956,N_22979);
nand U23168 (N_23168,N_22973,N_22939);
xor U23169 (N_23169,N_22813,N_22966);
or U23170 (N_23170,N_22872,N_22978);
nand U23171 (N_23171,N_22931,N_22916);
nor U23172 (N_23172,N_22926,N_22871);
xnor U23173 (N_23173,N_22811,N_22949);
xnor U23174 (N_23174,N_22975,N_22900);
and U23175 (N_23175,N_22901,N_22926);
and U23176 (N_23176,N_22816,N_22907);
nand U23177 (N_23177,N_22971,N_22805);
nand U23178 (N_23178,N_22820,N_22913);
nor U23179 (N_23179,N_22931,N_22947);
xor U23180 (N_23180,N_22941,N_22837);
or U23181 (N_23181,N_22807,N_22969);
or U23182 (N_23182,N_22866,N_22912);
xor U23183 (N_23183,N_22919,N_22827);
nor U23184 (N_23184,N_22995,N_22804);
and U23185 (N_23185,N_22869,N_22949);
and U23186 (N_23186,N_22815,N_22858);
nor U23187 (N_23187,N_22860,N_22914);
nor U23188 (N_23188,N_22982,N_22875);
or U23189 (N_23189,N_22981,N_22848);
and U23190 (N_23190,N_22844,N_22928);
and U23191 (N_23191,N_22824,N_22811);
nand U23192 (N_23192,N_22903,N_22872);
or U23193 (N_23193,N_22914,N_22972);
nor U23194 (N_23194,N_22982,N_22936);
or U23195 (N_23195,N_22920,N_22941);
or U23196 (N_23196,N_22839,N_22824);
xnor U23197 (N_23197,N_22994,N_22802);
and U23198 (N_23198,N_22977,N_22894);
and U23199 (N_23199,N_22944,N_22888);
and U23200 (N_23200,N_23037,N_23187);
xnor U23201 (N_23201,N_23023,N_23118);
and U23202 (N_23202,N_23174,N_23103);
xnor U23203 (N_23203,N_23102,N_23036);
nand U23204 (N_23204,N_23098,N_23123);
or U23205 (N_23205,N_23015,N_23128);
nor U23206 (N_23206,N_23010,N_23061);
nand U23207 (N_23207,N_23063,N_23134);
nand U23208 (N_23208,N_23044,N_23022);
xnor U23209 (N_23209,N_23009,N_23129);
or U23210 (N_23210,N_23004,N_23085);
xnor U23211 (N_23211,N_23016,N_23100);
xor U23212 (N_23212,N_23127,N_23124);
nor U23213 (N_23213,N_23165,N_23158);
xnor U23214 (N_23214,N_23183,N_23067);
nand U23215 (N_23215,N_23006,N_23079);
or U23216 (N_23216,N_23189,N_23081);
nor U23217 (N_23217,N_23088,N_23177);
and U23218 (N_23218,N_23047,N_23068);
or U23219 (N_23219,N_23052,N_23139);
nand U23220 (N_23220,N_23001,N_23126);
and U23221 (N_23221,N_23198,N_23115);
xnor U23222 (N_23222,N_23039,N_23024);
nand U23223 (N_23223,N_23005,N_23030);
nor U23224 (N_23224,N_23179,N_23144);
xnor U23225 (N_23225,N_23025,N_23114);
nand U23226 (N_23226,N_23190,N_23097);
xor U23227 (N_23227,N_23073,N_23192);
and U23228 (N_23228,N_23056,N_23136);
nand U23229 (N_23229,N_23096,N_23194);
nor U23230 (N_23230,N_23132,N_23191);
nand U23231 (N_23231,N_23125,N_23035);
xor U23232 (N_23232,N_23172,N_23029);
or U23233 (N_23233,N_23093,N_23094);
nand U23234 (N_23234,N_23046,N_23116);
nand U23235 (N_23235,N_23113,N_23012);
xnor U23236 (N_23236,N_23048,N_23184);
xor U23237 (N_23237,N_23185,N_23146);
nand U23238 (N_23238,N_23182,N_23060);
nor U23239 (N_23239,N_23087,N_23041);
nor U23240 (N_23240,N_23164,N_23080);
nor U23241 (N_23241,N_23059,N_23049);
or U23242 (N_23242,N_23178,N_23138);
nor U23243 (N_23243,N_23149,N_23090);
and U23244 (N_23244,N_23042,N_23021);
nor U23245 (N_23245,N_23122,N_23065);
nand U23246 (N_23246,N_23107,N_23014);
nand U23247 (N_23247,N_23167,N_23175);
and U23248 (N_23248,N_23109,N_23104);
nand U23249 (N_23249,N_23193,N_23147);
nor U23250 (N_23250,N_23101,N_23045);
nand U23251 (N_23251,N_23083,N_23160);
nand U23252 (N_23252,N_23033,N_23020);
xor U23253 (N_23253,N_23150,N_23055);
xnor U23254 (N_23254,N_23195,N_23130);
xor U23255 (N_23255,N_23121,N_23008);
or U23256 (N_23256,N_23075,N_23017);
or U23257 (N_23257,N_23141,N_23027);
nand U23258 (N_23258,N_23084,N_23119);
nand U23259 (N_23259,N_23013,N_23091);
nor U23260 (N_23260,N_23169,N_23162);
or U23261 (N_23261,N_23082,N_23040);
nor U23262 (N_23262,N_23011,N_23117);
or U23263 (N_23263,N_23066,N_23142);
or U23264 (N_23264,N_23070,N_23181);
or U23265 (N_23265,N_23007,N_23180);
nor U23266 (N_23266,N_23199,N_23161);
and U23267 (N_23267,N_23077,N_23086);
and U23268 (N_23268,N_23176,N_23153);
and U23269 (N_23269,N_23069,N_23131);
and U23270 (N_23270,N_23018,N_23143);
nand U23271 (N_23271,N_23038,N_23188);
nand U23272 (N_23272,N_23051,N_23032);
and U23273 (N_23273,N_23071,N_23111);
and U23274 (N_23274,N_23028,N_23050);
xor U23275 (N_23275,N_23057,N_23031);
and U23276 (N_23276,N_23151,N_23196);
nand U23277 (N_23277,N_23135,N_23078);
xor U23278 (N_23278,N_23034,N_23043);
or U23279 (N_23279,N_23154,N_23053);
xnor U23280 (N_23280,N_23019,N_23095);
nor U23281 (N_23281,N_23133,N_23062);
nor U23282 (N_23282,N_23173,N_23058);
xor U23283 (N_23283,N_23163,N_23076);
nand U23284 (N_23284,N_23148,N_23140);
nor U23285 (N_23285,N_23152,N_23000);
and U23286 (N_23286,N_23074,N_23072);
or U23287 (N_23287,N_23003,N_23157);
or U23288 (N_23288,N_23106,N_23092);
nor U23289 (N_23289,N_23108,N_23026);
nand U23290 (N_23290,N_23168,N_23155);
or U23291 (N_23291,N_23197,N_23171);
or U23292 (N_23292,N_23112,N_23054);
or U23293 (N_23293,N_23002,N_23186);
and U23294 (N_23294,N_23159,N_23166);
nor U23295 (N_23295,N_23105,N_23137);
nor U23296 (N_23296,N_23120,N_23156);
xnor U23297 (N_23297,N_23170,N_23064);
xor U23298 (N_23298,N_23145,N_23089);
xor U23299 (N_23299,N_23110,N_23099);
nor U23300 (N_23300,N_23068,N_23146);
and U23301 (N_23301,N_23034,N_23119);
nand U23302 (N_23302,N_23049,N_23005);
and U23303 (N_23303,N_23193,N_23166);
or U23304 (N_23304,N_23139,N_23043);
nor U23305 (N_23305,N_23031,N_23053);
nor U23306 (N_23306,N_23023,N_23111);
nor U23307 (N_23307,N_23197,N_23129);
or U23308 (N_23308,N_23033,N_23081);
nand U23309 (N_23309,N_23075,N_23175);
nand U23310 (N_23310,N_23177,N_23173);
nand U23311 (N_23311,N_23176,N_23185);
and U23312 (N_23312,N_23051,N_23187);
nand U23313 (N_23313,N_23016,N_23133);
or U23314 (N_23314,N_23192,N_23115);
xor U23315 (N_23315,N_23167,N_23042);
xnor U23316 (N_23316,N_23112,N_23067);
or U23317 (N_23317,N_23081,N_23097);
and U23318 (N_23318,N_23187,N_23192);
xnor U23319 (N_23319,N_23153,N_23102);
nor U23320 (N_23320,N_23161,N_23104);
nor U23321 (N_23321,N_23055,N_23192);
or U23322 (N_23322,N_23101,N_23097);
nand U23323 (N_23323,N_23180,N_23126);
nand U23324 (N_23324,N_23177,N_23130);
xor U23325 (N_23325,N_23159,N_23066);
xor U23326 (N_23326,N_23098,N_23044);
or U23327 (N_23327,N_23140,N_23004);
nand U23328 (N_23328,N_23071,N_23042);
nand U23329 (N_23329,N_23142,N_23005);
and U23330 (N_23330,N_23154,N_23001);
or U23331 (N_23331,N_23179,N_23195);
nand U23332 (N_23332,N_23031,N_23141);
nand U23333 (N_23333,N_23128,N_23063);
xnor U23334 (N_23334,N_23112,N_23187);
xnor U23335 (N_23335,N_23068,N_23086);
nand U23336 (N_23336,N_23180,N_23116);
or U23337 (N_23337,N_23190,N_23157);
or U23338 (N_23338,N_23028,N_23188);
nand U23339 (N_23339,N_23056,N_23152);
xnor U23340 (N_23340,N_23082,N_23053);
or U23341 (N_23341,N_23168,N_23058);
or U23342 (N_23342,N_23034,N_23130);
xnor U23343 (N_23343,N_23095,N_23132);
or U23344 (N_23344,N_23187,N_23030);
xnor U23345 (N_23345,N_23065,N_23121);
or U23346 (N_23346,N_23145,N_23066);
nand U23347 (N_23347,N_23009,N_23078);
and U23348 (N_23348,N_23098,N_23002);
nor U23349 (N_23349,N_23089,N_23050);
nand U23350 (N_23350,N_23165,N_23160);
nor U23351 (N_23351,N_23037,N_23068);
xnor U23352 (N_23352,N_23115,N_23057);
nand U23353 (N_23353,N_23042,N_23072);
xor U23354 (N_23354,N_23165,N_23034);
xnor U23355 (N_23355,N_23015,N_23035);
or U23356 (N_23356,N_23114,N_23121);
xnor U23357 (N_23357,N_23093,N_23159);
nor U23358 (N_23358,N_23131,N_23023);
or U23359 (N_23359,N_23072,N_23055);
nand U23360 (N_23360,N_23012,N_23124);
or U23361 (N_23361,N_23036,N_23009);
nor U23362 (N_23362,N_23164,N_23004);
xor U23363 (N_23363,N_23194,N_23011);
nor U23364 (N_23364,N_23000,N_23076);
or U23365 (N_23365,N_23190,N_23005);
nor U23366 (N_23366,N_23008,N_23051);
nand U23367 (N_23367,N_23172,N_23179);
nand U23368 (N_23368,N_23194,N_23057);
nand U23369 (N_23369,N_23061,N_23142);
and U23370 (N_23370,N_23124,N_23160);
nor U23371 (N_23371,N_23061,N_23176);
nand U23372 (N_23372,N_23077,N_23190);
nand U23373 (N_23373,N_23101,N_23009);
or U23374 (N_23374,N_23102,N_23096);
and U23375 (N_23375,N_23167,N_23153);
and U23376 (N_23376,N_23045,N_23070);
or U23377 (N_23377,N_23188,N_23010);
xor U23378 (N_23378,N_23090,N_23135);
and U23379 (N_23379,N_23175,N_23123);
xor U23380 (N_23380,N_23050,N_23055);
or U23381 (N_23381,N_23188,N_23127);
xor U23382 (N_23382,N_23080,N_23009);
xnor U23383 (N_23383,N_23083,N_23100);
and U23384 (N_23384,N_23111,N_23072);
nand U23385 (N_23385,N_23052,N_23013);
xnor U23386 (N_23386,N_23139,N_23053);
nor U23387 (N_23387,N_23093,N_23158);
nor U23388 (N_23388,N_23143,N_23190);
nor U23389 (N_23389,N_23052,N_23041);
xor U23390 (N_23390,N_23012,N_23071);
nand U23391 (N_23391,N_23046,N_23090);
or U23392 (N_23392,N_23095,N_23021);
or U23393 (N_23393,N_23152,N_23134);
nand U23394 (N_23394,N_23057,N_23146);
or U23395 (N_23395,N_23038,N_23190);
xnor U23396 (N_23396,N_23044,N_23020);
or U23397 (N_23397,N_23169,N_23135);
nand U23398 (N_23398,N_23119,N_23029);
nor U23399 (N_23399,N_23109,N_23150);
or U23400 (N_23400,N_23275,N_23379);
xor U23401 (N_23401,N_23362,N_23337);
and U23402 (N_23402,N_23267,N_23213);
or U23403 (N_23403,N_23228,N_23286);
nand U23404 (N_23404,N_23236,N_23377);
nor U23405 (N_23405,N_23391,N_23249);
nand U23406 (N_23406,N_23347,N_23322);
nand U23407 (N_23407,N_23247,N_23250);
nor U23408 (N_23408,N_23277,N_23332);
and U23409 (N_23409,N_23372,N_23309);
or U23410 (N_23410,N_23371,N_23387);
or U23411 (N_23411,N_23375,N_23283);
xor U23412 (N_23412,N_23308,N_23346);
xor U23413 (N_23413,N_23221,N_23384);
or U23414 (N_23414,N_23209,N_23208);
nand U23415 (N_23415,N_23356,N_23292);
and U23416 (N_23416,N_23380,N_23295);
nand U23417 (N_23417,N_23358,N_23211);
or U23418 (N_23418,N_23315,N_23271);
nor U23419 (N_23419,N_23293,N_23300);
and U23420 (N_23420,N_23280,N_23364);
and U23421 (N_23421,N_23298,N_23397);
nor U23422 (N_23422,N_23279,N_23386);
nand U23423 (N_23423,N_23239,N_23305);
or U23424 (N_23424,N_23307,N_23355);
nor U23425 (N_23425,N_23297,N_23222);
nor U23426 (N_23426,N_23312,N_23264);
xor U23427 (N_23427,N_23203,N_23288);
and U23428 (N_23428,N_23357,N_23234);
nand U23429 (N_23429,N_23302,N_23299);
and U23430 (N_23430,N_23255,N_23329);
or U23431 (N_23431,N_23219,N_23393);
or U23432 (N_23432,N_23254,N_23216);
or U23433 (N_23433,N_23323,N_23304);
nand U23434 (N_23434,N_23328,N_23217);
xor U23435 (N_23435,N_23349,N_23282);
and U23436 (N_23436,N_23206,N_23246);
xnor U23437 (N_23437,N_23338,N_23289);
nand U23438 (N_23438,N_23242,N_23301);
nor U23439 (N_23439,N_23240,N_23398);
nor U23440 (N_23440,N_23251,N_23265);
nand U23441 (N_23441,N_23274,N_23243);
xnor U23442 (N_23442,N_23260,N_23320);
nor U23443 (N_23443,N_23294,N_23248);
xor U23444 (N_23444,N_23369,N_23385);
xor U23445 (N_23445,N_23319,N_23218);
nor U23446 (N_23446,N_23335,N_23258);
or U23447 (N_23447,N_23359,N_23253);
nor U23448 (N_23448,N_23317,N_23245);
nor U23449 (N_23449,N_23310,N_23224);
nand U23450 (N_23450,N_23395,N_23365);
nand U23451 (N_23451,N_23363,N_23210);
nor U23452 (N_23452,N_23231,N_23326);
or U23453 (N_23453,N_23223,N_23204);
xor U23454 (N_23454,N_23202,N_23296);
or U23455 (N_23455,N_23284,N_23316);
or U23456 (N_23456,N_23360,N_23268);
nand U23457 (N_23457,N_23276,N_23287);
nor U23458 (N_23458,N_23321,N_23230);
or U23459 (N_23459,N_23256,N_23374);
or U23460 (N_23460,N_23200,N_23373);
nor U23461 (N_23461,N_23237,N_23348);
and U23462 (N_23462,N_23232,N_23383);
or U23463 (N_23463,N_23306,N_23318);
nor U23464 (N_23464,N_23388,N_23330);
nor U23465 (N_23465,N_23361,N_23311);
nor U23466 (N_23466,N_23342,N_23350);
nor U23467 (N_23467,N_23353,N_23207);
nand U23468 (N_23468,N_23229,N_23259);
nand U23469 (N_23469,N_23257,N_23394);
nor U23470 (N_23470,N_23220,N_23336);
nand U23471 (N_23471,N_23227,N_23341);
or U23472 (N_23472,N_23291,N_23376);
nor U23473 (N_23473,N_23366,N_23252);
xor U23474 (N_23474,N_23325,N_23269);
nor U23475 (N_23475,N_23238,N_23351);
xor U23476 (N_23476,N_23390,N_23345);
or U23477 (N_23477,N_23281,N_23314);
nand U23478 (N_23478,N_23333,N_23244);
nand U23479 (N_23479,N_23226,N_23225);
and U23480 (N_23480,N_23340,N_23233);
nor U23481 (N_23481,N_23313,N_23290);
xnor U23482 (N_23482,N_23339,N_23389);
xnor U23483 (N_23483,N_23327,N_23367);
xnor U23484 (N_23484,N_23278,N_23331);
nor U23485 (N_23485,N_23273,N_23334);
and U23486 (N_23486,N_23263,N_23399);
xor U23487 (N_23487,N_23378,N_23205);
nand U23488 (N_23488,N_23392,N_23381);
xnor U23489 (N_23489,N_23214,N_23368);
and U23490 (N_23490,N_23262,N_23235);
nand U23491 (N_23491,N_23212,N_23343);
nor U23492 (N_23492,N_23396,N_23215);
xnor U23493 (N_23493,N_23285,N_23352);
nor U23494 (N_23494,N_23261,N_23270);
nor U23495 (N_23495,N_23354,N_23344);
nor U23496 (N_23496,N_23272,N_23382);
and U23497 (N_23497,N_23303,N_23241);
nor U23498 (N_23498,N_23370,N_23266);
nand U23499 (N_23499,N_23201,N_23324);
xnor U23500 (N_23500,N_23397,N_23296);
and U23501 (N_23501,N_23381,N_23384);
nor U23502 (N_23502,N_23360,N_23390);
nand U23503 (N_23503,N_23216,N_23339);
xnor U23504 (N_23504,N_23319,N_23337);
nand U23505 (N_23505,N_23212,N_23281);
and U23506 (N_23506,N_23260,N_23285);
nor U23507 (N_23507,N_23349,N_23201);
xor U23508 (N_23508,N_23398,N_23266);
nand U23509 (N_23509,N_23356,N_23312);
or U23510 (N_23510,N_23396,N_23265);
xor U23511 (N_23511,N_23240,N_23341);
and U23512 (N_23512,N_23310,N_23309);
nand U23513 (N_23513,N_23262,N_23240);
nor U23514 (N_23514,N_23382,N_23209);
or U23515 (N_23515,N_23352,N_23368);
xor U23516 (N_23516,N_23223,N_23325);
or U23517 (N_23517,N_23226,N_23268);
xnor U23518 (N_23518,N_23265,N_23222);
xor U23519 (N_23519,N_23227,N_23382);
nor U23520 (N_23520,N_23350,N_23333);
or U23521 (N_23521,N_23313,N_23374);
xnor U23522 (N_23522,N_23250,N_23372);
nand U23523 (N_23523,N_23373,N_23264);
nor U23524 (N_23524,N_23203,N_23239);
xor U23525 (N_23525,N_23314,N_23390);
and U23526 (N_23526,N_23223,N_23219);
xor U23527 (N_23527,N_23247,N_23256);
and U23528 (N_23528,N_23374,N_23294);
xor U23529 (N_23529,N_23342,N_23366);
nor U23530 (N_23530,N_23213,N_23300);
xor U23531 (N_23531,N_23290,N_23220);
and U23532 (N_23532,N_23286,N_23332);
xor U23533 (N_23533,N_23397,N_23214);
nor U23534 (N_23534,N_23355,N_23238);
or U23535 (N_23535,N_23366,N_23351);
nand U23536 (N_23536,N_23216,N_23390);
nand U23537 (N_23537,N_23255,N_23319);
nor U23538 (N_23538,N_23263,N_23335);
and U23539 (N_23539,N_23373,N_23292);
nor U23540 (N_23540,N_23266,N_23209);
nor U23541 (N_23541,N_23279,N_23264);
nor U23542 (N_23542,N_23300,N_23243);
nor U23543 (N_23543,N_23375,N_23369);
and U23544 (N_23544,N_23300,N_23360);
nand U23545 (N_23545,N_23265,N_23282);
nor U23546 (N_23546,N_23293,N_23217);
and U23547 (N_23547,N_23382,N_23384);
nand U23548 (N_23548,N_23250,N_23225);
nand U23549 (N_23549,N_23383,N_23223);
and U23550 (N_23550,N_23387,N_23290);
nand U23551 (N_23551,N_23207,N_23358);
and U23552 (N_23552,N_23262,N_23209);
xor U23553 (N_23553,N_23228,N_23355);
nor U23554 (N_23554,N_23239,N_23301);
nand U23555 (N_23555,N_23249,N_23353);
xor U23556 (N_23556,N_23218,N_23233);
xor U23557 (N_23557,N_23238,N_23251);
nor U23558 (N_23558,N_23233,N_23315);
or U23559 (N_23559,N_23352,N_23394);
or U23560 (N_23560,N_23221,N_23313);
nor U23561 (N_23561,N_23342,N_23206);
xnor U23562 (N_23562,N_23281,N_23399);
xnor U23563 (N_23563,N_23323,N_23297);
or U23564 (N_23564,N_23207,N_23388);
and U23565 (N_23565,N_23281,N_23360);
and U23566 (N_23566,N_23326,N_23271);
xor U23567 (N_23567,N_23272,N_23334);
nor U23568 (N_23568,N_23310,N_23297);
xor U23569 (N_23569,N_23388,N_23225);
nor U23570 (N_23570,N_23235,N_23338);
nand U23571 (N_23571,N_23290,N_23325);
nand U23572 (N_23572,N_23295,N_23203);
xor U23573 (N_23573,N_23239,N_23398);
nor U23574 (N_23574,N_23328,N_23296);
nand U23575 (N_23575,N_23364,N_23345);
and U23576 (N_23576,N_23241,N_23332);
or U23577 (N_23577,N_23361,N_23347);
and U23578 (N_23578,N_23254,N_23307);
xnor U23579 (N_23579,N_23244,N_23309);
nand U23580 (N_23580,N_23286,N_23397);
nand U23581 (N_23581,N_23264,N_23242);
and U23582 (N_23582,N_23233,N_23226);
and U23583 (N_23583,N_23387,N_23361);
xor U23584 (N_23584,N_23301,N_23335);
and U23585 (N_23585,N_23275,N_23223);
and U23586 (N_23586,N_23266,N_23322);
xor U23587 (N_23587,N_23240,N_23377);
nor U23588 (N_23588,N_23225,N_23208);
nand U23589 (N_23589,N_23242,N_23391);
and U23590 (N_23590,N_23398,N_23227);
nand U23591 (N_23591,N_23359,N_23289);
nor U23592 (N_23592,N_23398,N_23276);
xnor U23593 (N_23593,N_23200,N_23226);
and U23594 (N_23594,N_23229,N_23246);
nand U23595 (N_23595,N_23397,N_23249);
and U23596 (N_23596,N_23386,N_23205);
nor U23597 (N_23597,N_23394,N_23258);
xnor U23598 (N_23598,N_23281,N_23356);
nand U23599 (N_23599,N_23235,N_23355);
xnor U23600 (N_23600,N_23414,N_23499);
or U23601 (N_23601,N_23445,N_23541);
and U23602 (N_23602,N_23454,N_23473);
xor U23603 (N_23603,N_23425,N_23578);
nand U23604 (N_23604,N_23467,N_23463);
xor U23605 (N_23605,N_23589,N_23462);
nor U23606 (N_23606,N_23479,N_23456);
and U23607 (N_23607,N_23549,N_23400);
and U23608 (N_23608,N_23553,N_23406);
nand U23609 (N_23609,N_23481,N_23452);
nand U23610 (N_23610,N_23519,N_23436);
nor U23611 (N_23611,N_23582,N_23573);
and U23612 (N_23612,N_23496,N_23548);
nor U23613 (N_23613,N_23470,N_23599);
nor U23614 (N_23614,N_23587,N_23528);
xnor U23615 (N_23615,N_23565,N_23444);
xor U23616 (N_23616,N_23505,N_23430);
or U23617 (N_23617,N_23408,N_23418);
and U23618 (N_23618,N_23506,N_23498);
xnor U23619 (N_23619,N_23596,N_23522);
xor U23620 (N_23620,N_23564,N_23434);
or U23621 (N_23621,N_23533,N_23568);
and U23622 (N_23622,N_23449,N_23560);
or U23623 (N_23623,N_23521,N_23459);
nor U23624 (N_23624,N_23551,N_23598);
or U23625 (N_23625,N_23590,N_23489);
nor U23626 (N_23626,N_23402,N_23588);
xor U23627 (N_23627,N_23442,N_23535);
xnor U23628 (N_23628,N_23439,N_23577);
nand U23629 (N_23629,N_23453,N_23433);
nand U23630 (N_23630,N_23404,N_23500);
or U23631 (N_23631,N_23552,N_23458);
nand U23632 (N_23632,N_23591,N_23483);
nor U23633 (N_23633,N_23477,N_23586);
xnor U23634 (N_23634,N_23469,N_23597);
nand U23635 (N_23635,N_23562,N_23474);
or U23636 (N_23636,N_23503,N_23464);
or U23637 (N_23637,N_23514,N_23416);
nor U23638 (N_23638,N_23450,N_23401);
nor U23639 (N_23639,N_23538,N_23545);
or U23640 (N_23640,N_23516,N_23572);
or U23641 (N_23641,N_23569,N_23525);
and U23642 (N_23642,N_23455,N_23494);
xor U23643 (N_23643,N_23508,N_23429);
xor U23644 (N_23644,N_23451,N_23446);
xor U23645 (N_23645,N_23515,N_23421);
and U23646 (N_23646,N_23540,N_23559);
xor U23647 (N_23647,N_23576,N_23490);
nor U23648 (N_23648,N_23593,N_23524);
and U23649 (N_23649,N_23413,N_23511);
nand U23650 (N_23650,N_23443,N_23571);
nor U23651 (N_23651,N_23512,N_23484);
nor U23652 (N_23652,N_23407,N_23428);
nand U23653 (N_23653,N_23448,N_23475);
and U23654 (N_23654,N_23476,N_23461);
or U23655 (N_23655,N_23495,N_23580);
or U23656 (N_23656,N_23544,N_23504);
xnor U23657 (N_23657,N_23513,N_23594);
xor U23658 (N_23658,N_23426,N_23547);
nand U23659 (N_23659,N_23447,N_23419);
nand U23660 (N_23660,N_23595,N_23563);
and U23661 (N_23661,N_23466,N_23412);
nor U23662 (N_23662,N_23537,N_23501);
nand U23663 (N_23663,N_23510,N_23435);
and U23664 (N_23664,N_23530,N_23584);
and U23665 (N_23665,N_23529,N_23542);
or U23666 (N_23666,N_23415,N_23480);
xor U23667 (N_23667,N_23536,N_23487);
and U23668 (N_23668,N_23583,N_23558);
xor U23669 (N_23669,N_23554,N_23485);
xnor U23670 (N_23670,N_23539,N_23523);
xnor U23671 (N_23671,N_23555,N_23592);
nand U23672 (N_23672,N_23437,N_23420);
and U23673 (N_23673,N_23431,N_23546);
and U23674 (N_23674,N_23465,N_23509);
xnor U23675 (N_23675,N_23492,N_23518);
or U23676 (N_23676,N_23417,N_23478);
nor U23677 (N_23677,N_23566,N_23432);
nor U23678 (N_23678,N_23422,N_23585);
or U23679 (N_23679,N_23410,N_23543);
xor U23680 (N_23680,N_23460,N_23532);
xnor U23681 (N_23681,N_23556,N_23424);
and U23682 (N_23682,N_23440,N_23423);
nor U23683 (N_23683,N_23561,N_23405);
and U23684 (N_23684,N_23493,N_23482);
and U23685 (N_23685,N_23517,N_23441);
xor U23686 (N_23686,N_23457,N_23471);
nand U23687 (N_23687,N_23579,N_23491);
nor U23688 (N_23688,N_23438,N_23574);
or U23689 (N_23689,N_23531,N_23570);
xor U23690 (N_23690,N_23427,N_23411);
xnor U23691 (N_23691,N_23468,N_23520);
xnor U23692 (N_23692,N_23575,N_23557);
nor U23693 (N_23693,N_23581,N_23507);
nor U23694 (N_23694,N_23497,N_23527);
nor U23695 (N_23695,N_23403,N_23534);
xnor U23696 (N_23696,N_23486,N_23409);
nor U23697 (N_23697,N_23526,N_23472);
or U23698 (N_23698,N_23502,N_23488);
nand U23699 (N_23699,N_23567,N_23550);
nand U23700 (N_23700,N_23527,N_23516);
nand U23701 (N_23701,N_23530,N_23482);
or U23702 (N_23702,N_23511,N_23508);
nand U23703 (N_23703,N_23415,N_23580);
nor U23704 (N_23704,N_23445,N_23442);
nor U23705 (N_23705,N_23511,N_23458);
or U23706 (N_23706,N_23589,N_23500);
xnor U23707 (N_23707,N_23515,N_23480);
or U23708 (N_23708,N_23456,N_23459);
xor U23709 (N_23709,N_23409,N_23579);
and U23710 (N_23710,N_23509,N_23442);
xnor U23711 (N_23711,N_23584,N_23422);
or U23712 (N_23712,N_23519,N_23506);
nor U23713 (N_23713,N_23403,N_23467);
xnor U23714 (N_23714,N_23530,N_23562);
nor U23715 (N_23715,N_23540,N_23464);
nand U23716 (N_23716,N_23416,N_23400);
xor U23717 (N_23717,N_23475,N_23459);
and U23718 (N_23718,N_23401,N_23453);
nor U23719 (N_23719,N_23582,N_23492);
or U23720 (N_23720,N_23596,N_23483);
or U23721 (N_23721,N_23468,N_23580);
nand U23722 (N_23722,N_23564,N_23494);
and U23723 (N_23723,N_23465,N_23510);
xor U23724 (N_23724,N_23524,N_23574);
nand U23725 (N_23725,N_23425,N_23506);
and U23726 (N_23726,N_23408,N_23456);
nand U23727 (N_23727,N_23566,N_23425);
nor U23728 (N_23728,N_23542,N_23520);
nor U23729 (N_23729,N_23593,N_23485);
xor U23730 (N_23730,N_23402,N_23515);
and U23731 (N_23731,N_23563,N_23461);
and U23732 (N_23732,N_23434,N_23588);
nand U23733 (N_23733,N_23595,N_23480);
nand U23734 (N_23734,N_23435,N_23517);
xor U23735 (N_23735,N_23435,N_23562);
xnor U23736 (N_23736,N_23467,N_23544);
or U23737 (N_23737,N_23440,N_23552);
xor U23738 (N_23738,N_23503,N_23437);
nor U23739 (N_23739,N_23404,N_23408);
nor U23740 (N_23740,N_23490,N_23429);
nand U23741 (N_23741,N_23471,N_23466);
nand U23742 (N_23742,N_23588,N_23459);
or U23743 (N_23743,N_23589,N_23508);
nor U23744 (N_23744,N_23511,N_23415);
xnor U23745 (N_23745,N_23408,N_23579);
nor U23746 (N_23746,N_23513,N_23455);
xor U23747 (N_23747,N_23582,N_23519);
xor U23748 (N_23748,N_23430,N_23515);
and U23749 (N_23749,N_23532,N_23470);
nand U23750 (N_23750,N_23552,N_23481);
nand U23751 (N_23751,N_23550,N_23598);
and U23752 (N_23752,N_23526,N_23463);
nor U23753 (N_23753,N_23558,N_23534);
or U23754 (N_23754,N_23438,N_23460);
or U23755 (N_23755,N_23502,N_23521);
or U23756 (N_23756,N_23478,N_23465);
nor U23757 (N_23757,N_23439,N_23432);
and U23758 (N_23758,N_23457,N_23415);
and U23759 (N_23759,N_23411,N_23440);
nor U23760 (N_23760,N_23552,N_23503);
and U23761 (N_23761,N_23490,N_23512);
nand U23762 (N_23762,N_23531,N_23566);
nor U23763 (N_23763,N_23426,N_23480);
nand U23764 (N_23764,N_23487,N_23486);
nor U23765 (N_23765,N_23408,N_23599);
nand U23766 (N_23766,N_23597,N_23491);
or U23767 (N_23767,N_23552,N_23542);
nor U23768 (N_23768,N_23533,N_23597);
xnor U23769 (N_23769,N_23558,N_23586);
nor U23770 (N_23770,N_23584,N_23582);
or U23771 (N_23771,N_23590,N_23486);
and U23772 (N_23772,N_23563,N_23531);
or U23773 (N_23773,N_23574,N_23539);
and U23774 (N_23774,N_23489,N_23513);
and U23775 (N_23775,N_23569,N_23452);
or U23776 (N_23776,N_23425,N_23542);
xor U23777 (N_23777,N_23492,N_23443);
xnor U23778 (N_23778,N_23598,N_23559);
or U23779 (N_23779,N_23583,N_23581);
and U23780 (N_23780,N_23556,N_23537);
and U23781 (N_23781,N_23521,N_23544);
nor U23782 (N_23782,N_23560,N_23445);
and U23783 (N_23783,N_23559,N_23494);
nand U23784 (N_23784,N_23476,N_23554);
and U23785 (N_23785,N_23467,N_23560);
nand U23786 (N_23786,N_23555,N_23504);
xnor U23787 (N_23787,N_23433,N_23551);
xor U23788 (N_23788,N_23498,N_23521);
nor U23789 (N_23789,N_23581,N_23500);
nand U23790 (N_23790,N_23497,N_23423);
or U23791 (N_23791,N_23458,N_23551);
or U23792 (N_23792,N_23403,N_23429);
xor U23793 (N_23793,N_23525,N_23458);
nor U23794 (N_23794,N_23436,N_23463);
xor U23795 (N_23795,N_23455,N_23426);
or U23796 (N_23796,N_23582,N_23456);
nand U23797 (N_23797,N_23465,N_23592);
xnor U23798 (N_23798,N_23424,N_23569);
or U23799 (N_23799,N_23554,N_23493);
and U23800 (N_23800,N_23667,N_23698);
xnor U23801 (N_23801,N_23776,N_23658);
nor U23802 (N_23802,N_23735,N_23700);
nand U23803 (N_23803,N_23651,N_23668);
nand U23804 (N_23804,N_23756,N_23665);
or U23805 (N_23805,N_23736,N_23683);
xor U23806 (N_23806,N_23708,N_23768);
or U23807 (N_23807,N_23704,N_23779);
nor U23808 (N_23808,N_23709,N_23721);
and U23809 (N_23809,N_23669,N_23797);
xor U23810 (N_23810,N_23688,N_23636);
and U23811 (N_23811,N_23793,N_23731);
xor U23812 (N_23812,N_23714,N_23650);
nand U23813 (N_23813,N_23607,N_23653);
nor U23814 (N_23814,N_23718,N_23766);
nor U23815 (N_23815,N_23646,N_23618);
xor U23816 (N_23816,N_23690,N_23716);
nor U23817 (N_23817,N_23678,N_23730);
and U23818 (N_23818,N_23712,N_23727);
nor U23819 (N_23819,N_23614,N_23626);
nor U23820 (N_23820,N_23620,N_23649);
or U23821 (N_23821,N_23640,N_23785);
and U23822 (N_23822,N_23654,N_23792);
or U23823 (N_23823,N_23799,N_23775);
xnor U23824 (N_23824,N_23770,N_23629);
or U23825 (N_23825,N_23719,N_23642);
nor U23826 (N_23826,N_23788,N_23624);
or U23827 (N_23827,N_23663,N_23764);
xnor U23828 (N_23828,N_23774,N_23782);
or U23829 (N_23829,N_23689,N_23790);
nand U23830 (N_23830,N_23726,N_23710);
and U23831 (N_23831,N_23701,N_23724);
nor U23832 (N_23832,N_23615,N_23632);
nand U23833 (N_23833,N_23659,N_23706);
nor U23834 (N_23834,N_23783,N_23621);
nand U23835 (N_23835,N_23773,N_23753);
or U23836 (N_23836,N_23630,N_23713);
and U23837 (N_23837,N_23674,N_23694);
nand U23838 (N_23838,N_23671,N_23778);
xnor U23839 (N_23839,N_23657,N_23670);
nor U23840 (N_23840,N_23639,N_23641);
and U23841 (N_23841,N_23613,N_23647);
xor U23842 (N_23842,N_23711,N_23787);
xor U23843 (N_23843,N_23611,N_23784);
and U23844 (N_23844,N_23677,N_23746);
nand U23845 (N_23845,N_23666,N_23699);
xnor U23846 (N_23846,N_23762,N_23656);
and U23847 (N_23847,N_23748,N_23728);
nor U23848 (N_23848,N_23794,N_23696);
or U23849 (N_23849,N_23686,N_23755);
or U23850 (N_23850,N_23743,N_23729);
nand U23851 (N_23851,N_23679,N_23601);
nor U23852 (N_23852,N_23625,N_23759);
nand U23853 (N_23853,N_23617,N_23765);
nor U23854 (N_23854,N_23702,N_23619);
xnor U23855 (N_23855,N_23744,N_23742);
and U23856 (N_23856,N_23623,N_23681);
nand U23857 (N_23857,N_23740,N_23780);
xnor U23858 (N_23858,N_23703,N_23761);
or U23859 (N_23859,N_23795,N_23644);
and U23860 (N_23860,N_23661,N_23687);
nand U23861 (N_23861,N_23691,N_23750);
nand U23862 (N_23862,N_23760,N_23628);
xor U23863 (N_23863,N_23786,N_23789);
nand U23864 (N_23864,N_23685,N_23637);
and U23865 (N_23865,N_23638,N_23692);
or U23866 (N_23866,N_23609,N_23734);
or U23867 (N_23867,N_23739,N_23732);
and U23868 (N_23868,N_23752,N_23664);
xor U23869 (N_23869,N_23643,N_23717);
xor U23870 (N_23870,N_23680,N_23715);
and U23871 (N_23871,N_23682,N_23738);
or U23872 (N_23872,N_23608,N_23747);
nor U23873 (N_23873,N_23791,N_23604);
xnor U23874 (N_23874,N_23769,N_23612);
nor U23875 (N_23875,N_23684,N_23648);
nand U23876 (N_23876,N_23749,N_23605);
and U23877 (N_23877,N_23737,N_23741);
or U23878 (N_23878,N_23722,N_23672);
nor U23879 (N_23879,N_23723,N_23600);
nor U23880 (N_23880,N_23733,N_23602);
and U23881 (N_23881,N_23662,N_23757);
and U23882 (N_23882,N_23627,N_23763);
or U23883 (N_23883,N_23758,N_23777);
or U23884 (N_23884,N_23631,N_23675);
nand U23885 (N_23885,N_23781,N_23645);
or U23886 (N_23886,N_23622,N_23652);
and U23887 (N_23887,N_23616,N_23673);
and U23888 (N_23888,N_23720,N_23798);
or U23889 (N_23889,N_23693,N_23676);
and U23890 (N_23890,N_23603,N_23633);
or U23891 (N_23891,N_23697,N_23655);
xor U23892 (N_23892,N_23634,N_23660);
nand U23893 (N_23893,N_23695,N_23754);
xnor U23894 (N_23894,N_23771,N_23635);
nor U23895 (N_23895,N_23745,N_23796);
and U23896 (N_23896,N_23751,N_23705);
nand U23897 (N_23897,N_23725,N_23610);
xnor U23898 (N_23898,N_23767,N_23772);
nor U23899 (N_23899,N_23606,N_23707);
xnor U23900 (N_23900,N_23663,N_23689);
nand U23901 (N_23901,N_23603,N_23738);
or U23902 (N_23902,N_23765,N_23729);
or U23903 (N_23903,N_23629,N_23685);
or U23904 (N_23904,N_23708,N_23633);
and U23905 (N_23905,N_23740,N_23706);
and U23906 (N_23906,N_23675,N_23785);
nand U23907 (N_23907,N_23626,N_23620);
and U23908 (N_23908,N_23758,N_23708);
nand U23909 (N_23909,N_23642,N_23715);
nand U23910 (N_23910,N_23711,N_23751);
nand U23911 (N_23911,N_23729,N_23667);
xor U23912 (N_23912,N_23711,N_23710);
or U23913 (N_23913,N_23624,N_23745);
nor U23914 (N_23914,N_23788,N_23696);
or U23915 (N_23915,N_23682,N_23770);
xor U23916 (N_23916,N_23624,N_23662);
and U23917 (N_23917,N_23674,N_23713);
and U23918 (N_23918,N_23669,N_23653);
and U23919 (N_23919,N_23664,N_23670);
or U23920 (N_23920,N_23776,N_23616);
nor U23921 (N_23921,N_23778,N_23739);
nor U23922 (N_23922,N_23785,N_23719);
nand U23923 (N_23923,N_23786,N_23793);
nor U23924 (N_23924,N_23674,N_23636);
nand U23925 (N_23925,N_23785,N_23748);
nor U23926 (N_23926,N_23773,N_23673);
nor U23927 (N_23927,N_23674,N_23718);
xnor U23928 (N_23928,N_23646,N_23721);
nand U23929 (N_23929,N_23727,N_23730);
xnor U23930 (N_23930,N_23755,N_23684);
nor U23931 (N_23931,N_23636,N_23728);
and U23932 (N_23932,N_23733,N_23634);
nor U23933 (N_23933,N_23779,N_23677);
xor U23934 (N_23934,N_23790,N_23704);
and U23935 (N_23935,N_23609,N_23601);
or U23936 (N_23936,N_23724,N_23689);
and U23937 (N_23937,N_23686,N_23778);
xnor U23938 (N_23938,N_23697,N_23625);
or U23939 (N_23939,N_23642,N_23690);
nor U23940 (N_23940,N_23614,N_23744);
xnor U23941 (N_23941,N_23667,N_23766);
xor U23942 (N_23942,N_23752,N_23613);
and U23943 (N_23943,N_23731,N_23779);
nand U23944 (N_23944,N_23765,N_23788);
xor U23945 (N_23945,N_23674,N_23622);
nor U23946 (N_23946,N_23729,N_23695);
xor U23947 (N_23947,N_23759,N_23621);
and U23948 (N_23948,N_23683,N_23601);
nor U23949 (N_23949,N_23775,N_23757);
nor U23950 (N_23950,N_23652,N_23657);
nor U23951 (N_23951,N_23744,N_23632);
and U23952 (N_23952,N_23729,N_23788);
nor U23953 (N_23953,N_23672,N_23707);
and U23954 (N_23954,N_23646,N_23785);
or U23955 (N_23955,N_23707,N_23764);
and U23956 (N_23956,N_23732,N_23622);
or U23957 (N_23957,N_23605,N_23764);
or U23958 (N_23958,N_23754,N_23716);
and U23959 (N_23959,N_23604,N_23648);
or U23960 (N_23960,N_23772,N_23729);
or U23961 (N_23961,N_23677,N_23699);
xnor U23962 (N_23962,N_23767,N_23738);
xor U23963 (N_23963,N_23713,N_23758);
nor U23964 (N_23964,N_23776,N_23716);
nand U23965 (N_23965,N_23659,N_23652);
or U23966 (N_23966,N_23762,N_23600);
xnor U23967 (N_23967,N_23674,N_23639);
nand U23968 (N_23968,N_23737,N_23749);
xor U23969 (N_23969,N_23692,N_23653);
and U23970 (N_23970,N_23775,N_23607);
xnor U23971 (N_23971,N_23707,N_23601);
xor U23972 (N_23972,N_23764,N_23622);
or U23973 (N_23973,N_23645,N_23753);
nor U23974 (N_23974,N_23732,N_23636);
or U23975 (N_23975,N_23724,N_23677);
or U23976 (N_23976,N_23682,N_23674);
nor U23977 (N_23977,N_23610,N_23675);
nand U23978 (N_23978,N_23749,N_23702);
nor U23979 (N_23979,N_23778,N_23725);
xnor U23980 (N_23980,N_23771,N_23764);
xnor U23981 (N_23981,N_23796,N_23709);
nand U23982 (N_23982,N_23792,N_23660);
nor U23983 (N_23983,N_23618,N_23731);
nand U23984 (N_23984,N_23774,N_23798);
xnor U23985 (N_23985,N_23776,N_23681);
and U23986 (N_23986,N_23785,N_23635);
and U23987 (N_23987,N_23620,N_23727);
nor U23988 (N_23988,N_23762,N_23758);
xnor U23989 (N_23989,N_23720,N_23672);
or U23990 (N_23990,N_23634,N_23724);
nor U23991 (N_23991,N_23793,N_23706);
or U23992 (N_23992,N_23616,N_23671);
and U23993 (N_23993,N_23660,N_23633);
nand U23994 (N_23994,N_23679,N_23674);
and U23995 (N_23995,N_23690,N_23710);
or U23996 (N_23996,N_23666,N_23702);
nand U23997 (N_23997,N_23739,N_23624);
and U23998 (N_23998,N_23777,N_23652);
xnor U23999 (N_23999,N_23729,N_23633);
xnor U24000 (N_24000,N_23866,N_23846);
nor U24001 (N_24001,N_23997,N_23826);
nand U24002 (N_24002,N_23863,N_23881);
or U24003 (N_24003,N_23808,N_23822);
or U24004 (N_24004,N_23967,N_23904);
or U24005 (N_24005,N_23841,N_23851);
nand U24006 (N_24006,N_23986,N_23943);
nor U24007 (N_24007,N_23999,N_23907);
nand U24008 (N_24008,N_23909,N_23804);
and U24009 (N_24009,N_23853,N_23963);
and U24010 (N_24010,N_23807,N_23940);
nor U24011 (N_24011,N_23875,N_23928);
xor U24012 (N_24012,N_23936,N_23805);
xnor U24013 (N_24013,N_23876,N_23947);
or U24014 (N_24014,N_23827,N_23960);
and U24015 (N_24015,N_23952,N_23954);
nor U24016 (N_24016,N_23932,N_23998);
and U24017 (N_24017,N_23994,N_23860);
nand U24018 (N_24018,N_23983,N_23914);
and U24019 (N_24019,N_23992,N_23981);
nand U24020 (N_24020,N_23942,N_23948);
nand U24021 (N_24021,N_23975,N_23938);
xnor U24022 (N_24022,N_23891,N_23859);
nand U24023 (N_24023,N_23973,N_23923);
nand U24024 (N_24024,N_23824,N_23957);
nor U24025 (N_24025,N_23856,N_23801);
nand U24026 (N_24026,N_23810,N_23872);
nor U24027 (N_24027,N_23982,N_23950);
and U24028 (N_24028,N_23831,N_23832);
or U24029 (N_24029,N_23955,N_23934);
nand U24030 (N_24030,N_23899,N_23953);
xnor U24031 (N_24031,N_23910,N_23916);
nand U24032 (N_24032,N_23877,N_23989);
nor U24033 (N_24033,N_23811,N_23951);
and U24034 (N_24034,N_23913,N_23864);
xnor U24035 (N_24035,N_23901,N_23918);
or U24036 (N_24036,N_23857,N_23930);
and U24037 (N_24037,N_23912,N_23883);
nor U24038 (N_24038,N_23897,N_23880);
xnor U24039 (N_24039,N_23813,N_23849);
xnor U24040 (N_24040,N_23976,N_23980);
and U24041 (N_24041,N_23821,N_23900);
nor U24042 (N_24042,N_23931,N_23803);
and U24043 (N_24043,N_23970,N_23979);
nand U24044 (N_24044,N_23991,N_23958);
nand U24045 (N_24045,N_23886,N_23987);
nand U24046 (N_24046,N_23902,N_23809);
or U24047 (N_24047,N_23917,N_23828);
and U24048 (N_24048,N_23838,N_23988);
or U24049 (N_24049,N_23926,N_23818);
or U24050 (N_24050,N_23946,N_23862);
xnor U24051 (N_24051,N_23819,N_23924);
nand U24052 (N_24052,N_23848,N_23905);
nor U24053 (N_24053,N_23996,N_23993);
nand U24054 (N_24054,N_23888,N_23839);
nand U24055 (N_24055,N_23929,N_23941);
nor U24056 (N_24056,N_23922,N_23817);
xor U24057 (N_24057,N_23816,N_23925);
or U24058 (N_24058,N_23815,N_23858);
nand U24059 (N_24059,N_23835,N_23800);
nor U24060 (N_24060,N_23966,N_23861);
and U24061 (N_24061,N_23995,N_23892);
nor U24062 (N_24062,N_23959,N_23812);
or U24063 (N_24063,N_23871,N_23830);
xnor U24064 (N_24064,N_23919,N_23906);
nor U24065 (N_24065,N_23898,N_23889);
nand U24066 (N_24066,N_23867,N_23874);
or U24067 (N_24067,N_23937,N_23814);
nor U24068 (N_24068,N_23911,N_23956);
nor U24069 (N_24069,N_23964,N_23969);
nand U24070 (N_24070,N_23961,N_23873);
and U24071 (N_24071,N_23921,N_23895);
and U24072 (N_24072,N_23882,N_23990);
xnor U24073 (N_24073,N_23985,N_23842);
nor U24074 (N_24074,N_23978,N_23939);
or U24075 (N_24075,N_23971,N_23845);
or U24076 (N_24076,N_23968,N_23868);
xnor U24077 (N_24077,N_23972,N_23977);
nor U24078 (N_24078,N_23962,N_23920);
nand U24079 (N_24079,N_23885,N_23974);
nor U24080 (N_24080,N_23844,N_23837);
xor U24081 (N_24081,N_23896,N_23878);
nor U24082 (N_24082,N_23820,N_23933);
nand U24083 (N_24083,N_23908,N_23829);
or U24084 (N_24084,N_23865,N_23927);
nand U24085 (N_24085,N_23945,N_23965);
xor U24086 (N_24086,N_23903,N_23949);
or U24087 (N_24087,N_23850,N_23935);
and U24088 (N_24088,N_23870,N_23806);
nor U24089 (N_24089,N_23915,N_23879);
and U24090 (N_24090,N_23825,N_23890);
xnor U24091 (N_24091,N_23847,N_23855);
xor U24092 (N_24092,N_23893,N_23823);
or U24093 (N_24093,N_23984,N_23884);
nor U24094 (N_24094,N_23833,N_23852);
xor U24095 (N_24095,N_23894,N_23869);
nor U24096 (N_24096,N_23802,N_23836);
and U24097 (N_24097,N_23887,N_23854);
or U24098 (N_24098,N_23834,N_23944);
nand U24099 (N_24099,N_23840,N_23843);
nor U24100 (N_24100,N_23886,N_23958);
and U24101 (N_24101,N_23954,N_23806);
nand U24102 (N_24102,N_23974,N_23865);
nor U24103 (N_24103,N_23824,N_23974);
or U24104 (N_24104,N_23865,N_23922);
and U24105 (N_24105,N_23983,N_23803);
nand U24106 (N_24106,N_23998,N_23818);
nand U24107 (N_24107,N_23877,N_23936);
and U24108 (N_24108,N_23891,N_23934);
nand U24109 (N_24109,N_23806,N_23838);
and U24110 (N_24110,N_23960,N_23955);
xor U24111 (N_24111,N_23885,N_23881);
or U24112 (N_24112,N_23870,N_23910);
nor U24113 (N_24113,N_23998,N_23952);
or U24114 (N_24114,N_23848,N_23918);
nand U24115 (N_24115,N_23937,N_23983);
nor U24116 (N_24116,N_23807,N_23980);
and U24117 (N_24117,N_23989,N_23936);
xor U24118 (N_24118,N_23839,N_23867);
xor U24119 (N_24119,N_23901,N_23838);
nor U24120 (N_24120,N_23871,N_23947);
xnor U24121 (N_24121,N_23938,N_23808);
xnor U24122 (N_24122,N_23826,N_23867);
xor U24123 (N_24123,N_23879,N_23977);
or U24124 (N_24124,N_23802,N_23843);
nor U24125 (N_24125,N_23990,N_23950);
nor U24126 (N_24126,N_23923,N_23846);
or U24127 (N_24127,N_23822,N_23828);
nand U24128 (N_24128,N_23984,N_23888);
and U24129 (N_24129,N_23913,N_23821);
and U24130 (N_24130,N_23933,N_23876);
nand U24131 (N_24131,N_23959,N_23827);
nand U24132 (N_24132,N_23877,N_23994);
and U24133 (N_24133,N_23914,N_23882);
or U24134 (N_24134,N_23871,N_23847);
or U24135 (N_24135,N_23985,N_23875);
nand U24136 (N_24136,N_23847,N_23895);
and U24137 (N_24137,N_23963,N_23998);
nand U24138 (N_24138,N_23830,N_23879);
or U24139 (N_24139,N_23800,N_23921);
nor U24140 (N_24140,N_23981,N_23971);
or U24141 (N_24141,N_23919,N_23844);
xor U24142 (N_24142,N_23874,N_23957);
nand U24143 (N_24143,N_23847,N_23978);
nand U24144 (N_24144,N_23876,N_23815);
and U24145 (N_24145,N_23962,N_23849);
nor U24146 (N_24146,N_23965,N_23878);
and U24147 (N_24147,N_23900,N_23893);
nand U24148 (N_24148,N_23816,N_23845);
or U24149 (N_24149,N_23813,N_23811);
and U24150 (N_24150,N_23989,N_23880);
xnor U24151 (N_24151,N_23934,N_23907);
nor U24152 (N_24152,N_23869,N_23898);
nand U24153 (N_24153,N_23921,N_23855);
nor U24154 (N_24154,N_23816,N_23880);
nor U24155 (N_24155,N_23981,N_23838);
and U24156 (N_24156,N_23860,N_23841);
xnor U24157 (N_24157,N_23927,N_23959);
nor U24158 (N_24158,N_23992,N_23861);
nor U24159 (N_24159,N_23835,N_23978);
xnor U24160 (N_24160,N_23869,N_23963);
and U24161 (N_24161,N_23946,N_23854);
and U24162 (N_24162,N_23944,N_23811);
xnor U24163 (N_24163,N_23859,N_23803);
nand U24164 (N_24164,N_23972,N_23945);
nor U24165 (N_24165,N_23955,N_23964);
nand U24166 (N_24166,N_23969,N_23983);
or U24167 (N_24167,N_23909,N_23818);
nor U24168 (N_24168,N_23855,N_23857);
or U24169 (N_24169,N_23976,N_23896);
nand U24170 (N_24170,N_23897,N_23962);
xor U24171 (N_24171,N_23979,N_23848);
and U24172 (N_24172,N_23906,N_23954);
and U24173 (N_24173,N_23951,N_23893);
xnor U24174 (N_24174,N_23931,N_23990);
xnor U24175 (N_24175,N_23915,N_23846);
xnor U24176 (N_24176,N_23917,N_23883);
nand U24177 (N_24177,N_23966,N_23906);
and U24178 (N_24178,N_23926,N_23985);
or U24179 (N_24179,N_23955,N_23966);
nor U24180 (N_24180,N_23909,N_23985);
or U24181 (N_24181,N_23890,N_23930);
nand U24182 (N_24182,N_23970,N_23820);
nand U24183 (N_24183,N_23921,N_23839);
nor U24184 (N_24184,N_23851,N_23845);
xor U24185 (N_24185,N_23865,N_23914);
xnor U24186 (N_24186,N_23826,N_23899);
nor U24187 (N_24187,N_23963,N_23884);
xor U24188 (N_24188,N_23939,N_23869);
or U24189 (N_24189,N_23866,N_23877);
or U24190 (N_24190,N_23957,N_23917);
or U24191 (N_24191,N_23955,N_23907);
xor U24192 (N_24192,N_23872,N_23845);
nand U24193 (N_24193,N_23917,N_23816);
nor U24194 (N_24194,N_23942,N_23984);
or U24195 (N_24195,N_23919,N_23878);
nand U24196 (N_24196,N_23911,N_23802);
or U24197 (N_24197,N_23823,N_23889);
or U24198 (N_24198,N_23875,N_23834);
xor U24199 (N_24199,N_23805,N_23838);
nor U24200 (N_24200,N_24044,N_24091);
or U24201 (N_24201,N_24162,N_24021);
or U24202 (N_24202,N_24001,N_24121);
nor U24203 (N_24203,N_24010,N_24078);
nand U24204 (N_24204,N_24163,N_24125);
nand U24205 (N_24205,N_24159,N_24011);
nand U24206 (N_24206,N_24122,N_24130);
nor U24207 (N_24207,N_24131,N_24156);
nor U24208 (N_24208,N_24185,N_24168);
and U24209 (N_24209,N_24190,N_24027);
and U24210 (N_24210,N_24057,N_24051);
or U24211 (N_24211,N_24107,N_24020);
nor U24212 (N_24212,N_24026,N_24158);
and U24213 (N_24213,N_24147,N_24157);
nor U24214 (N_24214,N_24087,N_24050);
nor U24215 (N_24215,N_24148,N_24053);
and U24216 (N_24216,N_24043,N_24003);
nor U24217 (N_24217,N_24128,N_24046);
or U24218 (N_24218,N_24136,N_24167);
nor U24219 (N_24219,N_24080,N_24041);
nor U24220 (N_24220,N_24047,N_24154);
nor U24221 (N_24221,N_24077,N_24113);
nor U24222 (N_24222,N_24144,N_24195);
xor U24223 (N_24223,N_24065,N_24112);
xnor U24224 (N_24224,N_24141,N_24110);
nor U24225 (N_24225,N_24104,N_24145);
nor U24226 (N_24226,N_24060,N_24038);
xnor U24227 (N_24227,N_24092,N_24064);
xor U24228 (N_24228,N_24007,N_24040);
and U24229 (N_24229,N_24172,N_24174);
and U24230 (N_24230,N_24149,N_24178);
nor U24231 (N_24231,N_24177,N_24096);
nor U24232 (N_24232,N_24164,N_24199);
or U24233 (N_24233,N_24189,N_24133);
xor U24234 (N_24234,N_24151,N_24032);
nand U24235 (N_24235,N_24018,N_24105);
nor U24236 (N_24236,N_24061,N_24187);
or U24237 (N_24237,N_24085,N_24033);
and U24238 (N_24238,N_24120,N_24153);
nor U24239 (N_24239,N_24002,N_24176);
nor U24240 (N_24240,N_24019,N_24037);
xor U24241 (N_24241,N_24028,N_24114);
and U24242 (N_24242,N_24170,N_24138);
or U24243 (N_24243,N_24143,N_24086);
or U24244 (N_24244,N_24070,N_24052);
or U24245 (N_24245,N_24031,N_24197);
xnor U24246 (N_24246,N_24059,N_24048);
nand U24247 (N_24247,N_24132,N_24062);
xnor U24248 (N_24248,N_24067,N_24179);
nand U24249 (N_24249,N_24108,N_24045);
xnor U24250 (N_24250,N_24022,N_24089);
and U24251 (N_24251,N_24036,N_24088);
xnor U24252 (N_24252,N_24135,N_24181);
xnor U24253 (N_24253,N_24063,N_24171);
xor U24254 (N_24254,N_24103,N_24023);
or U24255 (N_24255,N_24074,N_24123);
or U24256 (N_24256,N_24169,N_24069);
nor U24257 (N_24257,N_24008,N_24166);
or U24258 (N_24258,N_24198,N_24073);
xnor U24259 (N_24259,N_24175,N_24068);
and U24260 (N_24260,N_24116,N_24160);
nand U24261 (N_24261,N_24034,N_24014);
xnor U24262 (N_24262,N_24017,N_24058);
nor U24263 (N_24263,N_24106,N_24161);
and U24264 (N_24264,N_24094,N_24035);
or U24265 (N_24265,N_24193,N_24098);
and U24266 (N_24266,N_24173,N_24134);
or U24267 (N_24267,N_24140,N_24191);
and U24268 (N_24268,N_24102,N_24029);
nand U24269 (N_24269,N_24005,N_24071);
and U24270 (N_24270,N_24055,N_24186);
nor U24271 (N_24271,N_24081,N_24054);
nor U24272 (N_24272,N_24015,N_24115);
or U24273 (N_24273,N_24076,N_24016);
and U24274 (N_24274,N_24139,N_24109);
or U24275 (N_24275,N_24101,N_24129);
nand U24276 (N_24276,N_24004,N_24039);
xnor U24277 (N_24277,N_24099,N_24194);
or U24278 (N_24278,N_24009,N_24188);
or U24279 (N_24279,N_24180,N_24095);
and U24280 (N_24280,N_24072,N_24097);
nor U24281 (N_24281,N_24183,N_24118);
or U24282 (N_24282,N_24184,N_24127);
or U24283 (N_24283,N_24155,N_24049);
nor U24284 (N_24284,N_24042,N_24082);
xor U24285 (N_24285,N_24111,N_24152);
nor U24286 (N_24286,N_24090,N_24146);
and U24287 (N_24287,N_24030,N_24013);
xor U24288 (N_24288,N_24025,N_24066);
nand U24289 (N_24289,N_24093,N_24075);
xnor U24290 (N_24290,N_24196,N_24083);
nor U24291 (N_24291,N_24117,N_24142);
and U24292 (N_24292,N_24056,N_24182);
nor U24293 (N_24293,N_24006,N_24165);
and U24294 (N_24294,N_24012,N_24137);
nand U24295 (N_24295,N_24150,N_24079);
and U24296 (N_24296,N_24084,N_24192);
and U24297 (N_24297,N_24100,N_24024);
or U24298 (N_24298,N_24119,N_24124);
nor U24299 (N_24299,N_24000,N_24126);
or U24300 (N_24300,N_24189,N_24101);
nand U24301 (N_24301,N_24157,N_24129);
nor U24302 (N_24302,N_24166,N_24169);
or U24303 (N_24303,N_24040,N_24081);
nand U24304 (N_24304,N_24107,N_24090);
and U24305 (N_24305,N_24155,N_24127);
nor U24306 (N_24306,N_24103,N_24071);
nor U24307 (N_24307,N_24083,N_24011);
and U24308 (N_24308,N_24035,N_24188);
and U24309 (N_24309,N_24032,N_24116);
nand U24310 (N_24310,N_24189,N_24188);
xor U24311 (N_24311,N_24072,N_24022);
nand U24312 (N_24312,N_24142,N_24004);
or U24313 (N_24313,N_24044,N_24171);
nand U24314 (N_24314,N_24157,N_24143);
and U24315 (N_24315,N_24036,N_24121);
nand U24316 (N_24316,N_24159,N_24113);
nor U24317 (N_24317,N_24149,N_24110);
or U24318 (N_24318,N_24026,N_24010);
xor U24319 (N_24319,N_24084,N_24194);
xnor U24320 (N_24320,N_24096,N_24112);
nor U24321 (N_24321,N_24160,N_24036);
nor U24322 (N_24322,N_24012,N_24080);
and U24323 (N_24323,N_24025,N_24106);
nor U24324 (N_24324,N_24084,N_24054);
or U24325 (N_24325,N_24046,N_24037);
or U24326 (N_24326,N_24021,N_24042);
and U24327 (N_24327,N_24010,N_24064);
and U24328 (N_24328,N_24157,N_24124);
xor U24329 (N_24329,N_24022,N_24189);
or U24330 (N_24330,N_24150,N_24055);
and U24331 (N_24331,N_24135,N_24108);
or U24332 (N_24332,N_24103,N_24080);
xnor U24333 (N_24333,N_24179,N_24098);
xor U24334 (N_24334,N_24174,N_24065);
and U24335 (N_24335,N_24155,N_24139);
nand U24336 (N_24336,N_24151,N_24025);
xor U24337 (N_24337,N_24094,N_24050);
or U24338 (N_24338,N_24015,N_24161);
or U24339 (N_24339,N_24054,N_24075);
nor U24340 (N_24340,N_24178,N_24134);
and U24341 (N_24341,N_24164,N_24044);
xor U24342 (N_24342,N_24196,N_24135);
nor U24343 (N_24343,N_24027,N_24099);
nand U24344 (N_24344,N_24086,N_24121);
and U24345 (N_24345,N_24102,N_24002);
nand U24346 (N_24346,N_24056,N_24070);
nor U24347 (N_24347,N_24040,N_24198);
or U24348 (N_24348,N_24093,N_24082);
or U24349 (N_24349,N_24034,N_24106);
and U24350 (N_24350,N_24099,N_24009);
nand U24351 (N_24351,N_24015,N_24032);
nor U24352 (N_24352,N_24153,N_24085);
or U24353 (N_24353,N_24133,N_24111);
or U24354 (N_24354,N_24033,N_24112);
and U24355 (N_24355,N_24061,N_24096);
or U24356 (N_24356,N_24022,N_24170);
or U24357 (N_24357,N_24025,N_24076);
xnor U24358 (N_24358,N_24172,N_24063);
xnor U24359 (N_24359,N_24029,N_24157);
nand U24360 (N_24360,N_24140,N_24162);
nand U24361 (N_24361,N_24017,N_24036);
nand U24362 (N_24362,N_24131,N_24115);
or U24363 (N_24363,N_24087,N_24187);
or U24364 (N_24364,N_24044,N_24086);
or U24365 (N_24365,N_24117,N_24169);
and U24366 (N_24366,N_24113,N_24152);
xor U24367 (N_24367,N_24179,N_24117);
xor U24368 (N_24368,N_24053,N_24133);
and U24369 (N_24369,N_24116,N_24018);
or U24370 (N_24370,N_24183,N_24059);
nor U24371 (N_24371,N_24121,N_24189);
and U24372 (N_24372,N_24075,N_24087);
nor U24373 (N_24373,N_24069,N_24011);
xor U24374 (N_24374,N_24119,N_24015);
xor U24375 (N_24375,N_24138,N_24161);
and U24376 (N_24376,N_24195,N_24069);
and U24377 (N_24377,N_24173,N_24164);
nor U24378 (N_24378,N_24104,N_24011);
and U24379 (N_24379,N_24031,N_24138);
or U24380 (N_24380,N_24025,N_24075);
nor U24381 (N_24381,N_24125,N_24130);
nor U24382 (N_24382,N_24045,N_24189);
and U24383 (N_24383,N_24188,N_24058);
nor U24384 (N_24384,N_24101,N_24022);
nand U24385 (N_24385,N_24144,N_24059);
nor U24386 (N_24386,N_24084,N_24078);
nand U24387 (N_24387,N_24128,N_24189);
nand U24388 (N_24388,N_24075,N_24116);
xor U24389 (N_24389,N_24105,N_24188);
or U24390 (N_24390,N_24009,N_24054);
xnor U24391 (N_24391,N_24183,N_24131);
nand U24392 (N_24392,N_24144,N_24036);
or U24393 (N_24393,N_24137,N_24009);
and U24394 (N_24394,N_24004,N_24091);
or U24395 (N_24395,N_24104,N_24048);
nand U24396 (N_24396,N_24033,N_24132);
nand U24397 (N_24397,N_24056,N_24107);
nand U24398 (N_24398,N_24109,N_24098);
or U24399 (N_24399,N_24037,N_24172);
and U24400 (N_24400,N_24200,N_24363);
nor U24401 (N_24401,N_24215,N_24335);
xnor U24402 (N_24402,N_24264,N_24216);
nor U24403 (N_24403,N_24313,N_24337);
xor U24404 (N_24404,N_24360,N_24301);
and U24405 (N_24405,N_24329,N_24265);
xor U24406 (N_24406,N_24233,N_24386);
nor U24407 (N_24407,N_24280,N_24320);
nor U24408 (N_24408,N_24315,N_24366);
xnor U24409 (N_24409,N_24398,N_24255);
and U24410 (N_24410,N_24269,N_24312);
or U24411 (N_24411,N_24254,N_24227);
nand U24412 (N_24412,N_24244,N_24202);
nand U24413 (N_24413,N_24231,N_24205);
xor U24414 (N_24414,N_24362,N_24214);
nor U24415 (N_24415,N_24295,N_24395);
nor U24416 (N_24416,N_24234,N_24397);
and U24417 (N_24417,N_24352,N_24220);
xor U24418 (N_24418,N_24278,N_24350);
nor U24419 (N_24419,N_24399,N_24296);
and U24420 (N_24420,N_24341,N_24349);
and U24421 (N_24421,N_24380,N_24207);
and U24422 (N_24422,N_24257,N_24361);
or U24423 (N_24423,N_24245,N_24241);
nand U24424 (N_24424,N_24346,N_24336);
xor U24425 (N_24425,N_24388,N_24378);
nand U24426 (N_24426,N_24373,N_24317);
nor U24427 (N_24427,N_24275,N_24294);
xnor U24428 (N_24428,N_24298,N_24267);
nor U24429 (N_24429,N_24332,N_24288);
xnor U24430 (N_24430,N_24209,N_24271);
and U24431 (N_24431,N_24356,N_24225);
nor U24432 (N_24432,N_24310,N_24307);
nor U24433 (N_24433,N_24348,N_24321);
or U24434 (N_24434,N_24258,N_24289);
nand U24435 (N_24435,N_24291,N_24239);
nor U24436 (N_24436,N_24219,N_24224);
nand U24437 (N_24437,N_24268,N_24344);
and U24438 (N_24438,N_24287,N_24338);
and U24439 (N_24439,N_24389,N_24273);
xnor U24440 (N_24440,N_24203,N_24272);
or U24441 (N_24441,N_24355,N_24251);
and U24442 (N_24442,N_24342,N_24229);
or U24443 (N_24443,N_24262,N_24347);
and U24444 (N_24444,N_24247,N_24282);
and U24445 (N_24445,N_24327,N_24256);
nor U24446 (N_24446,N_24381,N_24367);
or U24447 (N_24447,N_24260,N_24324);
nor U24448 (N_24448,N_24331,N_24303);
and U24449 (N_24449,N_24333,N_24261);
xor U24450 (N_24450,N_24283,N_24369);
xor U24451 (N_24451,N_24240,N_24325);
or U24452 (N_24452,N_24354,N_24339);
nor U24453 (N_24453,N_24394,N_24249);
xnor U24454 (N_24454,N_24248,N_24235);
nand U24455 (N_24455,N_24392,N_24328);
or U24456 (N_24456,N_24322,N_24230);
or U24457 (N_24457,N_24326,N_24223);
nor U24458 (N_24458,N_24228,N_24204);
nand U24459 (N_24459,N_24218,N_24384);
xor U24460 (N_24460,N_24374,N_24221);
and U24461 (N_24461,N_24340,N_24285);
or U24462 (N_24462,N_24293,N_24246);
nor U24463 (N_24463,N_24372,N_24238);
or U24464 (N_24464,N_24243,N_24316);
or U24465 (N_24465,N_24211,N_24253);
or U24466 (N_24466,N_24353,N_24343);
xnor U24467 (N_24467,N_24277,N_24306);
nor U24468 (N_24468,N_24274,N_24299);
nor U24469 (N_24469,N_24370,N_24217);
nand U24470 (N_24470,N_24297,N_24377);
xor U24471 (N_24471,N_24387,N_24376);
or U24472 (N_24472,N_24292,N_24393);
nand U24473 (N_24473,N_24305,N_24252);
nor U24474 (N_24474,N_24323,N_24222);
nor U24475 (N_24475,N_24279,N_24212);
nor U24476 (N_24476,N_24213,N_24371);
xor U24477 (N_24477,N_24345,N_24270);
or U24478 (N_24478,N_24330,N_24368);
xnor U24479 (N_24479,N_24276,N_24304);
and U24480 (N_24480,N_24359,N_24311);
or U24481 (N_24481,N_24358,N_24302);
or U24482 (N_24482,N_24396,N_24206);
or U24483 (N_24483,N_24284,N_24390);
and U24484 (N_24484,N_24201,N_24263);
nand U24485 (N_24485,N_24308,N_24351);
nor U24486 (N_24486,N_24250,N_24266);
or U24487 (N_24487,N_24382,N_24383);
nor U24488 (N_24488,N_24309,N_24242);
or U24489 (N_24489,N_24237,N_24286);
or U24490 (N_24490,N_24226,N_24300);
xnor U24491 (N_24491,N_24365,N_24379);
nor U24492 (N_24492,N_24364,N_24357);
nand U24493 (N_24493,N_24236,N_24334);
and U24494 (N_24494,N_24210,N_24314);
xnor U24495 (N_24495,N_24290,N_24232);
nor U24496 (N_24496,N_24385,N_24208);
or U24497 (N_24497,N_24319,N_24259);
and U24498 (N_24498,N_24281,N_24391);
xor U24499 (N_24499,N_24375,N_24318);
or U24500 (N_24500,N_24236,N_24385);
xor U24501 (N_24501,N_24325,N_24265);
xor U24502 (N_24502,N_24394,N_24280);
or U24503 (N_24503,N_24257,N_24343);
or U24504 (N_24504,N_24302,N_24210);
nand U24505 (N_24505,N_24294,N_24387);
nor U24506 (N_24506,N_24382,N_24337);
or U24507 (N_24507,N_24373,N_24352);
and U24508 (N_24508,N_24246,N_24360);
nor U24509 (N_24509,N_24257,N_24261);
xnor U24510 (N_24510,N_24234,N_24368);
nand U24511 (N_24511,N_24265,N_24281);
nand U24512 (N_24512,N_24329,N_24267);
nor U24513 (N_24513,N_24248,N_24285);
nor U24514 (N_24514,N_24371,N_24241);
and U24515 (N_24515,N_24280,N_24324);
and U24516 (N_24516,N_24274,N_24389);
and U24517 (N_24517,N_24204,N_24243);
nand U24518 (N_24518,N_24231,N_24320);
nand U24519 (N_24519,N_24325,N_24201);
nand U24520 (N_24520,N_24249,N_24277);
nor U24521 (N_24521,N_24343,N_24360);
and U24522 (N_24522,N_24338,N_24243);
or U24523 (N_24523,N_24392,N_24310);
or U24524 (N_24524,N_24327,N_24399);
xnor U24525 (N_24525,N_24283,N_24321);
xnor U24526 (N_24526,N_24389,N_24372);
nand U24527 (N_24527,N_24372,N_24356);
and U24528 (N_24528,N_24392,N_24385);
nand U24529 (N_24529,N_24319,N_24368);
xor U24530 (N_24530,N_24383,N_24255);
and U24531 (N_24531,N_24254,N_24249);
nor U24532 (N_24532,N_24366,N_24293);
and U24533 (N_24533,N_24353,N_24231);
nand U24534 (N_24534,N_24263,N_24235);
nor U24535 (N_24535,N_24205,N_24336);
and U24536 (N_24536,N_24380,N_24390);
nor U24537 (N_24537,N_24353,N_24311);
nor U24538 (N_24538,N_24272,N_24264);
nor U24539 (N_24539,N_24340,N_24379);
or U24540 (N_24540,N_24343,N_24347);
and U24541 (N_24541,N_24284,N_24341);
xnor U24542 (N_24542,N_24383,N_24316);
nor U24543 (N_24543,N_24398,N_24261);
nor U24544 (N_24544,N_24224,N_24220);
xor U24545 (N_24545,N_24240,N_24250);
xnor U24546 (N_24546,N_24393,N_24256);
nand U24547 (N_24547,N_24319,N_24297);
nor U24548 (N_24548,N_24376,N_24230);
or U24549 (N_24549,N_24359,N_24305);
nor U24550 (N_24550,N_24223,N_24237);
xor U24551 (N_24551,N_24384,N_24284);
or U24552 (N_24552,N_24283,N_24398);
nor U24553 (N_24553,N_24391,N_24360);
nor U24554 (N_24554,N_24368,N_24265);
xor U24555 (N_24555,N_24386,N_24324);
nand U24556 (N_24556,N_24385,N_24302);
xnor U24557 (N_24557,N_24327,N_24325);
nor U24558 (N_24558,N_24317,N_24399);
nor U24559 (N_24559,N_24334,N_24328);
nor U24560 (N_24560,N_24327,N_24368);
or U24561 (N_24561,N_24397,N_24385);
or U24562 (N_24562,N_24366,N_24272);
xnor U24563 (N_24563,N_24329,N_24363);
xnor U24564 (N_24564,N_24254,N_24302);
xor U24565 (N_24565,N_24353,N_24373);
xnor U24566 (N_24566,N_24329,N_24266);
and U24567 (N_24567,N_24360,N_24202);
or U24568 (N_24568,N_24268,N_24301);
and U24569 (N_24569,N_24303,N_24315);
or U24570 (N_24570,N_24303,N_24381);
and U24571 (N_24571,N_24337,N_24201);
or U24572 (N_24572,N_24314,N_24290);
xor U24573 (N_24573,N_24231,N_24372);
or U24574 (N_24574,N_24379,N_24241);
and U24575 (N_24575,N_24374,N_24232);
nor U24576 (N_24576,N_24302,N_24332);
or U24577 (N_24577,N_24384,N_24221);
or U24578 (N_24578,N_24307,N_24326);
and U24579 (N_24579,N_24355,N_24209);
xnor U24580 (N_24580,N_24265,N_24328);
xnor U24581 (N_24581,N_24241,N_24275);
nand U24582 (N_24582,N_24329,N_24320);
or U24583 (N_24583,N_24260,N_24345);
xnor U24584 (N_24584,N_24334,N_24231);
xor U24585 (N_24585,N_24345,N_24223);
nor U24586 (N_24586,N_24273,N_24210);
nand U24587 (N_24587,N_24332,N_24343);
and U24588 (N_24588,N_24346,N_24218);
and U24589 (N_24589,N_24281,N_24214);
nor U24590 (N_24590,N_24349,N_24253);
nand U24591 (N_24591,N_24307,N_24378);
and U24592 (N_24592,N_24394,N_24202);
nand U24593 (N_24593,N_24389,N_24236);
xor U24594 (N_24594,N_24301,N_24318);
and U24595 (N_24595,N_24312,N_24287);
nand U24596 (N_24596,N_24315,N_24382);
or U24597 (N_24597,N_24231,N_24201);
xnor U24598 (N_24598,N_24256,N_24296);
and U24599 (N_24599,N_24220,N_24328);
nand U24600 (N_24600,N_24404,N_24415);
and U24601 (N_24601,N_24568,N_24527);
and U24602 (N_24602,N_24478,N_24438);
nand U24603 (N_24603,N_24544,N_24531);
nand U24604 (N_24604,N_24461,N_24471);
and U24605 (N_24605,N_24587,N_24402);
xnor U24606 (N_24606,N_24479,N_24542);
nor U24607 (N_24607,N_24485,N_24588);
and U24608 (N_24608,N_24424,N_24571);
nor U24609 (N_24609,N_24406,N_24495);
nand U24610 (N_24610,N_24463,N_24519);
xor U24611 (N_24611,N_24508,N_24462);
nand U24612 (N_24612,N_24559,N_24411);
xor U24613 (N_24613,N_24557,N_24432);
nor U24614 (N_24614,N_24558,N_24524);
nor U24615 (N_24615,N_24577,N_24448);
nand U24616 (N_24616,N_24476,N_24533);
or U24617 (N_24617,N_24430,N_24482);
nor U24618 (N_24618,N_24492,N_24589);
and U24619 (N_24619,N_24539,N_24453);
nor U24620 (N_24620,N_24468,N_24578);
xnor U24621 (N_24621,N_24521,N_24493);
xnor U24622 (N_24622,N_24477,N_24412);
or U24623 (N_24623,N_24565,N_24592);
nor U24624 (N_24624,N_24400,N_24525);
nor U24625 (N_24625,N_24553,N_24509);
nand U24626 (N_24626,N_24538,N_24503);
nand U24627 (N_24627,N_24446,N_24442);
nand U24628 (N_24628,N_24464,N_24431);
or U24629 (N_24629,N_24407,N_24408);
nand U24630 (N_24630,N_24403,N_24585);
or U24631 (N_24631,N_24497,N_24469);
xnor U24632 (N_24632,N_24466,N_24561);
xnor U24633 (N_24633,N_24459,N_24425);
xnor U24634 (N_24634,N_24575,N_24414);
and U24635 (N_24635,N_24455,N_24499);
nand U24636 (N_24636,N_24441,N_24489);
nor U24637 (N_24637,N_24502,N_24529);
xnor U24638 (N_24638,N_24473,N_24570);
nor U24639 (N_24639,N_24449,N_24599);
or U24640 (N_24640,N_24530,N_24593);
nor U24641 (N_24641,N_24549,N_24419);
xor U24642 (N_24642,N_24443,N_24423);
nand U24643 (N_24643,N_24436,N_24512);
and U24644 (N_24644,N_24594,N_24505);
nand U24645 (N_24645,N_24569,N_24450);
and U24646 (N_24646,N_24528,N_24566);
xor U24647 (N_24647,N_24456,N_24439);
xnor U24648 (N_24648,N_24546,N_24437);
nand U24649 (N_24649,N_24444,N_24551);
or U24650 (N_24650,N_24518,N_24548);
nor U24651 (N_24651,N_24435,N_24574);
and U24652 (N_24652,N_24516,N_24547);
xor U24653 (N_24653,N_24540,N_24418);
nor U24654 (N_24654,N_24554,N_24583);
nand U24655 (N_24655,N_24410,N_24433);
and U24656 (N_24656,N_24470,N_24401);
and U24657 (N_24657,N_24532,N_24452);
and U24658 (N_24658,N_24474,N_24564);
nor U24659 (N_24659,N_24465,N_24573);
xor U24660 (N_24660,N_24545,N_24413);
and U24661 (N_24661,N_24504,N_24445);
nand U24662 (N_24662,N_24597,N_24543);
nand U24663 (N_24663,N_24576,N_24496);
or U24664 (N_24664,N_24490,N_24460);
nand U24665 (N_24665,N_24417,N_24506);
nand U24666 (N_24666,N_24500,N_24429);
or U24667 (N_24667,N_24598,N_24494);
nor U24668 (N_24668,N_24567,N_24534);
xor U24669 (N_24669,N_24522,N_24486);
and U24670 (N_24670,N_24458,N_24491);
or U24671 (N_24671,N_24467,N_24472);
xor U24672 (N_24672,N_24526,N_24550);
and U24673 (N_24673,N_24584,N_24541);
nand U24674 (N_24674,N_24421,N_24562);
nand U24675 (N_24675,N_24513,N_24498);
nand U24676 (N_24676,N_24484,N_24427);
or U24677 (N_24677,N_24454,N_24409);
xor U24678 (N_24678,N_24451,N_24536);
xnor U24679 (N_24679,N_24537,N_24579);
xor U24680 (N_24680,N_24426,N_24483);
and U24681 (N_24681,N_24422,N_24535);
nor U24682 (N_24682,N_24501,N_24581);
nand U24683 (N_24683,N_24440,N_24507);
and U24684 (N_24684,N_24586,N_24428);
or U24685 (N_24685,N_24510,N_24580);
nor U24686 (N_24686,N_24556,N_24560);
or U24687 (N_24687,N_24457,N_24552);
nand U24688 (N_24688,N_24405,N_24480);
xor U24689 (N_24689,N_24572,N_24514);
xor U24690 (N_24690,N_24416,N_24596);
nand U24691 (N_24691,N_24488,N_24555);
and U24692 (N_24692,N_24434,N_24563);
xor U24693 (N_24693,N_24582,N_24511);
nor U24694 (N_24694,N_24590,N_24481);
nor U24695 (N_24695,N_24420,N_24447);
and U24696 (N_24696,N_24515,N_24523);
and U24697 (N_24697,N_24517,N_24591);
or U24698 (N_24698,N_24595,N_24487);
xnor U24699 (N_24699,N_24520,N_24475);
or U24700 (N_24700,N_24598,N_24536);
or U24701 (N_24701,N_24586,N_24591);
or U24702 (N_24702,N_24499,N_24584);
and U24703 (N_24703,N_24581,N_24569);
nor U24704 (N_24704,N_24586,N_24541);
or U24705 (N_24705,N_24557,N_24430);
nand U24706 (N_24706,N_24429,N_24510);
and U24707 (N_24707,N_24426,N_24408);
or U24708 (N_24708,N_24482,N_24438);
and U24709 (N_24709,N_24551,N_24452);
xor U24710 (N_24710,N_24444,N_24541);
xor U24711 (N_24711,N_24494,N_24528);
or U24712 (N_24712,N_24531,N_24529);
and U24713 (N_24713,N_24538,N_24470);
and U24714 (N_24714,N_24538,N_24429);
nor U24715 (N_24715,N_24485,N_24494);
or U24716 (N_24716,N_24478,N_24549);
nor U24717 (N_24717,N_24573,N_24530);
or U24718 (N_24718,N_24461,N_24500);
xnor U24719 (N_24719,N_24564,N_24574);
and U24720 (N_24720,N_24495,N_24518);
nor U24721 (N_24721,N_24585,N_24581);
or U24722 (N_24722,N_24503,N_24565);
nand U24723 (N_24723,N_24516,N_24591);
xor U24724 (N_24724,N_24432,N_24502);
and U24725 (N_24725,N_24442,N_24505);
nand U24726 (N_24726,N_24526,N_24448);
or U24727 (N_24727,N_24436,N_24465);
nand U24728 (N_24728,N_24448,N_24482);
and U24729 (N_24729,N_24569,N_24415);
nor U24730 (N_24730,N_24554,N_24496);
nand U24731 (N_24731,N_24434,N_24549);
or U24732 (N_24732,N_24494,N_24549);
and U24733 (N_24733,N_24462,N_24540);
and U24734 (N_24734,N_24499,N_24509);
nand U24735 (N_24735,N_24547,N_24536);
xor U24736 (N_24736,N_24572,N_24407);
or U24737 (N_24737,N_24553,N_24423);
xor U24738 (N_24738,N_24418,N_24583);
and U24739 (N_24739,N_24406,N_24491);
xnor U24740 (N_24740,N_24509,N_24599);
nand U24741 (N_24741,N_24472,N_24515);
xnor U24742 (N_24742,N_24489,N_24412);
and U24743 (N_24743,N_24456,N_24563);
or U24744 (N_24744,N_24560,N_24414);
or U24745 (N_24745,N_24583,N_24436);
nor U24746 (N_24746,N_24555,N_24486);
nor U24747 (N_24747,N_24435,N_24580);
or U24748 (N_24748,N_24553,N_24588);
nor U24749 (N_24749,N_24578,N_24430);
nand U24750 (N_24750,N_24427,N_24570);
nor U24751 (N_24751,N_24439,N_24433);
and U24752 (N_24752,N_24501,N_24579);
xnor U24753 (N_24753,N_24476,N_24446);
nor U24754 (N_24754,N_24570,N_24404);
xnor U24755 (N_24755,N_24583,N_24458);
or U24756 (N_24756,N_24530,N_24442);
nor U24757 (N_24757,N_24507,N_24569);
and U24758 (N_24758,N_24572,N_24523);
nor U24759 (N_24759,N_24417,N_24577);
or U24760 (N_24760,N_24514,N_24563);
nor U24761 (N_24761,N_24578,N_24476);
nor U24762 (N_24762,N_24488,N_24491);
and U24763 (N_24763,N_24592,N_24456);
nand U24764 (N_24764,N_24419,N_24431);
and U24765 (N_24765,N_24473,N_24431);
or U24766 (N_24766,N_24420,N_24405);
or U24767 (N_24767,N_24583,N_24435);
nor U24768 (N_24768,N_24436,N_24459);
nor U24769 (N_24769,N_24554,N_24573);
nand U24770 (N_24770,N_24567,N_24588);
or U24771 (N_24771,N_24563,N_24490);
or U24772 (N_24772,N_24517,N_24484);
and U24773 (N_24773,N_24533,N_24431);
or U24774 (N_24774,N_24503,N_24428);
or U24775 (N_24775,N_24452,N_24415);
and U24776 (N_24776,N_24506,N_24422);
nand U24777 (N_24777,N_24402,N_24540);
nor U24778 (N_24778,N_24514,N_24498);
or U24779 (N_24779,N_24546,N_24516);
or U24780 (N_24780,N_24591,N_24490);
or U24781 (N_24781,N_24454,N_24481);
xnor U24782 (N_24782,N_24546,N_24429);
or U24783 (N_24783,N_24480,N_24503);
nor U24784 (N_24784,N_24427,N_24572);
xor U24785 (N_24785,N_24592,N_24531);
nor U24786 (N_24786,N_24481,N_24537);
or U24787 (N_24787,N_24552,N_24559);
or U24788 (N_24788,N_24564,N_24466);
and U24789 (N_24789,N_24434,N_24520);
nor U24790 (N_24790,N_24543,N_24447);
or U24791 (N_24791,N_24510,N_24495);
xor U24792 (N_24792,N_24548,N_24450);
nand U24793 (N_24793,N_24449,N_24503);
nand U24794 (N_24794,N_24454,N_24553);
and U24795 (N_24795,N_24497,N_24475);
nand U24796 (N_24796,N_24588,N_24571);
nand U24797 (N_24797,N_24515,N_24405);
or U24798 (N_24798,N_24569,N_24479);
or U24799 (N_24799,N_24422,N_24576);
and U24800 (N_24800,N_24638,N_24725);
nand U24801 (N_24801,N_24628,N_24715);
or U24802 (N_24802,N_24615,N_24740);
xnor U24803 (N_24803,N_24609,N_24711);
or U24804 (N_24804,N_24660,N_24693);
nand U24805 (N_24805,N_24731,N_24643);
and U24806 (N_24806,N_24665,N_24644);
or U24807 (N_24807,N_24761,N_24699);
nand U24808 (N_24808,N_24616,N_24648);
and U24809 (N_24809,N_24694,N_24730);
and U24810 (N_24810,N_24784,N_24776);
nor U24811 (N_24811,N_24650,N_24696);
nor U24812 (N_24812,N_24637,N_24722);
xor U24813 (N_24813,N_24640,N_24619);
nand U24814 (N_24814,N_24797,N_24756);
nand U24815 (N_24815,N_24742,N_24709);
nor U24816 (N_24816,N_24630,N_24683);
and U24817 (N_24817,N_24703,N_24705);
nand U24818 (N_24818,N_24600,N_24765);
nor U24819 (N_24819,N_24758,N_24775);
nand U24820 (N_24820,N_24732,N_24713);
nand U24821 (N_24821,N_24627,N_24779);
and U24822 (N_24822,N_24608,N_24708);
xor U24823 (N_24823,N_24738,N_24624);
or U24824 (N_24824,N_24788,N_24743);
or U24825 (N_24825,N_24639,N_24706);
and U24826 (N_24826,N_24651,N_24714);
xnor U24827 (N_24827,N_24688,N_24757);
or U24828 (N_24828,N_24750,N_24659);
nor U24829 (N_24829,N_24717,N_24735);
or U24830 (N_24830,N_24718,N_24728);
or U24831 (N_24831,N_24759,N_24679);
and U24832 (N_24832,N_24768,N_24747);
or U24833 (N_24833,N_24766,N_24767);
and U24834 (N_24834,N_24701,N_24716);
and U24835 (N_24835,N_24607,N_24692);
nor U24836 (N_24836,N_24762,N_24700);
or U24837 (N_24837,N_24721,N_24791);
and U24838 (N_24838,N_24669,N_24666);
and U24839 (N_24839,N_24601,N_24686);
and U24840 (N_24840,N_24770,N_24667);
or U24841 (N_24841,N_24786,N_24745);
or U24842 (N_24842,N_24685,N_24622);
or U24843 (N_24843,N_24796,N_24687);
nand U24844 (N_24844,N_24654,N_24647);
or U24845 (N_24845,N_24729,N_24611);
xor U24846 (N_24846,N_24751,N_24668);
or U24847 (N_24847,N_24790,N_24748);
nor U24848 (N_24848,N_24646,N_24689);
or U24849 (N_24849,N_24602,N_24771);
nand U24850 (N_24850,N_24749,N_24641);
nand U24851 (N_24851,N_24678,N_24649);
nand U24852 (N_24852,N_24621,N_24795);
xor U24853 (N_24853,N_24617,N_24798);
xor U24854 (N_24854,N_24774,N_24769);
or U24855 (N_24855,N_24632,N_24642);
or U24856 (N_24856,N_24657,N_24746);
or U24857 (N_24857,N_24789,N_24612);
nor U24858 (N_24858,N_24671,N_24794);
nor U24859 (N_24859,N_24737,N_24606);
nand U24860 (N_24860,N_24661,N_24752);
or U24861 (N_24861,N_24623,N_24676);
or U24862 (N_24862,N_24781,N_24635);
and U24863 (N_24863,N_24614,N_24707);
nand U24864 (N_24864,N_24645,N_24773);
nand U24865 (N_24865,N_24658,N_24793);
or U24866 (N_24866,N_24618,N_24777);
xnor U24867 (N_24867,N_24613,N_24697);
nand U24868 (N_24868,N_24763,N_24670);
nor U24869 (N_24869,N_24673,N_24739);
nand U24870 (N_24870,N_24631,N_24655);
and U24871 (N_24871,N_24787,N_24799);
and U24872 (N_24872,N_24755,N_24672);
nand U24873 (N_24873,N_24682,N_24724);
nand U24874 (N_24874,N_24677,N_24690);
and U24875 (N_24875,N_24691,N_24782);
or U24876 (N_24876,N_24727,N_24626);
or U24877 (N_24877,N_24620,N_24663);
nand U24878 (N_24878,N_24726,N_24695);
nor U24879 (N_24879,N_24698,N_24772);
xor U24880 (N_24880,N_24733,N_24605);
or U24881 (N_24881,N_24744,N_24625);
and U24882 (N_24882,N_24610,N_24785);
nand U24883 (N_24883,N_24753,N_24719);
or U24884 (N_24884,N_24629,N_24684);
nand U24885 (N_24885,N_24656,N_24764);
or U24886 (N_24886,N_24792,N_24680);
or U24887 (N_24887,N_24652,N_24780);
xor U24888 (N_24888,N_24664,N_24778);
or U24889 (N_24889,N_24653,N_24741);
and U24890 (N_24890,N_24734,N_24675);
nor U24891 (N_24891,N_24754,N_24603);
nor U24892 (N_24892,N_24633,N_24783);
or U24893 (N_24893,N_24604,N_24674);
and U24894 (N_24894,N_24681,N_24710);
nand U24895 (N_24895,N_24704,N_24736);
xnor U24896 (N_24896,N_24636,N_24662);
nor U24897 (N_24897,N_24712,N_24760);
nor U24898 (N_24898,N_24723,N_24634);
nor U24899 (N_24899,N_24702,N_24720);
xnor U24900 (N_24900,N_24653,N_24715);
or U24901 (N_24901,N_24626,N_24720);
or U24902 (N_24902,N_24789,N_24674);
xnor U24903 (N_24903,N_24727,N_24631);
nor U24904 (N_24904,N_24758,N_24606);
nand U24905 (N_24905,N_24715,N_24710);
and U24906 (N_24906,N_24704,N_24703);
nor U24907 (N_24907,N_24621,N_24604);
and U24908 (N_24908,N_24715,N_24683);
and U24909 (N_24909,N_24744,N_24773);
or U24910 (N_24910,N_24774,N_24768);
and U24911 (N_24911,N_24733,N_24676);
or U24912 (N_24912,N_24763,N_24746);
xor U24913 (N_24913,N_24736,N_24739);
xor U24914 (N_24914,N_24640,N_24768);
or U24915 (N_24915,N_24649,N_24601);
xnor U24916 (N_24916,N_24672,N_24608);
xor U24917 (N_24917,N_24784,N_24714);
xnor U24918 (N_24918,N_24768,N_24739);
xor U24919 (N_24919,N_24660,N_24799);
nor U24920 (N_24920,N_24642,N_24755);
and U24921 (N_24921,N_24689,N_24654);
or U24922 (N_24922,N_24775,N_24768);
or U24923 (N_24923,N_24672,N_24605);
xor U24924 (N_24924,N_24634,N_24773);
and U24925 (N_24925,N_24618,N_24742);
or U24926 (N_24926,N_24791,N_24718);
or U24927 (N_24927,N_24677,N_24749);
nor U24928 (N_24928,N_24778,N_24760);
xor U24929 (N_24929,N_24699,N_24720);
and U24930 (N_24930,N_24764,N_24719);
or U24931 (N_24931,N_24684,N_24768);
nand U24932 (N_24932,N_24738,N_24755);
nand U24933 (N_24933,N_24686,N_24771);
xor U24934 (N_24934,N_24630,N_24659);
and U24935 (N_24935,N_24678,N_24762);
nand U24936 (N_24936,N_24793,N_24706);
or U24937 (N_24937,N_24613,N_24790);
or U24938 (N_24938,N_24769,N_24742);
xor U24939 (N_24939,N_24750,N_24642);
nand U24940 (N_24940,N_24620,N_24793);
nor U24941 (N_24941,N_24753,N_24712);
nand U24942 (N_24942,N_24611,N_24783);
and U24943 (N_24943,N_24743,N_24744);
and U24944 (N_24944,N_24708,N_24683);
and U24945 (N_24945,N_24699,N_24659);
and U24946 (N_24946,N_24780,N_24683);
nand U24947 (N_24947,N_24691,N_24715);
and U24948 (N_24948,N_24727,N_24624);
nor U24949 (N_24949,N_24617,N_24619);
nand U24950 (N_24950,N_24692,N_24721);
or U24951 (N_24951,N_24658,N_24778);
nand U24952 (N_24952,N_24690,N_24670);
nand U24953 (N_24953,N_24668,N_24775);
xnor U24954 (N_24954,N_24704,N_24647);
or U24955 (N_24955,N_24781,N_24750);
nor U24956 (N_24956,N_24780,N_24610);
and U24957 (N_24957,N_24744,N_24791);
xor U24958 (N_24958,N_24605,N_24787);
xnor U24959 (N_24959,N_24695,N_24678);
nand U24960 (N_24960,N_24730,N_24732);
nand U24961 (N_24961,N_24671,N_24759);
and U24962 (N_24962,N_24653,N_24669);
or U24963 (N_24963,N_24744,N_24603);
nor U24964 (N_24964,N_24604,N_24616);
nor U24965 (N_24965,N_24764,N_24784);
nor U24966 (N_24966,N_24786,N_24650);
nor U24967 (N_24967,N_24638,N_24669);
nand U24968 (N_24968,N_24664,N_24629);
or U24969 (N_24969,N_24704,N_24767);
nand U24970 (N_24970,N_24733,N_24753);
and U24971 (N_24971,N_24600,N_24648);
nor U24972 (N_24972,N_24704,N_24669);
nor U24973 (N_24973,N_24761,N_24780);
nand U24974 (N_24974,N_24657,N_24632);
and U24975 (N_24975,N_24693,N_24731);
nand U24976 (N_24976,N_24676,N_24636);
nor U24977 (N_24977,N_24755,N_24717);
or U24978 (N_24978,N_24699,N_24787);
and U24979 (N_24979,N_24698,N_24600);
and U24980 (N_24980,N_24621,N_24717);
nor U24981 (N_24981,N_24787,N_24615);
or U24982 (N_24982,N_24636,N_24715);
and U24983 (N_24983,N_24693,N_24697);
xnor U24984 (N_24984,N_24768,N_24605);
xnor U24985 (N_24985,N_24606,N_24697);
nor U24986 (N_24986,N_24701,N_24659);
nor U24987 (N_24987,N_24718,N_24629);
xnor U24988 (N_24988,N_24703,N_24706);
nor U24989 (N_24989,N_24748,N_24628);
nor U24990 (N_24990,N_24772,N_24620);
nand U24991 (N_24991,N_24749,N_24712);
and U24992 (N_24992,N_24600,N_24784);
nor U24993 (N_24993,N_24789,N_24703);
nor U24994 (N_24994,N_24768,N_24697);
nor U24995 (N_24995,N_24685,N_24719);
xnor U24996 (N_24996,N_24602,N_24617);
nand U24997 (N_24997,N_24774,N_24749);
or U24998 (N_24998,N_24642,N_24713);
nand U24999 (N_24999,N_24638,N_24642);
nand U25000 (N_25000,N_24944,N_24977);
or U25001 (N_25001,N_24889,N_24943);
or U25002 (N_25002,N_24954,N_24939);
or U25003 (N_25003,N_24905,N_24830);
or U25004 (N_25004,N_24911,N_24803);
or U25005 (N_25005,N_24927,N_24877);
nor U25006 (N_25006,N_24873,N_24956);
or U25007 (N_25007,N_24970,N_24916);
xor U25008 (N_25008,N_24884,N_24969);
nand U25009 (N_25009,N_24933,N_24824);
nand U25010 (N_25010,N_24965,N_24828);
nand U25011 (N_25011,N_24880,N_24957);
nor U25012 (N_25012,N_24895,N_24967);
nand U25013 (N_25013,N_24906,N_24855);
and U25014 (N_25014,N_24949,N_24899);
xnor U25015 (N_25015,N_24832,N_24932);
nand U25016 (N_25016,N_24851,N_24990);
nand U25017 (N_25017,N_24812,N_24839);
nand U25018 (N_25018,N_24842,N_24980);
and U25019 (N_25019,N_24940,N_24907);
and U25020 (N_25020,N_24883,N_24972);
nand U25021 (N_25021,N_24868,N_24885);
nand U25022 (N_25022,N_24925,N_24937);
nor U25023 (N_25023,N_24822,N_24867);
and U25024 (N_25024,N_24838,N_24856);
xor U25025 (N_25025,N_24919,N_24909);
or U25026 (N_25026,N_24931,N_24848);
and U25027 (N_25027,N_24902,N_24994);
nor U25028 (N_25028,N_24871,N_24934);
nand U25029 (N_25029,N_24805,N_24979);
nand U25030 (N_25030,N_24804,N_24807);
nor U25031 (N_25031,N_24893,N_24998);
nand U25032 (N_25032,N_24926,N_24922);
and U25033 (N_25033,N_24843,N_24904);
or U25034 (N_25034,N_24814,N_24879);
nand U25035 (N_25035,N_24862,N_24878);
or U25036 (N_25036,N_24890,N_24816);
nor U25037 (N_25037,N_24850,N_24975);
and U25038 (N_25038,N_24835,N_24858);
nand U25039 (N_25039,N_24935,N_24958);
or U25040 (N_25040,N_24959,N_24888);
xnor U25041 (N_25041,N_24984,N_24810);
and U25042 (N_25042,N_24903,N_24921);
xnor U25043 (N_25043,N_24817,N_24892);
and U25044 (N_25044,N_24923,N_24999);
or U25045 (N_25045,N_24968,N_24964);
xnor U25046 (N_25046,N_24955,N_24991);
xor U25047 (N_25047,N_24845,N_24981);
and U25048 (N_25048,N_24811,N_24930);
nor U25049 (N_25049,N_24861,N_24901);
and U25050 (N_25050,N_24813,N_24910);
and U25051 (N_25051,N_24971,N_24819);
or U25052 (N_25052,N_24894,N_24863);
nand U25053 (N_25053,N_24870,N_24900);
or U25054 (N_25054,N_24996,N_24898);
nor U25055 (N_25055,N_24806,N_24823);
xor U25056 (N_25056,N_24820,N_24874);
nor U25057 (N_25057,N_24865,N_24962);
and U25058 (N_25058,N_24946,N_24808);
xor U25059 (N_25059,N_24948,N_24936);
or U25060 (N_25060,N_24827,N_24860);
or U25061 (N_25061,N_24854,N_24876);
nand U25062 (N_25062,N_24815,N_24802);
or U25063 (N_25063,N_24995,N_24897);
nand U25064 (N_25064,N_24840,N_24866);
xnor U25065 (N_25065,N_24978,N_24844);
xnor U25066 (N_25066,N_24825,N_24831);
nand U25067 (N_25067,N_24809,N_24942);
or U25068 (N_25068,N_24872,N_24988);
xor U25069 (N_25069,N_24891,N_24915);
nor U25070 (N_25070,N_24821,N_24961);
nor U25071 (N_25071,N_24896,N_24974);
nand U25072 (N_25072,N_24952,N_24853);
nor U25073 (N_25073,N_24836,N_24881);
and U25074 (N_25074,N_24917,N_24947);
nand U25075 (N_25075,N_24875,N_24800);
nor U25076 (N_25076,N_24920,N_24993);
nor U25077 (N_25077,N_24857,N_24966);
and U25078 (N_25078,N_24989,N_24859);
nand U25079 (N_25079,N_24941,N_24997);
and U25080 (N_25080,N_24918,N_24960);
nand U25081 (N_25081,N_24887,N_24953);
nor U25082 (N_25082,N_24945,N_24976);
xnor U25083 (N_25083,N_24928,N_24864);
nand U25084 (N_25084,N_24837,N_24829);
xor U25085 (N_25085,N_24841,N_24882);
xor U25086 (N_25086,N_24938,N_24950);
nor U25087 (N_25087,N_24818,N_24914);
xnor U25088 (N_25088,N_24834,N_24985);
and U25089 (N_25089,N_24992,N_24924);
xor U25090 (N_25090,N_24886,N_24929);
nor U25091 (N_25091,N_24849,N_24913);
or U25092 (N_25092,N_24982,N_24973);
and U25093 (N_25093,N_24833,N_24983);
and U25094 (N_25094,N_24826,N_24986);
and U25095 (N_25095,N_24847,N_24963);
and U25096 (N_25096,N_24846,N_24852);
nand U25097 (N_25097,N_24987,N_24801);
and U25098 (N_25098,N_24912,N_24951);
or U25099 (N_25099,N_24908,N_24869);
and U25100 (N_25100,N_24892,N_24928);
nand U25101 (N_25101,N_24814,N_24946);
nor U25102 (N_25102,N_24966,N_24987);
or U25103 (N_25103,N_24826,N_24923);
and U25104 (N_25104,N_24927,N_24973);
xor U25105 (N_25105,N_24948,N_24950);
or U25106 (N_25106,N_24867,N_24926);
nor U25107 (N_25107,N_24985,N_24807);
nand U25108 (N_25108,N_24904,N_24943);
or U25109 (N_25109,N_24890,N_24800);
xor U25110 (N_25110,N_24855,N_24831);
or U25111 (N_25111,N_24969,N_24865);
nand U25112 (N_25112,N_24852,N_24913);
or U25113 (N_25113,N_24874,N_24881);
or U25114 (N_25114,N_24910,N_24870);
or U25115 (N_25115,N_24995,N_24998);
and U25116 (N_25116,N_24864,N_24806);
nor U25117 (N_25117,N_24930,N_24836);
nand U25118 (N_25118,N_24942,N_24944);
nor U25119 (N_25119,N_24974,N_24994);
and U25120 (N_25120,N_24974,N_24825);
xnor U25121 (N_25121,N_24895,N_24898);
or U25122 (N_25122,N_24985,N_24833);
nor U25123 (N_25123,N_24949,N_24897);
or U25124 (N_25124,N_24986,N_24803);
nor U25125 (N_25125,N_24970,N_24945);
nand U25126 (N_25126,N_24802,N_24914);
or U25127 (N_25127,N_24980,N_24814);
or U25128 (N_25128,N_24907,N_24891);
nor U25129 (N_25129,N_24907,N_24981);
or U25130 (N_25130,N_24862,N_24944);
and U25131 (N_25131,N_24994,N_24820);
or U25132 (N_25132,N_24971,N_24816);
and U25133 (N_25133,N_24953,N_24897);
or U25134 (N_25134,N_24965,N_24929);
xor U25135 (N_25135,N_24934,N_24841);
or U25136 (N_25136,N_24860,N_24919);
nand U25137 (N_25137,N_24869,N_24901);
xnor U25138 (N_25138,N_24834,N_24908);
and U25139 (N_25139,N_24889,N_24817);
and U25140 (N_25140,N_24863,N_24898);
and U25141 (N_25141,N_24830,N_24984);
nor U25142 (N_25142,N_24874,N_24908);
or U25143 (N_25143,N_24902,N_24962);
or U25144 (N_25144,N_24819,N_24962);
or U25145 (N_25145,N_24810,N_24895);
nand U25146 (N_25146,N_24886,N_24915);
nor U25147 (N_25147,N_24819,N_24878);
xnor U25148 (N_25148,N_24953,N_24991);
or U25149 (N_25149,N_24888,N_24966);
nand U25150 (N_25150,N_24855,N_24923);
and U25151 (N_25151,N_24948,N_24945);
nand U25152 (N_25152,N_24938,N_24853);
xnor U25153 (N_25153,N_24829,N_24883);
xnor U25154 (N_25154,N_24847,N_24969);
nor U25155 (N_25155,N_24814,N_24817);
nor U25156 (N_25156,N_24856,N_24892);
nor U25157 (N_25157,N_24803,N_24999);
and U25158 (N_25158,N_24859,N_24987);
and U25159 (N_25159,N_24920,N_24840);
nand U25160 (N_25160,N_24842,N_24834);
nor U25161 (N_25161,N_24836,N_24887);
and U25162 (N_25162,N_24919,N_24981);
xor U25163 (N_25163,N_24963,N_24873);
xor U25164 (N_25164,N_24821,N_24808);
xor U25165 (N_25165,N_24825,N_24843);
and U25166 (N_25166,N_24843,N_24967);
nor U25167 (N_25167,N_24821,N_24910);
or U25168 (N_25168,N_24801,N_24950);
xor U25169 (N_25169,N_24979,N_24904);
or U25170 (N_25170,N_24858,N_24956);
nor U25171 (N_25171,N_24921,N_24825);
xor U25172 (N_25172,N_24838,N_24999);
or U25173 (N_25173,N_24897,N_24979);
and U25174 (N_25174,N_24945,N_24831);
nor U25175 (N_25175,N_24840,N_24990);
or U25176 (N_25176,N_24945,N_24982);
nor U25177 (N_25177,N_24882,N_24982);
nand U25178 (N_25178,N_24871,N_24920);
or U25179 (N_25179,N_24881,N_24911);
xor U25180 (N_25180,N_24876,N_24888);
nand U25181 (N_25181,N_24995,N_24920);
nor U25182 (N_25182,N_24981,N_24911);
xnor U25183 (N_25183,N_24862,N_24892);
or U25184 (N_25184,N_24894,N_24903);
xor U25185 (N_25185,N_24846,N_24851);
nor U25186 (N_25186,N_24961,N_24926);
nand U25187 (N_25187,N_24911,N_24839);
or U25188 (N_25188,N_24975,N_24810);
nor U25189 (N_25189,N_24924,N_24844);
nor U25190 (N_25190,N_24988,N_24805);
nand U25191 (N_25191,N_24820,N_24945);
and U25192 (N_25192,N_24960,N_24938);
and U25193 (N_25193,N_24963,N_24916);
nor U25194 (N_25194,N_24876,N_24874);
xnor U25195 (N_25195,N_24864,N_24880);
xor U25196 (N_25196,N_24830,N_24865);
nand U25197 (N_25197,N_24958,N_24805);
nor U25198 (N_25198,N_24831,N_24865);
nor U25199 (N_25199,N_24813,N_24830);
or U25200 (N_25200,N_25153,N_25056);
xor U25201 (N_25201,N_25069,N_25101);
and U25202 (N_25202,N_25128,N_25031);
and U25203 (N_25203,N_25065,N_25079);
nor U25204 (N_25204,N_25085,N_25179);
nor U25205 (N_25205,N_25137,N_25162);
nand U25206 (N_25206,N_25189,N_25029);
nand U25207 (N_25207,N_25094,N_25064);
or U25208 (N_25208,N_25049,N_25026);
nor U25209 (N_25209,N_25195,N_25078);
xor U25210 (N_25210,N_25011,N_25135);
xnor U25211 (N_25211,N_25131,N_25111);
nand U25212 (N_25212,N_25199,N_25034);
nor U25213 (N_25213,N_25014,N_25132);
nor U25214 (N_25214,N_25068,N_25134);
nor U25215 (N_25215,N_25122,N_25010);
or U25216 (N_25216,N_25170,N_25192);
nand U25217 (N_25217,N_25114,N_25158);
xnor U25218 (N_25218,N_25177,N_25159);
nor U25219 (N_25219,N_25090,N_25144);
nand U25220 (N_25220,N_25006,N_25053);
and U25221 (N_25221,N_25166,N_25092);
xor U25222 (N_25222,N_25008,N_25002);
and U25223 (N_25223,N_25044,N_25015);
nor U25224 (N_25224,N_25130,N_25081);
xnor U25225 (N_25225,N_25022,N_25040);
nand U25226 (N_25226,N_25075,N_25074);
and U25227 (N_25227,N_25147,N_25196);
or U25228 (N_25228,N_25103,N_25186);
nand U25229 (N_25229,N_25060,N_25136);
nor U25230 (N_25230,N_25193,N_25073);
nor U25231 (N_25231,N_25183,N_25087);
nor U25232 (N_25232,N_25168,N_25003);
xnor U25233 (N_25233,N_25163,N_25188);
xnor U25234 (N_25234,N_25091,N_25184);
xor U25235 (N_25235,N_25061,N_25173);
or U25236 (N_25236,N_25139,N_25127);
or U25237 (N_25237,N_25093,N_25119);
nand U25238 (N_25238,N_25043,N_25080);
nor U25239 (N_25239,N_25005,N_25033);
nand U25240 (N_25240,N_25151,N_25187);
nor U25241 (N_25241,N_25165,N_25112);
and U25242 (N_25242,N_25150,N_25109);
and U25243 (N_25243,N_25190,N_25017);
or U25244 (N_25244,N_25146,N_25138);
nand U25245 (N_25245,N_25126,N_25012);
or U25246 (N_25246,N_25171,N_25095);
or U25247 (N_25247,N_25007,N_25066);
or U25248 (N_25248,N_25098,N_25077);
or U25249 (N_25249,N_25038,N_25105);
and U25250 (N_25250,N_25018,N_25164);
nor U25251 (N_25251,N_25039,N_25057);
nand U25252 (N_25252,N_25013,N_25133);
and U25253 (N_25253,N_25088,N_25113);
or U25254 (N_25254,N_25020,N_25021);
and U25255 (N_25255,N_25016,N_25048);
xor U25256 (N_25256,N_25055,N_25157);
nand U25257 (N_25257,N_25197,N_25161);
or U25258 (N_25258,N_25071,N_25028);
or U25259 (N_25259,N_25032,N_25045);
nor U25260 (N_25260,N_25096,N_25104);
xnor U25261 (N_25261,N_25072,N_25172);
and U25262 (N_25262,N_25052,N_25041);
or U25263 (N_25263,N_25149,N_25009);
nand U25264 (N_25264,N_25050,N_25115);
and U25265 (N_25265,N_25070,N_25102);
xnor U25266 (N_25266,N_25175,N_25194);
or U25267 (N_25267,N_25063,N_25140);
xnor U25268 (N_25268,N_25089,N_25023);
xor U25269 (N_25269,N_25120,N_25154);
or U25270 (N_25270,N_25051,N_25062);
nand U25271 (N_25271,N_25082,N_25110);
or U25272 (N_25272,N_25019,N_25116);
and U25273 (N_25273,N_25097,N_25123);
nor U25274 (N_25274,N_25106,N_25000);
xnor U25275 (N_25275,N_25155,N_25145);
or U25276 (N_25276,N_25037,N_25001);
xor U25277 (N_25277,N_25141,N_25185);
nand U25278 (N_25278,N_25125,N_25121);
and U25279 (N_25279,N_25076,N_25148);
nand U25280 (N_25280,N_25059,N_25047);
nor U25281 (N_25281,N_25124,N_25129);
and U25282 (N_25282,N_25099,N_25046);
xor U25283 (N_25283,N_25191,N_25178);
or U25284 (N_25284,N_25024,N_25004);
xnor U25285 (N_25285,N_25167,N_25058);
nand U25286 (N_25286,N_25117,N_25030);
xor U25287 (N_25287,N_25100,N_25107);
nor U25288 (N_25288,N_25198,N_25181);
xor U25289 (N_25289,N_25036,N_25160);
nand U25290 (N_25290,N_25143,N_25067);
nand U25291 (N_25291,N_25054,N_25142);
nor U25292 (N_25292,N_25156,N_25169);
nor U25293 (N_25293,N_25042,N_25182);
nor U25294 (N_25294,N_25152,N_25174);
and U25295 (N_25295,N_25118,N_25083);
and U25296 (N_25296,N_25027,N_25108);
nand U25297 (N_25297,N_25084,N_25180);
nand U25298 (N_25298,N_25035,N_25025);
or U25299 (N_25299,N_25176,N_25086);
nand U25300 (N_25300,N_25015,N_25048);
nand U25301 (N_25301,N_25155,N_25025);
or U25302 (N_25302,N_25048,N_25021);
or U25303 (N_25303,N_25076,N_25031);
or U25304 (N_25304,N_25146,N_25013);
nand U25305 (N_25305,N_25125,N_25057);
and U25306 (N_25306,N_25160,N_25014);
nand U25307 (N_25307,N_25045,N_25155);
nand U25308 (N_25308,N_25140,N_25073);
nor U25309 (N_25309,N_25152,N_25048);
and U25310 (N_25310,N_25118,N_25187);
xnor U25311 (N_25311,N_25092,N_25165);
nand U25312 (N_25312,N_25003,N_25174);
or U25313 (N_25313,N_25101,N_25118);
xnor U25314 (N_25314,N_25086,N_25093);
and U25315 (N_25315,N_25115,N_25117);
nand U25316 (N_25316,N_25155,N_25187);
xnor U25317 (N_25317,N_25011,N_25118);
or U25318 (N_25318,N_25019,N_25163);
or U25319 (N_25319,N_25052,N_25075);
xnor U25320 (N_25320,N_25087,N_25196);
xnor U25321 (N_25321,N_25013,N_25142);
or U25322 (N_25322,N_25091,N_25002);
and U25323 (N_25323,N_25059,N_25123);
or U25324 (N_25324,N_25132,N_25138);
and U25325 (N_25325,N_25022,N_25177);
nand U25326 (N_25326,N_25178,N_25155);
nand U25327 (N_25327,N_25035,N_25174);
xor U25328 (N_25328,N_25017,N_25042);
nor U25329 (N_25329,N_25193,N_25098);
nor U25330 (N_25330,N_25129,N_25005);
or U25331 (N_25331,N_25017,N_25094);
nand U25332 (N_25332,N_25183,N_25069);
nand U25333 (N_25333,N_25088,N_25161);
xnor U25334 (N_25334,N_25136,N_25126);
or U25335 (N_25335,N_25122,N_25192);
and U25336 (N_25336,N_25010,N_25180);
and U25337 (N_25337,N_25002,N_25046);
xor U25338 (N_25338,N_25133,N_25004);
or U25339 (N_25339,N_25110,N_25023);
nand U25340 (N_25340,N_25124,N_25090);
nand U25341 (N_25341,N_25102,N_25092);
nand U25342 (N_25342,N_25046,N_25057);
or U25343 (N_25343,N_25078,N_25141);
nor U25344 (N_25344,N_25088,N_25056);
and U25345 (N_25345,N_25131,N_25159);
or U25346 (N_25346,N_25071,N_25173);
nor U25347 (N_25347,N_25198,N_25074);
and U25348 (N_25348,N_25060,N_25085);
or U25349 (N_25349,N_25103,N_25179);
nor U25350 (N_25350,N_25014,N_25180);
or U25351 (N_25351,N_25183,N_25014);
nor U25352 (N_25352,N_25137,N_25014);
xor U25353 (N_25353,N_25095,N_25104);
nor U25354 (N_25354,N_25093,N_25195);
or U25355 (N_25355,N_25033,N_25149);
xor U25356 (N_25356,N_25052,N_25088);
nor U25357 (N_25357,N_25107,N_25186);
nand U25358 (N_25358,N_25175,N_25054);
and U25359 (N_25359,N_25172,N_25009);
or U25360 (N_25360,N_25086,N_25032);
nand U25361 (N_25361,N_25066,N_25075);
xnor U25362 (N_25362,N_25078,N_25156);
nand U25363 (N_25363,N_25137,N_25195);
and U25364 (N_25364,N_25140,N_25150);
nor U25365 (N_25365,N_25004,N_25087);
or U25366 (N_25366,N_25036,N_25051);
nand U25367 (N_25367,N_25126,N_25062);
and U25368 (N_25368,N_25062,N_25115);
or U25369 (N_25369,N_25190,N_25162);
nor U25370 (N_25370,N_25078,N_25159);
nand U25371 (N_25371,N_25124,N_25143);
nor U25372 (N_25372,N_25007,N_25005);
xor U25373 (N_25373,N_25014,N_25181);
nor U25374 (N_25374,N_25117,N_25186);
nor U25375 (N_25375,N_25039,N_25070);
nand U25376 (N_25376,N_25064,N_25063);
nand U25377 (N_25377,N_25072,N_25123);
xnor U25378 (N_25378,N_25135,N_25115);
nand U25379 (N_25379,N_25037,N_25158);
or U25380 (N_25380,N_25000,N_25197);
xnor U25381 (N_25381,N_25102,N_25121);
nor U25382 (N_25382,N_25084,N_25003);
xnor U25383 (N_25383,N_25165,N_25047);
or U25384 (N_25384,N_25149,N_25184);
xor U25385 (N_25385,N_25187,N_25173);
and U25386 (N_25386,N_25189,N_25175);
nand U25387 (N_25387,N_25041,N_25093);
nand U25388 (N_25388,N_25178,N_25098);
and U25389 (N_25389,N_25148,N_25110);
nor U25390 (N_25390,N_25171,N_25022);
xnor U25391 (N_25391,N_25161,N_25184);
xor U25392 (N_25392,N_25121,N_25150);
nor U25393 (N_25393,N_25110,N_25195);
nor U25394 (N_25394,N_25061,N_25095);
or U25395 (N_25395,N_25157,N_25093);
nor U25396 (N_25396,N_25060,N_25016);
xnor U25397 (N_25397,N_25125,N_25008);
xnor U25398 (N_25398,N_25148,N_25031);
nand U25399 (N_25399,N_25073,N_25085);
xnor U25400 (N_25400,N_25392,N_25364);
nor U25401 (N_25401,N_25371,N_25314);
xnor U25402 (N_25402,N_25246,N_25344);
and U25403 (N_25403,N_25249,N_25372);
nor U25404 (N_25404,N_25213,N_25339);
or U25405 (N_25405,N_25385,N_25329);
and U25406 (N_25406,N_25304,N_25370);
nand U25407 (N_25407,N_25218,N_25317);
and U25408 (N_25408,N_25353,N_25399);
and U25409 (N_25409,N_25315,N_25226);
nor U25410 (N_25410,N_25210,N_25281);
or U25411 (N_25411,N_25240,N_25328);
nand U25412 (N_25412,N_25336,N_25217);
and U25413 (N_25413,N_25268,N_25312);
nor U25414 (N_25414,N_25236,N_25238);
or U25415 (N_25415,N_25215,N_25365);
xor U25416 (N_25416,N_25342,N_25316);
nor U25417 (N_25417,N_25292,N_25397);
or U25418 (N_25418,N_25333,N_25224);
and U25419 (N_25419,N_25327,N_25274);
or U25420 (N_25420,N_25220,N_25320);
or U25421 (N_25421,N_25255,N_25338);
and U25422 (N_25422,N_25357,N_25299);
or U25423 (N_25423,N_25228,N_25256);
or U25424 (N_25424,N_25324,N_25258);
and U25425 (N_25425,N_25283,N_25261);
or U25426 (N_25426,N_25262,N_25376);
and U25427 (N_25427,N_25251,N_25343);
nand U25428 (N_25428,N_25241,N_25373);
xnor U25429 (N_25429,N_25347,N_25330);
or U25430 (N_25430,N_25264,N_25231);
and U25431 (N_25431,N_25289,N_25230);
or U25432 (N_25432,N_25259,N_25308);
and U25433 (N_25433,N_25222,N_25311);
nor U25434 (N_25434,N_25345,N_25273);
or U25435 (N_25435,N_25363,N_25216);
nor U25436 (N_25436,N_25252,N_25285);
nand U25437 (N_25437,N_25287,N_25243);
and U25438 (N_25438,N_25200,N_25300);
nor U25439 (N_25439,N_25284,N_25297);
and U25440 (N_25440,N_25279,N_25265);
and U25441 (N_25441,N_25248,N_25242);
or U25442 (N_25442,N_25302,N_25352);
or U25443 (N_25443,N_25391,N_25383);
or U25444 (N_25444,N_25233,N_25361);
nand U25445 (N_25445,N_25326,N_25354);
nor U25446 (N_25446,N_25367,N_25253);
nor U25447 (N_25447,N_25204,N_25319);
nor U25448 (N_25448,N_25334,N_25269);
nor U25449 (N_25449,N_25235,N_25305);
xnor U25450 (N_25450,N_25286,N_25267);
and U25451 (N_25451,N_25272,N_25207);
nor U25452 (N_25452,N_25332,N_25229);
nor U25453 (N_25453,N_25377,N_25375);
nor U25454 (N_25454,N_25201,N_25237);
nor U25455 (N_25455,N_25290,N_25394);
xnor U25456 (N_25456,N_25244,N_25395);
nand U25457 (N_25457,N_25227,N_25366);
nand U25458 (N_25458,N_25260,N_25348);
nand U25459 (N_25459,N_25296,N_25208);
xnor U25460 (N_25460,N_25380,N_25250);
and U25461 (N_25461,N_25379,N_25214);
nand U25462 (N_25462,N_25277,N_25387);
xor U25463 (N_25463,N_25203,N_25359);
and U25464 (N_25464,N_25303,N_25335);
nor U25465 (N_25465,N_25301,N_25356);
or U25466 (N_25466,N_25280,N_25288);
nor U25467 (N_25467,N_25358,N_25234);
or U25468 (N_25468,N_25398,N_25221);
xor U25469 (N_25469,N_25225,N_25325);
nor U25470 (N_25470,N_25396,N_25331);
and U25471 (N_25471,N_25205,N_25266);
nand U25472 (N_25472,N_25349,N_25275);
or U25473 (N_25473,N_25294,N_25389);
and U25474 (N_25474,N_25374,N_25378);
or U25475 (N_25475,N_25346,N_25382);
xnor U25476 (N_25476,N_25271,N_25341);
xor U25477 (N_25477,N_25270,N_25355);
and U25478 (N_25478,N_25351,N_25209);
or U25479 (N_25479,N_25337,N_25291);
and U25480 (N_25480,N_25295,N_25340);
and U25481 (N_25481,N_25368,N_25239);
or U25482 (N_25482,N_25257,N_25263);
nor U25483 (N_25483,N_25323,N_25212);
xnor U25484 (N_25484,N_25393,N_25219);
and U25485 (N_25485,N_25322,N_25381);
nor U25486 (N_25486,N_25362,N_25202);
xor U25487 (N_25487,N_25276,N_25388);
and U25488 (N_25488,N_25247,N_25386);
and U25489 (N_25489,N_25390,N_25321);
or U25490 (N_25490,N_25369,N_25298);
xnor U25491 (N_25491,N_25318,N_25360);
xor U25492 (N_25492,N_25282,N_25211);
xnor U25493 (N_25493,N_25223,N_25278);
nor U25494 (N_25494,N_25232,N_25313);
xor U25495 (N_25495,N_25309,N_25254);
xor U25496 (N_25496,N_25350,N_25245);
xor U25497 (N_25497,N_25206,N_25310);
nand U25498 (N_25498,N_25307,N_25293);
xnor U25499 (N_25499,N_25384,N_25306);
and U25500 (N_25500,N_25381,N_25395);
nor U25501 (N_25501,N_25313,N_25333);
xnor U25502 (N_25502,N_25214,N_25210);
xor U25503 (N_25503,N_25382,N_25344);
nor U25504 (N_25504,N_25302,N_25270);
nand U25505 (N_25505,N_25273,N_25302);
nor U25506 (N_25506,N_25300,N_25260);
xor U25507 (N_25507,N_25241,N_25272);
xor U25508 (N_25508,N_25234,N_25225);
nand U25509 (N_25509,N_25339,N_25377);
nand U25510 (N_25510,N_25268,N_25300);
nor U25511 (N_25511,N_25258,N_25238);
nor U25512 (N_25512,N_25326,N_25301);
and U25513 (N_25513,N_25284,N_25345);
nand U25514 (N_25514,N_25340,N_25223);
or U25515 (N_25515,N_25396,N_25359);
or U25516 (N_25516,N_25390,N_25341);
and U25517 (N_25517,N_25384,N_25269);
nor U25518 (N_25518,N_25326,N_25388);
nand U25519 (N_25519,N_25346,N_25333);
nor U25520 (N_25520,N_25302,N_25348);
and U25521 (N_25521,N_25337,N_25349);
or U25522 (N_25522,N_25217,N_25351);
xor U25523 (N_25523,N_25306,N_25215);
xor U25524 (N_25524,N_25384,N_25397);
xnor U25525 (N_25525,N_25370,N_25244);
or U25526 (N_25526,N_25243,N_25327);
nor U25527 (N_25527,N_25280,N_25290);
nor U25528 (N_25528,N_25287,N_25210);
xnor U25529 (N_25529,N_25387,N_25210);
and U25530 (N_25530,N_25392,N_25365);
nor U25531 (N_25531,N_25277,N_25358);
or U25532 (N_25532,N_25347,N_25354);
xnor U25533 (N_25533,N_25350,N_25275);
or U25534 (N_25534,N_25217,N_25318);
nand U25535 (N_25535,N_25376,N_25238);
and U25536 (N_25536,N_25331,N_25254);
nand U25537 (N_25537,N_25383,N_25349);
xor U25538 (N_25538,N_25366,N_25390);
nor U25539 (N_25539,N_25326,N_25345);
nand U25540 (N_25540,N_25243,N_25367);
nand U25541 (N_25541,N_25265,N_25351);
nand U25542 (N_25542,N_25258,N_25268);
nor U25543 (N_25543,N_25351,N_25315);
nand U25544 (N_25544,N_25220,N_25233);
or U25545 (N_25545,N_25280,N_25249);
and U25546 (N_25546,N_25244,N_25305);
or U25547 (N_25547,N_25326,N_25394);
and U25548 (N_25548,N_25393,N_25395);
nor U25549 (N_25549,N_25217,N_25369);
xor U25550 (N_25550,N_25289,N_25363);
nor U25551 (N_25551,N_25305,N_25321);
and U25552 (N_25552,N_25311,N_25309);
xor U25553 (N_25553,N_25338,N_25394);
or U25554 (N_25554,N_25333,N_25342);
and U25555 (N_25555,N_25292,N_25319);
or U25556 (N_25556,N_25387,N_25333);
nor U25557 (N_25557,N_25247,N_25394);
and U25558 (N_25558,N_25225,N_25256);
nor U25559 (N_25559,N_25216,N_25285);
nand U25560 (N_25560,N_25331,N_25281);
nor U25561 (N_25561,N_25253,N_25224);
nor U25562 (N_25562,N_25379,N_25317);
nand U25563 (N_25563,N_25364,N_25201);
xor U25564 (N_25564,N_25270,N_25372);
xor U25565 (N_25565,N_25247,N_25340);
xnor U25566 (N_25566,N_25382,N_25265);
nor U25567 (N_25567,N_25313,N_25388);
nand U25568 (N_25568,N_25332,N_25373);
nor U25569 (N_25569,N_25311,N_25327);
xnor U25570 (N_25570,N_25375,N_25361);
xnor U25571 (N_25571,N_25339,N_25217);
or U25572 (N_25572,N_25220,N_25297);
or U25573 (N_25573,N_25227,N_25383);
nand U25574 (N_25574,N_25359,N_25390);
or U25575 (N_25575,N_25272,N_25288);
and U25576 (N_25576,N_25337,N_25324);
nand U25577 (N_25577,N_25312,N_25304);
nand U25578 (N_25578,N_25216,N_25370);
nand U25579 (N_25579,N_25331,N_25256);
and U25580 (N_25580,N_25223,N_25222);
nor U25581 (N_25581,N_25268,N_25385);
xnor U25582 (N_25582,N_25204,N_25231);
nor U25583 (N_25583,N_25319,N_25315);
or U25584 (N_25584,N_25244,N_25230);
or U25585 (N_25585,N_25328,N_25323);
xnor U25586 (N_25586,N_25305,N_25260);
or U25587 (N_25587,N_25209,N_25254);
or U25588 (N_25588,N_25322,N_25262);
nand U25589 (N_25589,N_25272,N_25337);
nor U25590 (N_25590,N_25329,N_25360);
nand U25591 (N_25591,N_25268,N_25225);
xnor U25592 (N_25592,N_25227,N_25279);
or U25593 (N_25593,N_25213,N_25378);
or U25594 (N_25594,N_25271,N_25263);
or U25595 (N_25595,N_25276,N_25266);
and U25596 (N_25596,N_25206,N_25336);
xor U25597 (N_25597,N_25322,N_25275);
or U25598 (N_25598,N_25365,N_25355);
xnor U25599 (N_25599,N_25211,N_25218);
xor U25600 (N_25600,N_25440,N_25429);
xor U25601 (N_25601,N_25550,N_25479);
or U25602 (N_25602,N_25433,N_25453);
and U25603 (N_25603,N_25447,N_25452);
and U25604 (N_25604,N_25516,N_25512);
nand U25605 (N_25605,N_25408,N_25411);
nand U25606 (N_25606,N_25410,N_25533);
nor U25607 (N_25607,N_25458,N_25464);
or U25608 (N_25608,N_25445,N_25490);
xor U25609 (N_25609,N_25513,N_25559);
xnor U25610 (N_25610,N_25517,N_25427);
nand U25611 (N_25611,N_25463,N_25582);
nor U25612 (N_25612,N_25591,N_25483);
and U25613 (N_25613,N_25400,N_25540);
xnor U25614 (N_25614,N_25537,N_25567);
nand U25615 (N_25615,N_25545,N_25405);
nand U25616 (N_25616,N_25521,N_25572);
or U25617 (N_25617,N_25457,N_25450);
and U25618 (N_25618,N_25565,N_25546);
nor U25619 (N_25619,N_25486,N_25439);
nand U25620 (N_25620,N_25402,N_25588);
or U25621 (N_25621,N_25524,N_25414);
nand U25622 (N_25622,N_25469,N_25580);
and U25623 (N_25623,N_25503,N_25417);
nand U25624 (N_25624,N_25431,N_25574);
nor U25625 (N_25625,N_25554,N_25571);
or U25626 (N_25626,N_25534,N_25525);
nor U25627 (N_25627,N_25584,N_25530);
nand U25628 (N_25628,N_25573,N_25563);
or U25629 (N_25629,N_25598,N_25586);
nor U25630 (N_25630,N_25501,N_25462);
nor U25631 (N_25631,N_25555,N_25515);
and U25632 (N_25632,N_25575,N_25485);
or U25633 (N_25633,N_25599,N_25423);
nand U25634 (N_25634,N_25422,N_25587);
and U25635 (N_25635,N_25419,N_25560);
nor U25636 (N_25636,N_25549,N_25435);
nor U25637 (N_25637,N_25589,N_25441);
xnor U25638 (N_25638,N_25502,N_25558);
nand U25639 (N_25639,N_25562,N_25442);
nand U25640 (N_25640,N_25475,N_25413);
and U25641 (N_25641,N_25471,N_25594);
nand U25642 (N_25642,N_25528,N_25518);
xnor U25643 (N_25643,N_25566,N_25480);
or U25644 (N_25644,N_25454,N_25551);
xnor U25645 (N_25645,N_25428,N_25597);
nand U25646 (N_25646,N_25596,N_25478);
and U25647 (N_25647,N_25590,N_25465);
or U25648 (N_25648,N_25509,N_25544);
nor U25649 (N_25649,N_25552,N_25569);
nand U25650 (N_25650,N_25425,N_25407);
and U25651 (N_25651,N_25477,N_25522);
or U25652 (N_25652,N_25581,N_25496);
xnor U25653 (N_25653,N_25482,N_25493);
and U25654 (N_25654,N_25556,N_25514);
or U25655 (N_25655,N_25476,N_25424);
and U25656 (N_25656,N_25532,N_25430);
nor U25657 (N_25657,N_25561,N_25455);
nand U25658 (N_25658,N_25473,N_25459);
and U25659 (N_25659,N_25578,N_25487);
nor U25660 (N_25660,N_25474,N_25436);
nor U25661 (N_25661,N_25527,N_25461);
nand U25662 (N_25662,N_25470,N_25548);
and U25663 (N_25663,N_25499,N_25595);
xnor U25664 (N_25664,N_25507,N_25446);
or U25665 (N_25665,N_25508,N_25564);
and U25666 (N_25666,N_25404,N_25495);
nand U25667 (N_25667,N_25504,N_25531);
nand U25668 (N_25668,N_25494,N_25543);
nand U25669 (N_25669,N_25505,N_25570);
and U25670 (N_25670,N_25557,N_25438);
xor U25671 (N_25671,N_25497,N_25539);
nand U25672 (N_25672,N_25541,N_25466);
and U25673 (N_25673,N_25488,N_25510);
and U25674 (N_25674,N_25547,N_25526);
and U25675 (N_25675,N_25498,N_25536);
xnor U25676 (N_25676,N_25506,N_25535);
nor U25677 (N_25677,N_25500,N_25523);
xor U25678 (N_25678,N_25472,N_25443);
xor U25679 (N_25679,N_25401,N_25481);
nand U25680 (N_25680,N_25538,N_25491);
nor U25681 (N_25681,N_25418,N_25489);
nor U25682 (N_25682,N_25492,N_25511);
nor U25683 (N_25683,N_25520,N_25592);
xnor U25684 (N_25684,N_25593,N_25529);
xor U25685 (N_25685,N_25468,N_25406);
xnor U25686 (N_25686,N_25448,N_25460);
nor U25687 (N_25687,N_25409,N_25542);
and U25688 (N_25688,N_25412,N_25420);
and U25689 (N_25689,N_25467,N_25585);
xor U25690 (N_25690,N_25583,N_25415);
xor U25691 (N_25691,N_25426,N_25577);
nor U25692 (N_25692,N_25434,N_25444);
xnor U25693 (N_25693,N_25553,N_25451);
nor U25694 (N_25694,N_25576,N_25484);
nor U25695 (N_25695,N_25456,N_25568);
nor U25696 (N_25696,N_25579,N_25432);
or U25697 (N_25697,N_25519,N_25449);
nand U25698 (N_25698,N_25437,N_25421);
and U25699 (N_25699,N_25416,N_25403);
xnor U25700 (N_25700,N_25536,N_25438);
or U25701 (N_25701,N_25500,N_25487);
nor U25702 (N_25702,N_25551,N_25564);
and U25703 (N_25703,N_25583,N_25558);
xnor U25704 (N_25704,N_25469,N_25534);
nor U25705 (N_25705,N_25449,N_25442);
xor U25706 (N_25706,N_25433,N_25599);
xnor U25707 (N_25707,N_25550,N_25498);
or U25708 (N_25708,N_25527,N_25579);
nand U25709 (N_25709,N_25542,N_25552);
nand U25710 (N_25710,N_25540,N_25551);
or U25711 (N_25711,N_25586,N_25474);
nand U25712 (N_25712,N_25491,N_25466);
nor U25713 (N_25713,N_25435,N_25547);
and U25714 (N_25714,N_25466,N_25430);
nand U25715 (N_25715,N_25562,N_25429);
or U25716 (N_25716,N_25559,N_25436);
or U25717 (N_25717,N_25509,N_25466);
nor U25718 (N_25718,N_25445,N_25475);
xnor U25719 (N_25719,N_25460,N_25466);
and U25720 (N_25720,N_25435,N_25474);
xor U25721 (N_25721,N_25430,N_25569);
or U25722 (N_25722,N_25571,N_25513);
or U25723 (N_25723,N_25521,N_25488);
nor U25724 (N_25724,N_25583,N_25425);
and U25725 (N_25725,N_25588,N_25553);
xnor U25726 (N_25726,N_25517,N_25583);
nor U25727 (N_25727,N_25524,N_25440);
xnor U25728 (N_25728,N_25556,N_25472);
nand U25729 (N_25729,N_25475,N_25559);
nand U25730 (N_25730,N_25590,N_25533);
nand U25731 (N_25731,N_25551,N_25445);
nand U25732 (N_25732,N_25515,N_25554);
and U25733 (N_25733,N_25544,N_25465);
nor U25734 (N_25734,N_25454,N_25405);
and U25735 (N_25735,N_25541,N_25482);
and U25736 (N_25736,N_25521,N_25531);
or U25737 (N_25737,N_25452,N_25519);
nor U25738 (N_25738,N_25412,N_25422);
nor U25739 (N_25739,N_25543,N_25526);
and U25740 (N_25740,N_25578,N_25574);
and U25741 (N_25741,N_25460,N_25503);
nand U25742 (N_25742,N_25515,N_25418);
xnor U25743 (N_25743,N_25426,N_25514);
xor U25744 (N_25744,N_25485,N_25572);
nand U25745 (N_25745,N_25474,N_25509);
xnor U25746 (N_25746,N_25581,N_25543);
xnor U25747 (N_25747,N_25425,N_25527);
or U25748 (N_25748,N_25581,N_25414);
or U25749 (N_25749,N_25401,N_25457);
nand U25750 (N_25750,N_25546,N_25513);
and U25751 (N_25751,N_25544,N_25557);
or U25752 (N_25752,N_25521,N_25409);
nor U25753 (N_25753,N_25532,N_25537);
nor U25754 (N_25754,N_25533,N_25462);
nand U25755 (N_25755,N_25400,N_25402);
xor U25756 (N_25756,N_25570,N_25450);
nand U25757 (N_25757,N_25545,N_25543);
nor U25758 (N_25758,N_25470,N_25418);
nand U25759 (N_25759,N_25478,N_25541);
and U25760 (N_25760,N_25403,N_25578);
nand U25761 (N_25761,N_25470,N_25485);
and U25762 (N_25762,N_25418,N_25475);
and U25763 (N_25763,N_25514,N_25552);
xor U25764 (N_25764,N_25453,N_25519);
xnor U25765 (N_25765,N_25507,N_25532);
or U25766 (N_25766,N_25476,N_25521);
nor U25767 (N_25767,N_25527,N_25553);
xnor U25768 (N_25768,N_25494,N_25409);
or U25769 (N_25769,N_25488,N_25411);
and U25770 (N_25770,N_25427,N_25431);
xor U25771 (N_25771,N_25493,N_25579);
nor U25772 (N_25772,N_25564,N_25437);
or U25773 (N_25773,N_25578,N_25492);
or U25774 (N_25774,N_25518,N_25584);
nand U25775 (N_25775,N_25493,N_25581);
nand U25776 (N_25776,N_25597,N_25488);
nand U25777 (N_25777,N_25445,N_25411);
or U25778 (N_25778,N_25595,N_25438);
nand U25779 (N_25779,N_25516,N_25520);
xnor U25780 (N_25780,N_25573,N_25501);
and U25781 (N_25781,N_25589,N_25499);
nand U25782 (N_25782,N_25476,N_25531);
or U25783 (N_25783,N_25436,N_25510);
nor U25784 (N_25784,N_25442,N_25426);
nor U25785 (N_25785,N_25498,N_25489);
xnor U25786 (N_25786,N_25585,N_25502);
or U25787 (N_25787,N_25447,N_25424);
nand U25788 (N_25788,N_25507,N_25599);
nor U25789 (N_25789,N_25493,N_25569);
nor U25790 (N_25790,N_25526,N_25522);
nor U25791 (N_25791,N_25421,N_25553);
nand U25792 (N_25792,N_25484,N_25520);
or U25793 (N_25793,N_25458,N_25484);
nand U25794 (N_25794,N_25515,N_25575);
nand U25795 (N_25795,N_25555,N_25508);
nand U25796 (N_25796,N_25470,N_25509);
nor U25797 (N_25797,N_25546,N_25439);
nor U25798 (N_25798,N_25532,N_25556);
or U25799 (N_25799,N_25538,N_25578);
and U25800 (N_25800,N_25667,N_25658);
xor U25801 (N_25801,N_25645,N_25639);
xnor U25802 (N_25802,N_25782,N_25646);
or U25803 (N_25803,N_25792,N_25612);
or U25804 (N_25804,N_25758,N_25685);
nand U25805 (N_25805,N_25749,N_25738);
nor U25806 (N_25806,N_25743,N_25779);
nor U25807 (N_25807,N_25784,N_25729);
nor U25808 (N_25808,N_25671,N_25746);
and U25809 (N_25809,N_25772,N_25689);
nand U25810 (N_25810,N_25603,N_25630);
xor U25811 (N_25811,N_25794,N_25723);
xnor U25812 (N_25812,N_25715,N_25732);
xnor U25813 (N_25813,N_25619,N_25608);
nand U25814 (N_25814,N_25727,N_25662);
or U25815 (N_25815,N_25640,N_25678);
nor U25816 (N_25816,N_25707,N_25780);
nor U25817 (N_25817,N_25788,N_25759);
nand U25818 (N_25818,N_25720,N_25711);
nand U25819 (N_25819,N_25634,N_25781);
nor U25820 (N_25820,N_25740,N_25675);
nor U25821 (N_25821,N_25756,N_25760);
or U25822 (N_25822,N_25696,N_25726);
xor U25823 (N_25823,N_25752,N_25697);
and U25824 (N_25824,N_25631,N_25652);
nor U25825 (N_25825,N_25627,N_25773);
nor U25826 (N_25826,N_25648,N_25791);
nor U25827 (N_25827,N_25618,N_25763);
xnor U25828 (N_25828,N_25668,N_25702);
or U25829 (N_25829,N_25692,N_25680);
or U25830 (N_25830,N_25797,N_25602);
xnor U25831 (N_25831,N_25736,N_25786);
xor U25832 (N_25832,N_25796,N_25799);
and U25833 (N_25833,N_25638,N_25774);
nor U25834 (N_25834,N_25771,N_25798);
xor U25835 (N_25835,N_25664,N_25705);
xor U25836 (N_25836,N_25653,N_25694);
nor U25837 (N_25837,N_25670,N_25649);
and U25838 (N_25838,N_25703,N_25604);
xnor U25839 (N_25839,N_25714,N_25617);
or U25840 (N_25840,N_25725,N_25679);
nor U25841 (N_25841,N_25625,N_25641);
and U25842 (N_25842,N_25745,N_25693);
nand U25843 (N_25843,N_25783,N_25613);
and U25844 (N_25844,N_25721,N_25684);
nor U25845 (N_25845,N_25632,N_25644);
nor U25846 (N_25846,N_25778,N_25650);
and U25847 (N_25847,N_25691,N_25657);
and U25848 (N_25848,N_25708,N_25659);
and U25849 (N_25849,N_25739,N_25636);
and U25850 (N_25850,N_25751,N_25677);
xnor U25851 (N_25851,N_25734,N_25742);
nor U25852 (N_25852,N_25666,N_25795);
and U25853 (N_25853,N_25615,N_25624);
and U25854 (N_25854,N_25635,N_25610);
nand U25855 (N_25855,N_25651,N_25607);
or U25856 (N_25856,N_25704,N_25660);
nor U25857 (N_25857,N_25637,N_25755);
nor U25858 (N_25858,N_25601,N_25761);
and U25859 (N_25859,N_25750,N_25673);
xnor U25860 (N_25860,N_25767,N_25698);
xor U25861 (N_25861,N_25633,N_25661);
xor U25862 (N_25862,N_25728,N_25699);
and U25863 (N_25863,N_25765,N_25719);
and U25864 (N_25864,N_25777,N_25626);
and U25865 (N_25865,N_25656,N_25776);
nor U25866 (N_25866,N_25762,N_25716);
and U25867 (N_25867,N_25600,N_25616);
xor U25868 (N_25868,N_25672,N_25712);
nor U25869 (N_25869,N_25695,N_25775);
or U25870 (N_25870,N_25622,N_25713);
and U25871 (N_25871,N_25688,N_25787);
and U25872 (N_25872,N_25744,N_25676);
and U25873 (N_25873,N_25674,N_25690);
nand U25874 (N_25874,N_25754,N_25621);
nand U25875 (N_25875,N_25733,N_25709);
nor U25876 (N_25876,N_25669,N_25665);
and U25877 (N_25877,N_25741,N_25768);
or U25878 (N_25878,N_25647,N_25683);
xor U25879 (N_25879,N_25700,N_25682);
or U25880 (N_25880,N_25737,N_25785);
nor U25881 (N_25881,N_25718,N_25764);
nor U25882 (N_25882,N_25611,N_25717);
nand U25883 (N_25883,N_25628,N_25753);
or U25884 (N_25884,N_25731,N_25793);
xnor U25885 (N_25885,N_25642,N_25735);
or U25886 (N_25886,N_25663,N_25706);
xor U25887 (N_25887,N_25605,N_25757);
or U25888 (N_25888,N_25769,N_25681);
or U25889 (N_25889,N_25701,N_25790);
or U25890 (N_25890,N_25609,N_25748);
and U25891 (N_25891,N_25614,N_25606);
and U25892 (N_25892,N_25724,N_25687);
nor U25893 (N_25893,N_25654,N_25629);
nor U25894 (N_25894,N_25620,N_25789);
nor U25895 (N_25895,N_25730,N_25623);
and U25896 (N_25896,N_25722,N_25710);
nand U25897 (N_25897,N_25766,N_25643);
and U25898 (N_25898,N_25747,N_25770);
and U25899 (N_25899,N_25655,N_25686);
or U25900 (N_25900,N_25650,N_25661);
nor U25901 (N_25901,N_25762,N_25730);
xnor U25902 (N_25902,N_25784,N_25706);
or U25903 (N_25903,N_25660,N_25796);
nand U25904 (N_25904,N_25637,N_25608);
nor U25905 (N_25905,N_25660,N_25773);
or U25906 (N_25906,N_25672,N_25643);
nand U25907 (N_25907,N_25697,N_25643);
and U25908 (N_25908,N_25742,N_25601);
and U25909 (N_25909,N_25688,N_25607);
xor U25910 (N_25910,N_25618,N_25654);
nand U25911 (N_25911,N_25721,N_25630);
or U25912 (N_25912,N_25785,N_25659);
nor U25913 (N_25913,N_25728,N_25690);
and U25914 (N_25914,N_25600,N_25606);
and U25915 (N_25915,N_25672,N_25673);
or U25916 (N_25916,N_25614,N_25757);
or U25917 (N_25917,N_25716,N_25770);
nand U25918 (N_25918,N_25795,N_25675);
nor U25919 (N_25919,N_25785,N_25618);
xor U25920 (N_25920,N_25660,N_25736);
xor U25921 (N_25921,N_25750,N_25636);
nand U25922 (N_25922,N_25609,N_25675);
and U25923 (N_25923,N_25735,N_25773);
nand U25924 (N_25924,N_25711,N_25686);
nand U25925 (N_25925,N_25616,N_25797);
or U25926 (N_25926,N_25645,N_25623);
nand U25927 (N_25927,N_25669,N_25754);
xor U25928 (N_25928,N_25716,N_25690);
nand U25929 (N_25929,N_25656,N_25614);
or U25930 (N_25930,N_25608,N_25709);
nor U25931 (N_25931,N_25768,N_25795);
xnor U25932 (N_25932,N_25665,N_25796);
nand U25933 (N_25933,N_25714,N_25695);
or U25934 (N_25934,N_25749,N_25647);
and U25935 (N_25935,N_25665,N_25654);
or U25936 (N_25936,N_25709,N_25720);
nand U25937 (N_25937,N_25744,N_25718);
and U25938 (N_25938,N_25749,N_25710);
and U25939 (N_25939,N_25709,N_25667);
nand U25940 (N_25940,N_25685,N_25698);
or U25941 (N_25941,N_25747,N_25773);
nor U25942 (N_25942,N_25702,N_25674);
and U25943 (N_25943,N_25620,N_25621);
xnor U25944 (N_25944,N_25767,N_25656);
xnor U25945 (N_25945,N_25768,N_25702);
nor U25946 (N_25946,N_25704,N_25720);
nor U25947 (N_25947,N_25729,N_25704);
nor U25948 (N_25948,N_25772,N_25776);
xor U25949 (N_25949,N_25727,N_25708);
or U25950 (N_25950,N_25673,N_25762);
xnor U25951 (N_25951,N_25776,N_25693);
or U25952 (N_25952,N_25649,N_25607);
or U25953 (N_25953,N_25681,N_25624);
nand U25954 (N_25954,N_25762,N_25789);
and U25955 (N_25955,N_25774,N_25778);
and U25956 (N_25956,N_25668,N_25725);
or U25957 (N_25957,N_25791,N_25751);
or U25958 (N_25958,N_25767,N_25774);
or U25959 (N_25959,N_25665,N_25692);
nor U25960 (N_25960,N_25605,N_25740);
nor U25961 (N_25961,N_25738,N_25753);
nor U25962 (N_25962,N_25695,N_25657);
or U25963 (N_25963,N_25786,N_25636);
or U25964 (N_25964,N_25600,N_25741);
nand U25965 (N_25965,N_25631,N_25720);
nand U25966 (N_25966,N_25640,N_25708);
xor U25967 (N_25967,N_25763,N_25741);
nand U25968 (N_25968,N_25698,N_25611);
xnor U25969 (N_25969,N_25695,N_25634);
nor U25970 (N_25970,N_25677,N_25759);
nor U25971 (N_25971,N_25760,N_25749);
xor U25972 (N_25972,N_25757,N_25791);
nor U25973 (N_25973,N_25607,N_25728);
or U25974 (N_25974,N_25642,N_25733);
or U25975 (N_25975,N_25674,N_25776);
nor U25976 (N_25976,N_25738,N_25721);
nor U25977 (N_25977,N_25653,N_25735);
or U25978 (N_25978,N_25625,N_25720);
nand U25979 (N_25979,N_25753,N_25708);
nor U25980 (N_25980,N_25647,N_25696);
or U25981 (N_25981,N_25699,N_25718);
and U25982 (N_25982,N_25718,N_25600);
and U25983 (N_25983,N_25618,N_25732);
or U25984 (N_25984,N_25794,N_25607);
xnor U25985 (N_25985,N_25610,N_25662);
nor U25986 (N_25986,N_25644,N_25712);
nand U25987 (N_25987,N_25635,N_25623);
nand U25988 (N_25988,N_25634,N_25761);
nand U25989 (N_25989,N_25743,N_25788);
and U25990 (N_25990,N_25656,N_25759);
and U25991 (N_25991,N_25715,N_25778);
nor U25992 (N_25992,N_25615,N_25662);
nand U25993 (N_25993,N_25769,N_25747);
and U25994 (N_25994,N_25623,N_25601);
nand U25995 (N_25995,N_25782,N_25628);
nand U25996 (N_25996,N_25755,N_25611);
nand U25997 (N_25997,N_25798,N_25601);
or U25998 (N_25998,N_25655,N_25763);
nand U25999 (N_25999,N_25614,N_25721);
and U26000 (N_26000,N_25861,N_25813);
and U26001 (N_26001,N_25835,N_25933);
or U26002 (N_26002,N_25930,N_25836);
nor U26003 (N_26003,N_25804,N_25822);
or U26004 (N_26004,N_25906,N_25845);
and U26005 (N_26005,N_25849,N_25989);
xnor U26006 (N_26006,N_25946,N_25843);
or U26007 (N_26007,N_25840,N_25968);
and U26008 (N_26008,N_25934,N_25913);
nand U26009 (N_26009,N_25802,N_25868);
or U26010 (N_26010,N_25842,N_25931);
xor U26011 (N_26011,N_25898,N_25877);
xnor U26012 (N_26012,N_25872,N_25812);
or U26013 (N_26013,N_25884,N_25829);
and U26014 (N_26014,N_25928,N_25800);
nand U26015 (N_26015,N_25981,N_25823);
and U26016 (N_26016,N_25927,N_25808);
xnor U26017 (N_26017,N_25972,N_25962);
xor U26018 (N_26018,N_25963,N_25859);
or U26019 (N_26019,N_25866,N_25879);
or U26020 (N_26020,N_25937,N_25995);
nor U26021 (N_26021,N_25863,N_25892);
xor U26022 (N_26022,N_25851,N_25971);
nand U26023 (N_26023,N_25807,N_25926);
nor U26024 (N_26024,N_25905,N_25890);
nand U26025 (N_26025,N_25991,N_25824);
or U26026 (N_26026,N_25955,N_25816);
and U26027 (N_26027,N_25977,N_25894);
nor U26028 (N_26028,N_25875,N_25837);
xnor U26029 (N_26029,N_25860,N_25865);
and U26030 (N_26030,N_25904,N_25909);
and U26031 (N_26031,N_25952,N_25954);
and U26032 (N_26032,N_25878,N_25832);
nand U26033 (N_26033,N_25957,N_25965);
nand U26034 (N_26034,N_25847,N_25895);
xnor U26035 (N_26035,N_25925,N_25960);
and U26036 (N_26036,N_25964,N_25899);
xor U26037 (N_26037,N_25876,N_25817);
and U26038 (N_26038,N_25803,N_25915);
nor U26039 (N_26039,N_25929,N_25916);
and U26040 (N_26040,N_25914,N_25932);
xor U26041 (N_26041,N_25819,N_25844);
or U26042 (N_26042,N_25923,N_25867);
xor U26043 (N_26043,N_25940,N_25978);
nor U26044 (N_26044,N_25882,N_25982);
and U26045 (N_26045,N_25900,N_25936);
and U26046 (N_26046,N_25838,N_25880);
or U26047 (N_26047,N_25912,N_25959);
and U26048 (N_26048,N_25948,N_25881);
or U26049 (N_26049,N_25967,N_25987);
nand U26050 (N_26050,N_25821,N_25870);
or U26051 (N_26051,N_25846,N_25958);
nand U26052 (N_26052,N_25961,N_25801);
xor U26053 (N_26053,N_25918,N_25947);
nand U26054 (N_26054,N_25953,N_25887);
xor U26055 (N_26055,N_25970,N_25924);
and U26056 (N_26056,N_25980,N_25901);
or U26057 (N_26057,N_25984,N_25950);
nand U26058 (N_26058,N_25889,N_25862);
or U26059 (N_26059,N_25814,N_25854);
nand U26060 (N_26060,N_25922,N_25897);
or U26061 (N_26061,N_25852,N_25983);
nor U26062 (N_26062,N_25920,N_25805);
and U26063 (N_26063,N_25966,N_25839);
nor U26064 (N_26064,N_25919,N_25874);
and U26065 (N_26065,N_25818,N_25858);
nand U26066 (N_26066,N_25869,N_25806);
xor U26067 (N_26067,N_25942,N_25886);
nand U26068 (N_26068,N_25873,N_25990);
xnor U26069 (N_26069,N_25883,N_25848);
xnor U26070 (N_26070,N_25917,N_25949);
nor U26071 (N_26071,N_25888,N_25908);
nor U26072 (N_26072,N_25985,N_25864);
nor U26073 (N_26073,N_25855,N_25902);
and U26074 (N_26074,N_25871,N_25939);
nor U26075 (N_26075,N_25828,N_25885);
and U26076 (N_26076,N_25850,N_25999);
nand U26077 (N_26077,N_25833,N_25992);
nor U26078 (N_26078,N_25893,N_25945);
nor U26079 (N_26079,N_25911,N_25811);
or U26080 (N_26080,N_25810,N_25994);
and U26081 (N_26081,N_25943,N_25997);
xor U26082 (N_26082,N_25831,N_25841);
nor U26083 (N_26083,N_25975,N_25969);
or U26084 (N_26084,N_25974,N_25986);
nand U26085 (N_26085,N_25853,N_25903);
and U26086 (N_26086,N_25921,N_25907);
or U26087 (N_26087,N_25826,N_25941);
xnor U26088 (N_26088,N_25910,N_25988);
nor U26089 (N_26089,N_25896,N_25973);
nor U26090 (N_26090,N_25809,N_25834);
nor U26091 (N_26091,N_25993,N_25825);
xor U26092 (N_26092,N_25996,N_25976);
nand U26093 (N_26093,N_25956,N_25815);
and U26094 (N_26094,N_25951,N_25891);
xor U26095 (N_26095,N_25944,N_25827);
or U26096 (N_26096,N_25938,N_25830);
or U26097 (N_26097,N_25979,N_25935);
nor U26098 (N_26098,N_25820,N_25856);
nor U26099 (N_26099,N_25998,N_25857);
nor U26100 (N_26100,N_25813,N_25821);
xor U26101 (N_26101,N_25836,N_25829);
and U26102 (N_26102,N_25855,N_25931);
xor U26103 (N_26103,N_25833,N_25861);
and U26104 (N_26104,N_25996,N_25835);
or U26105 (N_26105,N_25955,N_25895);
nand U26106 (N_26106,N_25931,N_25816);
and U26107 (N_26107,N_25830,N_25903);
nor U26108 (N_26108,N_25993,N_25976);
or U26109 (N_26109,N_25806,N_25819);
nand U26110 (N_26110,N_25838,N_25934);
and U26111 (N_26111,N_25821,N_25946);
nor U26112 (N_26112,N_25891,N_25853);
xnor U26113 (N_26113,N_25833,N_25954);
nor U26114 (N_26114,N_25831,N_25865);
nand U26115 (N_26115,N_25968,N_25942);
nand U26116 (N_26116,N_25808,N_25824);
and U26117 (N_26117,N_25980,N_25915);
or U26118 (N_26118,N_25876,N_25938);
nand U26119 (N_26119,N_25871,N_25961);
nor U26120 (N_26120,N_25875,N_25856);
xnor U26121 (N_26121,N_25898,N_25835);
xnor U26122 (N_26122,N_25816,N_25919);
and U26123 (N_26123,N_25804,N_25814);
and U26124 (N_26124,N_25922,N_25892);
nor U26125 (N_26125,N_25913,N_25816);
nor U26126 (N_26126,N_25992,N_25880);
or U26127 (N_26127,N_25909,N_25962);
and U26128 (N_26128,N_25836,N_25957);
nor U26129 (N_26129,N_25971,N_25903);
nand U26130 (N_26130,N_25821,N_25968);
nor U26131 (N_26131,N_25921,N_25835);
or U26132 (N_26132,N_25801,N_25943);
and U26133 (N_26133,N_25879,N_25989);
nand U26134 (N_26134,N_25880,N_25943);
xnor U26135 (N_26135,N_25811,N_25906);
xnor U26136 (N_26136,N_25987,N_25893);
xor U26137 (N_26137,N_25980,N_25845);
nand U26138 (N_26138,N_25875,N_25901);
xnor U26139 (N_26139,N_25806,N_25892);
xor U26140 (N_26140,N_25870,N_25917);
nor U26141 (N_26141,N_25968,N_25827);
and U26142 (N_26142,N_25930,N_25949);
and U26143 (N_26143,N_25826,N_25940);
and U26144 (N_26144,N_25897,N_25830);
nand U26145 (N_26145,N_25977,N_25911);
or U26146 (N_26146,N_25911,N_25854);
nand U26147 (N_26147,N_25822,N_25861);
nor U26148 (N_26148,N_25915,N_25849);
xnor U26149 (N_26149,N_25807,N_25946);
xnor U26150 (N_26150,N_25906,N_25943);
xnor U26151 (N_26151,N_25883,N_25857);
nand U26152 (N_26152,N_25892,N_25856);
nor U26153 (N_26153,N_25992,N_25839);
xnor U26154 (N_26154,N_25848,N_25929);
nor U26155 (N_26155,N_25948,N_25986);
nand U26156 (N_26156,N_25825,N_25850);
nor U26157 (N_26157,N_25891,N_25970);
and U26158 (N_26158,N_25993,N_25922);
xor U26159 (N_26159,N_25834,N_25880);
nand U26160 (N_26160,N_25991,N_25959);
nor U26161 (N_26161,N_25809,N_25940);
nand U26162 (N_26162,N_25804,N_25970);
or U26163 (N_26163,N_25867,N_25821);
xnor U26164 (N_26164,N_25874,N_25860);
xor U26165 (N_26165,N_25848,N_25935);
and U26166 (N_26166,N_25927,N_25999);
and U26167 (N_26167,N_25806,N_25939);
nor U26168 (N_26168,N_25991,N_25823);
nor U26169 (N_26169,N_25892,N_25938);
and U26170 (N_26170,N_25929,N_25936);
nor U26171 (N_26171,N_25860,N_25911);
or U26172 (N_26172,N_25843,N_25811);
nand U26173 (N_26173,N_25848,N_25855);
nor U26174 (N_26174,N_25805,N_25810);
nor U26175 (N_26175,N_25885,N_25892);
or U26176 (N_26176,N_25857,N_25814);
nand U26177 (N_26177,N_25803,N_25997);
nand U26178 (N_26178,N_25900,N_25885);
nand U26179 (N_26179,N_25969,N_25828);
xor U26180 (N_26180,N_25864,N_25993);
or U26181 (N_26181,N_25993,N_25915);
nor U26182 (N_26182,N_25935,N_25859);
nor U26183 (N_26183,N_25963,N_25875);
and U26184 (N_26184,N_25809,N_25913);
xor U26185 (N_26185,N_25968,N_25847);
nand U26186 (N_26186,N_25887,N_25996);
nand U26187 (N_26187,N_25815,N_25934);
xor U26188 (N_26188,N_25809,N_25819);
or U26189 (N_26189,N_25987,N_25863);
nand U26190 (N_26190,N_25987,N_25872);
xnor U26191 (N_26191,N_25882,N_25908);
or U26192 (N_26192,N_25971,N_25804);
nand U26193 (N_26193,N_25826,N_25946);
and U26194 (N_26194,N_25824,N_25839);
nor U26195 (N_26195,N_25853,N_25910);
or U26196 (N_26196,N_25854,N_25959);
and U26197 (N_26197,N_25998,N_25950);
nand U26198 (N_26198,N_25837,N_25845);
nor U26199 (N_26199,N_25899,N_25879);
xnor U26200 (N_26200,N_26149,N_26115);
nand U26201 (N_26201,N_26062,N_26137);
nor U26202 (N_26202,N_26043,N_26045);
or U26203 (N_26203,N_26056,N_26155);
nor U26204 (N_26204,N_26144,N_26022);
xor U26205 (N_26205,N_26180,N_26027);
nor U26206 (N_26206,N_26194,N_26175);
nor U26207 (N_26207,N_26130,N_26023);
xnor U26208 (N_26208,N_26141,N_26104);
xor U26209 (N_26209,N_26121,N_26158);
nor U26210 (N_26210,N_26112,N_26109);
nor U26211 (N_26211,N_26165,N_26148);
nor U26212 (N_26212,N_26168,N_26116);
xor U26213 (N_26213,N_26100,N_26196);
and U26214 (N_26214,N_26054,N_26038);
nor U26215 (N_26215,N_26024,N_26199);
nor U26216 (N_26216,N_26004,N_26019);
nand U26217 (N_26217,N_26110,N_26150);
or U26218 (N_26218,N_26037,N_26154);
or U26219 (N_26219,N_26173,N_26162);
nor U26220 (N_26220,N_26092,N_26189);
and U26221 (N_26221,N_26103,N_26005);
xnor U26222 (N_26222,N_26076,N_26167);
and U26223 (N_26223,N_26094,N_26108);
and U26224 (N_26224,N_26081,N_26088);
nor U26225 (N_26225,N_26051,N_26073);
or U26226 (N_26226,N_26114,N_26067);
and U26227 (N_26227,N_26035,N_26010);
nand U26228 (N_26228,N_26063,N_26174);
and U26229 (N_26229,N_26084,N_26143);
nor U26230 (N_26230,N_26039,N_26183);
xor U26231 (N_26231,N_26011,N_26044);
nand U26232 (N_26232,N_26036,N_26138);
and U26233 (N_26233,N_26060,N_26042);
and U26234 (N_26234,N_26185,N_26193);
or U26235 (N_26235,N_26075,N_26157);
nor U26236 (N_26236,N_26025,N_26098);
nor U26237 (N_26237,N_26192,N_26026);
and U26238 (N_26238,N_26096,N_26120);
nor U26239 (N_26239,N_26047,N_26034);
nor U26240 (N_26240,N_26018,N_26013);
nor U26241 (N_26241,N_26085,N_26184);
nand U26242 (N_26242,N_26017,N_26099);
or U26243 (N_26243,N_26049,N_26140);
nor U26244 (N_26244,N_26113,N_26055);
or U26245 (N_26245,N_26117,N_26122);
or U26246 (N_26246,N_26007,N_26052);
nor U26247 (N_26247,N_26050,N_26021);
nand U26248 (N_26248,N_26068,N_26132);
xnor U26249 (N_26249,N_26032,N_26124);
xor U26250 (N_26250,N_26146,N_26069);
or U26251 (N_26251,N_26064,N_26135);
or U26252 (N_26252,N_26028,N_26079);
and U26253 (N_26253,N_26111,N_26160);
and U26254 (N_26254,N_26082,N_26153);
nand U26255 (N_26255,N_26061,N_26077);
xnor U26256 (N_26256,N_26123,N_26078);
or U26257 (N_26257,N_26172,N_26169);
or U26258 (N_26258,N_26131,N_26093);
xor U26259 (N_26259,N_26182,N_26118);
and U26260 (N_26260,N_26046,N_26087);
nand U26261 (N_26261,N_26074,N_26101);
nor U26262 (N_26262,N_26127,N_26072);
and U26263 (N_26263,N_26102,N_26191);
nand U26264 (N_26264,N_26136,N_26156);
and U26265 (N_26265,N_26000,N_26164);
xor U26266 (N_26266,N_26033,N_26090);
xor U26267 (N_26267,N_26097,N_26057);
xor U26268 (N_26268,N_26197,N_26142);
nand U26269 (N_26269,N_26041,N_26170);
or U26270 (N_26270,N_26016,N_26048);
nand U26271 (N_26271,N_26133,N_26029);
and U26272 (N_26272,N_26188,N_26128);
xor U26273 (N_26273,N_26040,N_26001);
nand U26274 (N_26274,N_26195,N_26080);
and U26275 (N_26275,N_26031,N_26105);
xnor U26276 (N_26276,N_26106,N_26178);
xnor U26277 (N_26277,N_26186,N_26179);
xnor U26278 (N_26278,N_26014,N_26009);
and U26279 (N_26279,N_26152,N_26145);
nand U26280 (N_26280,N_26002,N_26166);
xnor U26281 (N_26281,N_26161,N_26012);
nand U26282 (N_26282,N_26003,N_26171);
nor U26283 (N_26283,N_26151,N_26058);
xor U26284 (N_26284,N_26176,N_26139);
and U26285 (N_26285,N_26190,N_26187);
and U26286 (N_26286,N_26066,N_26008);
and U26287 (N_26287,N_26030,N_26089);
nor U26288 (N_26288,N_26006,N_26059);
nand U26289 (N_26289,N_26159,N_26125);
or U26290 (N_26290,N_26053,N_26095);
xnor U26291 (N_26291,N_26065,N_26163);
and U26292 (N_26292,N_26091,N_26086);
xnor U26293 (N_26293,N_26119,N_26071);
and U26294 (N_26294,N_26015,N_26147);
or U26295 (N_26295,N_26129,N_26126);
xor U26296 (N_26296,N_26020,N_26070);
or U26297 (N_26297,N_26134,N_26177);
or U26298 (N_26298,N_26107,N_26181);
nor U26299 (N_26299,N_26198,N_26083);
or U26300 (N_26300,N_26197,N_26126);
and U26301 (N_26301,N_26106,N_26024);
and U26302 (N_26302,N_26000,N_26144);
and U26303 (N_26303,N_26176,N_26000);
nor U26304 (N_26304,N_26173,N_26075);
or U26305 (N_26305,N_26154,N_26152);
or U26306 (N_26306,N_26014,N_26063);
and U26307 (N_26307,N_26197,N_26168);
nand U26308 (N_26308,N_26101,N_26007);
xor U26309 (N_26309,N_26146,N_26111);
nand U26310 (N_26310,N_26139,N_26080);
nand U26311 (N_26311,N_26019,N_26184);
nand U26312 (N_26312,N_26136,N_26153);
xor U26313 (N_26313,N_26007,N_26126);
nand U26314 (N_26314,N_26169,N_26077);
and U26315 (N_26315,N_26185,N_26103);
and U26316 (N_26316,N_26043,N_26114);
xor U26317 (N_26317,N_26197,N_26146);
and U26318 (N_26318,N_26188,N_26160);
nand U26319 (N_26319,N_26036,N_26037);
nand U26320 (N_26320,N_26196,N_26148);
nor U26321 (N_26321,N_26115,N_26170);
and U26322 (N_26322,N_26196,N_26120);
nor U26323 (N_26323,N_26112,N_26164);
nand U26324 (N_26324,N_26138,N_26044);
xor U26325 (N_26325,N_26111,N_26051);
nor U26326 (N_26326,N_26087,N_26176);
or U26327 (N_26327,N_26166,N_26138);
and U26328 (N_26328,N_26010,N_26102);
and U26329 (N_26329,N_26057,N_26093);
or U26330 (N_26330,N_26029,N_26074);
nand U26331 (N_26331,N_26114,N_26153);
nand U26332 (N_26332,N_26188,N_26028);
and U26333 (N_26333,N_26109,N_26121);
xnor U26334 (N_26334,N_26102,N_26107);
or U26335 (N_26335,N_26135,N_26129);
xnor U26336 (N_26336,N_26164,N_26187);
or U26337 (N_26337,N_26113,N_26073);
and U26338 (N_26338,N_26127,N_26115);
xor U26339 (N_26339,N_26078,N_26015);
nand U26340 (N_26340,N_26152,N_26175);
and U26341 (N_26341,N_26136,N_26193);
nor U26342 (N_26342,N_26165,N_26154);
xor U26343 (N_26343,N_26078,N_26147);
or U26344 (N_26344,N_26074,N_26020);
nand U26345 (N_26345,N_26147,N_26154);
nand U26346 (N_26346,N_26019,N_26169);
and U26347 (N_26347,N_26132,N_26025);
nor U26348 (N_26348,N_26028,N_26124);
xor U26349 (N_26349,N_26163,N_26037);
and U26350 (N_26350,N_26106,N_26122);
or U26351 (N_26351,N_26134,N_26085);
xor U26352 (N_26352,N_26035,N_26081);
nor U26353 (N_26353,N_26009,N_26095);
and U26354 (N_26354,N_26055,N_26084);
nand U26355 (N_26355,N_26144,N_26173);
and U26356 (N_26356,N_26037,N_26142);
and U26357 (N_26357,N_26147,N_26040);
xor U26358 (N_26358,N_26134,N_26169);
and U26359 (N_26359,N_26016,N_26003);
nand U26360 (N_26360,N_26189,N_26008);
nor U26361 (N_26361,N_26198,N_26182);
xor U26362 (N_26362,N_26151,N_26066);
xor U26363 (N_26363,N_26061,N_26105);
nand U26364 (N_26364,N_26092,N_26035);
or U26365 (N_26365,N_26188,N_26078);
xor U26366 (N_26366,N_26156,N_26115);
and U26367 (N_26367,N_26182,N_26105);
or U26368 (N_26368,N_26138,N_26006);
or U26369 (N_26369,N_26078,N_26067);
and U26370 (N_26370,N_26179,N_26039);
and U26371 (N_26371,N_26112,N_26005);
nand U26372 (N_26372,N_26143,N_26164);
nor U26373 (N_26373,N_26146,N_26057);
xor U26374 (N_26374,N_26058,N_26148);
xor U26375 (N_26375,N_26126,N_26059);
nand U26376 (N_26376,N_26143,N_26137);
nand U26377 (N_26377,N_26013,N_26003);
and U26378 (N_26378,N_26020,N_26089);
and U26379 (N_26379,N_26036,N_26092);
xor U26380 (N_26380,N_26115,N_26066);
nand U26381 (N_26381,N_26172,N_26187);
nand U26382 (N_26382,N_26172,N_26055);
or U26383 (N_26383,N_26120,N_26080);
or U26384 (N_26384,N_26082,N_26056);
xor U26385 (N_26385,N_26190,N_26097);
nor U26386 (N_26386,N_26068,N_26080);
xnor U26387 (N_26387,N_26081,N_26109);
nand U26388 (N_26388,N_26197,N_26109);
and U26389 (N_26389,N_26174,N_26037);
and U26390 (N_26390,N_26077,N_26041);
nand U26391 (N_26391,N_26066,N_26095);
or U26392 (N_26392,N_26173,N_26083);
or U26393 (N_26393,N_26134,N_26120);
nor U26394 (N_26394,N_26173,N_26003);
and U26395 (N_26395,N_26101,N_26190);
xor U26396 (N_26396,N_26131,N_26129);
or U26397 (N_26397,N_26029,N_26062);
nand U26398 (N_26398,N_26180,N_26128);
and U26399 (N_26399,N_26185,N_26067);
nand U26400 (N_26400,N_26217,N_26355);
nand U26401 (N_26401,N_26232,N_26302);
xnor U26402 (N_26402,N_26312,N_26349);
nand U26403 (N_26403,N_26222,N_26397);
nor U26404 (N_26404,N_26354,N_26282);
and U26405 (N_26405,N_26248,N_26311);
and U26406 (N_26406,N_26239,N_26321);
and U26407 (N_26407,N_26359,N_26267);
nor U26408 (N_26408,N_26203,N_26269);
or U26409 (N_26409,N_26244,N_26398);
xor U26410 (N_26410,N_26357,N_26292);
xnor U26411 (N_26411,N_26376,N_26242);
nand U26412 (N_26412,N_26298,N_26364);
xnor U26413 (N_26413,N_26257,N_26393);
nand U26414 (N_26414,N_26206,N_26294);
and U26415 (N_26415,N_26253,N_26366);
nand U26416 (N_26416,N_26327,N_26211);
nand U26417 (N_26417,N_26291,N_26209);
nor U26418 (N_26418,N_26389,N_26307);
nor U26419 (N_26419,N_26338,N_26262);
nor U26420 (N_26420,N_26286,N_26263);
xnor U26421 (N_26421,N_26275,N_26391);
nor U26422 (N_26422,N_26337,N_26396);
or U26423 (N_26423,N_26216,N_26334);
xor U26424 (N_26424,N_26207,N_26394);
xnor U26425 (N_26425,N_26383,N_26308);
xnor U26426 (N_26426,N_26245,N_26296);
nor U26427 (N_26427,N_26270,N_26310);
nand U26428 (N_26428,N_26212,N_26363);
xor U26429 (N_26429,N_26230,N_26317);
nand U26430 (N_26430,N_26237,N_26299);
nor U26431 (N_26431,N_26300,N_26367);
xnor U26432 (N_26432,N_26247,N_26276);
xor U26433 (N_26433,N_26304,N_26289);
xnor U26434 (N_26434,N_26271,N_26339);
nor U26435 (N_26435,N_26335,N_26372);
nand U26436 (N_26436,N_26384,N_26382);
nand U26437 (N_26437,N_26274,N_26221);
and U26438 (N_26438,N_26325,N_26280);
xnor U26439 (N_26439,N_26219,N_26256);
or U26440 (N_26440,N_26214,N_26234);
xor U26441 (N_26441,N_26224,N_26255);
and U26442 (N_26442,N_26265,N_26264);
or U26443 (N_26443,N_26322,N_26208);
nand U26444 (N_26444,N_26392,N_26227);
nor U26445 (N_26445,N_26233,N_26251);
nor U26446 (N_26446,N_26202,N_26326);
or U26447 (N_26447,N_26301,N_26315);
nand U26448 (N_26448,N_26371,N_26240);
and U26449 (N_26449,N_26381,N_26358);
xnor U26450 (N_26450,N_26318,N_26368);
nand U26451 (N_26451,N_26385,N_26395);
xor U26452 (N_26452,N_26342,N_26279);
xnor U26453 (N_26453,N_26213,N_26215);
and U26454 (N_26454,N_26343,N_26336);
or U26455 (N_26455,N_26399,N_26313);
xor U26456 (N_26456,N_26204,N_26375);
xnor U26457 (N_26457,N_26223,N_26387);
and U26458 (N_26458,N_26236,N_26362);
nor U26459 (N_26459,N_26330,N_26243);
and U26460 (N_26460,N_26361,N_26356);
or U26461 (N_26461,N_26285,N_26306);
xnor U26462 (N_26462,N_26210,N_26254);
nand U26463 (N_26463,N_26273,N_26297);
nand U26464 (N_26464,N_26218,N_26379);
or U26465 (N_26465,N_26378,N_26370);
nor U26466 (N_26466,N_26231,N_26341);
nor U26467 (N_26467,N_26246,N_26250);
or U26468 (N_26468,N_26347,N_26319);
nor U26469 (N_26469,N_26277,N_26205);
and U26470 (N_26470,N_26220,N_26260);
and U26471 (N_26471,N_26373,N_26346);
xor U26472 (N_26472,N_26351,N_26200);
or U26473 (N_26473,N_26331,N_26281);
and U26474 (N_26474,N_26390,N_26241);
and U26475 (N_26475,N_26258,N_26348);
and U26476 (N_26476,N_26287,N_26314);
nor U26477 (N_26477,N_26226,N_26268);
xor U26478 (N_26478,N_26238,N_26259);
and U26479 (N_26479,N_26261,N_26228);
nand U26480 (N_26480,N_26303,N_26266);
nor U26481 (N_26481,N_26235,N_26295);
nor U26482 (N_26482,N_26388,N_26290);
nor U26483 (N_26483,N_26305,N_26345);
and U26484 (N_26484,N_26201,N_26332);
and U26485 (N_26485,N_26320,N_26278);
xnor U26486 (N_26486,N_26340,N_26350);
nand U26487 (N_26487,N_26386,N_26249);
nor U26488 (N_26488,N_26365,N_26374);
nor U26489 (N_26489,N_26283,N_26369);
nand U26490 (N_26490,N_26252,N_26360);
xnor U26491 (N_26491,N_26272,N_26380);
nor U26492 (N_26492,N_26344,N_26352);
nand U26493 (N_26493,N_26324,N_26225);
nand U26494 (N_26494,N_26333,N_26329);
nor U26495 (N_26495,N_26316,N_26353);
xor U26496 (N_26496,N_26284,N_26328);
xor U26497 (N_26497,N_26377,N_26229);
xnor U26498 (N_26498,N_26323,N_26309);
or U26499 (N_26499,N_26293,N_26288);
nor U26500 (N_26500,N_26327,N_26317);
nand U26501 (N_26501,N_26216,N_26304);
nor U26502 (N_26502,N_26361,N_26287);
xor U26503 (N_26503,N_26236,N_26234);
xnor U26504 (N_26504,N_26379,N_26226);
xnor U26505 (N_26505,N_26210,N_26286);
or U26506 (N_26506,N_26239,N_26214);
or U26507 (N_26507,N_26205,N_26390);
nor U26508 (N_26508,N_26234,N_26258);
xor U26509 (N_26509,N_26308,N_26222);
xor U26510 (N_26510,N_26233,N_26219);
or U26511 (N_26511,N_26216,N_26298);
or U26512 (N_26512,N_26352,N_26388);
or U26513 (N_26513,N_26243,N_26278);
or U26514 (N_26514,N_26320,N_26295);
and U26515 (N_26515,N_26303,N_26201);
nand U26516 (N_26516,N_26393,N_26286);
and U26517 (N_26517,N_26213,N_26201);
nand U26518 (N_26518,N_26215,N_26241);
and U26519 (N_26519,N_26369,N_26294);
or U26520 (N_26520,N_26286,N_26302);
xor U26521 (N_26521,N_26244,N_26209);
or U26522 (N_26522,N_26272,N_26257);
xnor U26523 (N_26523,N_26241,N_26282);
or U26524 (N_26524,N_26380,N_26276);
nor U26525 (N_26525,N_26380,N_26257);
xor U26526 (N_26526,N_26254,N_26286);
and U26527 (N_26527,N_26228,N_26306);
nor U26528 (N_26528,N_26342,N_26212);
nand U26529 (N_26529,N_26295,N_26357);
xor U26530 (N_26530,N_26249,N_26310);
nand U26531 (N_26531,N_26322,N_26350);
or U26532 (N_26532,N_26370,N_26385);
nor U26533 (N_26533,N_26360,N_26366);
or U26534 (N_26534,N_26226,N_26292);
xor U26535 (N_26535,N_26308,N_26377);
and U26536 (N_26536,N_26273,N_26256);
and U26537 (N_26537,N_26347,N_26361);
nand U26538 (N_26538,N_26218,N_26262);
and U26539 (N_26539,N_26200,N_26327);
nand U26540 (N_26540,N_26224,N_26315);
nand U26541 (N_26541,N_26251,N_26243);
nand U26542 (N_26542,N_26272,N_26360);
and U26543 (N_26543,N_26245,N_26226);
nor U26544 (N_26544,N_26287,N_26261);
nor U26545 (N_26545,N_26312,N_26300);
nor U26546 (N_26546,N_26215,N_26340);
xnor U26547 (N_26547,N_26357,N_26283);
xnor U26548 (N_26548,N_26260,N_26399);
nor U26549 (N_26549,N_26224,N_26300);
nand U26550 (N_26550,N_26345,N_26223);
or U26551 (N_26551,N_26374,N_26241);
nor U26552 (N_26552,N_26224,N_26369);
nor U26553 (N_26553,N_26264,N_26209);
nand U26554 (N_26554,N_26332,N_26316);
nand U26555 (N_26555,N_26397,N_26240);
or U26556 (N_26556,N_26292,N_26297);
nand U26557 (N_26557,N_26243,N_26221);
and U26558 (N_26558,N_26330,N_26209);
or U26559 (N_26559,N_26268,N_26327);
nand U26560 (N_26560,N_26207,N_26246);
nand U26561 (N_26561,N_26263,N_26291);
and U26562 (N_26562,N_26361,N_26271);
xor U26563 (N_26563,N_26204,N_26352);
and U26564 (N_26564,N_26319,N_26277);
xnor U26565 (N_26565,N_26355,N_26240);
xnor U26566 (N_26566,N_26393,N_26224);
nor U26567 (N_26567,N_26215,N_26308);
nand U26568 (N_26568,N_26239,N_26262);
and U26569 (N_26569,N_26387,N_26282);
and U26570 (N_26570,N_26397,N_26364);
or U26571 (N_26571,N_26330,N_26381);
nor U26572 (N_26572,N_26301,N_26209);
xor U26573 (N_26573,N_26361,N_26329);
or U26574 (N_26574,N_26253,N_26227);
nor U26575 (N_26575,N_26361,N_26276);
and U26576 (N_26576,N_26262,N_26226);
nor U26577 (N_26577,N_26377,N_26231);
nand U26578 (N_26578,N_26331,N_26354);
nor U26579 (N_26579,N_26377,N_26297);
nand U26580 (N_26580,N_26348,N_26294);
nor U26581 (N_26581,N_26365,N_26384);
nand U26582 (N_26582,N_26230,N_26209);
and U26583 (N_26583,N_26303,N_26252);
and U26584 (N_26584,N_26367,N_26385);
or U26585 (N_26585,N_26329,N_26284);
or U26586 (N_26586,N_26312,N_26329);
and U26587 (N_26587,N_26399,N_26220);
or U26588 (N_26588,N_26275,N_26286);
and U26589 (N_26589,N_26355,N_26278);
nor U26590 (N_26590,N_26353,N_26380);
xor U26591 (N_26591,N_26390,N_26279);
nand U26592 (N_26592,N_26257,N_26309);
nor U26593 (N_26593,N_26201,N_26355);
and U26594 (N_26594,N_26388,N_26391);
nor U26595 (N_26595,N_26315,N_26247);
nor U26596 (N_26596,N_26304,N_26342);
or U26597 (N_26597,N_26348,N_26227);
nor U26598 (N_26598,N_26216,N_26253);
or U26599 (N_26599,N_26399,N_26283);
xor U26600 (N_26600,N_26492,N_26448);
nand U26601 (N_26601,N_26541,N_26575);
or U26602 (N_26602,N_26480,N_26520);
or U26603 (N_26603,N_26514,N_26435);
nor U26604 (N_26604,N_26451,N_26439);
or U26605 (N_26605,N_26573,N_26401);
or U26606 (N_26606,N_26499,N_26483);
nor U26607 (N_26607,N_26489,N_26449);
or U26608 (N_26608,N_26568,N_26402);
nor U26609 (N_26609,N_26570,N_26505);
xor U26610 (N_26610,N_26522,N_26513);
nor U26611 (N_26611,N_26488,N_26486);
and U26612 (N_26612,N_26478,N_26438);
nand U26613 (N_26613,N_26546,N_26458);
and U26614 (N_26614,N_26584,N_26574);
nor U26615 (N_26615,N_26554,N_26555);
nor U26616 (N_26616,N_26443,N_26504);
or U26617 (N_26617,N_26450,N_26490);
nor U26618 (N_26618,N_26571,N_26440);
and U26619 (N_26619,N_26510,N_26566);
nand U26620 (N_26620,N_26589,N_26547);
xnor U26621 (N_26621,N_26576,N_26494);
xor U26622 (N_26622,N_26412,N_26549);
nand U26623 (N_26623,N_26519,N_26508);
xor U26624 (N_26624,N_26423,N_26561);
nor U26625 (N_26625,N_26521,N_26594);
or U26626 (N_26626,N_26543,N_26456);
and U26627 (N_26627,N_26477,N_26411);
nor U26628 (N_26628,N_26461,N_26422);
nor U26629 (N_26629,N_26523,N_26471);
and U26630 (N_26630,N_26597,N_26403);
and U26631 (N_26631,N_26415,N_26537);
or U26632 (N_26632,N_26410,N_26503);
and U26633 (N_26633,N_26468,N_26563);
xnor U26634 (N_26634,N_26536,N_26445);
and U26635 (N_26635,N_26446,N_26473);
xnor U26636 (N_26636,N_26479,N_26587);
or U26637 (N_26637,N_26538,N_26404);
nor U26638 (N_26638,N_26407,N_26591);
or U26639 (N_26639,N_26557,N_26515);
and U26640 (N_26640,N_26484,N_26509);
nand U26641 (N_26641,N_26592,N_26485);
nor U26642 (N_26642,N_26436,N_26562);
nand U26643 (N_26643,N_26432,N_26596);
nand U26644 (N_26644,N_26497,N_26418);
xor U26645 (N_26645,N_26464,N_26463);
xnor U26646 (N_26646,N_26482,N_26586);
or U26647 (N_26647,N_26569,N_26465);
or U26648 (N_26648,N_26400,N_26472);
xnor U26649 (N_26649,N_26481,N_26512);
nor U26650 (N_26650,N_26579,N_26559);
and U26651 (N_26651,N_26491,N_26487);
and U26652 (N_26652,N_26518,N_26454);
nand U26653 (N_26653,N_26437,N_26409);
and U26654 (N_26654,N_26558,N_26539);
xor U26655 (N_26655,N_26553,N_26413);
or U26656 (N_26656,N_26556,N_26531);
and U26657 (N_26657,N_26598,N_26564);
nand U26658 (N_26658,N_26419,N_26476);
nor U26659 (N_26659,N_26593,N_26590);
or U26660 (N_26660,N_26421,N_26453);
or U26661 (N_26661,N_26517,N_26493);
or U26662 (N_26662,N_26572,N_26431);
or U26663 (N_26663,N_26424,N_26599);
and U26664 (N_26664,N_26567,N_26447);
and U26665 (N_26665,N_26474,N_26434);
nand U26666 (N_26666,N_26527,N_26416);
or U26667 (N_26667,N_26583,N_26582);
xnor U26668 (N_26668,N_26548,N_26414);
xor U26669 (N_26669,N_26469,N_26578);
xnor U26670 (N_26670,N_26550,N_26429);
xnor U26671 (N_26671,N_26405,N_26506);
and U26672 (N_26672,N_26552,N_26560);
xor U26673 (N_26673,N_26495,N_26501);
nand U26674 (N_26674,N_26580,N_26444);
nor U26675 (N_26675,N_26430,N_26475);
and U26676 (N_26676,N_26595,N_26542);
or U26677 (N_26677,N_26585,N_26500);
or U26678 (N_26678,N_26565,N_26530);
xor U26679 (N_26679,N_26452,N_26540);
and U26680 (N_26680,N_26545,N_26426);
xnor U26681 (N_26681,N_26525,N_26544);
nor U26682 (N_26682,N_26455,N_26526);
xor U26683 (N_26683,N_26459,N_26462);
or U26684 (N_26684,N_26408,N_26460);
and U26685 (N_26685,N_26441,N_26466);
xnor U26686 (N_26686,N_26507,N_26502);
nor U26687 (N_26687,N_26524,N_26420);
nor U26688 (N_26688,N_26535,N_26551);
nor U26689 (N_26689,N_26467,N_26533);
nand U26690 (N_26690,N_26534,N_26511);
nand U26691 (N_26691,N_26496,N_26529);
nor U26692 (N_26692,N_26427,N_26577);
nor U26693 (N_26693,N_26588,N_26442);
or U26694 (N_26694,N_26406,N_26428);
nand U26695 (N_26695,N_26433,N_26417);
or U26696 (N_26696,N_26470,N_26581);
and U26697 (N_26697,N_26498,N_26516);
or U26698 (N_26698,N_26532,N_26528);
nor U26699 (N_26699,N_26425,N_26457);
xnor U26700 (N_26700,N_26579,N_26539);
or U26701 (N_26701,N_26502,N_26559);
nor U26702 (N_26702,N_26577,N_26595);
nor U26703 (N_26703,N_26559,N_26516);
nand U26704 (N_26704,N_26592,N_26459);
nor U26705 (N_26705,N_26408,N_26598);
or U26706 (N_26706,N_26470,N_26449);
or U26707 (N_26707,N_26468,N_26488);
or U26708 (N_26708,N_26586,N_26556);
nand U26709 (N_26709,N_26533,N_26422);
nor U26710 (N_26710,N_26528,N_26586);
nand U26711 (N_26711,N_26509,N_26457);
or U26712 (N_26712,N_26440,N_26426);
nand U26713 (N_26713,N_26491,N_26596);
nor U26714 (N_26714,N_26455,N_26572);
xnor U26715 (N_26715,N_26407,N_26568);
and U26716 (N_26716,N_26582,N_26576);
and U26717 (N_26717,N_26408,N_26441);
or U26718 (N_26718,N_26496,N_26415);
or U26719 (N_26719,N_26501,N_26527);
and U26720 (N_26720,N_26592,N_26444);
nor U26721 (N_26721,N_26547,N_26525);
nand U26722 (N_26722,N_26556,N_26456);
or U26723 (N_26723,N_26567,N_26575);
xnor U26724 (N_26724,N_26591,N_26440);
and U26725 (N_26725,N_26550,N_26424);
or U26726 (N_26726,N_26462,N_26427);
nor U26727 (N_26727,N_26552,N_26547);
or U26728 (N_26728,N_26593,N_26478);
nor U26729 (N_26729,N_26532,N_26402);
or U26730 (N_26730,N_26473,N_26579);
and U26731 (N_26731,N_26420,N_26523);
xor U26732 (N_26732,N_26584,N_26465);
xnor U26733 (N_26733,N_26568,N_26566);
nand U26734 (N_26734,N_26484,N_26401);
and U26735 (N_26735,N_26499,N_26575);
nand U26736 (N_26736,N_26554,N_26580);
or U26737 (N_26737,N_26507,N_26446);
or U26738 (N_26738,N_26570,N_26485);
and U26739 (N_26739,N_26412,N_26417);
nand U26740 (N_26740,N_26426,N_26528);
xnor U26741 (N_26741,N_26446,N_26575);
nor U26742 (N_26742,N_26589,N_26437);
or U26743 (N_26743,N_26504,N_26535);
nand U26744 (N_26744,N_26418,N_26505);
or U26745 (N_26745,N_26433,N_26429);
nand U26746 (N_26746,N_26482,N_26552);
or U26747 (N_26747,N_26403,N_26569);
nand U26748 (N_26748,N_26527,N_26405);
nand U26749 (N_26749,N_26550,N_26449);
nand U26750 (N_26750,N_26539,N_26540);
nor U26751 (N_26751,N_26456,N_26538);
and U26752 (N_26752,N_26541,N_26594);
or U26753 (N_26753,N_26473,N_26451);
xnor U26754 (N_26754,N_26561,N_26557);
nand U26755 (N_26755,N_26598,N_26484);
and U26756 (N_26756,N_26487,N_26459);
nand U26757 (N_26757,N_26447,N_26475);
nand U26758 (N_26758,N_26425,N_26462);
nor U26759 (N_26759,N_26591,N_26495);
xor U26760 (N_26760,N_26486,N_26579);
nor U26761 (N_26761,N_26539,N_26473);
nor U26762 (N_26762,N_26569,N_26466);
xnor U26763 (N_26763,N_26401,N_26445);
xor U26764 (N_26764,N_26404,N_26524);
nand U26765 (N_26765,N_26490,N_26557);
nand U26766 (N_26766,N_26503,N_26464);
and U26767 (N_26767,N_26525,N_26521);
nand U26768 (N_26768,N_26505,N_26536);
nand U26769 (N_26769,N_26480,N_26423);
nor U26770 (N_26770,N_26581,N_26525);
xor U26771 (N_26771,N_26432,N_26533);
and U26772 (N_26772,N_26457,N_26599);
nand U26773 (N_26773,N_26495,N_26404);
and U26774 (N_26774,N_26467,N_26534);
nor U26775 (N_26775,N_26577,N_26457);
xor U26776 (N_26776,N_26438,N_26512);
or U26777 (N_26777,N_26569,N_26578);
nand U26778 (N_26778,N_26408,N_26462);
or U26779 (N_26779,N_26532,N_26533);
and U26780 (N_26780,N_26400,N_26467);
nand U26781 (N_26781,N_26473,N_26570);
nand U26782 (N_26782,N_26518,N_26509);
nor U26783 (N_26783,N_26496,N_26476);
or U26784 (N_26784,N_26593,N_26463);
xnor U26785 (N_26785,N_26503,N_26434);
or U26786 (N_26786,N_26467,N_26440);
and U26787 (N_26787,N_26418,N_26553);
nor U26788 (N_26788,N_26571,N_26531);
and U26789 (N_26789,N_26566,N_26458);
and U26790 (N_26790,N_26513,N_26409);
or U26791 (N_26791,N_26539,N_26436);
or U26792 (N_26792,N_26579,N_26571);
nor U26793 (N_26793,N_26460,N_26472);
or U26794 (N_26794,N_26423,N_26481);
xor U26795 (N_26795,N_26537,N_26571);
and U26796 (N_26796,N_26506,N_26514);
xor U26797 (N_26797,N_26534,N_26589);
xnor U26798 (N_26798,N_26454,N_26596);
or U26799 (N_26799,N_26476,N_26447);
xor U26800 (N_26800,N_26652,N_26760);
xor U26801 (N_26801,N_26762,N_26729);
and U26802 (N_26802,N_26797,N_26753);
nor U26803 (N_26803,N_26684,N_26693);
or U26804 (N_26804,N_26763,N_26791);
and U26805 (N_26805,N_26719,N_26728);
or U26806 (N_26806,N_26758,N_26750);
xnor U26807 (N_26807,N_26646,N_26783);
xnor U26808 (N_26808,N_26650,N_26632);
and U26809 (N_26809,N_26657,N_26681);
xor U26810 (N_26810,N_26606,N_26616);
or U26811 (N_26811,N_26672,N_26639);
nand U26812 (N_26812,N_26615,N_26757);
nand U26813 (N_26813,N_26779,N_26781);
and U26814 (N_26814,N_26723,N_26691);
xor U26815 (N_26815,N_26756,N_26747);
nand U26816 (N_26816,N_26739,N_26673);
nand U26817 (N_26817,N_26700,N_26789);
nor U26818 (N_26818,N_26622,N_26734);
xor U26819 (N_26819,N_26609,N_26655);
nand U26820 (N_26820,N_26707,N_26787);
xnor U26821 (N_26821,N_26661,N_26746);
and U26822 (N_26822,N_26735,N_26687);
xnor U26823 (N_26823,N_26648,N_26620);
nor U26824 (N_26824,N_26663,N_26738);
and U26825 (N_26825,N_26699,N_26714);
nand U26826 (N_26826,N_26614,N_26640);
nand U26827 (N_26827,N_26610,N_26694);
nand U26828 (N_26828,N_26647,N_26752);
xnor U26829 (N_26829,N_26755,N_26773);
and U26830 (N_26830,N_26618,N_26623);
nor U26831 (N_26831,N_26630,N_26769);
nand U26832 (N_26832,N_26730,N_26701);
xor U26833 (N_26833,N_26712,N_26659);
nor U26834 (N_26834,N_26705,N_26709);
xnor U26835 (N_26835,N_26676,N_26733);
or U26836 (N_26836,N_26764,N_26642);
and U26837 (N_26837,N_26748,N_26794);
or U26838 (N_26838,N_26708,N_26774);
and U26839 (N_26839,N_26771,N_26754);
or U26840 (N_26840,N_26625,N_26782);
nand U26841 (N_26841,N_26702,N_26660);
xor U26842 (N_26842,N_26703,N_26795);
nor U26843 (N_26843,N_26751,N_26766);
nand U26844 (N_26844,N_26613,N_26720);
xor U26845 (N_26845,N_26643,N_26692);
and U26846 (N_26846,N_26670,N_26780);
nor U26847 (N_26847,N_26724,N_26679);
or U26848 (N_26848,N_26674,N_26690);
xnor U26849 (N_26849,N_26678,N_26772);
nor U26850 (N_26850,N_26710,N_26775);
nor U26851 (N_26851,N_26665,N_26799);
xnor U26852 (N_26852,N_26677,N_26631);
and U26853 (N_26853,N_26745,N_26669);
nand U26854 (N_26854,N_26658,N_26731);
and U26855 (N_26855,N_26635,N_26706);
and U26856 (N_26856,N_26759,N_26718);
or U26857 (N_26857,N_26628,N_26736);
nor U26858 (N_26858,N_26770,N_26629);
nor U26859 (N_26859,N_26798,N_26689);
nor U26860 (N_26860,N_26634,N_26742);
or U26861 (N_26861,N_26641,N_26737);
nand U26862 (N_26862,N_26698,N_26656);
and U26863 (N_26863,N_26727,N_26683);
or U26864 (N_26864,N_26790,N_26685);
nand U26865 (N_26865,N_26675,N_26711);
or U26866 (N_26866,N_26668,N_26717);
and U26867 (N_26867,N_26666,N_26627);
nand U26868 (N_26868,N_26626,N_26662);
or U26869 (N_26869,N_26722,N_26637);
xor U26870 (N_26870,N_26778,N_26654);
nor U26871 (N_26871,N_26645,N_26761);
nor U26872 (N_26872,N_26741,N_26644);
or U26873 (N_26873,N_26768,N_26664);
and U26874 (N_26874,N_26686,N_26776);
and U26875 (N_26875,N_26633,N_26765);
and U26876 (N_26876,N_26788,N_26786);
nor U26877 (N_26877,N_26695,N_26680);
nor U26878 (N_26878,N_26621,N_26697);
or U26879 (N_26879,N_26604,N_26653);
xnor U26880 (N_26880,N_26721,N_26732);
nand U26881 (N_26881,N_26716,N_26671);
nand U26882 (N_26882,N_26744,N_26793);
nand U26883 (N_26883,N_26636,N_26651);
nand U26884 (N_26884,N_26605,N_26600);
or U26885 (N_26885,N_26624,N_26767);
nand U26886 (N_26886,N_26696,N_26784);
and U26887 (N_26887,N_26792,N_26785);
nand U26888 (N_26888,N_26612,N_26638);
and U26889 (N_26889,N_26607,N_26796);
or U26890 (N_26890,N_26601,N_26602);
nor U26891 (N_26891,N_26617,N_26608);
or U26892 (N_26892,N_26725,N_26743);
and U26893 (N_26893,N_26740,N_26688);
xor U26894 (N_26894,N_26667,N_26715);
and U26895 (N_26895,N_26619,N_26611);
nor U26896 (N_26896,N_26603,N_26726);
and U26897 (N_26897,N_26682,N_26713);
xor U26898 (N_26898,N_26777,N_26749);
nor U26899 (N_26899,N_26704,N_26649);
and U26900 (N_26900,N_26788,N_26621);
xor U26901 (N_26901,N_26725,N_26739);
xor U26902 (N_26902,N_26618,N_26770);
and U26903 (N_26903,N_26681,N_26680);
nor U26904 (N_26904,N_26711,N_26761);
nand U26905 (N_26905,N_26646,N_26716);
nand U26906 (N_26906,N_26742,N_26681);
or U26907 (N_26907,N_26604,N_26691);
xnor U26908 (N_26908,N_26780,N_26682);
or U26909 (N_26909,N_26741,N_26790);
xor U26910 (N_26910,N_26625,N_26760);
xor U26911 (N_26911,N_26764,N_26638);
or U26912 (N_26912,N_26695,N_26765);
or U26913 (N_26913,N_26706,N_26703);
and U26914 (N_26914,N_26674,N_26773);
nand U26915 (N_26915,N_26720,N_26705);
or U26916 (N_26916,N_26751,N_26765);
and U26917 (N_26917,N_26676,N_26716);
nor U26918 (N_26918,N_26733,N_26777);
xnor U26919 (N_26919,N_26625,N_26729);
xnor U26920 (N_26920,N_26760,N_26758);
xor U26921 (N_26921,N_26667,N_26635);
and U26922 (N_26922,N_26753,N_26689);
nand U26923 (N_26923,N_26670,N_26731);
or U26924 (N_26924,N_26644,N_26606);
or U26925 (N_26925,N_26760,N_26666);
or U26926 (N_26926,N_26605,N_26610);
or U26927 (N_26927,N_26793,N_26748);
nor U26928 (N_26928,N_26792,N_26748);
nand U26929 (N_26929,N_26606,N_26717);
and U26930 (N_26930,N_26789,N_26603);
xor U26931 (N_26931,N_26633,N_26716);
and U26932 (N_26932,N_26685,N_26713);
and U26933 (N_26933,N_26707,N_26600);
or U26934 (N_26934,N_26670,N_26616);
and U26935 (N_26935,N_26751,N_26767);
and U26936 (N_26936,N_26791,N_26698);
or U26937 (N_26937,N_26676,N_26728);
nor U26938 (N_26938,N_26675,N_26780);
and U26939 (N_26939,N_26735,N_26700);
nor U26940 (N_26940,N_26789,N_26691);
and U26941 (N_26941,N_26722,N_26604);
nand U26942 (N_26942,N_26700,N_26681);
xor U26943 (N_26943,N_26755,N_26767);
xnor U26944 (N_26944,N_26683,N_26789);
nor U26945 (N_26945,N_26644,N_26667);
xor U26946 (N_26946,N_26757,N_26734);
and U26947 (N_26947,N_26621,N_26762);
nor U26948 (N_26948,N_26653,N_26663);
nand U26949 (N_26949,N_26717,N_26635);
nand U26950 (N_26950,N_26657,N_26638);
or U26951 (N_26951,N_26604,N_26680);
nor U26952 (N_26952,N_26790,N_26773);
nor U26953 (N_26953,N_26793,N_26674);
and U26954 (N_26954,N_26722,N_26606);
nor U26955 (N_26955,N_26712,N_26795);
nand U26956 (N_26956,N_26630,N_26693);
xnor U26957 (N_26957,N_26734,N_26661);
xor U26958 (N_26958,N_26768,N_26663);
or U26959 (N_26959,N_26609,N_26671);
nor U26960 (N_26960,N_26771,N_26615);
nand U26961 (N_26961,N_26752,N_26608);
nand U26962 (N_26962,N_26745,N_26657);
or U26963 (N_26963,N_26638,N_26737);
nand U26964 (N_26964,N_26682,N_26665);
and U26965 (N_26965,N_26742,N_26635);
nor U26966 (N_26966,N_26733,N_26653);
nor U26967 (N_26967,N_26649,N_26791);
and U26968 (N_26968,N_26740,N_26787);
nand U26969 (N_26969,N_26606,N_26690);
nand U26970 (N_26970,N_26707,N_26626);
and U26971 (N_26971,N_26617,N_26720);
and U26972 (N_26972,N_26692,N_26689);
nand U26973 (N_26973,N_26782,N_26669);
nor U26974 (N_26974,N_26613,N_26774);
or U26975 (N_26975,N_26736,N_26677);
and U26976 (N_26976,N_26624,N_26739);
xnor U26977 (N_26977,N_26770,N_26603);
nor U26978 (N_26978,N_26654,N_26756);
nand U26979 (N_26979,N_26775,N_26771);
nand U26980 (N_26980,N_26747,N_26769);
xor U26981 (N_26981,N_26720,N_26767);
and U26982 (N_26982,N_26716,N_26710);
nor U26983 (N_26983,N_26773,N_26710);
nand U26984 (N_26984,N_26683,N_26618);
nand U26985 (N_26985,N_26615,N_26728);
nor U26986 (N_26986,N_26678,N_26665);
or U26987 (N_26987,N_26755,N_26690);
nand U26988 (N_26988,N_26625,N_26607);
nor U26989 (N_26989,N_26627,N_26714);
nor U26990 (N_26990,N_26727,N_26619);
nor U26991 (N_26991,N_26655,N_26716);
or U26992 (N_26992,N_26641,N_26728);
nand U26993 (N_26993,N_26633,N_26604);
nor U26994 (N_26994,N_26644,N_26611);
xnor U26995 (N_26995,N_26729,N_26794);
and U26996 (N_26996,N_26640,N_26667);
xor U26997 (N_26997,N_26627,N_26665);
nor U26998 (N_26998,N_26689,N_26629);
and U26999 (N_26999,N_26749,N_26769);
and U27000 (N_27000,N_26960,N_26876);
and U27001 (N_27001,N_26807,N_26889);
or U27002 (N_27002,N_26852,N_26821);
nor U27003 (N_27003,N_26816,N_26813);
nand U27004 (N_27004,N_26869,N_26820);
and U27005 (N_27005,N_26881,N_26861);
nand U27006 (N_27006,N_26837,N_26958);
nor U27007 (N_27007,N_26956,N_26809);
nand U27008 (N_27008,N_26953,N_26819);
nand U27009 (N_27009,N_26959,N_26843);
nor U27010 (N_27010,N_26871,N_26911);
and U27011 (N_27011,N_26831,N_26933);
nand U27012 (N_27012,N_26965,N_26914);
nor U27013 (N_27013,N_26894,N_26985);
xnor U27014 (N_27014,N_26921,N_26896);
and U27015 (N_27015,N_26815,N_26980);
xnor U27016 (N_27016,N_26878,N_26873);
and U27017 (N_27017,N_26903,N_26833);
nor U27018 (N_27018,N_26810,N_26818);
and U27019 (N_27019,N_26939,N_26936);
nand U27020 (N_27020,N_26899,N_26991);
or U27021 (N_27021,N_26966,N_26859);
xor U27022 (N_27022,N_26835,N_26864);
nor U27023 (N_27023,N_26986,N_26988);
or U27024 (N_27024,N_26895,N_26845);
nor U27025 (N_27025,N_26941,N_26997);
or U27026 (N_27026,N_26972,N_26981);
and U27027 (N_27027,N_26967,N_26901);
xor U27028 (N_27028,N_26961,N_26890);
nor U27029 (N_27029,N_26848,N_26908);
and U27030 (N_27030,N_26826,N_26806);
or U27031 (N_27031,N_26946,N_26948);
nand U27032 (N_27032,N_26917,N_26934);
and U27033 (N_27033,N_26858,N_26817);
or U27034 (N_27034,N_26919,N_26857);
xor U27035 (N_27035,N_26930,N_26954);
and U27036 (N_27036,N_26925,N_26916);
xor U27037 (N_27037,N_26990,N_26907);
nor U27038 (N_27038,N_26900,N_26830);
or U27039 (N_27039,N_26964,N_26824);
nand U27040 (N_27040,N_26846,N_26885);
nand U27041 (N_27041,N_26913,N_26850);
and U27042 (N_27042,N_26855,N_26923);
and U27043 (N_27043,N_26841,N_26992);
or U27044 (N_27044,N_26849,N_26942);
xor U27045 (N_27045,N_26893,N_26839);
or U27046 (N_27046,N_26822,N_26897);
xor U27047 (N_27047,N_26909,N_26867);
and U27048 (N_27048,N_26996,N_26874);
or U27049 (N_27049,N_26832,N_26882);
nand U27050 (N_27050,N_26993,N_26928);
or U27051 (N_27051,N_26863,N_26898);
nand U27052 (N_27052,N_26971,N_26834);
or U27053 (N_27053,N_26978,N_26929);
nor U27054 (N_27054,N_26987,N_26968);
nor U27055 (N_27055,N_26853,N_26924);
or U27056 (N_27056,N_26805,N_26982);
nand U27057 (N_27057,N_26868,N_26957);
and U27058 (N_27058,N_26998,N_26840);
nand U27059 (N_27059,N_26935,N_26989);
nor U27060 (N_27060,N_26938,N_26870);
nor U27061 (N_27061,N_26825,N_26962);
xnor U27062 (N_27062,N_26943,N_26844);
nand U27063 (N_27063,N_26951,N_26827);
nand U27064 (N_27064,N_26836,N_26976);
or U27065 (N_27065,N_26927,N_26872);
or U27066 (N_27066,N_26904,N_26866);
and U27067 (N_27067,N_26802,N_26950);
and U27068 (N_27068,N_26801,N_26888);
and U27069 (N_27069,N_26949,N_26877);
xnor U27070 (N_27070,N_26812,N_26884);
nor U27071 (N_27071,N_26995,N_26983);
or U27072 (N_27072,N_26979,N_26906);
or U27073 (N_27073,N_26838,N_26926);
nor U27074 (N_27074,N_26918,N_26800);
or U27075 (N_27075,N_26880,N_26851);
and U27076 (N_27076,N_26940,N_26811);
or U27077 (N_27077,N_26974,N_26883);
or U27078 (N_27078,N_26931,N_26905);
nand U27079 (N_27079,N_26975,N_26944);
or U27080 (N_27080,N_26860,N_26984);
nor U27081 (N_27081,N_26970,N_26847);
nor U27082 (N_27082,N_26823,N_26842);
nor U27083 (N_27083,N_26973,N_26945);
nand U27084 (N_27084,N_26994,N_26891);
nand U27085 (N_27085,N_26977,N_26910);
xnor U27086 (N_27086,N_26912,N_26922);
and U27087 (N_27087,N_26999,N_26932);
or U27088 (N_27088,N_26915,N_26963);
or U27089 (N_27089,N_26879,N_26902);
nor U27090 (N_27090,N_26804,N_26886);
and U27091 (N_27091,N_26969,N_26887);
xor U27092 (N_27092,N_26828,N_26808);
nand U27093 (N_27093,N_26892,N_26952);
nor U27094 (N_27094,N_26875,N_26947);
nor U27095 (N_27095,N_26814,N_26829);
nor U27096 (N_27096,N_26862,N_26937);
xor U27097 (N_27097,N_26865,N_26955);
nand U27098 (N_27098,N_26854,N_26856);
and U27099 (N_27099,N_26920,N_26803);
nand U27100 (N_27100,N_26930,N_26800);
and U27101 (N_27101,N_26907,N_26949);
nand U27102 (N_27102,N_26964,N_26830);
nor U27103 (N_27103,N_26841,N_26912);
nand U27104 (N_27104,N_26814,N_26956);
nand U27105 (N_27105,N_26823,N_26913);
and U27106 (N_27106,N_26846,N_26909);
or U27107 (N_27107,N_26986,N_26971);
xor U27108 (N_27108,N_26967,N_26854);
nand U27109 (N_27109,N_26875,N_26979);
xnor U27110 (N_27110,N_26845,N_26936);
or U27111 (N_27111,N_26913,N_26957);
nor U27112 (N_27112,N_26827,N_26886);
nor U27113 (N_27113,N_26936,N_26979);
xor U27114 (N_27114,N_26990,N_26830);
or U27115 (N_27115,N_26880,N_26845);
or U27116 (N_27116,N_26822,N_26874);
nor U27117 (N_27117,N_26860,N_26931);
or U27118 (N_27118,N_26947,N_26986);
xnor U27119 (N_27119,N_26927,N_26836);
nand U27120 (N_27120,N_26907,N_26841);
nand U27121 (N_27121,N_26869,N_26849);
nand U27122 (N_27122,N_26887,N_26987);
or U27123 (N_27123,N_26943,N_26835);
and U27124 (N_27124,N_26943,N_26877);
xnor U27125 (N_27125,N_26994,N_26918);
or U27126 (N_27126,N_26911,N_26850);
and U27127 (N_27127,N_26959,N_26881);
or U27128 (N_27128,N_26828,N_26805);
nor U27129 (N_27129,N_26815,N_26949);
nand U27130 (N_27130,N_26900,N_26964);
or U27131 (N_27131,N_26853,N_26879);
nor U27132 (N_27132,N_26867,N_26824);
nand U27133 (N_27133,N_26851,N_26884);
xnor U27134 (N_27134,N_26827,N_26988);
nand U27135 (N_27135,N_26937,N_26900);
and U27136 (N_27136,N_26974,N_26889);
or U27137 (N_27137,N_26983,N_26914);
xnor U27138 (N_27138,N_26905,N_26955);
nand U27139 (N_27139,N_26919,N_26879);
nand U27140 (N_27140,N_26833,N_26809);
nand U27141 (N_27141,N_26956,N_26862);
nor U27142 (N_27142,N_26831,N_26835);
and U27143 (N_27143,N_26969,N_26944);
xnor U27144 (N_27144,N_26920,N_26985);
nor U27145 (N_27145,N_26840,N_26992);
xor U27146 (N_27146,N_26909,N_26987);
and U27147 (N_27147,N_26915,N_26822);
nor U27148 (N_27148,N_26831,N_26979);
nand U27149 (N_27149,N_26820,N_26943);
xor U27150 (N_27150,N_26843,N_26898);
nand U27151 (N_27151,N_26893,N_26923);
nand U27152 (N_27152,N_26939,N_26800);
xor U27153 (N_27153,N_26970,N_26818);
and U27154 (N_27154,N_26833,N_26822);
xnor U27155 (N_27155,N_26849,N_26951);
xnor U27156 (N_27156,N_26809,N_26848);
and U27157 (N_27157,N_26966,N_26913);
nand U27158 (N_27158,N_26824,N_26825);
or U27159 (N_27159,N_26834,N_26928);
or U27160 (N_27160,N_26962,N_26912);
nand U27161 (N_27161,N_26916,N_26940);
xor U27162 (N_27162,N_26944,N_26940);
xnor U27163 (N_27163,N_26885,N_26818);
xnor U27164 (N_27164,N_26857,N_26840);
xnor U27165 (N_27165,N_26806,N_26988);
nor U27166 (N_27166,N_26955,N_26980);
xor U27167 (N_27167,N_26954,N_26907);
nand U27168 (N_27168,N_26912,N_26810);
or U27169 (N_27169,N_26929,N_26984);
xor U27170 (N_27170,N_26860,N_26831);
nor U27171 (N_27171,N_26876,N_26959);
xnor U27172 (N_27172,N_26899,N_26900);
xor U27173 (N_27173,N_26983,N_26854);
nor U27174 (N_27174,N_26934,N_26855);
nand U27175 (N_27175,N_26987,N_26871);
and U27176 (N_27176,N_26936,N_26924);
xor U27177 (N_27177,N_26977,N_26903);
nor U27178 (N_27178,N_26858,N_26829);
and U27179 (N_27179,N_26972,N_26863);
nand U27180 (N_27180,N_26932,N_26828);
nand U27181 (N_27181,N_26957,N_26821);
or U27182 (N_27182,N_26985,N_26995);
xnor U27183 (N_27183,N_26962,N_26862);
and U27184 (N_27184,N_26936,N_26857);
and U27185 (N_27185,N_26996,N_26833);
nand U27186 (N_27186,N_26993,N_26889);
nor U27187 (N_27187,N_26934,N_26882);
and U27188 (N_27188,N_26990,N_26801);
nand U27189 (N_27189,N_26979,N_26870);
and U27190 (N_27190,N_26902,N_26805);
xnor U27191 (N_27191,N_26811,N_26984);
nor U27192 (N_27192,N_26865,N_26936);
xor U27193 (N_27193,N_26967,N_26862);
or U27194 (N_27194,N_26832,N_26823);
xnor U27195 (N_27195,N_26890,N_26901);
nor U27196 (N_27196,N_26856,N_26918);
xnor U27197 (N_27197,N_26878,N_26850);
nor U27198 (N_27198,N_26996,N_26819);
nor U27199 (N_27199,N_26897,N_26961);
or U27200 (N_27200,N_27072,N_27053);
nor U27201 (N_27201,N_27086,N_27098);
nand U27202 (N_27202,N_27193,N_27005);
or U27203 (N_27203,N_27081,N_27032);
and U27204 (N_27204,N_27018,N_27139);
xor U27205 (N_27205,N_27191,N_27199);
and U27206 (N_27206,N_27177,N_27112);
and U27207 (N_27207,N_27154,N_27118);
nor U27208 (N_27208,N_27100,N_27007);
or U27209 (N_27209,N_27041,N_27025);
nor U27210 (N_27210,N_27026,N_27114);
or U27211 (N_27211,N_27158,N_27084);
xor U27212 (N_27212,N_27077,N_27124);
nand U27213 (N_27213,N_27131,N_27009);
xor U27214 (N_27214,N_27049,N_27014);
nand U27215 (N_27215,N_27165,N_27070);
and U27216 (N_27216,N_27195,N_27168);
or U27217 (N_27217,N_27024,N_27006);
and U27218 (N_27218,N_27121,N_27120);
xnor U27219 (N_27219,N_27178,N_27021);
or U27220 (N_27220,N_27093,N_27132);
xnor U27221 (N_27221,N_27159,N_27003);
or U27222 (N_27222,N_27185,N_27113);
nor U27223 (N_27223,N_27115,N_27088);
or U27224 (N_27224,N_27126,N_27022);
nand U27225 (N_27225,N_27054,N_27015);
xor U27226 (N_27226,N_27128,N_27004);
nor U27227 (N_27227,N_27042,N_27001);
nor U27228 (N_27228,N_27055,N_27076);
nor U27229 (N_27229,N_27052,N_27039);
and U27230 (N_27230,N_27000,N_27133);
nand U27231 (N_27231,N_27109,N_27148);
nand U27232 (N_27232,N_27074,N_27094);
nand U27233 (N_27233,N_27030,N_27157);
xor U27234 (N_27234,N_27012,N_27136);
or U27235 (N_27235,N_27187,N_27151);
and U27236 (N_27236,N_27057,N_27138);
or U27237 (N_27237,N_27082,N_27135);
nand U27238 (N_27238,N_27079,N_27170);
or U27239 (N_27239,N_27040,N_27174);
and U27240 (N_27240,N_27125,N_27104);
or U27241 (N_27241,N_27019,N_27069);
or U27242 (N_27242,N_27087,N_27176);
nor U27243 (N_27243,N_27036,N_27107);
nand U27244 (N_27244,N_27119,N_27198);
xnor U27245 (N_27245,N_27080,N_27181);
nor U27246 (N_27246,N_27099,N_27020);
or U27247 (N_27247,N_27134,N_27173);
nand U27248 (N_27248,N_27065,N_27043);
nor U27249 (N_27249,N_27016,N_27106);
xnor U27250 (N_27250,N_27184,N_27066);
nor U27251 (N_27251,N_27153,N_27156);
nor U27252 (N_27252,N_27145,N_27146);
and U27253 (N_27253,N_27078,N_27147);
xor U27254 (N_27254,N_27142,N_27117);
and U27255 (N_27255,N_27058,N_27108);
nand U27256 (N_27256,N_27038,N_27188);
nor U27257 (N_27257,N_27123,N_27051);
nor U27258 (N_27258,N_27048,N_27116);
and U27259 (N_27259,N_27169,N_27095);
or U27260 (N_27260,N_27162,N_27029);
and U27261 (N_27261,N_27105,N_27163);
nand U27262 (N_27262,N_27179,N_27127);
and U27263 (N_27263,N_27152,N_27149);
xnor U27264 (N_27264,N_27046,N_27182);
or U27265 (N_27265,N_27194,N_27155);
nand U27266 (N_27266,N_27037,N_27062);
xor U27267 (N_27267,N_27083,N_27150);
and U27268 (N_27268,N_27089,N_27050);
nand U27269 (N_27269,N_27137,N_27110);
nand U27270 (N_27270,N_27097,N_27180);
or U27271 (N_27271,N_27059,N_27060);
xnor U27272 (N_27272,N_27017,N_27023);
xor U27273 (N_27273,N_27091,N_27045);
nor U27274 (N_27274,N_27044,N_27027);
nor U27275 (N_27275,N_27102,N_27166);
and U27276 (N_27276,N_27171,N_27172);
or U27277 (N_27277,N_27103,N_27111);
nor U27278 (N_27278,N_27028,N_27010);
nand U27279 (N_27279,N_27061,N_27047);
and U27280 (N_27280,N_27130,N_27033);
nand U27281 (N_27281,N_27063,N_27141);
nor U27282 (N_27282,N_27068,N_27192);
nand U27283 (N_27283,N_27144,N_27064);
nand U27284 (N_27284,N_27034,N_27140);
nand U27285 (N_27285,N_27008,N_27122);
xor U27286 (N_27286,N_27143,N_27175);
xor U27287 (N_27287,N_27186,N_27071);
and U27288 (N_27288,N_27013,N_27096);
or U27289 (N_27289,N_27035,N_27011);
xnor U27290 (N_27290,N_27092,N_27090);
xnor U27291 (N_27291,N_27196,N_27161);
xnor U27292 (N_27292,N_27002,N_27075);
or U27293 (N_27293,N_27101,N_27164);
nand U27294 (N_27294,N_27067,N_27073);
and U27295 (N_27295,N_27129,N_27183);
and U27296 (N_27296,N_27056,N_27190);
xnor U27297 (N_27297,N_27189,N_27031);
or U27298 (N_27298,N_27085,N_27167);
or U27299 (N_27299,N_27197,N_27160);
or U27300 (N_27300,N_27056,N_27089);
and U27301 (N_27301,N_27157,N_27192);
and U27302 (N_27302,N_27032,N_27080);
nand U27303 (N_27303,N_27047,N_27078);
or U27304 (N_27304,N_27195,N_27093);
and U27305 (N_27305,N_27059,N_27156);
nand U27306 (N_27306,N_27081,N_27085);
nor U27307 (N_27307,N_27174,N_27058);
or U27308 (N_27308,N_27050,N_27052);
xor U27309 (N_27309,N_27139,N_27182);
nor U27310 (N_27310,N_27034,N_27027);
or U27311 (N_27311,N_27186,N_27085);
and U27312 (N_27312,N_27043,N_27081);
xor U27313 (N_27313,N_27152,N_27024);
or U27314 (N_27314,N_27020,N_27042);
and U27315 (N_27315,N_27107,N_27151);
xor U27316 (N_27316,N_27105,N_27060);
and U27317 (N_27317,N_27163,N_27031);
or U27318 (N_27318,N_27021,N_27167);
or U27319 (N_27319,N_27068,N_27195);
nor U27320 (N_27320,N_27068,N_27102);
nor U27321 (N_27321,N_27116,N_27108);
nor U27322 (N_27322,N_27022,N_27136);
and U27323 (N_27323,N_27176,N_27045);
nand U27324 (N_27324,N_27191,N_27047);
xor U27325 (N_27325,N_27106,N_27197);
nor U27326 (N_27326,N_27174,N_27018);
and U27327 (N_27327,N_27175,N_27081);
nand U27328 (N_27328,N_27075,N_27182);
nor U27329 (N_27329,N_27123,N_27124);
and U27330 (N_27330,N_27021,N_27104);
nor U27331 (N_27331,N_27164,N_27131);
nand U27332 (N_27332,N_27162,N_27052);
or U27333 (N_27333,N_27034,N_27165);
nor U27334 (N_27334,N_27130,N_27095);
nor U27335 (N_27335,N_27126,N_27061);
and U27336 (N_27336,N_27131,N_27178);
and U27337 (N_27337,N_27066,N_27029);
xnor U27338 (N_27338,N_27006,N_27011);
nand U27339 (N_27339,N_27100,N_27017);
nand U27340 (N_27340,N_27171,N_27145);
xnor U27341 (N_27341,N_27100,N_27131);
or U27342 (N_27342,N_27176,N_27129);
and U27343 (N_27343,N_27182,N_27070);
nor U27344 (N_27344,N_27184,N_27091);
nand U27345 (N_27345,N_27186,N_27059);
xor U27346 (N_27346,N_27120,N_27168);
nor U27347 (N_27347,N_27043,N_27006);
and U27348 (N_27348,N_27171,N_27030);
and U27349 (N_27349,N_27179,N_27140);
xnor U27350 (N_27350,N_27184,N_27046);
nand U27351 (N_27351,N_27172,N_27022);
xor U27352 (N_27352,N_27097,N_27118);
nor U27353 (N_27353,N_27014,N_27125);
nor U27354 (N_27354,N_27080,N_27075);
nor U27355 (N_27355,N_27070,N_27151);
or U27356 (N_27356,N_27012,N_27082);
xnor U27357 (N_27357,N_27082,N_27053);
or U27358 (N_27358,N_27133,N_27078);
xor U27359 (N_27359,N_27150,N_27068);
or U27360 (N_27360,N_27193,N_27069);
or U27361 (N_27361,N_27132,N_27006);
or U27362 (N_27362,N_27175,N_27034);
and U27363 (N_27363,N_27059,N_27138);
or U27364 (N_27364,N_27167,N_27046);
xor U27365 (N_27365,N_27171,N_27165);
or U27366 (N_27366,N_27195,N_27014);
nand U27367 (N_27367,N_27087,N_27114);
nor U27368 (N_27368,N_27087,N_27026);
nand U27369 (N_27369,N_27181,N_27044);
nor U27370 (N_27370,N_27021,N_27046);
and U27371 (N_27371,N_27154,N_27052);
and U27372 (N_27372,N_27136,N_27150);
and U27373 (N_27373,N_27162,N_27011);
nor U27374 (N_27374,N_27011,N_27191);
or U27375 (N_27375,N_27127,N_27158);
nand U27376 (N_27376,N_27136,N_27005);
nor U27377 (N_27377,N_27196,N_27048);
or U27378 (N_27378,N_27150,N_27064);
xnor U27379 (N_27379,N_27005,N_27047);
nor U27380 (N_27380,N_27167,N_27047);
and U27381 (N_27381,N_27085,N_27130);
nand U27382 (N_27382,N_27014,N_27165);
or U27383 (N_27383,N_27124,N_27140);
and U27384 (N_27384,N_27033,N_27017);
or U27385 (N_27385,N_27163,N_27094);
nor U27386 (N_27386,N_27129,N_27047);
and U27387 (N_27387,N_27188,N_27084);
nor U27388 (N_27388,N_27102,N_27011);
xnor U27389 (N_27389,N_27096,N_27048);
or U27390 (N_27390,N_27064,N_27092);
nor U27391 (N_27391,N_27199,N_27018);
and U27392 (N_27392,N_27028,N_27185);
and U27393 (N_27393,N_27144,N_27125);
or U27394 (N_27394,N_27113,N_27158);
xnor U27395 (N_27395,N_27164,N_27075);
and U27396 (N_27396,N_27028,N_27169);
xnor U27397 (N_27397,N_27128,N_27172);
nor U27398 (N_27398,N_27167,N_27079);
and U27399 (N_27399,N_27077,N_27048);
or U27400 (N_27400,N_27341,N_27359);
and U27401 (N_27401,N_27288,N_27360);
nor U27402 (N_27402,N_27228,N_27293);
nor U27403 (N_27403,N_27232,N_27213);
nand U27404 (N_27404,N_27371,N_27352);
and U27405 (N_27405,N_27308,N_27239);
nor U27406 (N_27406,N_27281,N_27255);
and U27407 (N_27407,N_27248,N_27350);
nand U27408 (N_27408,N_27209,N_27249);
or U27409 (N_27409,N_27253,N_27276);
xor U27410 (N_27410,N_27234,N_27212);
xnor U27411 (N_27411,N_27282,N_27317);
and U27412 (N_27412,N_27366,N_27292);
nand U27413 (N_27413,N_27378,N_27278);
nand U27414 (N_27414,N_27358,N_27349);
xnor U27415 (N_27415,N_27300,N_27285);
xnor U27416 (N_27416,N_27303,N_27398);
and U27417 (N_27417,N_27363,N_27345);
and U27418 (N_27418,N_27327,N_27319);
nand U27419 (N_27419,N_27214,N_27251);
nor U27420 (N_27420,N_27357,N_27268);
or U27421 (N_27421,N_27344,N_27325);
and U27422 (N_27422,N_27295,N_27339);
and U27423 (N_27423,N_27326,N_27254);
nand U27424 (N_27424,N_27338,N_27242);
or U27425 (N_27425,N_27312,N_27284);
xor U27426 (N_27426,N_27305,N_27205);
xor U27427 (N_27427,N_27369,N_27376);
or U27428 (N_27428,N_27310,N_27320);
or U27429 (N_27429,N_27279,N_27272);
or U27430 (N_27430,N_27348,N_27375);
xnor U27431 (N_27431,N_27260,N_27223);
nor U27432 (N_27432,N_27383,N_27216);
xor U27433 (N_27433,N_27315,N_27298);
or U27434 (N_27434,N_27393,N_27266);
or U27435 (N_27435,N_27217,N_27336);
and U27436 (N_27436,N_27335,N_27211);
or U27437 (N_27437,N_27238,N_27222);
xor U27438 (N_27438,N_27373,N_27215);
xor U27439 (N_27439,N_27334,N_27322);
or U27440 (N_27440,N_27311,N_27271);
nor U27441 (N_27441,N_27245,N_27200);
or U27442 (N_27442,N_27247,N_27246);
nor U27443 (N_27443,N_27269,N_27367);
nor U27444 (N_27444,N_27351,N_27356);
nand U27445 (N_27445,N_27289,N_27264);
nand U27446 (N_27446,N_27353,N_27390);
nor U27447 (N_27447,N_27202,N_27386);
nor U27448 (N_27448,N_27370,N_27394);
nor U27449 (N_27449,N_27226,N_27208);
nor U27450 (N_27450,N_27224,N_27297);
nor U27451 (N_27451,N_27291,N_27387);
nor U27452 (N_27452,N_27362,N_27250);
xor U27453 (N_27453,N_27231,N_27261);
and U27454 (N_27454,N_27275,N_27219);
or U27455 (N_27455,N_27267,N_27391);
and U27456 (N_27456,N_27230,N_27309);
nand U27457 (N_27457,N_27368,N_27354);
and U27458 (N_27458,N_27204,N_27385);
and U27459 (N_27459,N_27258,N_27330);
xnor U27460 (N_27460,N_27206,N_27361);
nor U27461 (N_27461,N_27381,N_27240);
xor U27462 (N_27462,N_27388,N_27286);
nand U27463 (N_27463,N_27233,N_27280);
nor U27464 (N_27464,N_27283,N_27379);
or U27465 (N_27465,N_27333,N_27220);
nand U27466 (N_27466,N_27244,N_27331);
xor U27467 (N_27467,N_27304,N_27287);
nand U27468 (N_27468,N_27301,N_27347);
or U27469 (N_27469,N_27340,N_27395);
nor U27470 (N_27470,N_27365,N_27377);
and U27471 (N_27471,N_27324,N_27364);
nor U27472 (N_27472,N_27316,N_27203);
nor U27473 (N_27473,N_27399,N_27396);
or U27474 (N_27474,N_27372,N_27397);
or U27475 (N_27475,N_27241,N_27290);
nor U27476 (N_27476,N_27307,N_27218);
nand U27477 (N_27477,N_27299,N_27389);
and U27478 (N_27478,N_27207,N_27229);
and U27479 (N_27479,N_27263,N_27256);
nor U27480 (N_27480,N_27296,N_27355);
xor U27481 (N_27481,N_27294,N_27265);
or U27482 (N_27482,N_27346,N_27227);
or U27483 (N_27483,N_27318,N_27392);
and U27484 (N_27484,N_27337,N_27328);
xnor U27485 (N_27485,N_27382,N_27313);
nand U27486 (N_27486,N_27321,N_27380);
or U27487 (N_27487,N_27374,N_27332);
or U27488 (N_27488,N_27210,N_27236);
and U27489 (N_27489,N_27235,N_27323);
and U27490 (N_27490,N_27252,N_27243);
nand U27491 (N_27491,N_27274,N_27302);
or U27492 (N_27492,N_27201,N_27221);
and U27493 (N_27493,N_27270,N_27342);
xor U27494 (N_27494,N_27343,N_27306);
nor U27495 (N_27495,N_27257,N_27237);
xnor U27496 (N_27496,N_27259,N_27314);
or U27497 (N_27497,N_27273,N_27225);
xor U27498 (N_27498,N_27277,N_27384);
and U27499 (N_27499,N_27329,N_27262);
nor U27500 (N_27500,N_27372,N_27366);
xnor U27501 (N_27501,N_27306,N_27313);
xnor U27502 (N_27502,N_27358,N_27203);
and U27503 (N_27503,N_27394,N_27379);
xor U27504 (N_27504,N_27272,N_27300);
nor U27505 (N_27505,N_27206,N_27251);
nand U27506 (N_27506,N_27389,N_27336);
or U27507 (N_27507,N_27208,N_27366);
nand U27508 (N_27508,N_27344,N_27214);
nand U27509 (N_27509,N_27391,N_27202);
and U27510 (N_27510,N_27353,N_27227);
nand U27511 (N_27511,N_27207,N_27336);
xnor U27512 (N_27512,N_27222,N_27327);
xnor U27513 (N_27513,N_27267,N_27288);
and U27514 (N_27514,N_27229,N_27291);
nand U27515 (N_27515,N_27327,N_27317);
nor U27516 (N_27516,N_27222,N_27365);
and U27517 (N_27517,N_27212,N_27374);
and U27518 (N_27518,N_27397,N_27282);
nand U27519 (N_27519,N_27238,N_27302);
or U27520 (N_27520,N_27391,N_27264);
or U27521 (N_27521,N_27375,N_27270);
xor U27522 (N_27522,N_27324,N_27391);
or U27523 (N_27523,N_27274,N_27209);
nor U27524 (N_27524,N_27330,N_27370);
nor U27525 (N_27525,N_27265,N_27273);
nand U27526 (N_27526,N_27288,N_27225);
nand U27527 (N_27527,N_27265,N_27200);
and U27528 (N_27528,N_27329,N_27293);
nor U27529 (N_27529,N_27389,N_27286);
and U27530 (N_27530,N_27250,N_27332);
and U27531 (N_27531,N_27352,N_27261);
xor U27532 (N_27532,N_27311,N_27220);
and U27533 (N_27533,N_27352,N_27364);
and U27534 (N_27534,N_27394,N_27377);
and U27535 (N_27535,N_27396,N_27386);
xnor U27536 (N_27536,N_27333,N_27319);
and U27537 (N_27537,N_27397,N_27252);
xor U27538 (N_27538,N_27345,N_27385);
nand U27539 (N_27539,N_27347,N_27298);
or U27540 (N_27540,N_27212,N_27355);
or U27541 (N_27541,N_27252,N_27262);
nand U27542 (N_27542,N_27221,N_27203);
or U27543 (N_27543,N_27219,N_27378);
xor U27544 (N_27544,N_27331,N_27351);
xnor U27545 (N_27545,N_27391,N_27339);
nor U27546 (N_27546,N_27283,N_27313);
nand U27547 (N_27547,N_27290,N_27270);
or U27548 (N_27548,N_27222,N_27333);
xnor U27549 (N_27549,N_27257,N_27290);
nor U27550 (N_27550,N_27257,N_27303);
nor U27551 (N_27551,N_27354,N_27269);
and U27552 (N_27552,N_27379,N_27262);
and U27553 (N_27553,N_27332,N_27214);
nand U27554 (N_27554,N_27271,N_27224);
and U27555 (N_27555,N_27337,N_27373);
xor U27556 (N_27556,N_27262,N_27279);
and U27557 (N_27557,N_27291,N_27357);
xnor U27558 (N_27558,N_27364,N_27397);
xor U27559 (N_27559,N_27238,N_27243);
or U27560 (N_27560,N_27243,N_27262);
xnor U27561 (N_27561,N_27335,N_27394);
xor U27562 (N_27562,N_27366,N_27248);
nand U27563 (N_27563,N_27244,N_27286);
or U27564 (N_27564,N_27203,N_27284);
nor U27565 (N_27565,N_27277,N_27259);
nor U27566 (N_27566,N_27347,N_27391);
or U27567 (N_27567,N_27275,N_27224);
and U27568 (N_27568,N_27255,N_27339);
xor U27569 (N_27569,N_27293,N_27206);
nor U27570 (N_27570,N_27209,N_27284);
nor U27571 (N_27571,N_27244,N_27262);
or U27572 (N_27572,N_27266,N_27301);
or U27573 (N_27573,N_27222,N_27360);
and U27574 (N_27574,N_27281,N_27356);
nor U27575 (N_27575,N_27321,N_27260);
or U27576 (N_27576,N_27342,N_27389);
nor U27577 (N_27577,N_27294,N_27301);
nand U27578 (N_27578,N_27332,N_27243);
or U27579 (N_27579,N_27231,N_27298);
and U27580 (N_27580,N_27389,N_27244);
xor U27581 (N_27581,N_27383,N_27354);
or U27582 (N_27582,N_27284,N_27288);
nand U27583 (N_27583,N_27340,N_27348);
and U27584 (N_27584,N_27268,N_27320);
nor U27585 (N_27585,N_27242,N_27232);
nor U27586 (N_27586,N_27316,N_27254);
and U27587 (N_27587,N_27368,N_27383);
nor U27588 (N_27588,N_27377,N_27217);
nand U27589 (N_27589,N_27244,N_27231);
xnor U27590 (N_27590,N_27334,N_27249);
nor U27591 (N_27591,N_27281,N_27301);
or U27592 (N_27592,N_27352,N_27321);
or U27593 (N_27593,N_27363,N_27334);
nand U27594 (N_27594,N_27229,N_27336);
xnor U27595 (N_27595,N_27278,N_27259);
xor U27596 (N_27596,N_27290,N_27317);
and U27597 (N_27597,N_27344,N_27219);
xnor U27598 (N_27598,N_27285,N_27222);
nor U27599 (N_27599,N_27374,N_27224);
xnor U27600 (N_27600,N_27592,N_27409);
nand U27601 (N_27601,N_27405,N_27426);
nor U27602 (N_27602,N_27581,N_27465);
or U27603 (N_27603,N_27499,N_27596);
nand U27604 (N_27604,N_27571,N_27563);
nor U27605 (N_27605,N_27521,N_27555);
xor U27606 (N_27606,N_27545,N_27515);
xnor U27607 (N_27607,N_27505,N_27480);
xor U27608 (N_27608,N_27501,N_27527);
or U27609 (N_27609,N_27458,N_27456);
xnor U27610 (N_27610,N_27554,N_27478);
or U27611 (N_27611,N_27489,N_27540);
nor U27612 (N_27612,N_27526,N_27512);
nand U27613 (N_27613,N_27446,N_27528);
nor U27614 (N_27614,N_27510,N_27536);
and U27615 (N_27615,N_27522,N_27552);
or U27616 (N_27616,N_27508,N_27543);
nand U27617 (N_27617,N_27408,N_27564);
or U27618 (N_27618,N_27578,N_27441);
nor U27619 (N_27619,N_27461,N_27460);
nand U27620 (N_27620,N_27407,N_27470);
nand U27621 (N_27621,N_27587,N_27491);
nand U27622 (N_27622,N_27556,N_27567);
nand U27623 (N_27623,N_27516,N_27582);
and U27624 (N_27624,N_27568,N_27422);
nand U27625 (N_27625,N_27463,N_27573);
and U27626 (N_27626,N_27503,N_27479);
or U27627 (N_27627,N_27448,N_27520);
nor U27628 (N_27628,N_27466,N_27544);
or U27629 (N_27629,N_27450,N_27496);
and U27630 (N_27630,N_27502,N_27588);
or U27631 (N_27631,N_27454,N_27432);
or U27632 (N_27632,N_27551,N_27420);
xor U27633 (N_27633,N_27506,N_27418);
or U27634 (N_27634,N_27597,N_27468);
or U27635 (N_27635,N_27590,N_27416);
or U27636 (N_27636,N_27434,N_27439);
and U27637 (N_27637,N_27451,N_27484);
xor U27638 (N_27638,N_27561,N_27403);
xor U27639 (N_27639,N_27531,N_27539);
nor U27640 (N_27640,N_27595,N_27433);
and U27641 (N_27641,N_27507,N_27594);
xor U27642 (N_27642,N_27449,N_27469);
or U27643 (N_27643,N_27438,N_27437);
nand U27644 (N_27644,N_27482,N_27428);
and U27645 (N_27645,N_27430,N_27411);
nor U27646 (N_27646,N_27589,N_27406);
nand U27647 (N_27647,N_27474,N_27517);
nor U27648 (N_27648,N_27523,N_27566);
or U27649 (N_27649,N_27445,N_27464);
nor U27650 (N_27650,N_27572,N_27574);
nand U27651 (N_27651,N_27562,N_27580);
xor U27652 (N_27652,N_27546,N_27443);
xnor U27653 (N_27653,N_27452,N_27534);
xnor U27654 (N_27654,N_27490,N_27593);
or U27655 (N_27655,N_27471,N_27419);
and U27656 (N_27656,N_27410,N_27511);
nand U27657 (N_27657,N_27475,N_27500);
nor U27658 (N_27658,N_27453,N_27569);
or U27659 (N_27659,N_27504,N_27598);
nor U27660 (N_27660,N_27467,N_27415);
xnor U27661 (N_27661,N_27591,N_27519);
and U27662 (N_27662,N_27525,N_27585);
or U27663 (N_27663,N_27542,N_27583);
and U27664 (N_27664,N_27404,N_27457);
or U27665 (N_27665,N_27518,N_27497);
nor U27666 (N_27666,N_27565,N_27462);
xor U27667 (N_27667,N_27401,N_27548);
xnor U27668 (N_27668,N_27485,N_27557);
xnor U27669 (N_27669,N_27486,N_27493);
and U27670 (N_27670,N_27514,N_27498);
nand U27671 (N_27671,N_27429,N_27413);
nor U27672 (N_27672,N_27442,N_27412);
or U27673 (N_27673,N_27559,N_27427);
and U27674 (N_27674,N_27477,N_27538);
nor U27675 (N_27675,N_27553,N_27547);
xnor U27676 (N_27676,N_27492,N_27535);
xnor U27677 (N_27677,N_27487,N_27481);
nand U27678 (N_27678,N_27575,N_27577);
and U27679 (N_27679,N_27440,N_27533);
nand U27680 (N_27680,N_27530,N_27400);
or U27681 (N_27681,N_27476,N_27560);
and U27682 (N_27682,N_27459,N_27550);
and U27683 (N_27683,N_27532,N_27435);
and U27684 (N_27684,N_27579,N_27488);
xnor U27685 (N_27685,N_27584,N_27509);
xor U27686 (N_27686,N_27423,N_27494);
nor U27687 (N_27687,N_27402,N_27549);
nand U27688 (N_27688,N_27436,N_27513);
nand U27689 (N_27689,N_27529,N_27473);
nor U27690 (N_27690,N_27444,N_27417);
nand U27691 (N_27691,N_27424,N_27425);
nor U27692 (N_27692,N_27495,N_27455);
xor U27693 (N_27693,N_27558,N_27472);
xor U27694 (N_27694,N_27431,N_27414);
and U27695 (N_27695,N_27483,N_27570);
nor U27696 (N_27696,N_27586,N_27599);
or U27697 (N_27697,N_27537,N_27541);
or U27698 (N_27698,N_27524,N_27447);
nand U27699 (N_27699,N_27576,N_27421);
or U27700 (N_27700,N_27506,N_27501);
nor U27701 (N_27701,N_27529,N_27466);
and U27702 (N_27702,N_27557,N_27509);
xnor U27703 (N_27703,N_27411,N_27594);
xor U27704 (N_27704,N_27519,N_27542);
xnor U27705 (N_27705,N_27471,N_27579);
or U27706 (N_27706,N_27412,N_27482);
nand U27707 (N_27707,N_27435,N_27412);
nand U27708 (N_27708,N_27449,N_27575);
and U27709 (N_27709,N_27466,N_27567);
or U27710 (N_27710,N_27578,N_27547);
nand U27711 (N_27711,N_27544,N_27586);
or U27712 (N_27712,N_27492,N_27527);
xnor U27713 (N_27713,N_27427,N_27494);
and U27714 (N_27714,N_27520,N_27483);
nand U27715 (N_27715,N_27483,N_27498);
nand U27716 (N_27716,N_27568,N_27548);
nor U27717 (N_27717,N_27511,N_27426);
xnor U27718 (N_27718,N_27572,N_27428);
nand U27719 (N_27719,N_27542,N_27409);
or U27720 (N_27720,N_27480,N_27474);
and U27721 (N_27721,N_27466,N_27598);
nor U27722 (N_27722,N_27594,N_27587);
or U27723 (N_27723,N_27530,N_27442);
and U27724 (N_27724,N_27542,N_27556);
nand U27725 (N_27725,N_27444,N_27481);
nand U27726 (N_27726,N_27566,N_27585);
or U27727 (N_27727,N_27505,N_27513);
and U27728 (N_27728,N_27520,N_27406);
and U27729 (N_27729,N_27536,N_27408);
nor U27730 (N_27730,N_27498,N_27561);
xnor U27731 (N_27731,N_27405,N_27517);
or U27732 (N_27732,N_27416,N_27497);
and U27733 (N_27733,N_27409,N_27422);
nor U27734 (N_27734,N_27436,N_27464);
and U27735 (N_27735,N_27590,N_27460);
or U27736 (N_27736,N_27570,N_27575);
and U27737 (N_27737,N_27522,N_27535);
and U27738 (N_27738,N_27435,N_27553);
and U27739 (N_27739,N_27542,N_27445);
and U27740 (N_27740,N_27552,N_27545);
xor U27741 (N_27741,N_27506,N_27575);
nand U27742 (N_27742,N_27452,N_27580);
nand U27743 (N_27743,N_27485,N_27438);
nor U27744 (N_27744,N_27460,N_27537);
and U27745 (N_27745,N_27535,N_27497);
nor U27746 (N_27746,N_27472,N_27491);
nand U27747 (N_27747,N_27521,N_27423);
xnor U27748 (N_27748,N_27595,N_27512);
xor U27749 (N_27749,N_27530,N_27476);
or U27750 (N_27750,N_27565,N_27443);
and U27751 (N_27751,N_27463,N_27554);
nor U27752 (N_27752,N_27578,N_27555);
nor U27753 (N_27753,N_27594,N_27469);
xor U27754 (N_27754,N_27489,N_27543);
and U27755 (N_27755,N_27428,N_27450);
nand U27756 (N_27756,N_27574,N_27596);
and U27757 (N_27757,N_27559,N_27570);
xnor U27758 (N_27758,N_27467,N_27468);
nor U27759 (N_27759,N_27465,N_27543);
and U27760 (N_27760,N_27480,N_27558);
nor U27761 (N_27761,N_27560,N_27537);
nand U27762 (N_27762,N_27579,N_27571);
or U27763 (N_27763,N_27598,N_27437);
xor U27764 (N_27764,N_27435,N_27444);
or U27765 (N_27765,N_27465,N_27416);
or U27766 (N_27766,N_27592,N_27483);
xor U27767 (N_27767,N_27503,N_27536);
nor U27768 (N_27768,N_27567,N_27434);
nor U27769 (N_27769,N_27409,N_27506);
and U27770 (N_27770,N_27469,N_27506);
nor U27771 (N_27771,N_27579,N_27481);
and U27772 (N_27772,N_27522,N_27486);
xnor U27773 (N_27773,N_27456,N_27495);
nand U27774 (N_27774,N_27524,N_27556);
nor U27775 (N_27775,N_27524,N_27404);
and U27776 (N_27776,N_27549,N_27417);
and U27777 (N_27777,N_27466,N_27427);
nand U27778 (N_27778,N_27479,N_27427);
and U27779 (N_27779,N_27443,N_27415);
or U27780 (N_27780,N_27428,N_27570);
nand U27781 (N_27781,N_27474,N_27580);
nor U27782 (N_27782,N_27554,N_27481);
xnor U27783 (N_27783,N_27589,N_27549);
nor U27784 (N_27784,N_27421,N_27536);
nor U27785 (N_27785,N_27578,N_27505);
xor U27786 (N_27786,N_27580,N_27456);
nand U27787 (N_27787,N_27591,N_27556);
and U27788 (N_27788,N_27413,N_27557);
nor U27789 (N_27789,N_27466,N_27422);
or U27790 (N_27790,N_27478,N_27574);
xor U27791 (N_27791,N_27441,N_27489);
xor U27792 (N_27792,N_27544,N_27552);
nand U27793 (N_27793,N_27477,N_27579);
or U27794 (N_27794,N_27578,N_27515);
xor U27795 (N_27795,N_27418,N_27449);
and U27796 (N_27796,N_27405,N_27432);
xor U27797 (N_27797,N_27470,N_27467);
xnor U27798 (N_27798,N_27548,N_27562);
and U27799 (N_27799,N_27562,N_27473);
or U27800 (N_27800,N_27739,N_27724);
nand U27801 (N_27801,N_27675,N_27779);
or U27802 (N_27802,N_27690,N_27617);
or U27803 (N_27803,N_27658,N_27758);
or U27804 (N_27804,N_27659,N_27694);
or U27805 (N_27805,N_27773,N_27640);
and U27806 (N_27806,N_27746,N_27627);
or U27807 (N_27807,N_27601,N_27767);
nand U27808 (N_27808,N_27700,N_27791);
nand U27809 (N_27809,N_27660,N_27693);
nor U27810 (N_27810,N_27705,N_27719);
nor U27811 (N_27811,N_27649,N_27768);
xor U27812 (N_27812,N_27682,N_27666);
nand U27813 (N_27813,N_27743,N_27657);
nand U27814 (N_27814,N_27684,N_27661);
and U27815 (N_27815,N_27790,N_27760);
or U27816 (N_27816,N_27706,N_27629);
or U27817 (N_27817,N_27685,N_27793);
nand U27818 (N_27818,N_27704,N_27643);
and U27819 (N_27819,N_27770,N_27678);
or U27820 (N_27820,N_27725,N_27784);
and U27821 (N_27821,N_27796,N_27618);
nand U27822 (N_27822,N_27736,N_27697);
xor U27823 (N_27823,N_27799,N_27783);
nand U27824 (N_27824,N_27703,N_27774);
nand U27825 (N_27825,N_27655,N_27639);
nor U27826 (N_27826,N_27707,N_27623);
xnor U27827 (N_27827,N_27789,N_27716);
or U27828 (N_27828,N_27794,N_27677);
or U27829 (N_27829,N_27651,N_27692);
nand U27830 (N_27830,N_27745,N_27727);
nor U27831 (N_27831,N_27734,N_27765);
and U27832 (N_27832,N_27709,N_27762);
or U27833 (N_27833,N_27645,N_27664);
nand U27834 (N_27834,N_27711,N_27720);
nor U27835 (N_27835,N_27747,N_27691);
nor U27836 (N_27836,N_27652,N_27624);
and U27837 (N_27837,N_27613,N_27728);
or U27838 (N_27838,N_27735,N_27607);
or U27839 (N_27839,N_27679,N_27619);
or U27840 (N_27840,N_27782,N_27680);
and U27841 (N_27841,N_27754,N_27688);
or U27842 (N_27842,N_27670,N_27781);
nand U27843 (N_27843,N_27798,N_27753);
nor U27844 (N_27844,N_27718,N_27778);
xnor U27845 (N_27845,N_27600,N_27638);
nor U27846 (N_27846,N_27750,N_27671);
nor U27847 (N_27847,N_27674,N_27775);
or U27848 (N_27848,N_27786,N_27737);
nand U27849 (N_27849,N_27702,N_27662);
or U27850 (N_27850,N_27656,N_27631);
and U27851 (N_27851,N_27712,N_27695);
nor U27852 (N_27852,N_27628,N_27733);
nor U27853 (N_27853,N_27771,N_27766);
and U27854 (N_27854,N_27654,N_27769);
and U27855 (N_27855,N_27797,N_27731);
nand U27856 (N_27856,N_27622,N_27792);
and U27857 (N_27857,N_27787,N_27641);
nor U27858 (N_27858,N_27681,N_27777);
nand U27859 (N_27859,N_27603,N_27650);
and U27860 (N_27860,N_27636,N_27633);
and U27861 (N_27861,N_27698,N_27673);
nor U27862 (N_27862,N_27708,N_27742);
xnor U27863 (N_27863,N_27756,N_27757);
nor U27864 (N_27864,N_27683,N_27780);
or U27865 (N_27865,N_27776,N_27621);
and U27866 (N_27866,N_27729,N_27625);
and U27867 (N_27867,N_27614,N_27665);
nor U27868 (N_27868,N_27772,N_27667);
or U27869 (N_27869,N_27676,N_27606);
nand U27870 (N_27870,N_27696,N_27630);
nand U27871 (N_27871,N_27726,N_27751);
and U27872 (N_27872,N_27668,N_27605);
xnor U27873 (N_27873,N_27795,N_27710);
and U27874 (N_27874,N_27608,N_27730);
nor U27875 (N_27875,N_27604,N_27744);
and U27876 (N_27876,N_27646,N_27602);
or U27877 (N_27877,N_27740,N_27722);
xnor U27878 (N_27878,N_27616,N_27612);
nand U27879 (N_27879,N_27669,N_27763);
nor U27880 (N_27880,N_27723,N_27715);
nor U27881 (N_27881,N_27755,N_27635);
nor U27882 (N_27882,N_27672,N_27748);
xor U27883 (N_27883,N_27689,N_27701);
or U27884 (N_27884,N_27761,N_27713);
nand U27885 (N_27885,N_27637,N_27741);
or U27886 (N_27886,N_27653,N_27610);
nand U27887 (N_27887,N_27714,N_27699);
xnor U27888 (N_27888,N_27644,N_27609);
nor U27889 (N_27889,N_27717,N_27615);
nand U27890 (N_27890,N_27749,N_27663);
xnor U27891 (N_27891,N_27648,N_27647);
nor U27892 (N_27892,N_27642,N_27785);
xnor U27893 (N_27893,N_27759,N_27632);
and U27894 (N_27894,N_27611,N_27686);
nor U27895 (N_27895,N_27764,N_27634);
nor U27896 (N_27896,N_27721,N_27738);
nor U27897 (N_27897,N_27620,N_27788);
xor U27898 (N_27898,N_27732,N_27687);
xor U27899 (N_27899,N_27626,N_27752);
nand U27900 (N_27900,N_27794,N_27624);
nor U27901 (N_27901,N_27629,N_27630);
nor U27902 (N_27902,N_27698,N_27666);
nor U27903 (N_27903,N_27655,N_27734);
nor U27904 (N_27904,N_27762,N_27726);
nor U27905 (N_27905,N_27749,N_27668);
nand U27906 (N_27906,N_27675,N_27785);
nand U27907 (N_27907,N_27695,N_27613);
nand U27908 (N_27908,N_27736,N_27790);
xnor U27909 (N_27909,N_27788,N_27781);
and U27910 (N_27910,N_27611,N_27776);
and U27911 (N_27911,N_27637,N_27606);
and U27912 (N_27912,N_27786,N_27731);
and U27913 (N_27913,N_27618,N_27747);
nand U27914 (N_27914,N_27634,N_27736);
and U27915 (N_27915,N_27659,N_27734);
nor U27916 (N_27916,N_27789,N_27765);
or U27917 (N_27917,N_27699,N_27629);
and U27918 (N_27918,N_27752,N_27704);
xor U27919 (N_27919,N_27606,N_27683);
xor U27920 (N_27920,N_27650,N_27617);
and U27921 (N_27921,N_27704,N_27608);
nor U27922 (N_27922,N_27746,N_27714);
nand U27923 (N_27923,N_27706,N_27665);
or U27924 (N_27924,N_27747,N_27744);
xnor U27925 (N_27925,N_27608,N_27751);
xor U27926 (N_27926,N_27733,N_27677);
and U27927 (N_27927,N_27709,N_27650);
nor U27928 (N_27928,N_27614,N_27609);
or U27929 (N_27929,N_27678,N_27773);
or U27930 (N_27930,N_27757,N_27680);
and U27931 (N_27931,N_27656,N_27798);
xor U27932 (N_27932,N_27671,N_27666);
nor U27933 (N_27933,N_27700,N_27631);
xor U27934 (N_27934,N_27666,N_27601);
nor U27935 (N_27935,N_27798,N_27770);
nor U27936 (N_27936,N_27717,N_27780);
xnor U27937 (N_27937,N_27739,N_27768);
and U27938 (N_27938,N_27694,N_27625);
or U27939 (N_27939,N_27703,N_27730);
and U27940 (N_27940,N_27615,N_27709);
and U27941 (N_27941,N_27724,N_27714);
nand U27942 (N_27942,N_27707,N_27762);
xor U27943 (N_27943,N_27659,N_27623);
nor U27944 (N_27944,N_27794,N_27634);
nand U27945 (N_27945,N_27661,N_27727);
xnor U27946 (N_27946,N_27723,N_27627);
nand U27947 (N_27947,N_27798,N_27713);
nand U27948 (N_27948,N_27645,N_27796);
and U27949 (N_27949,N_27742,N_27614);
or U27950 (N_27950,N_27724,N_27750);
and U27951 (N_27951,N_27688,N_27708);
xor U27952 (N_27952,N_27769,N_27718);
and U27953 (N_27953,N_27645,N_27748);
or U27954 (N_27954,N_27742,N_27799);
and U27955 (N_27955,N_27794,N_27704);
xor U27956 (N_27956,N_27689,N_27613);
nand U27957 (N_27957,N_27755,N_27768);
xnor U27958 (N_27958,N_27682,N_27610);
nand U27959 (N_27959,N_27701,N_27753);
nor U27960 (N_27960,N_27651,N_27687);
nand U27961 (N_27961,N_27732,N_27624);
nand U27962 (N_27962,N_27754,N_27795);
and U27963 (N_27963,N_27770,N_27609);
nor U27964 (N_27964,N_27675,N_27633);
nand U27965 (N_27965,N_27656,N_27787);
nor U27966 (N_27966,N_27684,N_27637);
nand U27967 (N_27967,N_27777,N_27643);
nor U27968 (N_27968,N_27770,N_27721);
nor U27969 (N_27969,N_27785,N_27789);
nor U27970 (N_27970,N_27719,N_27710);
nand U27971 (N_27971,N_27785,N_27701);
nand U27972 (N_27972,N_27621,N_27742);
or U27973 (N_27973,N_27640,N_27695);
and U27974 (N_27974,N_27780,N_27755);
nand U27975 (N_27975,N_27759,N_27789);
nand U27976 (N_27976,N_27613,N_27690);
nand U27977 (N_27977,N_27724,N_27600);
or U27978 (N_27978,N_27726,N_27720);
nand U27979 (N_27979,N_27758,N_27749);
and U27980 (N_27980,N_27775,N_27640);
or U27981 (N_27981,N_27743,N_27634);
xor U27982 (N_27982,N_27728,N_27789);
and U27983 (N_27983,N_27740,N_27677);
xnor U27984 (N_27984,N_27622,N_27640);
or U27985 (N_27985,N_27692,N_27752);
or U27986 (N_27986,N_27681,N_27799);
nand U27987 (N_27987,N_27604,N_27785);
xor U27988 (N_27988,N_27665,N_27764);
nand U27989 (N_27989,N_27698,N_27756);
and U27990 (N_27990,N_27602,N_27604);
xor U27991 (N_27991,N_27684,N_27682);
and U27992 (N_27992,N_27618,N_27606);
xnor U27993 (N_27993,N_27778,N_27610);
nand U27994 (N_27994,N_27763,N_27604);
nand U27995 (N_27995,N_27797,N_27746);
and U27996 (N_27996,N_27670,N_27720);
or U27997 (N_27997,N_27730,N_27754);
nand U27998 (N_27998,N_27793,N_27618);
xor U27999 (N_27999,N_27716,N_27648);
or U28000 (N_28000,N_27949,N_27897);
nor U28001 (N_28001,N_27907,N_27978);
xor U28002 (N_28002,N_27803,N_27915);
nand U28003 (N_28003,N_27989,N_27863);
nor U28004 (N_28004,N_27995,N_27976);
nor U28005 (N_28005,N_27974,N_27955);
xnor U28006 (N_28006,N_27925,N_27893);
xor U28007 (N_28007,N_27876,N_27873);
and U28008 (N_28008,N_27952,N_27832);
or U28009 (N_28009,N_27875,N_27850);
xnor U28010 (N_28010,N_27807,N_27862);
or U28011 (N_28011,N_27804,N_27835);
nand U28012 (N_28012,N_27855,N_27825);
xor U28013 (N_28013,N_27878,N_27840);
nand U28014 (N_28014,N_27919,N_27826);
nand U28015 (N_28015,N_27802,N_27951);
or U28016 (N_28016,N_27818,N_27821);
xnor U28017 (N_28017,N_27865,N_27911);
and U28018 (N_28018,N_27847,N_27932);
nor U28019 (N_28019,N_27819,N_27827);
xor U28020 (N_28020,N_27947,N_27861);
nand U28021 (N_28021,N_27894,N_27845);
nor U28022 (N_28022,N_27910,N_27813);
nor U28023 (N_28023,N_27954,N_27998);
or U28024 (N_28024,N_27872,N_27985);
or U28025 (N_28025,N_27880,N_27944);
nand U28026 (N_28026,N_27886,N_27814);
and U28027 (N_28027,N_27999,N_27990);
xor U28028 (N_28028,N_27896,N_27948);
or U28029 (N_28029,N_27820,N_27960);
xor U28030 (N_28030,N_27868,N_27902);
xor U28031 (N_28031,N_27913,N_27950);
nand U28032 (N_28032,N_27830,N_27882);
nor U28033 (N_28033,N_27953,N_27992);
nand U28034 (N_28034,N_27943,N_27899);
nor U28035 (N_28035,N_27846,N_27848);
nand U28036 (N_28036,N_27997,N_27933);
or U28037 (N_28037,N_27839,N_27986);
nor U28038 (N_28038,N_27929,N_27833);
xor U28039 (N_28039,N_27962,N_27972);
nor U28040 (N_28040,N_27810,N_27869);
or U28041 (N_28041,N_27969,N_27916);
nor U28042 (N_28042,N_27966,N_27900);
xor U28043 (N_28043,N_27898,N_27816);
and U28044 (N_28044,N_27815,N_27812);
or U28045 (N_28045,N_27852,N_27928);
and U28046 (N_28046,N_27866,N_27838);
nand U28047 (N_28047,N_27965,N_27977);
nand U28048 (N_28048,N_27936,N_27841);
or U28049 (N_28049,N_27888,N_27891);
and U28050 (N_28050,N_27856,N_27987);
nor U28051 (N_28051,N_27982,N_27889);
or U28052 (N_28052,N_27935,N_27946);
nand U28053 (N_28053,N_27924,N_27834);
and U28054 (N_28054,N_27828,N_27959);
or U28055 (N_28055,N_27945,N_27958);
nand U28056 (N_28056,N_27883,N_27851);
or U28057 (N_28057,N_27912,N_27906);
and U28058 (N_28058,N_27890,N_27901);
and U28059 (N_28059,N_27908,N_27979);
xnor U28060 (N_28060,N_27967,N_27808);
nand U28061 (N_28061,N_27991,N_27922);
nand U28062 (N_28062,N_27994,N_27817);
xnor U28063 (N_28063,N_27871,N_27975);
nor U28064 (N_28064,N_27983,N_27957);
and U28065 (N_28065,N_27971,N_27937);
and U28066 (N_28066,N_27874,N_27988);
and U28067 (N_28067,N_27927,N_27842);
nor U28068 (N_28068,N_27917,N_27973);
or U28069 (N_28069,N_27800,N_27941);
nor U28070 (N_28070,N_27805,N_27921);
nand U28071 (N_28071,N_27823,N_27864);
nor U28072 (N_28072,N_27956,N_27867);
nor U28073 (N_28073,N_27887,N_27831);
nor U28074 (N_28074,N_27843,N_27881);
nor U28075 (N_28075,N_27980,N_27892);
xnor U28076 (N_28076,N_27809,N_27844);
nand U28077 (N_28077,N_27858,N_27926);
xnor U28078 (N_28078,N_27879,N_27837);
nor U28079 (N_28079,N_27970,N_27918);
xnor U28080 (N_28080,N_27806,N_27860);
xor U28081 (N_28081,N_27909,N_27877);
and U28082 (N_28082,N_27829,N_27836);
or U28083 (N_28083,N_27904,N_27961);
xor U28084 (N_28084,N_27964,N_27993);
nand U28085 (N_28085,N_27968,N_27801);
nand U28086 (N_28086,N_27996,N_27859);
xor U28087 (N_28087,N_27811,N_27903);
nor U28088 (N_28088,N_27963,N_27857);
and U28089 (N_28089,N_27930,N_27923);
or U28090 (N_28090,N_27931,N_27942);
and U28091 (N_28091,N_27905,N_27914);
nor U28092 (N_28092,N_27884,N_27920);
or U28093 (N_28093,N_27984,N_27849);
xnor U28094 (N_28094,N_27885,N_27853);
nor U28095 (N_28095,N_27895,N_27938);
or U28096 (N_28096,N_27822,N_27870);
xor U28097 (N_28097,N_27981,N_27824);
nor U28098 (N_28098,N_27939,N_27854);
and U28099 (N_28099,N_27940,N_27934);
and U28100 (N_28100,N_27860,N_27874);
or U28101 (N_28101,N_27814,N_27912);
nand U28102 (N_28102,N_27912,N_27950);
and U28103 (N_28103,N_27897,N_27928);
nor U28104 (N_28104,N_27988,N_27891);
and U28105 (N_28105,N_27952,N_27874);
or U28106 (N_28106,N_27936,N_27955);
nand U28107 (N_28107,N_27835,N_27879);
xor U28108 (N_28108,N_27910,N_27907);
xor U28109 (N_28109,N_27925,N_27853);
or U28110 (N_28110,N_27815,N_27807);
and U28111 (N_28111,N_27938,N_27805);
and U28112 (N_28112,N_27816,N_27868);
xnor U28113 (N_28113,N_27877,N_27881);
and U28114 (N_28114,N_27995,N_27828);
xor U28115 (N_28115,N_27829,N_27827);
nand U28116 (N_28116,N_27918,N_27839);
nand U28117 (N_28117,N_27943,N_27850);
nor U28118 (N_28118,N_27876,N_27914);
nand U28119 (N_28119,N_27975,N_27862);
nor U28120 (N_28120,N_27863,N_27962);
nand U28121 (N_28121,N_27949,N_27962);
or U28122 (N_28122,N_27959,N_27854);
nor U28123 (N_28123,N_27958,N_27948);
xor U28124 (N_28124,N_27974,N_27813);
nor U28125 (N_28125,N_27933,N_27846);
nor U28126 (N_28126,N_27823,N_27944);
nor U28127 (N_28127,N_27967,N_27825);
and U28128 (N_28128,N_27996,N_27822);
xor U28129 (N_28129,N_27851,N_27930);
and U28130 (N_28130,N_27941,N_27846);
nor U28131 (N_28131,N_27940,N_27918);
xor U28132 (N_28132,N_27851,N_27800);
nor U28133 (N_28133,N_27830,N_27947);
nand U28134 (N_28134,N_27826,N_27935);
and U28135 (N_28135,N_27926,N_27840);
nor U28136 (N_28136,N_27904,N_27871);
xnor U28137 (N_28137,N_27882,N_27917);
or U28138 (N_28138,N_27918,N_27867);
or U28139 (N_28139,N_27877,N_27880);
xnor U28140 (N_28140,N_27879,N_27917);
nand U28141 (N_28141,N_27967,N_27931);
nor U28142 (N_28142,N_27929,N_27927);
nor U28143 (N_28143,N_27969,N_27844);
nor U28144 (N_28144,N_27995,N_27821);
nand U28145 (N_28145,N_27996,N_27868);
or U28146 (N_28146,N_27943,N_27835);
or U28147 (N_28147,N_27962,N_27867);
xnor U28148 (N_28148,N_27832,N_27956);
xnor U28149 (N_28149,N_27924,N_27974);
and U28150 (N_28150,N_27988,N_27930);
xor U28151 (N_28151,N_27871,N_27882);
xnor U28152 (N_28152,N_27927,N_27944);
xor U28153 (N_28153,N_27998,N_27811);
nand U28154 (N_28154,N_27971,N_27934);
nand U28155 (N_28155,N_27807,N_27913);
nor U28156 (N_28156,N_27992,N_27938);
nand U28157 (N_28157,N_27998,N_27986);
nor U28158 (N_28158,N_27916,N_27999);
nor U28159 (N_28159,N_27931,N_27821);
nor U28160 (N_28160,N_27948,N_27864);
nand U28161 (N_28161,N_27882,N_27839);
nor U28162 (N_28162,N_27893,N_27967);
or U28163 (N_28163,N_27888,N_27928);
and U28164 (N_28164,N_27945,N_27851);
xor U28165 (N_28165,N_27951,N_27835);
and U28166 (N_28166,N_27925,N_27846);
nor U28167 (N_28167,N_27808,N_27892);
or U28168 (N_28168,N_27845,N_27930);
or U28169 (N_28169,N_27884,N_27875);
and U28170 (N_28170,N_27873,N_27968);
and U28171 (N_28171,N_27888,N_27960);
nand U28172 (N_28172,N_27908,N_27878);
nand U28173 (N_28173,N_27946,N_27906);
nor U28174 (N_28174,N_27910,N_27987);
nor U28175 (N_28175,N_27898,N_27940);
or U28176 (N_28176,N_27857,N_27964);
nand U28177 (N_28177,N_27900,N_27874);
xor U28178 (N_28178,N_27912,N_27886);
nor U28179 (N_28179,N_27990,N_27846);
nor U28180 (N_28180,N_27975,N_27855);
xnor U28181 (N_28181,N_27998,N_27889);
or U28182 (N_28182,N_27852,N_27963);
nor U28183 (N_28183,N_27976,N_27932);
or U28184 (N_28184,N_27957,N_27968);
nor U28185 (N_28185,N_27927,N_27945);
or U28186 (N_28186,N_27987,N_27894);
xor U28187 (N_28187,N_27827,N_27929);
and U28188 (N_28188,N_27977,N_27841);
or U28189 (N_28189,N_27820,N_27824);
and U28190 (N_28190,N_27968,N_27944);
xnor U28191 (N_28191,N_27954,N_27952);
nor U28192 (N_28192,N_27960,N_27818);
nand U28193 (N_28193,N_27955,N_27845);
or U28194 (N_28194,N_27886,N_27852);
nand U28195 (N_28195,N_27920,N_27871);
or U28196 (N_28196,N_27860,N_27899);
nand U28197 (N_28197,N_27979,N_27896);
or U28198 (N_28198,N_27998,N_27979);
and U28199 (N_28199,N_27905,N_27921);
or U28200 (N_28200,N_28116,N_28038);
and U28201 (N_28201,N_28189,N_28058);
xor U28202 (N_28202,N_28142,N_28123);
nand U28203 (N_28203,N_28013,N_28104);
or U28204 (N_28204,N_28089,N_28087);
nand U28205 (N_28205,N_28128,N_28059);
xnor U28206 (N_28206,N_28039,N_28101);
nand U28207 (N_28207,N_28082,N_28199);
nor U28208 (N_28208,N_28085,N_28044);
xnor U28209 (N_28209,N_28029,N_28164);
or U28210 (N_28210,N_28017,N_28004);
nand U28211 (N_28211,N_28131,N_28025);
nand U28212 (N_28212,N_28172,N_28096);
nand U28213 (N_28213,N_28130,N_28122);
xnor U28214 (N_28214,N_28095,N_28014);
and U28215 (N_28215,N_28046,N_28099);
nor U28216 (N_28216,N_28185,N_28158);
and U28217 (N_28217,N_28175,N_28153);
nor U28218 (N_28218,N_28077,N_28160);
or U28219 (N_28219,N_28019,N_28000);
nand U28220 (N_28220,N_28042,N_28031);
and U28221 (N_28221,N_28147,N_28148);
or U28222 (N_28222,N_28071,N_28156);
nand U28223 (N_28223,N_28075,N_28145);
xnor U28224 (N_28224,N_28047,N_28143);
nand U28225 (N_28225,N_28001,N_28008);
nand U28226 (N_28226,N_28024,N_28149);
nand U28227 (N_28227,N_28093,N_28045);
or U28228 (N_28228,N_28003,N_28057);
and U28229 (N_28229,N_28178,N_28124);
nor U28230 (N_28230,N_28090,N_28140);
or U28231 (N_28231,N_28197,N_28068);
and U28232 (N_28232,N_28177,N_28138);
or U28233 (N_28233,N_28028,N_28115);
and U28234 (N_28234,N_28152,N_28135);
or U28235 (N_28235,N_28016,N_28168);
and U28236 (N_28236,N_28170,N_28186);
nor U28237 (N_28237,N_28091,N_28195);
xor U28238 (N_28238,N_28133,N_28056);
xnor U28239 (N_28239,N_28173,N_28103);
nor U28240 (N_28240,N_28063,N_28150);
xnor U28241 (N_28241,N_28078,N_28171);
xnor U28242 (N_28242,N_28129,N_28165);
xor U28243 (N_28243,N_28176,N_28036);
nor U28244 (N_28244,N_28119,N_28105);
or U28245 (N_28245,N_28073,N_28196);
nor U28246 (N_28246,N_28106,N_28050);
nand U28247 (N_28247,N_28030,N_28136);
or U28248 (N_28248,N_28169,N_28184);
or U28249 (N_28249,N_28162,N_28102);
nand U28250 (N_28250,N_28084,N_28190);
xnor U28251 (N_28251,N_28067,N_28194);
and U28252 (N_28252,N_28098,N_28074);
and U28253 (N_28253,N_28188,N_28021);
xor U28254 (N_28254,N_28035,N_28009);
nand U28255 (N_28255,N_28180,N_28015);
nor U28256 (N_28256,N_28048,N_28097);
or U28257 (N_28257,N_28061,N_28183);
and U28258 (N_28258,N_28052,N_28043);
or U28259 (N_28259,N_28094,N_28144);
and U28260 (N_28260,N_28053,N_28134);
and U28261 (N_28261,N_28191,N_28033);
nor U28262 (N_28262,N_28146,N_28080);
nand U28263 (N_28263,N_28086,N_28088);
xor U28264 (N_28264,N_28081,N_28065);
xnor U28265 (N_28265,N_28002,N_28079);
or U28266 (N_28266,N_28040,N_28159);
nor U28267 (N_28267,N_28127,N_28010);
and U28268 (N_28268,N_28041,N_28198);
nand U28269 (N_28269,N_28167,N_28064);
nand U28270 (N_28270,N_28126,N_28114);
nand U28271 (N_28271,N_28166,N_28117);
xnor U28272 (N_28272,N_28026,N_28192);
nand U28273 (N_28273,N_28108,N_28023);
and U28274 (N_28274,N_28137,N_28069);
or U28275 (N_28275,N_28032,N_28151);
and U28276 (N_28276,N_28020,N_28049);
and U28277 (N_28277,N_28139,N_28112);
and U28278 (N_28278,N_28181,N_28161);
and U28279 (N_28279,N_28007,N_28154);
nand U28280 (N_28280,N_28006,N_28083);
nand U28281 (N_28281,N_28076,N_28011);
nand U28282 (N_28282,N_28155,N_28022);
and U28283 (N_28283,N_28110,N_28070);
nand U28284 (N_28284,N_28055,N_28060);
nand U28285 (N_28285,N_28187,N_28027);
xnor U28286 (N_28286,N_28121,N_28034);
nand U28287 (N_28287,N_28193,N_28005);
nor U28288 (N_28288,N_28018,N_28012);
nor U28289 (N_28289,N_28141,N_28066);
xnor U28290 (N_28290,N_28107,N_28051);
or U28291 (N_28291,N_28118,N_28157);
xnor U28292 (N_28292,N_28100,N_28092);
xor U28293 (N_28293,N_28174,N_28037);
nand U28294 (N_28294,N_28132,N_28062);
nand U28295 (N_28295,N_28054,N_28163);
xnor U28296 (N_28296,N_28109,N_28179);
nor U28297 (N_28297,N_28072,N_28125);
xnor U28298 (N_28298,N_28120,N_28111);
nor U28299 (N_28299,N_28113,N_28182);
nand U28300 (N_28300,N_28033,N_28184);
and U28301 (N_28301,N_28015,N_28034);
or U28302 (N_28302,N_28131,N_28111);
or U28303 (N_28303,N_28159,N_28126);
or U28304 (N_28304,N_28166,N_28027);
nor U28305 (N_28305,N_28034,N_28010);
and U28306 (N_28306,N_28094,N_28001);
nand U28307 (N_28307,N_28042,N_28071);
nand U28308 (N_28308,N_28120,N_28060);
nand U28309 (N_28309,N_28047,N_28063);
and U28310 (N_28310,N_28059,N_28143);
xnor U28311 (N_28311,N_28093,N_28169);
nand U28312 (N_28312,N_28005,N_28155);
nor U28313 (N_28313,N_28128,N_28110);
nand U28314 (N_28314,N_28009,N_28165);
nand U28315 (N_28315,N_28034,N_28198);
nor U28316 (N_28316,N_28136,N_28194);
or U28317 (N_28317,N_28013,N_28113);
nor U28318 (N_28318,N_28092,N_28166);
nor U28319 (N_28319,N_28156,N_28056);
nor U28320 (N_28320,N_28182,N_28108);
nor U28321 (N_28321,N_28073,N_28045);
xnor U28322 (N_28322,N_28190,N_28168);
and U28323 (N_28323,N_28157,N_28179);
and U28324 (N_28324,N_28167,N_28153);
xnor U28325 (N_28325,N_28162,N_28037);
or U28326 (N_28326,N_28049,N_28000);
xor U28327 (N_28327,N_28073,N_28066);
nor U28328 (N_28328,N_28111,N_28164);
nand U28329 (N_28329,N_28182,N_28082);
xnor U28330 (N_28330,N_28040,N_28156);
xor U28331 (N_28331,N_28166,N_28038);
and U28332 (N_28332,N_28156,N_28074);
nand U28333 (N_28333,N_28073,N_28103);
or U28334 (N_28334,N_28079,N_28136);
nor U28335 (N_28335,N_28071,N_28165);
nand U28336 (N_28336,N_28082,N_28124);
and U28337 (N_28337,N_28083,N_28097);
nand U28338 (N_28338,N_28188,N_28108);
nand U28339 (N_28339,N_28110,N_28061);
xor U28340 (N_28340,N_28086,N_28112);
nand U28341 (N_28341,N_28036,N_28067);
nor U28342 (N_28342,N_28031,N_28095);
nor U28343 (N_28343,N_28171,N_28130);
and U28344 (N_28344,N_28032,N_28074);
nand U28345 (N_28345,N_28160,N_28110);
nor U28346 (N_28346,N_28001,N_28027);
and U28347 (N_28347,N_28142,N_28185);
xnor U28348 (N_28348,N_28154,N_28039);
nor U28349 (N_28349,N_28105,N_28127);
and U28350 (N_28350,N_28162,N_28123);
and U28351 (N_28351,N_28060,N_28012);
xnor U28352 (N_28352,N_28053,N_28158);
xor U28353 (N_28353,N_28099,N_28109);
or U28354 (N_28354,N_28121,N_28013);
nor U28355 (N_28355,N_28066,N_28134);
xor U28356 (N_28356,N_28074,N_28020);
and U28357 (N_28357,N_28071,N_28079);
and U28358 (N_28358,N_28070,N_28130);
nand U28359 (N_28359,N_28166,N_28188);
or U28360 (N_28360,N_28080,N_28014);
nand U28361 (N_28361,N_28124,N_28113);
or U28362 (N_28362,N_28101,N_28059);
nor U28363 (N_28363,N_28190,N_28095);
xnor U28364 (N_28364,N_28181,N_28135);
nand U28365 (N_28365,N_28045,N_28161);
or U28366 (N_28366,N_28071,N_28159);
and U28367 (N_28367,N_28024,N_28094);
and U28368 (N_28368,N_28085,N_28128);
nand U28369 (N_28369,N_28140,N_28039);
nor U28370 (N_28370,N_28134,N_28150);
nand U28371 (N_28371,N_28001,N_28058);
nor U28372 (N_28372,N_28026,N_28001);
xor U28373 (N_28373,N_28067,N_28020);
nand U28374 (N_28374,N_28179,N_28162);
and U28375 (N_28375,N_28187,N_28103);
or U28376 (N_28376,N_28002,N_28144);
nand U28377 (N_28377,N_28138,N_28087);
or U28378 (N_28378,N_28004,N_28133);
nand U28379 (N_28379,N_28131,N_28097);
and U28380 (N_28380,N_28098,N_28028);
or U28381 (N_28381,N_28060,N_28058);
and U28382 (N_28382,N_28104,N_28139);
and U28383 (N_28383,N_28026,N_28114);
nand U28384 (N_28384,N_28123,N_28037);
nor U28385 (N_28385,N_28054,N_28036);
nor U28386 (N_28386,N_28079,N_28095);
nand U28387 (N_28387,N_28071,N_28109);
and U28388 (N_28388,N_28015,N_28041);
or U28389 (N_28389,N_28083,N_28095);
and U28390 (N_28390,N_28046,N_28097);
or U28391 (N_28391,N_28108,N_28164);
or U28392 (N_28392,N_28188,N_28020);
or U28393 (N_28393,N_28181,N_28005);
nor U28394 (N_28394,N_28052,N_28031);
and U28395 (N_28395,N_28172,N_28082);
xor U28396 (N_28396,N_28019,N_28098);
nor U28397 (N_28397,N_28039,N_28005);
xnor U28398 (N_28398,N_28067,N_28018);
nand U28399 (N_28399,N_28066,N_28191);
or U28400 (N_28400,N_28315,N_28380);
xor U28401 (N_28401,N_28239,N_28382);
or U28402 (N_28402,N_28200,N_28219);
nor U28403 (N_28403,N_28374,N_28360);
nor U28404 (N_28404,N_28362,N_28359);
and U28405 (N_28405,N_28307,N_28371);
or U28406 (N_28406,N_28384,N_28289);
nor U28407 (N_28407,N_28265,N_28397);
or U28408 (N_28408,N_28332,N_28310);
or U28409 (N_28409,N_28295,N_28211);
nor U28410 (N_28410,N_28346,N_28262);
or U28411 (N_28411,N_28368,N_28301);
xor U28412 (N_28412,N_28398,N_28372);
and U28413 (N_28413,N_28280,N_28340);
or U28414 (N_28414,N_28223,N_28285);
xor U28415 (N_28415,N_28251,N_28358);
or U28416 (N_28416,N_28271,N_28274);
and U28417 (N_28417,N_28287,N_28296);
or U28418 (N_28418,N_28353,N_28238);
xnor U28419 (N_28419,N_28344,N_28290);
or U28420 (N_28420,N_28351,N_28385);
nor U28421 (N_28421,N_28395,N_28329);
xor U28422 (N_28422,N_28378,N_28396);
xor U28423 (N_28423,N_28331,N_28347);
and U28424 (N_28424,N_28282,N_28240);
nor U28425 (N_28425,N_28230,N_28377);
nand U28426 (N_28426,N_28294,N_28297);
nor U28427 (N_28427,N_28335,N_28257);
or U28428 (N_28428,N_28369,N_28291);
and U28429 (N_28429,N_28204,N_28298);
nor U28430 (N_28430,N_28330,N_28221);
nor U28431 (N_28431,N_28392,N_28365);
nor U28432 (N_28432,N_28341,N_28356);
nor U28433 (N_28433,N_28319,N_28383);
or U28434 (N_28434,N_28387,N_28318);
or U28435 (N_28435,N_28316,N_28250);
or U28436 (N_28436,N_28393,N_28370);
and U28437 (N_28437,N_28373,N_28352);
or U28438 (N_28438,N_28212,N_28336);
nand U28439 (N_28439,N_28270,N_28308);
nand U28440 (N_28440,N_28390,N_28288);
or U28441 (N_28441,N_28225,N_28361);
and U28442 (N_28442,N_28348,N_28245);
or U28443 (N_28443,N_28333,N_28364);
and U28444 (N_28444,N_28216,N_28305);
or U28445 (N_28445,N_28252,N_28268);
xnor U28446 (N_28446,N_28350,N_28321);
xnor U28447 (N_28447,N_28339,N_28325);
or U28448 (N_28448,N_28363,N_28312);
and U28449 (N_28449,N_28338,N_28284);
nor U28450 (N_28450,N_28311,N_28201);
or U28451 (N_28451,N_28300,N_28391);
nand U28452 (N_28452,N_28234,N_28242);
nor U28453 (N_28453,N_28233,N_28334);
nor U28454 (N_28454,N_28281,N_28226);
or U28455 (N_28455,N_28229,N_28254);
nor U28456 (N_28456,N_28210,N_28209);
and U28457 (N_28457,N_28279,N_28255);
nand U28458 (N_28458,N_28215,N_28342);
nor U28459 (N_28459,N_28266,N_28306);
and U28460 (N_28460,N_28203,N_28241);
and U28461 (N_28461,N_28246,N_28206);
and U28462 (N_28462,N_28317,N_28232);
xor U28463 (N_28463,N_28324,N_28328);
nand U28464 (N_28464,N_28278,N_28337);
nor U28465 (N_28465,N_28237,N_28236);
nor U28466 (N_28466,N_28264,N_28228);
and U28467 (N_28467,N_28320,N_28304);
and U28468 (N_28468,N_28309,N_28343);
nor U28469 (N_28469,N_28244,N_28202);
or U28470 (N_28470,N_28256,N_28222);
nand U28471 (N_28471,N_28224,N_28214);
and U28472 (N_28472,N_28355,N_28302);
and U28473 (N_28473,N_28213,N_28269);
nand U28474 (N_28474,N_28272,N_28379);
nand U28475 (N_28475,N_28235,N_28231);
and U28476 (N_28476,N_28207,N_28313);
and U28477 (N_28477,N_28263,N_28205);
or U28478 (N_28478,N_28261,N_28322);
or U28479 (N_28479,N_28275,N_28345);
nor U28480 (N_28480,N_28354,N_28293);
nor U28481 (N_28481,N_28386,N_28248);
nand U28482 (N_28482,N_28367,N_28276);
or U28483 (N_28483,N_28220,N_28208);
xnor U28484 (N_28484,N_28277,N_28327);
or U28485 (N_28485,N_28389,N_28349);
and U28486 (N_28486,N_28303,N_28399);
and U28487 (N_28487,N_28249,N_28381);
nand U28488 (N_28488,N_28326,N_28314);
nand U28489 (N_28489,N_28323,N_28267);
nor U28490 (N_28490,N_28299,N_28357);
or U28491 (N_28491,N_28260,N_28286);
nand U28492 (N_28492,N_28218,N_28227);
nand U28493 (N_28493,N_28366,N_28247);
xnor U28494 (N_28494,N_28243,N_28217);
or U28495 (N_28495,N_28273,N_28258);
xor U28496 (N_28496,N_28253,N_28388);
or U28497 (N_28497,N_28283,N_28394);
and U28498 (N_28498,N_28292,N_28376);
xor U28499 (N_28499,N_28375,N_28259);
or U28500 (N_28500,N_28290,N_28214);
nand U28501 (N_28501,N_28380,N_28206);
nor U28502 (N_28502,N_28391,N_28226);
and U28503 (N_28503,N_28351,N_28271);
nand U28504 (N_28504,N_28344,N_28268);
or U28505 (N_28505,N_28298,N_28279);
nor U28506 (N_28506,N_28349,N_28342);
nand U28507 (N_28507,N_28350,N_28369);
or U28508 (N_28508,N_28265,N_28248);
or U28509 (N_28509,N_28209,N_28390);
and U28510 (N_28510,N_28327,N_28240);
xor U28511 (N_28511,N_28317,N_28221);
or U28512 (N_28512,N_28290,N_28319);
or U28513 (N_28513,N_28279,N_28285);
and U28514 (N_28514,N_28293,N_28315);
nor U28515 (N_28515,N_28249,N_28344);
nor U28516 (N_28516,N_28384,N_28259);
nor U28517 (N_28517,N_28397,N_28298);
xnor U28518 (N_28518,N_28302,N_28357);
xnor U28519 (N_28519,N_28268,N_28317);
nand U28520 (N_28520,N_28373,N_28225);
nand U28521 (N_28521,N_28347,N_28329);
and U28522 (N_28522,N_28288,N_28214);
nor U28523 (N_28523,N_28237,N_28201);
and U28524 (N_28524,N_28361,N_28275);
xor U28525 (N_28525,N_28341,N_28344);
nand U28526 (N_28526,N_28312,N_28369);
xnor U28527 (N_28527,N_28263,N_28257);
nand U28528 (N_28528,N_28266,N_28344);
xnor U28529 (N_28529,N_28373,N_28272);
or U28530 (N_28530,N_28233,N_28218);
or U28531 (N_28531,N_28371,N_28245);
nand U28532 (N_28532,N_28205,N_28304);
nor U28533 (N_28533,N_28260,N_28300);
nand U28534 (N_28534,N_28272,N_28225);
xnor U28535 (N_28535,N_28290,N_28217);
and U28536 (N_28536,N_28204,N_28312);
and U28537 (N_28537,N_28214,N_28349);
xnor U28538 (N_28538,N_28341,N_28238);
nand U28539 (N_28539,N_28342,N_28345);
xnor U28540 (N_28540,N_28354,N_28218);
xor U28541 (N_28541,N_28389,N_28274);
xor U28542 (N_28542,N_28215,N_28255);
xnor U28543 (N_28543,N_28354,N_28335);
nor U28544 (N_28544,N_28368,N_28360);
nor U28545 (N_28545,N_28387,N_28269);
and U28546 (N_28546,N_28269,N_28334);
nor U28547 (N_28547,N_28327,N_28351);
or U28548 (N_28548,N_28344,N_28289);
nand U28549 (N_28549,N_28306,N_28399);
nand U28550 (N_28550,N_28235,N_28358);
or U28551 (N_28551,N_28387,N_28259);
and U28552 (N_28552,N_28395,N_28363);
nand U28553 (N_28553,N_28396,N_28219);
xnor U28554 (N_28554,N_28391,N_28346);
and U28555 (N_28555,N_28245,N_28241);
nand U28556 (N_28556,N_28295,N_28346);
nand U28557 (N_28557,N_28301,N_28399);
nand U28558 (N_28558,N_28394,N_28273);
or U28559 (N_28559,N_28395,N_28232);
and U28560 (N_28560,N_28265,N_28273);
or U28561 (N_28561,N_28345,N_28334);
xor U28562 (N_28562,N_28236,N_28391);
nand U28563 (N_28563,N_28399,N_28361);
and U28564 (N_28564,N_28332,N_28250);
xnor U28565 (N_28565,N_28373,N_28252);
nand U28566 (N_28566,N_28203,N_28291);
nor U28567 (N_28567,N_28287,N_28290);
nand U28568 (N_28568,N_28324,N_28334);
or U28569 (N_28569,N_28390,N_28215);
xnor U28570 (N_28570,N_28287,N_28350);
nor U28571 (N_28571,N_28202,N_28306);
xnor U28572 (N_28572,N_28396,N_28295);
xor U28573 (N_28573,N_28342,N_28207);
and U28574 (N_28574,N_28341,N_28286);
nand U28575 (N_28575,N_28254,N_28341);
nor U28576 (N_28576,N_28298,N_28259);
nor U28577 (N_28577,N_28380,N_28243);
or U28578 (N_28578,N_28388,N_28227);
xnor U28579 (N_28579,N_28371,N_28312);
and U28580 (N_28580,N_28253,N_28281);
and U28581 (N_28581,N_28239,N_28211);
nand U28582 (N_28582,N_28213,N_28278);
or U28583 (N_28583,N_28201,N_28241);
or U28584 (N_28584,N_28234,N_28266);
and U28585 (N_28585,N_28202,N_28273);
nand U28586 (N_28586,N_28314,N_28387);
xnor U28587 (N_28587,N_28211,N_28349);
nor U28588 (N_28588,N_28346,N_28352);
nor U28589 (N_28589,N_28308,N_28357);
xnor U28590 (N_28590,N_28249,N_28379);
xor U28591 (N_28591,N_28330,N_28273);
and U28592 (N_28592,N_28258,N_28386);
nor U28593 (N_28593,N_28220,N_28216);
nand U28594 (N_28594,N_28380,N_28343);
xor U28595 (N_28595,N_28266,N_28206);
nand U28596 (N_28596,N_28242,N_28207);
and U28597 (N_28597,N_28280,N_28260);
or U28598 (N_28598,N_28223,N_28352);
and U28599 (N_28599,N_28328,N_28395);
and U28600 (N_28600,N_28439,N_28440);
xnor U28601 (N_28601,N_28422,N_28420);
or U28602 (N_28602,N_28451,N_28494);
or U28603 (N_28603,N_28578,N_28542);
nand U28604 (N_28604,N_28586,N_28412);
nand U28605 (N_28605,N_28414,N_28455);
and U28606 (N_28606,N_28558,N_28538);
and U28607 (N_28607,N_28549,N_28596);
nor U28608 (N_28608,N_28444,N_28530);
xor U28609 (N_28609,N_28453,N_28488);
nor U28610 (N_28610,N_28524,N_28561);
nand U28611 (N_28611,N_28571,N_28501);
nand U28612 (N_28612,N_28469,N_28423);
nand U28613 (N_28613,N_28511,N_28431);
xnor U28614 (N_28614,N_28417,N_28519);
nor U28615 (N_28615,N_28534,N_28435);
nor U28616 (N_28616,N_28574,N_28535);
and U28617 (N_28617,N_28406,N_28464);
nand U28618 (N_28618,N_28556,N_28427);
or U28619 (N_28619,N_28506,N_28466);
or U28620 (N_28620,N_28569,N_28479);
nand U28621 (N_28621,N_28443,N_28410);
or U28622 (N_28622,N_28470,N_28409);
nor U28623 (N_28623,N_28438,N_28539);
nand U28624 (N_28624,N_28487,N_28518);
or U28625 (N_28625,N_28485,N_28421);
or U28626 (N_28626,N_28523,N_28594);
nor U28627 (N_28627,N_28588,N_28573);
nand U28628 (N_28628,N_28411,N_28545);
or U28629 (N_28629,N_28541,N_28459);
xor U28630 (N_28630,N_28424,N_28521);
nand U28631 (N_28631,N_28575,N_28477);
nor U28632 (N_28632,N_28567,N_28447);
xor U28633 (N_28633,N_28563,N_28408);
xnor U28634 (N_28634,N_28413,N_28513);
or U28635 (N_28635,N_28515,N_28590);
xnor U28636 (N_28636,N_28456,N_28436);
nand U28637 (N_28637,N_28517,N_28445);
nor U28638 (N_28638,N_28531,N_28560);
or U28639 (N_28639,N_28512,N_28576);
or U28640 (N_28640,N_28581,N_28587);
and U28641 (N_28641,N_28449,N_28403);
or U28642 (N_28642,N_28441,N_28529);
xor U28643 (N_28643,N_28500,N_28498);
nand U28644 (N_28644,N_28527,N_28593);
and U28645 (N_28645,N_28565,N_28559);
xnor U28646 (N_28646,N_28507,N_28404);
or U28647 (N_28647,N_28543,N_28481);
nor U28648 (N_28648,N_28599,N_28598);
nand U28649 (N_28649,N_28509,N_28514);
xor U28650 (N_28650,N_28448,N_28546);
nor U28651 (N_28651,N_28533,N_28475);
nor U28652 (N_28652,N_28497,N_28551);
nor U28653 (N_28653,N_28589,N_28555);
xnor U28654 (N_28654,N_28493,N_28597);
nor U28655 (N_28655,N_28547,N_28568);
xor U28656 (N_28656,N_28572,N_28548);
xnor U28657 (N_28657,N_28483,N_28508);
or U28658 (N_28658,N_28595,N_28536);
nor U28659 (N_28659,N_28416,N_28580);
and U28660 (N_28660,N_28489,N_28401);
nor U28661 (N_28661,N_28502,N_28584);
xnor U28662 (N_28662,N_28503,N_28537);
and U28663 (N_28663,N_28442,N_28462);
xnor U28664 (N_28664,N_28592,N_28405);
and U28665 (N_28665,N_28591,N_28554);
xor U28666 (N_28666,N_28532,N_28525);
and U28667 (N_28667,N_28450,N_28471);
or U28668 (N_28668,N_28486,N_28496);
or U28669 (N_28669,N_28419,N_28474);
or U28670 (N_28670,N_28430,N_28577);
xnor U28671 (N_28671,N_28472,N_28426);
xor U28672 (N_28672,N_28553,N_28562);
xor U28673 (N_28673,N_28467,N_28458);
nand U28674 (N_28674,N_28484,N_28402);
xnor U28675 (N_28675,N_28566,N_28540);
or U28676 (N_28676,N_28415,N_28418);
xor U28677 (N_28677,N_28491,N_28570);
or U28678 (N_28678,N_28473,N_28550);
or U28679 (N_28679,N_28476,N_28454);
nor U28680 (N_28680,N_28460,N_28425);
nand U28681 (N_28681,N_28482,N_28407);
nand U28682 (N_28682,N_28505,N_28579);
nand U28683 (N_28683,N_28526,N_28495);
or U28684 (N_28684,N_28490,N_28457);
nor U28685 (N_28685,N_28429,N_28557);
and U28686 (N_28686,N_28552,N_28504);
xnor U28687 (N_28687,N_28585,N_28461);
xnor U28688 (N_28688,N_28434,N_28437);
nor U28689 (N_28689,N_28522,N_28582);
nand U28690 (N_28690,N_28428,N_28465);
nor U28691 (N_28691,N_28516,N_28480);
nor U28692 (N_28692,N_28478,N_28544);
or U28693 (N_28693,N_28520,N_28468);
xor U28694 (N_28694,N_28400,N_28463);
nor U28695 (N_28695,N_28446,N_28583);
or U28696 (N_28696,N_28499,N_28433);
nand U28697 (N_28697,N_28510,N_28528);
xor U28698 (N_28698,N_28452,N_28564);
or U28699 (N_28699,N_28492,N_28432);
xnor U28700 (N_28700,N_28452,N_28540);
xor U28701 (N_28701,N_28487,N_28483);
and U28702 (N_28702,N_28458,N_28412);
xnor U28703 (N_28703,N_28570,N_28414);
nand U28704 (N_28704,N_28422,N_28407);
and U28705 (N_28705,N_28564,N_28430);
nor U28706 (N_28706,N_28571,N_28507);
and U28707 (N_28707,N_28547,N_28448);
and U28708 (N_28708,N_28520,N_28444);
and U28709 (N_28709,N_28417,N_28459);
nor U28710 (N_28710,N_28453,N_28589);
xor U28711 (N_28711,N_28558,N_28489);
nor U28712 (N_28712,N_28509,N_28504);
xnor U28713 (N_28713,N_28448,N_28414);
and U28714 (N_28714,N_28562,N_28485);
or U28715 (N_28715,N_28494,N_28543);
and U28716 (N_28716,N_28446,N_28440);
or U28717 (N_28717,N_28465,N_28517);
nand U28718 (N_28718,N_28592,N_28553);
or U28719 (N_28719,N_28525,N_28550);
nor U28720 (N_28720,N_28430,N_28583);
nand U28721 (N_28721,N_28435,N_28409);
nor U28722 (N_28722,N_28582,N_28484);
xnor U28723 (N_28723,N_28496,N_28562);
xor U28724 (N_28724,N_28462,N_28592);
nand U28725 (N_28725,N_28522,N_28590);
and U28726 (N_28726,N_28433,N_28594);
and U28727 (N_28727,N_28519,N_28445);
and U28728 (N_28728,N_28448,N_28594);
xor U28729 (N_28729,N_28511,N_28570);
nand U28730 (N_28730,N_28410,N_28457);
or U28731 (N_28731,N_28457,N_28572);
or U28732 (N_28732,N_28416,N_28527);
or U28733 (N_28733,N_28455,N_28412);
nor U28734 (N_28734,N_28483,N_28447);
xor U28735 (N_28735,N_28410,N_28560);
or U28736 (N_28736,N_28569,N_28587);
nor U28737 (N_28737,N_28512,N_28566);
xnor U28738 (N_28738,N_28473,N_28533);
nand U28739 (N_28739,N_28451,N_28575);
or U28740 (N_28740,N_28575,N_28550);
nor U28741 (N_28741,N_28475,N_28573);
nor U28742 (N_28742,N_28517,N_28475);
and U28743 (N_28743,N_28528,N_28566);
or U28744 (N_28744,N_28549,N_28401);
or U28745 (N_28745,N_28471,N_28439);
nand U28746 (N_28746,N_28569,N_28514);
and U28747 (N_28747,N_28417,N_28548);
xnor U28748 (N_28748,N_28435,N_28463);
nor U28749 (N_28749,N_28547,N_28559);
nor U28750 (N_28750,N_28430,N_28478);
and U28751 (N_28751,N_28513,N_28468);
xor U28752 (N_28752,N_28462,N_28491);
and U28753 (N_28753,N_28583,N_28482);
xnor U28754 (N_28754,N_28462,N_28565);
or U28755 (N_28755,N_28446,N_28462);
or U28756 (N_28756,N_28498,N_28538);
or U28757 (N_28757,N_28494,N_28542);
or U28758 (N_28758,N_28524,N_28447);
nor U28759 (N_28759,N_28467,N_28428);
xor U28760 (N_28760,N_28568,N_28446);
xnor U28761 (N_28761,N_28452,N_28544);
nor U28762 (N_28762,N_28573,N_28538);
and U28763 (N_28763,N_28530,N_28460);
xnor U28764 (N_28764,N_28573,N_28519);
and U28765 (N_28765,N_28414,N_28537);
or U28766 (N_28766,N_28565,N_28539);
and U28767 (N_28767,N_28488,N_28467);
nand U28768 (N_28768,N_28412,N_28404);
xnor U28769 (N_28769,N_28598,N_28512);
and U28770 (N_28770,N_28530,N_28485);
or U28771 (N_28771,N_28437,N_28512);
nand U28772 (N_28772,N_28502,N_28401);
or U28773 (N_28773,N_28480,N_28402);
xor U28774 (N_28774,N_28444,N_28572);
and U28775 (N_28775,N_28574,N_28550);
or U28776 (N_28776,N_28513,N_28526);
and U28777 (N_28777,N_28484,N_28423);
or U28778 (N_28778,N_28595,N_28512);
nand U28779 (N_28779,N_28553,N_28461);
nor U28780 (N_28780,N_28574,N_28542);
nor U28781 (N_28781,N_28582,N_28432);
nand U28782 (N_28782,N_28495,N_28556);
nand U28783 (N_28783,N_28589,N_28445);
xor U28784 (N_28784,N_28508,N_28455);
nand U28785 (N_28785,N_28437,N_28449);
xnor U28786 (N_28786,N_28507,N_28498);
xnor U28787 (N_28787,N_28472,N_28539);
and U28788 (N_28788,N_28407,N_28487);
nand U28789 (N_28789,N_28451,N_28568);
xnor U28790 (N_28790,N_28446,N_28567);
nor U28791 (N_28791,N_28547,N_28433);
and U28792 (N_28792,N_28575,N_28440);
xor U28793 (N_28793,N_28479,N_28539);
or U28794 (N_28794,N_28486,N_28552);
or U28795 (N_28795,N_28537,N_28422);
and U28796 (N_28796,N_28589,N_28411);
xor U28797 (N_28797,N_28530,N_28423);
nor U28798 (N_28798,N_28517,N_28508);
and U28799 (N_28799,N_28545,N_28514);
or U28800 (N_28800,N_28795,N_28617);
and U28801 (N_28801,N_28637,N_28621);
or U28802 (N_28802,N_28790,N_28748);
and U28803 (N_28803,N_28650,N_28709);
xor U28804 (N_28804,N_28777,N_28623);
or U28805 (N_28805,N_28604,N_28679);
xor U28806 (N_28806,N_28766,N_28715);
xnor U28807 (N_28807,N_28780,N_28734);
and U28808 (N_28808,N_28611,N_28770);
nand U28809 (N_28809,N_28671,N_28642);
xor U28810 (N_28810,N_28602,N_28782);
xnor U28811 (N_28811,N_28733,N_28784);
nor U28812 (N_28812,N_28614,N_28746);
or U28813 (N_28813,N_28740,N_28719);
nor U28814 (N_28814,N_28720,N_28696);
xor U28815 (N_28815,N_28764,N_28705);
or U28816 (N_28816,N_28796,N_28665);
nor U28817 (N_28817,N_28672,N_28669);
and U28818 (N_28818,N_28693,N_28613);
or U28819 (N_28819,N_28789,N_28749);
or U28820 (N_28820,N_28760,N_28646);
xnor U28821 (N_28821,N_28666,N_28683);
or U28822 (N_28822,N_28622,N_28771);
or U28823 (N_28823,N_28668,N_28767);
and U28824 (N_28824,N_28688,N_28768);
and U28825 (N_28825,N_28639,N_28712);
and U28826 (N_28826,N_28702,N_28649);
xnor U28827 (N_28827,N_28730,N_28644);
and U28828 (N_28828,N_28792,N_28676);
or U28829 (N_28829,N_28655,N_28721);
nand U28830 (N_28830,N_28663,N_28739);
nor U28831 (N_28831,N_28778,N_28774);
or U28832 (N_28832,N_28675,N_28660);
and U28833 (N_28833,N_28707,N_28605);
and U28834 (N_28834,N_28747,N_28603);
or U28835 (N_28835,N_28634,N_28610);
nand U28836 (N_28836,N_28692,N_28785);
and U28837 (N_28837,N_28742,N_28791);
and U28838 (N_28838,N_28787,N_28744);
or U28839 (N_28839,N_28697,N_28689);
nand U28840 (N_28840,N_28643,N_28648);
or U28841 (N_28841,N_28727,N_28662);
nor U28842 (N_28842,N_28761,N_28640);
and U28843 (N_28843,N_28651,N_28633);
nand U28844 (N_28844,N_28752,N_28684);
and U28845 (N_28845,N_28619,N_28728);
nor U28846 (N_28846,N_28670,N_28708);
nand U28847 (N_28847,N_28735,N_28714);
and U28848 (N_28848,N_28797,N_28608);
and U28849 (N_28849,N_28754,N_28731);
nand U28850 (N_28850,N_28741,N_28772);
or U28851 (N_28851,N_28677,N_28658);
xor U28852 (N_28852,N_28723,N_28757);
and U28853 (N_28853,N_28703,N_28762);
nand U28854 (N_28854,N_28638,N_28691);
and U28855 (N_28855,N_28701,N_28654);
nand U28856 (N_28856,N_28680,N_28729);
xor U28857 (N_28857,N_28626,N_28636);
and U28858 (N_28858,N_28758,N_28745);
xnor U28859 (N_28859,N_28716,N_28620);
nand U28860 (N_28860,N_28694,N_28710);
and U28861 (N_28861,N_28681,N_28738);
or U28862 (N_28862,N_28687,N_28600);
and U28863 (N_28863,N_28601,N_28632);
xor U28864 (N_28864,N_28664,N_28732);
and U28865 (N_28865,N_28661,N_28713);
nand U28866 (N_28866,N_28765,N_28773);
nand U28867 (N_28867,N_28775,N_28783);
or U28868 (N_28868,N_28674,N_28612);
and U28869 (N_28869,N_28625,N_28667);
nor U28870 (N_28870,N_28704,N_28779);
xor U28871 (N_28871,N_28627,N_28695);
or U28872 (N_28872,N_28641,N_28652);
xor U28873 (N_28873,N_28781,N_28717);
nand U28874 (N_28874,N_28615,N_28635);
nand U28875 (N_28875,N_28616,N_28678);
and U28876 (N_28876,N_28724,N_28685);
and U28877 (N_28877,N_28763,N_28743);
nand U28878 (N_28878,N_28759,N_28794);
or U28879 (N_28879,N_28618,N_28786);
nor U28880 (N_28880,N_28799,N_28645);
nand U28881 (N_28881,N_28659,N_28653);
nand U28882 (N_28882,N_28699,N_28751);
xor U28883 (N_28883,N_28722,N_28656);
xor U28884 (N_28884,N_28756,N_28769);
nand U28885 (N_28885,N_28686,N_28628);
and U28886 (N_28886,N_28682,N_28631);
nand U28887 (N_28887,N_28609,N_28698);
xnor U28888 (N_28888,N_28793,N_28750);
or U28889 (N_28889,N_28753,N_28606);
nor U28890 (N_28890,N_28736,N_28673);
and U28891 (N_28891,N_28718,N_28607);
and U28892 (N_28892,N_28647,N_28706);
or U28893 (N_28893,N_28737,N_28788);
xnor U28894 (N_28894,N_28726,N_28690);
xnor U28895 (N_28895,N_28798,N_28700);
nor U28896 (N_28896,N_28657,N_28711);
nor U28897 (N_28897,N_28630,N_28624);
nand U28898 (N_28898,N_28629,N_28755);
and U28899 (N_28899,N_28776,N_28725);
xnor U28900 (N_28900,N_28648,N_28611);
or U28901 (N_28901,N_28606,N_28651);
or U28902 (N_28902,N_28600,N_28689);
or U28903 (N_28903,N_28661,N_28759);
or U28904 (N_28904,N_28700,N_28693);
or U28905 (N_28905,N_28749,N_28651);
nand U28906 (N_28906,N_28615,N_28634);
nor U28907 (N_28907,N_28668,N_28757);
or U28908 (N_28908,N_28777,N_28787);
or U28909 (N_28909,N_28676,N_28619);
nand U28910 (N_28910,N_28683,N_28749);
or U28911 (N_28911,N_28718,N_28683);
nor U28912 (N_28912,N_28764,N_28610);
nand U28913 (N_28913,N_28658,N_28793);
nor U28914 (N_28914,N_28707,N_28607);
and U28915 (N_28915,N_28777,N_28665);
xor U28916 (N_28916,N_28797,N_28620);
or U28917 (N_28917,N_28625,N_28715);
or U28918 (N_28918,N_28707,N_28783);
or U28919 (N_28919,N_28745,N_28738);
or U28920 (N_28920,N_28696,N_28651);
nand U28921 (N_28921,N_28633,N_28629);
and U28922 (N_28922,N_28642,N_28647);
or U28923 (N_28923,N_28712,N_28624);
nor U28924 (N_28924,N_28616,N_28762);
or U28925 (N_28925,N_28666,N_28684);
and U28926 (N_28926,N_28646,N_28638);
and U28927 (N_28927,N_28740,N_28763);
and U28928 (N_28928,N_28715,N_28757);
xnor U28929 (N_28929,N_28683,N_28676);
nand U28930 (N_28930,N_28748,N_28634);
nand U28931 (N_28931,N_28673,N_28632);
xnor U28932 (N_28932,N_28632,N_28741);
xnor U28933 (N_28933,N_28630,N_28790);
and U28934 (N_28934,N_28616,N_28777);
nand U28935 (N_28935,N_28682,N_28723);
and U28936 (N_28936,N_28762,N_28781);
xnor U28937 (N_28937,N_28727,N_28626);
or U28938 (N_28938,N_28724,N_28618);
nor U28939 (N_28939,N_28609,N_28761);
and U28940 (N_28940,N_28792,N_28759);
or U28941 (N_28941,N_28736,N_28687);
nand U28942 (N_28942,N_28771,N_28746);
nand U28943 (N_28943,N_28628,N_28726);
or U28944 (N_28944,N_28643,N_28732);
nor U28945 (N_28945,N_28658,N_28645);
xnor U28946 (N_28946,N_28798,N_28718);
nand U28947 (N_28947,N_28773,N_28767);
nor U28948 (N_28948,N_28781,N_28625);
and U28949 (N_28949,N_28659,N_28642);
xnor U28950 (N_28950,N_28704,N_28644);
xnor U28951 (N_28951,N_28619,N_28763);
and U28952 (N_28952,N_28654,N_28648);
or U28953 (N_28953,N_28727,N_28678);
or U28954 (N_28954,N_28666,N_28621);
or U28955 (N_28955,N_28735,N_28797);
xnor U28956 (N_28956,N_28700,N_28710);
nor U28957 (N_28957,N_28677,N_28700);
nand U28958 (N_28958,N_28603,N_28743);
and U28959 (N_28959,N_28699,N_28655);
xor U28960 (N_28960,N_28653,N_28642);
nor U28961 (N_28961,N_28660,N_28776);
and U28962 (N_28962,N_28784,N_28712);
nor U28963 (N_28963,N_28693,N_28676);
nand U28964 (N_28964,N_28646,N_28673);
nor U28965 (N_28965,N_28657,N_28632);
nor U28966 (N_28966,N_28744,N_28607);
or U28967 (N_28967,N_28694,N_28657);
xnor U28968 (N_28968,N_28682,N_28784);
nand U28969 (N_28969,N_28628,N_28747);
nand U28970 (N_28970,N_28637,N_28715);
nor U28971 (N_28971,N_28674,N_28756);
nand U28972 (N_28972,N_28725,N_28661);
or U28973 (N_28973,N_28718,N_28645);
or U28974 (N_28974,N_28771,N_28640);
and U28975 (N_28975,N_28679,N_28744);
xor U28976 (N_28976,N_28632,N_28788);
nand U28977 (N_28977,N_28615,N_28799);
nor U28978 (N_28978,N_28727,N_28758);
nand U28979 (N_28979,N_28679,N_28799);
nor U28980 (N_28980,N_28623,N_28738);
and U28981 (N_28981,N_28674,N_28730);
or U28982 (N_28982,N_28755,N_28611);
nor U28983 (N_28983,N_28713,N_28729);
or U28984 (N_28984,N_28629,N_28616);
nor U28985 (N_28985,N_28733,N_28659);
xor U28986 (N_28986,N_28651,N_28637);
nand U28987 (N_28987,N_28608,N_28633);
nand U28988 (N_28988,N_28612,N_28642);
nand U28989 (N_28989,N_28748,N_28683);
xnor U28990 (N_28990,N_28746,N_28789);
nand U28991 (N_28991,N_28633,N_28721);
or U28992 (N_28992,N_28699,N_28723);
nor U28993 (N_28993,N_28643,N_28698);
xnor U28994 (N_28994,N_28609,N_28652);
and U28995 (N_28995,N_28631,N_28610);
or U28996 (N_28996,N_28783,N_28634);
xnor U28997 (N_28997,N_28619,N_28780);
or U28998 (N_28998,N_28761,N_28651);
and U28999 (N_28999,N_28711,N_28778);
and U29000 (N_29000,N_28959,N_28973);
nand U29001 (N_29001,N_28811,N_28995);
nand U29002 (N_29002,N_28933,N_28827);
nor U29003 (N_29003,N_28996,N_28856);
nor U29004 (N_29004,N_28805,N_28999);
nand U29005 (N_29005,N_28822,N_28879);
nor U29006 (N_29006,N_28828,N_28867);
nand U29007 (N_29007,N_28939,N_28887);
xnor U29008 (N_29008,N_28945,N_28894);
and U29009 (N_29009,N_28936,N_28941);
nor U29010 (N_29010,N_28870,N_28962);
nor U29011 (N_29011,N_28892,N_28967);
and U29012 (N_29012,N_28881,N_28917);
nand U29013 (N_29013,N_28970,N_28952);
nand U29014 (N_29014,N_28864,N_28880);
nand U29015 (N_29015,N_28985,N_28833);
nor U29016 (N_29016,N_28874,N_28901);
and U29017 (N_29017,N_28947,N_28853);
xnor U29018 (N_29018,N_28969,N_28807);
xor U29019 (N_29019,N_28826,N_28857);
and U29020 (N_29020,N_28940,N_28845);
nor U29021 (N_29021,N_28992,N_28994);
nand U29022 (N_29022,N_28860,N_28974);
and U29023 (N_29023,N_28844,N_28871);
and U29024 (N_29024,N_28913,N_28835);
xnor U29025 (N_29025,N_28953,N_28937);
and U29026 (N_29026,N_28868,N_28926);
nand U29027 (N_29027,N_28821,N_28841);
nor U29028 (N_29028,N_28989,N_28893);
nor U29029 (N_29029,N_28902,N_28804);
and U29030 (N_29030,N_28801,N_28924);
or U29031 (N_29031,N_28922,N_28943);
or U29032 (N_29032,N_28961,N_28908);
nand U29033 (N_29033,N_28912,N_28850);
xor U29034 (N_29034,N_28808,N_28965);
nor U29035 (N_29035,N_28983,N_28981);
nor U29036 (N_29036,N_28907,N_28971);
and U29037 (N_29037,N_28858,N_28998);
xnor U29038 (N_29038,N_28921,N_28928);
xor U29039 (N_29039,N_28800,N_28956);
nor U29040 (N_29040,N_28877,N_28823);
nand U29041 (N_29041,N_28869,N_28975);
nor U29042 (N_29042,N_28852,N_28839);
or U29043 (N_29043,N_28919,N_28979);
and U29044 (N_29044,N_28882,N_28863);
nand U29045 (N_29045,N_28829,N_28990);
nor U29046 (N_29046,N_28909,N_28972);
or U29047 (N_29047,N_28842,N_28813);
xor U29048 (N_29048,N_28840,N_28817);
xnor U29049 (N_29049,N_28923,N_28873);
xor U29050 (N_29050,N_28897,N_28889);
and U29051 (N_29051,N_28914,N_28866);
xor U29052 (N_29052,N_28906,N_28825);
and U29053 (N_29053,N_28946,N_28944);
nand U29054 (N_29054,N_28930,N_28831);
or U29055 (N_29055,N_28883,N_28949);
nand U29056 (N_29056,N_28925,N_28814);
xor U29057 (N_29057,N_28886,N_28935);
and U29058 (N_29058,N_28855,N_28832);
and U29059 (N_29059,N_28927,N_28932);
xnor U29060 (N_29060,N_28984,N_28891);
nand U29061 (N_29061,N_28875,N_28824);
or U29062 (N_29062,N_28951,N_28895);
and U29063 (N_29063,N_28978,N_28898);
nor U29064 (N_29064,N_28819,N_28888);
and U29065 (N_29065,N_28899,N_28818);
xor U29066 (N_29066,N_28834,N_28903);
nor U29067 (N_29067,N_28938,N_28896);
nand U29068 (N_29068,N_28987,N_28900);
xnor U29069 (N_29069,N_28986,N_28865);
or U29070 (N_29070,N_28843,N_28918);
or U29071 (N_29071,N_28812,N_28963);
xor U29072 (N_29072,N_28916,N_28997);
xnor U29073 (N_29073,N_28810,N_28876);
and U29074 (N_29074,N_28872,N_28960);
and U29075 (N_29075,N_28934,N_28830);
nor U29076 (N_29076,N_28851,N_28929);
nor U29077 (N_29077,N_28890,N_28920);
or U29078 (N_29078,N_28803,N_28809);
or U29079 (N_29079,N_28976,N_28957);
nor U29080 (N_29080,N_28982,N_28878);
xor U29081 (N_29081,N_28968,N_28848);
and U29082 (N_29082,N_28942,N_28910);
nor U29083 (N_29083,N_28993,N_28904);
xnor U29084 (N_29084,N_28980,N_28905);
nand U29085 (N_29085,N_28991,N_28862);
or U29086 (N_29086,N_28948,N_28849);
nand U29087 (N_29087,N_28964,N_28958);
and U29088 (N_29088,N_28838,N_28816);
nand U29089 (N_29089,N_28988,N_28911);
or U29090 (N_29090,N_28859,N_28847);
and U29091 (N_29091,N_28854,N_28806);
or U29092 (N_29092,N_28861,N_28815);
or U29093 (N_29093,N_28837,N_28955);
or U29094 (N_29094,N_28884,N_28977);
xnor U29095 (N_29095,N_28966,N_28915);
nand U29096 (N_29096,N_28820,N_28950);
and U29097 (N_29097,N_28836,N_28931);
and U29098 (N_29098,N_28802,N_28954);
xnor U29099 (N_29099,N_28885,N_28846);
nand U29100 (N_29100,N_28876,N_28995);
nand U29101 (N_29101,N_28911,N_28883);
xor U29102 (N_29102,N_28874,N_28867);
xor U29103 (N_29103,N_28882,N_28857);
and U29104 (N_29104,N_28834,N_28906);
xnor U29105 (N_29105,N_28942,N_28815);
and U29106 (N_29106,N_28824,N_28898);
nand U29107 (N_29107,N_28961,N_28974);
xnor U29108 (N_29108,N_28844,N_28885);
nand U29109 (N_29109,N_28923,N_28837);
nor U29110 (N_29110,N_28939,N_28882);
xnor U29111 (N_29111,N_28945,N_28954);
nor U29112 (N_29112,N_28963,N_28939);
nor U29113 (N_29113,N_28877,N_28957);
and U29114 (N_29114,N_28865,N_28867);
xor U29115 (N_29115,N_28875,N_28998);
and U29116 (N_29116,N_28862,N_28954);
nand U29117 (N_29117,N_28906,N_28895);
or U29118 (N_29118,N_28828,N_28891);
xor U29119 (N_29119,N_28883,N_28836);
nor U29120 (N_29120,N_28923,N_28972);
and U29121 (N_29121,N_28853,N_28884);
nand U29122 (N_29122,N_28897,N_28890);
nor U29123 (N_29123,N_28834,N_28846);
nand U29124 (N_29124,N_28947,N_28858);
nand U29125 (N_29125,N_28881,N_28836);
nor U29126 (N_29126,N_28946,N_28960);
nand U29127 (N_29127,N_28902,N_28903);
xnor U29128 (N_29128,N_28951,N_28905);
and U29129 (N_29129,N_28819,N_28856);
and U29130 (N_29130,N_28944,N_28970);
and U29131 (N_29131,N_28929,N_28871);
and U29132 (N_29132,N_28961,N_28835);
and U29133 (N_29133,N_28896,N_28969);
or U29134 (N_29134,N_28980,N_28880);
nor U29135 (N_29135,N_28822,N_28928);
nor U29136 (N_29136,N_28983,N_28957);
nand U29137 (N_29137,N_28908,N_28913);
xor U29138 (N_29138,N_28888,N_28922);
nor U29139 (N_29139,N_28974,N_28949);
nand U29140 (N_29140,N_28963,N_28871);
nand U29141 (N_29141,N_28850,N_28853);
xor U29142 (N_29142,N_28909,N_28989);
nand U29143 (N_29143,N_28925,N_28923);
nor U29144 (N_29144,N_28933,N_28831);
nand U29145 (N_29145,N_28818,N_28982);
nor U29146 (N_29146,N_28839,N_28871);
xor U29147 (N_29147,N_28870,N_28826);
nor U29148 (N_29148,N_28898,N_28998);
and U29149 (N_29149,N_28920,N_28983);
or U29150 (N_29150,N_28914,N_28926);
or U29151 (N_29151,N_28804,N_28933);
nor U29152 (N_29152,N_28866,N_28935);
and U29153 (N_29153,N_28838,N_28854);
xnor U29154 (N_29154,N_28905,N_28936);
nand U29155 (N_29155,N_28823,N_28809);
and U29156 (N_29156,N_28990,N_28918);
nand U29157 (N_29157,N_28813,N_28876);
xor U29158 (N_29158,N_28959,N_28859);
xor U29159 (N_29159,N_28937,N_28913);
xnor U29160 (N_29160,N_28844,N_28939);
nor U29161 (N_29161,N_28859,N_28851);
nor U29162 (N_29162,N_28944,N_28805);
nor U29163 (N_29163,N_28879,N_28823);
and U29164 (N_29164,N_28867,N_28839);
xnor U29165 (N_29165,N_28989,N_28824);
and U29166 (N_29166,N_28867,N_28957);
nor U29167 (N_29167,N_28972,N_28843);
nor U29168 (N_29168,N_28822,N_28859);
nand U29169 (N_29169,N_28874,N_28914);
xor U29170 (N_29170,N_28957,N_28879);
and U29171 (N_29171,N_28840,N_28889);
xnor U29172 (N_29172,N_28977,N_28865);
xnor U29173 (N_29173,N_28895,N_28876);
and U29174 (N_29174,N_28812,N_28880);
or U29175 (N_29175,N_28930,N_28953);
or U29176 (N_29176,N_28974,N_28840);
xor U29177 (N_29177,N_28890,N_28861);
nand U29178 (N_29178,N_28829,N_28957);
and U29179 (N_29179,N_28906,N_28946);
xnor U29180 (N_29180,N_28819,N_28806);
xnor U29181 (N_29181,N_28857,N_28956);
nor U29182 (N_29182,N_28846,N_28961);
xor U29183 (N_29183,N_28848,N_28962);
or U29184 (N_29184,N_28905,N_28946);
xnor U29185 (N_29185,N_28840,N_28994);
nand U29186 (N_29186,N_28913,N_28931);
nand U29187 (N_29187,N_28954,N_28864);
nor U29188 (N_29188,N_28926,N_28814);
nand U29189 (N_29189,N_28947,N_28812);
nand U29190 (N_29190,N_28866,N_28822);
nor U29191 (N_29191,N_28883,N_28978);
and U29192 (N_29192,N_28814,N_28859);
nand U29193 (N_29193,N_28826,N_28853);
nand U29194 (N_29194,N_28891,N_28801);
nor U29195 (N_29195,N_28973,N_28864);
nand U29196 (N_29196,N_28898,N_28919);
nor U29197 (N_29197,N_28966,N_28840);
xnor U29198 (N_29198,N_28894,N_28863);
nor U29199 (N_29199,N_28983,N_28826);
or U29200 (N_29200,N_29115,N_29079);
nand U29201 (N_29201,N_29144,N_29007);
or U29202 (N_29202,N_29005,N_29122);
xor U29203 (N_29203,N_29163,N_29178);
nor U29204 (N_29204,N_29128,N_29106);
and U29205 (N_29205,N_29065,N_29154);
and U29206 (N_29206,N_29158,N_29093);
and U29207 (N_29207,N_29074,N_29137);
nor U29208 (N_29208,N_29130,N_29001);
nor U29209 (N_29209,N_29120,N_29190);
nand U29210 (N_29210,N_29043,N_29057);
and U29211 (N_29211,N_29058,N_29047);
or U29212 (N_29212,N_29103,N_29126);
nor U29213 (N_29213,N_29002,N_29070);
or U29214 (N_29214,N_29037,N_29036);
or U29215 (N_29215,N_29114,N_29022);
or U29216 (N_29216,N_29033,N_29098);
xor U29217 (N_29217,N_29135,N_29092);
nor U29218 (N_29218,N_29134,N_29041);
nor U29219 (N_29219,N_29066,N_29083);
nor U29220 (N_29220,N_29054,N_29145);
nand U29221 (N_29221,N_29010,N_29089);
nand U29222 (N_29222,N_29131,N_29182);
nor U29223 (N_29223,N_29040,N_29188);
xnor U29224 (N_29224,N_29169,N_29082);
xor U29225 (N_29225,N_29111,N_29044);
and U29226 (N_29226,N_29081,N_29003);
nor U29227 (N_29227,N_29029,N_29095);
and U29228 (N_29228,N_29147,N_29053);
nand U29229 (N_29229,N_29170,N_29011);
or U29230 (N_29230,N_29113,N_29026);
and U29231 (N_29231,N_29195,N_29105);
nor U29232 (N_29232,N_29028,N_29175);
nor U29233 (N_29233,N_29075,N_29097);
xor U29234 (N_29234,N_29140,N_29156);
nor U29235 (N_29235,N_29031,N_29121);
nor U29236 (N_29236,N_29123,N_29024);
and U29237 (N_29237,N_29038,N_29072);
xor U29238 (N_29238,N_29149,N_29157);
xor U29239 (N_29239,N_29067,N_29160);
nor U29240 (N_29240,N_29166,N_29050);
and U29241 (N_29241,N_29185,N_29060);
nor U29242 (N_29242,N_29167,N_29018);
and U29243 (N_29243,N_29080,N_29136);
and U29244 (N_29244,N_29193,N_29168);
xor U29245 (N_29245,N_29000,N_29143);
xnor U29246 (N_29246,N_29153,N_29014);
and U29247 (N_29247,N_29129,N_29174);
nor U29248 (N_29248,N_29189,N_29090);
and U29249 (N_29249,N_29159,N_29025);
or U29250 (N_29250,N_29187,N_29078);
and U29251 (N_29251,N_29164,N_29198);
or U29252 (N_29252,N_29071,N_29116);
and U29253 (N_29253,N_29104,N_29096);
or U29254 (N_29254,N_29165,N_29196);
nor U29255 (N_29255,N_29112,N_29194);
nand U29256 (N_29256,N_29012,N_29176);
and U29257 (N_29257,N_29117,N_29046);
and U29258 (N_29258,N_29049,N_29177);
or U29259 (N_29259,N_29184,N_29133);
nor U29260 (N_29260,N_29077,N_29086);
nand U29261 (N_29261,N_29102,N_29155);
or U29262 (N_29262,N_29192,N_29042);
nor U29263 (N_29263,N_29199,N_29191);
nand U29264 (N_29264,N_29125,N_29052);
nand U29265 (N_29265,N_29013,N_29100);
nor U29266 (N_29266,N_29076,N_29055);
xor U29267 (N_29267,N_29179,N_29063);
and U29268 (N_29268,N_29146,N_29032);
and U29269 (N_29269,N_29056,N_29019);
nor U29270 (N_29270,N_29048,N_29020);
and U29271 (N_29271,N_29017,N_29101);
and U29272 (N_29272,N_29108,N_29087);
nand U29273 (N_29273,N_29132,N_29021);
nand U29274 (N_29274,N_29059,N_29069);
or U29275 (N_29275,N_29006,N_29027);
nand U29276 (N_29276,N_29061,N_29162);
or U29277 (N_29277,N_29139,N_29124);
nor U29278 (N_29278,N_29180,N_29039);
xnor U29279 (N_29279,N_29161,N_29142);
nor U29280 (N_29280,N_29152,N_29062);
nor U29281 (N_29281,N_29004,N_29119);
nor U29282 (N_29282,N_29141,N_29015);
xor U29283 (N_29283,N_29148,N_29009);
nor U29284 (N_29284,N_29030,N_29091);
or U29285 (N_29285,N_29183,N_29173);
nor U29286 (N_29286,N_29181,N_29150);
xnor U29287 (N_29287,N_29171,N_29045);
nand U29288 (N_29288,N_29094,N_29023);
xnor U29289 (N_29289,N_29186,N_29088);
nor U29290 (N_29290,N_29068,N_29109);
nor U29291 (N_29291,N_29064,N_29197);
nor U29292 (N_29292,N_29008,N_29099);
and U29293 (N_29293,N_29035,N_29085);
xor U29294 (N_29294,N_29073,N_29051);
or U29295 (N_29295,N_29084,N_29110);
nand U29296 (N_29296,N_29034,N_29127);
and U29297 (N_29297,N_29107,N_29118);
nor U29298 (N_29298,N_29016,N_29138);
nor U29299 (N_29299,N_29172,N_29151);
nor U29300 (N_29300,N_29101,N_29120);
xnor U29301 (N_29301,N_29008,N_29137);
xor U29302 (N_29302,N_29135,N_29107);
nand U29303 (N_29303,N_29179,N_29045);
or U29304 (N_29304,N_29183,N_29129);
xor U29305 (N_29305,N_29181,N_29182);
xor U29306 (N_29306,N_29184,N_29078);
or U29307 (N_29307,N_29125,N_29061);
nand U29308 (N_29308,N_29020,N_29169);
and U29309 (N_29309,N_29095,N_29022);
nor U29310 (N_29310,N_29083,N_29078);
xnor U29311 (N_29311,N_29134,N_29063);
or U29312 (N_29312,N_29191,N_29011);
nor U29313 (N_29313,N_29006,N_29164);
or U29314 (N_29314,N_29051,N_29046);
nor U29315 (N_29315,N_29125,N_29115);
and U29316 (N_29316,N_29168,N_29016);
nand U29317 (N_29317,N_29081,N_29181);
xnor U29318 (N_29318,N_29035,N_29076);
nor U29319 (N_29319,N_29167,N_29036);
nor U29320 (N_29320,N_29137,N_29004);
xor U29321 (N_29321,N_29184,N_29136);
nor U29322 (N_29322,N_29162,N_29082);
or U29323 (N_29323,N_29026,N_29096);
nor U29324 (N_29324,N_29033,N_29112);
nor U29325 (N_29325,N_29143,N_29037);
and U29326 (N_29326,N_29065,N_29073);
nor U29327 (N_29327,N_29126,N_29000);
and U29328 (N_29328,N_29166,N_29078);
or U29329 (N_29329,N_29112,N_29154);
nand U29330 (N_29330,N_29157,N_29108);
or U29331 (N_29331,N_29131,N_29139);
nand U29332 (N_29332,N_29182,N_29160);
nor U29333 (N_29333,N_29199,N_29101);
nor U29334 (N_29334,N_29145,N_29198);
or U29335 (N_29335,N_29026,N_29141);
nor U29336 (N_29336,N_29076,N_29019);
xor U29337 (N_29337,N_29092,N_29103);
or U29338 (N_29338,N_29190,N_29112);
or U29339 (N_29339,N_29016,N_29118);
or U29340 (N_29340,N_29011,N_29054);
nor U29341 (N_29341,N_29159,N_29034);
xor U29342 (N_29342,N_29142,N_29043);
nor U29343 (N_29343,N_29079,N_29132);
or U29344 (N_29344,N_29135,N_29123);
or U29345 (N_29345,N_29199,N_29118);
and U29346 (N_29346,N_29048,N_29186);
nor U29347 (N_29347,N_29103,N_29140);
nor U29348 (N_29348,N_29108,N_29006);
nand U29349 (N_29349,N_29111,N_29046);
and U29350 (N_29350,N_29051,N_29084);
and U29351 (N_29351,N_29106,N_29029);
and U29352 (N_29352,N_29074,N_29163);
xnor U29353 (N_29353,N_29192,N_29166);
xor U29354 (N_29354,N_29157,N_29088);
nor U29355 (N_29355,N_29171,N_29010);
nand U29356 (N_29356,N_29094,N_29163);
or U29357 (N_29357,N_29091,N_29021);
and U29358 (N_29358,N_29095,N_29016);
nand U29359 (N_29359,N_29064,N_29039);
and U29360 (N_29360,N_29122,N_29078);
nand U29361 (N_29361,N_29074,N_29135);
or U29362 (N_29362,N_29047,N_29103);
or U29363 (N_29363,N_29003,N_29109);
nor U29364 (N_29364,N_29147,N_29165);
nor U29365 (N_29365,N_29195,N_29022);
xnor U29366 (N_29366,N_29069,N_29024);
nor U29367 (N_29367,N_29006,N_29096);
and U29368 (N_29368,N_29047,N_29161);
nor U29369 (N_29369,N_29149,N_29026);
and U29370 (N_29370,N_29133,N_29091);
nor U29371 (N_29371,N_29183,N_29117);
and U29372 (N_29372,N_29093,N_29116);
nor U29373 (N_29373,N_29095,N_29162);
or U29374 (N_29374,N_29098,N_29045);
and U29375 (N_29375,N_29082,N_29084);
or U29376 (N_29376,N_29074,N_29050);
and U29377 (N_29377,N_29039,N_29191);
or U29378 (N_29378,N_29018,N_29171);
or U29379 (N_29379,N_29134,N_29127);
xor U29380 (N_29380,N_29138,N_29068);
or U29381 (N_29381,N_29014,N_29134);
or U29382 (N_29382,N_29094,N_29099);
xnor U29383 (N_29383,N_29185,N_29199);
nand U29384 (N_29384,N_29172,N_29148);
or U29385 (N_29385,N_29030,N_29128);
and U29386 (N_29386,N_29046,N_29106);
nand U29387 (N_29387,N_29081,N_29022);
nand U29388 (N_29388,N_29165,N_29092);
nand U29389 (N_29389,N_29074,N_29118);
and U29390 (N_29390,N_29148,N_29121);
or U29391 (N_29391,N_29138,N_29127);
nor U29392 (N_29392,N_29058,N_29091);
nand U29393 (N_29393,N_29099,N_29176);
and U29394 (N_29394,N_29133,N_29115);
nor U29395 (N_29395,N_29115,N_29044);
xor U29396 (N_29396,N_29160,N_29174);
or U29397 (N_29397,N_29188,N_29090);
and U29398 (N_29398,N_29199,N_29096);
nor U29399 (N_29399,N_29043,N_29060);
xor U29400 (N_29400,N_29285,N_29219);
nor U29401 (N_29401,N_29329,N_29349);
nor U29402 (N_29402,N_29236,N_29322);
nand U29403 (N_29403,N_29304,N_29237);
and U29404 (N_29404,N_29227,N_29280);
nand U29405 (N_29405,N_29374,N_29397);
and U29406 (N_29406,N_29294,N_29216);
or U29407 (N_29407,N_29261,N_29281);
nand U29408 (N_29408,N_29312,N_29346);
and U29409 (N_29409,N_29299,N_29303);
or U29410 (N_29410,N_29319,N_29362);
and U29411 (N_29411,N_29262,N_29300);
nor U29412 (N_29412,N_29347,N_29241);
nor U29413 (N_29413,N_29283,N_29222);
nor U29414 (N_29414,N_29291,N_29268);
nor U29415 (N_29415,N_29357,N_29399);
or U29416 (N_29416,N_29259,N_29325);
nor U29417 (N_29417,N_29214,N_29278);
and U29418 (N_29418,N_29260,N_29247);
nand U29419 (N_29419,N_29373,N_29257);
and U29420 (N_29420,N_29258,N_29209);
nand U29421 (N_29421,N_29213,N_29231);
and U29422 (N_29422,N_29244,N_29395);
nor U29423 (N_29423,N_29310,N_29384);
or U29424 (N_29424,N_29361,N_29343);
nor U29425 (N_29425,N_29314,N_29263);
xnor U29426 (N_29426,N_29345,N_29334);
nand U29427 (N_29427,N_29298,N_29243);
or U29428 (N_29428,N_29206,N_29210);
xnor U29429 (N_29429,N_29389,N_29321);
or U29430 (N_29430,N_29223,N_29335);
nand U29431 (N_29431,N_29306,N_29234);
xor U29432 (N_29432,N_29255,N_29324);
xor U29433 (N_29433,N_29352,N_29228);
and U29434 (N_29434,N_29390,N_29235);
nand U29435 (N_29435,N_29201,N_29264);
or U29436 (N_29436,N_29360,N_29383);
nor U29437 (N_29437,N_29368,N_29230);
nand U29438 (N_29438,N_29240,N_29363);
or U29439 (N_29439,N_29381,N_29256);
nor U29440 (N_29440,N_29203,N_29246);
and U29441 (N_29441,N_29317,N_29323);
nand U29442 (N_29442,N_29242,N_29250);
and U29443 (N_29443,N_29270,N_29356);
nor U29444 (N_29444,N_29202,N_29277);
and U29445 (N_29445,N_29251,N_29311);
xnor U29446 (N_29446,N_29287,N_29279);
or U29447 (N_29447,N_29269,N_29238);
xor U29448 (N_29448,N_29341,N_29318);
and U29449 (N_29449,N_29387,N_29286);
nor U29450 (N_29450,N_29232,N_29284);
xnor U29451 (N_29451,N_29315,N_29305);
or U29452 (N_29452,N_29328,N_29372);
and U29453 (N_29453,N_29375,N_29313);
or U29454 (N_29454,N_29377,N_29288);
and U29455 (N_29455,N_29394,N_29273);
nand U29456 (N_29456,N_29364,N_29386);
and U29457 (N_29457,N_29342,N_29393);
nor U29458 (N_29458,N_29379,N_29275);
nor U29459 (N_29459,N_29365,N_29391);
and U29460 (N_29460,N_29339,N_29371);
and U29461 (N_29461,N_29204,N_29239);
xor U29462 (N_29462,N_29370,N_29332);
nor U29463 (N_29463,N_29233,N_29296);
and U29464 (N_29464,N_29366,N_29308);
nor U29465 (N_29465,N_29336,N_29289);
nor U29466 (N_29466,N_29205,N_29224);
and U29467 (N_29467,N_29378,N_29354);
nand U29468 (N_29468,N_29307,N_29316);
xor U29469 (N_29469,N_29200,N_29327);
nand U29470 (N_29470,N_29309,N_29272);
or U29471 (N_29471,N_29271,N_29226);
xnor U29472 (N_29472,N_29208,N_29398);
or U29473 (N_29473,N_29282,N_29274);
nand U29474 (N_29474,N_29396,N_29266);
nand U29475 (N_29475,N_29292,N_29382);
nor U29476 (N_29476,N_29380,N_29326);
and U29477 (N_29477,N_29297,N_29249);
nor U29478 (N_29478,N_29344,N_29225);
or U29479 (N_29479,N_29295,N_29252);
or U29480 (N_29480,N_29348,N_29367);
nand U29481 (N_29481,N_29355,N_29359);
and U29482 (N_29482,N_29221,N_29350);
nand U29483 (N_29483,N_29385,N_29265);
xnor U29484 (N_29484,N_29215,N_29290);
and U29485 (N_29485,N_29330,N_29337);
xor U29486 (N_29486,N_29207,N_29320);
nor U29487 (N_29487,N_29229,N_29331);
xor U29488 (N_29488,N_29338,N_29211);
xor U29489 (N_29489,N_29254,N_29212);
xnor U29490 (N_29490,N_29392,N_29253);
xor U29491 (N_29491,N_29376,N_29217);
nand U29492 (N_29492,N_29358,N_29302);
or U29493 (N_29493,N_29340,N_29267);
nand U29494 (N_29494,N_29369,N_29293);
xor U29495 (N_29495,N_29301,N_29388);
and U29496 (N_29496,N_29248,N_29245);
or U29497 (N_29497,N_29333,N_29351);
nor U29498 (N_29498,N_29276,N_29353);
nor U29499 (N_29499,N_29218,N_29220);
and U29500 (N_29500,N_29237,N_29300);
nand U29501 (N_29501,N_29311,N_29252);
or U29502 (N_29502,N_29215,N_29207);
nand U29503 (N_29503,N_29269,N_29277);
nor U29504 (N_29504,N_29249,N_29242);
nand U29505 (N_29505,N_29227,N_29312);
nand U29506 (N_29506,N_29312,N_29352);
xor U29507 (N_29507,N_29376,N_29329);
or U29508 (N_29508,N_29364,N_29265);
nand U29509 (N_29509,N_29320,N_29376);
nor U29510 (N_29510,N_29382,N_29390);
nor U29511 (N_29511,N_29312,N_29318);
nor U29512 (N_29512,N_29298,N_29338);
nand U29513 (N_29513,N_29306,N_29273);
xnor U29514 (N_29514,N_29294,N_29274);
or U29515 (N_29515,N_29356,N_29263);
or U29516 (N_29516,N_29330,N_29279);
nor U29517 (N_29517,N_29208,N_29351);
xor U29518 (N_29518,N_29351,N_29349);
or U29519 (N_29519,N_29231,N_29380);
nand U29520 (N_29520,N_29238,N_29226);
nor U29521 (N_29521,N_29391,N_29362);
xnor U29522 (N_29522,N_29245,N_29310);
xnor U29523 (N_29523,N_29378,N_29326);
and U29524 (N_29524,N_29388,N_29387);
and U29525 (N_29525,N_29265,N_29230);
nor U29526 (N_29526,N_29236,N_29232);
xor U29527 (N_29527,N_29205,N_29225);
xor U29528 (N_29528,N_29350,N_29328);
nor U29529 (N_29529,N_29262,N_29215);
or U29530 (N_29530,N_29397,N_29327);
xnor U29531 (N_29531,N_29224,N_29299);
nand U29532 (N_29532,N_29329,N_29312);
nand U29533 (N_29533,N_29385,N_29386);
nor U29534 (N_29534,N_29238,N_29252);
and U29535 (N_29535,N_29266,N_29262);
or U29536 (N_29536,N_29221,N_29201);
and U29537 (N_29537,N_29202,N_29320);
nand U29538 (N_29538,N_29245,N_29262);
or U29539 (N_29539,N_29335,N_29345);
xor U29540 (N_29540,N_29308,N_29365);
xor U29541 (N_29541,N_29278,N_29203);
or U29542 (N_29542,N_29397,N_29273);
nand U29543 (N_29543,N_29302,N_29323);
and U29544 (N_29544,N_29359,N_29274);
and U29545 (N_29545,N_29363,N_29392);
nor U29546 (N_29546,N_29326,N_29363);
xor U29547 (N_29547,N_29273,N_29390);
nor U29548 (N_29548,N_29311,N_29387);
nand U29549 (N_29549,N_29307,N_29224);
and U29550 (N_29550,N_29225,N_29311);
nand U29551 (N_29551,N_29380,N_29277);
xnor U29552 (N_29552,N_29289,N_29250);
nor U29553 (N_29553,N_29294,N_29219);
nor U29554 (N_29554,N_29372,N_29394);
nand U29555 (N_29555,N_29365,N_29284);
nor U29556 (N_29556,N_29398,N_29368);
nand U29557 (N_29557,N_29232,N_29326);
and U29558 (N_29558,N_29344,N_29389);
or U29559 (N_29559,N_29381,N_29330);
or U29560 (N_29560,N_29286,N_29283);
nor U29561 (N_29561,N_29329,N_29306);
nor U29562 (N_29562,N_29202,N_29210);
and U29563 (N_29563,N_29327,N_29381);
xor U29564 (N_29564,N_29388,N_29302);
nand U29565 (N_29565,N_29383,N_29292);
nand U29566 (N_29566,N_29351,N_29202);
nor U29567 (N_29567,N_29376,N_29315);
nand U29568 (N_29568,N_29398,N_29374);
nor U29569 (N_29569,N_29292,N_29276);
or U29570 (N_29570,N_29389,N_29323);
or U29571 (N_29571,N_29360,N_29262);
nand U29572 (N_29572,N_29395,N_29325);
nand U29573 (N_29573,N_29355,N_29223);
nand U29574 (N_29574,N_29267,N_29211);
nand U29575 (N_29575,N_29211,N_29374);
nand U29576 (N_29576,N_29396,N_29361);
and U29577 (N_29577,N_29389,N_29239);
or U29578 (N_29578,N_29356,N_29277);
nand U29579 (N_29579,N_29348,N_29279);
or U29580 (N_29580,N_29334,N_29212);
or U29581 (N_29581,N_29247,N_29314);
xor U29582 (N_29582,N_29334,N_29265);
or U29583 (N_29583,N_29242,N_29345);
xnor U29584 (N_29584,N_29261,N_29286);
and U29585 (N_29585,N_29289,N_29238);
nor U29586 (N_29586,N_29351,N_29395);
and U29587 (N_29587,N_29365,N_29222);
and U29588 (N_29588,N_29240,N_29306);
nor U29589 (N_29589,N_29232,N_29243);
and U29590 (N_29590,N_29376,N_29360);
and U29591 (N_29591,N_29375,N_29298);
and U29592 (N_29592,N_29319,N_29279);
xnor U29593 (N_29593,N_29330,N_29364);
and U29594 (N_29594,N_29219,N_29296);
or U29595 (N_29595,N_29251,N_29340);
nor U29596 (N_29596,N_29292,N_29222);
or U29597 (N_29597,N_29242,N_29309);
and U29598 (N_29598,N_29286,N_29349);
xnor U29599 (N_29599,N_29362,N_29294);
or U29600 (N_29600,N_29456,N_29514);
xor U29601 (N_29601,N_29431,N_29411);
xor U29602 (N_29602,N_29533,N_29439);
and U29603 (N_29603,N_29459,N_29472);
nor U29604 (N_29604,N_29499,N_29429);
nand U29605 (N_29605,N_29490,N_29538);
nor U29606 (N_29606,N_29589,N_29495);
nand U29607 (N_29607,N_29583,N_29443);
or U29608 (N_29608,N_29572,N_29445);
nor U29609 (N_29609,N_29547,N_29436);
or U29610 (N_29610,N_29484,N_29470);
or U29611 (N_29611,N_29465,N_29506);
nand U29612 (N_29612,N_29502,N_29466);
and U29613 (N_29613,N_29414,N_29556);
or U29614 (N_29614,N_29468,N_29524);
xor U29615 (N_29615,N_29554,N_29534);
or U29616 (N_29616,N_29564,N_29575);
or U29617 (N_29617,N_29562,N_29508);
and U29618 (N_29618,N_29433,N_29475);
and U29619 (N_29619,N_29510,N_29457);
nand U29620 (N_29620,N_29413,N_29567);
xor U29621 (N_29621,N_29400,N_29594);
or U29622 (N_29622,N_29549,N_29550);
nand U29623 (N_29623,N_29535,N_29590);
nand U29624 (N_29624,N_29463,N_29428);
nor U29625 (N_29625,N_29512,N_29530);
xor U29626 (N_29626,N_29426,N_29476);
nor U29627 (N_29627,N_29487,N_29507);
or U29628 (N_29628,N_29541,N_29523);
nor U29629 (N_29629,N_29409,N_29489);
xor U29630 (N_29630,N_29473,N_29498);
or U29631 (N_29631,N_29454,N_29532);
nor U29632 (N_29632,N_29477,N_29559);
xnor U29633 (N_29633,N_29441,N_29452);
xnor U29634 (N_29634,N_29587,N_29555);
nor U29635 (N_29635,N_29460,N_29427);
xnor U29636 (N_29636,N_29513,N_29479);
and U29637 (N_29637,N_29561,N_29520);
nor U29638 (N_29638,N_29417,N_29503);
xor U29639 (N_29639,N_29406,N_29551);
nor U29640 (N_29640,N_29595,N_29596);
or U29641 (N_29641,N_29584,N_29416);
and U29642 (N_29642,N_29405,N_29599);
or U29643 (N_29643,N_29464,N_29423);
nand U29644 (N_29644,N_29424,N_29519);
nor U29645 (N_29645,N_29432,N_29467);
nor U29646 (N_29646,N_29412,N_29402);
and U29647 (N_29647,N_29580,N_29573);
and U29648 (N_29648,N_29453,N_29415);
xor U29649 (N_29649,N_29482,N_29557);
and U29650 (N_29650,N_29518,N_29435);
and U29651 (N_29651,N_29418,N_29592);
or U29652 (N_29652,N_29521,N_29545);
xnor U29653 (N_29653,N_29516,N_29537);
and U29654 (N_29654,N_29563,N_29568);
and U29655 (N_29655,N_29585,N_29419);
nand U29656 (N_29656,N_29544,N_29420);
xnor U29657 (N_29657,N_29548,N_29474);
xor U29658 (N_29658,N_29430,N_29449);
xor U29659 (N_29659,N_29522,N_29598);
or U29660 (N_29660,N_29597,N_29483);
nor U29661 (N_29661,N_29494,N_29408);
nand U29662 (N_29662,N_29438,N_29403);
nand U29663 (N_29663,N_29500,N_29488);
nor U29664 (N_29664,N_29511,N_29505);
or U29665 (N_29665,N_29491,N_29496);
xnor U29666 (N_29666,N_29434,N_29539);
nor U29667 (N_29667,N_29444,N_29586);
nand U29668 (N_29668,N_29478,N_29421);
nand U29669 (N_29669,N_29581,N_29455);
and U29670 (N_29670,N_29553,N_29566);
nand U29671 (N_29671,N_29558,N_29571);
and U29672 (N_29672,N_29579,N_29440);
or U29673 (N_29673,N_29570,N_29471);
and U29674 (N_29674,N_29536,N_29552);
and U29675 (N_29675,N_29577,N_29565);
nor U29676 (N_29676,N_29569,N_29458);
and U29677 (N_29677,N_29543,N_29492);
or U29678 (N_29678,N_29560,N_29401);
or U29679 (N_29679,N_29410,N_29504);
and U29680 (N_29680,N_29480,N_29407);
nand U29681 (N_29681,N_29461,N_29425);
nand U29682 (N_29682,N_29593,N_29515);
xnor U29683 (N_29683,N_29486,N_29442);
and U29684 (N_29684,N_29582,N_29448);
nor U29685 (N_29685,N_29447,N_29437);
and U29686 (N_29686,N_29497,N_29588);
nand U29687 (N_29687,N_29576,N_29469);
and U29688 (N_29688,N_29451,N_29446);
nor U29689 (N_29689,N_29462,N_29525);
xor U29690 (N_29690,N_29493,N_29578);
and U29691 (N_29691,N_29501,N_29542);
nand U29692 (N_29692,N_29528,N_29529);
and U29693 (N_29693,N_29526,N_29450);
and U29694 (N_29694,N_29485,N_29527);
nand U29695 (N_29695,N_29574,N_29509);
nand U29696 (N_29696,N_29481,N_29546);
nand U29697 (N_29697,N_29540,N_29517);
nand U29698 (N_29698,N_29591,N_29531);
xnor U29699 (N_29699,N_29422,N_29404);
or U29700 (N_29700,N_29413,N_29505);
and U29701 (N_29701,N_29557,N_29513);
xor U29702 (N_29702,N_29567,N_29547);
xnor U29703 (N_29703,N_29575,N_29441);
and U29704 (N_29704,N_29434,N_29498);
or U29705 (N_29705,N_29588,N_29455);
or U29706 (N_29706,N_29518,N_29469);
and U29707 (N_29707,N_29493,N_29449);
or U29708 (N_29708,N_29465,N_29462);
nand U29709 (N_29709,N_29478,N_29497);
or U29710 (N_29710,N_29545,N_29558);
or U29711 (N_29711,N_29561,N_29578);
or U29712 (N_29712,N_29443,N_29501);
nor U29713 (N_29713,N_29529,N_29458);
or U29714 (N_29714,N_29595,N_29579);
and U29715 (N_29715,N_29565,N_29487);
nor U29716 (N_29716,N_29547,N_29421);
or U29717 (N_29717,N_29555,N_29557);
xor U29718 (N_29718,N_29455,N_29420);
xnor U29719 (N_29719,N_29408,N_29536);
and U29720 (N_29720,N_29596,N_29528);
or U29721 (N_29721,N_29590,N_29448);
xor U29722 (N_29722,N_29574,N_29523);
and U29723 (N_29723,N_29452,N_29421);
nor U29724 (N_29724,N_29471,N_29559);
or U29725 (N_29725,N_29545,N_29472);
nand U29726 (N_29726,N_29484,N_29488);
nor U29727 (N_29727,N_29578,N_29487);
nor U29728 (N_29728,N_29596,N_29548);
xnor U29729 (N_29729,N_29559,N_29597);
and U29730 (N_29730,N_29490,N_29451);
and U29731 (N_29731,N_29592,N_29561);
and U29732 (N_29732,N_29406,N_29506);
nand U29733 (N_29733,N_29405,N_29555);
nand U29734 (N_29734,N_29494,N_29547);
nand U29735 (N_29735,N_29597,N_29409);
xnor U29736 (N_29736,N_29523,N_29597);
or U29737 (N_29737,N_29406,N_29555);
nand U29738 (N_29738,N_29470,N_29462);
nand U29739 (N_29739,N_29505,N_29544);
xor U29740 (N_29740,N_29451,N_29447);
nand U29741 (N_29741,N_29519,N_29447);
xnor U29742 (N_29742,N_29520,N_29439);
nor U29743 (N_29743,N_29452,N_29548);
xor U29744 (N_29744,N_29441,N_29529);
or U29745 (N_29745,N_29447,N_29494);
and U29746 (N_29746,N_29433,N_29464);
xnor U29747 (N_29747,N_29538,N_29420);
nor U29748 (N_29748,N_29490,N_29545);
nand U29749 (N_29749,N_29458,N_29599);
nand U29750 (N_29750,N_29487,N_29510);
xnor U29751 (N_29751,N_29419,N_29586);
xnor U29752 (N_29752,N_29588,N_29482);
nor U29753 (N_29753,N_29584,N_29535);
xnor U29754 (N_29754,N_29478,N_29431);
xor U29755 (N_29755,N_29564,N_29480);
xor U29756 (N_29756,N_29408,N_29485);
xnor U29757 (N_29757,N_29574,N_29419);
nand U29758 (N_29758,N_29442,N_29437);
nor U29759 (N_29759,N_29583,N_29508);
xor U29760 (N_29760,N_29504,N_29561);
and U29761 (N_29761,N_29540,N_29529);
nor U29762 (N_29762,N_29406,N_29491);
nand U29763 (N_29763,N_29438,N_29475);
nand U29764 (N_29764,N_29443,N_29559);
and U29765 (N_29765,N_29538,N_29553);
or U29766 (N_29766,N_29590,N_29409);
xor U29767 (N_29767,N_29516,N_29568);
or U29768 (N_29768,N_29583,N_29432);
nand U29769 (N_29769,N_29514,N_29583);
or U29770 (N_29770,N_29517,N_29498);
nor U29771 (N_29771,N_29563,N_29464);
nor U29772 (N_29772,N_29595,N_29496);
xor U29773 (N_29773,N_29402,N_29495);
and U29774 (N_29774,N_29409,N_29553);
nand U29775 (N_29775,N_29428,N_29410);
and U29776 (N_29776,N_29552,N_29510);
or U29777 (N_29777,N_29400,N_29528);
and U29778 (N_29778,N_29408,N_29515);
nor U29779 (N_29779,N_29557,N_29553);
and U29780 (N_29780,N_29506,N_29518);
nand U29781 (N_29781,N_29525,N_29416);
xnor U29782 (N_29782,N_29514,N_29460);
and U29783 (N_29783,N_29594,N_29438);
nor U29784 (N_29784,N_29444,N_29552);
and U29785 (N_29785,N_29512,N_29574);
xor U29786 (N_29786,N_29449,N_29533);
nand U29787 (N_29787,N_29524,N_29425);
nand U29788 (N_29788,N_29479,N_29420);
or U29789 (N_29789,N_29539,N_29460);
nand U29790 (N_29790,N_29437,N_29548);
xor U29791 (N_29791,N_29581,N_29566);
and U29792 (N_29792,N_29591,N_29473);
xor U29793 (N_29793,N_29470,N_29458);
xor U29794 (N_29794,N_29440,N_29589);
or U29795 (N_29795,N_29582,N_29544);
or U29796 (N_29796,N_29599,N_29438);
and U29797 (N_29797,N_29414,N_29492);
or U29798 (N_29798,N_29409,N_29562);
nor U29799 (N_29799,N_29455,N_29437);
nand U29800 (N_29800,N_29708,N_29700);
nor U29801 (N_29801,N_29673,N_29611);
or U29802 (N_29802,N_29765,N_29618);
nor U29803 (N_29803,N_29751,N_29769);
and U29804 (N_29804,N_29785,N_29647);
xor U29805 (N_29805,N_29691,N_29733);
nor U29806 (N_29806,N_29768,N_29688);
nor U29807 (N_29807,N_29645,N_29652);
nor U29808 (N_29808,N_29764,N_29713);
and U29809 (N_29809,N_29616,N_29723);
or U29810 (N_29810,N_29752,N_29629);
nand U29811 (N_29811,N_29672,N_29731);
xnor U29812 (N_29812,N_29690,N_29797);
nand U29813 (N_29813,N_29716,N_29658);
nor U29814 (N_29814,N_29681,N_29780);
nor U29815 (N_29815,N_29650,N_29620);
xor U29816 (N_29816,N_29683,N_29715);
or U29817 (N_29817,N_29721,N_29678);
and U29818 (N_29818,N_29726,N_29653);
nand U29819 (N_29819,N_29692,N_29682);
nor U29820 (N_29820,N_29722,N_29703);
nand U29821 (N_29821,N_29759,N_29632);
nand U29822 (N_29822,N_29791,N_29627);
nand U29823 (N_29823,N_29702,N_29792);
nor U29824 (N_29824,N_29656,N_29675);
xor U29825 (N_29825,N_29711,N_29767);
nor U29826 (N_29826,N_29739,N_29660);
and U29827 (N_29827,N_29728,N_29646);
xor U29828 (N_29828,N_29609,N_29617);
nand U29829 (N_29829,N_29744,N_29799);
nor U29830 (N_29830,N_29724,N_29770);
and U29831 (N_29831,N_29619,N_29635);
xor U29832 (N_29832,N_29608,N_29709);
nor U29833 (N_29833,N_29626,N_29694);
xnor U29834 (N_29834,N_29734,N_29699);
or U29835 (N_29835,N_29643,N_29718);
nor U29836 (N_29836,N_29735,N_29630);
nand U29837 (N_29837,N_29606,N_29605);
nor U29838 (N_29838,N_29644,N_29707);
nor U29839 (N_29839,N_29754,N_29679);
or U29840 (N_29840,N_29732,N_29693);
xnor U29841 (N_29841,N_29657,N_29771);
or U29842 (N_29842,N_29738,N_29763);
and U29843 (N_29843,N_29798,N_29669);
nor U29844 (N_29844,N_29612,N_29725);
xor U29845 (N_29845,N_29737,N_29659);
nand U29846 (N_29846,N_29637,N_29782);
nand U29847 (N_29847,N_29680,N_29685);
nor U29848 (N_29848,N_29787,N_29729);
or U29849 (N_29849,N_29636,N_29640);
and U29850 (N_29850,N_29776,N_29697);
or U29851 (N_29851,N_29642,N_29775);
and U29852 (N_29852,N_29651,N_29689);
xor U29853 (N_29853,N_29623,N_29662);
and U29854 (N_29854,N_29638,N_29753);
nor U29855 (N_29855,N_29670,N_29760);
xor U29856 (N_29856,N_29602,N_29757);
nand U29857 (N_29857,N_29793,N_29667);
and U29858 (N_29858,N_29796,N_29666);
xor U29859 (N_29859,N_29788,N_29600);
xor U29860 (N_29860,N_29712,N_29746);
or U29861 (N_29861,N_29668,N_29756);
and U29862 (N_29862,N_29701,N_29621);
and U29863 (N_29863,N_29761,N_29736);
nand U29864 (N_29864,N_29624,N_29661);
and U29865 (N_29865,N_29789,N_29622);
or U29866 (N_29866,N_29677,N_29698);
nor U29867 (N_29867,N_29654,N_29663);
nand U29868 (N_29868,N_29604,N_29634);
and U29869 (N_29869,N_29648,N_29784);
xnor U29870 (N_29870,N_29727,N_29706);
nand U29871 (N_29871,N_29649,N_29664);
nor U29872 (N_29872,N_29613,N_29686);
nor U29873 (N_29873,N_29783,N_29665);
and U29874 (N_29874,N_29773,N_29714);
nand U29875 (N_29875,N_29740,N_29601);
or U29876 (N_29876,N_29684,N_29743);
or U29877 (N_29877,N_29781,N_29614);
or U29878 (N_29878,N_29717,N_29631);
or U29879 (N_29879,N_29655,N_29696);
xnor U29880 (N_29880,N_29625,N_29676);
nand U29881 (N_29881,N_29720,N_29778);
nor U29882 (N_29882,N_29705,N_29790);
or U29883 (N_29883,N_29710,N_29687);
or U29884 (N_29884,N_29755,N_29674);
xnor U29885 (N_29885,N_29610,N_29730);
or U29886 (N_29886,N_29749,N_29786);
nor U29887 (N_29887,N_29741,N_29794);
nor U29888 (N_29888,N_29758,N_29719);
nand U29889 (N_29889,N_29671,N_29766);
or U29890 (N_29890,N_29628,N_29615);
and U29891 (N_29891,N_29779,N_29747);
nand U29892 (N_29892,N_29772,N_29633);
and U29893 (N_29893,N_29774,N_29607);
nor U29894 (N_29894,N_29762,N_29750);
nor U29895 (N_29895,N_29777,N_29641);
nor U29896 (N_29896,N_29639,N_29695);
and U29897 (N_29897,N_29704,N_29795);
xor U29898 (N_29898,N_29742,N_29603);
nand U29899 (N_29899,N_29745,N_29748);
and U29900 (N_29900,N_29720,N_29629);
and U29901 (N_29901,N_29712,N_29729);
nand U29902 (N_29902,N_29685,N_29730);
or U29903 (N_29903,N_29790,N_29719);
nand U29904 (N_29904,N_29722,N_29624);
or U29905 (N_29905,N_29607,N_29789);
or U29906 (N_29906,N_29613,N_29714);
nor U29907 (N_29907,N_29758,N_29675);
and U29908 (N_29908,N_29621,N_29796);
xnor U29909 (N_29909,N_29762,N_29636);
xor U29910 (N_29910,N_29692,N_29727);
xor U29911 (N_29911,N_29702,N_29663);
nand U29912 (N_29912,N_29690,N_29723);
xnor U29913 (N_29913,N_29727,N_29623);
nand U29914 (N_29914,N_29603,N_29757);
xnor U29915 (N_29915,N_29780,N_29645);
nand U29916 (N_29916,N_29644,N_29780);
and U29917 (N_29917,N_29776,N_29740);
xor U29918 (N_29918,N_29655,N_29680);
nand U29919 (N_29919,N_29748,N_29648);
or U29920 (N_29920,N_29654,N_29620);
and U29921 (N_29921,N_29663,N_29776);
nor U29922 (N_29922,N_29660,N_29675);
nand U29923 (N_29923,N_29602,N_29726);
nor U29924 (N_29924,N_29647,N_29721);
or U29925 (N_29925,N_29630,N_29783);
xor U29926 (N_29926,N_29673,N_29691);
or U29927 (N_29927,N_29684,N_29718);
or U29928 (N_29928,N_29636,N_29614);
xnor U29929 (N_29929,N_29635,N_29705);
or U29930 (N_29930,N_29779,N_29628);
xor U29931 (N_29931,N_29792,N_29718);
or U29932 (N_29932,N_29639,N_29732);
xnor U29933 (N_29933,N_29764,N_29621);
and U29934 (N_29934,N_29781,N_29623);
nor U29935 (N_29935,N_29767,N_29655);
nor U29936 (N_29936,N_29776,N_29603);
xor U29937 (N_29937,N_29603,N_29686);
or U29938 (N_29938,N_29770,N_29697);
nand U29939 (N_29939,N_29626,N_29695);
nand U29940 (N_29940,N_29768,N_29685);
or U29941 (N_29941,N_29640,N_29603);
nor U29942 (N_29942,N_29659,N_29704);
xor U29943 (N_29943,N_29752,N_29607);
nor U29944 (N_29944,N_29635,N_29676);
xor U29945 (N_29945,N_29698,N_29701);
nand U29946 (N_29946,N_29711,N_29734);
nor U29947 (N_29947,N_29623,N_29644);
or U29948 (N_29948,N_29716,N_29789);
nor U29949 (N_29949,N_29743,N_29654);
nand U29950 (N_29950,N_29636,N_29727);
nand U29951 (N_29951,N_29606,N_29662);
or U29952 (N_29952,N_29697,N_29682);
or U29953 (N_29953,N_29600,N_29687);
nor U29954 (N_29954,N_29643,N_29601);
and U29955 (N_29955,N_29709,N_29609);
xor U29956 (N_29956,N_29781,N_29721);
and U29957 (N_29957,N_29627,N_29624);
xnor U29958 (N_29958,N_29664,N_29768);
and U29959 (N_29959,N_29618,N_29631);
or U29960 (N_29960,N_29754,N_29661);
nor U29961 (N_29961,N_29627,N_29740);
or U29962 (N_29962,N_29727,N_29607);
or U29963 (N_29963,N_29694,N_29789);
nor U29964 (N_29964,N_29717,N_29617);
or U29965 (N_29965,N_29707,N_29673);
and U29966 (N_29966,N_29655,N_29641);
and U29967 (N_29967,N_29752,N_29710);
or U29968 (N_29968,N_29782,N_29733);
nor U29969 (N_29969,N_29636,N_29605);
nand U29970 (N_29970,N_29742,N_29722);
and U29971 (N_29971,N_29797,N_29628);
nand U29972 (N_29972,N_29772,N_29652);
nand U29973 (N_29973,N_29645,N_29730);
nand U29974 (N_29974,N_29631,N_29736);
and U29975 (N_29975,N_29730,N_29617);
or U29976 (N_29976,N_29769,N_29657);
nor U29977 (N_29977,N_29704,N_29677);
or U29978 (N_29978,N_29655,N_29784);
and U29979 (N_29979,N_29615,N_29683);
xnor U29980 (N_29980,N_29742,N_29778);
or U29981 (N_29981,N_29624,N_29693);
or U29982 (N_29982,N_29735,N_29768);
nor U29983 (N_29983,N_29774,N_29697);
nor U29984 (N_29984,N_29620,N_29630);
nor U29985 (N_29985,N_29685,N_29778);
or U29986 (N_29986,N_29691,N_29636);
nand U29987 (N_29987,N_29745,N_29771);
nand U29988 (N_29988,N_29777,N_29657);
and U29989 (N_29989,N_29695,N_29728);
nor U29990 (N_29990,N_29743,N_29685);
or U29991 (N_29991,N_29733,N_29685);
xnor U29992 (N_29992,N_29706,N_29603);
or U29993 (N_29993,N_29773,N_29735);
nor U29994 (N_29994,N_29694,N_29663);
or U29995 (N_29995,N_29615,N_29658);
nor U29996 (N_29996,N_29721,N_29626);
nor U29997 (N_29997,N_29784,N_29733);
and U29998 (N_29998,N_29643,N_29688);
or U29999 (N_29999,N_29613,N_29607);
or UO_0 (O_0,N_29866,N_29995);
xor UO_1 (O_1,N_29922,N_29855);
nor UO_2 (O_2,N_29972,N_29896);
xor UO_3 (O_3,N_29850,N_29973);
xor UO_4 (O_4,N_29942,N_29878);
or UO_5 (O_5,N_29981,N_29867);
and UO_6 (O_6,N_29858,N_29841);
nand UO_7 (O_7,N_29911,N_29929);
xor UO_8 (O_8,N_29950,N_29905);
xnor UO_9 (O_9,N_29868,N_29884);
or UO_10 (O_10,N_29829,N_29835);
or UO_11 (O_11,N_29849,N_29809);
xor UO_12 (O_12,N_29812,N_29979);
nand UO_13 (O_13,N_29803,N_29976);
nand UO_14 (O_14,N_29894,N_29864);
or UO_15 (O_15,N_29932,N_29933);
nor UO_16 (O_16,N_29984,N_29926);
nand UO_17 (O_17,N_29805,N_29957);
and UO_18 (O_18,N_29895,N_29808);
or UO_19 (O_19,N_29987,N_29980);
nor UO_20 (O_20,N_29997,N_29916);
nor UO_21 (O_21,N_29844,N_29924);
xnor UO_22 (O_22,N_29879,N_29820);
or UO_23 (O_23,N_29901,N_29876);
nand UO_24 (O_24,N_29970,N_29815);
nor UO_25 (O_25,N_29989,N_29821);
and UO_26 (O_26,N_29843,N_29983);
nand UO_27 (O_27,N_29898,N_29985);
xor UO_28 (O_28,N_29890,N_29943);
xnor UO_29 (O_29,N_29910,N_29802);
xnor UO_30 (O_30,N_29927,N_29838);
or UO_31 (O_31,N_29880,N_29920);
nand UO_32 (O_32,N_29847,N_29968);
nor UO_33 (O_33,N_29857,N_29800);
nand UO_34 (O_34,N_29801,N_29982);
or UO_35 (O_35,N_29830,N_29919);
or UO_36 (O_36,N_29885,N_29832);
and UO_37 (O_37,N_29934,N_29912);
and UO_38 (O_38,N_29966,N_29915);
and UO_39 (O_39,N_29917,N_29931);
xor UO_40 (O_40,N_29831,N_29967);
or UO_41 (O_41,N_29807,N_29854);
or UO_42 (O_42,N_29992,N_29804);
and UO_43 (O_43,N_29842,N_29865);
nand UO_44 (O_44,N_29948,N_29994);
nand UO_45 (O_45,N_29883,N_29998);
or UO_46 (O_46,N_29827,N_29814);
xor UO_47 (O_47,N_29881,N_29913);
nand UO_48 (O_48,N_29952,N_29840);
or UO_49 (O_49,N_29860,N_29999);
xnor UO_50 (O_50,N_29940,N_29899);
or UO_51 (O_51,N_29897,N_29834);
nor UO_52 (O_52,N_29875,N_29816);
or UO_53 (O_53,N_29941,N_29823);
or UO_54 (O_54,N_29818,N_29991);
nand UO_55 (O_55,N_29951,N_29975);
or UO_56 (O_56,N_29944,N_29887);
and UO_57 (O_57,N_29882,N_29811);
nand UO_58 (O_58,N_29974,N_29956);
nand UO_59 (O_59,N_29873,N_29977);
and UO_60 (O_60,N_29963,N_29969);
or UO_61 (O_61,N_29978,N_29862);
nor UO_62 (O_62,N_29871,N_29837);
or UO_63 (O_63,N_29958,N_29848);
xnor UO_64 (O_64,N_29824,N_29889);
nand UO_65 (O_65,N_29909,N_29921);
or UO_66 (O_66,N_29851,N_29961);
nand UO_67 (O_67,N_29953,N_29856);
or UO_68 (O_68,N_29877,N_29874);
nand UO_69 (O_69,N_29904,N_29936);
xor UO_70 (O_70,N_29907,N_29965);
xnor UO_71 (O_71,N_29861,N_29918);
nor UO_72 (O_72,N_29930,N_29993);
xnor UO_73 (O_73,N_29836,N_29819);
xor UO_74 (O_74,N_29886,N_29959);
nand UO_75 (O_75,N_29870,N_29954);
xnor UO_76 (O_76,N_29852,N_29908);
and UO_77 (O_77,N_29828,N_29817);
or UO_78 (O_78,N_29833,N_29955);
or UO_79 (O_79,N_29839,N_29988);
and UO_80 (O_80,N_29825,N_29888);
nand UO_81 (O_81,N_29949,N_29900);
or UO_82 (O_82,N_29902,N_29962);
nand UO_83 (O_83,N_29892,N_29945);
or UO_84 (O_84,N_29938,N_29964);
or UO_85 (O_85,N_29947,N_29813);
and UO_86 (O_86,N_29946,N_29971);
nor UO_87 (O_87,N_29822,N_29939);
nor UO_88 (O_88,N_29806,N_29960);
nand UO_89 (O_89,N_29928,N_29891);
nor UO_90 (O_90,N_29925,N_29986);
xnor UO_91 (O_91,N_29914,N_29859);
or UO_92 (O_92,N_29990,N_29863);
xnor UO_93 (O_93,N_29853,N_29845);
and UO_94 (O_94,N_29935,N_29923);
or UO_95 (O_95,N_29893,N_29826);
or UO_96 (O_96,N_29869,N_29937);
or UO_97 (O_97,N_29903,N_29906);
or UO_98 (O_98,N_29810,N_29872);
xnor UO_99 (O_99,N_29846,N_29996);
or UO_100 (O_100,N_29981,N_29926);
nand UO_101 (O_101,N_29984,N_29978);
nand UO_102 (O_102,N_29933,N_29911);
or UO_103 (O_103,N_29828,N_29916);
nand UO_104 (O_104,N_29962,N_29953);
nor UO_105 (O_105,N_29898,N_29963);
nand UO_106 (O_106,N_29822,N_29933);
xor UO_107 (O_107,N_29956,N_29805);
or UO_108 (O_108,N_29800,N_29994);
xnor UO_109 (O_109,N_29900,N_29926);
nor UO_110 (O_110,N_29849,N_29998);
and UO_111 (O_111,N_29896,N_29904);
nand UO_112 (O_112,N_29996,N_29819);
nor UO_113 (O_113,N_29963,N_29825);
xnor UO_114 (O_114,N_29990,N_29844);
nand UO_115 (O_115,N_29966,N_29908);
nor UO_116 (O_116,N_29933,N_29841);
nand UO_117 (O_117,N_29807,N_29915);
and UO_118 (O_118,N_29868,N_29858);
xnor UO_119 (O_119,N_29807,N_29839);
nor UO_120 (O_120,N_29864,N_29960);
and UO_121 (O_121,N_29881,N_29935);
or UO_122 (O_122,N_29898,N_29880);
and UO_123 (O_123,N_29944,N_29926);
nor UO_124 (O_124,N_29873,N_29943);
or UO_125 (O_125,N_29844,N_29891);
nor UO_126 (O_126,N_29969,N_29888);
xnor UO_127 (O_127,N_29872,N_29939);
xnor UO_128 (O_128,N_29895,N_29908);
nor UO_129 (O_129,N_29854,N_29819);
xnor UO_130 (O_130,N_29926,N_29960);
and UO_131 (O_131,N_29872,N_29899);
nor UO_132 (O_132,N_29871,N_29979);
and UO_133 (O_133,N_29828,N_29973);
nand UO_134 (O_134,N_29876,N_29803);
nor UO_135 (O_135,N_29908,N_29924);
xnor UO_136 (O_136,N_29822,N_29849);
or UO_137 (O_137,N_29865,N_29889);
and UO_138 (O_138,N_29833,N_29991);
xnor UO_139 (O_139,N_29913,N_29845);
and UO_140 (O_140,N_29841,N_29869);
xor UO_141 (O_141,N_29976,N_29972);
and UO_142 (O_142,N_29997,N_29833);
and UO_143 (O_143,N_29833,N_29971);
nand UO_144 (O_144,N_29977,N_29817);
xnor UO_145 (O_145,N_29899,N_29844);
nor UO_146 (O_146,N_29828,N_29821);
or UO_147 (O_147,N_29935,N_29879);
xnor UO_148 (O_148,N_29911,N_29934);
and UO_149 (O_149,N_29839,N_29969);
nand UO_150 (O_150,N_29929,N_29867);
and UO_151 (O_151,N_29961,N_29841);
nand UO_152 (O_152,N_29868,N_29807);
or UO_153 (O_153,N_29980,N_29813);
and UO_154 (O_154,N_29931,N_29934);
nand UO_155 (O_155,N_29921,N_29969);
xnor UO_156 (O_156,N_29945,N_29933);
and UO_157 (O_157,N_29956,N_29861);
and UO_158 (O_158,N_29998,N_29931);
nand UO_159 (O_159,N_29981,N_29816);
nor UO_160 (O_160,N_29945,N_29826);
or UO_161 (O_161,N_29884,N_29870);
and UO_162 (O_162,N_29900,N_29804);
or UO_163 (O_163,N_29992,N_29983);
nand UO_164 (O_164,N_29869,N_29892);
nand UO_165 (O_165,N_29861,N_29800);
and UO_166 (O_166,N_29811,N_29861);
nand UO_167 (O_167,N_29804,N_29888);
and UO_168 (O_168,N_29938,N_29909);
and UO_169 (O_169,N_29924,N_29883);
and UO_170 (O_170,N_29934,N_29952);
or UO_171 (O_171,N_29822,N_29881);
nand UO_172 (O_172,N_29938,N_29995);
xnor UO_173 (O_173,N_29837,N_29968);
nand UO_174 (O_174,N_29812,N_29923);
xor UO_175 (O_175,N_29927,N_29857);
or UO_176 (O_176,N_29937,N_29900);
xnor UO_177 (O_177,N_29940,N_29824);
xor UO_178 (O_178,N_29981,N_29845);
and UO_179 (O_179,N_29988,N_29802);
or UO_180 (O_180,N_29820,N_29876);
or UO_181 (O_181,N_29840,N_29824);
nand UO_182 (O_182,N_29863,N_29824);
nand UO_183 (O_183,N_29816,N_29943);
nor UO_184 (O_184,N_29912,N_29985);
xor UO_185 (O_185,N_29852,N_29905);
and UO_186 (O_186,N_29982,N_29987);
nand UO_187 (O_187,N_29989,N_29856);
or UO_188 (O_188,N_29924,N_29948);
and UO_189 (O_189,N_29996,N_29935);
nand UO_190 (O_190,N_29932,N_29850);
or UO_191 (O_191,N_29889,N_29982);
nand UO_192 (O_192,N_29915,N_29913);
nor UO_193 (O_193,N_29988,N_29976);
nand UO_194 (O_194,N_29863,N_29956);
xnor UO_195 (O_195,N_29818,N_29895);
and UO_196 (O_196,N_29832,N_29959);
xor UO_197 (O_197,N_29889,N_29863);
and UO_198 (O_198,N_29888,N_29975);
and UO_199 (O_199,N_29890,N_29913);
and UO_200 (O_200,N_29915,N_29819);
nand UO_201 (O_201,N_29821,N_29839);
nor UO_202 (O_202,N_29887,N_29853);
nor UO_203 (O_203,N_29860,N_29818);
or UO_204 (O_204,N_29885,N_29927);
and UO_205 (O_205,N_29828,N_29917);
nor UO_206 (O_206,N_29991,N_29863);
nor UO_207 (O_207,N_29827,N_29849);
and UO_208 (O_208,N_29850,N_29816);
or UO_209 (O_209,N_29928,N_29925);
and UO_210 (O_210,N_29915,N_29846);
nand UO_211 (O_211,N_29911,N_29983);
nor UO_212 (O_212,N_29873,N_29965);
xnor UO_213 (O_213,N_29919,N_29893);
xor UO_214 (O_214,N_29978,N_29860);
xnor UO_215 (O_215,N_29978,N_29832);
xor UO_216 (O_216,N_29825,N_29849);
nand UO_217 (O_217,N_29808,N_29956);
and UO_218 (O_218,N_29937,N_29814);
nor UO_219 (O_219,N_29822,N_29858);
nor UO_220 (O_220,N_29940,N_29876);
nand UO_221 (O_221,N_29948,N_29926);
xor UO_222 (O_222,N_29997,N_29967);
nand UO_223 (O_223,N_29832,N_29857);
nand UO_224 (O_224,N_29820,N_29871);
xnor UO_225 (O_225,N_29890,N_29951);
nor UO_226 (O_226,N_29949,N_29894);
xnor UO_227 (O_227,N_29842,N_29949);
xnor UO_228 (O_228,N_29819,N_29989);
or UO_229 (O_229,N_29950,N_29919);
nor UO_230 (O_230,N_29915,N_29805);
or UO_231 (O_231,N_29958,N_29935);
or UO_232 (O_232,N_29951,N_29820);
or UO_233 (O_233,N_29867,N_29885);
nor UO_234 (O_234,N_29810,N_29845);
xnor UO_235 (O_235,N_29955,N_29971);
nand UO_236 (O_236,N_29954,N_29873);
nor UO_237 (O_237,N_29814,N_29976);
nor UO_238 (O_238,N_29894,N_29904);
nor UO_239 (O_239,N_29916,N_29849);
and UO_240 (O_240,N_29855,N_29888);
and UO_241 (O_241,N_29962,N_29931);
xnor UO_242 (O_242,N_29968,N_29962);
and UO_243 (O_243,N_29833,N_29863);
xor UO_244 (O_244,N_29965,N_29845);
and UO_245 (O_245,N_29802,N_29977);
nand UO_246 (O_246,N_29978,N_29900);
xnor UO_247 (O_247,N_29912,N_29953);
xnor UO_248 (O_248,N_29913,N_29920);
nor UO_249 (O_249,N_29925,N_29862);
xor UO_250 (O_250,N_29850,N_29826);
or UO_251 (O_251,N_29815,N_29899);
nand UO_252 (O_252,N_29905,N_29912);
xor UO_253 (O_253,N_29832,N_29943);
xor UO_254 (O_254,N_29934,N_29893);
nand UO_255 (O_255,N_29987,N_29802);
or UO_256 (O_256,N_29901,N_29857);
nand UO_257 (O_257,N_29961,N_29804);
and UO_258 (O_258,N_29943,N_29801);
or UO_259 (O_259,N_29991,N_29868);
or UO_260 (O_260,N_29984,N_29967);
or UO_261 (O_261,N_29925,N_29926);
or UO_262 (O_262,N_29811,N_29821);
nand UO_263 (O_263,N_29908,N_29905);
and UO_264 (O_264,N_29809,N_29855);
nand UO_265 (O_265,N_29990,N_29957);
xor UO_266 (O_266,N_29973,N_29852);
and UO_267 (O_267,N_29809,N_29916);
and UO_268 (O_268,N_29987,N_29874);
and UO_269 (O_269,N_29900,N_29820);
xnor UO_270 (O_270,N_29894,N_29884);
nor UO_271 (O_271,N_29919,N_29925);
or UO_272 (O_272,N_29958,N_29952);
nor UO_273 (O_273,N_29882,N_29990);
nand UO_274 (O_274,N_29834,N_29904);
xor UO_275 (O_275,N_29892,N_29917);
and UO_276 (O_276,N_29918,N_29935);
nor UO_277 (O_277,N_29901,N_29882);
and UO_278 (O_278,N_29956,N_29920);
and UO_279 (O_279,N_29977,N_29911);
nand UO_280 (O_280,N_29874,N_29918);
nand UO_281 (O_281,N_29967,N_29900);
and UO_282 (O_282,N_29816,N_29980);
nand UO_283 (O_283,N_29840,N_29957);
xnor UO_284 (O_284,N_29945,N_29978);
nand UO_285 (O_285,N_29859,N_29855);
and UO_286 (O_286,N_29915,N_29878);
xnor UO_287 (O_287,N_29836,N_29971);
or UO_288 (O_288,N_29890,N_29933);
xor UO_289 (O_289,N_29870,N_29876);
and UO_290 (O_290,N_29934,N_29950);
nand UO_291 (O_291,N_29817,N_29970);
xnor UO_292 (O_292,N_29950,N_29984);
and UO_293 (O_293,N_29899,N_29910);
xor UO_294 (O_294,N_29813,N_29899);
nor UO_295 (O_295,N_29896,N_29800);
or UO_296 (O_296,N_29906,N_29965);
or UO_297 (O_297,N_29891,N_29832);
nor UO_298 (O_298,N_29975,N_29908);
nor UO_299 (O_299,N_29830,N_29935);
xnor UO_300 (O_300,N_29971,N_29998);
nand UO_301 (O_301,N_29865,N_29966);
and UO_302 (O_302,N_29913,N_29953);
nor UO_303 (O_303,N_29836,N_29901);
nor UO_304 (O_304,N_29816,N_29868);
nand UO_305 (O_305,N_29999,N_29875);
or UO_306 (O_306,N_29983,N_29979);
nor UO_307 (O_307,N_29822,N_29831);
nor UO_308 (O_308,N_29943,N_29846);
and UO_309 (O_309,N_29972,N_29954);
nor UO_310 (O_310,N_29819,N_29895);
and UO_311 (O_311,N_29934,N_29844);
nand UO_312 (O_312,N_29932,N_29967);
nor UO_313 (O_313,N_29812,N_29994);
or UO_314 (O_314,N_29892,N_29916);
xor UO_315 (O_315,N_29968,N_29812);
xor UO_316 (O_316,N_29986,N_29951);
and UO_317 (O_317,N_29908,N_29872);
nor UO_318 (O_318,N_29990,N_29803);
or UO_319 (O_319,N_29865,N_29890);
xor UO_320 (O_320,N_29896,N_29905);
nand UO_321 (O_321,N_29930,N_29827);
and UO_322 (O_322,N_29958,N_29807);
nor UO_323 (O_323,N_29982,N_29955);
xor UO_324 (O_324,N_29913,N_29891);
or UO_325 (O_325,N_29950,N_29829);
or UO_326 (O_326,N_29857,N_29844);
or UO_327 (O_327,N_29811,N_29855);
or UO_328 (O_328,N_29876,N_29969);
and UO_329 (O_329,N_29843,N_29953);
nor UO_330 (O_330,N_29961,N_29971);
nor UO_331 (O_331,N_29808,N_29830);
xor UO_332 (O_332,N_29935,N_29817);
nand UO_333 (O_333,N_29972,N_29894);
or UO_334 (O_334,N_29907,N_29942);
nand UO_335 (O_335,N_29984,N_29811);
nor UO_336 (O_336,N_29903,N_29872);
nand UO_337 (O_337,N_29882,N_29974);
nand UO_338 (O_338,N_29971,N_29917);
xor UO_339 (O_339,N_29889,N_29997);
or UO_340 (O_340,N_29958,N_29943);
nor UO_341 (O_341,N_29989,N_29913);
nor UO_342 (O_342,N_29843,N_29946);
nor UO_343 (O_343,N_29883,N_29877);
or UO_344 (O_344,N_29865,N_29841);
and UO_345 (O_345,N_29985,N_29989);
nand UO_346 (O_346,N_29851,N_29981);
nor UO_347 (O_347,N_29997,N_29919);
nor UO_348 (O_348,N_29855,N_29822);
nand UO_349 (O_349,N_29839,N_29987);
and UO_350 (O_350,N_29992,N_29926);
or UO_351 (O_351,N_29933,N_29966);
or UO_352 (O_352,N_29818,N_29901);
nor UO_353 (O_353,N_29870,N_29921);
and UO_354 (O_354,N_29881,N_29993);
nand UO_355 (O_355,N_29912,N_29831);
xnor UO_356 (O_356,N_29869,N_29950);
nand UO_357 (O_357,N_29978,N_29851);
and UO_358 (O_358,N_29858,N_29961);
and UO_359 (O_359,N_29841,N_29978);
nor UO_360 (O_360,N_29928,N_29800);
and UO_361 (O_361,N_29970,N_29829);
nor UO_362 (O_362,N_29944,N_29962);
and UO_363 (O_363,N_29886,N_29967);
nor UO_364 (O_364,N_29962,N_29829);
or UO_365 (O_365,N_29883,N_29825);
nor UO_366 (O_366,N_29826,N_29868);
and UO_367 (O_367,N_29960,N_29970);
nor UO_368 (O_368,N_29852,N_29894);
or UO_369 (O_369,N_29819,N_29822);
nand UO_370 (O_370,N_29932,N_29939);
or UO_371 (O_371,N_29989,N_29800);
nor UO_372 (O_372,N_29930,N_29893);
nand UO_373 (O_373,N_29978,N_29948);
nor UO_374 (O_374,N_29991,N_29809);
or UO_375 (O_375,N_29972,N_29855);
xnor UO_376 (O_376,N_29888,N_29856);
or UO_377 (O_377,N_29826,N_29831);
or UO_378 (O_378,N_29835,N_29957);
xnor UO_379 (O_379,N_29952,N_29966);
nand UO_380 (O_380,N_29804,N_29997);
or UO_381 (O_381,N_29994,N_29888);
nor UO_382 (O_382,N_29929,N_29914);
and UO_383 (O_383,N_29866,N_29883);
nor UO_384 (O_384,N_29814,N_29929);
nor UO_385 (O_385,N_29829,N_29999);
or UO_386 (O_386,N_29886,N_29828);
or UO_387 (O_387,N_29904,N_29966);
or UO_388 (O_388,N_29993,N_29982);
or UO_389 (O_389,N_29920,N_29970);
nand UO_390 (O_390,N_29969,N_29992);
xor UO_391 (O_391,N_29956,N_29833);
nand UO_392 (O_392,N_29872,N_29995);
and UO_393 (O_393,N_29929,N_29934);
and UO_394 (O_394,N_29826,N_29962);
nor UO_395 (O_395,N_29991,N_29931);
nand UO_396 (O_396,N_29845,N_29945);
xnor UO_397 (O_397,N_29852,N_29899);
xor UO_398 (O_398,N_29939,N_29991);
and UO_399 (O_399,N_29901,N_29881);
nor UO_400 (O_400,N_29892,N_29843);
or UO_401 (O_401,N_29909,N_29890);
or UO_402 (O_402,N_29905,N_29963);
or UO_403 (O_403,N_29948,N_29808);
nor UO_404 (O_404,N_29852,N_29924);
and UO_405 (O_405,N_29932,N_29893);
or UO_406 (O_406,N_29943,N_29859);
or UO_407 (O_407,N_29922,N_29905);
xor UO_408 (O_408,N_29810,N_29801);
or UO_409 (O_409,N_29901,N_29848);
nand UO_410 (O_410,N_29872,N_29948);
nor UO_411 (O_411,N_29848,N_29892);
xor UO_412 (O_412,N_29901,N_29811);
xor UO_413 (O_413,N_29861,N_29846);
or UO_414 (O_414,N_29992,N_29950);
nor UO_415 (O_415,N_29846,N_29869);
and UO_416 (O_416,N_29984,N_29898);
and UO_417 (O_417,N_29858,N_29906);
and UO_418 (O_418,N_29858,N_29879);
nand UO_419 (O_419,N_29880,N_29890);
xnor UO_420 (O_420,N_29974,N_29918);
nor UO_421 (O_421,N_29909,N_29817);
nand UO_422 (O_422,N_29852,N_29831);
xor UO_423 (O_423,N_29944,N_29852);
nor UO_424 (O_424,N_29800,N_29929);
nand UO_425 (O_425,N_29989,N_29994);
nand UO_426 (O_426,N_29995,N_29900);
or UO_427 (O_427,N_29921,N_29985);
xor UO_428 (O_428,N_29910,N_29952);
nor UO_429 (O_429,N_29952,N_29858);
nor UO_430 (O_430,N_29913,N_29812);
nand UO_431 (O_431,N_29833,N_29847);
nor UO_432 (O_432,N_29947,N_29961);
nor UO_433 (O_433,N_29859,N_29937);
xnor UO_434 (O_434,N_29961,N_29808);
nand UO_435 (O_435,N_29877,N_29985);
nand UO_436 (O_436,N_29882,N_29820);
nand UO_437 (O_437,N_29894,N_29845);
xor UO_438 (O_438,N_29874,N_29948);
nor UO_439 (O_439,N_29883,N_29824);
and UO_440 (O_440,N_29838,N_29981);
and UO_441 (O_441,N_29924,N_29941);
or UO_442 (O_442,N_29959,N_29960);
xor UO_443 (O_443,N_29974,N_29842);
nand UO_444 (O_444,N_29887,N_29831);
xnor UO_445 (O_445,N_29902,N_29955);
nor UO_446 (O_446,N_29819,N_29839);
or UO_447 (O_447,N_29949,N_29911);
nor UO_448 (O_448,N_29862,N_29908);
xnor UO_449 (O_449,N_29861,N_29943);
nor UO_450 (O_450,N_29953,N_29965);
and UO_451 (O_451,N_29970,N_29812);
nor UO_452 (O_452,N_29886,N_29822);
nand UO_453 (O_453,N_29944,N_29874);
nand UO_454 (O_454,N_29988,N_29800);
or UO_455 (O_455,N_29901,N_29802);
or UO_456 (O_456,N_29867,N_29976);
or UO_457 (O_457,N_29813,N_29961);
and UO_458 (O_458,N_29842,N_29939);
or UO_459 (O_459,N_29862,N_29928);
nor UO_460 (O_460,N_29871,N_29903);
nor UO_461 (O_461,N_29866,N_29893);
xor UO_462 (O_462,N_29907,N_29852);
nor UO_463 (O_463,N_29972,N_29813);
and UO_464 (O_464,N_29966,N_29853);
nand UO_465 (O_465,N_29968,N_29806);
or UO_466 (O_466,N_29834,N_29956);
or UO_467 (O_467,N_29911,N_29987);
and UO_468 (O_468,N_29876,N_29827);
xnor UO_469 (O_469,N_29900,N_29851);
nand UO_470 (O_470,N_29954,N_29919);
xnor UO_471 (O_471,N_29880,N_29904);
or UO_472 (O_472,N_29884,N_29935);
nand UO_473 (O_473,N_29830,N_29960);
nor UO_474 (O_474,N_29907,N_29929);
xnor UO_475 (O_475,N_29914,N_29948);
and UO_476 (O_476,N_29812,N_29884);
nand UO_477 (O_477,N_29935,N_29913);
or UO_478 (O_478,N_29959,N_29930);
nor UO_479 (O_479,N_29954,N_29854);
nor UO_480 (O_480,N_29801,N_29938);
or UO_481 (O_481,N_29965,N_29920);
nand UO_482 (O_482,N_29807,N_29806);
xor UO_483 (O_483,N_29962,N_29927);
and UO_484 (O_484,N_29893,N_29857);
nand UO_485 (O_485,N_29819,N_29807);
and UO_486 (O_486,N_29951,N_29834);
and UO_487 (O_487,N_29942,N_29962);
and UO_488 (O_488,N_29903,N_29907);
and UO_489 (O_489,N_29817,N_29991);
nor UO_490 (O_490,N_29837,N_29907);
xnor UO_491 (O_491,N_29904,N_29871);
nand UO_492 (O_492,N_29959,N_29880);
and UO_493 (O_493,N_29876,N_29999);
nor UO_494 (O_494,N_29840,N_29944);
xor UO_495 (O_495,N_29975,N_29964);
or UO_496 (O_496,N_29907,N_29876);
xor UO_497 (O_497,N_29901,N_29911);
xor UO_498 (O_498,N_29812,N_29881);
nand UO_499 (O_499,N_29879,N_29918);
nor UO_500 (O_500,N_29920,N_29906);
and UO_501 (O_501,N_29997,N_29871);
nand UO_502 (O_502,N_29848,N_29889);
and UO_503 (O_503,N_29991,N_29906);
xnor UO_504 (O_504,N_29867,N_29891);
nor UO_505 (O_505,N_29983,N_29891);
or UO_506 (O_506,N_29955,N_29944);
xnor UO_507 (O_507,N_29886,N_29880);
nand UO_508 (O_508,N_29995,N_29844);
or UO_509 (O_509,N_29837,N_29823);
nand UO_510 (O_510,N_29877,N_29976);
xor UO_511 (O_511,N_29807,N_29838);
xnor UO_512 (O_512,N_29871,N_29916);
or UO_513 (O_513,N_29874,N_29805);
nor UO_514 (O_514,N_29968,N_29924);
or UO_515 (O_515,N_29872,N_29936);
nor UO_516 (O_516,N_29883,N_29959);
xor UO_517 (O_517,N_29967,N_29888);
xor UO_518 (O_518,N_29871,N_29989);
or UO_519 (O_519,N_29927,N_29979);
nand UO_520 (O_520,N_29866,N_29836);
and UO_521 (O_521,N_29938,N_29866);
xnor UO_522 (O_522,N_29815,N_29935);
or UO_523 (O_523,N_29928,N_29932);
and UO_524 (O_524,N_29805,N_29925);
nand UO_525 (O_525,N_29930,N_29868);
and UO_526 (O_526,N_29932,N_29979);
and UO_527 (O_527,N_29864,N_29938);
nand UO_528 (O_528,N_29908,N_29857);
xnor UO_529 (O_529,N_29896,N_29960);
or UO_530 (O_530,N_29946,N_29889);
xnor UO_531 (O_531,N_29843,N_29924);
xor UO_532 (O_532,N_29863,N_29958);
xor UO_533 (O_533,N_29944,N_29986);
or UO_534 (O_534,N_29853,N_29861);
xor UO_535 (O_535,N_29880,N_29841);
nor UO_536 (O_536,N_29861,N_29881);
nand UO_537 (O_537,N_29914,N_29879);
nor UO_538 (O_538,N_29855,N_29812);
and UO_539 (O_539,N_29955,N_29975);
or UO_540 (O_540,N_29815,N_29986);
and UO_541 (O_541,N_29954,N_29978);
nand UO_542 (O_542,N_29886,N_29864);
nand UO_543 (O_543,N_29948,N_29935);
and UO_544 (O_544,N_29835,N_29812);
xnor UO_545 (O_545,N_29872,N_29847);
or UO_546 (O_546,N_29953,N_29859);
nand UO_547 (O_547,N_29947,N_29825);
and UO_548 (O_548,N_29804,N_29845);
and UO_549 (O_549,N_29926,N_29863);
nor UO_550 (O_550,N_29904,N_29997);
and UO_551 (O_551,N_29886,N_29830);
and UO_552 (O_552,N_29988,N_29952);
nor UO_553 (O_553,N_29879,N_29852);
xor UO_554 (O_554,N_29983,N_29845);
nand UO_555 (O_555,N_29950,N_29852);
nand UO_556 (O_556,N_29982,N_29811);
or UO_557 (O_557,N_29878,N_29985);
and UO_558 (O_558,N_29870,N_29888);
or UO_559 (O_559,N_29897,N_29903);
or UO_560 (O_560,N_29962,N_29869);
nand UO_561 (O_561,N_29905,N_29998);
nand UO_562 (O_562,N_29984,N_29851);
nor UO_563 (O_563,N_29909,N_29956);
nor UO_564 (O_564,N_29809,N_29962);
or UO_565 (O_565,N_29870,N_29922);
xor UO_566 (O_566,N_29944,N_29869);
nand UO_567 (O_567,N_29934,N_29921);
nor UO_568 (O_568,N_29943,N_29945);
xor UO_569 (O_569,N_29960,N_29805);
nand UO_570 (O_570,N_29859,N_29983);
or UO_571 (O_571,N_29833,N_29806);
xnor UO_572 (O_572,N_29867,N_29945);
and UO_573 (O_573,N_29815,N_29853);
and UO_574 (O_574,N_29946,N_29832);
and UO_575 (O_575,N_29958,N_29918);
xor UO_576 (O_576,N_29890,N_29939);
or UO_577 (O_577,N_29984,N_29943);
nand UO_578 (O_578,N_29835,N_29858);
xnor UO_579 (O_579,N_29818,N_29997);
and UO_580 (O_580,N_29973,N_29893);
nand UO_581 (O_581,N_29952,N_29950);
and UO_582 (O_582,N_29813,N_29883);
nand UO_583 (O_583,N_29887,N_29977);
and UO_584 (O_584,N_29884,N_29819);
and UO_585 (O_585,N_29814,N_29849);
nor UO_586 (O_586,N_29915,N_29916);
nand UO_587 (O_587,N_29947,N_29950);
nand UO_588 (O_588,N_29884,N_29942);
nand UO_589 (O_589,N_29842,N_29957);
xnor UO_590 (O_590,N_29908,N_29911);
xnor UO_591 (O_591,N_29859,N_29964);
nor UO_592 (O_592,N_29971,N_29923);
nand UO_593 (O_593,N_29886,N_29867);
or UO_594 (O_594,N_29841,N_29997);
xnor UO_595 (O_595,N_29816,N_29865);
or UO_596 (O_596,N_29814,N_29963);
xnor UO_597 (O_597,N_29838,N_29987);
and UO_598 (O_598,N_29827,N_29895);
or UO_599 (O_599,N_29886,N_29978);
nor UO_600 (O_600,N_29845,N_29811);
and UO_601 (O_601,N_29882,N_29996);
and UO_602 (O_602,N_29866,N_29903);
nand UO_603 (O_603,N_29851,N_29926);
nand UO_604 (O_604,N_29881,N_29949);
and UO_605 (O_605,N_29991,N_29952);
nor UO_606 (O_606,N_29983,N_29972);
and UO_607 (O_607,N_29976,N_29986);
nor UO_608 (O_608,N_29813,N_29827);
xor UO_609 (O_609,N_29826,N_29977);
and UO_610 (O_610,N_29971,N_29989);
xor UO_611 (O_611,N_29822,N_29974);
nand UO_612 (O_612,N_29997,N_29875);
xnor UO_613 (O_613,N_29966,N_29925);
or UO_614 (O_614,N_29942,N_29802);
nand UO_615 (O_615,N_29920,N_29916);
xnor UO_616 (O_616,N_29828,N_29809);
and UO_617 (O_617,N_29899,N_29893);
or UO_618 (O_618,N_29948,N_29830);
nor UO_619 (O_619,N_29816,N_29883);
xnor UO_620 (O_620,N_29970,N_29901);
xor UO_621 (O_621,N_29812,N_29897);
nor UO_622 (O_622,N_29975,N_29813);
nand UO_623 (O_623,N_29855,N_29979);
nand UO_624 (O_624,N_29870,N_29926);
xnor UO_625 (O_625,N_29971,N_29991);
nor UO_626 (O_626,N_29808,N_29926);
nand UO_627 (O_627,N_29964,N_29831);
nand UO_628 (O_628,N_29862,N_29868);
or UO_629 (O_629,N_29820,N_29969);
and UO_630 (O_630,N_29856,N_29886);
nand UO_631 (O_631,N_29854,N_29941);
and UO_632 (O_632,N_29885,N_29926);
xnor UO_633 (O_633,N_29930,N_29889);
nor UO_634 (O_634,N_29981,N_29992);
nor UO_635 (O_635,N_29854,N_29875);
nor UO_636 (O_636,N_29903,N_29804);
nand UO_637 (O_637,N_29947,N_29915);
nand UO_638 (O_638,N_29832,N_29869);
nand UO_639 (O_639,N_29809,N_29903);
or UO_640 (O_640,N_29844,N_29944);
xor UO_641 (O_641,N_29926,N_29967);
nand UO_642 (O_642,N_29815,N_29817);
nor UO_643 (O_643,N_29998,N_29847);
and UO_644 (O_644,N_29995,N_29829);
nor UO_645 (O_645,N_29991,N_29978);
or UO_646 (O_646,N_29943,N_29916);
xor UO_647 (O_647,N_29898,N_29975);
and UO_648 (O_648,N_29861,N_29831);
and UO_649 (O_649,N_29898,N_29801);
xor UO_650 (O_650,N_29850,N_29975);
and UO_651 (O_651,N_29814,N_29919);
xnor UO_652 (O_652,N_29844,N_29809);
or UO_653 (O_653,N_29887,N_29961);
nor UO_654 (O_654,N_29804,N_29919);
nand UO_655 (O_655,N_29873,N_29929);
and UO_656 (O_656,N_29808,N_29807);
or UO_657 (O_657,N_29980,N_29845);
and UO_658 (O_658,N_29866,N_29954);
xnor UO_659 (O_659,N_29921,N_29882);
nand UO_660 (O_660,N_29986,N_29854);
or UO_661 (O_661,N_29930,N_29821);
nor UO_662 (O_662,N_29944,N_29984);
nor UO_663 (O_663,N_29800,N_29824);
or UO_664 (O_664,N_29913,N_29836);
or UO_665 (O_665,N_29894,N_29878);
or UO_666 (O_666,N_29868,N_29808);
and UO_667 (O_667,N_29908,N_29825);
nand UO_668 (O_668,N_29889,N_29937);
nand UO_669 (O_669,N_29860,N_29835);
and UO_670 (O_670,N_29978,N_29867);
xor UO_671 (O_671,N_29925,N_29898);
and UO_672 (O_672,N_29810,N_29822);
nand UO_673 (O_673,N_29966,N_29982);
nand UO_674 (O_674,N_29986,N_29969);
nand UO_675 (O_675,N_29893,N_29812);
nor UO_676 (O_676,N_29904,N_29802);
xor UO_677 (O_677,N_29927,N_29894);
xnor UO_678 (O_678,N_29923,N_29879);
and UO_679 (O_679,N_29981,N_29805);
nor UO_680 (O_680,N_29994,N_29964);
or UO_681 (O_681,N_29844,N_29866);
nand UO_682 (O_682,N_29921,N_29806);
nor UO_683 (O_683,N_29917,N_29841);
nand UO_684 (O_684,N_29820,N_29832);
or UO_685 (O_685,N_29957,N_29864);
xnor UO_686 (O_686,N_29919,N_29985);
and UO_687 (O_687,N_29995,N_29834);
nor UO_688 (O_688,N_29849,N_29800);
xor UO_689 (O_689,N_29819,N_29850);
nor UO_690 (O_690,N_29994,N_29810);
xor UO_691 (O_691,N_29985,N_29869);
nand UO_692 (O_692,N_29940,N_29829);
nor UO_693 (O_693,N_29918,N_29813);
xor UO_694 (O_694,N_29858,N_29892);
nor UO_695 (O_695,N_29976,N_29941);
and UO_696 (O_696,N_29874,N_29863);
nor UO_697 (O_697,N_29847,N_29862);
or UO_698 (O_698,N_29841,N_29899);
and UO_699 (O_699,N_29824,N_29853);
nor UO_700 (O_700,N_29809,N_29802);
nor UO_701 (O_701,N_29992,N_29961);
or UO_702 (O_702,N_29938,N_29851);
or UO_703 (O_703,N_29988,N_29978);
nand UO_704 (O_704,N_29906,N_29899);
xnor UO_705 (O_705,N_29994,N_29976);
xor UO_706 (O_706,N_29965,N_29927);
nor UO_707 (O_707,N_29986,N_29899);
and UO_708 (O_708,N_29980,N_29825);
nand UO_709 (O_709,N_29961,N_29881);
nor UO_710 (O_710,N_29895,N_29930);
and UO_711 (O_711,N_29938,N_29894);
or UO_712 (O_712,N_29999,N_29868);
nand UO_713 (O_713,N_29971,N_29893);
nor UO_714 (O_714,N_29838,N_29937);
nand UO_715 (O_715,N_29877,N_29910);
and UO_716 (O_716,N_29966,N_29942);
or UO_717 (O_717,N_29805,N_29802);
nor UO_718 (O_718,N_29929,N_29865);
and UO_719 (O_719,N_29910,N_29941);
and UO_720 (O_720,N_29865,N_29898);
and UO_721 (O_721,N_29901,N_29923);
or UO_722 (O_722,N_29921,N_29912);
xor UO_723 (O_723,N_29984,N_29895);
nand UO_724 (O_724,N_29966,N_29990);
or UO_725 (O_725,N_29930,N_29852);
xor UO_726 (O_726,N_29884,N_29930);
and UO_727 (O_727,N_29927,N_29818);
or UO_728 (O_728,N_29981,N_29841);
and UO_729 (O_729,N_29870,N_29872);
xnor UO_730 (O_730,N_29819,N_29928);
nand UO_731 (O_731,N_29940,N_29862);
nand UO_732 (O_732,N_29979,N_29948);
nor UO_733 (O_733,N_29847,N_29897);
xor UO_734 (O_734,N_29809,N_29803);
or UO_735 (O_735,N_29864,N_29878);
and UO_736 (O_736,N_29829,N_29913);
nand UO_737 (O_737,N_29831,N_29950);
and UO_738 (O_738,N_29857,N_29905);
and UO_739 (O_739,N_29908,N_29832);
xor UO_740 (O_740,N_29894,N_29955);
nor UO_741 (O_741,N_29989,N_29925);
or UO_742 (O_742,N_29892,N_29835);
nor UO_743 (O_743,N_29899,N_29905);
nor UO_744 (O_744,N_29873,N_29979);
xor UO_745 (O_745,N_29910,N_29923);
nand UO_746 (O_746,N_29937,N_29977);
and UO_747 (O_747,N_29803,N_29933);
or UO_748 (O_748,N_29855,N_29827);
nor UO_749 (O_749,N_29863,N_29808);
xnor UO_750 (O_750,N_29943,N_29820);
or UO_751 (O_751,N_29981,N_29846);
or UO_752 (O_752,N_29823,N_29839);
nor UO_753 (O_753,N_29977,N_29984);
and UO_754 (O_754,N_29979,N_29978);
nor UO_755 (O_755,N_29815,N_29891);
and UO_756 (O_756,N_29980,N_29873);
and UO_757 (O_757,N_29802,N_29806);
and UO_758 (O_758,N_29883,N_29827);
xnor UO_759 (O_759,N_29813,N_29998);
and UO_760 (O_760,N_29917,N_29887);
nor UO_761 (O_761,N_29859,N_29826);
xor UO_762 (O_762,N_29975,N_29917);
and UO_763 (O_763,N_29945,N_29926);
or UO_764 (O_764,N_29976,N_29843);
nor UO_765 (O_765,N_29974,N_29969);
xor UO_766 (O_766,N_29872,N_29881);
nand UO_767 (O_767,N_29910,N_29844);
or UO_768 (O_768,N_29883,N_29876);
or UO_769 (O_769,N_29960,N_29808);
and UO_770 (O_770,N_29898,N_29828);
nor UO_771 (O_771,N_29811,N_29862);
or UO_772 (O_772,N_29878,N_29811);
nor UO_773 (O_773,N_29894,N_29828);
xnor UO_774 (O_774,N_29965,N_29801);
nor UO_775 (O_775,N_29813,N_29877);
or UO_776 (O_776,N_29970,N_29921);
and UO_777 (O_777,N_29948,N_29873);
xor UO_778 (O_778,N_29953,N_29944);
xor UO_779 (O_779,N_29954,N_29922);
and UO_780 (O_780,N_29831,N_29993);
xnor UO_781 (O_781,N_29935,N_29896);
nor UO_782 (O_782,N_29921,N_29800);
and UO_783 (O_783,N_29993,N_29926);
and UO_784 (O_784,N_29824,N_29911);
and UO_785 (O_785,N_29862,N_29971);
nor UO_786 (O_786,N_29894,N_29853);
and UO_787 (O_787,N_29823,N_29894);
nand UO_788 (O_788,N_29876,N_29802);
nor UO_789 (O_789,N_29847,N_29952);
xor UO_790 (O_790,N_29853,N_29895);
or UO_791 (O_791,N_29823,N_29915);
nor UO_792 (O_792,N_29985,N_29900);
nor UO_793 (O_793,N_29966,N_29947);
nor UO_794 (O_794,N_29838,N_29887);
nor UO_795 (O_795,N_29962,N_29833);
xnor UO_796 (O_796,N_29906,N_29987);
or UO_797 (O_797,N_29926,N_29957);
nor UO_798 (O_798,N_29874,N_29862);
xor UO_799 (O_799,N_29907,N_29800);
nor UO_800 (O_800,N_29919,N_29972);
xnor UO_801 (O_801,N_29939,N_29848);
xnor UO_802 (O_802,N_29889,N_29942);
nor UO_803 (O_803,N_29871,N_29848);
nor UO_804 (O_804,N_29896,N_29915);
and UO_805 (O_805,N_29873,N_29897);
or UO_806 (O_806,N_29937,N_29846);
and UO_807 (O_807,N_29916,N_29940);
nand UO_808 (O_808,N_29946,N_29943);
or UO_809 (O_809,N_29941,N_29871);
xor UO_810 (O_810,N_29910,N_29800);
or UO_811 (O_811,N_29811,N_29931);
nand UO_812 (O_812,N_29918,N_29952);
and UO_813 (O_813,N_29948,N_29919);
nor UO_814 (O_814,N_29881,N_29946);
nor UO_815 (O_815,N_29807,N_29877);
nor UO_816 (O_816,N_29899,N_29801);
xor UO_817 (O_817,N_29933,N_29969);
nor UO_818 (O_818,N_29898,N_29818);
xor UO_819 (O_819,N_29974,N_29959);
and UO_820 (O_820,N_29989,N_29810);
nor UO_821 (O_821,N_29812,N_29940);
nor UO_822 (O_822,N_29963,N_29853);
and UO_823 (O_823,N_29829,N_29907);
xnor UO_824 (O_824,N_29873,N_29937);
nor UO_825 (O_825,N_29848,N_29961);
nand UO_826 (O_826,N_29894,N_29959);
nand UO_827 (O_827,N_29801,N_29811);
xnor UO_828 (O_828,N_29996,N_29801);
and UO_829 (O_829,N_29904,N_29867);
and UO_830 (O_830,N_29862,N_29954);
nand UO_831 (O_831,N_29971,N_29802);
and UO_832 (O_832,N_29858,N_29937);
nand UO_833 (O_833,N_29848,N_29817);
xnor UO_834 (O_834,N_29971,N_29981);
or UO_835 (O_835,N_29821,N_29872);
xnor UO_836 (O_836,N_29878,N_29908);
nand UO_837 (O_837,N_29855,N_29807);
nor UO_838 (O_838,N_29847,N_29829);
or UO_839 (O_839,N_29814,N_29911);
xnor UO_840 (O_840,N_29880,N_29905);
and UO_841 (O_841,N_29946,N_29863);
nand UO_842 (O_842,N_29843,N_29826);
and UO_843 (O_843,N_29915,N_29857);
and UO_844 (O_844,N_29908,N_29926);
nor UO_845 (O_845,N_29942,N_29891);
or UO_846 (O_846,N_29826,N_29905);
nand UO_847 (O_847,N_29828,N_29876);
nor UO_848 (O_848,N_29891,N_29934);
xnor UO_849 (O_849,N_29962,N_29872);
nand UO_850 (O_850,N_29933,N_29823);
or UO_851 (O_851,N_29871,N_29867);
and UO_852 (O_852,N_29848,N_29927);
or UO_853 (O_853,N_29928,N_29846);
or UO_854 (O_854,N_29814,N_29872);
nand UO_855 (O_855,N_29975,N_29895);
and UO_856 (O_856,N_29910,N_29845);
xnor UO_857 (O_857,N_29815,N_29844);
nand UO_858 (O_858,N_29838,N_29897);
nand UO_859 (O_859,N_29873,N_29826);
nand UO_860 (O_860,N_29831,N_29844);
or UO_861 (O_861,N_29912,N_29859);
xnor UO_862 (O_862,N_29976,N_29974);
nand UO_863 (O_863,N_29961,N_29812);
or UO_864 (O_864,N_29981,N_29907);
nand UO_865 (O_865,N_29832,N_29997);
nor UO_866 (O_866,N_29984,N_29841);
nand UO_867 (O_867,N_29835,N_29946);
nor UO_868 (O_868,N_29872,N_29836);
nand UO_869 (O_869,N_29854,N_29882);
or UO_870 (O_870,N_29803,N_29935);
and UO_871 (O_871,N_29959,N_29829);
and UO_872 (O_872,N_29819,N_29971);
or UO_873 (O_873,N_29909,N_29953);
nor UO_874 (O_874,N_29962,N_29989);
or UO_875 (O_875,N_29953,N_29808);
nand UO_876 (O_876,N_29903,N_29913);
nand UO_877 (O_877,N_29991,N_29853);
or UO_878 (O_878,N_29936,N_29879);
and UO_879 (O_879,N_29822,N_29857);
xor UO_880 (O_880,N_29907,N_29922);
nor UO_881 (O_881,N_29876,N_29986);
nor UO_882 (O_882,N_29972,N_29844);
xor UO_883 (O_883,N_29899,N_29869);
xnor UO_884 (O_884,N_29885,N_29879);
xnor UO_885 (O_885,N_29896,N_29866);
xnor UO_886 (O_886,N_29993,N_29920);
and UO_887 (O_887,N_29989,N_29934);
xor UO_888 (O_888,N_29989,N_29883);
xnor UO_889 (O_889,N_29956,N_29896);
nor UO_890 (O_890,N_29876,N_29908);
xor UO_891 (O_891,N_29873,N_29909);
and UO_892 (O_892,N_29945,N_29823);
or UO_893 (O_893,N_29998,N_29936);
or UO_894 (O_894,N_29802,N_29867);
nor UO_895 (O_895,N_29826,N_29885);
nor UO_896 (O_896,N_29893,N_29900);
or UO_897 (O_897,N_29936,N_29980);
nand UO_898 (O_898,N_29859,N_29889);
xor UO_899 (O_899,N_29830,N_29993);
nor UO_900 (O_900,N_29829,N_29947);
or UO_901 (O_901,N_29814,N_29884);
nand UO_902 (O_902,N_29821,N_29835);
and UO_903 (O_903,N_29905,N_29966);
xor UO_904 (O_904,N_29973,N_29890);
xor UO_905 (O_905,N_29817,N_29804);
nand UO_906 (O_906,N_29958,N_29827);
or UO_907 (O_907,N_29838,N_29841);
nor UO_908 (O_908,N_29921,N_29979);
and UO_909 (O_909,N_29837,N_29901);
and UO_910 (O_910,N_29857,N_29895);
or UO_911 (O_911,N_29918,N_29844);
and UO_912 (O_912,N_29813,N_29893);
and UO_913 (O_913,N_29803,N_29893);
and UO_914 (O_914,N_29849,N_29973);
or UO_915 (O_915,N_29957,N_29953);
xor UO_916 (O_916,N_29807,N_29968);
xor UO_917 (O_917,N_29929,N_29877);
nor UO_918 (O_918,N_29980,N_29856);
or UO_919 (O_919,N_29923,N_29825);
nor UO_920 (O_920,N_29992,N_29836);
xnor UO_921 (O_921,N_29816,N_29808);
or UO_922 (O_922,N_29962,N_29911);
or UO_923 (O_923,N_29816,N_29914);
xor UO_924 (O_924,N_29990,N_29977);
nand UO_925 (O_925,N_29874,N_29904);
nor UO_926 (O_926,N_29991,N_29904);
xor UO_927 (O_927,N_29972,N_29881);
nand UO_928 (O_928,N_29896,N_29932);
and UO_929 (O_929,N_29995,N_29935);
nor UO_930 (O_930,N_29838,N_29945);
or UO_931 (O_931,N_29950,N_29967);
nor UO_932 (O_932,N_29866,N_29959);
xor UO_933 (O_933,N_29881,N_29858);
nor UO_934 (O_934,N_29801,N_29977);
xor UO_935 (O_935,N_29875,N_29965);
or UO_936 (O_936,N_29987,N_29988);
nor UO_937 (O_937,N_29847,N_29936);
xnor UO_938 (O_938,N_29995,N_29933);
xor UO_939 (O_939,N_29862,N_29871);
nand UO_940 (O_940,N_29923,N_29925);
nand UO_941 (O_941,N_29974,N_29944);
nand UO_942 (O_942,N_29955,N_29979);
and UO_943 (O_943,N_29827,N_29953);
and UO_944 (O_944,N_29875,N_29956);
or UO_945 (O_945,N_29804,N_29864);
nor UO_946 (O_946,N_29999,N_29975);
or UO_947 (O_947,N_29830,N_29809);
nor UO_948 (O_948,N_29934,N_29942);
and UO_949 (O_949,N_29958,N_29957);
nand UO_950 (O_950,N_29993,N_29880);
nor UO_951 (O_951,N_29926,N_29995);
nand UO_952 (O_952,N_29809,N_29873);
nand UO_953 (O_953,N_29989,N_29896);
nor UO_954 (O_954,N_29883,N_29895);
nand UO_955 (O_955,N_29894,N_29986);
xor UO_956 (O_956,N_29867,N_29965);
and UO_957 (O_957,N_29861,N_29920);
xnor UO_958 (O_958,N_29824,N_29857);
nor UO_959 (O_959,N_29982,N_29956);
or UO_960 (O_960,N_29856,N_29972);
nor UO_961 (O_961,N_29923,N_29975);
xor UO_962 (O_962,N_29983,N_29951);
or UO_963 (O_963,N_29962,N_29873);
xnor UO_964 (O_964,N_29810,N_29813);
or UO_965 (O_965,N_29988,N_29922);
nor UO_966 (O_966,N_29927,N_29808);
or UO_967 (O_967,N_29854,N_29983);
nor UO_968 (O_968,N_29993,N_29894);
or UO_969 (O_969,N_29828,N_29845);
and UO_970 (O_970,N_29892,N_29813);
xnor UO_971 (O_971,N_29873,N_29990);
nand UO_972 (O_972,N_29860,N_29863);
nand UO_973 (O_973,N_29825,N_29920);
xnor UO_974 (O_974,N_29809,N_29995);
or UO_975 (O_975,N_29855,N_29999);
nand UO_976 (O_976,N_29906,N_29831);
or UO_977 (O_977,N_29847,N_29967);
and UO_978 (O_978,N_29827,N_29918);
nor UO_979 (O_979,N_29875,N_29867);
xor UO_980 (O_980,N_29932,N_29876);
or UO_981 (O_981,N_29811,N_29896);
xnor UO_982 (O_982,N_29962,N_29804);
xnor UO_983 (O_983,N_29997,N_29956);
and UO_984 (O_984,N_29896,N_29925);
nor UO_985 (O_985,N_29835,N_29953);
xnor UO_986 (O_986,N_29999,N_29976);
xor UO_987 (O_987,N_29890,N_29907);
nand UO_988 (O_988,N_29814,N_29928);
xnor UO_989 (O_989,N_29866,N_29805);
and UO_990 (O_990,N_29995,N_29981);
xor UO_991 (O_991,N_29889,N_29866);
nor UO_992 (O_992,N_29932,N_29996);
nand UO_993 (O_993,N_29987,N_29883);
nand UO_994 (O_994,N_29978,N_29972);
or UO_995 (O_995,N_29840,N_29832);
or UO_996 (O_996,N_29923,N_29811);
nor UO_997 (O_997,N_29971,N_29905);
xnor UO_998 (O_998,N_29852,N_29834);
nor UO_999 (O_999,N_29947,N_29839);
nand UO_1000 (O_1000,N_29969,N_29996);
nand UO_1001 (O_1001,N_29891,N_29980);
xor UO_1002 (O_1002,N_29908,N_29880);
and UO_1003 (O_1003,N_29936,N_29826);
nor UO_1004 (O_1004,N_29888,N_29977);
or UO_1005 (O_1005,N_29953,N_29898);
or UO_1006 (O_1006,N_29965,N_29979);
or UO_1007 (O_1007,N_29899,N_29846);
or UO_1008 (O_1008,N_29948,N_29904);
nand UO_1009 (O_1009,N_29841,N_29941);
nor UO_1010 (O_1010,N_29826,N_29812);
nand UO_1011 (O_1011,N_29941,N_29894);
xor UO_1012 (O_1012,N_29957,N_29853);
and UO_1013 (O_1013,N_29808,N_29848);
or UO_1014 (O_1014,N_29821,N_29879);
nand UO_1015 (O_1015,N_29845,N_29904);
and UO_1016 (O_1016,N_29955,N_29849);
or UO_1017 (O_1017,N_29953,N_29976);
nor UO_1018 (O_1018,N_29858,N_29831);
nor UO_1019 (O_1019,N_29996,N_29921);
xor UO_1020 (O_1020,N_29901,N_29912);
nand UO_1021 (O_1021,N_29894,N_29819);
or UO_1022 (O_1022,N_29955,N_29805);
nand UO_1023 (O_1023,N_29943,N_29867);
xnor UO_1024 (O_1024,N_29872,N_29982);
xor UO_1025 (O_1025,N_29910,N_29938);
or UO_1026 (O_1026,N_29837,N_29805);
nand UO_1027 (O_1027,N_29905,N_29965);
and UO_1028 (O_1028,N_29939,N_29849);
or UO_1029 (O_1029,N_29961,N_29901);
xnor UO_1030 (O_1030,N_29850,N_29938);
or UO_1031 (O_1031,N_29855,N_29885);
or UO_1032 (O_1032,N_29996,N_29854);
and UO_1033 (O_1033,N_29832,N_29825);
nand UO_1034 (O_1034,N_29947,N_29930);
and UO_1035 (O_1035,N_29811,N_29912);
or UO_1036 (O_1036,N_29942,N_29997);
and UO_1037 (O_1037,N_29994,N_29980);
or UO_1038 (O_1038,N_29858,N_29842);
and UO_1039 (O_1039,N_29928,N_29902);
nor UO_1040 (O_1040,N_29897,N_29815);
or UO_1041 (O_1041,N_29953,N_29845);
nand UO_1042 (O_1042,N_29925,N_29992);
nand UO_1043 (O_1043,N_29847,N_29905);
and UO_1044 (O_1044,N_29984,N_29859);
xor UO_1045 (O_1045,N_29987,N_29963);
or UO_1046 (O_1046,N_29992,N_29976);
or UO_1047 (O_1047,N_29916,N_29957);
and UO_1048 (O_1048,N_29817,N_29925);
xnor UO_1049 (O_1049,N_29878,N_29943);
xor UO_1050 (O_1050,N_29907,N_29967);
nor UO_1051 (O_1051,N_29915,N_29967);
or UO_1052 (O_1052,N_29853,N_29968);
nor UO_1053 (O_1053,N_29823,N_29951);
or UO_1054 (O_1054,N_29990,N_29812);
or UO_1055 (O_1055,N_29920,N_29893);
xnor UO_1056 (O_1056,N_29812,N_29930);
and UO_1057 (O_1057,N_29967,N_29971);
nor UO_1058 (O_1058,N_29847,N_29945);
and UO_1059 (O_1059,N_29905,N_29906);
nor UO_1060 (O_1060,N_29999,N_29977);
xnor UO_1061 (O_1061,N_29903,N_29893);
and UO_1062 (O_1062,N_29942,N_29861);
xnor UO_1063 (O_1063,N_29840,N_29982);
nor UO_1064 (O_1064,N_29901,N_29898);
nand UO_1065 (O_1065,N_29939,N_29878);
and UO_1066 (O_1066,N_29885,N_29925);
or UO_1067 (O_1067,N_29890,N_29967);
nand UO_1068 (O_1068,N_29822,N_29975);
xor UO_1069 (O_1069,N_29867,N_29940);
nor UO_1070 (O_1070,N_29867,N_29907);
or UO_1071 (O_1071,N_29914,N_29965);
xnor UO_1072 (O_1072,N_29877,N_29998);
nor UO_1073 (O_1073,N_29907,N_29849);
and UO_1074 (O_1074,N_29844,N_29881);
nand UO_1075 (O_1075,N_29848,N_29936);
xor UO_1076 (O_1076,N_29901,N_29892);
nor UO_1077 (O_1077,N_29800,N_29823);
nor UO_1078 (O_1078,N_29906,N_29896);
or UO_1079 (O_1079,N_29937,N_29872);
nor UO_1080 (O_1080,N_29956,N_29917);
xor UO_1081 (O_1081,N_29907,N_29992);
nor UO_1082 (O_1082,N_29995,N_29906);
nor UO_1083 (O_1083,N_29939,N_29959);
or UO_1084 (O_1084,N_29883,N_29819);
and UO_1085 (O_1085,N_29833,N_29886);
nand UO_1086 (O_1086,N_29948,N_29897);
xor UO_1087 (O_1087,N_29921,N_29967);
or UO_1088 (O_1088,N_29843,N_29990);
and UO_1089 (O_1089,N_29977,N_29905);
nand UO_1090 (O_1090,N_29961,N_29934);
xor UO_1091 (O_1091,N_29928,N_29960);
nor UO_1092 (O_1092,N_29954,N_29965);
or UO_1093 (O_1093,N_29941,N_29822);
or UO_1094 (O_1094,N_29977,N_29920);
nor UO_1095 (O_1095,N_29883,N_29851);
nand UO_1096 (O_1096,N_29853,N_29946);
and UO_1097 (O_1097,N_29893,N_29846);
nor UO_1098 (O_1098,N_29950,N_29977);
xor UO_1099 (O_1099,N_29919,N_29916);
xor UO_1100 (O_1100,N_29993,N_29976);
nor UO_1101 (O_1101,N_29820,N_29840);
and UO_1102 (O_1102,N_29880,N_29971);
or UO_1103 (O_1103,N_29895,N_29835);
xnor UO_1104 (O_1104,N_29948,N_29878);
or UO_1105 (O_1105,N_29812,N_29924);
and UO_1106 (O_1106,N_29983,N_29980);
nand UO_1107 (O_1107,N_29967,N_29868);
and UO_1108 (O_1108,N_29969,N_29826);
or UO_1109 (O_1109,N_29856,N_29815);
nor UO_1110 (O_1110,N_29900,N_29922);
or UO_1111 (O_1111,N_29893,N_29914);
nand UO_1112 (O_1112,N_29890,N_29965);
or UO_1113 (O_1113,N_29924,N_29984);
or UO_1114 (O_1114,N_29878,N_29936);
or UO_1115 (O_1115,N_29903,N_29829);
and UO_1116 (O_1116,N_29806,N_29834);
xnor UO_1117 (O_1117,N_29963,N_29845);
xor UO_1118 (O_1118,N_29813,N_29895);
nor UO_1119 (O_1119,N_29835,N_29971);
or UO_1120 (O_1120,N_29947,N_29936);
nor UO_1121 (O_1121,N_29897,N_29922);
or UO_1122 (O_1122,N_29932,N_29922);
or UO_1123 (O_1123,N_29874,N_29825);
xnor UO_1124 (O_1124,N_29830,N_29964);
and UO_1125 (O_1125,N_29846,N_29897);
nand UO_1126 (O_1126,N_29965,N_29987);
or UO_1127 (O_1127,N_29844,N_29961);
or UO_1128 (O_1128,N_29825,N_29938);
and UO_1129 (O_1129,N_29877,N_29923);
xnor UO_1130 (O_1130,N_29834,N_29861);
nand UO_1131 (O_1131,N_29861,N_29990);
xnor UO_1132 (O_1132,N_29864,N_29828);
nor UO_1133 (O_1133,N_29870,N_29908);
or UO_1134 (O_1134,N_29970,N_29811);
or UO_1135 (O_1135,N_29996,N_29851);
nor UO_1136 (O_1136,N_29811,N_29839);
and UO_1137 (O_1137,N_29863,N_29979);
xor UO_1138 (O_1138,N_29827,N_29861);
and UO_1139 (O_1139,N_29906,N_29971);
and UO_1140 (O_1140,N_29837,N_29897);
or UO_1141 (O_1141,N_29898,N_29875);
nor UO_1142 (O_1142,N_29912,N_29868);
nor UO_1143 (O_1143,N_29851,N_29852);
and UO_1144 (O_1144,N_29914,N_29822);
and UO_1145 (O_1145,N_29886,N_29949);
nand UO_1146 (O_1146,N_29810,N_29815);
and UO_1147 (O_1147,N_29999,N_29816);
or UO_1148 (O_1148,N_29869,N_29990);
xnor UO_1149 (O_1149,N_29916,N_29844);
nand UO_1150 (O_1150,N_29967,N_29855);
or UO_1151 (O_1151,N_29977,N_29916);
xnor UO_1152 (O_1152,N_29805,N_29824);
or UO_1153 (O_1153,N_29863,N_29846);
xnor UO_1154 (O_1154,N_29938,N_29927);
and UO_1155 (O_1155,N_29968,N_29908);
nand UO_1156 (O_1156,N_29825,N_29806);
and UO_1157 (O_1157,N_29922,N_29858);
nor UO_1158 (O_1158,N_29882,N_29852);
nand UO_1159 (O_1159,N_29985,N_29969);
or UO_1160 (O_1160,N_29914,N_29943);
xor UO_1161 (O_1161,N_29999,N_29863);
or UO_1162 (O_1162,N_29805,N_29980);
and UO_1163 (O_1163,N_29813,N_29944);
nor UO_1164 (O_1164,N_29811,N_29817);
xnor UO_1165 (O_1165,N_29867,N_29922);
or UO_1166 (O_1166,N_29812,N_29877);
nor UO_1167 (O_1167,N_29993,N_29942);
or UO_1168 (O_1168,N_29833,N_29909);
xor UO_1169 (O_1169,N_29860,N_29966);
or UO_1170 (O_1170,N_29947,N_29896);
xor UO_1171 (O_1171,N_29864,N_29991);
or UO_1172 (O_1172,N_29896,N_29974);
and UO_1173 (O_1173,N_29991,N_29937);
nor UO_1174 (O_1174,N_29825,N_29917);
nand UO_1175 (O_1175,N_29837,N_29826);
nand UO_1176 (O_1176,N_29873,N_29998);
or UO_1177 (O_1177,N_29809,N_29839);
and UO_1178 (O_1178,N_29822,N_29943);
xor UO_1179 (O_1179,N_29931,N_29881);
or UO_1180 (O_1180,N_29934,N_29918);
or UO_1181 (O_1181,N_29901,N_29870);
and UO_1182 (O_1182,N_29822,N_29865);
and UO_1183 (O_1183,N_29970,N_29935);
nor UO_1184 (O_1184,N_29982,N_29997);
xor UO_1185 (O_1185,N_29840,N_29991);
nor UO_1186 (O_1186,N_29909,N_29997);
nor UO_1187 (O_1187,N_29849,N_29883);
and UO_1188 (O_1188,N_29824,N_29820);
nand UO_1189 (O_1189,N_29929,N_29816);
nand UO_1190 (O_1190,N_29947,N_29942);
xor UO_1191 (O_1191,N_29807,N_29867);
nor UO_1192 (O_1192,N_29917,N_29970);
and UO_1193 (O_1193,N_29991,N_29915);
or UO_1194 (O_1194,N_29914,N_29992);
xnor UO_1195 (O_1195,N_29860,N_29915);
xor UO_1196 (O_1196,N_29920,N_29863);
or UO_1197 (O_1197,N_29864,N_29946);
nor UO_1198 (O_1198,N_29885,N_29910);
or UO_1199 (O_1199,N_29961,N_29946);
xor UO_1200 (O_1200,N_29918,N_29814);
nand UO_1201 (O_1201,N_29886,N_29844);
nor UO_1202 (O_1202,N_29830,N_29861);
nor UO_1203 (O_1203,N_29963,N_29955);
or UO_1204 (O_1204,N_29910,N_29801);
nand UO_1205 (O_1205,N_29941,N_29954);
nand UO_1206 (O_1206,N_29881,N_29817);
xnor UO_1207 (O_1207,N_29871,N_29898);
and UO_1208 (O_1208,N_29981,N_29903);
xnor UO_1209 (O_1209,N_29983,N_29872);
or UO_1210 (O_1210,N_29843,N_29837);
or UO_1211 (O_1211,N_29997,N_29973);
nor UO_1212 (O_1212,N_29838,N_29951);
xor UO_1213 (O_1213,N_29989,N_29931);
nand UO_1214 (O_1214,N_29823,N_29938);
and UO_1215 (O_1215,N_29927,N_29989);
xnor UO_1216 (O_1216,N_29938,N_29855);
nor UO_1217 (O_1217,N_29874,N_29958);
nor UO_1218 (O_1218,N_29809,N_29881);
or UO_1219 (O_1219,N_29853,N_29955);
xnor UO_1220 (O_1220,N_29821,N_29969);
nand UO_1221 (O_1221,N_29819,N_29953);
nand UO_1222 (O_1222,N_29811,N_29871);
nor UO_1223 (O_1223,N_29953,N_29972);
xnor UO_1224 (O_1224,N_29890,N_29906);
or UO_1225 (O_1225,N_29908,N_29978);
and UO_1226 (O_1226,N_29870,N_29998);
and UO_1227 (O_1227,N_29834,N_29823);
and UO_1228 (O_1228,N_29885,N_29914);
nor UO_1229 (O_1229,N_29943,N_29831);
nor UO_1230 (O_1230,N_29845,N_29868);
nand UO_1231 (O_1231,N_29848,N_29973);
nand UO_1232 (O_1232,N_29985,N_29814);
nand UO_1233 (O_1233,N_29998,N_29909);
or UO_1234 (O_1234,N_29854,N_29870);
or UO_1235 (O_1235,N_29996,N_29904);
nor UO_1236 (O_1236,N_29882,N_29817);
and UO_1237 (O_1237,N_29870,N_29817);
or UO_1238 (O_1238,N_29951,N_29887);
xor UO_1239 (O_1239,N_29921,N_29896);
nor UO_1240 (O_1240,N_29884,N_29883);
xor UO_1241 (O_1241,N_29993,N_29825);
or UO_1242 (O_1242,N_29913,N_29998);
nand UO_1243 (O_1243,N_29883,N_29809);
nor UO_1244 (O_1244,N_29990,N_29845);
nor UO_1245 (O_1245,N_29947,N_29894);
and UO_1246 (O_1246,N_29887,N_29824);
nand UO_1247 (O_1247,N_29959,N_29913);
xor UO_1248 (O_1248,N_29885,N_29999);
nand UO_1249 (O_1249,N_29913,N_29900);
or UO_1250 (O_1250,N_29876,N_29808);
nand UO_1251 (O_1251,N_29985,N_29931);
nand UO_1252 (O_1252,N_29877,N_29837);
nand UO_1253 (O_1253,N_29815,N_29900);
nor UO_1254 (O_1254,N_29835,N_29856);
nand UO_1255 (O_1255,N_29904,N_29813);
or UO_1256 (O_1256,N_29912,N_29853);
xor UO_1257 (O_1257,N_29888,N_29993);
or UO_1258 (O_1258,N_29958,N_29822);
and UO_1259 (O_1259,N_29977,N_29883);
nor UO_1260 (O_1260,N_29854,N_29895);
nand UO_1261 (O_1261,N_29913,N_29901);
nand UO_1262 (O_1262,N_29979,N_29992);
and UO_1263 (O_1263,N_29954,N_29906);
nand UO_1264 (O_1264,N_29949,N_29859);
nand UO_1265 (O_1265,N_29852,N_29890);
or UO_1266 (O_1266,N_29811,N_29927);
nand UO_1267 (O_1267,N_29917,N_29913);
nand UO_1268 (O_1268,N_29828,N_29956);
nand UO_1269 (O_1269,N_29859,N_29825);
nand UO_1270 (O_1270,N_29926,N_29952);
nor UO_1271 (O_1271,N_29982,N_29833);
nand UO_1272 (O_1272,N_29805,N_29945);
and UO_1273 (O_1273,N_29821,N_29859);
nor UO_1274 (O_1274,N_29859,N_29965);
and UO_1275 (O_1275,N_29920,N_29820);
nand UO_1276 (O_1276,N_29877,N_29903);
nand UO_1277 (O_1277,N_29901,N_29900);
xor UO_1278 (O_1278,N_29987,N_29835);
nand UO_1279 (O_1279,N_29913,N_29885);
or UO_1280 (O_1280,N_29857,N_29863);
nand UO_1281 (O_1281,N_29924,N_29955);
or UO_1282 (O_1282,N_29964,N_29897);
and UO_1283 (O_1283,N_29869,N_29820);
or UO_1284 (O_1284,N_29829,N_29869);
or UO_1285 (O_1285,N_29997,N_29938);
or UO_1286 (O_1286,N_29886,N_29897);
xnor UO_1287 (O_1287,N_29949,N_29918);
and UO_1288 (O_1288,N_29915,N_29924);
or UO_1289 (O_1289,N_29886,N_29883);
nand UO_1290 (O_1290,N_29916,N_29835);
nor UO_1291 (O_1291,N_29857,N_29991);
xnor UO_1292 (O_1292,N_29999,N_29940);
or UO_1293 (O_1293,N_29853,N_29825);
and UO_1294 (O_1294,N_29918,N_29901);
or UO_1295 (O_1295,N_29854,N_29891);
nand UO_1296 (O_1296,N_29935,N_29864);
nand UO_1297 (O_1297,N_29991,N_29865);
xor UO_1298 (O_1298,N_29952,N_29898);
xnor UO_1299 (O_1299,N_29993,N_29919);
xor UO_1300 (O_1300,N_29855,N_29974);
and UO_1301 (O_1301,N_29904,N_29906);
nand UO_1302 (O_1302,N_29986,N_29811);
or UO_1303 (O_1303,N_29809,N_29934);
or UO_1304 (O_1304,N_29937,N_29845);
or UO_1305 (O_1305,N_29842,N_29994);
xnor UO_1306 (O_1306,N_29883,N_29930);
and UO_1307 (O_1307,N_29888,N_29866);
xnor UO_1308 (O_1308,N_29900,N_29853);
xnor UO_1309 (O_1309,N_29928,N_29892);
and UO_1310 (O_1310,N_29839,N_29843);
or UO_1311 (O_1311,N_29850,N_29987);
nand UO_1312 (O_1312,N_29948,N_29909);
nor UO_1313 (O_1313,N_29954,N_29886);
xor UO_1314 (O_1314,N_29887,N_29862);
xnor UO_1315 (O_1315,N_29869,N_29981);
xor UO_1316 (O_1316,N_29822,N_29814);
or UO_1317 (O_1317,N_29823,N_29950);
or UO_1318 (O_1318,N_29926,N_29817);
and UO_1319 (O_1319,N_29997,N_29899);
nor UO_1320 (O_1320,N_29957,N_29989);
nor UO_1321 (O_1321,N_29907,N_29879);
and UO_1322 (O_1322,N_29826,N_29909);
or UO_1323 (O_1323,N_29802,N_29956);
xnor UO_1324 (O_1324,N_29828,N_29957);
nor UO_1325 (O_1325,N_29985,N_29897);
or UO_1326 (O_1326,N_29886,N_29863);
nand UO_1327 (O_1327,N_29804,N_29984);
or UO_1328 (O_1328,N_29813,N_29862);
or UO_1329 (O_1329,N_29836,N_29808);
or UO_1330 (O_1330,N_29947,N_29921);
xor UO_1331 (O_1331,N_29919,N_29955);
xnor UO_1332 (O_1332,N_29901,N_29829);
nor UO_1333 (O_1333,N_29842,N_29935);
and UO_1334 (O_1334,N_29836,N_29899);
or UO_1335 (O_1335,N_29916,N_29822);
nor UO_1336 (O_1336,N_29900,N_29925);
and UO_1337 (O_1337,N_29821,N_29878);
and UO_1338 (O_1338,N_29904,N_29825);
or UO_1339 (O_1339,N_29899,N_29874);
nor UO_1340 (O_1340,N_29824,N_29827);
xnor UO_1341 (O_1341,N_29822,N_29875);
and UO_1342 (O_1342,N_29979,N_29944);
nor UO_1343 (O_1343,N_29976,N_29838);
nand UO_1344 (O_1344,N_29980,N_29858);
and UO_1345 (O_1345,N_29946,N_29866);
xnor UO_1346 (O_1346,N_29875,N_29804);
and UO_1347 (O_1347,N_29933,N_29991);
and UO_1348 (O_1348,N_29855,N_29930);
nor UO_1349 (O_1349,N_29895,N_29978);
or UO_1350 (O_1350,N_29980,N_29952);
nand UO_1351 (O_1351,N_29820,N_29933);
nor UO_1352 (O_1352,N_29836,N_29944);
nor UO_1353 (O_1353,N_29925,N_29895);
and UO_1354 (O_1354,N_29829,N_29863);
and UO_1355 (O_1355,N_29940,N_29944);
or UO_1356 (O_1356,N_29853,N_29892);
and UO_1357 (O_1357,N_29966,N_29821);
or UO_1358 (O_1358,N_29840,N_29826);
nand UO_1359 (O_1359,N_29930,N_29862);
xnor UO_1360 (O_1360,N_29923,N_29840);
xnor UO_1361 (O_1361,N_29886,N_29998);
nor UO_1362 (O_1362,N_29852,N_29932);
nor UO_1363 (O_1363,N_29900,N_29890);
xor UO_1364 (O_1364,N_29832,N_29969);
or UO_1365 (O_1365,N_29805,N_29971);
or UO_1366 (O_1366,N_29850,N_29839);
and UO_1367 (O_1367,N_29859,N_29900);
xnor UO_1368 (O_1368,N_29976,N_29856);
nor UO_1369 (O_1369,N_29859,N_29927);
xor UO_1370 (O_1370,N_29832,N_29866);
nand UO_1371 (O_1371,N_29928,N_29875);
and UO_1372 (O_1372,N_29957,N_29852);
nor UO_1373 (O_1373,N_29921,N_29952);
nand UO_1374 (O_1374,N_29841,N_29866);
and UO_1375 (O_1375,N_29942,N_29949);
xor UO_1376 (O_1376,N_29817,N_29966);
nor UO_1377 (O_1377,N_29867,N_29897);
and UO_1378 (O_1378,N_29935,N_29899);
nor UO_1379 (O_1379,N_29917,N_29827);
xnor UO_1380 (O_1380,N_29815,N_29887);
and UO_1381 (O_1381,N_29962,N_29965);
nor UO_1382 (O_1382,N_29911,N_29976);
nand UO_1383 (O_1383,N_29821,N_29924);
and UO_1384 (O_1384,N_29849,N_29984);
xor UO_1385 (O_1385,N_29938,N_29941);
nand UO_1386 (O_1386,N_29959,N_29992);
xor UO_1387 (O_1387,N_29819,N_29979);
xnor UO_1388 (O_1388,N_29810,N_29896);
nor UO_1389 (O_1389,N_29944,N_29997);
and UO_1390 (O_1390,N_29869,N_29946);
xnor UO_1391 (O_1391,N_29917,N_29979);
nor UO_1392 (O_1392,N_29828,N_29871);
or UO_1393 (O_1393,N_29866,N_29914);
nand UO_1394 (O_1394,N_29994,N_29910);
and UO_1395 (O_1395,N_29800,N_29895);
or UO_1396 (O_1396,N_29905,N_29918);
or UO_1397 (O_1397,N_29803,N_29916);
and UO_1398 (O_1398,N_29885,N_29827);
nand UO_1399 (O_1399,N_29972,N_29917);
and UO_1400 (O_1400,N_29942,N_29935);
nor UO_1401 (O_1401,N_29852,N_29840);
or UO_1402 (O_1402,N_29944,N_29925);
nor UO_1403 (O_1403,N_29936,N_29920);
and UO_1404 (O_1404,N_29989,N_29992);
xor UO_1405 (O_1405,N_29997,N_29837);
or UO_1406 (O_1406,N_29841,N_29806);
nor UO_1407 (O_1407,N_29854,N_29836);
nand UO_1408 (O_1408,N_29923,N_29861);
xor UO_1409 (O_1409,N_29873,N_29832);
xnor UO_1410 (O_1410,N_29874,N_29888);
nand UO_1411 (O_1411,N_29964,N_29850);
xnor UO_1412 (O_1412,N_29852,N_29847);
nand UO_1413 (O_1413,N_29869,N_29908);
or UO_1414 (O_1414,N_29898,N_29990);
nand UO_1415 (O_1415,N_29906,N_29822);
xnor UO_1416 (O_1416,N_29869,N_29826);
and UO_1417 (O_1417,N_29824,N_29920);
or UO_1418 (O_1418,N_29905,N_29840);
and UO_1419 (O_1419,N_29957,N_29927);
or UO_1420 (O_1420,N_29915,N_29982);
and UO_1421 (O_1421,N_29904,N_29882);
and UO_1422 (O_1422,N_29955,N_29886);
nor UO_1423 (O_1423,N_29925,N_29912);
or UO_1424 (O_1424,N_29980,N_29988);
xor UO_1425 (O_1425,N_29842,N_29835);
or UO_1426 (O_1426,N_29824,N_29917);
and UO_1427 (O_1427,N_29990,N_29849);
nor UO_1428 (O_1428,N_29867,N_29838);
or UO_1429 (O_1429,N_29934,N_29808);
xor UO_1430 (O_1430,N_29904,N_29926);
nor UO_1431 (O_1431,N_29966,N_29996);
nor UO_1432 (O_1432,N_29958,N_29817);
xnor UO_1433 (O_1433,N_29908,N_29922);
or UO_1434 (O_1434,N_29940,N_29929);
and UO_1435 (O_1435,N_29812,N_29916);
and UO_1436 (O_1436,N_29833,N_29882);
and UO_1437 (O_1437,N_29829,N_29846);
or UO_1438 (O_1438,N_29970,N_29987);
nor UO_1439 (O_1439,N_29831,N_29904);
nand UO_1440 (O_1440,N_29836,N_29993);
and UO_1441 (O_1441,N_29973,N_29858);
or UO_1442 (O_1442,N_29873,N_29907);
and UO_1443 (O_1443,N_29982,N_29891);
xor UO_1444 (O_1444,N_29880,N_29980);
and UO_1445 (O_1445,N_29935,N_29816);
or UO_1446 (O_1446,N_29947,N_29803);
nor UO_1447 (O_1447,N_29913,N_29966);
nand UO_1448 (O_1448,N_29859,N_29987);
nand UO_1449 (O_1449,N_29881,N_29885);
or UO_1450 (O_1450,N_29933,N_29908);
xor UO_1451 (O_1451,N_29928,N_29990);
and UO_1452 (O_1452,N_29942,N_29813);
or UO_1453 (O_1453,N_29967,N_29807);
or UO_1454 (O_1454,N_29906,N_29961);
or UO_1455 (O_1455,N_29992,N_29856);
nor UO_1456 (O_1456,N_29985,N_29947);
xor UO_1457 (O_1457,N_29934,N_29939);
nand UO_1458 (O_1458,N_29880,N_29816);
and UO_1459 (O_1459,N_29835,N_29927);
xnor UO_1460 (O_1460,N_29832,N_29819);
nor UO_1461 (O_1461,N_29845,N_29926);
nand UO_1462 (O_1462,N_29942,N_29969);
or UO_1463 (O_1463,N_29907,N_29928);
nand UO_1464 (O_1464,N_29811,N_29945);
nor UO_1465 (O_1465,N_29981,N_29852);
nand UO_1466 (O_1466,N_29897,N_29842);
nor UO_1467 (O_1467,N_29819,N_29908);
or UO_1468 (O_1468,N_29833,N_29850);
or UO_1469 (O_1469,N_29868,N_29897);
or UO_1470 (O_1470,N_29924,N_29825);
nand UO_1471 (O_1471,N_29964,N_29884);
or UO_1472 (O_1472,N_29959,N_29969);
and UO_1473 (O_1473,N_29940,N_29813);
or UO_1474 (O_1474,N_29983,N_29893);
and UO_1475 (O_1475,N_29932,N_29823);
nand UO_1476 (O_1476,N_29940,N_29917);
and UO_1477 (O_1477,N_29896,N_29948);
nor UO_1478 (O_1478,N_29991,N_29955);
xnor UO_1479 (O_1479,N_29913,N_29970);
nor UO_1480 (O_1480,N_29916,N_29840);
xnor UO_1481 (O_1481,N_29804,N_29918);
and UO_1482 (O_1482,N_29852,N_29898);
xor UO_1483 (O_1483,N_29908,N_29887);
and UO_1484 (O_1484,N_29855,N_29903);
xor UO_1485 (O_1485,N_29938,N_29828);
and UO_1486 (O_1486,N_29905,N_29850);
xnor UO_1487 (O_1487,N_29871,N_29891);
and UO_1488 (O_1488,N_29881,N_29998);
xnor UO_1489 (O_1489,N_29925,N_29924);
and UO_1490 (O_1490,N_29934,N_29964);
xor UO_1491 (O_1491,N_29841,N_29972);
and UO_1492 (O_1492,N_29903,N_29882);
and UO_1493 (O_1493,N_29834,N_29924);
xnor UO_1494 (O_1494,N_29916,N_29987);
or UO_1495 (O_1495,N_29862,N_29855);
nand UO_1496 (O_1496,N_29823,N_29892);
or UO_1497 (O_1497,N_29940,N_29961);
and UO_1498 (O_1498,N_29902,N_29894);
xnor UO_1499 (O_1499,N_29846,N_29963);
and UO_1500 (O_1500,N_29927,N_29914);
nor UO_1501 (O_1501,N_29909,N_29922);
nor UO_1502 (O_1502,N_29920,N_29894);
nand UO_1503 (O_1503,N_29848,N_29957);
and UO_1504 (O_1504,N_29810,N_29879);
or UO_1505 (O_1505,N_29918,N_29969);
nand UO_1506 (O_1506,N_29931,N_29876);
nand UO_1507 (O_1507,N_29822,N_29883);
nand UO_1508 (O_1508,N_29975,N_29869);
and UO_1509 (O_1509,N_29809,N_29924);
nor UO_1510 (O_1510,N_29814,N_29878);
or UO_1511 (O_1511,N_29847,N_29896);
and UO_1512 (O_1512,N_29919,N_29880);
nand UO_1513 (O_1513,N_29842,N_29864);
or UO_1514 (O_1514,N_29873,N_29833);
xnor UO_1515 (O_1515,N_29812,N_29921);
nor UO_1516 (O_1516,N_29970,N_29892);
nand UO_1517 (O_1517,N_29910,N_29830);
nor UO_1518 (O_1518,N_29867,N_29850);
xor UO_1519 (O_1519,N_29885,N_29940);
nand UO_1520 (O_1520,N_29945,N_29984);
and UO_1521 (O_1521,N_29847,N_29863);
and UO_1522 (O_1522,N_29893,N_29951);
nand UO_1523 (O_1523,N_29831,N_29972);
xnor UO_1524 (O_1524,N_29821,N_29938);
nor UO_1525 (O_1525,N_29919,N_29810);
nand UO_1526 (O_1526,N_29846,N_29988);
xnor UO_1527 (O_1527,N_29833,N_29972);
and UO_1528 (O_1528,N_29854,N_29873);
or UO_1529 (O_1529,N_29843,N_29884);
and UO_1530 (O_1530,N_29855,N_29803);
nand UO_1531 (O_1531,N_29846,N_29936);
or UO_1532 (O_1532,N_29982,N_29870);
or UO_1533 (O_1533,N_29931,N_29898);
nand UO_1534 (O_1534,N_29930,N_29861);
and UO_1535 (O_1535,N_29851,N_29947);
xor UO_1536 (O_1536,N_29921,N_29821);
and UO_1537 (O_1537,N_29973,N_29810);
or UO_1538 (O_1538,N_29804,N_29852);
xor UO_1539 (O_1539,N_29990,N_29920);
or UO_1540 (O_1540,N_29817,N_29957);
nand UO_1541 (O_1541,N_29986,N_29857);
nor UO_1542 (O_1542,N_29999,N_29838);
nor UO_1543 (O_1543,N_29828,N_29998);
nor UO_1544 (O_1544,N_29895,N_29850);
and UO_1545 (O_1545,N_29851,N_29842);
or UO_1546 (O_1546,N_29845,N_29911);
and UO_1547 (O_1547,N_29971,N_29999);
xor UO_1548 (O_1548,N_29939,N_29897);
or UO_1549 (O_1549,N_29945,N_29891);
nor UO_1550 (O_1550,N_29830,N_29877);
xor UO_1551 (O_1551,N_29848,N_29861);
xor UO_1552 (O_1552,N_29995,N_29968);
nand UO_1553 (O_1553,N_29964,N_29808);
and UO_1554 (O_1554,N_29993,N_29944);
or UO_1555 (O_1555,N_29819,N_29924);
and UO_1556 (O_1556,N_29923,N_29907);
nor UO_1557 (O_1557,N_29816,N_29884);
nand UO_1558 (O_1558,N_29985,N_29809);
xnor UO_1559 (O_1559,N_29883,N_29811);
or UO_1560 (O_1560,N_29986,N_29949);
nand UO_1561 (O_1561,N_29821,N_29955);
and UO_1562 (O_1562,N_29899,N_29983);
and UO_1563 (O_1563,N_29945,N_29968);
xnor UO_1564 (O_1564,N_29859,N_29928);
nand UO_1565 (O_1565,N_29916,N_29911);
nand UO_1566 (O_1566,N_29916,N_29864);
or UO_1567 (O_1567,N_29868,N_29854);
nor UO_1568 (O_1568,N_29963,N_29854);
or UO_1569 (O_1569,N_29838,N_29967);
nand UO_1570 (O_1570,N_29847,N_29930);
or UO_1571 (O_1571,N_29875,N_29937);
xor UO_1572 (O_1572,N_29935,N_29822);
nand UO_1573 (O_1573,N_29851,N_29933);
and UO_1574 (O_1574,N_29971,N_29844);
and UO_1575 (O_1575,N_29831,N_29879);
nor UO_1576 (O_1576,N_29839,N_29870);
nor UO_1577 (O_1577,N_29925,N_29904);
and UO_1578 (O_1578,N_29865,N_29844);
xnor UO_1579 (O_1579,N_29998,N_29921);
and UO_1580 (O_1580,N_29986,N_29927);
nand UO_1581 (O_1581,N_29976,N_29981);
nor UO_1582 (O_1582,N_29925,N_29831);
xor UO_1583 (O_1583,N_29953,N_29946);
nor UO_1584 (O_1584,N_29815,N_29968);
xor UO_1585 (O_1585,N_29876,N_29949);
nand UO_1586 (O_1586,N_29944,N_29954);
nor UO_1587 (O_1587,N_29902,N_29861);
nand UO_1588 (O_1588,N_29902,N_29927);
or UO_1589 (O_1589,N_29845,N_29863);
nor UO_1590 (O_1590,N_29887,N_29971);
or UO_1591 (O_1591,N_29914,N_29937);
nand UO_1592 (O_1592,N_29981,N_29956);
nand UO_1593 (O_1593,N_29983,N_29814);
nand UO_1594 (O_1594,N_29912,N_29816);
xor UO_1595 (O_1595,N_29853,N_29879);
or UO_1596 (O_1596,N_29833,N_29918);
and UO_1597 (O_1597,N_29835,N_29865);
xnor UO_1598 (O_1598,N_29914,N_29884);
and UO_1599 (O_1599,N_29902,N_29830);
nand UO_1600 (O_1600,N_29953,N_29956);
nor UO_1601 (O_1601,N_29841,N_29875);
xor UO_1602 (O_1602,N_29815,N_29883);
xor UO_1603 (O_1603,N_29902,N_29842);
and UO_1604 (O_1604,N_29836,N_29811);
or UO_1605 (O_1605,N_29846,N_29985);
or UO_1606 (O_1606,N_29923,N_29981);
or UO_1607 (O_1607,N_29850,N_29989);
nor UO_1608 (O_1608,N_29820,N_29826);
or UO_1609 (O_1609,N_29806,N_29989);
nor UO_1610 (O_1610,N_29970,N_29861);
xor UO_1611 (O_1611,N_29972,N_29998);
xnor UO_1612 (O_1612,N_29879,N_29889);
and UO_1613 (O_1613,N_29900,N_29920);
nor UO_1614 (O_1614,N_29865,N_29930);
or UO_1615 (O_1615,N_29830,N_29997);
xnor UO_1616 (O_1616,N_29844,N_29895);
or UO_1617 (O_1617,N_29990,N_29907);
and UO_1618 (O_1618,N_29880,N_29943);
and UO_1619 (O_1619,N_29906,N_29951);
or UO_1620 (O_1620,N_29817,N_29978);
or UO_1621 (O_1621,N_29947,N_29991);
nand UO_1622 (O_1622,N_29875,N_29990);
nor UO_1623 (O_1623,N_29832,N_29807);
xor UO_1624 (O_1624,N_29888,N_29822);
or UO_1625 (O_1625,N_29862,N_29809);
xnor UO_1626 (O_1626,N_29841,N_29989);
xnor UO_1627 (O_1627,N_29912,N_29913);
nand UO_1628 (O_1628,N_29905,N_29999);
nand UO_1629 (O_1629,N_29978,N_29942);
and UO_1630 (O_1630,N_29848,N_29999);
and UO_1631 (O_1631,N_29928,N_29810);
nand UO_1632 (O_1632,N_29863,N_29887);
and UO_1633 (O_1633,N_29968,N_29889);
or UO_1634 (O_1634,N_29940,N_29806);
and UO_1635 (O_1635,N_29971,N_29979);
nor UO_1636 (O_1636,N_29968,N_29981);
or UO_1637 (O_1637,N_29930,N_29878);
and UO_1638 (O_1638,N_29817,N_29904);
xnor UO_1639 (O_1639,N_29827,N_29807);
and UO_1640 (O_1640,N_29809,N_29825);
or UO_1641 (O_1641,N_29909,N_29940);
xnor UO_1642 (O_1642,N_29861,N_29973);
nor UO_1643 (O_1643,N_29990,N_29836);
or UO_1644 (O_1644,N_29998,N_29926);
nand UO_1645 (O_1645,N_29893,N_29863);
nor UO_1646 (O_1646,N_29827,N_29902);
nand UO_1647 (O_1647,N_29911,N_29812);
nor UO_1648 (O_1648,N_29983,N_29946);
nor UO_1649 (O_1649,N_29983,N_29944);
and UO_1650 (O_1650,N_29920,N_29917);
xor UO_1651 (O_1651,N_29831,N_29851);
and UO_1652 (O_1652,N_29831,N_29886);
nand UO_1653 (O_1653,N_29961,N_29888);
xnor UO_1654 (O_1654,N_29893,N_29871);
and UO_1655 (O_1655,N_29970,N_29964);
or UO_1656 (O_1656,N_29878,N_29918);
nor UO_1657 (O_1657,N_29974,N_29946);
nor UO_1658 (O_1658,N_29903,N_29819);
or UO_1659 (O_1659,N_29853,N_29990);
nor UO_1660 (O_1660,N_29991,N_29897);
nor UO_1661 (O_1661,N_29963,N_29954);
and UO_1662 (O_1662,N_29955,N_29878);
nand UO_1663 (O_1663,N_29910,N_29986);
and UO_1664 (O_1664,N_29867,N_29937);
or UO_1665 (O_1665,N_29981,N_29957);
nand UO_1666 (O_1666,N_29855,N_29942);
or UO_1667 (O_1667,N_29887,N_29847);
nor UO_1668 (O_1668,N_29862,N_29905);
and UO_1669 (O_1669,N_29914,N_29930);
or UO_1670 (O_1670,N_29917,N_29916);
nand UO_1671 (O_1671,N_29934,N_29940);
and UO_1672 (O_1672,N_29829,N_29986);
and UO_1673 (O_1673,N_29966,N_29951);
and UO_1674 (O_1674,N_29800,N_29960);
xnor UO_1675 (O_1675,N_29834,N_29894);
or UO_1676 (O_1676,N_29980,N_29804);
and UO_1677 (O_1677,N_29982,N_29843);
and UO_1678 (O_1678,N_29962,N_29940);
nand UO_1679 (O_1679,N_29990,N_29992);
nor UO_1680 (O_1680,N_29931,N_29899);
nor UO_1681 (O_1681,N_29858,N_29851);
nand UO_1682 (O_1682,N_29872,N_29831);
xnor UO_1683 (O_1683,N_29857,N_29815);
nor UO_1684 (O_1684,N_29804,N_29806);
and UO_1685 (O_1685,N_29926,N_29814);
xnor UO_1686 (O_1686,N_29846,N_29970);
nor UO_1687 (O_1687,N_29883,N_29872);
nand UO_1688 (O_1688,N_29807,N_29800);
or UO_1689 (O_1689,N_29854,N_29906);
nor UO_1690 (O_1690,N_29922,N_29817);
nor UO_1691 (O_1691,N_29954,N_29840);
or UO_1692 (O_1692,N_29850,N_29976);
or UO_1693 (O_1693,N_29875,N_29982);
or UO_1694 (O_1694,N_29909,N_29875);
or UO_1695 (O_1695,N_29800,N_29888);
xnor UO_1696 (O_1696,N_29968,N_29909);
xnor UO_1697 (O_1697,N_29952,N_29884);
nor UO_1698 (O_1698,N_29848,N_29974);
xor UO_1699 (O_1699,N_29871,N_29982);
nand UO_1700 (O_1700,N_29929,N_29840);
nand UO_1701 (O_1701,N_29925,N_29830);
nor UO_1702 (O_1702,N_29936,N_29873);
xnor UO_1703 (O_1703,N_29937,N_29907);
and UO_1704 (O_1704,N_29970,N_29832);
xnor UO_1705 (O_1705,N_29807,N_29955);
or UO_1706 (O_1706,N_29831,N_29819);
and UO_1707 (O_1707,N_29965,N_29974);
nor UO_1708 (O_1708,N_29913,N_29871);
xor UO_1709 (O_1709,N_29981,N_29843);
or UO_1710 (O_1710,N_29837,N_29894);
nand UO_1711 (O_1711,N_29935,N_29947);
nor UO_1712 (O_1712,N_29992,N_29900);
nor UO_1713 (O_1713,N_29838,N_29909);
xnor UO_1714 (O_1714,N_29968,N_29846);
or UO_1715 (O_1715,N_29863,N_29911);
and UO_1716 (O_1716,N_29920,N_29821);
nor UO_1717 (O_1717,N_29841,N_29839);
nor UO_1718 (O_1718,N_29963,N_29806);
nand UO_1719 (O_1719,N_29883,N_29952);
xor UO_1720 (O_1720,N_29959,N_29914);
nand UO_1721 (O_1721,N_29806,N_29863);
or UO_1722 (O_1722,N_29812,N_29890);
xnor UO_1723 (O_1723,N_29842,N_29874);
nand UO_1724 (O_1724,N_29825,N_29847);
or UO_1725 (O_1725,N_29954,N_29936);
or UO_1726 (O_1726,N_29827,N_29852);
and UO_1727 (O_1727,N_29955,N_29874);
nor UO_1728 (O_1728,N_29898,N_29883);
nand UO_1729 (O_1729,N_29936,N_29956);
and UO_1730 (O_1730,N_29893,N_29953);
or UO_1731 (O_1731,N_29972,N_29911);
nor UO_1732 (O_1732,N_29964,N_29946);
nor UO_1733 (O_1733,N_29939,N_29977);
xnor UO_1734 (O_1734,N_29898,N_29872);
or UO_1735 (O_1735,N_29935,N_29979);
xnor UO_1736 (O_1736,N_29971,N_29864);
xnor UO_1737 (O_1737,N_29917,N_29878);
nor UO_1738 (O_1738,N_29868,N_29818);
nand UO_1739 (O_1739,N_29841,N_29895);
and UO_1740 (O_1740,N_29978,N_29835);
nand UO_1741 (O_1741,N_29896,N_29910);
xnor UO_1742 (O_1742,N_29934,N_29938);
and UO_1743 (O_1743,N_29894,N_29871);
or UO_1744 (O_1744,N_29908,N_29838);
and UO_1745 (O_1745,N_29929,N_29924);
or UO_1746 (O_1746,N_29860,N_29988);
xor UO_1747 (O_1747,N_29855,N_29911);
and UO_1748 (O_1748,N_29989,N_29953);
nand UO_1749 (O_1749,N_29924,N_29874);
nor UO_1750 (O_1750,N_29916,N_29847);
or UO_1751 (O_1751,N_29954,N_29983);
nand UO_1752 (O_1752,N_29817,N_29906);
and UO_1753 (O_1753,N_29877,N_29988);
or UO_1754 (O_1754,N_29946,N_29919);
nand UO_1755 (O_1755,N_29932,N_29919);
or UO_1756 (O_1756,N_29928,N_29824);
or UO_1757 (O_1757,N_29854,N_29964);
nor UO_1758 (O_1758,N_29870,N_29981);
or UO_1759 (O_1759,N_29930,N_29849);
and UO_1760 (O_1760,N_29994,N_29921);
xor UO_1761 (O_1761,N_29834,N_29885);
or UO_1762 (O_1762,N_29835,N_29854);
xor UO_1763 (O_1763,N_29898,N_29947);
and UO_1764 (O_1764,N_29903,N_29834);
or UO_1765 (O_1765,N_29857,N_29963);
or UO_1766 (O_1766,N_29908,N_29999);
xor UO_1767 (O_1767,N_29830,N_29992);
xnor UO_1768 (O_1768,N_29807,N_29842);
or UO_1769 (O_1769,N_29839,N_29962);
or UO_1770 (O_1770,N_29940,N_29910);
xor UO_1771 (O_1771,N_29945,N_29985);
xor UO_1772 (O_1772,N_29838,N_29860);
nor UO_1773 (O_1773,N_29939,N_29935);
nor UO_1774 (O_1774,N_29904,N_29818);
nand UO_1775 (O_1775,N_29987,N_29855);
and UO_1776 (O_1776,N_29928,N_29956);
or UO_1777 (O_1777,N_29905,N_29898);
nand UO_1778 (O_1778,N_29812,N_29875);
nor UO_1779 (O_1779,N_29859,N_29898);
or UO_1780 (O_1780,N_29891,N_29939);
or UO_1781 (O_1781,N_29831,N_29896);
or UO_1782 (O_1782,N_29902,N_29891);
xnor UO_1783 (O_1783,N_29808,N_29954);
xor UO_1784 (O_1784,N_29813,N_29850);
xor UO_1785 (O_1785,N_29875,N_29897);
and UO_1786 (O_1786,N_29913,N_29973);
nand UO_1787 (O_1787,N_29941,N_29985);
and UO_1788 (O_1788,N_29959,N_29835);
xor UO_1789 (O_1789,N_29983,N_29819);
and UO_1790 (O_1790,N_29950,N_29988);
and UO_1791 (O_1791,N_29808,N_29944);
nand UO_1792 (O_1792,N_29975,N_29857);
nand UO_1793 (O_1793,N_29849,N_29838);
and UO_1794 (O_1794,N_29991,N_29851);
nand UO_1795 (O_1795,N_29834,N_29807);
nand UO_1796 (O_1796,N_29869,N_29889);
or UO_1797 (O_1797,N_29895,N_29979);
nand UO_1798 (O_1798,N_29956,N_29901);
nand UO_1799 (O_1799,N_29984,N_29970);
or UO_1800 (O_1800,N_29853,N_29803);
xnor UO_1801 (O_1801,N_29987,N_29893);
and UO_1802 (O_1802,N_29992,N_29881);
and UO_1803 (O_1803,N_29943,N_29938);
nor UO_1804 (O_1804,N_29991,N_29815);
xor UO_1805 (O_1805,N_29824,N_29877);
nor UO_1806 (O_1806,N_29875,N_29808);
nor UO_1807 (O_1807,N_29815,N_29987);
nand UO_1808 (O_1808,N_29885,N_29982);
nor UO_1809 (O_1809,N_29822,N_29884);
nor UO_1810 (O_1810,N_29962,N_29916);
and UO_1811 (O_1811,N_29909,N_29902);
nand UO_1812 (O_1812,N_29811,N_29851);
or UO_1813 (O_1813,N_29841,N_29918);
nor UO_1814 (O_1814,N_29896,N_29955);
or UO_1815 (O_1815,N_29891,N_29819);
xnor UO_1816 (O_1816,N_29910,N_29915);
nand UO_1817 (O_1817,N_29814,N_29916);
or UO_1818 (O_1818,N_29830,N_29967);
and UO_1819 (O_1819,N_29844,N_29945);
or UO_1820 (O_1820,N_29832,N_29801);
and UO_1821 (O_1821,N_29946,N_29985);
nand UO_1822 (O_1822,N_29978,N_29837);
nor UO_1823 (O_1823,N_29845,N_29942);
and UO_1824 (O_1824,N_29824,N_29921);
and UO_1825 (O_1825,N_29862,N_29831);
and UO_1826 (O_1826,N_29804,N_29857);
nor UO_1827 (O_1827,N_29898,N_29836);
nor UO_1828 (O_1828,N_29895,N_29910);
and UO_1829 (O_1829,N_29909,N_29923);
and UO_1830 (O_1830,N_29913,N_29877);
nand UO_1831 (O_1831,N_29834,N_29848);
nor UO_1832 (O_1832,N_29861,N_29935);
and UO_1833 (O_1833,N_29967,N_29885);
and UO_1834 (O_1834,N_29906,N_29946);
xor UO_1835 (O_1835,N_29872,N_29879);
nand UO_1836 (O_1836,N_29834,N_29976);
nand UO_1837 (O_1837,N_29873,N_29939);
and UO_1838 (O_1838,N_29921,N_29955);
xnor UO_1839 (O_1839,N_29894,N_29999);
nand UO_1840 (O_1840,N_29859,N_29936);
nor UO_1841 (O_1841,N_29927,N_29840);
nand UO_1842 (O_1842,N_29993,N_29887);
and UO_1843 (O_1843,N_29876,N_29836);
xnor UO_1844 (O_1844,N_29977,N_29859);
nor UO_1845 (O_1845,N_29932,N_29808);
nor UO_1846 (O_1846,N_29839,N_29836);
and UO_1847 (O_1847,N_29986,N_29808);
nand UO_1848 (O_1848,N_29922,N_29971);
nand UO_1849 (O_1849,N_29908,N_29861);
and UO_1850 (O_1850,N_29916,N_29951);
xor UO_1851 (O_1851,N_29866,N_29834);
nor UO_1852 (O_1852,N_29849,N_29879);
nor UO_1853 (O_1853,N_29887,N_29832);
xor UO_1854 (O_1854,N_29837,N_29900);
nand UO_1855 (O_1855,N_29907,N_29927);
nor UO_1856 (O_1856,N_29817,N_29806);
nand UO_1857 (O_1857,N_29816,N_29971);
and UO_1858 (O_1858,N_29898,N_29939);
nand UO_1859 (O_1859,N_29950,N_29837);
or UO_1860 (O_1860,N_29952,N_29824);
or UO_1861 (O_1861,N_29933,N_29807);
nor UO_1862 (O_1862,N_29961,N_29826);
nor UO_1863 (O_1863,N_29911,N_29923);
xnor UO_1864 (O_1864,N_29907,N_29920);
nand UO_1865 (O_1865,N_29942,N_29965);
nand UO_1866 (O_1866,N_29840,N_29800);
xnor UO_1867 (O_1867,N_29973,N_29946);
nand UO_1868 (O_1868,N_29815,N_29838);
xnor UO_1869 (O_1869,N_29801,N_29890);
or UO_1870 (O_1870,N_29802,N_29931);
or UO_1871 (O_1871,N_29974,N_29844);
or UO_1872 (O_1872,N_29828,N_29861);
nand UO_1873 (O_1873,N_29929,N_29848);
xor UO_1874 (O_1874,N_29869,N_29945);
or UO_1875 (O_1875,N_29883,N_29973);
xnor UO_1876 (O_1876,N_29881,N_29839);
nand UO_1877 (O_1877,N_29847,N_29954);
xnor UO_1878 (O_1878,N_29973,N_29809);
and UO_1879 (O_1879,N_29846,N_29976);
nor UO_1880 (O_1880,N_29937,N_29879);
and UO_1881 (O_1881,N_29944,N_29861);
and UO_1882 (O_1882,N_29874,N_29963);
xor UO_1883 (O_1883,N_29922,N_29947);
nor UO_1884 (O_1884,N_29868,N_29825);
nand UO_1885 (O_1885,N_29907,N_29998);
nand UO_1886 (O_1886,N_29939,N_29964);
and UO_1887 (O_1887,N_29993,N_29800);
xor UO_1888 (O_1888,N_29939,N_29835);
xnor UO_1889 (O_1889,N_29917,N_29978);
or UO_1890 (O_1890,N_29895,N_29882);
and UO_1891 (O_1891,N_29925,N_29878);
nor UO_1892 (O_1892,N_29899,N_29961);
nor UO_1893 (O_1893,N_29875,N_29836);
nand UO_1894 (O_1894,N_29974,N_29827);
nor UO_1895 (O_1895,N_29960,N_29815);
nor UO_1896 (O_1896,N_29808,N_29847);
nand UO_1897 (O_1897,N_29954,N_29807);
or UO_1898 (O_1898,N_29829,N_29906);
and UO_1899 (O_1899,N_29958,N_29830);
nor UO_1900 (O_1900,N_29809,N_29958);
and UO_1901 (O_1901,N_29881,N_29962);
nor UO_1902 (O_1902,N_29989,N_29805);
and UO_1903 (O_1903,N_29815,N_29915);
or UO_1904 (O_1904,N_29851,N_29973);
nand UO_1905 (O_1905,N_29923,N_29928);
and UO_1906 (O_1906,N_29870,N_29890);
and UO_1907 (O_1907,N_29872,N_29864);
or UO_1908 (O_1908,N_29812,N_29937);
nor UO_1909 (O_1909,N_29890,N_29889);
or UO_1910 (O_1910,N_29832,N_29994);
nand UO_1911 (O_1911,N_29999,N_29943);
or UO_1912 (O_1912,N_29804,N_29818);
xor UO_1913 (O_1913,N_29831,N_29919);
and UO_1914 (O_1914,N_29875,N_29866);
and UO_1915 (O_1915,N_29865,N_29922);
nor UO_1916 (O_1916,N_29900,N_29807);
and UO_1917 (O_1917,N_29943,N_29972);
xor UO_1918 (O_1918,N_29969,N_29961);
nand UO_1919 (O_1919,N_29881,N_29936);
xor UO_1920 (O_1920,N_29854,N_29879);
xnor UO_1921 (O_1921,N_29893,N_29963);
and UO_1922 (O_1922,N_29974,N_29869);
nor UO_1923 (O_1923,N_29948,N_29947);
and UO_1924 (O_1924,N_29813,N_29858);
xnor UO_1925 (O_1925,N_29822,N_29961);
or UO_1926 (O_1926,N_29859,N_29926);
or UO_1927 (O_1927,N_29904,N_29962);
or UO_1928 (O_1928,N_29966,N_29884);
xnor UO_1929 (O_1929,N_29999,N_29881);
and UO_1930 (O_1930,N_29811,N_29990);
nand UO_1931 (O_1931,N_29866,N_29862);
and UO_1932 (O_1932,N_29829,N_29899);
or UO_1933 (O_1933,N_29953,N_29991);
and UO_1934 (O_1934,N_29999,N_29929);
nor UO_1935 (O_1935,N_29958,N_29812);
nor UO_1936 (O_1936,N_29924,N_29872);
and UO_1937 (O_1937,N_29965,N_29985);
xor UO_1938 (O_1938,N_29954,N_29988);
xor UO_1939 (O_1939,N_29942,N_29876);
nor UO_1940 (O_1940,N_29973,N_29995);
and UO_1941 (O_1941,N_29985,N_29929);
nor UO_1942 (O_1942,N_29914,N_29843);
nand UO_1943 (O_1943,N_29929,N_29921);
nor UO_1944 (O_1944,N_29901,N_29816);
xnor UO_1945 (O_1945,N_29914,N_29875);
nand UO_1946 (O_1946,N_29939,N_29947);
xor UO_1947 (O_1947,N_29941,N_29851);
xnor UO_1948 (O_1948,N_29903,N_29983);
or UO_1949 (O_1949,N_29857,N_29875);
nand UO_1950 (O_1950,N_29890,N_29805);
nand UO_1951 (O_1951,N_29802,N_29980);
and UO_1952 (O_1952,N_29959,N_29893);
or UO_1953 (O_1953,N_29884,N_29945);
nand UO_1954 (O_1954,N_29983,N_29883);
and UO_1955 (O_1955,N_29951,N_29830);
nor UO_1956 (O_1956,N_29985,N_29815);
nand UO_1957 (O_1957,N_29906,N_29843);
or UO_1958 (O_1958,N_29990,N_29980);
nor UO_1959 (O_1959,N_29820,N_29863);
xnor UO_1960 (O_1960,N_29921,N_29964);
and UO_1961 (O_1961,N_29867,N_29855);
nand UO_1962 (O_1962,N_29875,N_29948);
xor UO_1963 (O_1963,N_29976,N_29861);
xnor UO_1964 (O_1964,N_29939,N_29950);
or UO_1965 (O_1965,N_29881,N_29932);
xnor UO_1966 (O_1966,N_29846,N_29864);
xnor UO_1967 (O_1967,N_29825,N_29939);
and UO_1968 (O_1968,N_29841,N_29876);
or UO_1969 (O_1969,N_29940,N_29826);
and UO_1970 (O_1970,N_29984,N_29893);
or UO_1971 (O_1971,N_29884,N_29971);
and UO_1972 (O_1972,N_29954,N_29959);
nor UO_1973 (O_1973,N_29848,N_29998);
and UO_1974 (O_1974,N_29980,N_29862);
or UO_1975 (O_1975,N_29841,N_29898);
xor UO_1976 (O_1976,N_29967,N_29837);
nor UO_1977 (O_1977,N_29886,N_29986);
or UO_1978 (O_1978,N_29888,N_29820);
and UO_1979 (O_1979,N_29989,N_29835);
xor UO_1980 (O_1980,N_29907,N_29863);
nor UO_1981 (O_1981,N_29815,N_29904);
xnor UO_1982 (O_1982,N_29819,N_29858);
xor UO_1983 (O_1983,N_29813,N_29922);
nand UO_1984 (O_1984,N_29879,N_29866);
or UO_1985 (O_1985,N_29994,N_29951);
xnor UO_1986 (O_1986,N_29818,N_29827);
and UO_1987 (O_1987,N_29963,N_29997);
or UO_1988 (O_1988,N_29932,N_29946);
and UO_1989 (O_1989,N_29920,N_29912);
nand UO_1990 (O_1990,N_29967,N_29995);
and UO_1991 (O_1991,N_29915,N_29997);
or UO_1992 (O_1992,N_29870,N_29971);
nor UO_1993 (O_1993,N_29856,N_29825);
and UO_1994 (O_1994,N_29808,N_29842);
nand UO_1995 (O_1995,N_29943,N_29874);
xnor UO_1996 (O_1996,N_29869,N_29896);
xor UO_1997 (O_1997,N_29885,N_29955);
and UO_1998 (O_1998,N_29952,N_29879);
and UO_1999 (O_1999,N_29847,N_29818);
nor UO_2000 (O_2000,N_29982,N_29921);
or UO_2001 (O_2001,N_29812,N_29971);
or UO_2002 (O_2002,N_29808,N_29952);
nand UO_2003 (O_2003,N_29974,N_29958);
xor UO_2004 (O_2004,N_29997,N_29914);
nand UO_2005 (O_2005,N_29866,N_29810);
xnor UO_2006 (O_2006,N_29835,N_29861);
and UO_2007 (O_2007,N_29836,N_29832);
xnor UO_2008 (O_2008,N_29834,N_29809);
and UO_2009 (O_2009,N_29834,N_29926);
nor UO_2010 (O_2010,N_29846,N_29868);
nand UO_2011 (O_2011,N_29812,N_29947);
nand UO_2012 (O_2012,N_29902,N_29831);
or UO_2013 (O_2013,N_29924,N_29882);
and UO_2014 (O_2014,N_29983,N_29842);
or UO_2015 (O_2015,N_29996,N_29869);
and UO_2016 (O_2016,N_29829,N_29943);
and UO_2017 (O_2017,N_29967,N_29814);
nor UO_2018 (O_2018,N_29983,N_29958);
nand UO_2019 (O_2019,N_29982,N_29936);
xor UO_2020 (O_2020,N_29899,N_29827);
or UO_2021 (O_2021,N_29843,N_29885);
xnor UO_2022 (O_2022,N_29867,N_29883);
xnor UO_2023 (O_2023,N_29830,N_29999);
or UO_2024 (O_2024,N_29937,N_29995);
nand UO_2025 (O_2025,N_29821,N_29850);
or UO_2026 (O_2026,N_29823,N_29897);
nand UO_2027 (O_2027,N_29958,N_29821);
xor UO_2028 (O_2028,N_29932,N_29951);
or UO_2029 (O_2029,N_29989,N_29848);
xnor UO_2030 (O_2030,N_29942,N_29926);
or UO_2031 (O_2031,N_29935,N_29983);
and UO_2032 (O_2032,N_29947,N_29889);
xnor UO_2033 (O_2033,N_29920,N_29951);
and UO_2034 (O_2034,N_29856,N_29857);
nand UO_2035 (O_2035,N_29977,N_29951);
nor UO_2036 (O_2036,N_29951,N_29926);
nor UO_2037 (O_2037,N_29852,N_29942);
or UO_2038 (O_2038,N_29804,N_29977);
nand UO_2039 (O_2039,N_29899,N_29855);
xnor UO_2040 (O_2040,N_29841,N_29867);
nand UO_2041 (O_2041,N_29893,N_29923);
and UO_2042 (O_2042,N_29899,N_29923);
xnor UO_2043 (O_2043,N_29984,N_29866);
xnor UO_2044 (O_2044,N_29942,N_29951);
nor UO_2045 (O_2045,N_29981,N_29965);
nor UO_2046 (O_2046,N_29831,N_29891);
xor UO_2047 (O_2047,N_29891,N_29920);
nand UO_2048 (O_2048,N_29833,N_29928);
xor UO_2049 (O_2049,N_29873,N_29851);
or UO_2050 (O_2050,N_29883,N_29978);
and UO_2051 (O_2051,N_29972,N_29879);
nand UO_2052 (O_2052,N_29870,N_29813);
or UO_2053 (O_2053,N_29820,N_29806);
nand UO_2054 (O_2054,N_29834,N_29888);
nor UO_2055 (O_2055,N_29908,N_29849);
nor UO_2056 (O_2056,N_29971,N_29980);
and UO_2057 (O_2057,N_29919,N_29917);
xnor UO_2058 (O_2058,N_29896,N_29885);
and UO_2059 (O_2059,N_29803,N_29813);
and UO_2060 (O_2060,N_29840,N_29895);
and UO_2061 (O_2061,N_29918,N_29821);
nand UO_2062 (O_2062,N_29868,N_29860);
xnor UO_2063 (O_2063,N_29833,N_29981);
nand UO_2064 (O_2064,N_29825,N_29914);
xor UO_2065 (O_2065,N_29908,N_29915);
and UO_2066 (O_2066,N_29911,N_29984);
xnor UO_2067 (O_2067,N_29945,N_29956);
and UO_2068 (O_2068,N_29808,N_29878);
or UO_2069 (O_2069,N_29973,N_29853);
xor UO_2070 (O_2070,N_29935,N_29810);
and UO_2071 (O_2071,N_29853,N_29818);
or UO_2072 (O_2072,N_29895,N_29935);
xnor UO_2073 (O_2073,N_29857,N_29965);
nor UO_2074 (O_2074,N_29881,N_29988);
nor UO_2075 (O_2075,N_29947,N_29920);
nand UO_2076 (O_2076,N_29815,N_29947);
and UO_2077 (O_2077,N_29942,N_29916);
nand UO_2078 (O_2078,N_29894,N_29953);
and UO_2079 (O_2079,N_29802,N_29908);
or UO_2080 (O_2080,N_29873,N_29904);
xnor UO_2081 (O_2081,N_29917,N_29935);
xor UO_2082 (O_2082,N_29850,N_29855);
and UO_2083 (O_2083,N_29996,N_29826);
xnor UO_2084 (O_2084,N_29881,N_29821);
nor UO_2085 (O_2085,N_29860,N_29949);
xnor UO_2086 (O_2086,N_29986,N_29983);
or UO_2087 (O_2087,N_29956,N_29962);
nor UO_2088 (O_2088,N_29887,N_29839);
xnor UO_2089 (O_2089,N_29817,N_29915);
and UO_2090 (O_2090,N_29925,N_29961);
nand UO_2091 (O_2091,N_29964,N_29845);
or UO_2092 (O_2092,N_29870,N_29800);
or UO_2093 (O_2093,N_29896,N_29892);
nor UO_2094 (O_2094,N_29851,N_29946);
and UO_2095 (O_2095,N_29961,N_29827);
nand UO_2096 (O_2096,N_29862,N_29948);
nor UO_2097 (O_2097,N_29803,N_29919);
or UO_2098 (O_2098,N_29860,N_29920);
and UO_2099 (O_2099,N_29863,N_29943);
nand UO_2100 (O_2100,N_29872,N_29904);
and UO_2101 (O_2101,N_29839,N_29873);
and UO_2102 (O_2102,N_29850,N_29851);
nor UO_2103 (O_2103,N_29998,N_29946);
nor UO_2104 (O_2104,N_29954,N_29838);
and UO_2105 (O_2105,N_29892,N_29987);
or UO_2106 (O_2106,N_29893,N_29842);
or UO_2107 (O_2107,N_29823,N_29869);
nor UO_2108 (O_2108,N_29875,N_29819);
nor UO_2109 (O_2109,N_29804,N_29948);
and UO_2110 (O_2110,N_29973,N_29935);
or UO_2111 (O_2111,N_29948,N_29961);
or UO_2112 (O_2112,N_29952,N_29936);
nand UO_2113 (O_2113,N_29971,N_29924);
xnor UO_2114 (O_2114,N_29957,N_29914);
xor UO_2115 (O_2115,N_29927,N_29855);
nand UO_2116 (O_2116,N_29929,N_29950);
nand UO_2117 (O_2117,N_29807,N_29803);
or UO_2118 (O_2118,N_29937,N_29824);
xor UO_2119 (O_2119,N_29875,N_29861);
nand UO_2120 (O_2120,N_29968,N_29898);
or UO_2121 (O_2121,N_29846,N_29839);
and UO_2122 (O_2122,N_29858,N_29988);
xor UO_2123 (O_2123,N_29942,N_29890);
nand UO_2124 (O_2124,N_29904,N_29942);
nand UO_2125 (O_2125,N_29844,N_29869);
nand UO_2126 (O_2126,N_29829,N_29894);
nand UO_2127 (O_2127,N_29996,N_29973);
nor UO_2128 (O_2128,N_29970,N_29814);
and UO_2129 (O_2129,N_29925,N_29939);
and UO_2130 (O_2130,N_29847,N_29963);
nor UO_2131 (O_2131,N_29901,N_29850);
nand UO_2132 (O_2132,N_29940,N_29952);
nand UO_2133 (O_2133,N_29911,N_29816);
or UO_2134 (O_2134,N_29904,N_29870);
nand UO_2135 (O_2135,N_29861,N_29926);
nand UO_2136 (O_2136,N_29832,N_29972);
nor UO_2137 (O_2137,N_29989,N_29921);
or UO_2138 (O_2138,N_29823,N_29961);
or UO_2139 (O_2139,N_29855,N_29849);
and UO_2140 (O_2140,N_29844,N_29978);
xor UO_2141 (O_2141,N_29922,N_29877);
nand UO_2142 (O_2142,N_29814,N_29996);
or UO_2143 (O_2143,N_29977,N_29956);
and UO_2144 (O_2144,N_29981,N_29878);
or UO_2145 (O_2145,N_29820,N_29889);
xnor UO_2146 (O_2146,N_29890,N_29854);
or UO_2147 (O_2147,N_29915,N_29858);
nor UO_2148 (O_2148,N_29969,N_29837);
and UO_2149 (O_2149,N_29837,N_29938);
nor UO_2150 (O_2150,N_29950,N_29912);
or UO_2151 (O_2151,N_29847,N_29977);
or UO_2152 (O_2152,N_29851,N_29944);
and UO_2153 (O_2153,N_29894,N_29830);
nand UO_2154 (O_2154,N_29967,N_29990);
nor UO_2155 (O_2155,N_29834,N_29837);
or UO_2156 (O_2156,N_29860,N_29848);
nor UO_2157 (O_2157,N_29994,N_29898);
nand UO_2158 (O_2158,N_29920,N_29980);
nand UO_2159 (O_2159,N_29901,N_29973);
or UO_2160 (O_2160,N_29997,N_29995);
nand UO_2161 (O_2161,N_29927,N_29969);
and UO_2162 (O_2162,N_29805,N_29848);
xnor UO_2163 (O_2163,N_29836,N_29860);
nand UO_2164 (O_2164,N_29876,N_29916);
or UO_2165 (O_2165,N_29838,N_29840);
nor UO_2166 (O_2166,N_29804,N_29978);
or UO_2167 (O_2167,N_29806,N_29998);
nand UO_2168 (O_2168,N_29831,N_29837);
nor UO_2169 (O_2169,N_29880,N_29902);
and UO_2170 (O_2170,N_29973,N_29920);
or UO_2171 (O_2171,N_29990,N_29983);
and UO_2172 (O_2172,N_29813,N_29818);
nor UO_2173 (O_2173,N_29921,N_29999);
nor UO_2174 (O_2174,N_29979,N_29806);
nor UO_2175 (O_2175,N_29922,N_29896);
nand UO_2176 (O_2176,N_29814,N_29880);
or UO_2177 (O_2177,N_29830,N_29913);
and UO_2178 (O_2178,N_29932,N_29824);
xor UO_2179 (O_2179,N_29927,N_29866);
or UO_2180 (O_2180,N_29937,N_29828);
or UO_2181 (O_2181,N_29913,N_29926);
xnor UO_2182 (O_2182,N_29929,N_29916);
or UO_2183 (O_2183,N_29831,N_29930);
xnor UO_2184 (O_2184,N_29901,N_29972);
nor UO_2185 (O_2185,N_29852,N_29846);
and UO_2186 (O_2186,N_29895,N_29929);
xor UO_2187 (O_2187,N_29866,N_29856);
nand UO_2188 (O_2188,N_29853,N_29807);
or UO_2189 (O_2189,N_29814,N_29819);
xnor UO_2190 (O_2190,N_29993,N_29900);
or UO_2191 (O_2191,N_29931,N_29845);
nor UO_2192 (O_2192,N_29936,N_29894);
nor UO_2193 (O_2193,N_29889,N_29977);
and UO_2194 (O_2194,N_29895,N_29811);
xnor UO_2195 (O_2195,N_29890,N_29827);
xor UO_2196 (O_2196,N_29846,N_29841);
nor UO_2197 (O_2197,N_29838,N_29971);
nor UO_2198 (O_2198,N_29932,N_29913);
and UO_2199 (O_2199,N_29802,N_29953);
xnor UO_2200 (O_2200,N_29972,N_29865);
nand UO_2201 (O_2201,N_29950,N_29854);
xor UO_2202 (O_2202,N_29959,N_29961);
nor UO_2203 (O_2203,N_29998,N_29947);
nor UO_2204 (O_2204,N_29817,N_29885);
and UO_2205 (O_2205,N_29966,N_29956);
or UO_2206 (O_2206,N_29860,N_29987);
or UO_2207 (O_2207,N_29937,N_29980);
nor UO_2208 (O_2208,N_29989,N_29936);
nand UO_2209 (O_2209,N_29994,N_29963);
xnor UO_2210 (O_2210,N_29807,N_29941);
xnor UO_2211 (O_2211,N_29891,N_29814);
nor UO_2212 (O_2212,N_29972,N_29962);
xnor UO_2213 (O_2213,N_29885,N_29916);
and UO_2214 (O_2214,N_29811,N_29881);
nand UO_2215 (O_2215,N_29890,N_29969);
xor UO_2216 (O_2216,N_29891,N_29858);
or UO_2217 (O_2217,N_29918,N_29802);
or UO_2218 (O_2218,N_29833,N_29899);
xor UO_2219 (O_2219,N_29987,N_29806);
nor UO_2220 (O_2220,N_29916,N_29936);
nor UO_2221 (O_2221,N_29984,N_29900);
or UO_2222 (O_2222,N_29966,N_29989);
xor UO_2223 (O_2223,N_29941,N_29874);
nor UO_2224 (O_2224,N_29991,N_29802);
nor UO_2225 (O_2225,N_29804,N_29974);
nand UO_2226 (O_2226,N_29953,N_29942);
xor UO_2227 (O_2227,N_29986,N_29800);
nor UO_2228 (O_2228,N_29809,N_29864);
nand UO_2229 (O_2229,N_29942,N_29811);
nand UO_2230 (O_2230,N_29851,N_29964);
nor UO_2231 (O_2231,N_29972,N_29922);
nor UO_2232 (O_2232,N_29948,N_29912);
nand UO_2233 (O_2233,N_29837,N_29986);
and UO_2234 (O_2234,N_29932,N_29925);
or UO_2235 (O_2235,N_29954,N_29879);
nand UO_2236 (O_2236,N_29912,N_29988);
nor UO_2237 (O_2237,N_29974,N_29807);
nor UO_2238 (O_2238,N_29861,N_29957);
xnor UO_2239 (O_2239,N_29824,N_29864);
xnor UO_2240 (O_2240,N_29821,N_29861);
or UO_2241 (O_2241,N_29982,N_29981);
nor UO_2242 (O_2242,N_29896,N_29881);
nand UO_2243 (O_2243,N_29966,N_29866);
nor UO_2244 (O_2244,N_29921,N_29991);
and UO_2245 (O_2245,N_29916,N_29806);
xnor UO_2246 (O_2246,N_29824,N_29929);
and UO_2247 (O_2247,N_29997,N_29800);
nor UO_2248 (O_2248,N_29818,N_29943);
nand UO_2249 (O_2249,N_29844,N_29877);
nor UO_2250 (O_2250,N_29862,N_29853);
xor UO_2251 (O_2251,N_29889,N_29874);
or UO_2252 (O_2252,N_29947,N_29973);
and UO_2253 (O_2253,N_29917,N_29811);
xnor UO_2254 (O_2254,N_29971,N_29814);
xnor UO_2255 (O_2255,N_29963,N_29950);
and UO_2256 (O_2256,N_29990,N_29998);
and UO_2257 (O_2257,N_29890,N_29803);
or UO_2258 (O_2258,N_29842,N_29920);
nand UO_2259 (O_2259,N_29917,N_29928);
xor UO_2260 (O_2260,N_29923,N_29991);
nand UO_2261 (O_2261,N_29881,N_29840);
or UO_2262 (O_2262,N_29824,N_29819);
or UO_2263 (O_2263,N_29837,N_29916);
and UO_2264 (O_2264,N_29946,N_29839);
and UO_2265 (O_2265,N_29848,N_29956);
or UO_2266 (O_2266,N_29952,N_29911);
or UO_2267 (O_2267,N_29973,N_29837);
xnor UO_2268 (O_2268,N_29952,N_29833);
or UO_2269 (O_2269,N_29927,N_29870);
and UO_2270 (O_2270,N_29868,N_29806);
xnor UO_2271 (O_2271,N_29961,N_29878);
xor UO_2272 (O_2272,N_29802,N_29937);
nor UO_2273 (O_2273,N_29829,N_29861);
nor UO_2274 (O_2274,N_29901,N_29984);
nor UO_2275 (O_2275,N_29996,N_29887);
or UO_2276 (O_2276,N_29817,N_29893);
xor UO_2277 (O_2277,N_29828,N_29872);
xor UO_2278 (O_2278,N_29925,N_29851);
and UO_2279 (O_2279,N_29851,N_29804);
and UO_2280 (O_2280,N_29870,N_29985);
nor UO_2281 (O_2281,N_29853,N_29985);
nand UO_2282 (O_2282,N_29900,N_29876);
xnor UO_2283 (O_2283,N_29802,N_29891);
or UO_2284 (O_2284,N_29830,N_29885);
xnor UO_2285 (O_2285,N_29990,N_29918);
xnor UO_2286 (O_2286,N_29974,N_29836);
xnor UO_2287 (O_2287,N_29950,N_29856);
xor UO_2288 (O_2288,N_29946,N_29842);
or UO_2289 (O_2289,N_29933,N_29973);
xnor UO_2290 (O_2290,N_29806,N_29997);
nand UO_2291 (O_2291,N_29853,N_29833);
and UO_2292 (O_2292,N_29980,N_29829);
xor UO_2293 (O_2293,N_29991,N_29927);
or UO_2294 (O_2294,N_29873,N_29888);
xor UO_2295 (O_2295,N_29818,N_29807);
xnor UO_2296 (O_2296,N_29859,N_29996);
nor UO_2297 (O_2297,N_29856,N_29986);
nand UO_2298 (O_2298,N_29907,N_29801);
nor UO_2299 (O_2299,N_29871,N_29863);
and UO_2300 (O_2300,N_29832,N_29854);
xnor UO_2301 (O_2301,N_29910,N_29920);
nor UO_2302 (O_2302,N_29972,N_29827);
nor UO_2303 (O_2303,N_29814,N_29954);
nor UO_2304 (O_2304,N_29929,N_29882);
nand UO_2305 (O_2305,N_29978,N_29941);
or UO_2306 (O_2306,N_29810,N_29892);
and UO_2307 (O_2307,N_29884,N_29949);
and UO_2308 (O_2308,N_29955,N_29892);
and UO_2309 (O_2309,N_29831,N_29976);
xnor UO_2310 (O_2310,N_29917,N_29837);
nor UO_2311 (O_2311,N_29895,N_29940);
or UO_2312 (O_2312,N_29939,N_29870);
nand UO_2313 (O_2313,N_29827,N_29832);
and UO_2314 (O_2314,N_29933,N_29844);
or UO_2315 (O_2315,N_29988,N_29962);
xnor UO_2316 (O_2316,N_29888,N_29957);
nor UO_2317 (O_2317,N_29999,N_29864);
and UO_2318 (O_2318,N_29996,N_29813);
nor UO_2319 (O_2319,N_29924,N_29830);
or UO_2320 (O_2320,N_29862,N_29999);
or UO_2321 (O_2321,N_29894,N_29935);
nor UO_2322 (O_2322,N_29839,N_29977);
nand UO_2323 (O_2323,N_29893,N_29944);
and UO_2324 (O_2324,N_29825,N_29812);
and UO_2325 (O_2325,N_29877,N_29970);
and UO_2326 (O_2326,N_29853,N_29932);
or UO_2327 (O_2327,N_29811,N_29890);
xnor UO_2328 (O_2328,N_29987,N_29999);
or UO_2329 (O_2329,N_29958,N_29905);
nand UO_2330 (O_2330,N_29985,N_29861);
and UO_2331 (O_2331,N_29857,N_29981);
nand UO_2332 (O_2332,N_29871,N_29830);
or UO_2333 (O_2333,N_29961,N_29993);
and UO_2334 (O_2334,N_29968,N_29992);
nand UO_2335 (O_2335,N_29952,N_29993);
nor UO_2336 (O_2336,N_29981,N_29806);
nand UO_2337 (O_2337,N_29917,N_29859);
or UO_2338 (O_2338,N_29941,N_29907);
nor UO_2339 (O_2339,N_29803,N_29993);
and UO_2340 (O_2340,N_29947,N_29835);
nor UO_2341 (O_2341,N_29831,N_29867);
nand UO_2342 (O_2342,N_29820,N_29913);
or UO_2343 (O_2343,N_29833,N_29824);
xor UO_2344 (O_2344,N_29814,N_29875);
or UO_2345 (O_2345,N_29828,N_29838);
nand UO_2346 (O_2346,N_29915,N_29921);
nor UO_2347 (O_2347,N_29970,N_29943);
and UO_2348 (O_2348,N_29837,N_29952);
xnor UO_2349 (O_2349,N_29917,N_29830);
nand UO_2350 (O_2350,N_29956,N_29886);
and UO_2351 (O_2351,N_29893,N_29945);
xor UO_2352 (O_2352,N_29944,N_29911);
nand UO_2353 (O_2353,N_29808,N_29826);
xor UO_2354 (O_2354,N_29862,N_29921);
nor UO_2355 (O_2355,N_29818,N_29881);
and UO_2356 (O_2356,N_29828,N_29829);
xor UO_2357 (O_2357,N_29815,N_29919);
xnor UO_2358 (O_2358,N_29885,N_29928);
xor UO_2359 (O_2359,N_29846,N_29837);
nand UO_2360 (O_2360,N_29981,N_29945);
or UO_2361 (O_2361,N_29901,N_29982);
and UO_2362 (O_2362,N_29955,N_29856);
nor UO_2363 (O_2363,N_29867,N_29876);
or UO_2364 (O_2364,N_29846,N_29880);
xor UO_2365 (O_2365,N_29881,N_29899);
nor UO_2366 (O_2366,N_29921,N_29950);
nand UO_2367 (O_2367,N_29822,N_29833);
xnor UO_2368 (O_2368,N_29971,N_29888);
xnor UO_2369 (O_2369,N_29991,N_29899);
and UO_2370 (O_2370,N_29854,N_29909);
and UO_2371 (O_2371,N_29889,N_29955);
xnor UO_2372 (O_2372,N_29801,N_29805);
nand UO_2373 (O_2373,N_29984,N_29840);
nand UO_2374 (O_2374,N_29813,N_29915);
xor UO_2375 (O_2375,N_29964,N_29980);
nand UO_2376 (O_2376,N_29974,N_29975);
and UO_2377 (O_2377,N_29916,N_29858);
or UO_2378 (O_2378,N_29883,N_29901);
or UO_2379 (O_2379,N_29854,N_29939);
xnor UO_2380 (O_2380,N_29952,N_29801);
nor UO_2381 (O_2381,N_29837,N_29830);
or UO_2382 (O_2382,N_29963,N_29864);
or UO_2383 (O_2383,N_29829,N_29930);
xor UO_2384 (O_2384,N_29825,N_29887);
xor UO_2385 (O_2385,N_29838,N_29992);
nor UO_2386 (O_2386,N_29859,N_29836);
nand UO_2387 (O_2387,N_29978,N_29918);
nand UO_2388 (O_2388,N_29945,N_29806);
xnor UO_2389 (O_2389,N_29949,N_29924);
xor UO_2390 (O_2390,N_29959,N_29955);
or UO_2391 (O_2391,N_29928,N_29945);
xnor UO_2392 (O_2392,N_29932,N_29875);
nor UO_2393 (O_2393,N_29948,N_29927);
and UO_2394 (O_2394,N_29978,N_29814);
xnor UO_2395 (O_2395,N_29960,N_29964);
nand UO_2396 (O_2396,N_29990,N_29890);
nand UO_2397 (O_2397,N_29815,N_29903);
nor UO_2398 (O_2398,N_29929,N_29815);
nand UO_2399 (O_2399,N_29824,N_29908);
xnor UO_2400 (O_2400,N_29912,N_29938);
or UO_2401 (O_2401,N_29891,N_29958);
nor UO_2402 (O_2402,N_29991,N_29889);
or UO_2403 (O_2403,N_29839,N_29855);
nor UO_2404 (O_2404,N_29823,N_29885);
or UO_2405 (O_2405,N_29838,N_29938);
or UO_2406 (O_2406,N_29829,N_29817);
and UO_2407 (O_2407,N_29856,N_29869);
and UO_2408 (O_2408,N_29816,N_29872);
xor UO_2409 (O_2409,N_29961,N_29883);
or UO_2410 (O_2410,N_29933,N_29992);
nand UO_2411 (O_2411,N_29922,N_29961);
or UO_2412 (O_2412,N_29889,N_29860);
and UO_2413 (O_2413,N_29898,N_29911);
nand UO_2414 (O_2414,N_29994,N_29962);
or UO_2415 (O_2415,N_29866,N_29997);
nor UO_2416 (O_2416,N_29804,N_29963);
or UO_2417 (O_2417,N_29899,N_29929);
xor UO_2418 (O_2418,N_29833,N_29887);
or UO_2419 (O_2419,N_29934,N_29913);
or UO_2420 (O_2420,N_29841,N_29988);
nand UO_2421 (O_2421,N_29898,N_29922);
or UO_2422 (O_2422,N_29987,N_29827);
nand UO_2423 (O_2423,N_29880,N_29804);
xnor UO_2424 (O_2424,N_29928,N_29964);
nor UO_2425 (O_2425,N_29803,N_29978);
and UO_2426 (O_2426,N_29942,N_29972);
nor UO_2427 (O_2427,N_29971,N_29821);
and UO_2428 (O_2428,N_29991,N_29948);
or UO_2429 (O_2429,N_29938,N_29982);
nand UO_2430 (O_2430,N_29884,N_29917);
nand UO_2431 (O_2431,N_29892,N_29847);
nor UO_2432 (O_2432,N_29977,N_29880);
and UO_2433 (O_2433,N_29818,N_29986);
or UO_2434 (O_2434,N_29862,N_29885);
and UO_2435 (O_2435,N_29940,N_29945);
xor UO_2436 (O_2436,N_29945,N_29931);
and UO_2437 (O_2437,N_29956,N_29850);
nand UO_2438 (O_2438,N_29870,N_29968);
xor UO_2439 (O_2439,N_29854,N_29861);
or UO_2440 (O_2440,N_29887,N_29823);
nand UO_2441 (O_2441,N_29803,N_29806);
or UO_2442 (O_2442,N_29935,N_29908);
nor UO_2443 (O_2443,N_29958,N_29846);
and UO_2444 (O_2444,N_29991,N_29958);
nor UO_2445 (O_2445,N_29824,N_29898);
xnor UO_2446 (O_2446,N_29972,N_29916);
and UO_2447 (O_2447,N_29989,N_29947);
nor UO_2448 (O_2448,N_29888,N_29826);
or UO_2449 (O_2449,N_29877,N_29860);
and UO_2450 (O_2450,N_29986,N_29803);
and UO_2451 (O_2451,N_29911,N_29964);
xnor UO_2452 (O_2452,N_29985,N_29899);
nand UO_2453 (O_2453,N_29902,N_29944);
or UO_2454 (O_2454,N_29947,N_29877);
and UO_2455 (O_2455,N_29845,N_29881);
and UO_2456 (O_2456,N_29903,N_29901);
or UO_2457 (O_2457,N_29857,N_29947);
nor UO_2458 (O_2458,N_29952,N_29825);
nor UO_2459 (O_2459,N_29839,N_29972);
xor UO_2460 (O_2460,N_29901,N_29880);
or UO_2461 (O_2461,N_29905,N_29818);
or UO_2462 (O_2462,N_29820,N_29827);
and UO_2463 (O_2463,N_29837,N_29860);
nand UO_2464 (O_2464,N_29864,N_29868);
nand UO_2465 (O_2465,N_29915,N_29847);
and UO_2466 (O_2466,N_29932,N_29825);
nand UO_2467 (O_2467,N_29925,N_29897);
nor UO_2468 (O_2468,N_29801,N_29883);
or UO_2469 (O_2469,N_29966,N_29856);
and UO_2470 (O_2470,N_29887,N_29859);
and UO_2471 (O_2471,N_29965,N_29904);
nor UO_2472 (O_2472,N_29951,N_29991);
or UO_2473 (O_2473,N_29953,N_29958);
and UO_2474 (O_2474,N_29981,N_29854);
nor UO_2475 (O_2475,N_29952,N_29838);
and UO_2476 (O_2476,N_29961,N_29845);
nor UO_2477 (O_2477,N_29924,N_29982);
nor UO_2478 (O_2478,N_29853,N_29943);
or UO_2479 (O_2479,N_29834,N_29882);
or UO_2480 (O_2480,N_29849,N_29895);
xnor UO_2481 (O_2481,N_29989,N_29919);
nand UO_2482 (O_2482,N_29973,N_29904);
nand UO_2483 (O_2483,N_29828,N_29997);
nor UO_2484 (O_2484,N_29866,N_29881);
nand UO_2485 (O_2485,N_29837,N_29915);
xnor UO_2486 (O_2486,N_29892,N_29849);
and UO_2487 (O_2487,N_29804,N_29869);
and UO_2488 (O_2488,N_29867,N_29888);
and UO_2489 (O_2489,N_29868,N_29944);
xor UO_2490 (O_2490,N_29826,N_29991);
xor UO_2491 (O_2491,N_29958,N_29955);
xor UO_2492 (O_2492,N_29894,N_29897);
or UO_2493 (O_2493,N_29965,N_29809);
nand UO_2494 (O_2494,N_29943,N_29964);
and UO_2495 (O_2495,N_29900,N_29971);
or UO_2496 (O_2496,N_29826,N_29875);
nor UO_2497 (O_2497,N_29914,N_29910);
or UO_2498 (O_2498,N_29807,N_29949);
nand UO_2499 (O_2499,N_29935,N_29806);
and UO_2500 (O_2500,N_29862,N_29981);
and UO_2501 (O_2501,N_29968,N_29937);
and UO_2502 (O_2502,N_29854,N_29960);
nor UO_2503 (O_2503,N_29883,N_29812);
nor UO_2504 (O_2504,N_29959,N_29844);
nor UO_2505 (O_2505,N_29808,N_29810);
or UO_2506 (O_2506,N_29809,N_29856);
nand UO_2507 (O_2507,N_29962,N_29892);
and UO_2508 (O_2508,N_29882,N_29986);
nor UO_2509 (O_2509,N_29929,N_29926);
xnor UO_2510 (O_2510,N_29958,N_29939);
nand UO_2511 (O_2511,N_29835,N_29870);
nand UO_2512 (O_2512,N_29825,N_29910);
nand UO_2513 (O_2513,N_29858,N_29990);
nand UO_2514 (O_2514,N_29919,N_29827);
and UO_2515 (O_2515,N_29896,N_29868);
and UO_2516 (O_2516,N_29990,N_29987);
xor UO_2517 (O_2517,N_29889,N_29872);
and UO_2518 (O_2518,N_29975,N_29889);
nand UO_2519 (O_2519,N_29963,N_29881);
nand UO_2520 (O_2520,N_29887,N_29810);
xnor UO_2521 (O_2521,N_29965,N_29957);
nand UO_2522 (O_2522,N_29803,N_29908);
or UO_2523 (O_2523,N_29864,N_29990);
nor UO_2524 (O_2524,N_29916,N_29905);
nand UO_2525 (O_2525,N_29807,N_29971);
or UO_2526 (O_2526,N_29822,N_29984);
xnor UO_2527 (O_2527,N_29882,N_29954);
nand UO_2528 (O_2528,N_29912,N_29883);
nor UO_2529 (O_2529,N_29845,N_29807);
nor UO_2530 (O_2530,N_29988,N_29966);
nor UO_2531 (O_2531,N_29917,N_29842);
xor UO_2532 (O_2532,N_29886,N_29926);
nor UO_2533 (O_2533,N_29999,N_29968);
or UO_2534 (O_2534,N_29946,N_29806);
nor UO_2535 (O_2535,N_29987,N_29881);
nand UO_2536 (O_2536,N_29905,N_29935);
xnor UO_2537 (O_2537,N_29852,N_29900);
or UO_2538 (O_2538,N_29881,N_29807);
nand UO_2539 (O_2539,N_29969,N_29856);
nor UO_2540 (O_2540,N_29954,N_29950);
nand UO_2541 (O_2541,N_29954,N_29924);
or UO_2542 (O_2542,N_29867,N_29866);
nand UO_2543 (O_2543,N_29930,N_29892);
nand UO_2544 (O_2544,N_29876,N_29877);
and UO_2545 (O_2545,N_29854,N_29965);
or UO_2546 (O_2546,N_29802,N_29967);
or UO_2547 (O_2547,N_29960,N_29901);
xnor UO_2548 (O_2548,N_29890,N_29992);
or UO_2549 (O_2549,N_29807,N_29916);
xor UO_2550 (O_2550,N_29891,N_29821);
nor UO_2551 (O_2551,N_29996,N_29950);
xor UO_2552 (O_2552,N_29886,N_29874);
xor UO_2553 (O_2553,N_29815,N_29961);
nand UO_2554 (O_2554,N_29847,N_29922);
nand UO_2555 (O_2555,N_29957,N_29949);
or UO_2556 (O_2556,N_29971,N_29933);
nand UO_2557 (O_2557,N_29820,N_29958);
and UO_2558 (O_2558,N_29855,N_29926);
xor UO_2559 (O_2559,N_29855,N_29864);
xor UO_2560 (O_2560,N_29848,N_29965);
and UO_2561 (O_2561,N_29825,N_29845);
and UO_2562 (O_2562,N_29991,N_29875);
xnor UO_2563 (O_2563,N_29885,N_29918);
nor UO_2564 (O_2564,N_29872,N_29878);
or UO_2565 (O_2565,N_29976,N_29909);
xor UO_2566 (O_2566,N_29977,N_29968);
xor UO_2567 (O_2567,N_29978,N_29846);
nor UO_2568 (O_2568,N_29993,N_29917);
nand UO_2569 (O_2569,N_29850,N_29869);
or UO_2570 (O_2570,N_29949,N_29872);
xor UO_2571 (O_2571,N_29877,N_29868);
nor UO_2572 (O_2572,N_29990,N_29949);
or UO_2573 (O_2573,N_29917,N_29879);
or UO_2574 (O_2574,N_29964,N_29875);
or UO_2575 (O_2575,N_29900,N_29821);
nor UO_2576 (O_2576,N_29883,N_29929);
nor UO_2577 (O_2577,N_29984,N_29976);
or UO_2578 (O_2578,N_29981,N_29996);
and UO_2579 (O_2579,N_29803,N_29814);
or UO_2580 (O_2580,N_29982,N_29944);
xor UO_2581 (O_2581,N_29859,N_29862);
and UO_2582 (O_2582,N_29996,N_29959);
nor UO_2583 (O_2583,N_29953,N_29996);
and UO_2584 (O_2584,N_29816,N_29978);
xnor UO_2585 (O_2585,N_29862,N_29889);
nor UO_2586 (O_2586,N_29892,N_29903);
and UO_2587 (O_2587,N_29938,N_29996);
nor UO_2588 (O_2588,N_29996,N_29855);
nor UO_2589 (O_2589,N_29835,N_29855);
or UO_2590 (O_2590,N_29849,N_29888);
nand UO_2591 (O_2591,N_29996,N_29805);
nand UO_2592 (O_2592,N_29925,N_29907);
nor UO_2593 (O_2593,N_29861,N_29998);
or UO_2594 (O_2594,N_29893,N_29824);
or UO_2595 (O_2595,N_29848,N_29801);
or UO_2596 (O_2596,N_29922,N_29857);
and UO_2597 (O_2597,N_29931,N_29901);
nand UO_2598 (O_2598,N_29846,N_29828);
and UO_2599 (O_2599,N_29801,N_29860);
and UO_2600 (O_2600,N_29991,N_29936);
or UO_2601 (O_2601,N_29909,N_29889);
or UO_2602 (O_2602,N_29840,N_29813);
and UO_2603 (O_2603,N_29991,N_29957);
xor UO_2604 (O_2604,N_29984,N_29982);
nor UO_2605 (O_2605,N_29936,N_29900);
and UO_2606 (O_2606,N_29882,N_29873);
nor UO_2607 (O_2607,N_29830,N_29963);
nor UO_2608 (O_2608,N_29856,N_29841);
nand UO_2609 (O_2609,N_29917,N_29927);
and UO_2610 (O_2610,N_29969,N_29810);
and UO_2611 (O_2611,N_29987,N_29946);
and UO_2612 (O_2612,N_29978,N_29892);
nor UO_2613 (O_2613,N_29982,N_29876);
nor UO_2614 (O_2614,N_29844,N_29900);
nor UO_2615 (O_2615,N_29947,N_29905);
nor UO_2616 (O_2616,N_29904,N_29913);
nand UO_2617 (O_2617,N_29921,N_29981);
nor UO_2618 (O_2618,N_29861,N_29857);
nor UO_2619 (O_2619,N_29875,N_29949);
xor UO_2620 (O_2620,N_29918,N_29825);
xor UO_2621 (O_2621,N_29959,N_29897);
xor UO_2622 (O_2622,N_29806,N_29983);
or UO_2623 (O_2623,N_29865,N_29977);
or UO_2624 (O_2624,N_29844,N_29816);
nor UO_2625 (O_2625,N_29811,N_29869);
nand UO_2626 (O_2626,N_29827,N_29878);
xor UO_2627 (O_2627,N_29923,N_29800);
nor UO_2628 (O_2628,N_29977,N_29853);
or UO_2629 (O_2629,N_29815,N_29992);
nor UO_2630 (O_2630,N_29877,N_29842);
xor UO_2631 (O_2631,N_29859,N_29875);
and UO_2632 (O_2632,N_29914,N_29802);
or UO_2633 (O_2633,N_29895,N_29865);
and UO_2634 (O_2634,N_29982,N_29929);
or UO_2635 (O_2635,N_29923,N_29963);
nor UO_2636 (O_2636,N_29816,N_29867);
and UO_2637 (O_2637,N_29831,N_29986);
or UO_2638 (O_2638,N_29824,N_29882);
nor UO_2639 (O_2639,N_29927,N_29963);
nand UO_2640 (O_2640,N_29949,N_29953);
nor UO_2641 (O_2641,N_29995,N_29892);
and UO_2642 (O_2642,N_29865,N_29805);
nor UO_2643 (O_2643,N_29820,N_29845);
xor UO_2644 (O_2644,N_29882,N_29917);
nor UO_2645 (O_2645,N_29911,N_29947);
and UO_2646 (O_2646,N_29973,N_29943);
nand UO_2647 (O_2647,N_29875,N_29945);
nor UO_2648 (O_2648,N_29811,N_29999);
or UO_2649 (O_2649,N_29933,N_29907);
and UO_2650 (O_2650,N_29826,N_29916);
and UO_2651 (O_2651,N_29876,N_29920);
nand UO_2652 (O_2652,N_29896,N_29954);
xnor UO_2653 (O_2653,N_29899,N_29990);
nor UO_2654 (O_2654,N_29962,N_29878);
and UO_2655 (O_2655,N_29946,N_29909);
nand UO_2656 (O_2656,N_29967,N_29993);
xor UO_2657 (O_2657,N_29921,N_29844);
or UO_2658 (O_2658,N_29865,N_29803);
or UO_2659 (O_2659,N_29961,N_29835);
xor UO_2660 (O_2660,N_29966,N_29844);
and UO_2661 (O_2661,N_29845,N_29829);
nor UO_2662 (O_2662,N_29880,N_29913);
xnor UO_2663 (O_2663,N_29934,N_29838);
and UO_2664 (O_2664,N_29925,N_29871);
nor UO_2665 (O_2665,N_29978,N_29929);
xor UO_2666 (O_2666,N_29866,N_29916);
nor UO_2667 (O_2667,N_29838,N_29965);
or UO_2668 (O_2668,N_29873,N_29822);
or UO_2669 (O_2669,N_29941,N_29900);
nor UO_2670 (O_2670,N_29824,N_29852);
xor UO_2671 (O_2671,N_29833,N_29935);
nor UO_2672 (O_2672,N_29981,N_29818);
or UO_2673 (O_2673,N_29986,N_29874);
nand UO_2674 (O_2674,N_29969,N_29818);
and UO_2675 (O_2675,N_29941,N_29957);
and UO_2676 (O_2676,N_29980,N_29842);
nor UO_2677 (O_2677,N_29825,N_29906);
nand UO_2678 (O_2678,N_29863,N_29875);
or UO_2679 (O_2679,N_29980,N_29914);
and UO_2680 (O_2680,N_29815,N_29902);
and UO_2681 (O_2681,N_29859,N_29802);
nor UO_2682 (O_2682,N_29909,N_29878);
and UO_2683 (O_2683,N_29945,N_29883);
xor UO_2684 (O_2684,N_29908,N_29996);
xor UO_2685 (O_2685,N_29911,N_29843);
nand UO_2686 (O_2686,N_29936,N_29898);
and UO_2687 (O_2687,N_29809,N_29970);
nor UO_2688 (O_2688,N_29924,N_29877);
or UO_2689 (O_2689,N_29923,N_29998);
nand UO_2690 (O_2690,N_29870,N_29929);
xor UO_2691 (O_2691,N_29847,N_29837);
xor UO_2692 (O_2692,N_29822,N_29801);
nand UO_2693 (O_2693,N_29929,N_29993);
nand UO_2694 (O_2694,N_29901,N_29909);
or UO_2695 (O_2695,N_29942,N_29870);
or UO_2696 (O_2696,N_29874,N_29966);
xor UO_2697 (O_2697,N_29909,N_29917);
xor UO_2698 (O_2698,N_29852,N_29993);
and UO_2699 (O_2699,N_29874,N_29881);
nand UO_2700 (O_2700,N_29925,N_29815);
and UO_2701 (O_2701,N_29967,N_29810);
nand UO_2702 (O_2702,N_29984,N_29886);
nor UO_2703 (O_2703,N_29885,N_29888);
xnor UO_2704 (O_2704,N_29869,N_29971);
xnor UO_2705 (O_2705,N_29861,N_29813);
and UO_2706 (O_2706,N_29890,N_29835);
and UO_2707 (O_2707,N_29849,N_29966);
and UO_2708 (O_2708,N_29801,N_29930);
xor UO_2709 (O_2709,N_29889,N_29893);
or UO_2710 (O_2710,N_29957,N_29946);
xor UO_2711 (O_2711,N_29856,N_29910);
and UO_2712 (O_2712,N_29990,N_29846);
nand UO_2713 (O_2713,N_29837,N_29975);
nand UO_2714 (O_2714,N_29999,N_29817);
and UO_2715 (O_2715,N_29849,N_29844);
nand UO_2716 (O_2716,N_29896,N_29813);
nor UO_2717 (O_2717,N_29862,N_29800);
nor UO_2718 (O_2718,N_29806,N_29805);
nand UO_2719 (O_2719,N_29880,N_29999);
nand UO_2720 (O_2720,N_29986,N_29995);
nor UO_2721 (O_2721,N_29962,N_29982);
and UO_2722 (O_2722,N_29962,N_29924);
and UO_2723 (O_2723,N_29858,N_29982);
nor UO_2724 (O_2724,N_29938,N_29918);
and UO_2725 (O_2725,N_29956,N_29849);
and UO_2726 (O_2726,N_29839,N_29963);
nor UO_2727 (O_2727,N_29816,N_29823);
nand UO_2728 (O_2728,N_29959,N_29945);
nand UO_2729 (O_2729,N_29919,N_29912);
xnor UO_2730 (O_2730,N_29857,N_29850);
xor UO_2731 (O_2731,N_29828,N_29935);
and UO_2732 (O_2732,N_29978,N_29864);
or UO_2733 (O_2733,N_29933,N_29956);
nand UO_2734 (O_2734,N_29893,N_29967);
nor UO_2735 (O_2735,N_29825,N_29831);
and UO_2736 (O_2736,N_29980,N_29899);
and UO_2737 (O_2737,N_29917,N_29953);
or UO_2738 (O_2738,N_29841,N_29821);
and UO_2739 (O_2739,N_29986,N_29851);
nand UO_2740 (O_2740,N_29868,N_29875);
nand UO_2741 (O_2741,N_29830,N_29852);
or UO_2742 (O_2742,N_29809,N_29982);
nand UO_2743 (O_2743,N_29979,N_29949);
xnor UO_2744 (O_2744,N_29931,N_29941);
or UO_2745 (O_2745,N_29907,N_29939);
or UO_2746 (O_2746,N_29848,N_29925);
nor UO_2747 (O_2747,N_29914,N_29836);
nor UO_2748 (O_2748,N_29950,N_29886);
or UO_2749 (O_2749,N_29912,N_29893);
or UO_2750 (O_2750,N_29949,N_29998);
xor UO_2751 (O_2751,N_29814,N_29949);
and UO_2752 (O_2752,N_29900,N_29996);
nand UO_2753 (O_2753,N_29984,N_29946);
and UO_2754 (O_2754,N_29847,N_29902);
or UO_2755 (O_2755,N_29871,N_29976);
xnor UO_2756 (O_2756,N_29888,N_29882);
or UO_2757 (O_2757,N_29848,N_29930);
or UO_2758 (O_2758,N_29950,N_29804);
nand UO_2759 (O_2759,N_29837,N_29884);
xor UO_2760 (O_2760,N_29922,N_29914);
nand UO_2761 (O_2761,N_29882,N_29950);
nand UO_2762 (O_2762,N_29864,N_29867);
and UO_2763 (O_2763,N_29804,N_29993);
nand UO_2764 (O_2764,N_29954,N_29842);
and UO_2765 (O_2765,N_29865,N_29887);
and UO_2766 (O_2766,N_29973,N_29839);
and UO_2767 (O_2767,N_29852,N_29909);
and UO_2768 (O_2768,N_29976,N_29857);
nand UO_2769 (O_2769,N_29993,N_29808);
or UO_2770 (O_2770,N_29874,N_29983);
nor UO_2771 (O_2771,N_29914,N_29964);
or UO_2772 (O_2772,N_29883,N_29957);
and UO_2773 (O_2773,N_29980,N_29870);
nor UO_2774 (O_2774,N_29827,N_29934);
nor UO_2775 (O_2775,N_29900,N_29898);
and UO_2776 (O_2776,N_29955,N_29903);
xor UO_2777 (O_2777,N_29931,N_29834);
or UO_2778 (O_2778,N_29811,N_29900);
or UO_2779 (O_2779,N_29992,N_29928);
nand UO_2780 (O_2780,N_29835,N_29936);
and UO_2781 (O_2781,N_29933,N_29839);
nor UO_2782 (O_2782,N_29953,N_29815);
nor UO_2783 (O_2783,N_29860,N_29855);
or UO_2784 (O_2784,N_29802,N_29922);
or UO_2785 (O_2785,N_29907,N_29898);
nand UO_2786 (O_2786,N_29900,N_29848);
nor UO_2787 (O_2787,N_29901,N_29844);
nand UO_2788 (O_2788,N_29886,N_29960);
nand UO_2789 (O_2789,N_29974,N_29814);
and UO_2790 (O_2790,N_29912,N_29805);
or UO_2791 (O_2791,N_29823,N_29812);
nand UO_2792 (O_2792,N_29893,N_29905);
nand UO_2793 (O_2793,N_29975,N_29872);
xnor UO_2794 (O_2794,N_29808,N_29857);
nor UO_2795 (O_2795,N_29980,N_29953);
nand UO_2796 (O_2796,N_29817,N_29928);
or UO_2797 (O_2797,N_29803,N_29872);
and UO_2798 (O_2798,N_29838,N_29932);
xnor UO_2799 (O_2799,N_29880,N_29873);
or UO_2800 (O_2800,N_29885,N_29966);
nor UO_2801 (O_2801,N_29898,N_29853);
or UO_2802 (O_2802,N_29925,N_29813);
nand UO_2803 (O_2803,N_29928,N_29838);
and UO_2804 (O_2804,N_29959,N_29874);
nor UO_2805 (O_2805,N_29971,N_29911);
xor UO_2806 (O_2806,N_29861,N_29882);
or UO_2807 (O_2807,N_29811,N_29948);
and UO_2808 (O_2808,N_29810,N_29884);
and UO_2809 (O_2809,N_29990,N_29835);
and UO_2810 (O_2810,N_29807,N_29910);
xor UO_2811 (O_2811,N_29984,N_29996);
nor UO_2812 (O_2812,N_29806,N_29891);
nor UO_2813 (O_2813,N_29826,N_29870);
xor UO_2814 (O_2814,N_29859,N_29959);
xnor UO_2815 (O_2815,N_29811,N_29952);
nor UO_2816 (O_2816,N_29963,N_29915);
nand UO_2817 (O_2817,N_29814,N_29842);
nor UO_2818 (O_2818,N_29891,N_29843);
nand UO_2819 (O_2819,N_29864,N_29836);
and UO_2820 (O_2820,N_29901,N_29820);
xnor UO_2821 (O_2821,N_29936,N_29896);
nor UO_2822 (O_2822,N_29830,N_29867);
xnor UO_2823 (O_2823,N_29896,N_29984);
nand UO_2824 (O_2824,N_29913,N_29865);
xnor UO_2825 (O_2825,N_29990,N_29996);
xnor UO_2826 (O_2826,N_29820,N_29843);
and UO_2827 (O_2827,N_29838,N_29885);
and UO_2828 (O_2828,N_29813,N_29881);
xor UO_2829 (O_2829,N_29841,N_29829);
xnor UO_2830 (O_2830,N_29991,N_29924);
nand UO_2831 (O_2831,N_29992,N_29996);
or UO_2832 (O_2832,N_29884,N_29990);
or UO_2833 (O_2833,N_29859,N_29857);
xor UO_2834 (O_2834,N_29873,N_29940);
nor UO_2835 (O_2835,N_29975,N_29817);
and UO_2836 (O_2836,N_29948,N_29892);
and UO_2837 (O_2837,N_29955,N_29858);
nand UO_2838 (O_2838,N_29828,N_29928);
nand UO_2839 (O_2839,N_29807,N_29990);
or UO_2840 (O_2840,N_29875,N_29858);
nor UO_2841 (O_2841,N_29831,N_29857);
nand UO_2842 (O_2842,N_29825,N_29855);
nor UO_2843 (O_2843,N_29835,N_29886);
nand UO_2844 (O_2844,N_29895,N_29833);
or UO_2845 (O_2845,N_29903,N_29946);
or UO_2846 (O_2846,N_29850,N_29814);
nand UO_2847 (O_2847,N_29912,N_29978);
xnor UO_2848 (O_2848,N_29944,N_29870);
and UO_2849 (O_2849,N_29963,N_29933);
and UO_2850 (O_2850,N_29907,N_29931);
nand UO_2851 (O_2851,N_29921,N_29956);
or UO_2852 (O_2852,N_29996,N_29941);
or UO_2853 (O_2853,N_29901,N_29966);
nor UO_2854 (O_2854,N_29987,N_29821);
or UO_2855 (O_2855,N_29979,N_29859);
and UO_2856 (O_2856,N_29865,N_29900);
xnor UO_2857 (O_2857,N_29926,N_29982);
xnor UO_2858 (O_2858,N_29896,N_29894);
xnor UO_2859 (O_2859,N_29833,N_29901);
and UO_2860 (O_2860,N_29939,N_29834);
xor UO_2861 (O_2861,N_29886,N_29806);
nor UO_2862 (O_2862,N_29851,N_29897);
or UO_2863 (O_2863,N_29930,N_29963);
or UO_2864 (O_2864,N_29845,N_29995);
xnor UO_2865 (O_2865,N_29926,N_29876);
xnor UO_2866 (O_2866,N_29867,N_29961);
or UO_2867 (O_2867,N_29855,N_29817);
xor UO_2868 (O_2868,N_29989,N_29951);
or UO_2869 (O_2869,N_29916,N_29843);
nor UO_2870 (O_2870,N_29887,N_29814);
and UO_2871 (O_2871,N_29878,N_29853);
nand UO_2872 (O_2872,N_29887,N_29884);
xnor UO_2873 (O_2873,N_29902,N_29991);
xor UO_2874 (O_2874,N_29804,N_29836);
nand UO_2875 (O_2875,N_29942,N_29963);
xor UO_2876 (O_2876,N_29924,N_29970);
nand UO_2877 (O_2877,N_29821,N_29819);
nor UO_2878 (O_2878,N_29921,N_29861);
and UO_2879 (O_2879,N_29982,N_29931);
xnor UO_2880 (O_2880,N_29818,N_29964);
or UO_2881 (O_2881,N_29819,N_29886);
or UO_2882 (O_2882,N_29852,N_29814);
nand UO_2883 (O_2883,N_29946,N_29925);
nor UO_2884 (O_2884,N_29967,N_29824);
nand UO_2885 (O_2885,N_29979,N_29868);
and UO_2886 (O_2886,N_29936,N_29964);
and UO_2887 (O_2887,N_29962,N_29990);
nor UO_2888 (O_2888,N_29947,N_29901);
nor UO_2889 (O_2889,N_29815,N_29843);
nor UO_2890 (O_2890,N_29905,N_29940);
nand UO_2891 (O_2891,N_29923,N_29849);
nand UO_2892 (O_2892,N_29989,N_29893);
xor UO_2893 (O_2893,N_29946,N_29890);
nor UO_2894 (O_2894,N_29862,N_29846);
nand UO_2895 (O_2895,N_29854,N_29863);
and UO_2896 (O_2896,N_29874,N_29934);
nand UO_2897 (O_2897,N_29892,N_29956);
nor UO_2898 (O_2898,N_29950,N_29965);
xor UO_2899 (O_2899,N_29942,N_29977);
nand UO_2900 (O_2900,N_29852,N_29821);
or UO_2901 (O_2901,N_29864,N_29879);
xor UO_2902 (O_2902,N_29885,N_29891);
nand UO_2903 (O_2903,N_29932,N_29847);
xnor UO_2904 (O_2904,N_29859,N_29916);
and UO_2905 (O_2905,N_29888,N_29960);
nor UO_2906 (O_2906,N_29827,N_29888);
nor UO_2907 (O_2907,N_29959,N_29935);
nor UO_2908 (O_2908,N_29847,N_29804);
xor UO_2909 (O_2909,N_29957,N_29829);
or UO_2910 (O_2910,N_29955,N_29950);
nand UO_2911 (O_2911,N_29821,N_29876);
and UO_2912 (O_2912,N_29972,N_29970);
and UO_2913 (O_2913,N_29956,N_29836);
xnor UO_2914 (O_2914,N_29986,N_29812);
nand UO_2915 (O_2915,N_29984,N_29930);
xor UO_2916 (O_2916,N_29812,N_29843);
or UO_2917 (O_2917,N_29991,N_29841);
xor UO_2918 (O_2918,N_29911,N_29805);
nand UO_2919 (O_2919,N_29974,N_29917);
and UO_2920 (O_2920,N_29842,N_29833);
xor UO_2921 (O_2921,N_29979,N_29982);
nor UO_2922 (O_2922,N_29832,N_29867);
nor UO_2923 (O_2923,N_29954,N_29987);
or UO_2924 (O_2924,N_29879,N_29878);
and UO_2925 (O_2925,N_29887,N_29856);
nor UO_2926 (O_2926,N_29879,N_29953);
xnor UO_2927 (O_2927,N_29875,N_29877);
and UO_2928 (O_2928,N_29916,N_29985);
xor UO_2929 (O_2929,N_29945,N_29851);
nor UO_2930 (O_2930,N_29993,N_29885);
xor UO_2931 (O_2931,N_29955,N_29811);
xnor UO_2932 (O_2932,N_29822,N_29915);
and UO_2933 (O_2933,N_29809,N_29935);
nor UO_2934 (O_2934,N_29907,N_29888);
nor UO_2935 (O_2935,N_29831,N_29878);
or UO_2936 (O_2936,N_29913,N_29807);
or UO_2937 (O_2937,N_29840,N_29981);
xnor UO_2938 (O_2938,N_29873,N_29821);
or UO_2939 (O_2939,N_29924,N_29888);
nor UO_2940 (O_2940,N_29929,N_29864);
nor UO_2941 (O_2941,N_29987,N_29871);
and UO_2942 (O_2942,N_29897,N_29967);
and UO_2943 (O_2943,N_29886,N_29931);
and UO_2944 (O_2944,N_29999,N_29967);
and UO_2945 (O_2945,N_29874,N_29827);
or UO_2946 (O_2946,N_29913,N_29898);
or UO_2947 (O_2947,N_29800,N_29925);
or UO_2948 (O_2948,N_29841,N_29833);
xor UO_2949 (O_2949,N_29803,N_29867);
and UO_2950 (O_2950,N_29873,N_29834);
or UO_2951 (O_2951,N_29998,N_29866);
and UO_2952 (O_2952,N_29986,N_29929);
nand UO_2953 (O_2953,N_29829,N_29945);
xor UO_2954 (O_2954,N_29856,N_29895);
nand UO_2955 (O_2955,N_29922,N_29882);
or UO_2956 (O_2956,N_29945,N_29907);
and UO_2957 (O_2957,N_29878,N_29854);
nor UO_2958 (O_2958,N_29813,N_29966);
xnor UO_2959 (O_2959,N_29852,N_29976);
nand UO_2960 (O_2960,N_29916,N_29870);
xnor UO_2961 (O_2961,N_29836,N_29807);
nor UO_2962 (O_2962,N_29911,N_29876);
or UO_2963 (O_2963,N_29987,N_29828);
nor UO_2964 (O_2964,N_29833,N_29879);
nand UO_2965 (O_2965,N_29923,N_29929);
nor UO_2966 (O_2966,N_29830,N_29817);
nand UO_2967 (O_2967,N_29979,N_29919);
xnor UO_2968 (O_2968,N_29923,N_29896);
and UO_2969 (O_2969,N_29993,N_29833);
or UO_2970 (O_2970,N_29840,N_29841);
nand UO_2971 (O_2971,N_29918,N_29837);
nor UO_2972 (O_2972,N_29933,N_29898);
nand UO_2973 (O_2973,N_29950,N_29815);
xor UO_2974 (O_2974,N_29975,N_29942);
xor UO_2975 (O_2975,N_29835,N_29967);
nand UO_2976 (O_2976,N_29895,N_29858);
nor UO_2977 (O_2977,N_29944,N_29850);
xor UO_2978 (O_2978,N_29986,N_29994);
nand UO_2979 (O_2979,N_29839,N_29832);
or UO_2980 (O_2980,N_29830,N_29961);
or UO_2981 (O_2981,N_29931,N_29867);
and UO_2982 (O_2982,N_29804,N_29965);
or UO_2983 (O_2983,N_29848,N_29915);
xor UO_2984 (O_2984,N_29872,N_29902);
and UO_2985 (O_2985,N_29814,N_29885);
and UO_2986 (O_2986,N_29993,N_29992);
nand UO_2987 (O_2987,N_29979,N_29841);
xnor UO_2988 (O_2988,N_29848,N_29985);
nor UO_2989 (O_2989,N_29857,N_29937);
and UO_2990 (O_2990,N_29953,N_29936);
nand UO_2991 (O_2991,N_29831,N_29944);
or UO_2992 (O_2992,N_29928,N_29841);
and UO_2993 (O_2993,N_29871,N_29869);
and UO_2994 (O_2994,N_29917,N_29875);
and UO_2995 (O_2995,N_29938,N_29936);
nor UO_2996 (O_2996,N_29933,N_29955);
or UO_2997 (O_2997,N_29819,N_29889);
nor UO_2998 (O_2998,N_29890,N_29844);
nand UO_2999 (O_2999,N_29913,N_29837);
xnor UO_3000 (O_3000,N_29933,N_29927);
or UO_3001 (O_3001,N_29808,N_29991);
or UO_3002 (O_3002,N_29947,N_29996);
nor UO_3003 (O_3003,N_29948,N_29931);
and UO_3004 (O_3004,N_29950,N_29899);
nor UO_3005 (O_3005,N_29877,N_29909);
or UO_3006 (O_3006,N_29975,N_29827);
nand UO_3007 (O_3007,N_29849,N_29856);
or UO_3008 (O_3008,N_29803,N_29881);
nor UO_3009 (O_3009,N_29980,N_29910);
nand UO_3010 (O_3010,N_29805,N_29807);
nand UO_3011 (O_3011,N_29924,N_29994);
or UO_3012 (O_3012,N_29818,N_29917);
or UO_3013 (O_3013,N_29948,N_29934);
xnor UO_3014 (O_3014,N_29941,N_29898);
or UO_3015 (O_3015,N_29859,N_29823);
xor UO_3016 (O_3016,N_29838,N_29868);
and UO_3017 (O_3017,N_29916,N_29856);
nor UO_3018 (O_3018,N_29812,N_29852);
nor UO_3019 (O_3019,N_29886,N_29918);
or UO_3020 (O_3020,N_29979,N_29963);
xnor UO_3021 (O_3021,N_29806,N_29922);
or UO_3022 (O_3022,N_29819,N_29892);
xnor UO_3023 (O_3023,N_29916,N_29969);
nand UO_3024 (O_3024,N_29914,N_29803);
nand UO_3025 (O_3025,N_29870,N_29828);
and UO_3026 (O_3026,N_29934,N_29899);
xor UO_3027 (O_3027,N_29847,N_29912);
nor UO_3028 (O_3028,N_29890,N_29903);
and UO_3029 (O_3029,N_29872,N_29984);
and UO_3030 (O_3030,N_29976,N_29835);
nand UO_3031 (O_3031,N_29845,N_29938);
and UO_3032 (O_3032,N_29803,N_29823);
and UO_3033 (O_3033,N_29841,N_29987);
and UO_3034 (O_3034,N_29905,N_29988);
xor UO_3035 (O_3035,N_29883,N_29870);
nor UO_3036 (O_3036,N_29994,N_29870);
and UO_3037 (O_3037,N_29802,N_29821);
xnor UO_3038 (O_3038,N_29920,N_29921);
or UO_3039 (O_3039,N_29882,N_29940);
xnor UO_3040 (O_3040,N_29837,N_29828);
nand UO_3041 (O_3041,N_29896,N_29807);
nor UO_3042 (O_3042,N_29800,N_29935);
xnor UO_3043 (O_3043,N_29908,N_29812);
xor UO_3044 (O_3044,N_29849,N_29859);
nand UO_3045 (O_3045,N_29992,N_29868);
nand UO_3046 (O_3046,N_29921,N_29924);
or UO_3047 (O_3047,N_29890,N_29821);
xor UO_3048 (O_3048,N_29899,N_29904);
or UO_3049 (O_3049,N_29821,N_29975);
and UO_3050 (O_3050,N_29957,N_29984);
nor UO_3051 (O_3051,N_29989,N_29993);
nor UO_3052 (O_3052,N_29814,N_29957);
nand UO_3053 (O_3053,N_29978,N_29849);
nand UO_3054 (O_3054,N_29882,N_29900);
xor UO_3055 (O_3055,N_29935,N_29838);
nand UO_3056 (O_3056,N_29900,N_29918);
nand UO_3057 (O_3057,N_29895,N_29944);
or UO_3058 (O_3058,N_29852,N_29902);
nor UO_3059 (O_3059,N_29979,N_29996);
nand UO_3060 (O_3060,N_29966,N_29976);
or UO_3061 (O_3061,N_29909,N_29894);
and UO_3062 (O_3062,N_29924,N_29967);
and UO_3063 (O_3063,N_29833,N_29821);
nand UO_3064 (O_3064,N_29879,N_29875);
xor UO_3065 (O_3065,N_29903,N_29942);
nor UO_3066 (O_3066,N_29809,N_29876);
and UO_3067 (O_3067,N_29993,N_29921);
and UO_3068 (O_3068,N_29973,N_29964);
and UO_3069 (O_3069,N_29840,N_29878);
nand UO_3070 (O_3070,N_29925,N_29863);
or UO_3071 (O_3071,N_29865,N_29917);
xor UO_3072 (O_3072,N_29991,N_29913);
and UO_3073 (O_3073,N_29932,N_29992);
xnor UO_3074 (O_3074,N_29807,N_29851);
nand UO_3075 (O_3075,N_29984,N_29876);
xnor UO_3076 (O_3076,N_29806,N_29938);
nor UO_3077 (O_3077,N_29825,N_29884);
or UO_3078 (O_3078,N_29936,N_29819);
or UO_3079 (O_3079,N_29845,N_29971);
or UO_3080 (O_3080,N_29974,N_29921);
xnor UO_3081 (O_3081,N_29958,N_29945);
nor UO_3082 (O_3082,N_29939,N_29829);
xor UO_3083 (O_3083,N_29811,N_29879);
and UO_3084 (O_3084,N_29982,N_29886);
nand UO_3085 (O_3085,N_29928,N_29825);
nor UO_3086 (O_3086,N_29900,N_29944);
xor UO_3087 (O_3087,N_29892,N_29897);
nand UO_3088 (O_3088,N_29963,N_29993);
nand UO_3089 (O_3089,N_29964,N_29951);
and UO_3090 (O_3090,N_29991,N_29954);
xor UO_3091 (O_3091,N_29832,N_29852);
nand UO_3092 (O_3092,N_29808,N_29969);
or UO_3093 (O_3093,N_29935,N_29856);
xor UO_3094 (O_3094,N_29895,N_29953);
xor UO_3095 (O_3095,N_29867,N_29833);
nor UO_3096 (O_3096,N_29933,N_29934);
or UO_3097 (O_3097,N_29839,N_29966);
nor UO_3098 (O_3098,N_29918,N_29989);
nor UO_3099 (O_3099,N_29828,N_29976);
or UO_3100 (O_3100,N_29880,N_29879);
nor UO_3101 (O_3101,N_29916,N_29989);
nor UO_3102 (O_3102,N_29989,N_29865);
and UO_3103 (O_3103,N_29943,N_29824);
or UO_3104 (O_3104,N_29896,N_29802);
and UO_3105 (O_3105,N_29969,N_29991);
xnor UO_3106 (O_3106,N_29839,N_29840);
xnor UO_3107 (O_3107,N_29989,N_29969);
xor UO_3108 (O_3108,N_29879,N_29969);
and UO_3109 (O_3109,N_29817,N_29846);
xnor UO_3110 (O_3110,N_29827,N_29840);
nand UO_3111 (O_3111,N_29997,N_29962);
nand UO_3112 (O_3112,N_29961,N_29950);
nand UO_3113 (O_3113,N_29942,N_29918);
or UO_3114 (O_3114,N_29877,N_29891);
nor UO_3115 (O_3115,N_29866,N_29907);
or UO_3116 (O_3116,N_29956,N_29930);
nand UO_3117 (O_3117,N_29828,N_29824);
and UO_3118 (O_3118,N_29962,N_29834);
nor UO_3119 (O_3119,N_29928,N_29980);
nand UO_3120 (O_3120,N_29870,N_29886);
or UO_3121 (O_3121,N_29861,N_29994);
and UO_3122 (O_3122,N_29874,N_29887);
nand UO_3123 (O_3123,N_29812,N_29819);
nor UO_3124 (O_3124,N_29966,N_29983);
nand UO_3125 (O_3125,N_29840,N_29876);
nor UO_3126 (O_3126,N_29952,N_29814);
or UO_3127 (O_3127,N_29951,N_29822);
and UO_3128 (O_3128,N_29939,N_29982);
xor UO_3129 (O_3129,N_29847,N_29988);
or UO_3130 (O_3130,N_29999,N_29963);
nand UO_3131 (O_3131,N_29844,N_29862);
xor UO_3132 (O_3132,N_29860,N_29891);
nand UO_3133 (O_3133,N_29962,N_29903);
or UO_3134 (O_3134,N_29884,N_29956);
and UO_3135 (O_3135,N_29832,N_29844);
nand UO_3136 (O_3136,N_29932,N_29807);
and UO_3137 (O_3137,N_29833,N_29921);
nand UO_3138 (O_3138,N_29935,N_29967);
xor UO_3139 (O_3139,N_29900,N_29938);
xnor UO_3140 (O_3140,N_29922,N_29887);
nand UO_3141 (O_3141,N_29992,N_29962);
or UO_3142 (O_3142,N_29811,N_29977);
xor UO_3143 (O_3143,N_29849,N_29854);
nand UO_3144 (O_3144,N_29878,N_29910);
and UO_3145 (O_3145,N_29844,N_29821);
nor UO_3146 (O_3146,N_29904,N_29822);
and UO_3147 (O_3147,N_29919,N_29855);
nor UO_3148 (O_3148,N_29825,N_29953);
and UO_3149 (O_3149,N_29859,N_29884);
nand UO_3150 (O_3150,N_29901,N_29823);
nand UO_3151 (O_3151,N_29841,N_29800);
nor UO_3152 (O_3152,N_29845,N_29956);
xnor UO_3153 (O_3153,N_29866,N_29939);
or UO_3154 (O_3154,N_29800,N_29845);
xor UO_3155 (O_3155,N_29974,N_29891);
or UO_3156 (O_3156,N_29878,N_29889);
xor UO_3157 (O_3157,N_29812,N_29869);
or UO_3158 (O_3158,N_29878,N_29870);
nand UO_3159 (O_3159,N_29906,N_29863);
nand UO_3160 (O_3160,N_29868,N_29922);
and UO_3161 (O_3161,N_29843,N_29872);
nor UO_3162 (O_3162,N_29867,N_29849);
nor UO_3163 (O_3163,N_29881,N_29942);
and UO_3164 (O_3164,N_29810,N_29992);
xnor UO_3165 (O_3165,N_29912,N_29830);
nor UO_3166 (O_3166,N_29899,N_29847);
and UO_3167 (O_3167,N_29920,N_29803);
xnor UO_3168 (O_3168,N_29918,N_29840);
nand UO_3169 (O_3169,N_29983,N_29999);
nand UO_3170 (O_3170,N_29917,N_29939);
and UO_3171 (O_3171,N_29923,N_29856);
nor UO_3172 (O_3172,N_29963,N_29910);
xnor UO_3173 (O_3173,N_29819,N_29937);
xnor UO_3174 (O_3174,N_29813,N_29853);
xor UO_3175 (O_3175,N_29982,N_29897);
nor UO_3176 (O_3176,N_29987,N_29801);
or UO_3177 (O_3177,N_29948,N_29890);
nor UO_3178 (O_3178,N_29983,N_29825);
xor UO_3179 (O_3179,N_29844,N_29977);
xor UO_3180 (O_3180,N_29956,N_29972);
and UO_3181 (O_3181,N_29949,N_29812);
or UO_3182 (O_3182,N_29939,N_29846);
xnor UO_3183 (O_3183,N_29956,N_29851);
nor UO_3184 (O_3184,N_29986,N_29912);
nand UO_3185 (O_3185,N_29860,N_29929);
and UO_3186 (O_3186,N_29857,N_29874);
nor UO_3187 (O_3187,N_29998,N_29978);
xnor UO_3188 (O_3188,N_29982,N_29991);
xor UO_3189 (O_3189,N_29980,N_29951);
nor UO_3190 (O_3190,N_29809,N_29821);
nand UO_3191 (O_3191,N_29952,N_29998);
xor UO_3192 (O_3192,N_29969,N_29966);
nor UO_3193 (O_3193,N_29809,N_29983);
nand UO_3194 (O_3194,N_29980,N_29801);
nor UO_3195 (O_3195,N_29863,N_29928);
xnor UO_3196 (O_3196,N_29964,N_29932);
xor UO_3197 (O_3197,N_29813,N_29936);
xnor UO_3198 (O_3198,N_29984,N_29965);
nand UO_3199 (O_3199,N_29859,N_29908);
nand UO_3200 (O_3200,N_29946,N_29989);
or UO_3201 (O_3201,N_29942,N_29938);
nor UO_3202 (O_3202,N_29985,N_29826);
or UO_3203 (O_3203,N_29830,N_29860);
nand UO_3204 (O_3204,N_29891,N_29973);
xnor UO_3205 (O_3205,N_29861,N_29966);
nor UO_3206 (O_3206,N_29819,N_29869);
nor UO_3207 (O_3207,N_29911,N_29994);
and UO_3208 (O_3208,N_29923,N_29897);
or UO_3209 (O_3209,N_29949,N_29864);
and UO_3210 (O_3210,N_29974,N_29957);
nor UO_3211 (O_3211,N_29983,N_29948);
nor UO_3212 (O_3212,N_29923,N_29987);
xnor UO_3213 (O_3213,N_29806,N_29964);
xnor UO_3214 (O_3214,N_29932,N_29948);
xnor UO_3215 (O_3215,N_29810,N_29806);
nand UO_3216 (O_3216,N_29824,N_29975);
nor UO_3217 (O_3217,N_29820,N_29916);
and UO_3218 (O_3218,N_29831,N_29958);
and UO_3219 (O_3219,N_29928,N_29914);
or UO_3220 (O_3220,N_29860,N_29903);
nor UO_3221 (O_3221,N_29857,N_29801);
and UO_3222 (O_3222,N_29975,N_29873);
and UO_3223 (O_3223,N_29880,N_29972);
xor UO_3224 (O_3224,N_29882,N_29998);
or UO_3225 (O_3225,N_29913,N_29827);
and UO_3226 (O_3226,N_29917,N_29977);
and UO_3227 (O_3227,N_29833,N_29888);
nand UO_3228 (O_3228,N_29806,N_29991);
nand UO_3229 (O_3229,N_29866,N_29967);
nand UO_3230 (O_3230,N_29892,N_29815);
and UO_3231 (O_3231,N_29948,N_29807);
or UO_3232 (O_3232,N_29900,N_29972);
or UO_3233 (O_3233,N_29816,N_29959);
nand UO_3234 (O_3234,N_29966,N_29957);
nor UO_3235 (O_3235,N_29877,N_29921);
or UO_3236 (O_3236,N_29828,N_29965);
xnor UO_3237 (O_3237,N_29872,N_29926);
or UO_3238 (O_3238,N_29926,N_29947);
or UO_3239 (O_3239,N_29938,N_29947);
xor UO_3240 (O_3240,N_29987,N_29948);
nor UO_3241 (O_3241,N_29892,N_29964);
or UO_3242 (O_3242,N_29844,N_29911);
nor UO_3243 (O_3243,N_29976,N_29830);
nand UO_3244 (O_3244,N_29843,N_29999);
nor UO_3245 (O_3245,N_29964,N_29877);
nor UO_3246 (O_3246,N_29940,N_29814);
nor UO_3247 (O_3247,N_29933,N_29964);
or UO_3248 (O_3248,N_29940,N_29846);
and UO_3249 (O_3249,N_29880,N_29875);
nand UO_3250 (O_3250,N_29980,N_29893);
nor UO_3251 (O_3251,N_29867,N_29813);
nor UO_3252 (O_3252,N_29814,N_29835);
nand UO_3253 (O_3253,N_29910,N_29840);
xnor UO_3254 (O_3254,N_29971,N_29983);
and UO_3255 (O_3255,N_29998,N_29932);
nand UO_3256 (O_3256,N_29879,N_29938);
nand UO_3257 (O_3257,N_29867,N_29865);
or UO_3258 (O_3258,N_29803,N_29885);
or UO_3259 (O_3259,N_29888,N_29928);
and UO_3260 (O_3260,N_29860,N_29879);
nand UO_3261 (O_3261,N_29803,N_29971);
or UO_3262 (O_3262,N_29913,N_29874);
or UO_3263 (O_3263,N_29947,N_29986);
xnor UO_3264 (O_3264,N_29851,N_29894);
or UO_3265 (O_3265,N_29990,N_29833);
or UO_3266 (O_3266,N_29817,N_29832);
nor UO_3267 (O_3267,N_29911,N_29997);
or UO_3268 (O_3268,N_29855,N_29990);
nor UO_3269 (O_3269,N_29892,N_29834);
or UO_3270 (O_3270,N_29930,N_29962);
nor UO_3271 (O_3271,N_29862,N_29927);
xor UO_3272 (O_3272,N_29865,N_29868);
xnor UO_3273 (O_3273,N_29842,N_29875);
nand UO_3274 (O_3274,N_29811,N_29983);
nor UO_3275 (O_3275,N_29987,N_29959);
nand UO_3276 (O_3276,N_29963,N_29941);
nand UO_3277 (O_3277,N_29939,N_29840);
and UO_3278 (O_3278,N_29847,N_29992);
or UO_3279 (O_3279,N_29855,N_29915);
and UO_3280 (O_3280,N_29889,N_29915);
nand UO_3281 (O_3281,N_29952,N_29877);
or UO_3282 (O_3282,N_29898,N_29810);
xor UO_3283 (O_3283,N_29904,N_29887);
xnor UO_3284 (O_3284,N_29807,N_29863);
xnor UO_3285 (O_3285,N_29821,N_29804);
xnor UO_3286 (O_3286,N_29884,N_29950);
nor UO_3287 (O_3287,N_29986,N_29955);
and UO_3288 (O_3288,N_29928,N_29986);
or UO_3289 (O_3289,N_29945,N_29824);
nand UO_3290 (O_3290,N_29862,N_29979);
nor UO_3291 (O_3291,N_29875,N_29984);
nor UO_3292 (O_3292,N_29862,N_29968);
xor UO_3293 (O_3293,N_29884,N_29803);
nand UO_3294 (O_3294,N_29891,N_29872);
xnor UO_3295 (O_3295,N_29842,N_29894);
xnor UO_3296 (O_3296,N_29891,N_29908);
nor UO_3297 (O_3297,N_29934,N_29904);
or UO_3298 (O_3298,N_29827,N_29946);
nor UO_3299 (O_3299,N_29882,N_29967);
nand UO_3300 (O_3300,N_29985,N_29975);
nor UO_3301 (O_3301,N_29976,N_29842);
nand UO_3302 (O_3302,N_29820,N_29918);
nand UO_3303 (O_3303,N_29902,N_29918);
and UO_3304 (O_3304,N_29925,N_29901);
nor UO_3305 (O_3305,N_29969,N_29886);
xor UO_3306 (O_3306,N_29989,N_29861);
nand UO_3307 (O_3307,N_29803,N_29938);
xor UO_3308 (O_3308,N_29968,N_29963);
and UO_3309 (O_3309,N_29979,N_29864);
and UO_3310 (O_3310,N_29849,N_29865);
and UO_3311 (O_3311,N_29948,N_29818);
xor UO_3312 (O_3312,N_29853,N_29886);
xnor UO_3313 (O_3313,N_29818,N_29829);
xor UO_3314 (O_3314,N_29901,N_29988);
xnor UO_3315 (O_3315,N_29820,N_29878);
or UO_3316 (O_3316,N_29856,N_29978);
and UO_3317 (O_3317,N_29910,N_29949);
and UO_3318 (O_3318,N_29994,N_29985);
xor UO_3319 (O_3319,N_29805,N_29898);
nor UO_3320 (O_3320,N_29954,N_29848);
xnor UO_3321 (O_3321,N_29878,N_29899);
nor UO_3322 (O_3322,N_29803,N_29977);
or UO_3323 (O_3323,N_29980,N_29883);
nor UO_3324 (O_3324,N_29887,N_29958);
nand UO_3325 (O_3325,N_29825,N_29881);
xor UO_3326 (O_3326,N_29809,N_29923);
and UO_3327 (O_3327,N_29848,N_29919);
or UO_3328 (O_3328,N_29930,N_29833);
nor UO_3329 (O_3329,N_29937,N_29987);
nor UO_3330 (O_3330,N_29819,N_29826);
or UO_3331 (O_3331,N_29813,N_29973);
and UO_3332 (O_3332,N_29951,N_29839);
or UO_3333 (O_3333,N_29887,N_29966);
nor UO_3334 (O_3334,N_29821,N_29950);
nand UO_3335 (O_3335,N_29946,N_29844);
nand UO_3336 (O_3336,N_29977,N_29929);
xor UO_3337 (O_3337,N_29936,N_29856);
and UO_3338 (O_3338,N_29910,N_29847);
xor UO_3339 (O_3339,N_29959,N_29892);
nand UO_3340 (O_3340,N_29824,N_29959);
or UO_3341 (O_3341,N_29851,N_29863);
xor UO_3342 (O_3342,N_29972,N_29964);
or UO_3343 (O_3343,N_29925,N_29920);
and UO_3344 (O_3344,N_29975,N_29835);
xnor UO_3345 (O_3345,N_29837,N_29821);
and UO_3346 (O_3346,N_29898,N_29973);
xor UO_3347 (O_3347,N_29803,N_29958);
nand UO_3348 (O_3348,N_29900,N_29845);
and UO_3349 (O_3349,N_29994,N_29865);
or UO_3350 (O_3350,N_29898,N_29820);
and UO_3351 (O_3351,N_29870,N_29972);
nor UO_3352 (O_3352,N_29848,N_29972);
xor UO_3353 (O_3353,N_29881,N_29887);
nand UO_3354 (O_3354,N_29910,N_29968);
or UO_3355 (O_3355,N_29837,N_29889);
nand UO_3356 (O_3356,N_29959,N_29984);
nand UO_3357 (O_3357,N_29891,N_29882);
xnor UO_3358 (O_3358,N_29898,N_29856);
or UO_3359 (O_3359,N_29896,N_29978);
nor UO_3360 (O_3360,N_29963,N_29937);
xor UO_3361 (O_3361,N_29908,N_29983);
xnor UO_3362 (O_3362,N_29929,N_29831);
xnor UO_3363 (O_3363,N_29857,N_29852);
or UO_3364 (O_3364,N_29863,N_29901);
or UO_3365 (O_3365,N_29874,N_29954);
nand UO_3366 (O_3366,N_29873,N_29993);
nand UO_3367 (O_3367,N_29807,N_29872);
or UO_3368 (O_3368,N_29922,N_29884);
nand UO_3369 (O_3369,N_29910,N_29997);
xor UO_3370 (O_3370,N_29868,N_29890);
or UO_3371 (O_3371,N_29908,N_29977);
xnor UO_3372 (O_3372,N_29819,N_29942);
and UO_3373 (O_3373,N_29995,N_29904);
nor UO_3374 (O_3374,N_29870,N_29973);
and UO_3375 (O_3375,N_29912,N_29976);
xnor UO_3376 (O_3376,N_29892,N_29873);
and UO_3377 (O_3377,N_29827,N_29893);
xor UO_3378 (O_3378,N_29894,N_29833);
nor UO_3379 (O_3379,N_29882,N_29890);
xnor UO_3380 (O_3380,N_29953,N_29884);
and UO_3381 (O_3381,N_29958,N_29985);
nand UO_3382 (O_3382,N_29985,N_29986);
xnor UO_3383 (O_3383,N_29906,N_29922);
or UO_3384 (O_3384,N_29950,N_29974);
nor UO_3385 (O_3385,N_29817,N_29800);
xnor UO_3386 (O_3386,N_29957,N_29976);
nor UO_3387 (O_3387,N_29945,N_29848);
nor UO_3388 (O_3388,N_29991,N_29880);
nand UO_3389 (O_3389,N_29839,N_29923);
nand UO_3390 (O_3390,N_29927,N_29939);
and UO_3391 (O_3391,N_29850,N_29909);
xnor UO_3392 (O_3392,N_29865,N_29980);
or UO_3393 (O_3393,N_29813,N_29898);
xnor UO_3394 (O_3394,N_29944,N_29820);
and UO_3395 (O_3395,N_29998,N_29950);
and UO_3396 (O_3396,N_29979,N_29824);
and UO_3397 (O_3397,N_29931,N_29981);
nand UO_3398 (O_3398,N_29966,N_29986);
xor UO_3399 (O_3399,N_29807,N_29934);
nor UO_3400 (O_3400,N_29868,N_29962);
nor UO_3401 (O_3401,N_29884,N_29912);
xnor UO_3402 (O_3402,N_29899,N_29987);
nand UO_3403 (O_3403,N_29928,N_29903);
or UO_3404 (O_3404,N_29905,N_29931);
or UO_3405 (O_3405,N_29887,N_29916);
nor UO_3406 (O_3406,N_29972,N_29889);
nor UO_3407 (O_3407,N_29971,N_29949);
xor UO_3408 (O_3408,N_29986,N_29834);
xor UO_3409 (O_3409,N_29951,N_29911);
nand UO_3410 (O_3410,N_29924,N_29956);
xnor UO_3411 (O_3411,N_29815,N_29880);
xor UO_3412 (O_3412,N_29860,N_29841);
xor UO_3413 (O_3413,N_29908,N_29888);
xor UO_3414 (O_3414,N_29903,N_29876);
nand UO_3415 (O_3415,N_29815,N_29909);
or UO_3416 (O_3416,N_29964,N_29885);
xnor UO_3417 (O_3417,N_29949,N_29809);
xor UO_3418 (O_3418,N_29863,N_29975);
or UO_3419 (O_3419,N_29889,N_29880);
and UO_3420 (O_3420,N_29884,N_29896);
or UO_3421 (O_3421,N_29887,N_29981);
nand UO_3422 (O_3422,N_29845,N_29952);
and UO_3423 (O_3423,N_29868,N_29984);
nor UO_3424 (O_3424,N_29877,N_29931);
nor UO_3425 (O_3425,N_29895,N_29894);
nor UO_3426 (O_3426,N_29822,N_29994);
or UO_3427 (O_3427,N_29860,N_29957);
and UO_3428 (O_3428,N_29926,N_29819);
nor UO_3429 (O_3429,N_29870,N_29899);
and UO_3430 (O_3430,N_29866,N_29934);
or UO_3431 (O_3431,N_29890,N_29997);
or UO_3432 (O_3432,N_29996,N_29877);
nor UO_3433 (O_3433,N_29817,N_29802);
xor UO_3434 (O_3434,N_29823,N_29904);
xor UO_3435 (O_3435,N_29880,N_29992);
nor UO_3436 (O_3436,N_29924,N_29806);
or UO_3437 (O_3437,N_29880,N_29949);
and UO_3438 (O_3438,N_29839,N_29856);
nand UO_3439 (O_3439,N_29865,N_29974);
nor UO_3440 (O_3440,N_29847,N_29856);
nor UO_3441 (O_3441,N_29835,N_29968);
nand UO_3442 (O_3442,N_29854,N_29938);
nand UO_3443 (O_3443,N_29803,N_29972);
or UO_3444 (O_3444,N_29937,N_29926);
or UO_3445 (O_3445,N_29914,N_29970);
or UO_3446 (O_3446,N_29985,N_29800);
xnor UO_3447 (O_3447,N_29928,N_29896);
nor UO_3448 (O_3448,N_29857,N_29954);
nand UO_3449 (O_3449,N_29821,N_29970);
nand UO_3450 (O_3450,N_29823,N_29868);
or UO_3451 (O_3451,N_29942,N_29883);
nand UO_3452 (O_3452,N_29890,N_29964);
xor UO_3453 (O_3453,N_29885,N_29807);
or UO_3454 (O_3454,N_29878,N_29935);
and UO_3455 (O_3455,N_29938,N_29817);
xnor UO_3456 (O_3456,N_29901,N_29803);
nor UO_3457 (O_3457,N_29913,N_29826);
xor UO_3458 (O_3458,N_29853,N_29962);
or UO_3459 (O_3459,N_29936,N_29966);
nor UO_3460 (O_3460,N_29857,N_29978);
nand UO_3461 (O_3461,N_29977,N_29997);
nor UO_3462 (O_3462,N_29960,N_29904);
xor UO_3463 (O_3463,N_29923,N_29980);
nor UO_3464 (O_3464,N_29980,N_29828);
nand UO_3465 (O_3465,N_29879,N_29945);
nand UO_3466 (O_3466,N_29801,N_29870);
and UO_3467 (O_3467,N_29834,N_29880);
nor UO_3468 (O_3468,N_29875,N_29946);
nand UO_3469 (O_3469,N_29842,N_29979);
or UO_3470 (O_3470,N_29840,N_29979);
xor UO_3471 (O_3471,N_29941,N_29868);
and UO_3472 (O_3472,N_29936,N_29815);
and UO_3473 (O_3473,N_29811,N_29993);
or UO_3474 (O_3474,N_29945,N_29814);
nor UO_3475 (O_3475,N_29967,N_29965);
xnor UO_3476 (O_3476,N_29941,N_29812);
or UO_3477 (O_3477,N_29874,N_29837);
xnor UO_3478 (O_3478,N_29813,N_29910);
or UO_3479 (O_3479,N_29887,N_29956);
or UO_3480 (O_3480,N_29882,N_29906);
or UO_3481 (O_3481,N_29828,N_29807);
nor UO_3482 (O_3482,N_29952,N_29954);
and UO_3483 (O_3483,N_29883,N_29999);
nand UO_3484 (O_3484,N_29880,N_29912);
nand UO_3485 (O_3485,N_29934,N_29858);
or UO_3486 (O_3486,N_29877,N_29848);
nor UO_3487 (O_3487,N_29993,N_29827);
or UO_3488 (O_3488,N_29952,N_29888);
nand UO_3489 (O_3489,N_29863,N_29974);
and UO_3490 (O_3490,N_29852,N_29841);
and UO_3491 (O_3491,N_29936,N_29917);
nor UO_3492 (O_3492,N_29952,N_29827);
and UO_3493 (O_3493,N_29835,N_29923);
and UO_3494 (O_3494,N_29891,N_29857);
xor UO_3495 (O_3495,N_29930,N_29971);
and UO_3496 (O_3496,N_29849,N_29872);
xnor UO_3497 (O_3497,N_29959,N_29904);
or UO_3498 (O_3498,N_29993,N_29918);
and UO_3499 (O_3499,N_29967,N_29943);
endmodule