module basic_500_3000_500_60_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_433,In_61);
nor U1 (N_1,In_20,In_89);
nor U2 (N_2,In_470,In_267);
nand U3 (N_3,In_312,In_357);
nor U4 (N_4,In_60,In_485);
nor U5 (N_5,In_283,In_145);
nand U6 (N_6,In_184,In_420);
or U7 (N_7,In_275,In_362);
xnor U8 (N_8,In_278,In_74);
nor U9 (N_9,In_187,In_28);
and U10 (N_10,In_301,In_150);
or U11 (N_11,In_345,In_498);
nor U12 (N_12,In_288,In_271);
nor U13 (N_13,In_156,In_442);
xor U14 (N_14,In_26,In_298);
xnor U15 (N_15,In_192,In_22);
xnor U16 (N_16,In_475,In_306);
xnor U17 (N_17,In_354,In_372);
and U18 (N_18,In_255,In_396);
xnor U19 (N_19,In_1,In_101);
nand U20 (N_20,In_347,In_139);
and U21 (N_21,In_33,In_34);
nor U22 (N_22,In_118,In_166);
and U23 (N_23,In_438,In_422);
xnor U24 (N_24,In_45,In_141);
and U25 (N_25,In_258,In_41);
or U26 (N_26,In_398,In_457);
nand U27 (N_27,In_127,In_331);
or U28 (N_28,In_387,In_488);
xor U29 (N_29,In_296,In_450);
nor U30 (N_30,In_463,In_379);
nor U31 (N_31,In_399,In_176);
or U32 (N_32,In_106,In_79);
nor U33 (N_33,In_429,In_226);
xor U34 (N_34,In_124,In_229);
nand U35 (N_35,In_400,In_234);
nand U36 (N_36,In_369,In_427);
xor U37 (N_37,In_410,In_448);
or U38 (N_38,In_201,In_227);
nor U39 (N_39,In_460,In_388);
and U40 (N_40,In_297,In_143);
or U41 (N_41,In_277,In_204);
xor U42 (N_42,In_374,In_92);
nand U43 (N_43,In_295,In_479);
nand U44 (N_44,In_65,In_445);
or U45 (N_45,In_196,In_38);
xor U46 (N_46,In_392,In_373);
nand U47 (N_47,In_224,In_161);
nand U48 (N_48,In_254,In_253);
xnor U49 (N_49,In_160,In_85);
xor U50 (N_50,In_18,In_363);
nor U51 (N_51,In_42,In_66);
nand U52 (N_52,In_134,In_282);
or U53 (N_53,In_167,In_169);
or U54 (N_54,In_165,In_402);
and U55 (N_55,In_123,In_37);
nor U56 (N_56,In_129,In_366);
nor U57 (N_57,In_29,In_495);
nand U58 (N_58,In_483,In_71);
xor U59 (N_59,In_337,In_452);
or U60 (N_60,In_413,In_342);
or U61 (N_61,In_261,In_385);
or U62 (N_62,In_19,In_352);
or U63 (N_63,In_191,In_408);
nor U64 (N_64,In_246,In_95);
and U65 (N_65,In_451,In_406);
and U66 (N_66,In_480,In_177);
xor U67 (N_67,In_25,In_5);
or U68 (N_68,In_104,N_19);
or U69 (N_69,In_232,In_286);
nor U70 (N_70,N_11,In_497);
nand U71 (N_71,In_222,In_235);
or U72 (N_72,In_98,In_76);
xor U73 (N_73,In_87,In_437);
nor U74 (N_74,In_21,In_17);
or U75 (N_75,In_12,In_307);
nand U76 (N_76,In_305,In_395);
or U77 (N_77,N_31,In_308);
and U78 (N_78,In_97,In_158);
nor U79 (N_79,In_208,In_237);
xor U80 (N_80,In_52,In_455);
nand U81 (N_81,In_325,In_233);
and U82 (N_82,In_202,In_404);
or U83 (N_83,In_188,In_30);
nor U84 (N_84,In_172,In_310);
and U85 (N_85,In_424,In_471);
nor U86 (N_86,In_211,N_20);
xnor U87 (N_87,In_23,N_0);
and U88 (N_88,In_39,In_209);
or U89 (N_89,In_54,In_14);
xor U90 (N_90,In_40,In_371);
nand U91 (N_91,In_327,N_46);
nor U92 (N_92,In_287,In_454);
nand U93 (N_93,In_317,In_130);
or U94 (N_94,In_225,In_193);
nor U95 (N_95,In_320,In_4);
nor U96 (N_96,N_43,In_238);
xor U97 (N_97,In_491,In_185);
nand U98 (N_98,In_493,In_403);
and U99 (N_99,In_351,N_7);
or U100 (N_100,In_249,In_272);
or U101 (N_101,In_121,In_142);
xor U102 (N_102,In_153,In_439);
nor U103 (N_103,In_333,N_63);
and U104 (N_104,In_370,In_252);
nand U105 (N_105,N_51,In_266);
nor U106 (N_106,In_302,N_33);
xnor U107 (N_107,In_175,In_6);
nand U108 (N_108,In_205,In_280);
nand U109 (N_109,In_279,In_384);
or U110 (N_110,In_242,In_416);
nor U111 (N_111,In_414,N_86);
xnor U112 (N_112,In_195,In_447);
xor U113 (N_113,In_263,N_23);
nand U114 (N_114,In_199,In_55);
nand U115 (N_115,In_376,In_340);
nor U116 (N_116,In_334,In_31);
and U117 (N_117,In_350,N_88);
or U118 (N_118,In_113,In_268);
nand U119 (N_119,In_46,In_149);
nand U120 (N_120,In_368,In_7);
nand U121 (N_121,In_323,In_215);
nor U122 (N_122,In_247,N_1);
or U123 (N_123,In_217,In_173);
nor U124 (N_124,In_183,N_27);
xor U125 (N_125,N_72,In_294);
or U126 (N_126,N_59,In_122);
nor U127 (N_127,In_428,In_443);
nor U128 (N_128,In_499,In_221);
xor U129 (N_129,In_43,In_421);
nor U130 (N_130,In_117,In_140);
nor U131 (N_131,In_8,In_494);
and U132 (N_132,In_311,N_29);
xor U133 (N_133,In_180,In_231);
nand U134 (N_134,In_162,In_259);
nor U135 (N_135,In_83,In_353);
nand U136 (N_136,N_74,In_423);
nor U137 (N_137,In_315,In_84);
nor U138 (N_138,In_289,In_174);
nor U139 (N_139,In_344,In_382);
and U140 (N_140,In_212,In_412);
nor U141 (N_141,In_484,In_240);
and U142 (N_142,In_159,In_446);
nor U143 (N_143,In_250,In_461);
xnor U144 (N_144,In_314,In_481);
and U145 (N_145,In_62,In_88);
and U146 (N_146,In_330,In_133);
or U147 (N_147,In_322,In_67);
nand U148 (N_148,In_380,N_4);
xor U149 (N_149,N_54,In_91);
xnor U150 (N_150,N_87,In_207);
xor U151 (N_151,In_418,In_332);
and U152 (N_152,N_144,In_291);
xor U153 (N_153,In_273,N_137);
nor U154 (N_154,N_123,In_440);
or U155 (N_155,In_151,In_270);
nand U156 (N_156,In_94,In_15);
nor U157 (N_157,N_79,N_121);
and U158 (N_158,In_397,In_147);
nor U159 (N_159,N_119,In_16);
xnor U160 (N_160,In_329,In_346);
or U161 (N_161,In_339,In_256);
nor U162 (N_162,In_190,N_77);
or U163 (N_163,In_276,N_149);
xor U164 (N_164,N_84,In_119);
and U165 (N_165,In_103,In_482);
and U166 (N_166,N_115,In_72);
nand U167 (N_167,In_115,In_319);
xnor U168 (N_168,N_132,N_65);
or U169 (N_169,In_462,In_415);
nand U170 (N_170,N_129,In_241);
xnor U171 (N_171,In_401,N_140);
nor U172 (N_172,In_220,N_21);
nor U173 (N_173,In_148,In_300);
or U174 (N_174,In_49,In_472);
nor U175 (N_175,N_142,N_101);
and U176 (N_176,In_383,In_274);
and U177 (N_177,In_114,In_431);
xnor U178 (N_178,In_367,In_3);
or U179 (N_179,N_85,N_66);
or U180 (N_180,In_186,In_108);
or U181 (N_181,N_112,In_244);
and U182 (N_182,In_248,In_131);
and U183 (N_183,N_39,In_228);
xor U184 (N_184,In_27,N_69);
or U185 (N_185,N_56,In_377);
nand U186 (N_186,N_98,N_143);
or U187 (N_187,In_394,N_130);
nor U188 (N_188,In_170,In_63);
and U189 (N_189,N_95,In_343);
nor U190 (N_190,In_100,In_390);
nor U191 (N_191,In_435,N_17);
xnor U192 (N_192,N_92,In_181);
nand U193 (N_193,In_360,In_171);
nand U194 (N_194,In_135,In_381);
nand U195 (N_195,In_473,N_128);
nor U196 (N_196,In_138,In_348);
and U197 (N_197,In_157,N_103);
nand U198 (N_198,N_24,N_122);
and U199 (N_199,In_290,In_86);
nand U200 (N_200,N_100,N_195);
or U201 (N_201,In_281,N_168);
and U202 (N_202,N_18,N_164);
xnor U203 (N_203,In_361,N_81);
xor U204 (N_204,N_16,In_164);
xnor U205 (N_205,N_45,N_171);
nor U206 (N_206,In_105,In_299);
or U207 (N_207,In_53,In_99);
nand U208 (N_208,In_236,In_68);
or U209 (N_209,N_25,N_93);
or U210 (N_210,N_189,In_467);
or U211 (N_211,In_78,In_73);
nand U212 (N_212,N_47,N_188);
nand U213 (N_213,N_52,N_179);
and U214 (N_214,In_349,N_64);
xor U215 (N_215,In_378,In_11);
nor U216 (N_216,N_180,N_127);
or U217 (N_217,In_203,In_364);
or U218 (N_218,N_60,In_321);
xor U219 (N_219,In_57,In_216);
and U220 (N_220,N_68,N_134);
nand U221 (N_221,N_174,In_476);
and U222 (N_222,In_107,In_116);
and U223 (N_223,N_106,N_78);
nor U224 (N_224,In_260,In_419);
nor U225 (N_225,In_110,N_139);
nor U226 (N_226,In_449,In_464);
and U227 (N_227,In_13,In_292);
and U228 (N_228,In_47,In_64);
or U229 (N_229,In_386,In_411);
nor U230 (N_230,In_210,In_474);
or U231 (N_231,N_48,In_486);
xnor U232 (N_232,In_69,N_186);
nor U233 (N_233,N_50,N_146);
and U234 (N_234,In_441,N_159);
xor U235 (N_235,N_111,In_432);
and U236 (N_236,N_133,In_313);
and U237 (N_237,N_99,In_178);
nand U238 (N_238,In_223,In_405);
xnor U239 (N_239,In_96,In_50);
and U240 (N_240,N_113,In_214);
and U241 (N_241,In_444,In_358);
nand U242 (N_242,N_35,In_407);
and U243 (N_243,In_218,In_375);
nand U244 (N_244,N_9,N_161);
xor U245 (N_245,N_102,In_239);
xnor U246 (N_246,In_243,N_104);
and U247 (N_247,In_77,N_124);
or U248 (N_248,In_265,N_61);
nor U249 (N_249,In_262,In_409);
or U250 (N_250,In_90,In_466);
nor U251 (N_251,N_40,In_426);
nor U252 (N_252,N_212,In_303);
or U253 (N_253,N_155,N_90);
nand U254 (N_254,N_105,N_145);
or U255 (N_255,N_190,N_125);
xor U256 (N_256,N_131,In_355);
and U257 (N_257,N_37,N_217);
or U258 (N_258,N_248,In_93);
or U259 (N_259,N_2,N_141);
xnor U260 (N_260,N_96,N_183);
xnor U261 (N_261,N_58,In_146);
and U262 (N_262,In_168,In_2);
nor U263 (N_263,In_75,N_182);
or U264 (N_264,In_436,In_179);
or U265 (N_265,In_120,In_144);
xor U266 (N_266,In_9,N_216);
nand U267 (N_267,N_169,N_185);
and U268 (N_268,N_230,N_80);
or U269 (N_269,N_196,N_234);
xor U270 (N_270,N_14,N_201);
nor U271 (N_271,In_359,In_304);
nor U272 (N_272,In_35,N_205);
or U273 (N_273,In_487,N_211);
xor U274 (N_274,N_206,In_285);
or U275 (N_275,N_181,N_108);
nor U276 (N_276,In_219,In_132);
and U277 (N_277,In_430,N_244);
xor U278 (N_278,N_22,N_178);
nand U279 (N_279,N_148,N_162);
nor U280 (N_280,In_365,In_111);
and U281 (N_281,In_48,N_135);
or U282 (N_282,N_28,N_76);
xnor U283 (N_283,In_257,N_231);
xnor U284 (N_284,N_15,N_71);
xnor U285 (N_285,N_153,N_218);
xnor U286 (N_286,N_163,N_191);
or U287 (N_287,In_309,N_34);
or U288 (N_288,N_110,In_417);
nor U289 (N_289,In_341,In_469);
nor U290 (N_290,N_207,N_89);
or U291 (N_291,N_221,In_200);
or U292 (N_292,N_91,In_458);
nand U293 (N_293,N_57,N_42);
and U294 (N_294,In_389,N_245);
nand U295 (N_295,In_82,N_235);
nand U296 (N_296,N_32,N_203);
nor U297 (N_297,N_55,N_233);
nand U298 (N_298,In_56,N_120);
and U299 (N_299,In_477,In_338);
or U300 (N_300,N_167,In_32);
nand U301 (N_301,N_194,In_70);
xor U302 (N_302,N_200,In_316);
or U303 (N_303,N_243,N_267);
xor U304 (N_304,In_324,In_126);
nand U305 (N_305,N_242,In_59);
and U306 (N_306,In_293,In_0);
xnor U307 (N_307,N_70,In_24);
nand U308 (N_308,N_213,N_223);
and U309 (N_309,N_271,N_294);
xnor U310 (N_310,N_249,In_492);
nor U311 (N_311,N_270,In_81);
nand U312 (N_312,In_36,In_197);
or U313 (N_313,N_293,In_182);
nand U314 (N_314,In_264,N_287);
nor U315 (N_315,In_112,N_256);
and U316 (N_316,In_496,N_227);
xnor U317 (N_317,In_154,In_51);
or U318 (N_318,N_41,In_198);
or U319 (N_319,N_266,N_214);
and U320 (N_320,N_275,N_150);
nor U321 (N_321,In_468,N_193);
nand U322 (N_322,N_151,In_102);
and U323 (N_323,N_263,N_187);
xor U324 (N_324,N_177,N_49);
nor U325 (N_325,N_192,N_289);
or U326 (N_326,N_225,N_278);
and U327 (N_327,In_163,In_80);
nor U328 (N_328,N_75,N_67);
nor U329 (N_329,N_209,N_117);
nand U330 (N_330,N_298,N_38);
nor U331 (N_331,N_296,N_288);
xor U332 (N_332,N_158,N_82);
nor U333 (N_333,N_228,N_97);
nor U334 (N_334,N_274,N_284);
and U335 (N_335,N_239,In_465);
nor U336 (N_336,N_157,N_247);
or U337 (N_337,N_238,In_425);
xnor U338 (N_338,N_10,N_114);
nand U339 (N_339,N_12,N_172);
and U340 (N_340,In_155,N_184);
and U341 (N_341,N_255,N_109);
nor U342 (N_342,In_230,In_326);
or U343 (N_343,N_254,N_208);
nand U344 (N_344,In_459,N_240);
xnor U345 (N_345,N_290,N_265);
and U346 (N_346,N_26,N_283);
or U347 (N_347,N_202,N_138);
nor U348 (N_348,N_237,N_295);
and U349 (N_349,In_336,N_5);
and U350 (N_350,N_340,N_337);
nor U351 (N_351,N_303,N_241);
or U352 (N_352,N_13,N_313);
and U353 (N_353,N_314,N_166);
and U354 (N_354,N_344,N_292);
or U355 (N_355,In_44,In_194);
and U356 (N_356,N_154,In_391);
nor U357 (N_357,In_490,N_160);
nand U358 (N_358,In_58,N_229);
nor U359 (N_359,N_318,N_316);
nor U360 (N_360,N_308,N_199);
and U361 (N_361,N_94,In_269);
nor U362 (N_362,N_269,N_152);
or U363 (N_363,N_62,N_330);
nand U364 (N_364,N_252,N_324);
nand U365 (N_365,N_220,N_197);
nor U366 (N_366,N_328,N_338);
xor U367 (N_367,N_334,N_349);
and U368 (N_368,N_6,N_281);
nand U369 (N_369,N_348,N_332);
nand U370 (N_370,N_170,N_280);
nor U371 (N_371,N_258,N_326);
nand U372 (N_372,In_284,N_321);
and U373 (N_373,N_310,N_272);
or U374 (N_374,N_333,N_219);
xnor U375 (N_375,N_302,N_325);
or U376 (N_376,In_478,N_53);
or U377 (N_377,N_279,In_335);
nor U378 (N_378,N_107,N_210);
or U379 (N_379,N_232,In_189);
xor U380 (N_380,N_336,N_304);
nand U381 (N_381,In_328,In_434);
or U382 (N_382,In_356,N_299);
nor U383 (N_383,N_329,N_277);
nand U384 (N_384,In_456,In_137);
nand U385 (N_385,N_250,N_317);
or U386 (N_386,N_339,N_307);
xnor U387 (N_387,N_260,In_489);
or U388 (N_388,N_215,In_213);
nor U389 (N_389,In_136,N_236);
nor U390 (N_390,N_305,N_286);
nand U391 (N_391,In_128,In_393);
xor U392 (N_392,N_331,In_453);
nor U393 (N_393,N_306,N_347);
and U394 (N_394,N_297,N_176);
and U395 (N_395,In_125,N_315);
nand U396 (N_396,N_345,N_116);
nand U397 (N_397,N_301,N_327);
and U398 (N_398,N_282,N_204);
nor U399 (N_399,In_318,N_147);
and U400 (N_400,N_361,In_206);
nand U401 (N_401,N_352,N_300);
and U402 (N_402,N_262,N_118);
and U403 (N_403,N_388,N_136);
and U404 (N_404,In_152,N_253);
nor U405 (N_405,N_378,N_396);
or U406 (N_406,N_322,In_10);
nand U407 (N_407,N_382,N_368);
nand U408 (N_408,N_83,N_3);
nand U409 (N_409,N_398,N_391);
nand U410 (N_410,N_273,N_360);
nor U411 (N_411,N_198,N_367);
or U412 (N_412,N_389,N_369);
and U413 (N_413,N_359,N_246);
and U414 (N_414,N_357,N_261);
nor U415 (N_415,N_393,N_251);
or U416 (N_416,N_355,N_354);
xnor U417 (N_417,N_311,N_309);
nand U418 (N_418,N_399,N_165);
nand U419 (N_419,N_385,N_30);
and U420 (N_420,N_370,N_374);
nand U421 (N_421,N_222,N_381);
and U422 (N_422,In_245,N_371);
and U423 (N_423,N_312,N_364);
xor U424 (N_424,N_365,N_175);
nor U425 (N_425,N_335,N_351);
xor U426 (N_426,N_341,N_346);
and U427 (N_427,N_377,N_372);
xnor U428 (N_428,N_342,N_320);
nand U429 (N_429,N_397,N_319);
and U430 (N_430,N_224,In_251);
and U431 (N_431,N_44,N_379);
nand U432 (N_432,N_257,N_259);
and U433 (N_433,N_264,N_375);
nand U434 (N_434,N_362,N_126);
nand U435 (N_435,N_390,N_226);
and U436 (N_436,N_358,N_291);
nor U437 (N_437,N_392,N_353);
nand U438 (N_438,N_394,N_343);
nand U439 (N_439,N_386,N_285);
nor U440 (N_440,N_395,N_380);
nand U441 (N_441,N_323,N_384);
and U442 (N_442,N_73,In_109);
nor U443 (N_443,N_373,N_363);
xnor U444 (N_444,N_376,N_383);
xor U445 (N_445,N_356,N_350);
nand U446 (N_446,N_156,N_387);
or U447 (N_447,N_173,N_8);
xor U448 (N_448,N_268,N_36);
nor U449 (N_449,N_276,N_366);
nand U450 (N_450,N_425,N_448);
nor U451 (N_451,N_427,N_429);
and U452 (N_452,N_421,N_406);
or U453 (N_453,N_435,N_409);
and U454 (N_454,N_400,N_423);
nand U455 (N_455,N_424,N_432);
or U456 (N_456,N_439,N_441);
and U457 (N_457,N_420,N_415);
xnor U458 (N_458,N_428,N_440);
and U459 (N_459,N_402,N_422);
nand U460 (N_460,N_412,N_417);
or U461 (N_461,N_401,N_446);
xor U462 (N_462,N_405,N_403);
xnor U463 (N_463,N_419,N_426);
xnor U464 (N_464,N_431,N_416);
nand U465 (N_465,N_436,N_430);
xor U466 (N_466,N_434,N_418);
nor U467 (N_467,N_413,N_442);
nand U468 (N_468,N_437,N_443);
xor U469 (N_469,N_444,N_438);
nor U470 (N_470,N_404,N_445);
and U471 (N_471,N_407,N_411);
or U472 (N_472,N_408,N_449);
or U473 (N_473,N_433,N_447);
and U474 (N_474,N_410,N_414);
nor U475 (N_475,N_430,N_402);
or U476 (N_476,N_403,N_440);
or U477 (N_477,N_402,N_424);
nand U478 (N_478,N_436,N_433);
and U479 (N_479,N_443,N_421);
or U480 (N_480,N_433,N_403);
or U481 (N_481,N_408,N_426);
nand U482 (N_482,N_445,N_412);
xor U483 (N_483,N_446,N_416);
or U484 (N_484,N_406,N_408);
and U485 (N_485,N_413,N_436);
and U486 (N_486,N_438,N_402);
xnor U487 (N_487,N_417,N_411);
or U488 (N_488,N_423,N_412);
xnor U489 (N_489,N_448,N_444);
xor U490 (N_490,N_449,N_429);
nor U491 (N_491,N_416,N_428);
or U492 (N_492,N_445,N_401);
nor U493 (N_493,N_401,N_441);
xnor U494 (N_494,N_408,N_429);
or U495 (N_495,N_431,N_445);
nor U496 (N_496,N_408,N_424);
and U497 (N_497,N_420,N_409);
nand U498 (N_498,N_425,N_429);
and U499 (N_499,N_422,N_417);
xnor U500 (N_500,N_474,N_464);
nand U501 (N_501,N_454,N_460);
and U502 (N_502,N_473,N_461);
nor U503 (N_503,N_468,N_485);
and U504 (N_504,N_486,N_457);
and U505 (N_505,N_496,N_497);
xnor U506 (N_506,N_479,N_491);
nor U507 (N_507,N_482,N_453);
nor U508 (N_508,N_470,N_488);
or U509 (N_509,N_467,N_475);
nand U510 (N_510,N_459,N_456);
xnor U511 (N_511,N_493,N_498);
xor U512 (N_512,N_451,N_499);
or U513 (N_513,N_494,N_469);
and U514 (N_514,N_484,N_480);
and U515 (N_515,N_458,N_495);
nand U516 (N_516,N_490,N_492);
xnor U517 (N_517,N_483,N_465);
or U518 (N_518,N_478,N_463);
and U519 (N_519,N_487,N_471);
and U520 (N_520,N_481,N_462);
and U521 (N_521,N_476,N_489);
or U522 (N_522,N_455,N_466);
xnor U523 (N_523,N_452,N_450);
nand U524 (N_524,N_477,N_472);
xnor U525 (N_525,N_455,N_481);
nand U526 (N_526,N_453,N_495);
or U527 (N_527,N_495,N_486);
nand U528 (N_528,N_493,N_452);
and U529 (N_529,N_463,N_498);
and U530 (N_530,N_483,N_492);
xor U531 (N_531,N_472,N_451);
xnor U532 (N_532,N_453,N_470);
and U533 (N_533,N_488,N_463);
nor U534 (N_534,N_496,N_498);
xor U535 (N_535,N_496,N_473);
nor U536 (N_536,N_481,N_453);
nand U537 (N_537,N_470,N_497);
nor U538 (N_538,N_459,N_460);
nand U539 (N_539,N_495,N_469);
nand U540 (N_540,N_495,N_450);
and U541 (N_541,N_499,N_459);
and U542 (N_542,N_489,N_452);
nand U543 (N_543,N_498,N_489);
xor U544 (N_544,N_468,N_469);
xnor U545 (N_545,N_461,N_488);
or U546 (N_546,N_464,N_488);
and U547 (N_547,N_474,N_466);
xnor U548 (N_548,N_451,N_465);
nand U549 (N_549,N_486,N_459);
or U550 (N_550,N_511,N_505);
and U551 (N_551,N_533,N_532);
or U552 (N_552,N_536,N_500);
nand U553 (N_553,N_529,N_502);
and U554 (N_554,N_540,N_528);
nor U555 (N_555,N_546,N_544);
and U556 (N_556,N_545,N_534);
nand U557 (N_557,N_522,N_501);
and U558 (N_558,N_503,N_510);
xnor U559 (N_559,N_538,N_508);
nor U560 (N_560,N_515,N_524);
xnor U561 (N_561,N_543,N_517);
and U562 (N_562,N_514,N_542);
nand U563 (N_563,N_521,N_504);
or U564 (N_564,N_527,N_530);
nor U565 (N_565,N_525,N_537);
and U566 (N_566,N_519,N_548);
nand U567 (N_567,N_549,N_516);
or U568 (N_568,N_547,N_535);
xnor U569 (N_569,N_513,N_509);
xnor U570 (N_570,N_506,N_523);
nand U571 (N_571,N_512,N_539);
and U572 (N_572,N_541,N_518);
xor U573 (N_573,N_531,N_507);
nor U574 (N_574,N_526,N_520);
and U575 (N_575,N_539,N_537);
nand U576 (N_576,N_509,N_511);
xnor U577 (N_577,N_522,N_518);
nor U578 (N_578,N_548,N_518);
and U579 (N_579,N_512,N_508);
or U580 (N_580,N_536,N_504);
or U581 (N_581,N_528,N_522);
or U582 (N_582,N_513,N_521);
and U583 (N_583,N_507,N_532);
and U584 (N_584,N_531,N_540);
xor U585 (N_585,N_503,N_501);
xor U586 (N_586,N_506,N_501);
nor U587 (N_587,N_530,N_540);
nor U588 (N_588,N_536,N_519);
and U589 (N_589,N_503,N_513);
or U590 (N_590,N_509,N_542);
nor U591 (N_591,N_549,N_538);
and U592 (N_592,N_506,N_526);
nand U593 (N_593,N_523,N_528);
nand U594 (N_594,N_507,N_542);
nand U595 (N_595,N_503,N_545);
nand U596 (N_596,N_522,N_549);
xor U597 (N_597,N_547,N_524);
or U598 (N_598,N_515,N_527);
nor U599 (N_599,N_533,N_502);
nand U600 (N_600,N_572,N_584);
xor U601 (N_601,N_597,N_579);
nand U602 (N_602,N_589,N_552);
nand U603 (N_603,N_565,N_553);
and U604 (N_604,N_592,N_594);
nand U605 (N_605,N_568,N_587);
nand U606 (N_606,N_566,N_570);
or U607 (N_607,N_580,N_581);
nor U608 (N_608,N_582,N_551);
xor U609 (N_609,N_586,N_567);
or U610 (N_610,N_596,N_598);
and U611 (N_611,N_556,N_558);
nand U612 (N_612,N_554,N_588);
and U613 (N_613,N_569,N_575);
nor U614 (N_614,N_590,N_577);
xor U615 (N_615,N_573,N_595);
xnor U616 (N_616,N_574,N_583);
xnor U617 (N_617,N_560,N_561);
xnor U618 (N_618,N_576,N_571);
or U619 (N_619,N_591,N_550);
or U620 (N_620,N_578,N_585);
and U621 (N_621,N_557,N_562);
nor U622 (N_622,N_555,N_559);
and U623 (N_623,N_564,N_593);
nand U624 (N_624,N_563,N_599);
nand U625 (N_625,N_558,N_565);
nor U626 (N_626,N_572,N_555);
nor U627 (N_627,N_562,N_558);
and U628 (N_628,N_572,N_599);
xnor U629 (N_629,N_568,N_582);
nand U630 (N_630,N_590,N_567);
and U631 (N_631,N_558,N_572);
or U632 (N_632,N_597,N_565);
nand U633 (N_633,N_591,N_559);
nor U634 (N_634,N_565,N_578);
xnor U635 (N_635,N_579,N_556);
and U636 (N_636,N_576,N_560);
and U637 (N_637,N_575,N_598);
xor U638 (N_638,N_556,N_553);
or U639 (N_639,N_551,N_571);
xnor U640 (N_640,N_558,N_576);
and U641 (N_641,N_567,N_591);
nand U642 (N_642,N_571,N_591);
nand U643 (N_643,N_583,N_550);
xor U644 (N_644,N_596,N_573);
or U645 (N_645,N_595,N_555);
or U646 (N_646,N_586,N_590);
and U647 (N_647,N_585,N_557);
or U648 (N_648,N_559,N_598);
nand U649 (N_649,N_599,N_568);
xor U650 (N_650,N_641,N_605);
nand U651 (N_651,N_645,N_639);
nor U652 (N_652,N_618,N_625);
xor U653 (N_653,N_606,N_635);
and U654 (N_654,N_611,N_604);
nand U655 (N_655,N_621,N_649);
nor U656 (N_656,N_640,N_629);
nor U657 (N_657,N_624,N_610);
nor U658 (N_658,N_647,N_638);
and U659 (N_659,N_648,N_630);
or U660 (N_660,N_643,N_633);
xor U661 (N_661,N_631,N_607);
and U662 (N_662,N_632,N_620);
nor U663 (N_663,N_636,N_637);
nand U664 (N_664,N_622,N_627);
nand U665 (N_665,N_628,N_619);
and U666 (N_666,N_615,N_613);
nand U667 (N_667,N_602,N_634);
or U668 (N_668,N_616,N_603);
xor U669 (N_669,N_612,N_608);
or U670 (N_670,N_623,N_642);
or U671 (N_671,N_617,N_626);
or U672 (N_672,N_614,N_601);
nand U673 (N_673,N_646,N_609);
nand U674 (N_674,N_644,N_600);
xor U675 (N_675,N_607,N_627);
or U676 (N_676,N_601,N_649);
or U677 (N_677,N_639,N_619);
and U678 (N_678,N_602,N_644);
or U679 (N_679,N_643,N_605);
nand U680 (N_680,N_623,N_608);
xor U681 (N_681,N_646,N_624);
and U682 (N_682,N_613,N_635);
nand U683 (N_683,N_630,N_645);
nor U684 (N_684,N_634,N_614);
nor U685 (N_685,N_632,N_609);
xor U686 (N_686,N_631,N_602);
or U687 (N_687,N_637,N_633);
nor U688 (N_688,N_612,N_624);
nor U689 (N_689,N_627,N_629);
nand U690 (N_690,N_613,N_620);
nor U691 (N_691,N_600,N_605);
nand U692 (N_692,N_613,N_639);
and U693 (N_693,N_631,N_633);
nand U694 (N_694,N_600,N_611);
xor U695 (N_695,N_602,N_647);
xor U696 (N_696,N_602,N_606);
or U697 (N_697,N_622,N_642);
and U698 (N_698,N_623,N_626);
xor U699 (N_699,N_616,N_601);
xor U700 (N_700,N_669,N_677);
nor U701 (N_701,N_685,N_661);
and U702 (N_702,N_692,N_660);
or U703 (N_703,N_650,N_699);
nor U704 (N_704,N_687,N_680);
or U705 (N_705,N_670,N_690);
nand U706 (N_706,N_683,N_689);
or U707 (N_707,N_686,N_658);
nor U708 (N_708,N_674,N_672);
and U709 (N_709,N_691,N_681);
xor U710 (N_710,N_676,N_652);
and U711 (N_711,N_651,N_696);
nand U712 (N_712,N_679,N_693);
xor U713 (N_713,N_665,N_671);
and U714 (N_714,N_656,N_675);
and U715 (N_715,N_664,N_655);
xnor U716 (N_716,N_667,N_666);
and U717 (N_717,N_663,N_662);
or U718 (N_718,N_697,N_695);
and U719 (N_719,N_694,N_673);
nand U720 (N_720,N_688,N_668);
xor U721 (N_721,N_698,N_653);
nand U722 (N_722,N_657,N_678);
and U723 (N_723,N_654,N_682);
xor U724 (N_724,N_684,N_659);
and U725 (N_725,N_654,N_668);
and U726 (N_726,N_653,N_672);
or U727 (N_727,N_680,N_688);
xnor U728 (N_728,N_686,N_661);
or U729 (N_729,N_696,N_691);
nor U730 (N_730,N_655,N_662);
nor U731 (N_731,N_688,N_695);
xor U732 (N_732,N_651,N_669);
xnor U733 (N_733,N_686,N_668);
xnor U734 (N_734,N_667,N_684);
nand U735 (N_735,N_674,N_693);
nand U736 (N_736,N_657,N_679);
or U737 (N_737,N_657,N_675);
nor U738 (N_738,N_686,N_662);
nand U739 (N_739,N_668,N_666);
nor U740 (N_740,N_673,N_690);
or U741 (N_741,N_680,N_661);
nand U742 (N_742,N_651,N_662);
nand U743 (N_743,N_670,N_657);
or U744 (N_744,N_681,N_654);
xnor U745 (N_745,N_692,N_676);
nor U746 (N_746,N_664,N_658);
and U747 (N_747,N_691,N_673);
xnor U748 (N_748,N_698,N_673);
or U749 (N_749,N_657,N_667);
nand U750 (N_750,N_749,N_714);
or U751 (N_751,N_710,N_702);
or U752 (N_752,N_730,N_744);
xnor U753 (N_753,N_706,N_739);
nor U754 (N_754,N_712,N_707);
nand U755 (N_755,N_742,N_715);
nor U756 (N_756,N_713,N_704);
or U757 (N_757,N_711,N_720);
nand U758 (N_758,N_731,N_732);
nand U759 (N_759,N_716,N_722);
and U760 (N_760,N_723,N_747);
or U761 (N_761,N_738,N_703);
nand U762 (N_762,N_726,N_740);
xnor U763 (N_763,N_721,N_735);
nor U764 (N_764,N_717,N_748);
nand U765 (N_765,N_746,N_708);
or U766 (N_766,N_743,N_737);
nor U767 (N_767,N_724,N_700);
nand U768 (N_768,N_736,N_745);
nand U769 (N_769,N_727,N_728);
nor U770 (N_770,N_718,N_719);
and U771 (N_771,N_701,N_729);
xnor U772 (N_772,N_734,N_725);
nor U773 (N_773,N_741,N_705);
nor U774 (N_774,N_733,N_709);
and U775 (N_775,N_740,N_704);
nand U776 (N_776,N_732,N_718);
nor U777 (N_777,N_718,N_733);
nor U778 (N_778,N_746,N_747);
nand U779 (N_779,N_738,N_728);
xnor U780 (N_780,N_731,N_725);
or U781 (N_781,N_716,N_736);
nand U782 (N_782,N_722,N_745);
nor U783 (N_783,N_723,N_700);
or U784 (N_784,N_704,N_714);
nor U785 (N_785,N_717,N_700);
xor U786 (N_786,N_724,N_748);
xnor U787 (N_787,N_748,N_737);
nand U788 (N_788,N_718,N_737);
nand U789 (N_789,N_717,N_742);
and U790 (N_790,N_718,N_744);
nand U791 (N_791,N_743,N_733);
nor U792 (N_792,N_729,N_719);
or U793 (N_793,N_748,N_713);
and U794 (N_794,N_748,N_702);
xnor U795 (N_795,N_721,N_737);
nand U796 (N_796,N_748,N_726);
nand U797 (N_797,N_737,N_702);
and U798 (N_798,N_701,N_728);
or U799 (N_799,N_746,N_737);
nor U800 (N_800,N_766,N_772);
xnor U801 (N_801,N_786,N_751);
nor U802 (N_802,N_782,N_799);
and U803 (N_803,N_756,N_776);
nand U804 (N_804,N_778,N_784);
xor U805 (N_805,N_754,N_774);
nand U806 (N_806,N_768,N_753);
nor U807 (N_807,N_762,N_761);
nand U808 (N_808,N_755,N_791);
nor U809 (N_809,N_794,N_773);
and U810 (N_810,N_758,N_783);
and U811 (N_811,N_764,N_790);
xor U812 (N_812,N_779,N_788);
or U813 (N_813,N_785,N_789);
and U814 (N_814,N_792,N_770);
nand U815 (N_815,N_771,N_777);
and U816 (N_816,N_793,N_797);
and U817 (N_817,N_763,N_750);
nor U818 (N_818,N_796,N_760);
or U819 (N_819,N_795,N_775);
nand U820 (N_820,N_767,N_781);
and U821 (N_821,N_787,N_769);
xor U822 (N_822,N_780,N_757);
and U823 (N_823,N_765,N_759);
xnor U824 (N_824,N_752,N_798);
and U825 (N_825,N_788,N_790);
nand U826 (N_826,N_798,N_787);
and U827 (N_827,N_773,N_785);
nand U828 (N_828,N_760,N_762);
xnor U829 (N_829,N_768,N_778);
nand U830 (N_830,N_797,N_782);
and U831 (N_831,N_778,N_798);
xor U832 (N_832,N_797,N_751);
or U833 (N_833,N_794,N_777);
and U834 (N_834,N_756,N_772);
nor U835 (N_835,N_796,N_761);
nor U836 (N_836,N_768,N_793);
xnor U837 (N_837,N_774,N_796);
nand U838 (N_838,N_753,N_754);
xnor U839 (N_839,N_793,N_780);
nor U840 (N_840,N_768,N_797);
nand U841 (N_841,N_776,N_765);
and U842 (N_842,N_765,N_775);
and U843 (N_843,N_756,N_790);
nor U844 (N_844,N_790,N_775);
xor U845 (N_845,N_789,N_780);
or U846 (N_846,N_758,N_798);
or U847 (N_847,N_784,N_781);
xnor U848 (N_848,N_772,N_788);
nor U849 (N_849,N_771,N_757);
or U850 (N_850,N_841,N_846);
xor U851 (N_851,N_842,N_806);
nand U852 (N_852,N_819,N_839);
nor U853 (N_853,N_828,N_803);
xor U854 (N_854,N_836,N_840);
xnor U855 (N_855,N_843,N_834);
xor U856 (N_856,N_824,N_845);
and U857 (N_857,N_800,N_832);
or U858 (N_858,N_807,N_829);
and U859 (N_859,N_847,N_826);
nor U860 (N_860,N_814,N_825);
nand U861 (N_861,N_823,N_817);
nor U862 (N_862,N_849,N_822);
nor U863 (N_863,N_801,N_830);
nor U864 (N_864,N_810,N_833);
nor U865 (N_865,N_805,N_848);
nand U866 (N_866,N_812,N_815);
nor U867 (N_867,N_816,N_844);
nand U868 (N_868,N_813,N_827);
and U869 (N_869,N_837,N_838);
and U870 (N_870,N_818,N_835);
or U871 (N_871,N_821,N_809);
xnor U872 (N_872,N_811,N_808);
nand U873 (N_873,N_804,N_802);
nor U874 (N_874,N_820,N_831);
and U875 (N_875,N_830,N_817);
or U876 (N_876,N_847,N_835);
xnor U877 (N_877,N_827,N_849);
xnor U878 (N_878,N_843,N_816);
xor U879 (N_879,N_839,N_809);
and U880 (N_880,N_817,N_843);
nand U881 (N_881,N_808,N_806);
nor U882 (N_882,N_812,N_811);
xnor U883 (N_883,N_806,N_801);
nand U884 (N_884,N_802,N_803);
or U885 (N_885,N_835,N_823);
xnor U886 (N_886,N_826,N_805);
xnor U887 (N_887,N_806,N_834);
xor U888 (N_888,N_807,N_847);
or U889 (N_889,N_832,N_835);
nor U890 (N_890,N_815,N_811);
or U891 (N_891,N_834,N_825);
or U892 (N_892,N_847,N_838);
and U893 (N_893,N_849,N_811);
xor U894 (N_894,N_839,N_847);
nor U895 (N_895,N_843,N_807);
nor U896 (N_896,N_806,N_824);
or U897 (N_897,N_838,N_808);
or U898 (N_898,N_829,N_817);
and U899 (N_899,N_817,N_808);
nand U900 (N_900,N_889,N_898);
xnor U901 (N_901,N_855,N_861);
nand U902 (N_902,N_869,N_874);
or U903 (N_903,N_875,N_876);
nand U904 (N_904,N_899,N_894);
nand U905 (N_905,N_862,N_892);
nand U906 (N_906,N_860,N_878);
nand U907 (N_907,N_882,N_851);
xnor U908 (N_908,N_853,N_852);
and U909 (N_909,N_888,N_856);
xnor U910 (N_910,N_873,N_871);
nand U911 (N_911,N_893,N_895);
and U912 (N_912,N_890,N_872);
nor U913 (N_913,N_891,N_857);
or U914 (N_914,N_896,N_864);
nand U915 (N_915,N_866,N_863);
nor U916 (N_916,N_850,N_880);
and U917 (N_917,N_897,N_886);
nand U918 (N_918,N_881,N_877);
xnor U919 (N_919,N_859,N_879);
nor U920 (N_920,N_867,N_868);
and U921 (N_921,N_885,N_865);
and U922 (N_922,N_884,N_887);
xor U923 (N_923,N_870,N_883);
or U924 (N_924,N_858,N_854);
nand U925 (N_925,N_895,N_871);
xnor U926 (N_926,N_851,N_894);
nand U927 (N_927,N_887,N_881);
and U928 (N_928,N_851,N_860);
xnor U929 (N_929,N_891,N_885);
xor U930 (N_930,N_879,N_898);
nand U931 (N_931,N_859,N_895);
or U932 (N_932,N_875,N_895);
nand U933 (N_933,N_860,N_884);
xnor U934 (N_934,N_898,N_867);
and U935 (N_935,N_856,N_855);
nand U936 (N_936,N_852,N_888);
or U937 (N_937,N_883,N_871);
xor U938 (N_938,N_879,N_865);
nor U939 (N_939,N_895,N_868);
nor U940 (N_940,N_866,N_875);
or U941 (N_941,N_872,N_859);
xnor U942 (N_942,N_874,N_870);
nand U943 (N_943,N_884,N_858);
and U944 (N_944,N_852,N_861);
or U945 (N_945,N_878,N_888);
xor U946 (N_946,N_859,N_891);
or U947 (N_947,N_871,N_898);
and U948 (N_948,N_862,N_896);
nand U949 (N_949,N_876,N_860);
and U950 (N_950,N_936,N_902);
xnor U951 (N_951,N_937,N_948);
xnor U952 (N_952,N_921,N_949);
or U953 (N_953,N_939,N_926);
xor U954 (N_954,N_944,N_947);
or U955 (N_955,N_901,N_930);
and U956 (N_956,N_943,N_941);
nor U957 (N_957,N_940,N_903);
and U958 (N_958,N_917,N_924);
xor U959 (N_959,N_928,N_932);
nor U960 (N_960,N_918,N_908);
and U961 (N_961,N_905,N_909);
nand U962 (N_962,N_922,N_927);
or U963 (N_963,N_910,N_914);
and U964 (N_964,N_911,N_915);
nor U965 (N_965,N_935,N_934);
or U966 (N_966,N_931,N_938);
and U967 (N_967,N_907,N_942);
xor U968 (N_968,N_906,N_913);
nand U969 (N_969,N_916,N_925);
or U970 (N_970,N_912,N_919);
nand U971 (N_971,N_923,N_920);
xnor U972 (N_972,N_929,N_946);
nand U973 (N_973,N_900,N_904);
nand U974 (N_974,N_945,N_933);
nor U975 (N_975,N_930,N_917);
or U976 (N_976,N_932,N_935);
or U977 (N_977,N_921,N_917);
nand U978 (N_978,N_938,N_940);
nor U979 (N_979,N_941,N_921);
nor U980 (N_980,N_940,N_947);
nor U981 (N_981,N_943,N_946);
nand U982 (N_982,N_905,N_906);
or U983 (N_983,N_921,N_928);
nand U984 (N_984,N_937,N_901);
nand U985 (N_985,N_928,N_926);
xor U986 (N_986,N_939,N_944);
nand U987 (N_987,N_949,N_926);
nor U988 (N_988,N_923,N_947);
or U989 (N_989,N_923,N_943);
nor U990 (N_990,N_905,N_926);
nor U991 (N_991,N_922,N_920);
and U992 (N_992,N_929,N_908);
or U993 (N_993,N_949,N_929);
and U994 (N_994,N_930,N_910);
xnor U995 (N_995,N_947,N_900);
xor U996 (N_996,N_944,N_930);
or U997 (N_997,N_926,N_916);
nand U998 (N_998,N_935,N_941);
nor U999 (N_999,N_905,N_939);
or U1000 (N_1000,N_967,N_980);
and U1001 (N_1001,N_969,N_962);
xnor U1002 (N_1002,N_977,N_979);
or U1003 (N_1003,N_987,N_995);
or U1004 (N_1004,N_958,N_990);
and U1005 (N_1005,N_981,N_965);
or U1006 (N_1006,N_974,N_955);
nor U1007 (N_1007,N_957,N_970);
nand U1008 (N_1008,N_971,N_973);
nand U1009 (N_1009,N_993,N_978);
nand U1010 (N_1010,N_997,N_983);
nor U1011 (N_1011,N_972,N_963);
xnor U1012 (N_1012,N_992,N_960);
or U1013 (N_1013,N_952,N_951);
xnor U1014 (N_1014,N_982,N_998);
or U1015 (N_1015,N_984,N_996);
nand U1016 (N_1016,N_989,N_966);
nor U1017 (N_1017,N_956,N_988);
nand U1018 (N_1018,N_953,N_964);
xnor U1019 (N_1019,N_994,N_975);
or U1020 (N_1020,N_986,N_976);
xnor U1021 (N_1021,N_999,N_985);
nand U1022 (N_1022,N_991,N_961);
and U1023 (N_1023,N_950,N_968);
nand U1024 (N_1024,N_954,N_959);
nand U1025 (N_1025,N_971,N_950);
and U1026 (N_1026,N_985,N_956);
xnor U1027 (N_1027,N_991,N_951);
nand U1028 (N_1028,N_993,N_950);
nor U1029 (N_1029,N_978,N_954);
xor U1030 (N_1030,N_967,N_987);
or U1031 (N_1031,N_995,N_993);
and U1032 (N_1032,N_983,N_970);
nand U1033 (N_1033,N_992,N_954);
nand U1034 (N_1034,N_952,N_997);
or U1035 (N_1035,N_963,N_984);
or U1036 (N_1036,N_965,N_990);
xor U1037 (N_1037,N_961,N_965);
or U1038 (N_1038,N_979,N_952);
or U1039 (N_1039,N_951,N_959);
xor U1040 (N_1040,N_958,N_998);
or U1041 (N_1041,N_967,N_969);
or U1042 (N_1042,N_953,N_984);
nor U1043 (N_1043,N_980,N_955);
or U1044 (N_1044,N_973,N_962);
nand U1045 (N_1045,N_954,N_967);
nor U1046 (N_1046,N_992,N_978);
and U1047 (N_1047,N_992,N_984);
nor U1048 (N_1048,N_950,N_988);
or U1049 (N_1049,N_989,N_978);
or U1050 (N_1050,N_1041,N_1034);
nor U1051 (N_1051,N_1014,N_1039);
nor U1052 (N_1052,N_1020,N_1038);
xnor U1053 (N_1053,N_1001,N_1036);
xnor U1054 (N_1054,N_1025,N_1030);
or U1055 (N_1055,N_1049,N_1045);
nor U1056 (N_1056,N_1007,N_1016);
nand U1057 (N_1057,N_1005,N_1003);
xnor U1058 (N_1058,N_1009,N_1040);
nor U1059 (N_1059,N_1017,N_1033);
xnor U1060 (N_1060,N_1031,N_1013);
nand U1061 (N_1061,N_1019,N_1006);
xnor U1062 (N_1062,N_1023,N_1002);
xnor U1063 (N_1063,N_1018,N_1027);
or U1064 (N_1064,N_1011,N_1012);
and U1065 (N_1065,N_1044,N_1035);
or U1066 (N_1066,N_1024,N_1021);
or U1067 (N_1067,N_1046,N_1037);
nand U1068 (N_1068,N_1015,N_1026);
nor U1069 (N_1069,N_1043,N_1029);
nor U1070 (N_1070,N_1010,N_1042);
or U1071 (N_1071,N_1032,N_1004);
and U1072 (N_1072,N_1022,N_1008);
and U1073 (N_1073,N_1048,N_1028);
nand U1074 (N_1074,N_1000,N_1047);
or U1075 (N_1075,N_1044,N_1046);
xnor U1076 (N_1076,N_1021,N_1033);
xor U1077 (N_1077,N_1015,N_1038);
nand U1078 (N_1078,N_1002,N_1027);
and U1079 (N_1079,N_1021,N_1042);
and U1080 (N_1080,N_1049,N_1047);
nand U1081 (N_1081,N_1000,N_1039);
xor U1082 (N_1082,N_1005,N_1031);
xor U1083 (N_1083,N_1009,N_1031);
and U1084 (N_1084,N_1019,N_1014);
and U1085 (N_1085,N_1037,N_1027);
and U1086 (N_1086,N_1013,N_1029);
nor U1087 (N_1087,N_1030,N_1012);
and U1088 (N_1088,N_1037,N_1048);
and U1089 (N_1089,N_1014,N_1001);
nor U1090 (N_1090,N_1002,N_1043);
nor U1091 (N_1091,N_1011,N_1043);
nor U1092 (N_1092,N_1045,N_1006);
nand U1093 (N_1093,N_1020,N_1014);
nor U1094 (N_1094,N_1025,N_1046);
nor U1095 (N_1095,N_1025,N_1022);
and U1096 (N_1096,N_1037,N_1049);
and U1097 (N_1097,N_1007,N_1032);
nor U1098 (N_1098,N_1049,N_1012);
or U1099 (N_1099,N_1036,N_1045);
or U1100 (N_1100,N_1071,N_1075);
xor U1101 (N_1101,N_1069,N_1083);
and U1102 (N_1102,N_1099,N_1096);
nor U1103 (N_1103,N_1094,N_1066);
and U1104 (N_1104,N_1087,N_1090);
and U1105 (N_1105,N_1062,N_1091);
nor U1106 (N_1106,N_1074,N_1052);
and U1107 (N_1107,N_1061,N_1080);
or U1108 (N_1108,N_1073,N_1076);
nor U1109 (N_1109,N_1086,N_1068);
and U1110 (N_1110,N_1079,N_1051);
nor U1111 (N_1111,N_1098,N_1053);
nor U1112 (N_1112,N_1092,N_1067);
nand U1113 (N_1113,N_1059,N_1082);
or U1114 (N_1114,N_1055,N_1070);
or U1115 (N_1115,N_1093,N_1089);
nand U1116 (N_1116,N_1064,N_1060);
nand U1117 (N_1117,N_1084,N_1058);
and U1118 (N_1118,N_1057,N_1056);
or U1119 (N_1119,N_1072,N_1065);
or U1120 (N_1120,N_1063,N_1050);
xor U1121 (N_1121,N_1077,N_1081);
nand U1122 (N_1122,N_1054,N_1085);
xnor U1123 (N_1123,N_1097,N_1095);
nor U1124 (N_1124,N_1088,N_1078);
or U1125 (N_1125,N_1078,N_1052);
and U1126 (N_1126,N_1064,N_1075);
and U1127 (N_1127,N_1059,N_1078);
xnor U1128 (N_1128,N_1091,N_1085);
and U1129 (N_1129,N_1052,N_1073);
nand U1130 (N_1130,N_1085,N_1077);
xnor U1131 (N_1131,N_1093,N_1087);
nor U1132 (N_1132,N_1095,N_1098);
xor U1133 (N_1133,N_1086,N_1069);
and U1134 (N_1134,N_1096,N_1071);
xor U1135 (N_1135,N_1073,N_1092);
and U1136 (N_1136,N_1058,N_1096);
or U1137 (N_1137,N_1088,N_1084);
or U1138 (N_1138,N_1074,N_1051);
or U1139 (N_1139,N_1097,N_1094);
and U1140 (N_1140,N_1073,N_1074);
and U1141 (N_1141,N_1069,N_1082);
xnor U1142 (N_1142,N_1077,N_1062);
or U1143 (N_1143,N_1083,N_1081);
nand U1144 (N_1144,N_1055,N_1097);
xnor U1145 (N_1145,N_1061,N_1073);
and U1146 (N_1146,N_1073,N_1081);
nand U1147 (N_1147,N_1076,N_1079);
xnor U1148 (N_1148,N_1078,N_1054);
nor U1149 (N_1149,N_1064,N_1094);
and U1150 (N_1150,N_1146,N_1119);
nand U1151 (N_1151,N_1137,N_1113);
and U1152 (N_1152,N_1106,N_1108);
and U1153 (N_1153,N_1143,N_1118);
or U1154 (N_1154,N_1122,N_1134);
nor U1155 (N_1155,N_1110,N_1131);
and U1156 (N_1156,N_1132,N_1123);
nor U1157 (N_1157,N_1136,N_1140);
nor U1158 (N_1158,N_1124,N_1149);
nand U1159 (N_1159,N_1126,N_1148);
and U1160 (N_1160,N_1142,N_1121);
xnor U1161 (N_1161,N_1109,N_1111);
nor U1162 (N_1162,N_1128,N_1133);
and U1163 (N_1163,N_1129,N_1138);
nand U1164 (N_1164,N_1112,N_1120);
and U1165 (N_1165,N_1114,N_1141);
or U1166 (N_1166,N_1102,N_1104);
nor U1167 (N_1167,N_1116,N_1107);
nand U1168 (N_1168,N_1115,N_1147);
xnor U1169 (N_1169,N_1105,N_1135);
nor U1170 (N_1170,N_1117,N_1103);
xor U1171 (N_1171,N_1130,N_1144);
or U1172 (N_1172,N_1100,N_1101);
nand U1173 (N_1173,N_1127,N_1145);
nor U1174 (N_1174,N_1125,N_1139);
nor U1175 (N_1175,N_1146,N_1111);
nand U1176 (N_1176,N_1123,N_1111);
xor U1177 (N_1177,N_1127,N_1133);
nor U1178 (N_1178,N_1145,N_1126);
nor U1179 (N_1179,N_1100,N_1106);
or U1180 (N_1180,N_1134,N_1141);
or U1181 (N_1181,N_1129,N_1141);
and U1182 (N_1182,N_1140,N_1109);
xor U1183 (N_1183,N_1112,N_1128);
nand U1184 (N_1184,N_1124,N_1128);
and U1185 (N_1185,N_1106,N_1103);
nand U1186 (N_1186,N_1101,N_1135);
xnor U1187 (N_1187,N_1102,N_1141);
xor U1188 (N_1188,N_1108,N_1147);
and U1189 (N_1189,N_1112,N_1114);
nor U1190 (N_1190,N_1113,N_1100);
xor U1191 (N_1191,N_1108,N_1110);
xor U1192 (N_1192,N_1142,N_1149);
or U1193 (N_1193,N_1120,N_1121);
xor U1194 (N_1194,N_1105,N_1141);
xor U1195 (N_1195,N_1101,N_1146);
nand U1196 (N_1196,N_1125,N_1131);
or U1197 (N_1197,N_1132,N_1145);
xnor U1198 (N_1198,N_1124,N_1125);
nor U1199 (N_1199,N_1124,N_1146);
and U1200 (N_1200,N_1188,N_1176);
nand U1201 (N_1201,N_1165,N_1192);
or U1202 (N_1202,N_1155,N_1181);
and U1203 (N_1203,N_1193,N_1191);
and U1204 (N_1204,N_1158,N_1185);
or U1205 (N_1205,N_1177,N_1167);
xor U1206 (N_1206,N_1164,N_1163);
or U1207 (N_1207,N_1162,N_1189);
xor U1208 (N_1208,N_1173,N_1156);
nor U1209 (N_1209,N_1187,N_1153);
nor U1210 (N_1210,N_1184,N_1150);
nor U1211 (N_1211,N_1199,N_1194);
and U1212 (N_1212,N_1197,N_1157);
xor U1213 (N_1213,N_1198,N_1179);
and U1214 (N_1214,N_1174,N_1168);
nor U1215 (N_1215,N_1196,N_1190);
nor U1216 (N_1216,N_1186,N_1159);
or U1217 (N_1217,N_1178,N_1169);
or U1218 (N_1218,N_1154,N_1166);
xnor U1219 (N_1219,N_1180,N_1172);
xnor U1220 (N_1220,N_1171,N_1175);
nor U1221 (N_1221,N_1170,N_1151);
nor U1222 (N_1222,N_1183,N_1160);
nand U1223 (N_1223,N_1182,N_1161);
and U1224 (N_1224,N_1195,N_1152);
and U1225 (N_1225,N_1174,N_1161);
or U1226 (N_1226,N_1171,N_1182);
or U1227 (N_1227,N_1192,N_1195);
nor U1228 (N_1228,N_1167,N_1187);
nand U1229 (N_1229,N_1161,N_1150);
or U1230 (N_1230,N_1150,N_1185);
xor U1231 (N_1231,N_1150,N_1162);
xor U1232 (N_1232,N_1197,N_1196);
nand U1233 (N_1233,N_1157,N_1151);
nor U1234 (N_1234,N_1185,N_1189);
xnor U1235 (N_1235,N_1199,N_1171);
nor U1236 (N_1236,N_1165,N_1154);
nand U1237 (N_1237,N_1181,N_1157);
xnor U1238 (N_1238,N_1181,N_1187);
nand U1239 (N_1239,N_1180,N_1166);
nand U1240 (N_1240,N_1175,N_1153);
xor U1241 (N_1241,N_1160,N_1189);
nor U1242 (N_1242,N_1191,N_1179);
xnor U1243 (N_1243,N_1199,N_1183);
or U1244 (N_1244,N_1198,N_1158);
xor U1245 (N_1245,N_1165,N_1179);
or U1246 (N_1246,N_1165,N_1177);
nand U1247 (N_1247,N_1197,N_1160);
and U1248 (N_1248,N_1182,N_1175);
or U1249 (N_1249,N_1168,N_1171);
nand U1250 (N_1250,N_1222,N_1202);
nor U1251 (N_1251,N_1210,N_1241);
nor U1252 (N_1252,N_1234,N_1218);
xor U1253 (N_1253,N_1220,N_1200);
xor U1254 (N_1254,N_1215,N_1208);
nor U1255 (N_1255,N_1242,N_1236);
nand U1256 (N_1256,N_1227,N_1226);
nand U1257 (N_1257,N_1211,N_1206);
xor U1258 (N_1258,N_1230,N_1209);
xor U1259 (N_1259,N_1229,N_1232);
and U1260 (N_1260,N_1225,N_1213);
xnor U1261 (N_1261,N_1245,N_1244);
and U1262 (N_1262,N_1239,N_1216);
nor U1263 (N_1263,N_1212,N_1228);
nand U1264 (N_1264,N_1203,N_1237);
nand U1265 (N_1265,N_1235,N_1233);
or U1266 (N_1266,N_1231,N_1238);
xnor U1267 (N_1267,N_1221,N_1240);
and U1268 (N_1268,N_1207,N_1205);
nor U1269 (N_1269,N_1219,N_1243);
or U1270 (N_1270,N_1204,N_1248);
and U1271 (N_1271,N_1217,N_1201);
xnor U1272 (N_1272,N_1249,N_1214);
or U1273 (N_1273,N_1223,N_1224);
nand U1274 (N_1274,N_1247,N_1246);
xor U1275 (N_1275,N_1217,N_1200);
xor U1276 (N_1276,N_1203,N_1226);
and U1277 (N_1277,N_1208,N_1211);
or U1278 (N_1278,N_1203,N_1235);
nor U1279 (N_1279,N_1232,N_1220);
nand U1280 (N_1280,N_1242,N_1234);
xor U1281 (N_1281,N_1206,N_1230);
nand U1282 (N_1282,N_1222,N_1220);
or U1283 (N_1283,N_1212,N_1220);
or U1284 (N_1284,N_1234,N_1244);
nor U1285 (N_1285,N_1242,N_1218);
nor U1286 (N_1286,N_1201,N_1230);
nor U1287 (N_1287,N_1225,N_1201);
or U1288 (N_1288,N_1204,N_1211);
or U1289 (N_1289,N_1206,N_1232);
nand U1290 (N_1290,N_1236,N_1214);
or U1291 (N_1291,N_1204,N_1202);
nand U1292 (N_1292,N_1205,N_1235);
nor U1293 (N_1293,N_1246,N_1237);
and U1294 (N_1294,N_1210,N_1220);
or U1295 (N_1295,N_1230,N_1218);
nor U1296 (N_1296,N_1200,N_1242);
xnor U1297 (N_1297,N_1204,N_1224);
nor U1298 (N_1298,N_1233,N_1225);
nand U1299 (N_1299,N_1208,N_1213);
or U1300 (N_1300,N_1296,N_1268);
xor U1301 (N_1301,N_1292,N_1257);
nand U1302 (N_1302,N_1277,N_1283);
nand U1303 (N_1303,N_1265,N_1297);
or U1304 (N_1304,N_1280,N_1267);
xnor U1305 (N_1305,N_1295,N_1278);
xnor U1306 (N_1306,N_1270,N_1293);
xor U1307 (N_1307,N_1282,N_1259);
and U1308 (N_1308,N_1284,N_1298);
xnor U1309 (N_1309,N_1287,N_1281);
xor U1310 (N_1310,N_1262,N_1254);
nand U1311 (N_1311,N_1285,N_1290);
nand U1312 (N_1312,N_1266,N_1286);
or U1313 (N_1313,N_1255,N_1252);
nor U1314 (N_1314,N_1299,N_1263);
or U1315 (N_1315,N_1253,N_1258);
xnor U1316 (N_1316,N_1272,N_1289);
nor U1317 (N_1317,N_1291,N_1256);
xnor U1318 (N_1318,N_1261,N_1294);
or U1319 (N_1319,N_1276,N_1279);
nand U1320 (N_1320,N_1260,N_1271);
xor U1321 (N_1321,N_1250,N_1275);
and U1322 (N_1322,N_1269,N_1251);
nor U1323 (N_1323,N_1273,N_1274);
and U1324 (N_1324,N_1264,N_1288);
xor U1325 (N_1325,N_1256,N_1258);
and U1326 (N_1326,N_1250,N_1274);
xnor U1327 (N_1327,N_1274,N_1277);
nand U1328 (N_1328,N_1268,N_1285);
and U1329 (N_1329,N_1285,N_1273);
nor U1330 (N_1330,N_1252,N_1269);
and U1331 (N_1331,N_1280,N_1270);
nor U1332 (N_1332,N_1251,N_1277);
xor U1333 (N_1333,N_1270,N_1285);
or U1334 (N_1334,N_1264,N_1296);
or U1335 (N_1335,N_1292,N_1285);
nand U1336 (N_1336,N_1263,N_1268);
or U1337 (N_1337,N_1279,N_1282);
nand U1338 (N_1338,N_1297,N_1290);
xor U1339 (N_1339,N_1257,N_1286);
and U1340 (N_1340,N_1266,N_1292);
or U1341 (N_1341,N_1292,N_1274);
nor U1342 (N_1342,N_1262,N_1276);
or U1343 (N_1343,N_1253,N_1287);
xor U1344 (N_1344,N_1293,N_1274);
and U1345 (N_1345,N_1288,N_1291);
nand U1346 (N_1346,N_1256,N_1254);
nor U1347 (N_1347,N_1290,N_1280);
xnor U1348 (N_1348,N_1272,N_1285);
nand U1349 (N_1349,N_1266,N_1289);
nand U1350 (N_1350,N_1338,N_1312);
or U1351 (N_1351,N_1343,N_1347);
or U1352 (N_1352,N_1321,N_1327);
xor U1353 (N_1353,N_1335,N_1313);
and U1354 (N_1354,N_1341,N_1305);
xnor U1355 (N_1355,N_1345,N_1346);
or U1356 (N_1356,N_1334,N_1331);
and U1357 (N_1357,N_1307,N_1337);
xnor U1358 (N_1358,N_1332,N_1309);
and U1359 (N_1359,N_1310,N_1315);
xnor U1360 (N_1360,N_1328,N_1317);
or U1361 (N_1361,N_1318,N_1336);
nand U1362 (N_1362,N_1340,N_1304);
nor U1363 (N_1363,N_1323,N_1329);
and U1364 (N_1364,N_1314,N_1306);
nor U1365 (N_1365,N_1348,N_1330);
or U1366 (N_1366,N_1311,N_1333);
or U1367 (N_1367,N_1301,N_1342);
xor U1368 (N_1368,N_1349,N_1319);
and U1369 (N_1369,N_1324,N_1302);
xor U1370 (N_1370,N_1316,N_1325);
and U1371 (N_1371,N_1320,N_1322);
or U1372 (N_1372,N_1300,N_1339);
nor U1373 (N_1373,N_1344,N_1326);
xnor U1374 (N_1374,N_1303,N_1308);
nor U1375 (N_1375,N_1322,N_1323);
and U1376 (N_1376,N_1324,N_1322);
or U1377 (N_1377,N_1329,N_1324);
or U1378 (N_1378,N_1308,N_1325);
nand U1379 (N_1379,N_1307,N_1303);
nor U1380 (N_1380,N_1326,N_1320);
or U1381 (N_1381,N_1347,N_1329);
or U1382 (N_1382,N_1328,N_1345);
nor U1383 (N_1383,N_1307,N_1333);
xnor U1384 (N_1384,N_1331,N_1328);
or U1385 (N_1385,N_1330,N_1326);
nor U1386 (N_1386,N_1308,N_1332);
nand U1387 (N_1387,N_1314,N_1329);
nor U1388 (N_1388,N_1326,N_1305);
xnor U1389 (N_1389,N_1346,N_1325);
and U1390 (N_1390,N_1331,N_1336);
nand U1391 (N_1391,N_1300,N_1305);
xor U1392 (N_1392,N_1332,N_1307);
nand U1393 (N_1393,N_1306,N_1331);
nand U1394 (N_1394,N_1328,N_1338);
or U1395 (N_1395,N_1306,N_1304);
xnor U1396 (N_1396,N_1306,N_1348);
and U1397 (N_1397,N_1324,N_1335);
and U1398 (N_1398,N_1313,N_1348);
and U1399 (N_1399,N_1318,N_1319);
nor U1400 (N_1400,N_1398,N_1369);
xor U1401 (N_1401,N_1352,N_1360);
nand U1402 (N_1402,N_1351,N_1386);
and U1403 (N_1403,N_1359,N_1374);
nand U1404 (N_1404,N_1370,N_1378);
nor U1405 (N_1405,N_1399,N_1373);
or U1406 (N_1406,N_1364,N_1387);
nand U1407 (N_1407,N_1354,N_1397);
and U1408 (N_1408,N_1372,N_1389);
nor U1409 (N_1409,N_1358,N_1366);
and U1410 (N_1410,N_1383,N_1391);
nor U1411 (N_1411,N_1356,N_1367);
or U1412 (N_1412,N_1394,N_1368);
nor U1413 (N_1413,N_1382,N_1392);
nand U1414 (N_1414,N_1362,N_1355);
nor U1415 (N_1415,N_1396,N_1371);
or U1416 (N_1416,N_1390,N_1375);
nor U1417 (N_1417,N_1361,N_1357);
or U1418 (N_1418,N_1376,N_1377);
and U1419 (N_1419,N_1380,N_1350);
and U1420 (N_1420,N_1379,N_1393);
and U1421 (N_1421,N_1353,N_1381);
xnor U1422 (N_1422,N_1363,N_1395);
nand U1423 (N_1423,N_1365,N_1385);
nor U1424 (N_1424,N_1388,N_1384);
nor U1425 (N_1425,N_1376,N_1359);
and U1426 (N_1426,N_1388,N_1355);
xor U1427 (N_1427,N_1361,N_1399);
xor U1428 (N_1428,N_1373,N_1388);
xor U1429 (N_1429,N_1354,N_1355);
and U1430 (N_1430,N_1361,N_1381);
or U1431 (N_1431,N_1368,N_1355);
or U1432 (N_1432,N_1377,N_1396);
xor U1433 (N_1433,N_1399,N_1365);
xor U1434 (N_1434,N_1358,N_1379);
nor U1435 (N_1435,N_1378,N_1362);
and U1436 (N_1436,N_1357,N_1351);
or U1437 (N_1437,N_1396,N_1394);
or U1438 (N_1438,N_1383,N_1362);
or U1439 (N_1439,N_1351,N_1395);
and U1440 (N_1440,N_1361,N_1389);
or U1441 (N_1441,N_1399,N_1378);
nor U1442 (N_1442,N_1391,N_1384);
nand U1443 (N_1443,N_1371,N_1386);
and U1444 (N_1444,N_1370,N_1366);
nor U1445 (N_1445,N_1372,N_1377);
or U1446 (N_1446,N_1369,N_1391);
xnor U1447 (N_1447,N_1391,N_1364);
nand U1448 (N_1448,N_1361,N_1377);
xnor U1449 (N_1449,N_1351,N_1363);
xnor U1450 (N_1450,N_1440,N_1446);
and U1451 (N_1451,N_1445,N_1420);
nand U1452 (N_1452,N_1427,N_1403);
and U1453 (N_1453,N_1400,N_1449);
or U1454 (N_1454,N_1439,N_1441);
or U1455 (N_1455,N_1435,N_1434);
and U1456 (N_1456,N_1417,N_1405);
nor U1457 (N_1457,N_1415,N_1423);
xor U1458 (N_1458,N_1424,N_1443);
or U1459 (N_1459,N_1407,N_1419);
nand U1460 (N_1460,N_1425,N_1404);
xnor U1461 (N_1461,N_1401,N_1448);
or U1462 (N_1462,N_1428,N_1431);
and U1463 (N_1463,N_1421,N_1408);
nand U1464 (N_1464,N_1422,N_1444);
nor U1465 (N_1465,N_1433,N_1411);
nand U1466 (N_1466,N_1414,N_1413);
nor U1467 (N_1467,N_1406,N_1436);
nor U1468 (N_1468,N_1437,N_1442);
nand U1469 (N_1469,N_1402,N_1438);
nor U1470 (N_1470,N_1429,N_1416);
nor U1471 (N_1471,N_1432,N_1412);
or U1472 (N_1472,N_1447,N_1409);
or U1473 (N_1473,N_1426,N_1430);
and U1474 (N_1474,N_1418,N_1410);
xor U1475 (N_1475,N_1408,N_1404);
and U1476 (N_1476,N_1429,N_1417);
nor U1477 (N_1477,N_1408,N_1415);
xor U1478 (N_1478,N_1409,N_1400);
or U1479 (N_1479,N_1428,N_1439);
nand U1480 (N_1480,N_1432,N_1419);
nand U1481 (N_1481,N_1424,N_1431);
or U1482 (N_1482,N_1443,N_1404);
xor U1483 (N_1483,N_1439,N_1419);
or U1484 (N_1484,N_1442,N_1407);
nand U1485 (N_1485,N_1416,N_1446);
nor U1486 (N_1486,N_1434,N_1414);
xnor U1487 (N_1487,N_1442,N_1426);
xnor U1488 (N_1488,N_1418,N_1432);
xor U1489 (N_1489,N_1441,N_1444);
xor U1490 (N_1490,N_1429,N_1442);
xor U1491 (N_1491,N_1427,N_1444);
nand U1492 (N_1492,N_1427,N_1441);
nand U1493 (N_1493,N_1432,N_1438);
and U1494 (N_1494,N_1403,N_1436);
nand U1495 (N_1495,N_1421,N_1424);
nor U1496 (N_1496,N_1406,N_1425);
xor U1497 (N_1497,N_1408,N_1423);
and U1498 (N_1498,N_1431,N_1445);
nand U1499 (N_1499,N_1438,N_1431);
xor U1500 (N_1500,N_1476,N_1462);
or U1501 (N_1501,N_1479,N_1468);
nor U1502 (N_1502,N_1460,N_1493);
nor U1503 (N_1503,N_1474,N_1475);
or U1504 (N_1504,N_1488,N_1465);
nor U1505 (N_1505,N_1470,N_1489);
nand U1506 (N_1506,N_1452,N_1458);
xnor U1507 (N_1507,N_1497,N_1469);
or U1508 (N_1508,N_1492,N_1454);
xor U1509 (N_1509,N_1451,N_1498);
xnor U1510 (N_1510,N_1459,N_1486);
nor U1511 (N_1511,N_1463,N_1487);
nor U1512 (N_1512,N_1483,N_1467);
nor U1513 (N_1513,N_1464,N_1499);
xor U1514 (N_1514,N_1485,N_1490);
nor U1515 (N_1515,N_1480,N_1478);
or U1516 (N_1516,N_1461,N_1481);
nor U1517 (N_1517,N_1457,N_1491);
nor U1518 (N_1518,N_1472,N_1471);
nor U1519 (N_1519,N_1453,N_1484);
nor U1520 (N_1520,N_1494,N_1466);
or U1521 (N_1521,N_1450,N_1455);
and U1522 (N_1522,N_1482,N_1496);
and U1523 (N_1523,N_1495,N_1473);
nand U1524 (N_1524,N_1477,N_1456);
or U1525 (N_1525,N_1480,N_1465);
or U1526 (N_1526,N_1466,N_1482);
nand U1527 (N_1527,N_1465,N_1499);
nand U1528 (N_1528,N_1465,N_1463);
and U1529 (N_1529,N_1477,N_1463);
xnor U1530 (N_1530,N_1451,N_1454);
or U1531 (N_1531,N_1493,N_1489);
or U1532 (N_1532,N_1473,N_1469);
nor U1533 (N_1533,N_1487,N_1476);
nand U1534 (N_1534,N_1456,N_1459);
xnor U1535 (N_1535,N_1496,N_1464);
and U1536 (N_1536,N_1493,N_1481);
or U1537 (N_1537,N_1472,N_1452);
or U1538 (N_1538,N_1498,N_1471);
xor U1539 (N_1539,N_1496,N_1466);
xor U1540 (N_1540,N_1464,N_1458);
and U1541 (N_1541,N_1466,N_1452);
xor U1542 (N_1542,N_1457,N_1463);
nor U1543 (N_1543,N_1462,N_1479);
and U1544 (N_1544,N_1483,N_1462);
or U1545 (N_1545,N_1458,N_1487);
and U1546 (N_1546,N_1467,N_1498);
nand U1547 (N_1547,N_1458,N_1455);
nor U1548 (N_1548,N_1476,N_1488);
xnor U1549 (N_1549,N_1462,N_1457);
and U1550 (N_1550,N_1510,N_1530);
and U1551 (N_1551,N_1528,N_1514);
nor U1552 (N_1552,N_1521,N_1520);
xnor U1553 (N_1553,N_1546,N_1541);
nand U1554 (N_1554,N_1517,N_1544);
xor U1555 (N_1555,N_1522,N_1545);
nor U1556 (N_1556,N_1509,N_1540);
or U1557 (N_1557,N_1529,N_1536);
and U1558 (N_1558,N_1548,N_1523);
nor U1559 (N_1559,N_1501,N_1527);
nand U1560 (N_1560,N_1519,N_1502);
nor U1561 (N_1561,N_1518,N_1539);
xor U1562 (N_1562,N_1512,N_1538);
and U1563 (N_1563,N_1533,N_1531);
or U1564 (N_1564,N_1513,N_1535);
or U1565 (N_1565,N_1543,N_1505);
nor U1566 (N_1566,N_1524,N_1504);
and U1567 (N_1567,N_1503,N_1515);
nor U1568 (N_1568,N_1525,N_1542);
or U1569 (N_1569,N_1537,N_1507);
and U1570 (N_1570,N_1532,N_1549);
xor U1571 (N_1571,N_1508,N_1534);
nor U1572 (N_1572,N_1500,N_1506);
xnor U1573 (N_1573,N_1516,N_1526);
nand U1574 (N_1574,N_1511,N_1547);
nand U1575 (N_1575,N_1507,N_1543);
or U1576 (N_1576,N_1525,N_1543);
xor U1577 (N_1577,N_1534,N_1503);
nor U1578 (N_1578,N_1521,N_1514);
nor U1579 (N_1579,N_1519,N_1540);
or U1580 (N_1580,N_1540,N_1545);
nor U1581 (N_1581,N_1515,N_1510);
or U1582 (N_1582,N_1516,N_1519);
and U1583 (N_1583,N_1549,N_1533);
nor U1584 (N_1584,N_1534,N_1527);
or U1585 (N_1585,N_1549,N_1509);
nand U1586 (N_1586,N_1547,N_1527);
xor U1587 (N_1587,N_1544,N_1533);
nand U1588 (N_1588,N_1525,N_1532);
nand U1589 (N_1589,N_1547,N_1524);
nand U1590 (N_1590,N_1547,N_1548);
and U1591 (N_1591,N_1547,N_1514);
or U1592 (N_1592,N_1542,N_1514);
or U1593 (N_1593,N_1544,N_1509);
nand U1594 (N_1594,N_1512,N_1531);
or U1595 (N_1595,N_1527,N_1518);
and U1596 (N_1596,N_1534,N_1517);
nor U1597 (N_1597,N_1536,N_1539);
xor U1598 (N_1598,N_1548,N_1549);
or U1599 (N_1599,N_1506,N_1531);
or U1600 (N_1600,N_1566,N_1583);
nand U1601 (N_1601,N_1554,N_1596);
nor U1602 (N_1602,N_1559,N_1565);
and U1603 (N_1603,N_1581,N_1589);
or U1604 (N_1604,N_1571,N_1569);
or U1605 (N_1605,N_1579,N_1597);
or U1606 (N_1606,N_1560,N_1578);
and U1607 (N_1607,N_1555,N_1592);
or U1608 (N_1608,N_1550,N_1598);
nand U1609 (N_1609,N_1572,N_1568);
xnor U1610 (N_1610,N_1599,N_1576);
xnor U1611 (N_1611,N_1593,N_1558);
nand U1612 (N_1612,N_1595,N_1574);
nand U1613 (N_1613,N_1594,N_1573);
xnor U1614 (N_1614,N_1587,N_1588);
xor U1615 (N_1615,N_1575,N_1590);
or U1616 (N_1616,N_1584,N_1556);
or U1617 (N_1617,N_1567,N_1563);
or U1618 (N_1618,N_1577,N_1562);
xor U1619 (N_1619,N_1586,N_1557);
nor U1620 (N_1620,N_1553,N_1585);
or U1621 (N_1621,N_1591,N_1551);
nor U1622 (N_1622,N_1564,N_1582);
nor U1623 (N_1623,N_1561,N_1570);
and U1624 (N_1624,N_1580,N_1552);
xnor U1625 (N_1625,N_1567,N_1578);
xnor U1626 (N_1626,N_1569,N_1575);
and U1627 (N_1627,N_1573,N_1583);
or U1628 (N_1628,N_1559,N_1596);
or U1629 (N_1629,N_1593,N_1595);
nor U1630 (N_1630,N_1586,N_1569);
nor U1631 (N_1631,N_1551,N_1582);
nor U1632 (N_1632,N_1588,N_1562);
xnor U1633 (N_1633,N_1576,N_1580);
nor U1634 (N_1634,N_1592,N_1582);
xnor U1635 (N_1635,N_1580,N_1562);
and U1636 (N_1636,N_1557,N_1577);
nand U1637 (N_1637,N_1595,N_1570);
nor U1638 (N_1638,N_1551,N_1552);
nor U1639 (N_1639,N_1559,N_1560);
nand U1640 (N_1640,N_1580,N_1558);
xor U1641 (N_1641,N_1578,N_1572);
nand U1642 (N_1642,N_1579,N_1561);
and U1643 (N_1643,N_1591,N_1590);
xor U1644 (N_1644,N_1560,N_1585);
or U1645 (N_1645,N_1561,N_1595);
nand U1646 (N_1646,N_1563,N_1566);
nor U1647 (N_1647,N_1591,N_1598);
nand U1648 (N_1648,N_1594,N_1592);
and U1649 (N_1649,N_1597,N_1594);
or U1650 (N_1650,N_1623,N_1614);
nor U1651 (N_1651,N_1606,N_1625);
xnor U1652 (N_1652,N_1602,N_1607);
or U1653 (N_1653,N_1646,N_1643);
nor U1654 (N_1654,N_1638,N_1619);
or U1655 (N_1655,N_1605,N_1627);
and U1656 (N_1656,N_1620,N_1629);
xor U1657 (N_1657,N_1648,N_1610);
or U1658 (N_1658,N_1616,N_1631);
xnor U1659 (N_1659,N_1647,N_1642);
nor U1660 (N_1660,N_1644,N_1608);
xnor U1661 (N_1661,N_1601,N_1626);
nor U1662 (N_1662,N_1604,N_1612);
xor U1663 (N_1663,N_1618,N_1649);
nand U1664 (N_1664,N_1632,N_1637);
and U1665 (N_1665,N_1634,N_1636);
nor U1666 (N_1666,N_1635,N_1621);
and U1667 (N_1667,N_1624,N_1630);
xor U1668 (N_1668,N_1639,N_1617);
nor U1669 (N_1669,N_1609,N_1622);
xor U1670 (N_1670,N_1640,N_1633);
and U1671 (N_1671,N_1611,N_1628);
xnor U1672 (N_1672,N_1600,N_1613);
and U1673 (N_1673,N_1641,N_1645);
nand U1674 (N_1674,N_1603,N_1615);
or U1675 (N_1675,N_1640,N_1645);
and U1676 (N_1676,N_1643,N_1615);
or U1677 (N_1677,N_1623,N_1632);
nor U1678 (N_1678,N_1622,N_1635);
nor U1679 (N_1679,N_1600,N_1627);
and U1680 (N_1680,N_1618,N_1605);
nand U1681 (N_1681,N_1639,N_1648);
nand U1682 (N_1682,N_1638,N_1605);
xor U1683 (N_1683,N_1633,N_1644);
and U1684 (N_1684,N_1618,N_1636);
nand U1685 (N_1685,N_1631,N_1629);
and U1686 (N_1686,N_1629,N_1630);
nor U1687 (N_1687,N_1647,N_1628);
nor U1688 (N_1688,N_1609,N_1644);
nor U1689 (N_1689,N_1640,N_1630);
and U1690 (N_1690,N_1636,N_1625);
nor U1691 (N_1691,N_1630,N_1649);
nor U1692 (N_1692,N_1640,N_1616);
and U1693 (N_1693,N_1640,N_1636);
and U1694 (N_1694,N_1646,N_1601);
nor U1695 (N_1695,N_1640,N_1607);
and U1696 (N_1696,N_1643,N_1608);
nor U1697 (N_1697,N_1617,N_1630);
nand U1698 (N_1698,N_1641,N_1648);
or U1699 (N_1699,N_1623,N_1634);
or U1700 (N_1700,N_1697,N_1664);
nor U1701 (N_1701,N_1681,N_1670);
nand U1702 (N_1702,N_1696,N_1673);
nand U1703 (N_1703,N_1655,N_1684);
and U1704 (N_1704,N_1687,N_1667);
xor U1705 (N_1705,N_1686,N_1698);
nor U1706 (N_1706,N_1660,N_1683);
or U1707 (N_1707,N_1662,N_1663);
and U1708 (N_1708,N_1651,N_1679);
or U1709 (N_1709,N_1650,N_1676);
nand U1710 (N_1710,N_1672,N_1661);
or U1711 (N_1711,N_1685,N_1654);
nor U1712 (N_1712,N_1653,N_1671);
nor U1713 (N_1713,N_1652,N_1674);
nor U1714 (N_1714,N_1665,N_1668);
nand U1715 (N_1715,N_1692,N_1689);
or U1716 (N_1716,N_1694,N_1680);
and U1717 (N_1717,N_1691,N_1677);
nor U1718 (N_1718,N_1666,N_1657);
nand U1719 (N_1719,N_1695,N_1659);
nand U1720 (N_1720,N_1699,N_1658);
nor U1721 (N_1721,N_1688,N_1678);
nor U1722 (N_1722,N_1656,N_1669);
or U1723 (N_1723,N_1690,N_1693);
and U1724 (N_1724,N_1682,N_1675);
nand U1725 (N_1725,N_1668,N_1691);
nand U1726 (N_1726,N_1653,N_1685);
or U1727 (N_1727,N_1665,N_1653);
nor U1728 (N_1728,N_1663,N_1691);
and U1729 (N_1729,N_1683,N_1661);
or U1730 (N_1730,N_1696,N_1678);
nand U1731 (N_1731,N_1658,N_1698);
nor U1732 (N_1732,N_1685,N_1698);
xor U1733 (N_1733,N_1670,N_1678);
xor U1734 (N_1734,N_1650,N_1684);
nor U1735 (N_1735,N_1656,N_1655);
nand U1736 (N_1736,N_1655,N_1682);
nand U1737 (N_1737,N_1651,N_1695);
xnor U1738 (N_1738,N_1659,N_1667);
nor U1739 (N_1739,N_1674,N_1675);
or U1740 (N_1740,N_1676,N_1678);
nor U1741 (N_1741,N_1674,N_1655);
nand U1742 (N_1742,N_1666,N_1685);
nor U1743 (N_1743,N_1688,N_1686);
xnor U1744 (N_1744,N_1679,N_1694);
nand U1745 (N_1745,N_1672,N_1687);
xor U1746 (N_1746,N_1677,N_1655);
xor U1747 (N_1747,N_1662,N_1658);
nand U1748 (N_1748,N_1673,N_1694);
nand U1749 (N_1749,N_1689,N_1658);
and U1750 (N_1750,N_1733,N_1718);
xnor U1751 (N_1751,N_1716,N_1705);
and U1752 (N_1752,N_1709,N_1746);
or U1753 (N_1753,N_1744,N_1725);
nand U1754 (N_1754,N_1743,N_1714);
xor U1755 (N_1755,N_1708,N_1735);
or U1756 (N_1756,N_1707,N_1749);
nand U1757 (N_1757,N_1702,N_1711);
nand U1758 (N_1758,N_1739,N_1738);
nand U1759 (N_1759,N_1745,N_1713);
xnor U1760 (N_1760,N_1701,N_1730);
or U1761 (N_1761,N_1715,N_1727);
or U1762 (N_1762,N_1720,N_1726);
xnor U1763 (N_1763,N_1721,N_1747);
xnor U1764 (N_1764,N_1724,N_1742);
nor U1765 (N_1765,N_1700,N_1740);
or U1766 (N_1766,N_1706,N_1736);
xnor U1767 (N_1767,N_1703,N_1728);
xnor U1768 (N_1768,N_1741,N_1737);
xnor U1769 (N_1769,N_1732,N_1723);
or U1770 (N_1770,N_1710,N_1729);
xnor U1771 (N_1771,N_1734,N_1717);
or U1772 (N_1772,N_1731,N_1719);
and U1773 (N_1773,N_1712,N_1704);
or U1774 (N_1774,N_1748,N_1722);
nor U1775 (N_1775,N_1717,N_1700);
and U1776 (N_1776,N_1707,N_1722);
nand U1777 (N_1777,N_1707,N_1720);
xnor U1778 (N_1778,N_1734,N_1732);
nor U1779 (N_1779,N_1739,N_1723);
nand U1780 (N_1780,N_1710,N_1715);
nor U1781 (N_1781,N_1701,N_1719);
nand U1782 (N_1782,N_1712,N_1724);
nor U1783 (N_1783,N_1731,N_1718);
or U1784 (N_1784,N_1731,N_1743);
or U1785 (N_1785,N_1743,N_1732);
nor U1786 (N_1786,N_1722,N_1724);
nand U1787 (N_1787,N_1708,N_1739);
nor U1788 (N_1788,N_1731,N_1705);
nor U1789 (N_1789,N_1701,N_1729);
nor U1790 (N_1790,N_1711,N_1722);
or U1791 (N_1791,N_1748,N_1726);
or U1792 (N_1792,N_1749,N_1720);
and U1793 (N_1793,N_1724,N_1730);
nor U1794 (N_1794,N_1727,N_1719);
nor U1795 (N_1795,N_1720,N_1721);
and U1796 (N_1796,N_1716,N_1717);
nor U1797 (N_1797,N_1721,N_1714);
xor U1798 (N_1798,N_1737,N_1702);
nand U1799 (N_1799,N_1732,N_1702);
xnor U1800 (N_1800,N_1780,N_1792);
nor U1801 (N_1801,N_1791,N_1777);
or U1802 (N_1802,N_1754,N_1783);
and U1803 (N_1803,N_1752,N_1750);
and U1804 (N_1804,N_1790,N_1781);
nand U1805 (N_1805,N_1789,N_1765);
nand U1806 (N_1806,N_1766,N_1753);
nor U1807 (N_1807,N_1776,N_1755);
and U1808 (N_1808,N_1772,N_1771);
or U1809 (N_1809,N_1759,N_1785);
nor U1810 (N_1810,N_1795,N_1793);
nor U1811 (N_1811,N_1775,N_1784);
nor U1812 (N_1812,N_1762,N_1769);
and U1813 (N_1813,N_1782,N_1767);
and U1814 (N_1814,N_1751,N_1758);
xor U1815 (N_1815,N_1773,N_1768);
or U1816 (N_1816,N_1797,N_1761);
nand U1817 (N_1817,N_1799,N_1779);
or U1818 (N_1818,N_1770,N_1757);
or U1819 (N_1819,N_1778,N_1788);
xor U1820 (N_1820,N_1798,N_1786);
or U1821 (N_1821,N_1796,N_1763);
nor U1822 (N_1822,N_1764,N_1760);
nor U1823 (N_1823,N_1787,N_1756);
nand U1824 (N_1824,N_1794,N_1774);
nor U1825 (N_1825,N_1773,N_1780);
and U1826 (N_1826,N_1755,N_1773);
xor U1827 (N_1827,N_1784,N_1778);
xor U1828 (N_1828,N_1753,N_1792);
and U1829 (N_1829,N_1769,N_1768);
and U1830 (N_1830,N_1774,N_1754);
nand U1831 (N_1831,N_1799,N_1763);
xnor U1832 (N_1832,N_1756,N_1751);
nor U1833 (N_1833,N_1768,N_1762);
xor U1834 (N_1834,N_1758,N_1784);
nand U1835 (N_1835,N_1768,N_1797);
nor U1836 (N_1836,N_1784,N_1756);
or U1837 (N_1837,N_1798,N_1760);
xnor U1838 (N_1838,N_1790,N_1795);
nor U1839 (N_1839,N_1788,N_1775);
nor U1840 (N_1840,N_1786,N_1781);
nand U1841 (N_1841,N_1786,N_1771);
and U1842 (N_1842,N_1792,N_1760);
nor U1843 (N_1843,N_1750,N_1755);
nand U1844 (N_1844,N_1798,N_1779);
nor U1845 (N_1845,N_1756,N_1776);
xnor U1846 (N_1846,N_1791,N_1796);
nand U1847 (N_1847,N_1776,N_1764);
xor U1848 (N_1848,N_1799,N_1760);
or U1849 (N_1849,N_1760,N_1756);
nor U1850 (N_1850,N_1823,N_1828);
nor U1851 (N_1851,N_1801,N_1802);
nor U1852 (N_1852,N_1837,N_1836);
nor U1853 (N_1853,N_1808,N_1844);
nand U1854 (N_1854,N_1835,N_1831);
or U1855 (N_1855,N_1834,N_1820);
or U1856 (N_1856,N_1805,N_1811);
or U1857 (N_1857,N_1814,N_1848);
nor U1858 (N_1858,N_1839,N_1847);
or U1859 (N_1859,N_1809,N_1812);
and U1860 (N_1860,N_1818,N_1819);
xnor U1861 (N_1861,N_1842,N_1813);
or U1862 (N_1862,N_1832,N_1817);
or U1863 (N_1863,N_1810,N_1843);
xnor U1864 (N_1864,N_1833,N_1845);
xnor U1865 (N_1865,N_1846,N_1821);
xor U1866 (N_1866,N_1830,N_1826);
nor U1867 (N_1867,N_1849,N_1807);
nand U1868 (N_1868,N_1841,N_1815);
nand U1869 (N_1869,N_1816,N_1824);
nor U1870 (N_1870,N_1800,N_1827);
and U1871 (N_1871,N_1804,N_1838);
and U1872 (N_1872,N_1840,N_1829);
or U1873 (N_1873,N_1803,N_1825);
or U1874 (N_1874,N_1822,N_1806);
and U1875 (N_1875,N_1833,N_1820);
or U1876 (N_1876,N_1807,N_1836);
nand U1877 (N_1877,N_1836,N_1833);
xnor U1878 (N_1878,N_1812,N_1831);
xnor U1879 (N_1879,N_1812,N_1840);
nor U1880 (N_1880,N_1812,N_1801);
nor U1881 (N_1881,N_1828,N_1811);
or U1882 (N_1882,N_1816,N_1838);
nor U1883 (N_1883,N_1844,N_1821);
or U1884 (N_1884,N_1806,N_1823);
and U1885 (N_1885,N_1846,N_1829);
nor U1886 (N_1886,N_1840,N_1825);
nor U1887 (N_1887,N_1841,N_1807);
or U1888 (N_1888,N_1810,N_1802);
or U1889 (N_1889,N_1823,N_1821);
nor U1890 (N_1890,N_1816,N_1829);
or U1891 (N_1891,N_1802,N_1846);
xnor U1892 (N_1892,N_1844,N_1816);
and U1893 (N_1893,N_1808,N_1814);
and U1894 (N_1894,N_1818,N_1844);
or U1895 (N_1895,N_1815,N_1808);
nor U1896 (N_1896,N_1820,N_1835);
nor U1897 (N_1897,N_1831,N_1846);
xor U1898 (N_1898,N_1810,N_1800);
and U1899 (N_1899,N_1824,N_1841);
nor U1900 (N_1900,N_1869,N_1857);
and U1901 (N_1901,N_1875,N_1864);
or U1902 (N_1902,N_1880,N_1887);
xor U1903 (N_1903,N_1893,N_1899);
xor U1904 (N_1904,N_1872,N_1876);
and U1905 (N_1905,N_1854,N_1895);
nand U1906 (N_1906,N_1858,N_1860);
and U1907 (N_1907,N_1891,N_1881);
and U1908 (N_1908,N_1850,N_1863);
nor U1909 (N_1909,N_1878,N_1861);
or U1910 (N_1910,N_1883,N_1884);
nand U1911 (N_1911,N_1885,N_1886);
or U1912 (N_1912,N_1877,N_1853);
or U1913 (N_1913,N_1874,N_1871);
nand U1914 (N_1914,N_1894,N_1898);
and U1915 (N_1915,N_1892,N_1867);
or U1916 (N_1916,N_1866,N_1879);
nand U1917 (N_1917,N_1851,N_1855);
xor U1918 (N_1918,N_1888,N_1896);
nor U1919 (N_1919,N_1859,N_1889);
xor U1920 (N_1920,N_1890,N_1852);
nor U1921 (N_1921,N_1870,N_1865);
or U1922 (N_1922,N_1868,N_1882);
and U1923 (N_1923,N_1862,N_1873);
or U1924 (N_1924,N_1897,N_1856);
xnor U1925 (N_1925,N_1850,N_1884);
nand U1926 (N_1926,N_1855,N_1861);
xnor U1927 (N_1927,N_1852,N_1875);
and U1928 (N_1928,N_1882,N_1898);
and U1929 (N_1929,N_1870,N_1897);
nand U1930 (N_1930,N_1882,N_1884);
or U1931 (N_1931,N_1866,N_1873);
nand U1932 (N_1932,N_1855,N_1870);
and U1933 (N_1933,N_1896,N_1882);
or U1934 (N_1934,N_1851,N_1861);
or U1935 (N_1935,N_1878,N_1851);
and U1936 (N_1936,N_1872,N_1897);
xnor U1937 (N_1937,N_1869,N_1880);
nor U1938 (N_1938,N_1891,N_1868);
nand U1939 (N_1939,N_1879,N_1877);
nor U1940 (N_1940,N_1892,N_1871);
and U1941 (N_1941,N_1893,N_1873);
nor U1942 (N_1942,N_1865,N_1866);
nor U1943 (N_1943,N_1855,N_1899);
nor U1944 (N_1944,N_1859,N_1882);
nand U1945 (N_1945,N_1896,N_1850);
xnor U1946 (N_1946,N_1851,N_1866);
and U1947 (N_1947,N_1865,N_1880);
nor U1948 (N_1948,N_1855,N_1856);
and U1949 (N_1949,N_1893,N_1860);
and U1950 (N_1950,N_1935,N_1937);
xnor U1951 (N_1951,N_1929,N_1938);
and U1952 (N_1952,N_1924,N_1948);
xor U1953 (N_1953,N_1916,N_1946);
nand U1954 (N_1954,N_1903,N_1902);
nand U1955 (N_1955,N_1945,N_1904);
nor U1956 (N_1956,N_1905,N_1914);
xnor U1957 (N_1957,N_1931,N_1910);
xnor U1958 (N_1958,N_1934,N_1930);
and U1959 (N_1959,N_1920,N_1927);
nor U1960 (N_1960,N_1928,N_1909);
and U1961 (N_1961,N_1944,N_1923);
and U1962 (N_1962,N_1925,N_1918);
and U1963 (N_1963,N_1939,N_1943);
nand U1964 (N_1964,N_1917,N_1932);
nor U1965 (N_1965,N_1913,N_1911);
or U1966 (N_1966,N_1926,N_1906);
or U1967 (N_1967,N_1942,N_1907);
xnor U1968 (N_1968,N_1933,N_1941);
nand U1969 (N_1969,N_1940,N_1901);
nor U1970 (N_1970,N_1912,N_1915);
and U1971 (N_1971,N_1947,N_1900);
and U1972 (N_1972,N_1908,N_1921);
or U1973 (N_1973,N_1919,N_1949);
or U1974 (N_1974,N_1922,N_1936);
nand U1975 (N_1975,N_1917,N_1946);
xnor U1976 (N_1976,N_1931,N_1942);
nor U1977 (N_1977,N_1909,N_1939);
or U1978 (N_1978,N_1944,N_1939);
nor U1979 (N_1979,N_1918,N_1917);
xor U1980 (N_1980,N_1919,N_1905);
or U1981 (N_1981,N_1904,N_1929);
xor U1982 (N_1982,N_1901,N_1903);
xnor U1983 (N_1983,N_1935,N_1905);
and U1984 (N_1984,N_1901,N_1904);
or U1985 (N_1985,N_1935,N_1933);
nor U1986 (N_1986,N_1940,N_1900);
or U1987 (N_1987,N_1943,N_1948);
or U1988 (N_1988,N_1911,N_1907);
and U1989 (N_1989,N_1932,N_1928);
or U1990 (N_1990,N_1910,N_1949);
xor U1991 (N_1991,N_1900,N_1946);
nand U1992 (N_1992,N_1931,N_1908);
nor U1993 (N_1993,N_1931,N_1935);
xor U1994 (N_1994,N_1928,N_1900);
nand U1995 (N_1995,N_1938,N_1945);
nor U1996 (N_1996,N_1947,N_1942);
xor U1997 (N_1997,N_1948,N_1936);
xor U1998 (N_1998,N_1917,N_1926);
nand U1999 (N_1999,N_1937,N_1927);
xnor U2000 (N_2000,N_1968,N_1979);
xnor U2001 (N_2001,N_1953,N_1963);
xor U2002 (N_2002,N_1996,N_1955);
and U2003 (N_2003,N_1998,N_1978);
nand U2004 (N_2004,N_1966,N_1991);
nand U2005 (N_2005,N_1990,N_1983);
xnor U2006 (N_2006,N_1962,N_1975);
xor U2007 (N_2007,N_1980,N_1997);
and U2008 (N_2008,N_1972,N_1977);
and U2009 (N_2009,N_1992,N_1965);
xnor U2010 (N_2010,N_1952,N_1951);
nor U2011 (N_2011,N_1989,N_1986);
nand U2012 (N_2012,N_1988,N_1957);
nand U2013 (N_2013,N_1987,N_1956);
nor U2014 (N_2014,N_1961,N_1981);
or U2015 (N_2015,N_1982,N_1954);
and U2016 (N_2016,N_1959,N_1993);
and U2017 (N_2017,N_1950,N_1973);
and U2018 (N_2018,N_1971,N_1967);
or U2019 (N_2019,N_1970,N_1974);
or U2020 (N_2020,N_1999,N_1964);
nor U2021 (N_2021,N_1985,N_1969);
or U2022 (N_2022,N_1958,N_1995);
xor U2023 (N_2023,N_1960,N_1994);
and U2024 (N_2024,N_1976,N_1984);
nand U2025 (N_2025,N_1995,N_1989);
and U2026 (N_2026,N_1962,N_1999);
and U2027 (N_2027,N_1982,N_1968);
xor U2028 (N_2028,N_1997,N_1966);
nand U2029 (N_2029,N_1962,N_1950);
or U2030 (N_2030,N_1995,N_1987);
nand U2031 (N_2031,N_1963,N_1987);
and U2032 (N_2032,N_1960,N_1973);
and U2033 (N_2033,N_1986,N_1961);
nand U2034 (N_2034,N_1968,N_1999);
xor U2035 (N_2035,N_1954,N_1986);
xnor U2036 (N_2036,N_1956,N_1961);
or U2037 (N_2037,N_1980,N_1985);
xor U2038 (N_2038,N_1958,N_1985);
nand U2039 (N_2039,N_1974,N_1992);
and U2040 (N_2040,N_1993,N_1964);
nand U2041 (N_2041,N_1989,N_1996);
or U2042 (N_2042,N_1958,N_1992);
nand U2043 (N_2043,N_1997,N_1953);
nor U2044 (N_2044,N_1953,N_1989);
nor U2045 (N_2045,N_1954,N_1956);
nor U2046 (N_2046,N_1950,N_1956);
and U2047 (N_2047,N_1983,N_1998);
or U2048 (N_2048,N_1950,N_1985);
and U2049 (N_2049,N_1992,N_1984);
and U2050 (N_2050,N_2032,N_2014);
xor U2051 (N_2051,N_2041,N_2043);
nor U2052 (N_2052,N_2017,N_2016);
nor U2053 (N_2053,N_2040,N_2013);
or U2054 (N_2054,N_2006,N_2024);
xnor U2055 (N_2055,N_2005,N_2046);
or U2056 (N_2056,N_2012,N_2007);
nor U2057 (N_2057,N_2033,N_2034);
and U2058 (N_2058,N_2027,N_2042);
nor U2059 (N_2059,N_2037,N_2023);
nor U2060 (N_2060,N_2047,N_2018);
xnor U2061 (N_2061,N_2029,N_2044);
xnor U2062 (N_2062,N_2035,N_2004);
nor U2063 (N_2063,N_2045,N_2021);
xnor U2064 (N_2064,N_2020,N_2011);
xnor U2065 (N_2065,N_2030,N_2001);
xor U2066 (N_2066,N_2049,N_2019);
nor U2067 (N_2067,N_2028,N_2022);
or U2068 (N_2068,N_2038,N_2000);
nor U2069 (N_2069,N_2039,N_2009);
xnor U2070 (N_2070,N_2002,N_2036);
xnor U2071 (N_2071,N_2003,N_2008);
nand U2072 (N_2072,N_2025,N_2031);
or U2073 (N_2073,N_2048,N_2015);
xor U2074 (N_2074,N_2026,N_2010);
nand U2075 (N_2075,N_2020,N_2003);
xor U2076 (N_2076,N_2037,N_2007);
xnor U2077 (N_2077,N_2016,N_2045);
xor U2078 (N_2078,N_2040,N_2037);
nand U2079 (N_2079,N_2029,N_2038);
xor U2080 (N_2080,N_2004,N_2045);
nand U2081 (N_2081,N_2004,N_2021);
nand U2082 (N_2082,N_2009,N_2003);
or U2083 (N_2083,N_2012,N_2024);
nand U2084 (N_2084,N_2008,N_2028);
or U2085 (N_2085,N_2044,N_2007);
nor U2086 (N_2086,N_2022,N_2008);
xnor U2087 (N_2087,N_2011,N_2016);
nand U2088 (N_2088,N_2018,N_2035);
and U2089 (N_2089,N_2008,N_2026);
xor U2090 (N_2090,N_2007,N_2021);
nor U2091 (N_2091,N_2033,N_2006);
nand U2092 (N_2092,N_2048,N_2003);
nor U2093 (N_2093,N_2038,N_2003);
nand U2094 (N_2094,N_2031,N_2009);
nand U2095 (N_2095,N_2023,N_2024);
and U2096 (N_2096,N_2043,N_2024);
or U2097 (N_2097,N_2039,N_2030);
nand U2098 (N_2098,N_2020,N_2046);
or U2099 (N_2099,N_2044,N_2033);
nor U2100 (N_2100,N_2050,N_2069);
nor U2101 (N_2101,N_2092,N_2079);
and U2102 (N_2102,N_2064,N_2076);
or U2103 (N_2103,N_2058,N_2089);
nor U2104 (N_2104,N_2096,N_2072);
nand U2105 (N_2105,N_2077,N_2057);
or U2106 (N_2106,N_2082,N_2071);
or U2107 (N_2107,N_2083,N_2098);
nand U2108 (N_2108,N_2051,N_2060);
and U2109 (N_2109,N_2081,N_2097);
or U2110 (N_2110,N_2090,N_2056);
and U2111 (N_2111,N_2087,N_2070);
xnor U2112 (N_2112,N_2088,N_2073);
nor U2113 (N_2113,N_2095,N_2094);
xnor U2114 (N_2114,N_2068,N_2075);
xor U2115 (N_2115,N_2093,N_2061);
nor U2116 (N_2116,N_2062,N_2084);
and U2117 (N_2117,N_2065,N_2052);
and U2118 (N_2118,N_2053,N_2085);
nand U2119 (N_2119,N_2078,N_2091);
nand U2120 (N_2120,N_2055,N_2067);
or U2121 (N_2121,N_2086,N_2054);
nor U2122 (N_2122,N_2063,N_2080);
nor U2123 (N_2123,N_2066,N_2059);
xnor U2124 (N_2124,N_2099,N_2074);
or U2125 (N_2125,N_2051,N_2093);
and U2126 (N_2126,N_2065,N_2076);
nand U2127 (N_2127,N_2083,N_2057);
nor U2128 (N_2128,N_2068,N_2095);
or U2129 (N_2129,N_2051,N_2077);
and U2130 (N_2130,N_2054,N_2098);
or U2131 (N_2131,N_2056,N_2098);
nand U2132 (N_2132,N_2069,N_2095);
xor U2133 (N_2133,N_2065,N_2084);
nor U2134 (N_2134,N_2073,N_2070);
nor U2135 (N_2135,N_2093,N_2060);
nand U2136 (N_2136,N_2080,N_2051);
nor U2137 (N_2137,N_2062,N_2051);
and U2138 (N_2138,N_2057,N_2052);
xor U2139 (N_2139,N_2059,N_2083);
and U2140 (N_2140,N_2068,N_2073);
xnor U2141 (N_2141,N_2073,N_2062);
and U2142 (N_2142,N_2077,N_2070);
xnor U2143 (N_2143,N_2099,N_2091);
xor U2144 (N_2144,N_2069,N_2079);
xnor U2145 (N_2145,N_2058,N_2088);
xnor U2146 (N_2146,N_2050,N_2054);
xnor U2147 (N_2147,N_2089,N_2078);
nand U2148 (N_2148,N_2065,N_2087);
xnor U2149 (N_2149,N_2092,N_2060);
and U2150 (N_2150,N_2119,N_2126);
or U2151 (N_2151,N_2105,N_2113);
nand U2152 (N_2152,N_2120,N_2124);
and U2153 (N_2153,N_2141,N_2115);
and U2154 (N_2154,N_2125,N_2136);
and U2155 (N_2155,N_2145,N_2122);
or U2156 (N_2156,N_2146,N_2108);
or U2157 (N_2157,N_2101,N_2111);
or U2158 (N_2158,N_2133,N_2127);
nor U2159 (N_2159,N_2109,N_2144);
xnor U2160 (N_2160,N_2102,N_2131);
xnor U2161 (N_2161,N_2142,N_2147);
xor U2162 (N_2162,N_2134,N_2132);
nor U2163 (N_2163,N_2138,N_2135);
or U2164 (N_2164,N_2103,N_2148);
xnor U2165 (N_2165,N_2117,N_2104);
or U2166 (N_2166,N_2121,N_2128);
and U2167 (N_2167,N_2130,N_2116);
or U2168 (N_2168,N_2137,N_2100);
xnor U2169 (N_2169,N_2123,N_2129);
xor U2170 (N_2170,N_2149,N_2110);
nand U2171 (N_2171,N_2112,N_2118);
nor U2172 (N_2172,N_2139,N_2140);
nor U2173 (N_2173,N_2107,N_2114);
xor U2174 (N_2174,N_2143,N_2106);
and U2175 (N_2175,N_2142,N_2129);
xnor U2176 (N_2176,N_2117,N_2141);
and U2177 (N_2177,N_2113,N_2142);
or U2178 (N_2178,N_2141,N_2113);
and U2179 (N_2179,N_2117,N_2122);
or U2180 (N_2180,N_2142,N_2106);
and U2181 (N_2181,N_2120,N_2140);
nand U2182 (N_2182,N_2101,N_2135);
or U2183 (N_2183,N_2134,N_2119);
and U2184 (N_2184,N_2129,N_2145);
and U2185 (N_2185,N_2138,N_2117);
and U2186 (N_2186,N_2121,N_2110);
xnor U2187 (N_2187,N_2113,N_2104);
or U2188 (N_2188,N_2134,N_2114);
nor U2189 (N_2189,N_2134,N_2147);
xnor U2190 (N_2190,N_2141,N_2108);
nor U2191 (N_2191,N_2111,N_2110);
xor U2192 (N_2192,N_2115,N_2118);
and U2193 (N_2193,N_2103,N_2137);
nor U2194 (N_2194,N_2101,N_2139);
nor U2195 (N_2195,N_2127,N_2138);
xor U2196 (N_2196,N_2113,N_2109);
or U2197 (N_2197,N_2143,N_2113);
and U2198 (N_2198,N_2111,N_2135);
and U2199 (N_2199,N_2146,N_2110);
or U2200 (N_2200,N_2184,N_2175);
nand U2201 (N_2201,N_2151,N_2179);
or U2202 (N_2202,N_2181,N_2190);
or U2203 (N_2203,N_2195,N_2160);
and U2204 (N_2204,N_2177,N_2188);
or U2205 (N_2205,N_2187,N_2162);
and U2206 (N_2206,N_2166,N_2168);
and U2207 (N_2207,N_2164,N_2173);
xnor U2208 (N_2208,N_2154,N_2197);
or U2209 (N_2209,N_2186,N_2153);
xor U2210 (N_2210,N_2159,N_2152);
nor U2211 (N_2211,N_2198,N_2171);
and U2212 (N_2212,N_2196,N_2150);
nand U2213 (N_2213,N_2157,N_2189);
or U2214 (N_2214,N_2155,N_2180);
or U2215 (N_2215,N_2169,N_2182);
or U2216 (N_2216,N_2176,N_2167);
or U2217 (N_2217,N_2194,N_2192);
xor U2218 (N_2218,N_2165,N_2178);
nand U2219 (N_2219,N_2156,N_2191);
or U2220 (N_2220,N_2199,N_2158);
or U2221 (N_2221,N_2174,N_2163);
xnor U2222 (N_2222,N_2183,N_2185);
nand U2223 (N_2223,N_2172,N_2161);
xnor U2224 (N_2224,N_2170,N_2193);
and U2225 (N_2225,N_2182,N_2167);
and U2226 (N_2226,N_2184,N_2165);
and U2227 (N_2227,N_2156,N_2170);
nor U2228 (N_2228,N_2179,N_2199);
nand U2229 (N_2229,N_2173,N_2189);
and U2230 (N_2230,N_2176,N_2179);
xor U2231 (N_2231,N_2183,N_2179);
and U2232 (N_2232,N_2175,N_2176);
nor U2233 (N_2233,N_2176,N_2185);
xor U2234 (N_2234,N_2192,N_2184);
xor U2235 (N_2235,N_2163,N_2179);
and U2236 (N_2236,N_2171,N_2193);
nand U2237 (N_2237,N_2175,N_2180);
or U2238 (N_2238,N_2165,N_2154);
or U2239 (N_2239,N_2163,N_2178);
or U2240 (N_2240,N_2185,N_2156);
and U2241 (N_2241,N_2181,N_2155);
xnor U2242 (N_2242,N_2183,N_2190);
xnor U2243 (N_2243,N_2158,N_2185);
and U2244 (N_2244,N_2154,N_2199);
and U2245 (N_2245,N_2159,N_2175);
and U2246 (N_2246,N_2188,N_2175);
and U2247 (N_2247,N_2171,N_2160);
xor U2248 (N_2248,N_2168,N_2190);
or U2249 (N_2249,N_2170,N_2196);
or U2250 (N_2250,N_2213,N_2208);
nor U2251 (N_2251,N_2211,N_2233);
and U2252 (N_2252,N_2242,N_2214);
xnor U2253 (N_2253,N_2247,N_2222);
or U2254 (N_2254,N_2217,N_2200);
nand U2255 (N_2255,N_2236,N_2203);
nor U2256 (N_2256,N_2237,N_2238);
nand U2257 (N_2257,N_2202,N_2219);
nor U2258 (N_2258,N_2230,N_2224);
nand U2259 (N_2259,N_2209,N_2204);
xnor U2260 (N_2260,N_2212,N_2234);
and U2261 (N_2261,N_2221,N_2246);
or U2262 (N_2262,N_2218,N_2229);
nand U2263 (N_2263,N_2216,N_2220);
nand U2264 (N_2264,N_2244,N_2232);
or U2265 (N_2265,N_2210,N_2215);
or U2266 (N_2266,N_2207,N_2231);
nand U2267 (N_2267,N_2235,N_2201);
and U2268 (N_2268,N_2245,N_2227);
nand U2269 (N_2269,N_2248,N_2228);
or U2270 (N_2270,N_2240,N_2205);
nor U2271 (N_2271,N_2239,N_2241);
nor U2272 (N_2272,N_2249,N_2223);
nand U2273 (N_2273,N_2243,N_2226);
nor U2274 (N_2274,N_2225,N_2206);
xnor U2275 (N_2275,N_2211,N_2225);
nor U2276 (N_2276,N_2205,N_2218);
nor U2277 (N_2277,N_2232,N_2245);
nor U2278 (N_2278,N_2247,N_2213);
or U2279 (N_2279,N_2209,N_2237);
xor U2280 (N_2280,N_2222,N_2242);
nand U2281 (N_2281,N_2205,N_2235);
nor U2282 (N_2282,N_2243,N_2211);
xnor U2283 (N_2283,N_2212,N_2246);
xor U2284 (N_2284,N_2243,N_2246);
xor U2285 (N_2285,N_2207,N_2205);
nor U2286 (N_2286,N_2248,N_2224);
and U2287 (N_2287,N_2226,N_2238);
and U2288 (N_2288,N_2249,N_2229);
nand U2289 (N_2289,N_2211,N_2240);
nor U2290 (N_2290,N_2200,N_2232);
or U2291 (N_2291,N_2232,N_2222);
nor U2292 (N_2292,N_2214,N_2244);
nand U2293 (N_2293,N_2218,N_2246);
and U2294 (N_2294,N_2222,N_2207);
nand U2295 (N_2295,N_2230,N_2244);
nand U2296 (N_2296,N_2203,N_2219);
nand U2297 (N_2297,N_2202,N_2215);
or U2298 (N_2298,N_2220,N_2233);
and U2299 (N_2299,N_2243,N_2205);
and U2300 (N_2300,N_2293,N_2253);
and U2301 (N_2301,N_2281,N_2263);
xnor U2302 (N_2302,N_2286,N_2299);
xor U2303 (N_2303,N_2298,N_2290);
nor U2304 (N_2304,N_2297,N_2265);
or U2305 (N_2305,N_2260,N_2291);
nor U2306 (N_2306,N_2256,N_2285);
xor U2307 (N_2307,N_2278,N_2289);
and U2308 (N_2308,N_2270,N_2267);
nand U2309 (N_2309,N_2251,N_2250);
nor U2310 (N_2310,N_2268,N_2271);
nor U2311 (N_2311,N_2294,N_2287);
xnor U2312 (N_2312,N_2277,N_2292);
xor U2313 (N_2313,N_2266,N_2275);
and U2314 (N_2314,N_2295,N_2279);
xnor U2315 (N_2315,N_2269,N_2259);
or U2316 (N_2316,N_2261,N_2283);
xor U2317 (N_2317,N_2296,N_2282);
and U2318 (N_2318,N_2284,N_2258);
nor U2319 (N_2319,N_2257,N_2262);
nor U2320 (N_2320,N_2264,N_2254);
xnor U2321 (N_2321,N_2274,N_2280);
nand U2322 (N_2322,N_2252,N_2273);
xor U2323 (N_2323,N_2272,N_2288);
xnor U2324 (N_2324,N_2276,N_2255);
xnor U2325 (N_2325,N_2290,N_2252);
or U2326 (N_2326,N_2263,N_2273);
nand U2327 (N_2327,N_2254,N_2294);
or U2328 (N_2328,N_2283,N_2286);
or U2329 (N_2329,N_2294,N_2255);
or U2330 (N_2330,N_2298,N_2281);
and U2331 (N_2331,N_2289,N_2266);
nand U2332 (N_2332,N_2272,N_2285);
nor U2333 (N_2333,N_2288,N_2286);
nand U2334 (N_2334,N_2273,N_2256);
xor U2335 (N_2335,N_2270,N_2268);
nand U2336 (N_2336,N_2279,N_2270);
and U2337 (N_2337,N_2258,N_2294);
xnor U2338 (N_2338,N_2252,N_2250);
xor U2339 (N_2339,N_2254,N_2297);
nand U2340 (N_2340,N_2299,N_2264);
and U2341 (N_2341,N_2287,N_2277);
and U2342 (N_2342,N_2282,N_2276);
nor U2343 (N_2343,N_2276,N_2277);
nand U2344 (N_2344,N_2285,N_2286);
and U2345 (N_2345,N_2250,N_2280);
xor U2346 (N_2346,N_2293,N_2272);
and U2347 (N_2347,N_2268,N_2269);
or U2348 (N_2348,N_2283,N_2263);
nand U2349 (N_2349,N_2250,N_2270);
and U2350 (N_2350,N_2323,N_2325);
nand U2351 (N_2351,N_2347,N_2333);
nand U2352 (N_2352,N_2337,N_2343);
xnor U2353 (N_2353,N_2334,N_2324);
nor U2354 (N_2354,N_2316,N_2311);
nand U2355 (N_2355,N_2305,N_2319);
xnor U2356 (N_2356,N_2338,N_2300);
xnor U2357 (N_2357,N_2329,N_2312);
and U2358 (N_2358,N_2315,N_2340);
and U2359 (N_2359,N_2332,N_2321);
xnor U2360 (N_2360,N_2339,N_2307);
xor U2361 (N_2361,N_2308,N_2304);
xor U2362 (N_2362,N_2322,N_2330);
xor U2363 (N_2363,N_2302,N_2344);
nand U2364 (N_2364,N_2314,N_2301);
or U2365 (N_2365,N_2336,N_2309);
nand U2366 (N_2366,N_2313,N_2317);
or U2367 (N_2367,N_2318,N_2306);
nor U2368 (N_2368,N_2345,N_2303);
nand U2369 (N_2369,N_2328,N_2320);
xor U2370 (N_2370,N_2335,N_2310);
or U2371 (N_2371,N_2348,N_2326);
nor U2372 (N_2372,N_2327,N_2341);
xor U2373 (N_2373,N_2342,N_2349);
nand U2374 (N_2374,N_2331,N_2346);
nand U2375 (N_2375,N_2335,N_2336);
or U2376 (N_2376,N_2303,N_2336);
and U2377 (N_2377,N_2308,N_2306);
xnor U2378 (N_2378,N_2306,N_2348);
nand U2379 (N_2379,N_2339,N_2337);
or U2380 (N_2380,N_2324,N_2317);
xor U2381 (N_2381,N_2302,N_2323);
nand U2382 (N_2382,N_2325,N_2338);
xor U2383 (N_2383,N_2312,N_2334);
xor U2384 (N_2384,N_2313,N_2306);
nor U2385 (N_2385,N_2335,N_2309);
or U2386 (N_2386,N_2308,N_2342);
nor U2387 (N_2387,N_2307,N_2324);
or U2388 (N_2388,N_2333,N_2306);
nand U2389 (N_2389,N_2305,N_2335);
nand U2390 (N_2390,N_2302,N_2301);
xor U2391 (N_2391,N_2349,N_2302);
nor U2392 (N_2392,N_2311,N_2340);
or U2393 (N_2393,N_2319,N_2328);
nand U2394 (N_2394,N_2330,N_2334);
or U2395 (N_2395,N_2314,N_2338);
or U2396 (N_2396,N_2317,N_2334);
and U2397 (N_2397,N_2339,N_2317);
xor U2398 (N_2398,N_2323,N_2317);
nand U2399 (N_2399,N_2316,N_2336);
nand U2400 (N_2400,N_2368,N_2377);
nand U2401 (N_2401,N_2384,N_2369);
or U2402 (N_2402,N_2353,N_2394);
nand U2403 (N_2403,N_2395,N_2373);
nand U2404 (N_2404,N_2392,N_2350);
nor U2405 (N_2405,N_2362,N_2357);
nand U2406 (N_2406,N_2390,N_2383);
and U2407 (N_2407,N_2355,N_2376);
nor U2408 (N_2408,N_2371,N_2378);
and U2409 (N_2409,N_2397,N_2372);
nand U2410 (N_2410,N_2379,N_2367);
xnor U2411 (N_2411,N_2354,N_2389);
xnor U2412 (N_2412,N_2366,N_2380);
and U2413 (N_2413,N_2388,N_2358);
or U2414 (N_2414,N_2370,N_2396);
xnor U2415 (N_2415,N_2374,N_2351);
nor U2416 (N_2416,N_2382,N_2398);
nor U2417 (N_2417,N_2352,N_2391);
nand U2418 (N_2418,N_2386,N_2356);
nor U2419 (N_2419,N_2375,N_2381);
or U2420 (N_2420,N_2385,N_2359);
nor U2421 (N_2421,N_2364,N_2361);
nand U2422 (N_2422,N_2387,N_2360);
xnor U2423 (N_2423,N_2399,N_2365);
nor U2424 (N_2424,N_2363,N_2393);
xor U2425 (N_2425,N_2382,N_2360);
or U2426 (N_2426,N_2396,N_2365);
nand U2427 (N_2427,N_2381,N_2377);
xor U2428 (N_2428,N_2389,N_2352);
xor U2429 (N_2429,N_2382,N_2397);
nor U2430 (N_2430,N_2353,N_2352);
nor U2431 (N_2431,N_2396,N_2350);
nor U2432 (N_2432,N_2373,N_2355);
or U2433 (N_2433,N_2362,N_2363);
nand U2434 (N_2434,N_2390,N_2355);
or U2435 (N_2435,N_2355,N_2384);
and U2436 (N_2436,N_2360,N_2355);
xor U2437 (N_2437,N_2386,N_2362);
or U2438 (N_2438,N_2354,N_2399);
or U2439 (N_2439,N_2373,N_2359);
xnor U2440 (N_2440,N_2371,N_2390);
nor U2441 (N_2441,N_2377,N_2385);
xor U2442 (N_2442,N_2395,N_2363);
or U2443 (N_2443,N_2385,N_2391);
xnor U2444 (N_2444,N_2365,N_2380);
or U2445 (N_2445,N_2353,N_2382);
and U2446 (N_2446,N_2356,N_2384);
xnor U2447 (N_2447,N_2373,N_2376);
nand U2448 (N_2448,N_2394,N_2389);
nand U2449 (N_2449,N_2394,N_2364);
and U2450 (N_2450,N_2425,N_2428);
nor U2451 (N_2451,N_2434,N_2423);
nand U2452 (N_2452,N_2430,N_2444);
nor U2453 (N_2453,N_2422,N_2403);
or U2454 (N_2454,N_2417,N_2424);
nor U2455 (N_2455,N_2415,N_2438);
xor U2456 (N_2456,N_2446,N_2420);
and U2457 (N_2457,N_2414,N_2413);
xnor U2458 (N_2458,N_2448,N_2447);
or U2459 (N_2459,N_2432,N_2402);
xnor U2460 (N_2460,N_2429,N_2400);
and U2461 (N_2461,N_2419,N_2436);
or U2462 (N_2462,N_2426,N_2439);
xnor U2463 (N_2463,N_2449,N_2431);
xnor U2464 (N_2464,N_2411,N_2416);
xnor U2465 (N_2465,N_2407,N_2401);
and U2466 (N_2466,N_2435,N_2405);
nor U2467 (N_2467,N_2409,N_2410);
nor U2468 (N_2468,N_2408,N_2427);
xnor U2469 (N_2469,N_2406,N_2421);
xnor U2470 (N_2470,N_2433,N_2445);
xnor U2471 (N_2471,N_2443,N_2437);
nand U2472 (N_2472,N_2442,N_2404);
xor U2473 (N_2473,N_2412,N_2441);
xnor U2474 (N_2474,N_2418,N_2440);
or U2475 (N_2475,N_2438,N_2405);
nor U2476 (N_2476,N_2405,N_2414);
nor U2477 (N_2477,N_2447,N_2432);
xor U2478 (N_2478,N_2432,N_2437);
xor U2479 (N_2479,N_2412,N_2406);
nand U2480 (N_2480,N_2430,N_2402);
nand U2481 (N_2481,N_2419,N_2422);
xor U2482 (N_2482,N_2439,N_2417);
nand U2483 (N_2483,N_2442,N_2449);
or U2484 (N_2484,N_2424,N_2439);
or U2485 (N_2485,N_2443,N_2448);
nor U2486 (N_2486,N_2436,N_2431);
nor U2487 (N_2487,N_2437,N_2414);
xor U2488 (N_2488,N_2401,N_2405);
xor U2489 (N_2489,N_2430,N_2408);
or U2490 (N_2490,N_2416,N_2423);
nand U2491 (N_2491,N_2420,N_2437);
or U2492 (N_2492,N_2416,N_2443);
nand U2493 (N_2493,N_2438,N_2445);
nand U2494 (N_2494,N_2416,N_2432);
nand U2495 (N_2495,N_2417,N_2441);
nand U2496 (N_2496,N_2427,N_2448);
nand U2497 (N_2497,N_2402,N_2416);
xnor U2498 (N_2498,N_2441,N_2430);
and U2499 (N_2499,N_2423,N_2442);
xnor U2500 (N_2500,N_2452,N_2465);
and U2501 (N_2501,N_2453,N_2490);
or U2502 (N_2502,N_2456,N_2497);
or U2503 (N_2503,N_2473,N_2478);
xnor U2504 (N_2504,N_2467,N_2464);
and U2505 (N_2505,N_2450,N_2487);
nand U2506 (N_2506,N_2462,N_2484);
nand U2507 (N_2507,N_2458,N_2483);
and U2508 (N_2508,N_2474,N_2481);
xor U2509 (N_2509,N_2455,N_2482);
nand U2510 (N_2510,N_2461,N_2493);
nand U2511 (N_2511,N_2480,N_2498);
nand U2512 (N_2512,N_2475,N_2470);
and U2513 (N_2513,N_2460,N_2496);
xor U2514 (N_2514,N_2491,N_2466);
nor U2515 (N_2515,N_2488,N_2479);
nor U2516 (N_2516,N_2451,N_2477);
nor U2517 (N_2517,N_2476,N_2463);
nand U2518 (N_2518,N_2486,N_2492);
and U2519 (N_2519,N_2469,N_2454);
nor U2520 (N_2520,N_2495,N_2499);
nor U2521 (N_2521,N_2485,N_2459);
xnor U2522 (N_2522,N_2471,N_2468);
and U2523 (N_2523,N_2472,N_2457);
nor U2524 (N_2524,N_2489,N_2494);
xor U2525 (N_2525,N_2486,N_2490);
nand U2526 (N_2526,N_2497,N_2490);
nor U2527 (N_2527,N_2487,N_2468);
or U2528 (N_2528,N_2480,N_2455);
and U2529 (N_2529,N_2454,N_2479);
nand U2530 (N_2530,N_2450,N_2466);
and U2531 (N_2531,N_2459,N_2467);
and U2532 (N_2532,N_2471,N_2458);
nor U2533 (N_2533,N_2488,N_2478);
and U2534 (N_2534,N_2460,N_2490);
nor U2535 (N_2535,N_2490,N_2463);
xnor U2536 (N_2536,N_2482,N_2458);
and U2537 (N_2537,N_2452,N_2475);
xor U2538 (N_2538,N_2451,N_2453);
and U2539 (N_2539,N_2455,N_2462);
xnor U2540 (N_2540,N_2479,N_2463);
or U2541 (N_2541,N_2484,N_2470);
xnor U2542 (N_2542,N_2456,N_2460);
and U2543 (N_2543,N_2497,N_2464);
xor U2544 (N_2544,N_2464,N_2470);
xor U2545 (N_2545,N_2491,N_2489);
nand U2546 (N_2546,N_2496,N_2476);
or U2547 (N_2547,N_2477,N_2470);
or U2548 (N_2548,N_2473,N_2466);
xor U2549 (N_2549,N_2489,N_2450);
and U2550 (N_2550,N_2519,N_2539);
nand U2551 (N_2551,N_2535,N_2546);
xor U2552 (N_2552,N_2523,N_2533);
xnor U2553 (N_2553,N_2508,N_2547);
or U2554 (N_2554,N_2540,N_2527);
nor U2555 (N_2555,N_2536,N_2515);
and U2556 (N_2556,N_2520,N_2518);
xnor U2557 (N_2557,N_2500,N_2538);
nand U2558 (N_2558,N_2501,N_2521);
and U2559 (N_2559,N_2530,N_2509);
nand U2560 (N_2560,N_2534,N_2517);
nor U2561 (N_2561,N_2528,N_2516);
nand U2562 (N_2562,N_2513,N_2545);
or U2563 (N_2563,N_2537,N_2504);
nor U2564 (N_2564,N_2503,N_2524);
nand U2565 (N_2565,N_2505,N_2548);
and U2566 (N_2566,N_2502,N_2514);
xor U2567 (N_2567,N_2529,N_2506);
xor U2568 (N_2568,N_2522,N_2511);
nand U2569 (N_2569,N_2525,N_2543);
or U2570 (N_2570,N_2532,N_2541);
or U2571 (N_2571,N_2544,N_2549);
or U2572 (N_2572,N_2542,N_2510);
or U2573 (N_2573,N_2531,N_2526);
nor U2574 (N_2574,N_2512,N_2507);
or U2575 (N_2575,N_2501,N_2544);
xnor U2576 (N_2576,N_2537,N_2549);
and U2577 (N_2577,N_2502,N_2544);
or U2578 (N_2578,N_2545,N_2508);
nor U2579 (N_2579,N_2521,N_2523);
xnor U2580 (N_2580,N_2512,N_2525);
and U2581 (N_2581,N_2539,N_2523);
and U2582 (N_2582,N_2509,N_2540);
nor U2583 (N_2583,N_2547,N_2534);
nor U2584 (N_2584,N_2540,N_2535);
xor U2585 (N_2585,N_2538,N_2518);
xnor U2586 (N_2586,N_2530,N_2502);
nand U2587 (N_2587,N_2503,N_2516);
and U2588 (N_2588,N_2511,N_2503);
nand U2589 (N_2589,N_2516,N_2511);
xnor U2590 (N_2590,N_2511,N_2512);
or U2591 (N_2591,N_2516,N_2510);
xor U2592 (N_2592,N_2538,N_2534);
and U2593 (N_2593,N_2549,N_2538);
nand U2594 (N_2594,N_2512,N_2524);
nor U2595 (N_2595,N_2546,N_2543);
or U2596 (N_2596,N_2504,N_2548);
nor U2597 (N_2597,N_2538,N_2514);
and U2598 (N_2598,N_2535,N_2539);
and U2599 (N_2599,N_2532,N_2517);
nand U2600 (N_2600,N_2556,N_2555);
and U2601 (N_2601,N_2557,N_2559);
nand U2602 (N_2602,N_2558,N_2599);
nand U2603 (N_2603,N_2581,N_2578);
or U2604 (N_2604,N_2565,N_2596);
or U2605 (N_2605,N_2593,N_2572);
and U2606 (N_2606,N_2588,N_2564);
nor U2607 (N_2607,N_2554,N_2550);
nand U2608 (N_2608,N_2582,N_2598);
and U2609 (N_2609,N_2567,N_2586);
nor U2610 (N_2610,N_2560,N_2577);
xnor U2611 (N_2611,N_2566,N_2592);
xor U2612 (N_2612,N_2568,N_2579);
and U2613 (N_2613,N_2569,N_2584);
nand U2614 (N_2614,N_2571,N_2551);
and U2615 (N_2615,N_2574,N_2591);
nand U2616 (N_2616,N_2597,N_2553);
and U2617 (N_2617,N_2563,N_2590);
nand U2618 (N_2618,N_2583,N_2562);
xnor U2619 (N_2619,N_2552,N_2561);
and U2620 (N_2620,N_2575,N_2580);
xnor U2621 (N_2621,N_2576,N_2587);
or U2622 (N_2622,N_2595,N_2573);
and U2623 (N_2623,N_2585,N_2594);
or U2624 (N_2624,N_2589,N_2570);
nand U2625 (N_2625,N_2563,N_2551);
and U2626 (N_2626,N_2564,N_2587);
or U2627 (N_2627,N_2595,N_2575);
or U2628 (N_2628,N_2567,N_2575);
nor U2629 (N_2629,N_2556,N_2588);
nor U2630 (N_2630,N_2581,N_2582);
nor U2631 (N_2631,N_2567,N_2598);
nor U2632 (N_2632,N_2558,N_2577);
or U2633 (N_2633,N_2586,N_2584);
nor U2634 (N_2634,N_2580,N_2570);
or U2635 (N_2635,N_2582,N_2597);
nand U2636 (N_2636,N_2584,N_2595);
nand U2637 (N_2637,N_2561,N_2599);
or U2638 (N_2638,N_2583,N_2551);
nand U2639 (N_2639,N_2596,N_2588);
nor U2640 (N_2640,N_2556,N_2580);
or U2641 (N_2641,N_2598,N_2581);
nand U2642 (N_2642,N_2585,N_2563);
nor U2643 (N_2643,N_2567,N_2556);
nor U2644 (N_2644,N_2577,N_2574);
or U2645 (N_2645,N_2565,N_2569);
xor U2646 (N_2646,N_2558,N_2564);
and U2647 (N_2647,N_2572,N_2573);
nor U2648 (N_2648,N_2599,N_2580);
nand U2649 (N_2649,N_2572,N_2599);
nor U2650 (N_2650,N_2635,N_2637);
and U2651 (N_2651,N_2647,N_2631);
nor U2652 (N_2652,N_2633,N_2607);
nor U2653 (N_2653,N_2612,N_2615);
xor U2654 (N_2654,N_2608,N_2643);
or U2655 (N_2655,N_2625,N_2623);
xnor U2656 (N_2656,N_2644,N_2601);
nand U2657 (N_2657,N_2626,N_2609);
nand U2658 (N_2658,N_2632,N_2638);
nor U2659 (N_2659,N_2619,N_2645);
or U2660 (N_2660,N_2603,N_2622);
xor U2661 (N_2661,N_2613,N_2628);
and U2662 (N_2662,N_2642,N_2627);
xnor U2663 (N_2663,N_2614,N_2639);
and U2664 (N_2664,N_2634,N_2602);
and U2665 (N_2665,N_2616,N_2641);
nor U2666 (N_2666,N_2629,N_2624);
nand U2667 (N_2667,N_2621,N_2600);
and U2668 (N_2668,N_2620,N_2649);
nor U2669 (N_2669,N_2605,N_2606);
and U2670 (N_2670,N_2617,N_2610);
or U2671 (N_2671,N_2636,N_2646);
xor U2672 (N_2672,N_2618,N_2611);
and U2673 (N_2673,N_2640,N_2630);
xor U2674 (N_2674,N_2648,N_2604);
and U2675 (N_2675,N_2616,N_2614);
and U2676 (N_2676,N_2612,N_2635);
xnor U2677 (N_2677,N_2616,N_2624);
nand U2678 (N_2678,N_2629,N_2633);
and U2679 (N_2679,N_2613,N_2626);
xnor U2680 (N_2680,N_2618,N_2609);
xor U2681 (N_2681,N_2632,N_2642);
nor U2682 (N_2682,N_2640,N_2605);
and U2683 (N_2683,N_2632,N_2603);
nand U2684 (N_2684,N_2623,N_2636);
xor U2685 (N_2685,N_2639,N_2633);
nor U2686 (N_2686,N_2643,N_2609);
and U2687 (N_2687,N_2641,N_2635);
nand U2688 (N_2688,N_2640,N_2637);
xor U2689 (N_2689,N_2619,N_2602);
nor U2690 (N_2690,N_2619,N_2629);
xor U2691 (N_2691,N_2620,N_2601);
and U2692 (N_2692,N_2609,N_2646);
nand U2693 (N_2693,N_2638,N_2600);
nand U2694 (N_2694,N_2637,N_2609);
nand U2695 (N_2695,N_2615,N_2618);
nand U2696 (N_2696,N_2642,N_2646);
or U2697 (N_2697,N_2637,N_2621);
xnor U2698 (N_2698,N_2612,N_2631);
nor U2699 (N_2699,N_2645,N_2614);
and U2700 (N_2700,N_2654,N_2668);
xor U2701 (N_2701,N_2691,N_2672);
nand U2702 (N_2702,N_2675,N_2669);
and U2703 (N_2703,N_2680,N_2673);
xnor U2704 (N_2704,N_2666,N_2699);
or U2705 (N_2705,N_2653,N_2671);
nand U2706 (N_2706,N_2698,N_2650);
xor U2707 (N_2707,N_2693,N_2690);
xor U2708 (N_2708,N_2682,N_2679);
xnor U2709 (N_2709,N_2664,N_2695);
nand U2710 (N_2710,N_2697,N_2660);
and U2711 (N_2711,N_2687,N_2696);
nand U2712 (N_2712,N_2677,N_2658);
xnor U2713 (N_2713,N_2657,N_2655);
and U2714 (N_2714,N_2678,N_2689);
nand U2715 (N_2715,N_2692,N_2681);
and U2716 (N_2716,N_2656,N_2676);
nand U2717 (N_2717,N_2667,N_2651);
or U2718 (N_2718,N_2663,N_2670);
or U2719 (N_2719,N_2674,N_2662);
nor U2720 (N_2720,N_2686,N_2665);
nor U2721 (N_2721,N_2685,N_2652);
xnor U2722 (N_2722,N_2694,N_2661);
nand U2723 (N_2723,N_2659,N_2684);
and U2724 (N_2724,N_2683,N_2688);
nand U2725 (N_2725,N_2686,N_2658);
or U2726 (N_2726,N_2689,N_2666);
nor U2727 (N_2727,N_2691,N_2653);
nor U2728 (N_2728,N_2682,N_2691);
and U2729 (N_2729,N_2696,N_2670);
or U2730 (N_2730,N_2693,N_2684);
nand U2731 (N_2731,N_2682,N_2690);
and U2732 (N_2732,N_2655,N_2695);
and U2733 (N_2733,N_2676,N_2688);
and U2734 (N_2734,N_2682,N_2663);
nor U2735 (N_2735,N_2666,N_2651);
or U2736 (N_2736,N_2650,N_2691);
or U2737 (N_2737,N_2686,N_2654);
xor U2738 (N_2738,N_2694,N_2692);
nor U2739 (N_2739,N_2688,N_2653);
nor U2740 (N_2740,N_2694,N_2680);
or U2741 (N_2741,N_2675,N_2679);
xor U2742 (N_2742,N_2699,N_2661);
nand U2743 (N_2743,N_2671,N_2687);
xor U2744 (N_2744,N_2664,N_2653);
xnor U2745 (N_2745,N_2665,N_2664);
nor U2746 (N_2746,N_2674,N_2656);
nand U2747 (N_2747,N_2671,N_2698);
nor U2748 (N_2748,N_2674,N_2666);
xor U2749 (N_2749,N_2677,N_2678);
nor U2750 (N_2750,N_2722,N_2719);
and U2751 (N_2751,N_2737,N_2733);
or U2752 (N_2752,N_2701,N_2723);
or U2753 (N_2753,N_2747,N_2736);
and U2754 (N_2754,N_2741,N_2749);
or U2755 (N_2755,N_2727,N_2725);
xnor U2756 (N_2756,N_2717,N_2718);
nand U2757 (N_2757,N_2707,N_2726);
nor U2758 (N_2758,N_2724,N_2740);
nand U2759 (N_2759,N_2710,N_2709);
nand U2760 (N_2760,N_2700,N_2730);
nand U2761 (N_2761,N_2721,N_2716);
and U2762 (N_2762,N_2745,N_2704);
nor U2763 (N_2763,N_2706,N_2744);
xor U2764 (N_2764,N_2729,N_2732);
and U2765 (N_2765,N_2734,N_2748);
or U2766 (N_2766,N_2731,N_2702);
or U2767 (N_2767,N_2720,N_2742);
nand U2768 (N_2768,N_2743,N_2746);
nor U2769 (N_2769,N_2712,N_2705);
xor U2770 (N_2770,N_2735,N_2703);
xnor U2771 (N_2771,N_2715,N_2714);
xor U2772 (N_2772,N_2738,N_2739);
nor U2773 (N_2773,N_2711,N_2728);
or U2774 (N_2774,N_2713,N_2708);
nand U2775 (N_2775,N_2729,N_2725);
xnor U2776 (N_2776,N_2710,N_2742);
xnor U2777 (N_2777,N_2734,N_2713);
and U2778 (N_2778,N_2729,N_2700);
nand U2779 (N_2779,N_2738,N_2736);
nand U2780 (N_2780,N_2709,N_2729);
and U2781 (N_2781,N_2709,N_2715);
xnor U2782 (N_2782,N_2703,N_2700);
or U2783 (N_2783,N_2730,N_2704);
or U2784 (N_2784,N_2706,N_2709);
nand U2785 (N_2785,N_2735,N_2737);
or U2786 (N_2786,N_2736,N_2723);
or U2787 (N_2787,N_2736,N_2743);
nand U2788 (N_2788,N_2701,N_2745);
and U2789 (N_2789,N_2713,N_2701);
or U2790 (N_2790,N_2705,N_2742);
nand U2791 (N_2791,N_2742,N_2736);
nor U2792 (N_2792,N_2721,N_2703);
xor U2793 (N_2793,N_2700,N_2734);
xnor U2794 (N_2794,N_2735,N_2718);
or U2795 (N_2795,N_2713,N_2720);
nand U2796 (N_2796,N_2713,N_2738);
nand U2797 (N_2797,N_2734,N_2720);
and U2798 (N_2798,N_2706,N_2710);
or U2799 (N_2799,N_2720,N_2717);
nand U2800 (N_2800,N_2760,N_2785);
nand U2801 (N_2801,N_2766,N_2778);
or U2802 (N_2802,N_2757,N_2754);
xor U2803 (N_2803,N_2782,N_2765);
nand U2804 (N_2804,N_2753,N_2799);
nand U2805 (N_2805,N_2789,N_2786);
and U2806 (N_2806,N_2784,N_2772);
xor U2807 (N_2807,N_2780,N_2792);
xor U2808 (N_2808,N_2769,N_2770);
xor U2809 (N_2809,N_2751,N_2768);
or U2810 (N_2810,N_2763,N_2779);
nand U2811 (N_2811,N_2795,N_2759);
or U2812 (N_2812,N_2756,N_2787);
nand U2813 (N_2813,N_2750,N_2798);
nor U2814 (N_2814,N_2773,N_2762);
nand U2815 (N_2815,N_2752,N_2774);
xnor U2816 (N_2816,N_2764,N_2758);
nand U2817 (N_2817,N_2796,N_2755);
and U2818 (N_2818,N_2776,N_2777);
xnor U2819 (N_2819,N_2793,N_2797);
nand U2820 (N_2820,N_2790,N_2783);
nand U2821 (N_2821,N_2771,N_2794);
nor U2822 (N_2822,N_2791,N_2775);
and U2823 (N_2823,N_2761,N_2767);
nand U2824 (N_2824,N_2788,N_2781);
or U2825 (N_2825,N_2781,N_2777);
and U2826 (N_2826,N_2774,N_2798);
xor U2827 (N_2827,N_2767,N_2768);
xnor U2828 (N_2828,N_2799,N_2763);
nand U2829 (N_2829,N_2791,N_2794);
or U2830 (N_2830,N_2780,N_2767);
and U2831 (N_2831,N_2762,N_2784);
xnor U2832 (N_2832,N_2783,N_2772);
and U2833 (N_2833,N_2774,N_2779);
and U2834 (N_2834,N_2758,N_2752);
xnor U2835 (N_2835,N_2758,N_2799);
nor U2836 (N_2836,N_2767,N_2764);
nor U2837 (N_2837,N_2771,N_2785);
and U2838 (N_2838,N_2798,N_2762);
and U2839 (N_2839,N_2787,N_2769);
and U2840 (N_2840,N_2777,N_2764);
or U2841 (N_2841,N_2763,N_2783);
xnor U2842 (N_2842,N_2768,N_2786);
or U2843 (N_2843,N_2754,N_2795);
xnor U2844 (N_2844,N_2797,N_2785);
and U2845 (N_2845,N_2768,N_2790);
nor U2846 (N_2846,N_2770,N_2773);
nand U2847 (N_2847,N_2785,N_2765);
and U2848 (N_2848,N_2769,N_2757);
and U2849 (N_2849,N_2781,N_2766);
xnor U2850 (N_2850,N_2811,N_2834);
and U2851 (N_2851,N_2832,N_2810);
or U2852 (N_2852,N_2829,N_2833);
xnor U2853 (N_2853,N_2827,N_2822);
nor U2854 (N_2854,N_2806,N_2813);
nand U2855 (N_2855,N_2817,N_2809);
xnor U2856 (N_2856,N_2802,N_2845);
nand U2857 (N_2857,N_2808,N_2803);
nor U2858 (N_2858,N_2831,N_2805);
or U2859 (N_2859,N_2815,N_2819);
nand U2860 (N_2860,N_2814,N_2830);
xnor U2861 (N_2861,N_2844,N_2816);
xnor U2862 (N_2862,N_2821,N_2820);
xnor U2863 (N_2863,N_2837,N_2842);
nand U2864 (N_2864,N_2801,N_2818);
nor U2865 (N_2865,N_2843,N_2841);
and U2866 (N_2866,N_2826,N_2823);
and U2867 (N_2867,N_2846,N_2835);
nand U2868 (N_2868,N_2840,N_2836);
or U2869 (N_2869,N_2828,N_2825);
and U2870 (N_2870,N_2849,N_2824);
or U2871 (N_2871,N_2812,N_2839);
nor U2872 (N_2872,N_2847,N_2800);
nor U2873 (N_2873,N_2807,N_2848);
xor U2874 (N_2874,N_2804,N_2838);
nor U2875 (N_2875,N_2825,N_2810);
nand U2876 (N_2876,N_2808,N_2802);
and U2877 (N_2877,N_2812,N_2814);
or U2878 (N_2878,N_2836,N_2801);
and U2879 (N_2879,N_2818,N_2833);
xnor U2880 (N_2880,N_2825,N_2833);
nor U2881 (N_2881,N_2815,N_2817);
and U2882 (N_2882,N_2846,N_2847);
and U2883 (N_2883,N_2816,N_2819);
or U2884 (N_2884,N_2809,N_2830);
nor U2885 (N_2885,N_2830,N_2849);
nor U2886 (N_2886,N_2819,N_2811);
xor U2887 (N_2887,N_2818,N_2806);
and U2888 (N_2888,N_2817,N_2849);
nor U2889 (N_2889,N_2801,N_2839);
and U2890 (N_2890,N_2804,N_2830);
nand U2891 (N_2891,N_2829,N_2823);
xnor U2892 (N_2892,N_2841,N_2835);
and U2893 (N_2893,N_2810,N_2819);
and U2894 (N_2894,N_2813,N_2831);
nand U2895 (N_2895,N_2820,N_2819);
xor U2896 (N_2896,N_2842,N_2814);
or U2897 (N_2897,N_2801,N_2814);
and U2898 (N_2898,N_2823,N_2812);
xnor U2899 (N_2899,N_2849,N_2843);
nand U2900 (N_2900,N_2870,N_2861);
or U2901 (N_2901,N_2879,N_2852);
or U2902 (N_2902,N_2873,N_2860);
xor U2903 (N_2903,N_2871,N_2855);
xor U2904 (N_2904,N_2898,N_2869);
or U2905 (N_2905,N_2888,N_2857);
nand U2906 (N_2906,N_2864,N_2892);
nor U2907 (N_2907,N_2899,N_2876);
nor U2908 (N_2908,N_2885,N_2897);
nand U2909 (N_2909,N_2887,N_2877);
nor U2910 (N_2910,N_2896,N_2866);
and U2911 (N_2911,N_2889,N_2880);
xor U2912 (N_2912,N_2850,N_2878);
nand U2913 (N_2913,N_2851,N_2854);
nor U2914 (N_2914,N_2858,N_2874);
or U2915 (N_2915,N_2859,N_2883);
or U2916 (N_2916,N_2886,N_2891);
or U2917 (N_2917,N_2875,N_2884);
and U2918 (N_2918,N_2863,N_2893);
or U2919 (N_2919,N_2881,N_2895);
nor U2920 (N_2920,N_2853,N_2856);
or U2921 (N_2921,N_2868,N_2867);
nand U2922 (N_2922,N_2894,N_2882);
or U2923 (N_2923,N_2865,N_2890);
xor U2924 (N_2924,N_2862,N_2872);
nor U2925 (N_2925,N_2894,N_2881);
or U2926 (N_2926,N_2853,N_2896);
or U2927 (N_2927,N_2882,N_2864);
and U2928 (N_2928,N_2862,N_2890);
xor U2929 (N_2929,N_2873,N_2877);
nand U2930 (N_2930,N_2878,N_2890);
or U2931 (N_2931,N_2861,N_2886);
xnor U2932 (N_2932,N_2870,N_2860);
nor U2933 (N_2933,N_2867,N_2876);
nor U2934 (N_2934,N_2891,N_2876);
xor U2935 (N_2935,N_2879,N_2869);
and U2936 (N_2936,N_2897,N_2855);
and U2937 (N_2937,N_2876,N_2886);
or U2938 (N_2938,N_2870,N_2868);
nor U2939 (N_2939,N_2877,N_2885);
nor U2940 (N_2940,N_2873,N_2857);
nand U2941 (N_2941,N_2898,N_2875);
xnor U2942 (N_2942,N_2877,N_2853);
and U2943 (N_2943,N_2896,N_2854);
and U2944 (N_2944,N_2853,N_2886);
nand U2945 (N_2945,N_2898,N_2856);
and U2946 (N_2946,N_2872,N_2889);
nand U2947 (N_2947,N_2855,N_2854);
nand U2948 (N_2948,N_2888,N_2867);
or U2949 (N_2949,N_2859,N_2853);
or U2950 (N_2950,N_2918,N_2920);
nand U2951 (N_2951,N_2925,N_2939);
and U2952 (N_2952,N_2938,N_2933);
nor U2953 (N_2953,N_2935,N_2926);
and U2954 (N_2954,N_2936,N_2911);
or U2955 (N_2955,N_2900,N_2921);
nand U2956 (N_2956,N_2902,N_2905);
nor U2957 (N_2957,N_2931,N_2941);
or U2958 (N_2958,N_2906,N_2901);
or U2959 (N_2959,N_2912,N_2948);
or U2960 (N_2960,N_2947,N_2930);
nand U2961 (N_2961,N_2915,N_2919);
nand U2962 (N_2962,N_2916,N_2907);
or U2963 (N_2963,N_2913,N_2903);
nor U2964 (N_2964,N_2928,N_2946);
xnor U2965 (N_2965,N_2909,N_2943);
nor U2966 (N_2966,N_2917,N_2914);
nand U2967 (N_2967,N_2929,N_2942);
xor U2968 (N_2968,N_2932,N_2922);
and U2969 (N_2969,N_2924,N_2949);
or U2970 (N_2970,N_2945,N_2908);
and U2971 (N_2971,N_2904,N_2934);
nor U2972 (N_2972,N_2923,N_2940);
or U2973 (N_2973,N_2944,N_2937);
and U2974 (N_2974,N_2910,N_2927);
and U2975 (N_2975,N_2912,N_2908);
or U2976 (N_2976,N_2938,N_2942);
and U2977 (N_2977,N_2946,N_2925);
xnor U2978 (N_2978,N_2933,N_2939);
xor U2979 (N_2979,N_2927,N_2904);
nand U2980 (N_2980,N_2933,N_2908);
and U2981 (N_2981,N_2919,N_2926);
and U2982 (N_2982,N_2931,N_2937);
xor U2983 (N_2983,N_2927,N_2920);
or U2984 (N_2984,N_2949,N_2918);
nor U2985 (N_2985,N_2918,N_2905);
and U2986 (N_2986,N_2934,N_2937);
xnor U2987 (N_2987,N_2944,N_2925);
or U2988 (N_2988,N_2931,N_2900);
or U2989 (N_2989,N_2926,N_2921);
xor U2990 (N_2990,N_2921,N_2946);
nand U2991 (N_2991,N_2913,N_2925);
nor U2992 (N_2992,N_2925,N_2924);
nand U2993 (N_2993,N_2936,N_2902);
nand U2994 (N_2994,N_2918,N_2946);
and U2995 (N_2995,N_2937,N_2913);
or U2996 (N_2996,N_2905,N_2933);
and U2997 (N_2997,N_2942,N_2934);
and U2998 (N_2998,N_2949,N_2901);
nand U2999 (N_2999,N_2948,N_2910);
or UO_0 (O_0,N_2974,N_2966);
or UO_1 (O_1,N_2997,N_2968);
nor UO_2 (O_2,N_2950,N_2976);
xnor UO_3 (O_3,N_2989,N_2951);
or UO_4 (O_4,N_2981,N_2965);
xnor UO_5 (O_5,N_2978,N_2987);
nand UO_6 (O_6,N_2962,N_2990);
xnor UO_7 (O_7,N_2956,N_2961);
or UO_8 (O_8,N_2993,N_2992);
xor UO_9 (O_9,N_2986,N_2973);
or UO_10 (O_10,N_2991,N_2963);
and UO_11 (O_11,N_2975,N_2985);
and UO_12 (O_12,N_2977,N_2984);
xor UO_13 (O_13,N_2952,N_2955);
nor UO_14 (O_14,N_2999,N_2954);
nand UO_15 (O_15,N_2994,N_2988);
nor UO_16 (O_16,N_2970,N_2983);
and UO_17 (O_17,N_2957,N_2979);
and UO_18 (O_18,N_2995,N_2958);
or UO_19 (O_19,N_2960,N_2980);
nor UO_20 (O_20,N_2971,N_2967);
nand UO_21 (O_21,N_2964,N_2959);
and UO_22 (O_22,N_2972,N_2982);
or UO_23 (O_23,N_2996,N_2969);
or UO_24 (O_24,N_2998,N_2953);
or UO_25 (O_25,N_2996,N_2990);
nor UO_26 (O_26,N_2994,N_2987);
nand UO_27 (O_27,N_2963,N_2961);
nand UO_28 (O_28,N_2981,N_2958);
nor UO_29 (O_29,N_2973,N_2998);
and UO_30 (O_30,N_2983,N_2995);
nor UO_31 (O_31,N_2955,N_2979);
nand UO_32 (O_32,N_2951,N_2984);
nand UO_33 (O_33,N_2954,N_2992);
or UO_34 (O_34,N_2985,N_2957);
nand UO_35 (O_35,N_2963,N_2992);
or UO_36 (O_36,N_2999,N_2970);
nand UO_37 (O_37,N_2968,N_2990);
or UO_38 (O_38,N_2982,N_2951);
and UO_39 (O_39,N_2981,N_2961);
or UO_40 (O_40,N_2986,N_2966);
and UO_41 (O_41,N_2953,N_2971);
and UO_42 (O_42,N_2972,N_2997);
or UO_43 (O_43,N_2984,N_2955);
nand UO_44 (O_44,N_2971,N_2969);
nor UO_45 (O_45,N_2967,N_2983);
or UO_46 (O_46,N_2996,N_2951);
nand UO_47 (O_47,N_2975,N_2974);
and UO_48 (O_48,N_2981,N_2970);
or UO_49 (O_49,N_2960,N_2953);
or UO_50 (O_50,N_2993,N_2985);
nand UO_51 (O_51,N_2988,N_2980);
xnor UO_52 (O_52,N_2980,N_2952);
xor UO_53 (O_53,N_2968,N_2969);
and UO_54 (O_54,N_2997,N_2959);
nor UO_55 (O_55,N_2950,N_2973);
or UO_56 (O_56,N_2975,N_2959);
xnor UO_57 (O_57,N_2976,N_2962);
and UO_58 (O_58,N_2983,N_2950);
nor UO_59 (O_59,N_2956,N_2973);
or UO_60 (O_60,N_2950,N_2975);
nor UO_61 (O_61,N_2958,N_2951);
nand UO_62 (O_62,N_2950,N_2986);
or UO_63 (O_63,N_2991,N_2990);
nor UO_64 (O_64,N_2959,N_2982);
nor UO_65 (O_65,N_2985,N_2994);
or UO_66 (O_66,N_2993,N_2990);
nor UO_67 (O_67,N_2967,N_2956);
nand UO_68 (O_68,N_2984,N_2998);
nand UO_69 (O_69,N_2968,N_2979);
nand UO_70 (O_70,N_2995,N_2963);
xnor UO_71 (O_71,N_2959,N_2979);
nand UO_72 (O_72,N_2972,N_2970);
nor UO_73 (O_73,N_2959,N_2998);
xnor UO_74 (O_74,N_2986,N_2983);
nor UO_75 (O_75,N_2966,N_2955);
and UO_76 (O_76,N_2999,N_2956);
and UO_77 (O_77,N_2973,N_2955);
and UO_78 (O_78,N_2998,N_2980);
nor UO_79 (O_79,N_2975,N_2984);
nor UO_80 (O_80,N_2961,N_2998);
and UO_81 (O_81,N_2968,N_2985);
nor UO_82 (O_82,N_2951,N_2962);
or UO_83 (O_83,N_2995,N_2970);
nand UO_84 (O_84,N_2963,N_2967);
or UO_85 (O_85,N_2978,N_2980);
nand UO_86 (O_86,N_2986,N_2958);
or UO_87 (O_87,N_2975,N_2999);
nor UO_88 (O_88,N_2959,N_2956);
xnor UO_89 (O_89,N_2993,N_2972);
nand UO_90 (O_90,N_2968,N_2988);
and UO_91 (O_91,N_2953,N_2984);
or UO_92 (O_92,N_2979,N_2985);
nand UO_93 (O_93,N_2951,N_2994);
nand UO_94 (O_94,N_2968,N_2963);
xnor UO_95 (O_95,N_2989,N_2963);
and UO_96 (O_96,N_2993,N_2986);
xnor UO_97 (O_97,N_2970,N_2961);
nor UO_98 (O_98,N_2963,N_2959);
and UO_99 (O_99,N_2983,N_2965);
xor UO_100 (O_100,N_2998,N_2979);
nand UO_101 (O_101,N_2952,N_2975);
and UO_102 (O_102,N_2990,N_2984);
nand UO_103 (O_103,N_2972,N_2981);
and UO_104 (O_104,N_2998,N_2994);
xor UO_105 (O_105,N_2956,N_2984);
nand UO_106 (O_106,N_2977,N_2994);
nor UO_107 (O_107,N_2976,N_2985);
and UO_108 (O_108,N_2968,N_2989);
nand UO_109 (O_109,N_2975,N_2962);
or UO_110 (O_110,N_2953,N_2978);
nor UO_111 (O_111,N_2962,N_2964);
nand UO_112 (O_112,N_2976,N_2958);
xor UO_113 (O_113,N_2957,N_2950);
xor UO_114 (O_114,N_2978,N_2993);
and UO_115 (O_115,N_2954,N_2970);
or UO_116 (O_116,N_2988,N_2964);
nand UO_117 (O_117,N_2977,N_2992);
or UO_118 (O_118,N_2987,N_2955);
nand UO_119 (O_119,N_2960,N_2999);
nand UO_120 (O_120,N_2984,N_2992);
xnor UO_121 (O_121,N_2999,N_2994);
nand UO_122 (O_122,N_2996,N_2957);
and UO_123 (O_123,N_2999,N_2977);
and UO_124 (O_124,N_2990,N_2957);
nor UO_125 (O_125,N_2987,N_2958);
or UO_126 (O_126,N_2984,N_2968);
or UO_127 (O_127,N_2966,N_2992);
nor UO_128 (O_128,N_2993,N_2983);
xnor UO_129 (O_129,N_2988,N_2971);
and UO_130 (O_130,N_2970,N_2953);
nand UO_131 (O_131,N_2963,N_2984);
or UO_132 (O_132,N_2952,N_2982);
nor UO_133 (O_133,N_2991,N_2961);
or UO_134 (O_134,N_2976,N_2984);
or UO_135 (O_135,N_2976,N_2986);
and UO_136 (O_136,N_2979,N_2956);
nor UO_137 (O_137,N_2955,N_2980);
nor UO_138 (O_138,N_2950,N_2954);
nand UO_139 (O_139,N_2962,N_2991);
and UO_140 (O_140,N_2997,N_2957);
nand UO_141 (O_141,N_2968,N_2954);
and UO_142 (O_142,N_2957,N_2969);
nand UO_143 (O_143,N_2955,N_2990);
xnor UO_144 (O_144,N_2972,N_2989);
and UO_145 (O_145,N_2999,N_2950);
nor UO_146 (O_146,N_2954,N_2959);
and UO_147 (O_147,N_2954,N_2985);
and UO_148 (O_148,N_2999,N_2974);
xor UO_149 (O_149,N_2985,N_2961);
nand UO_150 (O_150,N_2997,N_2987);
nor UO_151 (O_151,N_2956,N_2977);
nor UO_152 (O_152,N_2989,N_2996);
nand UO_153 (O_153,N_2973,N_2991);
xor UO_154 (O_154,N_2977,N_2978);
and UO_155 (O_155,N_2962,N_2997);
xnor UO_156 (O_156,N_2999,N_2969);
and UO_157 (O_157,N_2951,N_2991);
nor UO_158 (O_158,N_2963,N_2970);
nand UO_159 (O_159,N_2999,N_2988);
nor UO_160 (O_160,N_2996,N_2961);
or UO_161 (O_161,N_2991,N_2986);
nand UO_162 (O_162,N_2981,N_2986);
xnor UO_163 (O_163,N_2962,N_2973);
and UO_164 (O_164,N_2981,N_2963);
nand UO_165 (O_165,N_2990,N_2997);
nand UO_166 (O_166,N_2978,N_2955);
or UO_167 (O_167,N_2960,N_2996);
or UO_168 (O_168,N_2969,N_2958);
xor UO_169 (O_169,N_2992,N_2955);
xnor UO_170 (O_170,N_2959,N_2994);
nor UO_171 (O_171,N_2999,N_2958);
or UO_172 (O_172,N_2956,N_2953);
nand UO_173 (O_173,N_2956,N_2955);
and UO_174 (O_174,N_2965,N_2964);
nor UO_175 (O_175,N_2977,N_2968);
xnor UO_176 (O_176,N_2980,N_2951);
nor UO_177 (O_177,N_2996,N_2992);
or UO_178 (O_178,N_2954,N_2995);
nor UO_179 (O_179,N_2977,N_2975);
and UO_180 (O_180,N_2951,N_2998);
nand UO_181 (O_181,N_2982,N_2978);
nor UO_182 (O_182,N_2966,N_2993);
nor UO_183 (O_183,N_2975,N_2978);
nand UO_184 (O_184,N_2955,N_2970);
nand UO_185 (O_185,N_2957,N_2977);
nand UO_186 (O_186,N_2974,N_2958);
and UO_187 (O_187,N_2979,N_2954);
nand UO_188 (O_188,N_2971,N_2991);
nor UO_189 (O_189,N_2974,N_2983);
nor UO_190 (O_190,N_2957,N_2986);
and UO_191 (O_191,N_2956,N_2987);
xor UO_192 (O_192,N_2965,N_2975);
nor UO_193 (O_193,N_2992,N_2968);
nor UO_194 (O_194,N_2982,N_2997);
xnor UO_195 (O_195,N_2995,N_2957);
or UO_196 (O_196,N_2958,N_2962);
nor UO_197 (O_197,N_2978,N_2989);
nand UO_198 (O_198,N_2955,N_2960);
or UO_199 (O_199,N_2960,N_2951);
xnor UO_200 (O_200,N_2961,N_2993);
or UO_201 (O_201,N_2965,N_2985);
and UO_202 (O_202,N_2952,N_2951);
and UO_203 (O_203,N_2983,N_2988);
nor UO_204 (O_204,N_2956,N_2958);
and UO_205 (O_205,N_2983,N_2957);
and UO_206 (O_206,N_2958,N_2971);
nand UO_207 (O_207,N_2973,N_2978);
nand UO_208 (O_208,N_2970,N_2973);
and UO_209 (O_209,N_2995,N_2972);
nor UO_210 (O_210,N_2975,N_2992);
nor UO_211 (O_211,N_2986,N_2982);
nand UO_212 (O_212,N_2954,N_2989);
nor UO_213 (O_213,N_2963,N_2957);
or UO_214 (O_214,N_2979,N_2980);
xor UO_215 (O_215,N_2971,N_2995);
or UO_216 (O_216,N_2951,N_2986);
and UO_217 (O_217,N_2994,N_2970);
xnor UO_218 (O_218,N_2988,N_2985);
xor UO_219 (O_219,N_2952,N_2999);
nor UO_220 (O_220,N_2986,N_2969);
xnor UO_221 (O_221,N_2969,N_2993);
nor UO_222 (O_222,N_2991,N_2965);
and UO_223 (O_223,N_2981,N_2968);
nand UO_224 (O_224,N_2955,N_2999);
or UO_225 (O_225,N_2987,N_2959);
or UO_226 (O_226,N_2953,N_2976);
and UO_227 (O_227,N_2965,N_2966);
or UO_228 (O_228,N_2986,N_2980);
nor UO_229 (O_229,N_2987,N_2954);
and UO_230 (O_230,N_2997,N_2954);
nand UO_231 (O_231,N_2981,N_2989);
nor UO_232 (O_232,N_2950,N_2959);
nand UO_233 (O_233,N_2976,N_2973);
nand UO_234 (O_234,N_2967,N_2991);
and UO_235 (O_235,N_2961,N_2978);
and UO_236 (O_236,N_2983,N_2987);
and UO_237 (O_237,N_2950,N_2968);
or UO_238 (O_238,N_2958,N_2966);
or UO_239 (O_239,N_2981,N_2977);
and UO_240 (O_240,N_2996,N_2970);
nor UO_241 (O_241,N_2959,N_2995);
or UO_242 (O_242,N_2978,N_2954);
nor UO_243 (O_243,N_2967,N_2982);
nor UO_244 (O_244,N_2987,N_2979);
nand UO_245 (O_245,N_2992,N_2980);
and UO_246 (O_246,N_2972,N_2956);
nand UO_247 (O_247,N_2958,N_2977);
or UO_248 (O_248,N_2995,N_2965);
nor UO_249 (O_249,N_2950,N_2965);
xnor UO_250 (O_250,N_2993,N_2955);
xnor UO_251 (O_251,N_2963,N_2975);
nor UO_252 (O_252,N_2965,N_2980);
nand UO_253 (O_253,N_2972,N_2969);
nand UO_254 (O_254,N_2998,N_2965);
xor UO_255 (O_255,N_2981,N_2952);
or UO_256 (O_256,N_2984,N_2954);
or UO_257 (O_257,N_2983,N_2966);
and UO_258 (O_258,N_2981,N_2973);
and UO_259 (O_259,N_2959,N_2981);
or UO_260 (O_260,N_2989,N_2952);
nand UO_261 (O_261,N_2952,N_2964);
nor UO_262 (O_262,N_2952,N_2993);
and UO_263 (O_263,N_2966,N_2960);
nand UO_264 (O_264,N_2960,N_2976);
or UO_265 (O_265,N_2974,N_2972);
or UO_266 (O_266,N_2988,N_2955);
or UO_267 (O_267,N_2995,N_2980);
nor UO_268 (O_268,N_2967,N_2973);
nor UO_269 (O_269,N_2983,N_2990);
nor UO_270 (O_270,N_2971,N_2974);
and UO_271 (O_271,N_2959,N_2971);
and UO_272 (O_272,N_2987,N_2973);
xnor UO_273 (O_273,N_2962,N_2992);
xnor UO_274 (O_274,N_2961,N_2989);
xnor UO_275 (O_275,N_2956,N_2950);
xnor UO_276 (O_276,N_2964,N_2953);
or UO_277 (O_277,N_2962,N_2956);
nand UO_278 (O_278,N_2964,N_2993);
nor UO_279 (O_279,N_2952,N_2961);
nor UO_280 (O_280,N_2998,N_2983);
and UO_281 (O_281,N_2966,N_2962);
nand UO_282 (O_282,N_2960,N_2985);
nor UO_283 (O_283,N_2965,N_2958);
and UO_284 (O_284,N_2990,N_2961);
and UO_285 (O_285,N_2983,N_2976);
or UO_286 (O_286,N_2991,N_2977);
nor UO_287 (O_287,N_2958,N_2970);
and UO_288 (O_288,N_2968,N_2975);
or UO_289 (O_289,N_2976,N_2955);
nand UO_290 (O_290,N_2950,N_2970);
and UO_291 (O_291,N_2991,N_2989);
nor UO_292 (O_292,N_2982,N_2974);
xnor UO_293 (O_293,N_2980,N_2990);
nand UO_294 (O_294,N_2993,N_2981);
nand UO_295 (O_295,N_2988,N_2996);
or UO_296 (O_296,N_2971,N_2964);
and UO_297 (O_297,N_2980,N_2957);
or UO_298 (O_298,N_2976,N_2977);
xnor UO_299 (O_299,N_2963,N_2956);
and UO_300 (O_300,N_2961,N_2969);
nor UO_301 (O_301,N_2962,N_2957);
nand UO_302 (O_302,N_2986,N_2989);
nand UO_303 (O_303,N_2970,N_2982);
xor UO_304 (O_304,N_2954,N_2988);
xor UO_305 (O_305,N_2988,N_2972);
and UO_306 (O_306,N_2979,N_2953);
and UO_307 (O_307,N_2950,N_2996);
nor UO_308 (O_308,N_2971,N_2989);
xnor UO_309 (O_309,N_2983,N_2999);
xor UO_310 (O_310,N_2998,N_2977);
xnor UO_311 (O_311,N_2989,N_2969);
xnor UO_312 (O_312,N_2960,N_2994);
nor UO_313 (O_313,N_2978,N_2969);
nor UO_314 (O_314,N_2995,N_2975);
and UO_315 (O_315,N_2960,N_2971);
nand UO_316 (O_316,N_2997,N_2971);
or UO_317 (O_317,N_2994,N_2991);
nand UO_318 (O_318,N_2955,N_2997);
xnor UO_319 (O_319,N_2967,N_2960);
xor UO_320 (O_320,N_2973,N_2984);
or UO_321 (O_321,N_2991,N_2968);
nand UO_322 (O_322,N_2974,N_2955);
nand UO_323 (O_323,N_2995,N_2964);
and UO_324 (O_324,N_2964,N_2989);
and UO_325 (O_325,N_2960,N_2975);
nand UO_326 (O_326,N_2953,N_2996);
nand UO_327 (O_327,N_2985,N_2956);
xnor UO_328 (O_328,N_2980,N_2962);
nand UO_329 (O_329,N_2976,N_2999);
xnor UO_330 (O_330,N_2950,N_2990);
nand UO_331 (O_331,N_2963,N_2951);
or UO_332 (O_332,N_2996,N_2980);
nor UO_333 (O_333,N_2997,N_2974);
xor UO_334 (O_334,N_2959,N_2965);
or UO_335 (O_335,N_2974,N_2979);
xnor UO_336 (O_336,N_2975,N_2993);
xor UO_337 (O_337,N_2971,N_2956);
nor UO_338 (O_338,N_2974,N_2956);
nor UO_339 (O_339,N_2967,N_2975);
and UO_340 (O_340,N_2987,N_2976);
and UO_341 (O_341,N_2971,N_2950);
nor UO_342 (O_342,N_2983,N_2996);
or UO_343 (O_343,N_2987,N_2984);
nand UO_344 (O_344,N_2998,N_2969);
or UO_345 (O_345,N_2987,N_2992);
and UO_346 (O_346,N_2956,N_2965);
and UO_347 (O_347,N_2995,N_2967);
nor UO_348 (O_348,N_2988,N_2950);
xor UO_349 (O_349,N_2992,N_2967);
xnor UO_350 (O_350,N_2958,N_2983);
and UO_351 (O_351,N_2974,N_2998);
xor UO_352 (O_352,N_2970,N_2976);
nand UO_353 (O_353,N_2961,N_2966);
nor UO_354 (O_354,N_2985,N_2958);
and UO_355 (O_355,N_2957,N_2964);
or UO_356 (O_356,N_2965,N_2951);
or UO_357 (O_357,N_2951,N_2961);
and UO_358 (O_358,N_2995,N_2985);
and UO_359 (O_359,N_2967,N_2962);
and UO_360 (O_360,N_2975,N_2983);
nand UO_361 (O_361,N_2997,N_2989);
nand UO_362 (O_362,N_2961,N_2995);
nor UO_363 (O_363,N_2960,N_2995);
nand UO_364 (O_364,N_2981,N_2964);
and UO_365 (O_365,N_2953,N_2995);
nor UO_366 (O_366,N_2954,N_2981);
nand UO_367 (O_367,N_2950,N_2963);
nand UO_368 (O_368,N_2980,N_2981);
nor UO_369 (O_369,N_2951,N_2974);
and UO_370 (O_370,N_2973,N_2953);
and UO_371 (O_371,N_2959,N_2980);
nor UO_372 (O_372,N_2961,N_2950);
xnor UO_373 (O_373,N_2970,N_2951);
and UO_374 (O_374,N_2975,N_2973);
xnor UO_375 (O_375,N_2988,N_2998);
xor UO_376 (O_376,N_2989,N_2979);
and UO_377 (O_377,N_2962,N_2981);
nor UO_378 (O_378,N_2989,N_2960);
and UO_379 (O_379,N_2982,N_2998);
nand UO_380 (O_380,N_2969,N_2959);
nor UO_381 (O_381,N_2964,N_2992);
nor UO_382 (O_382,N_2971,N_2973);
or UO_383 (O_383,N_2990,N_2986);
nand UO_384 (O_384,N_2971,N_2980);
xnor UO_385 (O_385,N_2987,N_2967);
or UO_386 (O_386,N_2964,N_2951);
and UO_387 (O_387,N_2955,N_2971);
nand UO_388 (O_388,N_2991,N_2953);
nor UO_389 (O_389,N_2977,N_2954);
nand UO_390 (O_390,N_2971,N_2993);
nand UO_391 (O_391,N_2958,N_2955);
xnor UO_392 (O_392,N_2961,N_2984);
nand UO_393 (O_393,N_2974,N_2961);
nor UO_394 (O_394,N_2990,N_2981);
xor UO_395 (O_395,N_2960,N_2987);
xnor UO_396 (O_396,N_2973,N_2983);
or UO_397 (O_397,N_2989,N_2999);
nand UO_398 (O_398,N_2954,N_2951);
xnor UO_399 (O_399,N_2969,N_2981);
nor UO_400 (O_400,N_2951,N_2988);
xor UO_401 (O_401,N_2990,N_2973);
nor UO_402 (O_402,N_2980,N_2983);
nand UO_403 (O_403,N_2958,N_2993);
nor UO_404 (O_404,N_2979,N_2988);
nand UO_405 (O_405,N_2974,N_2965);
nand UO_406 (O_406,N_2984,N_2995);
xnor UO_407 (O_407,N_2984,N_2959);
and UO_408 (O_408,N_2953,N_2957);
and UO_409 (O_409,N_2978,N_2998);
nand UO_410 (O_410,N_2982,N_2971);
nor UO_411 (O_411,N_2961,N_2980);
xnor UO_412 (O_412,N_2992,N_2956);
nor UO_413 (O_413,N_2952,N_2958);
and UO_414 (O_414,N_2977,N_2993);
nor UO_415 (O_415,N_2960,N_2998);
nor UO_416 (O_416,N_2974,N_2976);
nand UO_417 (O_417,N_2962,N_2985);
nand UO_418 (O_418,N_2963,N_2979);
nand UO_419 (O_419,N_2988,N_2991);
and UO_420 (O_420,N_2995,N_2981);
and UO_421 (O_421,N_2997,N_2981);
nor UO_422 (O_422,N_2998,N_2972);
nor UO_423 (O_423,N_2954,N_2963);
nor UO_424 (O_424,N_2982,N_2965);
nand UO_425 (O_425,N_2950,N_2962);
and UO_426 (O_426,N_2969,N_2974);
nor UO_427 (O_427,N_2993,N_2996);
nor UO_428 (O_428,N_2977,N_2970);
xnor UO_429 (O_429,N_2999,N_2986);
nor UO_430 (O_430,N_2989,N_2995);
nand UO_431 (O_431,N_2957,N_2991);
or UO_432 (O_432,N_2966,N_2989);
and UO_433 (O_433,N_2978,N_2965);
nor UO_434 (O_434,N_2974,N_2957);
xor UO_435 (O_435,N_2978,N_2996);
or UO_436 (O_436,N_2984,N_2983);
or UO_437 (O_437,N_2967,N_2976);
nand UO_438 (O_438,N_2971,N_2978);
xnor UO_439 (O_439,N_2992,N_2994);
nand UO_440 (O_440,N_2999,N_2951);
xor UO_441 (O_441,N_2950,N_2989);
xor UO_442 (O_442,N_2982,N_2996);
and UO_443 (O_443,N_2959,N_2993);
nor UO_444 (O_444,N_2973,N_2959);
or UO_445 (O_445,N_2956,N_2978);
and UO_446 (O_446,N_2997,N_2963);
or UO_447 (O_447,N_2996,N_2995);
or UO_448 (O_448,N_2981,N_2991);
xor UO_449 (O_449,N_2979,N_2999);
nand UO_450 (O_450,N_2978,N_2995);
or UO_451 (O_451,N_2973,N_2963);
nor UO_452 (O_452,N_2965,N_2969);
or UO_453 (O_453,N_2966,N_2972);
and UO_454 (O_454,N_2990,N_2989);
xor UO_455 (O_455,N_2968,N_2967);
and UO_456 (O_456,N_2950,N_2951);
nand UO_457 (O_457,N_2970,N_2991);
nand UO_458 (O_458,N_2957,N_2972);
nor UO_459 (O_459,N_2996,N_2958);
and UO_460 (O_460,N_2950,N_2994);
or UO_461 (O_461,N_2991,N_2982);
and UO_462 (O_462,N_2970,N_2990);
and UO_463 (O_463,N_2974,N_2953);
nand UO_464 (O_464,N_2954,N_2960);
nor UO_465 (O_465,N_2951,N_2959);
nor UO_466 (O_466,N_2968,N_2960);
nor UO_467 (O_467,N_2974,N_2977);
or UO_468 (O_468,N_2976,N_2965);
nor UO_469 (O_469,N_2984,N_2970);
xor UO_470 (O_470,N_2994,N_2966);
and UO_471 (O_471,N_2979,N_2961);
xnor UO_472 (O_472,N_2958,N_2989);
or UO_473 (O_473,N_2978,N_2997);
and UO_474 (O_474,N_2995,N_2976);
xor UO_475 (O_475,N_2979,N_2951);
xor UO_476 (O_476,N_2958,N_2964);
xor UO_477 (O_477,N_2994,N_2963);
nor UO_478 (O_478,N_2998,N_2968);
nand UO_479 (O_479,N_2955,N_2951);
nor UO_480 (O_480,N_2952,N_2985);
xnor UO_481 (O_481,N_2969,N_2983);
xor UO_482 (O_482,N_2972,N_2955);
or UO_483 (O_483,N_2980,N_2964);
nor UO_484 (O_484,N_2960,N_2984);
and UO_485 (O_485,N_2973,N_2980);
nor UO_486 (O_486,N_2972,N_2986);
and UO_487 (O_487,N_2966,N_2963);
xnor UO_488 (O_488,N_2967,N_2999);
nor UO_489 (O_489,N_2978,N_2983);
nor UO_490 (O_490,N_2964,N_2999);
and UO_491 (O_491,N_2990,N_2954);
nor UO_492 (O_492,N_2964,N_2985);
xor UO_493 (O_493,N_2968,N_2982);
nor UO_494 (O_494,N_2994,N_2956);
xor UO_495 (O_495,N_2954,N_2957);
and UO_496 (O_496,N_2991,N_2992);
nand UO_497 (O_497,N_2963,N_2958);
or UO_498 (O_498,N_2999,N_2984);
and UO_499 (O_499,N_2987,N_2999);
endmodule