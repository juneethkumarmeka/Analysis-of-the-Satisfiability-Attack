module basic_750_5000_1000_10_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_347,In_407);
xnor U1 (N_1,In_205,In_148);
xnor U2 (N_2,In_312,In_482);
nor U3 (N_3,In_523,In_399);
and U4 (N_4,In_216,In_643);
xnor U5 (N_5,In_35,In_34);
xnor U6 (N_6,In_470,In_17);
or U7 (N_7,In_406,In_446);
or U8 (N_8,In_481,In_211);
nor U9 (N_9,In_129,In_542);
nor U10 (N_10,In_716,In_84);
nand U11 (N_11,In_280,In_311);
or U12 (N_12,In_702,In_251);
nor U13 (N_13,In_83,In_75);
nor U14 (N_14,In_387,In_108);
and U15 (N_15,In_241,In_263);
or U16 (N_16,In_398,In_372);
or U17 (N_17,In_171,In_541);
nor U18 (N_18,In_537,In_1);
or U19 (N_19,In_209,In_385);
nand U20 (N_20,In_32,In_690);
nor U21 (N_21,In_156,In_441);
or U22 (N_22,In_722,In_46);
xor U23 (N_23,In_103,In_87);
xor U24 (N_24,In_310,In_726);
xor U25 (N_25,In_400,In_730);
xor U26 (N_26,In_324,In_501);
nor U27 (N_27,In_498,In_160);
or U28 (N_28,In_326,In_689);
or U29 (N_29,In_141,In_25);
and U30 (N_30,In_601,In_612);
nand U31 (N_31,In_546,In_54);
nand U32 (N_32,In_193,In_40);
xnor U33 (N_33,In_710,In_414);
xor U34 (N_34,In_637,In_404);
xor U35 (N_35,In_717,In_262);
nand U36 (N_36,In_529,In_6);
nand U37 (N_37,In_439,In_272);
and U38 (N_38,In_465,In_195);
or U39 (N_39,In_668,In_673);
nor U40 (N_40,In_729,In_471);
nor U41 (N_41,In_639,In_433);
or U42 (N_42,In_686,In_685);
xnor U43 (N_43,In_519,In_238);
nor U44 (N_44,In_580,In_724);
nand U45 (N_45,In_602,In_342);
nand U46 (N_46,In_248,In_692);
nand U47 (N_47,In_436,In_506);
nor U48 (N_48,In_571,In_19);
and U49 (N_49,In_192,In_423);
and U50 (N_50,In_57,In_288);
nor U51 (N_51,In_58,In_588);
nand U52 (N_52,In_328,In_499);
xor U53 (N_53,In_666,In_239);
and U54 (N_54,In_510,In_53);
or U55 (N_55,In_101,In_178);
nand U56 (N_56,In_349,In_344);
xnor U57 (N_57,In_552,In_449);
nor U58 (N_58,In_67,In_247);
nor U59 (N_59,In_606,In_595);
and U60 (N_60,In_687,In_389);
and U61 (N_61,In_56,In_59);
nor U62 (N_62,In_187,In_151);
or U63 (N_63,In_120,In_382);
nor U64 (N_64,In_496,In_731);
xnor U65 (N_65,In_528,In_567);
xor U66 (N_66,In_380,In_313);
nand U67 (N_67,In_617,In_467);
and U68 (N_68,In_593,In_253);
xor U69 (N_69,In_170,In_268);
or U70 (N_70,In_144,In_719);
or U71 (N_71,In_503,In_627);
or U72 (N_72,In_577,In_426);
xnor U73 (N_73,In_275,In_116);
and U74 (N_74,In_424,In_374);
and U75 (N_75,In_37,In_462);
or U76 (N_76,In_409,In_284);
nand U77 (N_77,In_125,In_747);
nand U78 (N_78,In_479,In_740);
and U79 (N_79,In_508,In_51);
or U80 (N_80,In_712,In_442);
xor U81 (N_81,In_222,In_42);
nand U82 (N_82,In_381,In_278);
or U83 (N_83,In_444,In_106);
or U84 (N_84,In_30,In_180);
nand U85 (N_85,In_458,In_60);
or U86 (N_86,In_340,In_354);
or U87 (N_87,In_118,In_708);
and U88 (N_88,In_653,In_391);
xor U89 (N_89,In_491,In_212);
nor U90 (N_90,In_314,In_597);
nor U91 (N_91,In_361,In_276);
nor U92 (N_92,In_266,In_483);
nand U93 (N_93,In_675,In_24);
and U94 (N_94,In_49,In_246);
xnor U95 (N_95,In_664,In_565);
xnor U96 (N_96,In_111,In_680);
or U97 (N_97,In_319,In_723);
nand U98 (N_98,In_706,In_469);
or U99 (N_99,In_402,In_512);
and U100 (N_100,In_514,In_676);
and U101 (N_101,In_360,In_243);
xor U102 (N_102,In_656,In_375);
or U103 (N_103,In_448,In_438);
and U104 (N_104,In_581,In_614);
or U105 (N_105,In_226,In_590);
and U106 (N_106,In_245,In_478);
nand U107 (N_107,In_415,In_149);
and U108 (N_108,In_66,In_366);
and U109 (N_109,In_143,In_81);
nand U110 (N_110,In_392,In_383);
and U111 (N_111,In_490,In_718);
nor U112 (N_112,In_48,In_335);
xnor U113 (N_113,In_88,In_566);
or U114 (N_114,In_453,In_126);
nand U115 (N_115,In_123,In_74);
or U116 (N_116,In_488,In_713);
and U117 (N_117,In_397,In_329);
and U118 (N_118,In_408,In_511);
xnor U119 (N_119,In_269,In_667);
nor U120 (N_120,In_557,In_231);
and U121 (N_121,In_544,In_412);
nand U122 (N_122,In_330,In_715);
or U123 (N_123,In_283,In_620);
xor U124 (N_124,In_215,In_420);
or U125 (N_125,In_197,In_301);
nand U126 (N_126,In_64,In_474);
nand U127 (N_127,In_91,In_300);
and U128 (N_128,In_102,In_331);
nor U129 (N_129,In_658,In_682);
nor U130 (N_130,In_8,In_427);
or U131 (N_131,In_435,In_634);
and U132 (N_132,In_210,In_454);
or U133 (N_133,In_672,In_459);
or U134 (N_134,In_279,In_201);
xor U135 (N_135,In_316,In_534);
nand U136 (N_136,In_22,In_651);
xor U137 (N_137,In_332,In_703);
nor U138 (N_138,In_299,In_505);
xnor U139 (N_139,In_357,In_455);
and U140 (N_140,In_368,In_362);
xnor U141 (N_141,In_62,In_737);
xor U142 (N_142,In_36,In_353);
xnor U143 (N_143,In_677,In_486);
and U144 (N_144,In_237,In_377);
nor U145 (N_145,In_286,In_699);
nand U146 (N_146,In_630,In_256);
nor U147 (N_147,In_52,In_622);
and U148 (N_148,In_561,In_521);
xnor U149 (N_149,In_12,In_520);
xnor U150 (N_150,In_204,In_31);
or U151 (N_151,In_531,In_161);
or U152 (N_152,In_700,In_303);
nor U153 (N_153,In_670,In_198);
and U154 (N_154,In_738,In_683);
nor U155 (N_155,In_104,In_485);
and U156 (N_156,In_274,In_367);
xnor U157 (N_157,In_290,In_176);
and U158 (N_158,In_564,In_70);
or U159 (N_159,In_665,In_648);
or U160 (N_160,In_96,In_562);
and U161 (N_161,In_550,In_218);
nor U162 (N_162,In_135,In_475);
nor U163 (N_163,In_270,In_629);
nor U164 (N_164,In_646,In_321);
xor U165 (N_165,In_618,In_563);
or U166 (N_166,In_9,In_255);
xor U167 (N_167,In_749,In_364);
nand U168 (N_168,In_250,In_652);
xnor U169 (N_169,In_80,In_181);
xnor U170 (N_170,In_177,In_336);
nor U171 (N_171,In_99,In_466);
and U172 (N_172,In_277,In_242);
and U173 (N_173,In_356,In_191);
and U174 (N_174,In_492,In_282);
and U175 (N_175,In_139,In_572);
or U176 (N_176,In_741,In_662);
xnor U177 (N_177,In_227,In_421);
nor U178 (N_178,In_500,In_663);
nand U179 (N_179,In_203,In_232);
or U180 (N_180,In_184,In_234);
nor U181 (N_181,In_384,In_172);
nand U182 (N_182,In_616,In_405);
xnor U183 (N_183,In_432,In_76);
xnor U184 (N_184,In_431,In_480);
xnor U185 (N_185,In_39,In_655);
or U186 (N_186,In_654,In_249);
and U187 (N_187,In_320,In_14);
nor U188 (N_188,In_635,In_507);
and U189 (N_189,In_418,In_259);
or U190 (N_190,In_661,In_549);
nor U191 (N_191,In_18,In_701);
and U192 (N_192,In_569,In_173);
nand U193 (N_193,In_584,In_697);
nor U194 (N_194,In_355,In_124);
nor U195 (N_195,In_90,In_625);
or U196 (N_196,In_166,In_61);
and U197 (N_197,In_633,In_649);
nor U198 (N_198,In_113,In_709);
nand U199 (N_199,In_413,In_230);
nor U200 (N_200,In_307,In_711);
and U201 (N_201,In_285,In_305);
xor U202 (N_202,In_33,In_93);
and U203 (N_203,In_457,In_207);
nand U204 (N_204,In_146,In_681);
xor U205 (N_205,In_575,In_591);
xor U206 (N_206,In_348,In_164);
or U207 (N_207,In_744,In_189);
nand U208 (N_208,In_725,In_188);
or U209 (N_209,In_23,In_38);
and U210 (N_210,In_532,In_153);
or U211 (N_211,In_257,In_273);
nor U212 (N_212,In_609,In_742);
or U213 (N_213,In_97,In_621);
or U214 (N_214,In_174,In_105);
nor U215 (N_215,In_518,In_659);
and U216 (N_216,In_573,In_15);
nand U217 (N_217,In_114,In_167);
nand U218 (N_218,In_401,In_169);
or U219 (N_219,In_352,In_434);
xor U220 (N_220,In_592,In_261);
nand U221 (N_221,In_27,In_3);
and U222 (N_222,In_396,In_430);
xor U223 (N_223,In_502,In_628);
nor U224 (N_224,In_345,In_554);
and U225 (N_225,In_678,In_533);
or U226 (N_226,In_522,In_517);
or U227 (N_227,In_509,In_254);
xnor U228 (N_228,In_493,In_115);
xor U229 (N_229,In_460,In_746);
xor U230 (N_230,In_632,In_217);
xnor U231 (N_231,In_535,In_79);
nand U232 (N_232,In_732,In_315);
nor U233 (N_233,In_395,In_536);
or U234 (N_234,In_252,In_736);
and U235 (N_235,In_295,In_745);
and U236 (N_236,In_688,In_26);
and U237 (N_237,In_44,In_68);
and U238 (N_238,In_556,In_696);
nor U239 (N_239,In_147,In_271);
nand U240 (N_240,In_223,In_568);
nand U241 (N_241,In_7,In_570);
xor U242 (N_242,In_165,In_155);
or U243 (N_243,In_350,In_175);
nand U244 (N_244,In_162,In_267);
xor U245 (N_245,In_0,In_640);
or U246 (N_246,In_379,In_428);
nor U247 (N_247,In_596,In_43);
xnor U248 (N_248,In_309,In_393);
nor U249 (N_249,In_589,In_11);
nand U250 (N_250,In_89,In_369);
and U251 (N_251,In_186,In_497);
or U252 (N_252,In_464,In_647);
xor U253 (N_253,In_638,In_450);
or U254 (N_254,In_657,In_202);
or U255 (N_255,In_463,In_728);
nor U256 (N_256,In_194,In_206);
xor U257 (N_257,In_142,In_631);
xnor U258 (N_258,In_440,In_338);
and U259 (N_259,In_461,In_548);
nand U260 (N_260,In_425,In_45);
or U261 (N_261,In_671,In_323);
nand U262 (N_262,In_555,In_65);
xor U263 (N_263,In_137,In_733);
or U264 (N_264,In_626,In_513);
nor U265 (N_265,In_327,In_390);
xnor U266 (N_266,In_2,In_660);
nor U267 (N_267,In_574,In_322);
or U268 (N_268,In_610,In_587);
xor U269 (N_269,In_50,In_603);
nand U270 (N_270,In_585,In_473);
nor U271 (N_271,In_452,In_55);
or U272 (N_272,In_468,In_107);
or U273 (N_273,In_443,In_28);
or U274 (N_274,In_302,In_5);
and U275 (N_275,In_240,In_669);
nor U276 (N_276,In_644,In_705);
or U277 (N_277,In_553,In_200);
nor U278 (N_278,In_583,In_182);
nand U279 (N_279,In_526,In_339);
nand U280 (N_280,In_378,In_636);
or U281 (N_281,In_112,In_117);
and U282 (N_282,In_41,In_196);
nand U283 (N_283,In_29,In_403);
nand U284 (N_284,In_138,In_82);
or U285 (N_285,In_208,In_236);
nand U286 (N_286,In_333,In_394);
or U287 (N_287,In_297,In_641);
and U288 (N_288,In_152,In_346);
nand U289 (N_289,In_388,In_158);
nand U290 (N_290,In_605,In_410);
nor U291 (N_291,In_371,In_608);
nor U292 (N_292,In_219,In_698);
nand U293 (N_293,In_365,In_221);
or U294 (N_294,In_607,In_235);
or U295 (N_295,In_20,In_71);
or U296 (N_296,In_363,In_613);
or U297 (N_297,In_13,In_472);
xnor U298 (N_298,In_130,In_69);
or U299 (N_299,In_359,In_225);
nor U300 (N_300,In_695,In_586);
nand U301 (N_301,In_183,In_727);
nand U302 (N_302,In_539,In_748);
or U303 (N_303,In_411,In_264);
nor U304 (N_304,In_376,In_619);
or U305 (N_305,In_576,In_707);
or U306 (N_306,In_140,In_95);
nand U307 (N_307,In_373,In_445);
nand U308 (N_308,In_145,In_720);
or U309 (N_309,In_495,In_128);
nor U310 (N_310,In_296,In_150);
xor U311 (N_311,In_693,In_127);
and U312 (N_312,In_611,In_598);
xor U313 (N_313,In_624,In_704);
nand U314 (N_314,In_370,In_642);
nand U315 (N_315,In_298,In_265);
or U316 (N_316,In_220,In_4);
xnor U317 (N_317,In_419,In_122);
nand U318 (N_318,In_674,In_92);
nand U319 (N_319,In_47,In_163);
nand U320 (N_320,In_594,In_94);
or U321 (N_321,In_599,In_213);
xor U322 (N_322,In_98,In_615);
nor U323 (N_323,In_560,In_291);
or U324 (N_324,In_551,In_190);
nor U325 (N_325,In_429,In_734);
nand U326 (N_326,In_154,In_131);
nor U327 (N_327,In_86,In_527);
or U328 (N_328,In_386,In_487);
and U329 (N_329,In_159,In_524);
xnor U330 (N_330,In_179,In_294);
and U331 (N_331,In_735,In_292);
xor U332 (N_332,In_437,In_317);
nand U333 (N_333,In_489,In_229);
or U334 (N_334,In_358,In_228);
or U335 (N_335,In_306,In_281);
nor U336 (N_336,In_504,In_739);
nor U337 (N_337,In_224,In_287);
nand U338 (N_338,In_516,In_119);
xnor U339 (N_339,In_714,In_318);
nor U340 (N_340,In_477,In_258);
or U341 (N_341,In_85,In_417);
and U342 (N_342,In_78,In_545);
nor U343 (N_343,In_73,In_293);
or U344 (N_344,In_304,In_77);
xor U345 (N_345,In_559,In_494);
nor U346 (N_346,In_645,In_132);
nor U347 (N_347,In_341,In_16);
nand U348 (N_348,In_543,In_743);
nor U349 (N_349,In_456,In_558);
or U350 (N_350,In_600,In_63);
xor U351 (N_351,In_525,In_351);
nand U352 (N_352,In_133,In_110);
or U353 (N_353,In_260,In_308);
xnor U354 (N_354,In_289,In_579);
nand U355 (N_355,In_325,In_121);
xnor U356 (N_356,In_476,In_157);
or U357 (N_357,In_721,In_679);
nor U358 (N_358,In_10,In_582);
or U359 (N_359,In_233,In_214);
nor U360 (N_360,In_334,In_484);
nand U361 (N_361,In_604,In_540);
nand U362 (N_362,In_416,In_530);
nor U363 (N_363,In_650,In_694);
and U364 (N_364,In_451,In_515);
and U365 (N_365,In_72,In_168);
and U366 (N_366,In_691,In_623);
xor U367 (N_367,In_337,In_538);
and U368 (N_368,In_547,In_185);
or U369 (N_369,In_578,In_343);
nand U370 (N_370,In_136,In_447);
xor U371 (N_371,In_199,In_244);
and U372 (N_372,In_134,In_21);
nor U373 (N_373,In_422,In_100);
and U374 (N_374,In_109,In_684);
or U375 (N_375,In_546,In_622);
and U376 (N_376,In_67,In_519);
or U377 (N_377,In_59,In_468);
nor U378 (N_378,In_348,In_336);
nor U379 (N_379,In_624,In_463);
nand U380 (N_380,In_120,In_688);
or U381 (N_381,In_360,In_71);
and U382 (N_382,In_702,In_199);
nor U383 (N_383,In_463,In_312);
xor U384 (N_384,In_338,In_360);
nor U385 (N_385,In_448,In_741);
xor U386 (N_386,In_125,In_13);
nand U387 (N_387,In_97,In_739);
xor U388 (N_388,In_214,In_471);
nand U389 (N_389,In_227,In_625);
nor U390 (N_390,In_555,In_225);
nor U391 (N_391,In_253,In_26);
or U392 (N_392,In_28,In_392);
or U393 (N_393,In_101,In_538);
or U394 (N_394,In_7,In_314);
xor U395 (N_395,In_669,In_109);
and U396 (N_396,In_715,In_137);
nand U397 (N_397,In_357,In_259);
nor U398 (N_398,In_417,In_200);
nor U399 (N_399,In_407,In_132);
nand U400 (N_400,In_326,In_305);
and U401 (N_401,In_451,In_475);
nand U402 (N_402,In_403,In_226);
nand U403 (N_403,In_637,In_490);
xnor U404 (N_404,In_284,In_337);
nand U405 (N_405,In_223,In_729);
nand U406 (N_406,In_61,In_344);
nand U407 (N_407,In_0,In_429);
nand U408 (N_408,In_176,In_453);
xnor U409 (N_409,In_509,In_124);
nand U410 (N_410,In_616,In_481);
nor U411 (N_411,In_615,In_612);
nor U412 (N_412,In_279,In_269);
nor U413 (N_413,In_352,In_313);
nor U414 (N_414,In_718,In_418);
or U415 (N_415,In_247,In_622);
and U416 (N_416,In_275,In_469);
xnor U417 (N_417,In_149,In_89);
nand U418 (N_418,In_546,In_438);
and U419 (N_419,In_197,In_13);
and U420 (N_420,In_169,In_598);
and U421 (N_421,In_263,In_502);
xnor U422 (N_422,In_304,In_35);
and U423 (N_423,In_355,In_401);
and U424 (N_424,In_612,In_15);
or U425 (N_425,In_360,In_254);
nor U426 (N_426,In_158,In_113);
nand U427 (N_427,In_67,In_671);
nand U428 (N_428,In_595,In_173);
and U429 (N_429,In_4,In_344);
nand U430 (N_430,In_580,In_199);
and U431 (N_431,In_310,In_733);
nand U432 (N_432,In_688,In_730);
nor U433 (N_433,In_476,In_581);
nand U434 (N_434,In_256,In_310);
and U435 (N_435,In_465,In_108);
nor U436 (N_436,In_543,In_246);
xnor U437 (N_437,In_520,In_244);
and U438 (N_438,In_622,In_168);
nor U439 (N_439,In_577,In_19);
nand U440 (N_440,In_123,In_257);
xor U441 (N_441,In_438,In_185);
and U442 (N_442,In_738,In_14);
nand U443 (N_443,In_292,In_606);
and U444 (N_444,In_266,In_573);
nand U445 (N_445,In_659,In_399);
nand U446 (N_446,In_491,In_412);
and U447 (N_447,In_276,In_414);
nor U448 (N_448,In_606,In_371);
nor U449 (N_449,In_147,In_135);
and U450 (N_450,In_109,In_628);
or U451 (N_451,In_481,In_652);
or U452 (N_452,In_552,In_674);
nor U453 (N_453,In_583,In_298);
nand U454 (N_454,In_256,In_32);
xnor U455 (N_455,In_689,In_308);
nand U456 (N_456,In_292,In_298);
or U457 (N_457,In_122,In_691);
xnor U458 (N_458,In_596,In_483);
nand U459 (N_459,In_27,In_501);
nor U460 (N_460,In_561,In_724);
nor U461 (N_461,In_327,In_699);
xnor U462 (N_462,In_682,In_131);
xor U463 (N_463,In_711,In_133);
or U464 (N_464,In_173,In_92);
xnor U465 (N_465,In_618,In_692);
nand U466 (N_466,In_189,In_362);
or U467 (N_467,In_119,In_56);
or U468 (N_468,In_186,In_743);
or U469 (N_469,In_710,In_333);
nand U470 (N_470,In_685,In_176);
xor U471 (N_471,In_84,In_647);
or U472 (N_472,In_321,In_39);
nor U473 (N_473,In_461,In_734);
nor U474 (N_474,In_170,In_371);
and U475 (N_475,In_376,In_341);
xnor U476 (N_476,In_430,In_623);
nand U477 (N_477,In_696,In_170);
or U478 (N_478,In_423,In_223);
nor U479 (N_479,In_216,In_323);
or U480 (N_480,In_436,In_51);
and U481 (N_481,In_174,In_402);
xnor U482 (N_482,In_101,In_194);
nor U483 (N_483,In_401,In_737);
and U484 (N_484,In_6,In_191);
xnor U485 (N_485,In_67,In_683);
xor U486 (N_486,In_405,In_52);
nand U487 (N_487,In_442,In_410);
nand U488 (N_488,In_237,In_637);
and U489 (N_489,In_503,In_743);
or U490 (N_490,In_487,In_122);
nor U491 (N_491,In_75,In_270);
or U492 (N_492,In_237,In_388);
nor U493 (N_493,In_324,In_47);
nor U494 (N_494,In_553,In_379);
and U495 (N_495,In_545,In_590);
xor U496 (N_496,In_93,In_299);
xor U497 (N_497,In_579,In_571);
xnor U498 (N_498,In_40,In_565);
nor U499 (N_499,In_278,In_495);
nand U500 (N_500,N_425,N_201);
nor U501 (N_501,N_390,N_331);
xor U502 (N_502,N_463,N_89);
nand U503 (N_503,N_184,N_256);
and U504 (N_504,N_357,N_55);
and U505 (N_505,N_235,N_282);
nand U506 (N_506,N_494,N_56);
nor U507 (N_507,N_229,N_43);
nand U508 (N_508,N_105,N_400);
nand U509 (N_509,N_467,N_382);
xor U510 (N_510,N_372,N_413);
or U511 (N_511,N_140,N_130);
nand U512 (N_512,N_216,N_176);
nand U513 (N_513,N_471,N_335);
and U514 (N_514,N_198,N_220);
xnor U515 (N_515,N_320,N_142);
or U516 (N_516,N_383,N_394);
nor U517 (N_517,N_211,N_40);
or U518 (N_518,N_444,N_48);
nor U519 (N_519,N_202,N_294);
or U520 (N_520,N_241,N_173);
nor U521 (N_521,N_94,N_285);
and U522 (N_522,N_481,N_496);
or U523 (N_523,N_454,N_59);
nand U524 (N_524,N_364,N_412);
or U525 (N_525,N_106,N_486);
nor U526 (N_526,N_139,N_230);
nand U527 (N_527,N_146,N_458);
or U528 (N_528,N_380,N_87);
or U529 (N_529,N_245,N_278);
or U530 (N_530,N_460,N_189);
xor U531 (N_531,N_70,N_276);
and U532 (N_532,N_118,N_354);
nand U533 (N_533,N_293,N_416);
nand U534 (N_534,N_117,N_208);
or U535 (N_535,N_369,N_407);
xor U536 (N_536,N_295,N_150);
nand U537 (N_537,N_356,N_300);
and U538 (N_538,N_6,N_95);
nand U539 (N_539,N_258,N_313);
xnor U540 (N_540,N_397,N_341);
nor U541 (N_541,N_363,N_61);
and U542 (N_542,N_422,N_418);
nor U543 (N_543,N_327,N_482);
nand U544 (N_544,N_314,N_443);
xor U545 (N_545,N_339,N_274);
and U546 (N_546,N_451,N_286);
nand U547 (N_547,N_31,N_428);
and U548 (N_548,N_54,N_79);
xor U549 (N_549,N_232,N_238);
nor U550 (N_550,N_22,N_343);
xnor U551 (N_551,N_207,N_442);
xor U552 (N_552,N_495,N_392);
or U553 (N_553,N_99,N_464);
or U554 (N_554,N_69,N_4);
and U555 (N_555,N_361,N_309);
and U556 (N_556,N_26,N_161);
nand U557 (N_557,N_445,N_455);
nand U558 (N_558,N_476,N_132);
nor U559 (N_559,N_93,N_103);
and U560 (N_560,N_20,N_0);
xnor U561 (N_561,N_223,N_299);
and U562 (N_562,N_164,N_439);
nor U563 (N_563,N_109,N_315);
or U564 (N_564,N_127,N_65);
or U565 (N_565,N_209,N_166);
or U566 (N_566,N_264,N_144);
nand U567 (N_567,N_270,N_427);
nand U568 (N_568,N_218,N_57);
and U569 (N_569,N_108,N_1);
and U570 (N_570,N_206,N_483);
nand U571 (N_571,N_183,N_424);
xor U572 (N_572,N_280,N_462);
xnor U573 (N_573,N_91,N_178);
nand U574 (N_574,N_247,N_347);
or U575 (N_575,N_39,N_373);
nand U576 (N_576,N_15,N_171);
nor U577 (N_577,N_11,N_312);
nor U578 (N_578,N_461,N_302);
nand U579 (N_579,N_135,N_259);
nor U580 (N_580,N_113,N_37);
and U581 (N_581,N_440,N_352);
nand U582 (N_582,N_158,N_88);
xnor U583 (N_583,N_52,N_346);
nand U584 (N_584,N_194,N_355);
nand U585 (N_585,N_83,N_35);
nor U586 (N_586,N_466,N_30);
or U587 (N_587,N_449,N_136);
xor U588 (N_588,N_175,N_233);
xnor U589 (N_589,N_333,N_351);
and U590 (N_590,N_475,N_119);
xor U591 (N_591,N_47,N_401);
or U592 (N_592,N_155,N_226);
and U593 (N_593,N_435,N_367);
and U594 (N_594,N_237,N_303);
nor U595 (N_595,N_268,N_433);
or U596 (N_596,N_51,N_46);
nor U597 (N_597,N_254,N_344);
or U598 (N_598,N_212,N_485);
xnor U599 (N_599,N_114,N_358);
xor U600 (N_600,N_370,N_441);
or U601 (N_601,N_408,N_472);
nand U602 (N_602,N_298,N_214);
or U603 (N_603,N_44,N_159);
nand U604 (N_604,N_246,N_239);
xnor U605 (N_605,N_97,N_348);
nand U606 (N_606,N_228,N_17);
xor U607 (N_607,N_7,N_371);
nand U608 (N_608,N_430,N_253);
or U609 (N_609,N_38,N_126);
xor U610 (N_610,N_272,N_334);
nor U611 (N_611,N_321,N_337);
or U612 (N_612,N_250,N_14);
nor U613 (N_613,N_297,N_203);
or U614 (N_614,N_328,N_145);
or U615 (N_615,N_24,N_340);
xor U616 (N_616,N_167,N_62);
xnor U617 (N_617,N_498,N_169);
and U618 (N_618,N_307,N_499);
nor U619 (N_619,N_248,N_429);
xnor U620 (N_620,N_195,N_102);
or U621 (N_621,N_421,N_152);
and U622 (N_622,N_468,N_73);
or U623 (N_623,N_100,N_310);
nor U624 (N_624,N_411,N_205);
xor U625 (N_625,N_32,N_260);
nor U626 (N_626,N_116,N_359);
xnor U627 (N_627,N_234,N_275);
nor U628 (N_628,N_283,N_465);
nand U629 (N_629,N_279,N_375);
xnor U630 (N_630,N_185,N_188);
nor U631 (N_631,N_490,N_419);
xor U632 (N_632,N_23,N_165);
xor U633 (N_633,N_456,N_317);
or U634 (N_634,N_329,N_487);
or U635 (N_635,N_437,N_284);
nor U636 (N_636,N_410,N_33);
nand U637 (N_637,N_19,N_82);
nor U638 (N_638,N_148,N_72);
xnor U639 (N_639,N_269,N_18);
and U640 (N_640,N_409,N_292);
nand U641 (N_641,N_332,N_306);
or U642 (N_642,N_160,N_104);
and U643 (N_643,N_273,N_191);
or U644 (N_644,N_377,N_376);
xor U645 (N_645,N_395,N_21);
and U646 (N_646,N_385,N_389);
xnor U647 (N_647,N_8,N_244);
xor U648 (N_648,N_338,N_393);
nand U649 (N_649,N_53,N_265);
xnor U650 (N_650,N_289,N_81);
and U651 (N_651,N_174,N_42);
and U652 (N_652,N_342,N_252);
nand U653 (N_653,N_12,N_10);
nand U654 (N_654,N_484,N_489);
nor U655 (N_655,N_243,N_365);
nand U656 (N_656,N_379,N_177);
xor U657 (N_657,N_224,N_438);
or U658 (N_658,N_98,N_326);
and U659 (N_659,N_128,N_225);
xnor U660 (N_660,N_398,N_324);
xor U661 (N_661,N_50,N_141);
and U662 (N_662,N_151,N_316);
and U663 (N_663,N_196,N_34);
nor U664 (N_664,N_125,N_362);
xor U665 (N_665,N_448,N_101);
nor U666 (N_666,N_162,N_345);
nor U667 (N_667,N_107,N_213);
and U668 (N_668,N_63,N_488);
nand U669 (N_669,N_129,N_493);
or U670 (N_670,N_3,N_112);
or U671 (N_671,N_305,N_124);
or U672 (N_672,N_210,N_96);
and U673 (N_673,N_262,N_25);
xor U674 (N_674,N_450,N_193);
and U675 (N_675,N_49,N_68);
nor U676 (N_676,N_156,N_350);
xnor U677 (N_677,N_478,N_28);
nor U678 (N_678,N_222,N_479);
nand U679 (N_679,N_255,N_497);
and U680 (N_680,N_5,N_296);
or U681 (N_681,N_368,N_227);
and U682 (N_682,N_90,N_374);
and U683 (N_683,N_349,N_192);
nand U684 (N_684,N_287,N_41);
nor U685 (N_685,N_45,N_153);
and U686 (N_686,N_353,N_257);
and U687 (N_687,N_131,N_215);
nor U688 (N_688,N_491,N_120);
nor U689 (N_689,N_271,N_301);
nand U690 (N_690,N_381,N_71);
and U691 (N_691,N_423,N_122);
nor U692 (N_692,N_446,N_414);
nor U693 (N_693,N_66,N_304);
and U694 (N_694,N_182,N_434);
nand U695 (N_695,N_263,N_403);
nor U696 (N_696,N_76,N_74);
nand U697 (N_697,N_186,N_180);
or U698 (N_698,N_204,N_431);
nor U699 (N_699,N_134,N_84);
and U700 (N_700,N_154,N_447);
nor U701 (N_701,N_123,N_404);
and U702 (N_702,N_170,N_179);
nor U703 (N_703,N_322,N_457);
and U704 (N_704,N_366,N_149);
nor U705 (N_705,N_147,N_29);
or U706 (N_706,N_288,N_399);
nor U707 (N_707,N_281,N_402);
nand U708 (N_708,N_308,N_388);
xor U709 (N_709,N_330,N_453);
or U710 (N_710,N_78,N_384);
and U711 (N_711,N_217,N_323);
and U712 (N_712,N_406,N_311);
or U713 (N_713,N_240,N_415);
nand U714 (N_714,N_473,N_277);
xnor U715 (N_715,N_231,N_133);
and U716 (N_716,N_291,N_16);
xor U717 (N_717,N_236,N_290);
xnor U718 (N_718,N_378,N_432);
nor U719 (N_719,N_110,N_60);
and U720 (N_720,N_266,N_121);
nor U721 (N_721,N_85,N_426);
xnor U722 (N_722,N_477,N_436);
or U723 (N_723,N_172,N_9);
nand U724 (N_724,N_480,N_115);
and U725 (N_725,N_80,N_469);
nor U726 (N_726,N_386,N_181);
or U727 (N_727,N_242,N_138);
and U728 (N_728,N_219,N_470);
nand U729 (N_729,N_199,N_86);
nor U730 (N_730,N_163,N_221);
nor U731 (N_731,N_27,N_197);
nand U732 (N_732,N_249,N_452);
nand U733 (N_733,N_143,N_267);
xor U734 (N_734,N_92,N_111);
xor U735 (N_735,N_137,N_157);
nand U736 (N_736,N_474,N_387);
nand U737 (N_737,N_325,N_261);
and U738 (N_738,N_405,N_58);
and U739 (N_739,N_396,N_67);
and U740 (N_740,N_200,N_75);
or U741 (N_741,N_417,N_459);
or U742 (N_742,N_492,N_2);
nand U743 (N_743,N_420,N_360);
nor U744 (N_744,N_36,N_190);
nor U745 (N_745,N_318,N_187);
and U746 (N_746,N_391,N_64);
or U747 (N_747,N_77,N_251);
and U748 (N_748,N_319,N_336);
nand U749 (N_749,N_168,N_13);
nand U750 (N_750,N_19,N_359);
or U751 (N_751,N_19,N_441);
nand U752 (N_752,N_439,N_432);
or U753 (N_753,N_63,N_107);
xnor U754 (N_754,N_251,N_75);
nand U755 (N_755,N_389,N_300);
and U756 (N_756,N_181,N_257);
or U757 (N_757,N_206,N_217);
nand U758 (N_758,N_497,N_422);
or U759 (N_759,N_248,N_418);
and U760 (N_760,N_463,N_484);
and U761 (N_761,N_205,N_315);
nor U762 (N_762,N_121,N_192);
or U763 (N_763,N_237,N_25);
or U764 (N_764,N_164,N_204);
and U765 (N_765,N_167,N_207);
and U766 (N_766,N_268,N_212);
nand U767 (N_767,N_29,N_421);
nor U768 (N_768,N_309,N_244);
xor U769 (N_769,N_306,N_178);
and U770 (N_770,N_383,N_152);
and U771 (N_771,N_126,N_338);
or U772 (N_772,N_273,N_124);
nand U773 (N_773,N_297,N_166);
and U774 (N_774,N_48,N_356);
nand U775 (N_775,N_94,N_297);
xor U776 (N_776,N_331,N_444);
and U777 (N_777,N_351,N_94);
or U778 (N_778,N_75,N_33);
nor U779 (N_779,N_63,N_70);
nor U780 (N_780,N_267,N_144);
or U781 (N_781,N_85,N_408);
nand U782 (N_782,N_225,N_433);
xor U783 (N_783,N_403,N_82);
nor U784 (N_784,N_409,N_71);
nor U785 (N_785,N_251,N_182);
and U786 (N_786,N_447,N_450);
nor U787 (N_787,N_483,N_315);
or U788 (N_788,N_390,N_69);
or U789 (N_789,N_471,N_417);
and U790 (N_790,N_456,N_423);
and U791 (N_791,N_403,N_86);
nor U792 (N_792,N_448,N_275);
and U793 (N_793,N_232,N_441);
and U794 (N_794,N_440,N_222);
and U795 (N_795,N_475,N_420);
nor U796 (N_796,N_394,N_345);
nor U797 (N_797,N_108,N_100);
and U798 (N_798,N_296,N_34);
nor U799 (N_799,N_416,N_111);
nand U800 (N_800,N_384,N_89);
or U801 (N_801,N_14,N_365);
xnor U802 (N_802,N_367,N_345);
nand U803 (N_803,N_291,N_463);
nand U804 (N_804,N_142,N_241);
or U805 (N_805,N_147,N_126);
nor U806 (N_806,N_131,N_0);
xnor U807 (N_807,N_440,N_467);
nor U808 (N_808,N_144,N_26);
nor U809 (N_809,N_62,N_316);
nand U810 (N_810,N_289,N_157);
nand U811 (N_811,N_225,N_301);
nand U812 (N_812,N_327,N_13);
and U813 (N_813,N_244,N_495);
nor U814 (N_814,N_71,N_202);
nand U815 (N_815,N_165,N_266);
nor U816 (N_816,N_226,N_94);
xor U817 (N_817,N_433,N_132);
and U818 (N_818,N_53,N_24);
xor U819 (N_819,N_426,N_67);
or U820 (N_820,N_142,N_76);
xnor U821 (N_821,N_345,N_100);
and U822 (N_822,N_458,N_338);
or U823 (N_823,N_497,N_73);
and U824 (N_824,N_127,N_473);
nor U825 (N_825,N_134,N_64);
nand U826 (N_826,N_263,N_30);
nand U827 (N_827,N_397,N_35);
nand U828 (N_828,N_343,N_23);
nor U829 (N_829,N_145,N_109);
nor U830 (N_830,N_413,N_260);
nand U831 (N_831,N_187,N_307);
nor U832 (N_832,N_330,N_174);
or U833 (N_833,N_5,N_113);
or U834 (N_834,N_296,N_313);
nor U835 (N_835,N_314,N_259);
or U836 (N_836,N_17,N_207);
xnor U837 (N_837,N_255,N_296);
xnor U838 (N_838,N_302,N_132);
nor U839 (N_839,N_176,N_186);
or U840 (N_840,N_171,N_433);
nand U841 (N_841,N_38,N_237);
or U842 (N_842,N_316,N_39);
nand U843 (N_843,N_238,N_407);
and U844 (N_844,N_348,N_356);
and U845 (N_845,N_82,N_271);
nor U846 (N_846,N_119,N_138);
nor U847 (N_847,N_118,N_347);
and U848 (N_848,N_50,N_31);
nand U849 (N_849,N_52,N_213);
nor U850 (N_850,N_149,N_375);
nand U851 (N_851,N_450,N_89);
or U852 (N_852,N_382,N_435);
xor U853 (N_853,N_204,N_385);
and U854 (N_854,N_5,N_22);
and U855 (N_855,N_149,N_182);
nand U856 (N_856,N_106,N_184);
nand U857 (N_857,N_237,N_134);
or U858 (N_858,N_238,N_99);
and U859 (N_859,N_179,N_58);
nand U860 (N_860,N_361,N_154);
nand U861 (N_861,N_471,N_42);
nor U862 (N_862,N_165,N_380);
xnor U863 (N_863,N_345,N_26);
and U864 (N_864,N_27,N_479);
nor U865 (N_865,N_170,N_173);
xor U866 (N_866,N_316,N_391);
or U867 (N_867,N_87,N_178);
nand U868 (N_868,N_315,N_270);
xnor U869 (N_869,N_358,N_490);
nand U870 (N_870,N_300,N_333);
xnor U871 (N_871,N_172,N_265);
and U872 (N_872,N_219,N_38);
or U873 (N_873,N_68,N_16);
nor U874 (N_874,N_186,N_18);
and U875 (N_875,N_339,N_81);
nor U876 (N_876,N_432,N_435);
nand U877 (N_877,N_248,N_171);
xnor U878 (N_878,N_2,N_217);
nand U879 (N_879,N_427,N_299);
xor U880 (N_880,N_363,N_439);
nor U881 (N_881,N_403,N_270);
nand U882 (N_882,N_161,N_273);
nor U883 (N_883,N_67,N_250);
and U884 (N_884,N_54,N_17);
nor U885 (N_885,N_285,N_35);
nand U886 (N_886,N_2,N_255);
xor U887 (N_887,N_327,N_125);
and U888 (N_888,N_45,N_433);
and U889 (N_889,N_367,N_400);
xnor U890 (N_890,N_407,N_385);
nor U891 (N_891,N_206,N_410);
nand U892 (N_892,N_88,N_389);
xor U893 (N_893,N_450,N_50);
nor U894 (N_894,N_30,N_213);
and U895 (N_895,N_64,N_147);
or U896 (N_896,N_380,N_359);
and U897 (N_897,N_443,N_56);
xor U898 (N_898,N_245,N_493);
and U899 (N_899,N_154,N_368);
or U900 (N_900,N_284,N_5);
nor U901 (N_901,N_134,N_72);
nor U902 (N_902,N_491,N_183);
nor U903 (N_903,N_409,N_164);
or U904 (N_904,N_187,N_439);
nor U905 (N_905,N_466,N_368);
or U906 (N_906,N_438,N_280);
nand U907 (N_907,N_54,N_228);
nand U908 (N_908,N_374,N_300);
and U909 (N_909,N_3,N_422);
and U910 (N_910,N_66,N_333);
and U911 (N_911,N_60,N_34);
nand U912 (N_912,N_48,N_61);
nor U913 (N_913,N_401,N_168);
nor U914 (N_914,N_247,N_405);
nor U915 (N_915,N_294,N_94);
xor U916 (N_916,N_392,N_489);
or U917 (N_917,N_270,N_82);
nand U918 (N_918,N_84,N_204);
and U919 (N_919,N_353,N_398);
and U920 (N_920,N_7,N_353);
xnor U921 (N_921,N_388,N_327);
and U922 (N_922,N_482,N_138);
and U923 (N_923,N_83,N_130);
or U924 (N_924,N_173,N_289);
nand U925 (N_925,N_100,N_4);
nand U926 (N_926,N_388,N_448);
and U927 (N_927,N_382,N_267);
or U928 (N_928,N_215,N_227);
nand U929 (N_929,N_60,N_344);
nor U930 (N_930,N_59,N_155);
nand U931 (N_931,N_297,N_178);
xnor U932 (N_932,N_140,N_308);
and U933 (N_933,N_418,N_403);
xnor U934 (N_934,N_172,N_361);
and U935 (N_935,N_183,N_187);
nand U936 (N_936,N_191,N_383);
or U937 (N_937,N_120,N_401);
or U938 (N_938,N_438,N_316);
nor U939 (N_939,N_72,N_307);
and U940 (N_940,N_203,N_69);
xnor U941 (N_941,N_43,N_218);
and U942 (N_942,N_227,N_358);
xor U943 (N_943,N_170,N_41);
nand U944 (N_944,N_185,N_486);
and U945 (N_945,N_271,N_417);
nor U946 (N_946,N_402,N_290);
and U947 (N_947,N_2,N_27);
and U948 (N_948,N_493,N_377);
nand U949 (N_949,N_219,N_325);
and U950 (N_950,N_286,N_350);
nor U951 (N_951,N_37,N_489);
nor U952 (N_952,N_429,N_96);
nand U953 (N_953,N_395,N_145);
and U954 (N_954,N_362,N_363);
nand U955 (N_955,N_236,N_337);
and U956 (N_956,N_441,N_495);
nor U957 (N_957,N_401,N_260);
nor U958 (N_958,N_90,N_312);
xor U959 (N_959,N_221,N_412);
nor U960 (N_960,N_217,N_239);
nor U961 (N_961,N_259,N_223);
and U962 (N_962,N_22,N_151);
nor U963 (N_963,N_153,N_191);
nor U964 (N_964,N_173,N_357);
or U965 (N_965,N_12,N_257);
nor U966 (N_966,N_58,N_79);
and U967 (N_967,N_215,N_290);
nand U968 (N_968,N_416,N_169);
and U969 (N_969,N_166,N_39);
nand U970 (N_970,N_58,N_239);
and U971 (N_971,N_492,N_85);
nor U972 (N_972,N_98,N_432);
xor U973 (N_973,N_314,N_135);
xnor U974 (N_974,N_139,N_144);
xor U975 (N_975,N_329,N_144);
and U976 (N_976,N_240,N_142);
nand U977 (N_977,N_353,N_393);
xor U978 (N_978,N_182,N_197);
or U979 (N_979,N_125,N_305);
or U980 (N_980,N_178,N_0);
and U981 (N_981,N_216,N_482);
nand U982 (N_982,N_349,N_246);
nand U983 (N_983,N_466,N_369);
nor U984 (N_984,N_337,N_211);
nor U985 (N_985,N_384,N_477);
xor U986 (N_986,N_150,N_362);
nand U987 (N_987,N_217,N_356);
nor U988 (N_988,N_186,N_341);
and U989 (N_989,N_151,N_137);
nand U990 (N_990,N_248,N_257);
nand U991 (N_991,N_463,N_247);
xnor U992 (N_992,N_494,N_53);
nor U993 (N_993,N_241,N_299);
and U994 (N_994,N_154,N_250);
nor U995 (N_995,N_294,N_36);
and U996 (N_996,N_362,N_186);
xnor U997 (N_997,N_215,N_40);
and U998 (N_998,N_116,N_9);
or U999 (N_999,N_45,N_248);
and U1000 (N_1000,N_950,N_892);
nand U1001 (N_1001,N_941,N_986);
nor U1002 (N_1002,N_824,N_863);
or U1003 (N_1003,N_921,N_785);
nor U1004 (N_1004,N_981,N_911);
or U1005 (N_1005,N_775,N_508);
or U1006 (N_1006,N_881,N_586);
nand U1007 (N_1007,N_695,N_731);
xor U1008 (N_1008,N_673,N_700);
nand U1009 (N_1009,N_676,N_520);
or U1010 (N_1010,N_900,N_701);
and U1011 (N_1011,N_728,N_823);
nand U1012 (N_1012,N_766,N_947);
nor U1013 (N_1013,N_760,N_996);
nor U1014 (N_1014,N_524,N_562);
and U1015 (N_1015,N_968,N_674);
xor U1016 (N_1016,N_641,N_706);
and U1017 (N_1017,N_747,N_935);
and U1018 (N_1018,N_604,N_544);
nand U1019 (N_1019,N_737,N_710);
or U1020 (N_1020,N_519,N_540);
nand U1021 (N_1021,N_750,N_952);
xnor U1022 (N_1022,N_912,N_565);
or U1023 (N_1023,N_969,N_727);
nand U1024 (N_1024,N_790,N_847);
xor U1025 (N_1025,N_511,N_533);
or U1026 (N_1026,N_662,N_815);
or U1027 (N_1027,N_970,N_739);
xor U1028 (N_1028,N_705,N_738);
nand U1029 (N_1029,N_828,N_596);
xnor U1030 (N_1030,N_630,N_987);
xnor U1031 (N_1031,N_825,N_834);
nand U1032 (N_1032,N_749,N_769);
nand U1033 (N_1033,N_851,N_814);
nor U1034 (N_1034,N_504,N_580);
nor U1035 (N_1035,N_648,N_647);
xor U1036 (N_1036,N_835,N_751);
nand U1037 (N_1037,N_598,N_894);
xor U1038 (N_1038,N_726,N_839);
xnor U1039 (N_1039,N_628,N_669);
nor U1040 (N_1040,N_658,N_956);
xnor U1041 (N_1041,N_521,N_666);
xor U1042 (N_1042,N_649,N_548);
nor U1043 (N_1043,N_882,N_550);
xor U1044 (N_1044,N_840,N_682);
xor U1045 (N_1045,N_584,N_846);
xnor U1046 (N_1046,N_858,N_691);
nand U1047 (N_1047,N_717,N_998);
nor U1048 (N_1048,N_855,N_670);
or U1049 (N_1049,N_964,N_867);
and U1050 (N_1050,N_925,N_745);
or U1051 (N_1051,N_889,N_780);
and U1052 (N_1052,N_553,N_777);
nor U1053 (N_1053,N_665,N_595);
and U1054 (N_1054,N_594,N_612);
and U1055 (N_1055,N_686,N_767);
nand U1056 (N_1056,N_856,N_746);
xnor U1057 (N_1057,N_690,N_973);
xnor U1058 (N_1058,N_983,N_875);
nor U1059 (N_1059,N_714,N_923);
nand U1060 (N_1060,N_518,N_854);
and U1061 (N_1061,N_574,N_551);
xnor U1062 (N_1062,N_979,N_664);
nand U1063 (N_1063,N_978,N_868);
nand U1064 (N_1064,N_633,N_689);
or U1065 (N_1065,N_906,N_536);
or U1066 (N_1066,N_771,N_940);
nand U1067 (N_1067,N_933,N_954);
xor U1068 (N_1068,N_903,N_743);
xnor U1069 (N_1069,N_988,N_608);
or U1070 (N_1070,N_801,N_861);
xor U1071 (N_1071,N_937,N_784);
nor U1072 (N_1072,N_786,N_715);
or U1073 (N_1073,N_687,N_902);
or U1074 (N_1074,N_946,N_819);
nand U1075 (N_1075,N_585,N_898);
or U1076 (N_1076,N_837,N_927);
or U1077 (N_1077,N_614,N_741);
nor U1078 (N_1078,N_527,N_566);
xnor U1079 (N_1079,N_572,N_781);
or U1080 (N_1080,N_554,N_908);
xnor U1081 (N_1081,N_829,N_993);
nand U1082 (N_1082,N_953,N_799);
and U1083 (N_1083,N_713,N_939);
xnor U1084 (N_1084,N_958,N_995);
xor U1085 (N_1085,N_582,N_914);
or U1086 (N_1086,N_643,N_768);
xor U1087 (N_1087,N_859,N_545);
or U1088 (N_1088,N_600,N_619);
nor U1089 (N_1089,N_500,N_513);
xor U1090 (N_1090,N_560,N_629);
and U1091 (N_1091,N_822,N_593);
or U1092 (N_1092,N_721,N_677);
nand U1093 (N_1093,N_556,N_796);
or U1094 (N_1094,N_678,N_736);
or U1095 (N_1095,N_999,N_989);
nor U1096 (N_1096,N_878,N_934);
xnor U1097 (N_1097,N_729,N_657);
and U1098 (N_1098,N_755,N_510);
nand U1099 (N_1099,N_888,N_546);
nor U1100 (N_1100,N_871,N_588);
nand U1101 (N_1101,N_984,N_845);
xnor U1102 (N_1102,N_752,N_779);
xnor U1103 (N_1103,N_748,N_734);
nand U1104 (N_1104,N_803,N_931);
nand U1105 (N_1105,N_564,N_636);
xor U1106 (N_1106,N_764,N_797);
or U1107 (N_1107,N_971,N_506);
xnor U1108 (N_1108,N_756,N_836);
nor U1109 (N_1109,N_724,N_872);
nand U1110 (N_1110,N_622,N_592);
and U1111 (N_1111,N_758,N_907);
or U1112 (N_1112,N_638,N_735);
nand U1113 (N_1113,N_512,N_963);
and U1114 (N_1114,N_916,N_656);
nor U1115 (N_1115,N_708,N_639);
xnor U1116 (N_1116,N_770,N_928);
xnor U1117 (N_1117,N_692,N_936);
and U1118 (N_1118,N_555,N_515);
nand U1119 (N_1119,N_601,N_930);
xor U1120 (N_1120,N_891,N_826);
xor U1121 (N_1121,N_659,N_651);
and U1122 (N_1122,N_661,N_529);
or U1123 (N_1123,N_842,N_507);
nor U1124 (N_1124,N_722,N_757);
nor U1125 (N_1125,N_955,N_531);
xnor U1126 (N_1126,N_660,N_697);
xor U1127 (N_1127,N_509,N_617);
xnor U1128 (N_1128,N_597,N_838);
or U1129 (N_1129,N_578,N_631);
nand U1130 (N_1130,N_806,N_698);
xor U1131 (N_1131,N_704,N_563);
xnor U1132 (N_1132,N_541,N_609);
xor U1133 (N_1133,N_853,N_865);
xor U1134 (N_1134,N_547,N_812);
nand U1135 (N_1135,N_613,N_709);
or U1136 (N_1136,N_573,N_904);
or U1137 (N_1137,N_929,N_603);
nand U1138 (N_1138,N_577,N_793);
nor U1139 (N_1139,N_778,N_605);
nand U1140 (N_1140,N_849,N_794);
nand U1141 (N_1141,N_681,N_943);
and U1142 (N_1142,N_791,N_977);
nand U1143 (N_1143,N_589,N_542);
nor U1144 (N_1144,N_808,N_644);
or U1145 (N_1145,N_632,N_606);
or U1146 (N_1146,N_569,N_890);
nor U1147 (N_1147,N_517,N_762);
or U1148 (N_1148,N_528,N_850);
or U1149 (N_1149,N_831,N_537);
and U1150 (N_1150,N_693,N_707);
or U1151 (N_1151,N_730,N_844);
nor U1152 (N_1152,N_864,N_811);
and U1153 (N_1153,N_848,N_913);
nor U1154 (N_1154,N_539,N_897);
nand U1155 (N_1155,N_942,N_920);
or U1156 (N_1156,N_744,N_880);
or U1157 (N_1157,N_652,N_552);
nand U1158 (N_1158,N_821,N_945);
nand U1159 (N_1159,N_869,N_866);
nor U1160 (N_1160,N_841,N_774);
xnor U1161 (N_1161,N_980,N_813);
and U1162 (N_1162,N_602,N_718);
and U1163 (N_1163,N_966,N_830);
nor U1164 (N_1164,N_663,N_901);
or U1165 (N_1165,N_800,N_982);
or U1166 (N_1166,N_655,N_874);
nor U1167 (N_1167,N_761,N_616);
and U1168 (N_1168,N_623,N_514);
nand U1169 (N_1169,N_763,N_523);
nand U1170 (N_1170,N_772,N_792);
xor U1171 (N_1171,N_571,N_557);
and U1172 (N_1172,N_976,N_538);
and U1173 (N_1173,N_716,N_576);
xnor U1174 (N_1174,N_570,N_615);
or U1175 (N_1175,N_885,N_932);
xor U1176 (N_1176,N_587,N_625);
and U1177 (N_1177,N_759,N_675);
or U1178 (N_1178,N_962,N_640);
or U1179 (N_1179,N_627,N_960);
nand U1180 (N_1180,N_642,N_694);
nand U1181 (N_1181,N_702,N_820);
xnor U1182 (N_1182,N_985,N_918);
xor U1183 (N_1183,N_624,N_910);
nand U1184 (N_1184,N_862,N_575);
and U1185 (N_1185,N_883,N_719);
xor U1186 (N_1186,N_733,N_611);
xor U1187 (N_1187,N_668,N_712);
nor U1188 (N_1188,N_672,N_526);
or U1189 (N_1189,N_899,N_599);
nor U1190 (N_1190,N_650,N_637);
or U1191 (N_1191,N_591,N_967);
and U1192 (N_1192,N_787,N_620);
and U1193 (N_1193,N_997,N_558);
nor U1194 (N_1194,N_680,N_805);
xnor U1195 (N_1195,N_543,N_798);
xor U1196 (N_1196,N_503,N_974);
xnor U1197 (N_1197,N_684,N_991);
and U1198 (N_1198,N_505,N_893);
or U1199 (N_1199,N_568,N_919);
or U1200 (N_1200,N_896,N_688);
nand U1201 (N_1201,N_696,N_948);
nand U1202 (N_1202,N_534,N_961);
and U1203 (N_1203,N_938,N_817);
and U1204 (N_1204,N_549,N_809);
or U1205 (N_1205,N_559,N_501);
nor U1206 (N_1206,N_765,N_732);
or U1207 (N_1207,N_949,N_959);
xnor U1208 (N_1208,N_789,N_516);
or U1209 (N_1209,N_951,N_532);
nor U1210 (N_1210,N_754,N_990);
nor U1211 (N_1211,N_992,N_843);
xnor U1212 (N_1212,N_965,N_957);
nand U1213 (N_1213,N_788,N_646);
nor U1214 (N_1214,N_818,N_782);
xor U1215 (N_1215,N_567,N_667);
and U1216 (N_1216,N_645,N_804);
nor U1217 (N_1217,N_909,N_579);
nand U1218 (N_1218,N_530,N_924);
nand U1219 (N_1219,N_725,N_895);
nand U1220 (N_1220,N_583,N_525);
nand U1221 (N_1221,N_886,N_740);
xor U1222 (N_1222,N_753,N_635);
or U1223 (N_1223,N_502,N_610);
nor U1224 (N_1224,N_802,N_994);
xnor U1225 (N_1225,N_742,N_535);
and U1226 (N_1226,N_783,N_679);
nand U1227 (N_1227,N_723,N_877);
and U1228 (N_1228,N_522,N_876);
or U1229 (N_1229,N_654,N_773);
xor U1230 (N_1230,N_926,N_621);
and U1231 (N_1231,N_870,N_816);
or U1232 (N_1232,N_873,N_879);
xnor U1233 (N_1233,N_922,N_683);
or U1234 (N_1234,N_860,N_917);
nor U1235 (N_1235,N_972,N_699);
nand U1236 (N_1236,N_852,N_671);
nor U1237 (N_1237,N_810,N_703);
nor U1238 (N_1238,N_833,N_561);
and U1239 (N_1239,N_720,N_581);
or U1240 (N_1240,N_807,N_618);
or U1241 (N_1241,N_975,N_944);
and U1242 (N_1242,N_832,N_887);
or U1243 (N_1243,N_884,N_607);
and U1244 (N_1244,N_795,N_915);
or U1245 (N_1245,N_685,N_776);
and U1246 (N_1246,N_905,N_590);
or U1247 (N_1247,N_711,N_626);
or U1248 (N_1248,N_634,N_827);
xnor U1249 (N_1249,N_653,N_857);
and U1250 (N_1250,N_998,N_559);
nand U1251 (N_1251,N_874,N_693);
nand U1252 (N_1252,N_893,N_853);
and U1253 (N_1253,N_880,N_633);
nand U1254 (N_1254,N_670,N_992);
xor U1255 (N_1255,N_572,N_974);
and U1256 (N_1256,N_697,N_790);
nand U1257 (N_1257,N_696,N_705);
xor U1258 (N_1258,N_932,N_603);
nor U1259 (N_1259,N_695,N_679);
and U1260 (N_1260,N_642,N_853);
nand U1261 (N_1261,N_763,N_938);
nand U1262 (N_1262,N_562,N_823);
or U1263 (N_1263,N_784,N_969);
or U1264 (N_1264,N_649,N_990);
or U1265 (N_1265,N_857,N_922);
nand U1266 (N_1266,N_647,N_620);
and U1267 (N_1267,N_944,N_749);
or U1268 (N_1268,N_727,N_659);
nor U1269 (N_1269,N_592,N_727);
or U1270 (N_1270,N_598,N_905);
nand U1271 (N_1271,N_723,N_508);
xor U1272 (N_1272,N_537,N_708);
or U1273 (N_1273,N_806,N_545);
and U1274 (N_1274,N_850,N_712);
xnor U1275 (N_1275,N_527,N_858);
or U1276 (N_1276,N_523,N_518);
nand U1277 (N_1277,N_689,N_686);
nand U1278 (N_1278,N_509,N_829);
xnor U1279 (N_1279,N_517,N_813);
and U1280 (N_1280,N_778,N_733);
nor U1281 (N_1281,N_980,N_682);
or U1282 (N_1282,N_552,N_669);
xor U1283 (N_1283,N_582,N_526);
or U1284 (N_1284,N_565,N_902);
and U1285 (N_1285,N_780,N_813);
or U1286 (N_1286,N_506,N_810);
or U1287 (N_1287,N_806,N_870);
nor U1288 (N_1288,N_691,N_614);
or U1289 (N_1289,N_578,N_616);
or U1290 (N_1290,N_626,N_884);
nor U1291 (N_1291,N_680,N_621);
xnor U1292 (N_1292,N_896,N_639);
nor U1293 (N_1293,N_899,N_975);
nand U1294 (N_1294,N_734,N_866);
xor U1295 (N_1295,N_864,N_501);
nor U1296 (N_1296,N_808,N_914);
and U1297 (N_1297,N_770,N_613);
nor U1298 (N_1298,N_823,N_905);
or U1299 (N_1299,N_563,N_660);
nand U1300 (N_1300,N_992,N_706);
xor U1301 (N_1301,N_568,N_576);
and U1302 (N_1302,N_601,N_877);
and U1303 (N_1303,N_855,N_586);
or U1304 (N_1304,N_518,N_772);
or U1305 (N_1305,N_685,N_710);
or U1306 (N_1306,N_956,N_762);
nand U1307 (N_1307,N_697,N_724);
nand U1308 (N_1308,N_550,N_628);
xor U1309 (N_1309,N_520,N_703);
or U1310 (N_1310,N_640,N_789);
nor U1311 (N_1311,N_514,N_842);
or U1312 (N_1312,N_645,N_570);
or U1313 (N_1313,N_644,N_742);
or U1314 (N_1314,N_668,N_998);
or U1315 (N_1315,N_769,N_621);
xor U1316 (N_1316,N_711,N_553);
nand U1317 (N_1317,N_865,N_742);
or U1318 (N_1318,N_867,N_587);
xor U1319 (N_1319,N_720,N_910);
or U1320 (N_1320,N_847,N_987);
nand U1321 (N_1321,N_645,N_625);
nor U1322 (N_1322,N_937,N_875);
nor U1323 (N_1323,N_749,N_742);
and U1324 (N_1324,N_591,N_782);
or U1325 (N_1325,N_949,N_624);
and U1326 (N_1326,N_835,N_530);
and U1327 (N_1327,N_806,N_764);
and U1328 (N_1328,N_719,N_665);
nor U1329 (N_1329,N_556,N_826);
xnor U1330 (N_1330,N_968,N_850);
or U1331 (N_1331,N_699,N_903);
and U1332 (N_1332,N_841,N_915);
nand U1333 (N_1333,N_796,N_924);
or U1334 (N_1334,N_775,N_975);
nand U1335 (N_1335,N_915,N_692);
or U1336 (N_1336,N_974,N_665);
xnor U1337 (N_1337,N_660,N_528);
nand U1338 (N_1338,N_594,N_588);
nor U1339 (N_1339,N_855,N_663);
nand U1340 (N_1340,N_822,N_574);
xor U1341 (N_1341,N_898,N_915);
nand U1342 (N_1342,N_637,N_679);
nor U1343 (N_1343,N_533,N_928);
xor U1344 (N_1344,N_926,N_986);
and U1345 (N_1345,N_736,N_698);
nand U1346 (N_1346,N_954,N_590);
nor U1347 (N_1347,N_675,N_775);
xnor U1348 (N_1348,N_538,N_677);
and U1349 (N_1349,N_535,N_837);
nor U1350 (N_1350,N_956,N_782);
xor U1351 (N_1351,N_740,N_738);
and U1352 (N_1352,N_862,N_877);
and U1353 (N_1353,N_735,N_557);
nand U1354 (N_1354,N_687,N_569);
nor U1355 (N_1355,N_963,N_977);
xnor U1356 (N_1356,N_961,N_906);
nor U1357 (N_1357,N_927,N_508);
or U1358 (N_1358,N_665,N_672);
nand U1359 (N_1359,N_796,N_527);
nor U1360 (N_1360,N_710,N_693);
or U1361 (N_1361,N_790,N_738);
and U1362 (N_1362,N_866,N_873);
and U1363 (N_1363,N_705,N_708);
and U1364 (N_1364,N_767,N_782);
nor U1365 (N_1365,N_928,N_509);
or U1366 (N_1366,N_581,N_564);
or U1367 (N_1367,N_785,N_866);
nand U1368 (N_1368,N_628,N_632);
nand U1369 (N_1369,N_716,N_963);
xor U1370 (N_1370,N_698,N_674);
and U1371 (N_1371,N_606,N_562);
xor U1372 (N_1372,N_873,N_691);
xor U1373 (N_1373,N_815,N_961);
nand U1374 (N_1374,N_697,N_913);
and U1375 (N_1375,N_718,N_903);
nand U1376 (N_1376,N_687,N_700);
xor U1377 (N_1377,N_782,N_816);
nand U1378 (N_1378,N_547,N_817);
or U1379 (N_1379,N_985,N_823);
nand U1380 (N_1380,N_503,N_837);
and U1381 (N_1381,N_524,N_999);
xnor U1382 (N_1382,N_508,N_588);
and U1383 (N_1383,N_511,N_708);
xor U1384 (N_1384,N_819,N_849);
and U1385 (N_1385,N_572,N_854);
nor U1386 (N_1386,N_861,N_686);
and U1387 (N_1387,N_570,N_676);
nand U1388 (N_1388,N_584,N_875);
or U1389 (N_1389,N_801,N_901);
nand U1390 (N_1390,N_544,N_851);
nand U1391 (N_1391,N_821,N_769);
nand U1392 (N_1392,N_599,N_914);
or U1393 (N_1393,N_956,N_721);
or U1394 (N_1394,N_600,N_979);
nand U1395 (N_1395,N_881,N_716);
nand U1396 (N_1396,N_831,N_811);
and U1397 (N_1397,N_526,N_606);
nand U1398 (N_1398,N_980,N_519);
and U1399 (N_1399,N_568,N_932);
or U1400 (N_1400,N_764,N_837);
or U1401 (N_1401,N_683,N_841);
nand U1402 (N_1402,N_698,N_788);
nor U1403 (N_1403,N_890,N_555);
and U1404 (N_1404,N_620,N_649);
nor U1405 (N_1405,N_865,N_545);
nand U1406 (N_1406,N_875,N_508);
nand U1407 (N_1407,N_791,N_982);
xnor U1408 (N_1408,N_934,N_883);
or U1409 (N_1409,N_882,N_830);
nor U1410 (N_1410,N_541,N_561);
nand U1411 (N_1411,N_828,N_509);
and U1412 (N_1412,N_941,N_764);
nor U1413 (N_1413,N_873,N_658);
nor U1414 (N_1414,N_645,N_618);
nand U1415 (N_1415,N_790,N_834);
nor U1416 (N_1416,N_876,N_826);
nand U1417 (N_1417,N_925,N_561);
or U1418 (N_1418,N_848,N_505);
nor U1419 (N_1419,N_911,N_957);
nor U1420 (N_1420,N_547,N_666);
xor U1421 (N_1421,N_938,N_772);
nand U1422 (N_1422,N_552,N_845);
nand U1423 (N_1423,N_700,N_838);
nand U1424 (N_1424,N_583,N_608);
xor U1425 (N_1425,N_895,N_647);
nand U1426 (N_1426,N_851,N_703);
xor U1427 (N_1427,N_794,N_784);
or U1428 (N_1428,N_748,N_666);
xor U1429 (N_1429,N_912,N_654);
or U1430 (N_1430,N_702,N_519);
xor U1431 (N_1431,N_778,N_630);
nand U1432 (N_1432,N_646,N_919);
and U1433 (N_1433,N_526,N_629);
or U1434 (N_1434,N_556,N_655);
xor U1435 (N_1435,N_955,N_583);
or U1436 (N_1436,N_687,N_608);
or U1437 (N_1437,N_650,N_669);
and U1438 (N_1438,N_880,N_948);
nand U1439 (N_1439,N_752,N_977);
xnor U1440 (N_1440,N_955,N_730);
nand U1441 (N_1441,N_986,N_703);
and U1442 (N_1442,N_778,N_658);
xnor U1443 (N_1443,N_939,N_651);
nand U1444 (N_1444,N_599,N_542);
nor U1445 (N_1445,N_716,N_908);
nand U1446 (N_1446,N_520,N_985);
nor U1447 (N_1447,N_756,N_658);
nor U1448 (N_1448,N_509,N_565);
or U1449 (N_1449,N_608,N_501);
nor U1450 (N_1450,N_697,N_882);
nand U1451 (N_1451,N_645,N_888);
or U1452 (N_1452,N_759,N_509);
nand U1453 (N_1453,N_760,N_958);
xor U1454 (N_1454,N_730,N_770);
xnor U1455 (N_1455,N_762,N_931);
xor U1456 (N_1456,N_729,N_594);
nand U1457 (N_1457,N_726,N_795);
and U1458 (N_1458,N_910,N_593);
and U1459 (N_1459,N_561,N_799);
nand U1460 (N_1460,N_504,N_930);
or U1461 (N_1461,N_770,N_965);
or U1462 (N_1462,N_915,N_875);
nor U1463 (N_1463,N_531,N_897);
or U1464 (N_1464,N_718,N_591);
nand U1465 (N_1465,N_979,N_528);
nand U1466 (N_1466,N_948,N_563);
or U1467 (N_1467,N_694,N_625);
xnor U1468 (N_1468,N_968,N_846);
nand U1469 (N_1469,N_669,N_994);
nor U1470 (N_1470,N_997,N_830);
or U1471 (N_1471,N_912,N_553);
nand U1472 (N_1472,N_791,N_900);
and U1473 (N_1473,N_623,N_710);
nand U1474 (N_1474,N_974,N_760);
and U1475 (N_1475,N_631,N_901);
nand U1476 (N_1476,N_642,N_784);
nor U1477 (N_1477,N_602,N_836);
or U1478 (N_1478,N_906,N_528);
xnor U1479 (N_1479,N_526,N_624);
nor U1480 (N_1480,N_779,N_863);
xor U1481 (N_1481,N_940,N_697);
nor U1482 (N_1482,N_682,N_695);
nand U1483 (N_1483,N_965,N_524);
xor U1484 (N_1484,N_626,N_713);
and U1485 (N_1485,N_854,N_593);
xor U1486 (N_1486,N_863,N_930);
nand U1487 (N_1487,N_641,N_521);
nand U1488 (N_1488,N_767,N_674);
nor U1489 (N_1489,N_909,N_873);
nand U1490 (N_1490,N_720,N_644);
nor U1491 (N_1491,N_908,N_782);
nor U1492 (N_1492,N_634,N_818);
or U1493 (N_1493,N_614,N_912);
xor U1494 (N_1494,N_523,N_820);
and U1495 (N_1495,N_836,N_802);
or U1496 (N_1496,N_741,N_697);
and U1497 (N_1497,N_928,N_781);
xnor U1498 (N_1498,N_849,N_771);
and U1499 (N_1499,N_680,N_686);
nand U1500 (N_1500,N_1232,N_1160);
nand U1501 (N_1501,N_1279,N_1294);
xor U1502 (N_1502,N_1375,N_1283);
nand U1503 (N_1503,N_1423,N_1034);
xor U1504 (N_1504,N_1201,N_1449);
nor U1505 (N_1505,N_1311,N_1139);
nand U1506 (N_1506,N_1257,N_1255);
and U1507 (N_1507,N_1024,N_1284);
xor U1508 (N_1508,N_1282,N_1061);
nand U1509 (N_1509,N_1421,N_1238);
nor U1510 (N_1510,N_1137,N_1098);
xnor U1511 (N_1511,N_1356,N_1253);
and U1512 (N_1512,N_1101,N_1230);
xnor U1513 (N_1513,N_1393,N_1179);
or U1514 (N_1514,N_1142,N_1207);
and U1515 (N_1515,N_1145,N_1310);
xnor U1516 (N_1516,N_1005,N_1026);
xor U1517 (N_1517,N_1380,N_1184);
and U1518 (N_1518,N_1397,N_1196);
nor U1519 (N_1519,N_1409,N_1116);
and U1520 (N_1520,N_1468,N_1267);
or U1521 (N_1521,N_1308,N_1008);
or U1522 (N_1522,N_1335,N_1086);
or U1523 (N_1523,N_1062,N_1228);
nand U1524 (N_1524,N_1293,N_1346);
xnor U1525 (N_1525,N_1241,N_1334);
or U1526 (N_1526,N_1129,N_1268);
nand U1527 (N_1527,N_1149,N_1189);
and U1528 (N_1528,N_1432,N_1474);
nor U1529 (N_1529,N_1254,N_1373);
or U1530 (N_1530,N_1491,N_1433);
and U1531 (N_1531,N_1422,N_1464);
xor U1532 (N_1532,N_1322,N_1091);
or U1533 (N_1533,N_1042,N_1394);
or U1534 (N_1534,N_1362,N_1389);
xor U1535 (N_1535,N_1437,N_1262);
nand U1536 (N_1536,N_1195,N_1066);
xor U1537 (N_1537,N_1001,N_1047);
nand U1538 (N_1538,N_1332,N_1471);
and U1539 (N_1539,N_1320,N_1014);
or U1540 (N_1540,N_1285,N_1203);
and U1541 (N_1541,N_1440,N_1004);
and U1542 (N_1542,N_1465,N_1469);
or U1543 (N_1543,N_1260,N_1043);
nor U1544 (N_1544,N_1456,N_1118);
xor U1545 (N_1545,N_1455,N_1426);
xnor U1546 (N_1546,N_1068,N_1109);
nand U1547 (N_1547,N_1256,N_1488);
or U1548 (N_1548,N_1172,N_1171);
nor U1549 (N_1549,N_1300,N_1457);
nand U1550 (N_1550,N_1476,N_1462);
and U1551 (N_1551,N_1038,N_1057);
or U1552 (N_1552,N_1286,N_1071);
nand U1553 (N_1553,N_1099,N_1336);
nor U1554 (N_1554,N_1127,N_1446);
nor U1555 (N_1555,N_1454,N_1208);
nand U1556 (N_1556,N_1291,N_1309);
nor U1557 (N_1557,N_1002,N_1448);
or U1558 (N_1558,N_1401,N_1095);
nand U1559 (N_1559,N_1176,N_1221);
nand U1560 (N_1560,N_1453,N_1178);
or U1561 (N_1561,N_1242,N_1417);
and U1562 (N_1562,N_1399,N_1411);
nand U1563 (N_1563,N_1390,N_1317);
nor U1564 (N_1564,N_1094,N_1213);
or U1565 (N_1565,N_1050,N_1313);
xnor U1566 (N_1566,N_1261,N_1202);
and U1567 (N_1567,N_1191,N_1133);
and U1568 (N_1568,N_1022,N_1297);
or U1569 (N_1569,N_1188,N_1111);
nor U1570 (N_1570,N_1359,N_1036);
nor U1571 (N_1571,N_1117,N_1307);
and U1572 (N_1572,N_1248,N_1106);
or U1573 (N_1573,N_1452,N_1429);
xnor U1574 (N_1574,N_1377,N_1447);
nand U1575 (N_1575,N_1156,N_1170);
or U1576 (N_1576,N_1342,N_1020);
xor U1577 (N_1577,N_1444,N_1326);
nand U1578 (N_1578,N_1089,N_1372);
or U1579 (N_1579,N_1150,N_1466);
nand U1580 (N_1580,N_1030,N_1358);
or U1581 (N_1581,N_1143,N_1110);
and U1582 (N_1582,N_1306,N_1288);
nand U1583 (N_1583,N_1384,N_1271);
and U1584 (N_1584,N_1367,N_1054);
and U1585 (N_1585,N_1000,N_1475);
and U1586 (N_1586,N_1371,N_1124);
and U1587 (N_1587,N_1410,N_1161);
and U1588 (N_1588,N_1439,N_1220);
or U1589 (N_1589,N_1169,N_1056);
nand U1590 (N_1590,N_1460,N_1263);
nor U1591 (N_1591,N_1090,N_1425);
nor U1592 (N_1592,N_1274,N_1481);
or U1593 (N_1593,N_1374,N_1205);
or U1594 (N_1594,N_1214,N_1197);
and U1595 (N_1595,N_1325,N_1082);
or U1596 (N_1596,N_1032,N_1360);
xor U1597 (N_1597,N_1289,N_1236);
nor U1598 (N_1598,N_1391,N_1340);
nor U1599 (N_1599,N_1102,N_1158);
nand U1600 (N_1600,N_1212,N_1219);
and U1601 (N_1601,N_1199,N_1079);
xnor U1602 (N_1602,N_1107,N_1244);
or U1603 (N_1603,N_1281,N_1157);
or U1604 (N_1604,N_1459,N_1187);
or U1605 (N_1605,N_1120,N_1035);
nor U1606 (N_1606,N_1364,N_1315);
xnor U1607 (N_1607,N_1412,N_1060);
nor U1608 (N_1608,N_1162,N_1361);
and U1609 (N_1609,N_1163,N_1108);
nor U1610 (N_1610,N_1470,N_1173);
or U1611 (N_1611,N_1251,N_1318);
or U1612 (N_1612,N_1381,N_1063);
nor U1613 (N_1613,N_1119,N_1302);
nor U1614 (N_1614,N_1324,N_1065);
xor U1615 (N_1615,N_1216,N_1418);
nor U1616 (N_1616,N_1458,N_1339);
nor U1617 (N_1617,N_1200,N_1328);
xor U1618 (N_1618,N_1085,N_1100);
nand U1619 (N_1619,N_1303,N_1442);
nand U1620 (N_1620,N_1338,N_1366);
or U1621 (N_1621,N_1369,N_1175);
and U1622 (N_1622,N_1217,N_1105);
nand U1623 (N_1623,N_1019,N_1227);
or U1624 (N_1624,N_1441,N_1070);
or U1625 (N_1625,N_1438,N_1273);
nor U1626 (N_1626,N_1155,N_1134);
or U1627 (N_1627,N_1296,N_1017);
xor U1628 (N_1628,N_1074,N_1400);
nor U1629 (N_1629,N_1445,N_1420);
nor U1630 (N_1630,N_1395,N_1353);
xnor U1631 (N_1631,N_1270,N_1486);
and U1632 (N_1632,N_1333,N_1323);
nor U1633 (N_1633,N_1136,N_1477);
and U1634 (N_1634,N_1473,N_1180);
nor U1635 (N_1635,N_1235,N_1088);
xor U1636 (N_1636,N_1121,N_1144);
nand U1637 (N_1637,N_1276,N_1352);
nand U1638 (N_1638,N_1392,N_1246);
nor U1639 (N_1639,N_1048,N_1402);
or U1640 (N_1640,N_1405,N_1018);
xnor U1641 (N_1641,N_1430,N_1113);
nor U1642 (N_1642,N_1093,N_1037);
xnor U1643 (N_1643,N_1015,N_1168);
nor U1644 (N_1644,N_1406,N_1316);
or U1645 (N_1645,N_1206,N_1354);
and U1646 (N_1646,N_1349,N_1097);
or U1647 (N_1647,N_1436,N_1275);
nand U1648 (N_1648,N_1039,N_1130);
nand U1649 (N_1649,N_1321,N_1029);
nor U1650 (N_1650,N_1081,N_1419);
nand U1651 (N_1651,N_1427,N_1450);
nand U1652 (N_1652,N_1278,N_1343);
xor U1653 (N_1653,N_1483,N_1495);
nor U1654 (N_1654,N_1041,N_1479);
or U1655 (N_1655,N_1148,N_1166);
and U1656 (N_1656,N_1415,N_1104);
and U1657 (N_1657,N_1290,N_1482);
and U1658 (N_1658,N_1478,N_1264);
or U1659 (N_1659,N_1295,N_1341);
xor U1660 (N_1660,N_1265,N_1126);
or U1661 (N_1661,N_1087,N_1379);
nand U1662 (N_1662,N_1499,N_1234);
and U1663 (N_1663,N_1186,N_1141);
xor U1664 (N_1664,N_1193,N_1027);
nor U1665 (N_1665,N_1301,N_1407);
nor U1666 (N_1666,N_1078,N_1492);
nor U1667 (N_1667,N_1073,N_1040);
xor U1668 (N_1668,N_1204,N_1329);
nand U1669 (N_1669,N_1434,N_1092);
nor U1670 (N_1670,N_1226,N_1348);
xnor U1671 (N_1671,N_1028,N_1122);
nand U1672 (N_1672,N_1055,N_1404);
or U1673 (N_1673,N_1327,N_1490);
nor U1674 (N_1674,N_1387,N_1239);
nand U1675 (N_1675,N_1125,N_1123);
xor U1676 (N_1676,N_1077,N_1132);
xor U1677 (N_1677,N_1215,N_1331);
nor U1678 (N_1678,N_1167,N_1233);
xor U1679 (N_1679,N_1031,N_1461);
xnor U1680 (N_1680,N_1319,N_1185);
xnor U1681 (N_1681,N_1064,N_1210);
nor U1682 (N_1682,N_1006,N_1051);
and U1683 (N_1683,N_1067,N_1272);
nand U1684 (N_1684,N_1467,N_1059);
nand U1685 (N_1685,N_1231,N_1192);
xor U1686 (N_1686,N_1140,N_1007);
nor U1687 (N_1687,N_1218,N_1223);
and U1688 (N_1688,N_1045,N_1046);
and U1689 (N_1689,N_1131,N_1003);
xnor U1690 (N_1690,N_1096,N_1396);
nor U1691 (N_1691,N_1484,N_1194);
nor U1692 (N_1692,N_1128,N_1330);
nand U1693 (N_1693,N_1365,N_1266);
and U1694 (N_1694,N_1382,N_1388);
nand U1695 (N_1695,N_1198,N_1351);
nor U1696 (N_1696,N_1414,N_1135);
nand U1697 (N_1697,N_1152,N_1069);
nor U1698 (N_1698,N_1428,N_1280);
nand U1699 (N_1699,N_1368,N_1181);
nor U1700 (N_1700,N_1190,N_1012);
nor U1701 (N_1701,N_1451,N_1165);
nand U1702 (N_1702,N_1370,N_1347);
and U1703 (N_1703,N_1084,N_1403);
or U1704 (N_1704,N_1416,N_1072);
or U1705 (N_1705,N_1016,N_1463);
nor U1706 (N_1706,N_1487,N_1304);
nand U1707 (N_1707,N_1378,N_1269);
nor U1708 (N_1708,N_1258,N_1112);
nand U1709 (N_1709,N_1224,N_1247);
or U1710 (N_1710,N_1376,N_1115);
and U1711 (N_1711,N_1277,N_1147);
nand U1712 (N_1712,N_1496,N_1146);
xor U1713 (N_1713,N_1010,N_1252);
nor U1714 (N_1714,N_1497,N_1314);
and U1715 (N_1715,N_1485,N_1080);
and U1716 (N_1716,N_1498,N_1209);
and U1717 (N_1717,N_1183,N_1211);
xor U1718 (N_1718,N_1052,N_1493);
nor U1719 (N_1719,N_1025,N_1049);
xor U1720 (N_1720,N_1250,N_1259);
or U1721 (N_1721,N_1355,N_1413);
nand U1722 (N_1722,N_1229,N_1103);
nor U1723 (N_1723,N_1058,N_1114);
nor U1724 (N_1724,N_1177,N_1305);
and U1725 (N_1725,N_1408,N_1292);
nand U1726 (N_1726,N_1299,N_1245);
and U1727 (N_1727,N_1011,N_1443);
nor U1728 (N_1728,N_1350,N_1287);
xor U1729 (N_1729,N_1009,N_1153);
and U1730 (N_1730,N_1075,N_1386);
nor U1731 (N_1731,N_1385,N_1159);
xor U1732 (N_1732,N_1472,N_1013);
and U1733 (N_1733,N_1044,N_1424);
and U1734 (N_1734,N_1344,N_1383);
nand U1735 (N_1735,N_1494,N_1151);
xor U1736 (N_1736,N_1033,N_1431);
nor U1737 (N_1737,N_1398,N_1363);
nand U1738 (N_1738,N_1237,N_1312);
nand U1739 (N_1739,N_1337,N_1225);
nor U1740 (N_1740,N_1053,N_1021);
nor U1741 (N_1741,N_1480,N_1164);
or U1742 (N_1742,N_1076,N_1023);
and U1743 (N_1743,N_1249,N_1222);
xnor U1744 (N_1744,N_1345,N_1243);
nor U1745 (N_1745,N_1298,N_1489);
xnor U1746 (N_1746,N_1083,N_1357);
nor U1747 (N_1747,N_1435,N_1182);
and U1748 (N_1748,N_1174,N_1154);
nor U1749 (N_1749,N_1240,N_1138);
xnor U1750 (N_1750,N_1169,N_1310);
nand U1751 (N_1751,N_1183,N_1039);
nor U1752 (N_1752,N_1059,N_1317);
and U1753 (N_1753,N_1089,N_1378);
and U1754 (N_1754,N_1409,N_1451);
and U1755 (N_1755,N_1470,N_1235);
xor U1756 (N_1756,N_1089,N_1000);
and U1757 (N_1757,N_1276,N_1247);
nand U1758 (N_1758,N_1230,N_1020);
or U1759 (N_1759,N_1393,N_1143);
and U1760 (N_1760,N_1409,N_1287);
nor U1761 (N_1761,N_1491,N_1489);
or U1762 (N_1762,N_1459,N_1212);
nand U1763 (N_1763,N_1224,N_1216);
xnor U1764 (N_1764,N_1279,N_1185);
nand U1765 (N_1765,N_1059,N_1014);
nand U1766 (N_1766,N_1184,N_1089);
or U1767 (N_1767,N_1391,N_1095);
xor U1768 (N_1768,N_1008,N_1053);
xnor U1769 (N_1769,N_1203,N_1023);
or U1770 (N_1770,N_1409,N_1152);
or U1771 (N_1771,N_1217,N_1166);
nor U1772 (N_1772,N_1050,N_1431);
nand U1773 (N_1773,N_1059,N_1282);
and U1774 (N_1774,N_1255,N_1076);
nand U1775 (N_1775,N_1026,N_1018);
and U1776 (N_1776,N_1213,N_1017);
nor U1777 (N_1777,N_1121,N_1459);
or U1778 (N_1778,N_1162,N_1125);
xnor U1779 (N_1779,N_1402,N_1208);
xor U1780 (N_1780,N_1418,N_1212);
nand U1781 (N_1781,N_1295,N_1127);
nand U1782 (N_1782,N_1485,N_1069);
and U1783 (N_1783,N_1082,N_1149);
and U1784 (N_1784,N_1374,N_1264);
and U1785 (N_1785,N_1318,N_1452);
nand U1786 (N_1786,N_1183,N_1318);
or U1787 (N_1787,N_1414,N_1208);
nand U1788 (N_1788,N_1383,N_1234);
nand U1789 (N_1789,N_1317,N_1222);
nor U1790 (N_1790,N_1372,N_1348);
and U1791 (N_1791,N_1456,N_1266);
nand U1792 (N_1792,N_1105,N_1393);
and U1793 (N_1793,N_1378,N_1299);
or U1794 (N_1794,N_1005,N_1124);
nand U1795 (N_1795,N_1136,N_1327);
nand U1796 (N_1796,N_1149,N_1414);
and U1797 (N_1797,N_1174,N_1044);
nor U1798 (N_1798,N_1073,N_1184);
and U1799 (N_1799,N_1499,N_1041);
nor U1800 (N_1800,N_1470,N_1107);
nand U1801 (N_1801,N_1134,N_1054);
xnor U1802 (N_1802,N_1305,N_1141);
and U1803 (N_1803,N_1166,N_1250);
nor U1804 (N_1804,N_1016,N_1104);
or U1805 (N_1805,N_1039,N_1096);
and U1806 (N_1806,N_1152,N_1321);
or U1807 (N_1807,N_1197,N_1120);
xnor U1808 (N_1808,N_1143,N_1408);
and U1809 (N_1809,N_1358,N_1113);
nor U1810 (N_1810,N_1464,N_1020);
and U1811 (N_1811,N_1353,N_1235);
nor U1812 (N_1812,N_1490,N_1245);
or U1813 (N_1813,N_1078,N_1278);
nor U1814 (N_1814,N_1443,N_1452);
and U1815 (N_1815,N_1253,N_1172);
and U1816 (N_1816,N_1182,N_1028);
xor U1817 (N_1817,N_1056,N_1143);
or U1818 (N_1818,N_1496,N_1093);
nand U1819 (N_1819,N_1348,N_1292);
and U1820 (N_1820,N_1012,N_1135);
or U1821 (N_1821,N_1358,N_1311);
and U1822 (N_1822,N_1026,N_1369);
xnor U1823 (N_1823,N_1243,N_1492);
or U1824 (N_1824,N_1329,N_1419);
xor U1825 (N_1825,N_1435,N_1457);
or U1826 (N_1826,N_1490,N_1275);
and U1827 (N_1827,N_1325,N_1131);
and U1828 (N_1828,N_1297,N_1410);
nand U1829 (N_1829,N_1424,N_1215);
nor U1830 (N_1830,N_1446,N_1232);
nor U1831 (N_1831,N_1294,N_1031);
or U1832 (N_1832,N_1122,N_1063);
nand U1833 (N_1833,N_1166,N_1433);
nand U1834 (N_1834,N_1277,N_1461);
nor U1835 (N_1835,N_1188,N_1015);
nor U1836 (N_1836,N_1159,N_1183);
or U1837 (N_1837,N_1240,N_1379);
xnor U1838 (N_1838,N_1034,N_1496);
xor U1839 (N_1839,N_1119,N_1209);
nor U1840 (N_1840,N_1059,N_1411);
and U1841 (N_1841,N_1165,N_1402);
nand U1842 (N_1842,N_1372,N_1019);
and U1843 (N_1843,N_1057,N_1420);
or U1844 (N_1844,N_1186,N_1373);
and U1845 (N_1845,N_1007,N_1037);
and U1846 (N_1846,N_1391,N_1415);
xnor U1847 (N_1847,N_1006,N_1043);
xor U1848 (N_1848,N_1263,N_1137);
nand U1849 (N_1849,N_1218,N_1098);
xor U1850 (N_1850,N_1084,N_1252);
nand U1851 (N_1851,N_1478,N_1092);
xnor U1852 (N_1852,N_1499,N_1296);
nand U1853 (N_1853,N_1269,N_1472);
xor U1854 (N_1854,N_1020,N_1313);
nand U1855 (N_1855,N_1255,N_1003);
and U1856 (N_1856,N_1253,N_1191);
nor U1857 (N_1857,N_1381,N_1353);
or U1858 (N_1858,N_1257,N_1317);
xor U1859 (N_1859,N_1039,N_1117);
or U1860 (N_1860,N_1045,N_1067);
nor U1861 (N_1861,N_1249,N_1397);
or U1862 (N_1862,N_1129,N_1238);
xor U1863 (N_1863,N_1117,N_1261);
nand U1864 (N_1864,N_1486,N_1169);
xnor U1865 (N_1865,N_1260,N_1208);
nor U1866 (N_1866,N_1432,N_1401);
xor U1867 (N_1867,N_1133,N_1452);
nand U1868 (N_1868,N_1291,N_1494);
or U1869 (N_1869,N_1317,N_1205);
or U1870 (N_1870,N_1292,N_1447);
and U1871 (N_1871,N_1110,N_1267);
xnor U1872 (N_1872,N_1061,N_1395);
or U1873 (N_1873,N_1038,N_1112);
or U1874 (N_1874,N_1079,N_1235);
and U1875 (N_1875,N_1287,N_1232);
nand U1876 (N_1876,N_1420,N_1040);
xnor U1877 (N_1877,N_1061,N_1353);
nand U1878 (N_1878,N_1164,N_1388);
nor U1879 (N_1879,N_1277,N_1256);
or U1880 (N_1880,N_1497,N_1082);
or U1881 (N_1881,N_1366,N_1247);
or U1882 (N_1882,N_1010,N_1004);
xnor U1883 (N_1883,N_1073,N_1441);
xnor U1884 (N_1884,N_1203,N_1413);
and U1885 (N_1885,N_1412,N_1375);
or U1886 (N_1886,N_1366,N_1356);
and U1887 (N_1887,N_1196,N_1130);
or U1888 (N_1888,N_1043,N_1497);
nand U1889 (N_1889,N_1080,N_1164);
xnor U1890 (N_1890,N_1154,N_1336);
nand U1891 (N_1891,N_1075,N_1230);
xnor U1892 (N_1892,N_1384,N_1403);
xnor U1893 (N_1893,N_1391,N_1371);
xor U1894 (N_1894,N_1241,N_1273);
nor U1895 (N_1895,N_1124,N_1131);
and U1896 (N_1896,N_1417,N_1005);
nand U1897 (N_1897,N_1320,N_1170);
or U1898 (N_1898,N_1098,N_1082);
or U1899 (N_1899,N_1038,N_1178);
xor U1900 (N_1900,N_1360,N_1247);
xor U1901 (N_1901,N_1138,N_1394);
or U1902 (N_1902,N_1381,N_1296);
nor U1903 (N_1903,N_1390,N_1173);
or U1904 (N_1904,N_1438,N_1108);
or U1905 (N_1905,N_1347,N_1101);
or U1906 (N_1906,N_1029,N_1486);
nor U1907 (N_1907,N_1464,N_1112);
nor U1908 (N_1908,N_1151,N_1034);
nor U1909 (N_1909,N_1049,N_1334);
and U1910 (N_1910,N_1136,N_1261);
nor U1911 (N_1911,N_1476,N_1488);
nand U1912 (N_1912,N_1074,N_1397);
nand U1913 (N_1913,N_1354,N_1260);
nor U1914 (N_1914,N_1270,N_1027);
or U1915 (N_1915,N_1453,N_1337);
nand U1916 (N_1916,N_1282,N_1195);
and U1917 (N_1917,N_1014,N_1490);
xor U1918 (N_1918,N_1432,N_1319);
xor U1919 (N_1919,N_1306,N_1305);
nor U1920 (N_1920,N_1138,N_1317);
nand U1921 (N_1921,N_1419,N_1182);
nand U1922 (N_1922,N_1280,N_1078);
and U1923 (N_1923,N_1243,N_1421);
and U1924 (N_1924,N_1018,N_1368);
or U1925 (N_1925,N_1138,N_1043);
or U1926 (N_1926,N_1274,N_1219);
and U1927 (N_1927,N_1432,N_1426);
and U1928 (N_1928,N_1447,N_1281);
xnor U1929 (N_1929,N_1430,N_1468);
xor U1930 (N_1930,N_1443,N_1051);
nand U1931 (N_1931,N_1041,N_1488);
nor U1932 (N_1932,N_1050,N_1468);
nand U1933 (N_1933,N_1191,N_1068);
nand U1934 (N_1934,N_1351,N_1360);
or U1935 (N_1935,N_1337,N_1054);
nand U1936 (N_1936,N_1105,N_1480);
or U1937 (N_1937,N_1029,N_1328);
nand U1938 (N_1938,N_1289,N_1119);
xor U1939 (N_1939,N_1085,N_1425);
nor U1940 (N_1940,N_1367,N_1387);
xor U1941 (N_1941,N_1120,N_1195);
xor U1942 (N_1942,N_1237,N_1297);
xnor U1943 (N_1943,N_1241,N_1097);
nand U1944 (N_1944,N_1395,N_1113);
or U1945 (N_1945,N_1174,N_1039);
xor U1946 (N_1946,N_1014,N_1002);
and U1947 (N_1947,N_1306,N_1403);
or U1948 (N_1948,N_1128,N_1054);
and U1949 (N_1949,N_1459,N_1363);
or U1950 (N_1950,N_1082,N_1031);
nor U1951 (N_1951,N_1082,N_1105);
nand U1952 (N_1952,N_1476,N_1115);
and U1953 (N_1953,N_1380,N_1015);
nand U1954 (N_1954,N_1301,N_1481);
nor U1955 (N_1955,N_1391,N_1151);
nand U1956 (N_1956,N_1075,N_1037);
xor U1957 (N_1957,N_1044,N_1007);
or U1958 (N_1958,N_1220,N_1006);
nor U1959 (N_1959,N_1411,N_1295);
nor U1960 (N_1960,N_1416,N_1323);
and U1961 (N_1961,N_1088,N_1439);
nand U1962 (N_1962,N_1267,N_1235);
and U1963 (N_1963,N_1406,N_1462);
or U1964 (N_1964,N_1319,N_1472);
xor U1965 (N_1965,N_1441,N_1149);
xnor U1966 (N_1966,N_1268,N_1177);
and U1967 (N_1967,N_1262,N_1030);
nand U1968 (N_1968,N_1213,N_1493);
nand U1969 (N_1969,N_1047,N_1371);
or U1970 (N_1970,N_1397,N_1090);
nor U1971 (N_1971,N_1353,N_1219);
nand U1972 (N_1972,N_1450,N_1082);
or U1973 (N_1973,N_1385,N_1035);
nand U1974 (N_1974,N_1465,N_1104);
and U1975 (N_1975,N_1226,N_1165);
nor U1976 (N_1976,N_1341,N_1079);
and U1977 (N_1977,N_1015,N_1128);
nor U1978 (N_1978,N_1246,N_1326);
or U1979 (N_1979,N_1007,N_1372);
xnor U1980 (N_1980,N_1335,N_1485);
and U1981 (N_1981,N_1357,N_1251);
or U1982 (N_1982,N_1343,N_1128);
xor U1983 (N_1983,N_1307,N_1416);
and U1984 (N_1984,N_1018,N_1359);
and U1985 (N_1985,N_1061,N_1041);
and U1986 (N_1986,N_1079,N_1415);
xor U1987 (N_1987,N_1114,N_1044);
nor U1988 (N_1988,N_1340,N_1061);
nand U1989 (N_1989,N_1294,N_1142);
nor U1990 (N_1990,N_1415,N_1118);
or U1991 (N_1991,N_1038,N_1175);
nand U1992 (N_1992,N_1214,N_1066);
xor U1993 (N_1993,N_1245,N_1454);
nand U1994 (N_1994,N_1214,N_1176);
or U1995 (N_1995,N_1405,N_1012);
nand U1996 (N_1996,N_1074,N_1283);
nand U1997 (N_1997,N_1460,N_1201);
xnor U1998 (N_1998,N_1471,N_1061);
nand U1999 (N_1999,N_1028,N_1450);
nor U2000 (N_2000,N_1669,N_1528);
or U2001 (N_2001,N_1960,N_1809);
nor U2002 (N_2002,N_1780,N_1842);
nor U2003 (N_2003,N_1638,N_1525);
nand U2004 (N_2004,N_1844,N_1590);
or U2005 (N_2005,N_1831,N_1683);
xor U2006 (N_2006,N_1561,N_1794);
and U2007 (N_2007,N_1978,N_1962);
nand U2008 (N_2008,N_1724,N_1657);
xnor U2009 (N_2009,N_1503,N_1856);
nor U2010 (N_2010,N_1565,N_1951);
nand U2011 (N_2011,N_1887,N_1621);
nand U2012 (N_2012,N_1769,N_1548);
nand U2013 (N_2013,N_1571,N_1612);
xor U2014 (N_2014,N_1942,N_1852);
nor U2015 (N_2015,N_1554,N_1510);
nor U2016 (N_2016,N_1727,N_1505);
nand U2017 (N_2017,N_1775,N_1904);
and U2018 (N_2018,N_1720,N_1758);
nor U2019 (N_2019,N_1729,N_1757);
nand U2020 (N_2020,N_1784,N_1599);
or U2021 (N_2021,N_1982,N_1882);
or U2022 (N_2022,N_1923,N_1540);
nand U2023 (N_2023,N_1736,N_1667);
xor U2024 (N_2024,N_1989,N_1631);
nor U2025 (N_2025,N_1628,N_1739);
or U2026 (N_2026,N_1833,N_1584);
nor U2027 (N_2027,N_1568,N_1897);
and U2028 (N_2028,N_1557,N_1594);
and U2029 (N_2029,N_1973,N_1577);
nor U2030 (N_2030,N_1998,N_1542);
nand U2031 (N_2031,N_1947,N_1801);
nand U2032 (N_2032,N_1603,N_1911);
or U2033 (N_2033,N_1795,N_1846);
xnor U2034 (N_2034,N_1688,N_1839);
nor U2035 (N_2035,N_1545,N_1710);
nand U2036 (N_2036,N_1546,N_1777);
or U2037 (N_2037,N_1910,N_1734);
and U2038 (N_2038,N_1807,N_1779);
or U2039 (N_2039,N_1949,N_1712);
nor U2040 (N_2040,N_1964,N_1664);
xor U2041 (N_2041,N_1679,N_1682);
or U2042 (N_2042,N_1551,N_1886);
or U2043 (N_2043,N_1931,N_1576);
and U2044 (N_2044,N_1908,N_1976);
and U2045 (N_2045,N_1847,N_1627);
nand U2046 (N_2046,N_1836,N_1765);
and U2047 (N_2047,N_1953,N_1637);
nor U2048 (N_2048,N_1553,N_1957);
nor U2049 (N_2049,N_1971,N_1803);
xnor U2050 (N_2050,N_1604,N_1587);
or U2051 (N_2051,N_1614,N_1578);
or U2052 (N_2052,N_1741,N_1527);
and U2053 (N_2053,N_1963,N_1977);
nor U2054 (N_2054,N_1630,N_1871);
and U2055 (N_2055,N_1992,N_1566);
nor U2056 (N_2056,N_1644,N_1737);
and U2057 (N_2057,N_1997,N_1918);
nand U2058 (N_2058,N_1832,N_1752);
nand U2059 (N_2059,N_1671,N_1952);
and U2060 (N_2060,N_1533,N_1941);
or U2061 (N_2061,N_1880,N_1735);
nor U2062 (N_2062,N_1896,N_1754);
or U2063 (N_2063,N_1790,N_1948);
or U2064 (N_2064,N_1733,N_1793);
xor U2065 (N_2065,N_1912,N_1648);
nand U2066 (N_2066,N_1586,N_1980);
and U2067 (N_2067,N_1656,N_1675);
nor U2068 (N_2068,N_1514,N_1519);
or U2069 (N_2069,N_1802,N_1874);
xnor U2070 (N_2070,N_1969,N_1863);
nand U2071 (N_2071,N_1626,N_1579);
nand U2072 (N_2072,N_1691,N_1804);
or U2073 (N_2073,N_1526,N_1892);
nand U2074 (N_2074,N_1649,N_1569);
or U2075 (N_2075,N_1745,N_1618);
xnor U2076 (N_2076,N_1702,N_1524);
nor U2077 (N_2077,N_1991,N_1820);
or U2078 (N_2078,N_1925,N_1532);
nor U2079 (N_2079,N_1550,N_1926);
and U2080 (N_2080,N_1985,N_1861);
or U2081 (N_2081,N_1721,N_1860);
or U2082 (N_2082,N_1749,N_1591);
nor U2083 (N_2083,N_1708,N_1890);
nor U2084 (N_2084,N_1995,N_1642);
and U2085 (N_2085,N_1523,N_1956);
nor U2086 (N_2086,N_1835,N_1929);
or U2087 (N_2087,N_1913,N_1994);
xnor U2088 (N_2088,N_1654,N_1789);
nor U2089 (N_2089,N_1544,N_1785);
nand U2090 (N_2090,N_1845,N_1814);
or U2091 (N_2091,N_1870,N_1560);
nor U2092 (N_2092,N_1866,N_1703);
and U2093 (N_2093,N_1643,N_1965);
nor U2094 (N_2094,N_1744,N_1879);
xor U2095 (N_2095,N_1776,N_1601);
or U2096 (N_2096,N_1853,N_1888);
or U2097 (N_2097,N_1828,N_1782);
nor U2098 (N_2098,N_1827,N_1954);
nor U2099 (N_2099,N_1837,N_1635);
nand U2100 (N_2100,N_1796,N_1536);
and U2101 (N_2101,N_1676,N_1958);
nand U2102 (N_2102,N_1816,N_1822);
nor U2103 (N_2103,N_1522,N_1570);
xor U2104 (N_2104,N_1812,N_1917);
nand U2105 (N_2105,N_1602,N_1786);
and U2106 (N_2106,N_1981,N_1558);
or U2107 (N_2107,N_1838,N_1694);
nor U2108 (N_2108,N_1932,N_1959);
nand U2109 (N_2109,N_1502,N_1662);
and U2110 (N_2110,N_1759,N_1541);
nand U2111 (N_2111,N_1996,N_1848);
nor U2112 (N_2112,N_1849,N_1993);
nor U2113 (N_2113,N_1567,N_1945);
and U2114 (N_2114,N_1755,N_1593);
or U2115 (N_2115,N_1915,N_1583);
or U2116 (N_2116,N_1680,N_1620);
nor U2117 (N_2117,N_1661,N_1508);
or U2118 (N_2118,N_1990,N_1747);
nor U2119 (N_2119,N_1501,N_1883);
xnor U2120 (N_2120,N_1500,N_1711);
nor U2121 (N_2121,N_1746,N_1800);
xor U2122 (N_2122,N_1823,N_1850);
and U2123 (N_2123,N_1921,N_1718);
and U2124 (N_2124,N_1608,N_1686);
or U2125 (N_2125,N_1666,N_1658);
xnor U2126 (N_2126,N_1770,N_1588);
and U2127 (N_2127,N_1819,N_1824);
nand U2128 (N_2128,N_1698,N_1613);
nor U2129 (N_2129,N_1885,N_1513);
or U2130 (N_2130,N_1791,N_1826);
or U2131 (N_2131,N_1723,N_1884);
xnor U2132 (N_2132,N_1673,N_1650);
and U2133 (N_2133,N_1970,N_1936);
and U2134 (N_2134,N_1697,N_1625);
and U2135 (N_2135,N_1868,N_1955);
and U2136 (N_2136,N_1899,N_1950);
nor U2137 (N_2137,N_1813,N_1968);
nor U2138 (N_2138,N_1629,N_1891);
nor U2139 (N_2139,N_1877,N_1670);
or U2140 (N_2140,N_1520,N_1987);
nand U2141 (N_2141,N_1855,N_1895);
or U2142 (N_2142,N_1534,N_1924);
or U2143 (N_2143,N_1592,N_1574);
nor U2144 (N_2144,N_1766,N_1873);
nor U2145 (N_2145,N_1716,N_1700);
or U2146 (N_2146,N_1699,N_1646);
and U2147 (N_2147,N_1685,N_1641);
nor U2148 (N_2148,N_1684,N_1974);
nand U2149 (N_2149,N_1660,N_1783);
nand U2150 (N_2150,N_1851,N_1655);
nand U2151 (N_2151,N_1640,N_1916);
xnor U2152 (N_2152,N_1862,N_1652);
or U2153 (N_2153,N_1872,N_1909);
nand U2154 (N_2154,N_1606,N_1805);
or U2155 (N_2155,N_1999,N_1552);
nor U2156 (N_2156,N_1830,N_1772);
nand U2157 (N_2157,N_1748,N_1537);
nor U2158 (N_2158,N_1902,N_1659);
xor U2159 (N_2159,N_1573,N_1943);
nor U2160 (N_2160,N_1529,N_1778);
nor U2161 (N_2161,N_1653,N_1818);
nor U2162 (N_2162,N_1869,N_1647);
or U2163 (N_2163,N_1768,N_1753);
xnor U2164 (N_2164,N_1798,N_1972);
nor U2165 (N_2165,N_1773,N_1905);
xor U2166 (N_2166,N_1539,N_1701);
nand U2167 (N_2167,N_1616,N_1933);
xnor U2168 (N_2168,N_1967,N_1674);
xnor U2169 (N_2169,N_1840,N_1750);
xor U2170 (N_2170,N_1854,N_1731);
xnor U2171 (N_2171,N_1562,N_1507);
and U2172 (N_2172,N_1817,N_1645);
xnor U2173 (N_2173,N_1572,N_1815);
nor U2174 (N_2174,N_1531,N_1864);
nor U2175 (N_2175,N_1582,N_1668);
or U2176 (N_2176,N_1857,N_1761);
xnor U2177 (N_2177,N_1610,N_1564);
or U2178 (N_2178,N_1920,N_1781);
or U2179 (N_2179,N_1611,N_1651);
or U2180 (N_2180,N_1764,N_1984);
and U2181 (N_2181,N_1549,N_1693);
xnor U2182 (N_2182,N_1615,N_1760);
nor U2183 (N_2183,N_1979,N_1961);
nand U2184 (N_2184,N_1907,N_1829);
and U2185 (N_2185,N_1939,N_1900);
or U2186 (N_2186,N_1728,N_1726);
nand U2187 (N_2187,N_1555,N_1563);
and U2188 (N_2188,N_1713,N_1988);
nor U2189 (N_2189,N_1681,N_1517);
nor U2190 (N_2190,N_1751,N_1535);
nand U2191 (N_2191,N_1799,N_1547);
nand U2192 (N_2192,N_1623,N_1821);
nor U2193 (N_2193,N_1806,N_1763);
nor U2194 (N_2194,N_1986,N_1639);
nor U2195 (N_2195,N_1690,N_1927);
nand U2196 (N_2196,N_1930,N_1707);
nor U2197 (N_2197,N_1944,N_1919);
and U2198 (N_2198,N_1717,N_1934);
and U2199 (N_2199,N_1538,N_1940);
xnor U2200 (N_2200,N_1678,N_1622);
nand U2201 (N_2201,N_1865,N_1903);
or U2202 (N_2202,N_1633,N_1714);
xnor U2203 (N_2203,N_1893,N_1894);
and U2204 (N_2204,N_1867,N_1946);
xnor U2205 (N_2205,N_1787,N_1889);
and U2206 (N_2206,N_1983,N_1730);
nor U2207 (N_2207,N_1875,N_1521);
nor U2208 (N_2208,N_1738,N_1935);
and U2209 (N_2209,N_1859,N_1843);
and U2210 (N_2210,N_1743,N_1922);
and U2211 (N_2211,N_1704,N_1504);
and U2212 (N_2212,N_1695,N_1619);
nor U2213 (N_2213,N_1632,N_1636);
nor U2214 (N_2214,N_1692,N_1609);
and U2215 (N_2215,N_1715,N_1901);
nor U2216 (N_2216,N_1788,N_1677);
nand U2217 (N_2217,N_1575,N_1530);
nor U2218 (N_2218,N_1585,N_1825);
nand U2219 (N_2219,N_1595,N_1810);
nor U2220 (N_2220,N_1580,N_1878);
and U2221 (N_2221,N_1811,N_1774);
and U2222 (N_2222,N_1512,N_1515);
nor U2223 (N_2223,N_1858,N_1881);
and U2224 (N_2224,N_1597,N_1841);
xor U2225 (N_2225,N_1732,N_1687);
and U2226 (N_2226,N_1672,N_1756);
nor U2227 (N_2227,N_1975,N_1581);
xor U2228 (N_2228,N_1966,N_1876);
nand U2229 (N_2229,N_1665,N_1634);
or U2230 (N_2230,N_1598,N_1938);
xnor U2231 (N_2231,N_1589,N_1722);
nor U2232 (N_2232,N_1559,N_1705);
xnor U2233 (N_2233,N_1725,N_1617);
and U2234 (N_2234,N_1797,N_1719);
nor U2235 (N_2235,N_1511,N_1663);
nor U2236 (N_2236,N_1509,N_1543);
or U2237 (N_2237,N_1808,N_1762);
nor U2238 (N_2238,N_1928,N_1689);
nor U2239 (N_2239,N_1767,N_1600);
and U2240 (N_2240,N_1709,N_1834);
or U2241 (N_2241,N_1914,N_1624);
nand U2242 (N_2242,N_1696,N_1596);
or U2243 (N_2243,N_1740,N_1937);
or U2244 (N_2244,N_1516,N_1898);
and U2245 (N_2245,N_1771,N_1556);
nand U2246 (N_2246,N_1906,N_1607);
and U2247 (N_2247,N_1518,N_1506);
nor U2248 (N_2248,N_1792,N_1605);
xor U2249 (N_2249,N_1742,N_1706);
xnor U2250 (N_2250,N_1898,N_1667);
xor U2251 (N_2251,N_1676,N_1518);
or U2252 (N_2252,N_1912,N_1517);
nand U2253 (N_2253,N_1646,N_1586);
nand U2254 (N_2254,N_1581,N_1654);
nor U2255 (N_2255,N_1978,N_1543);
nor U2256 (N_2256,N_1872,N_1810);
and U2257 (N_2257,N_1678,N_1581);
or U2258 (N_2258,N_1556,N_1731);
or U2259 (N_2259,N_1513,N_1742);
or U2260 (N_2260,N_1783,N_1937);
nand U2261 (N_2261,N_1704,N_1790);
and U2262 (N_2262,N_1997,N_1815);
nor U2263 (N_2263,N_1728,N_1681);
and U2264 (N_2264,N_1646,N_1950);
nor U2265 (N_2265,N_1967,N_1758);
nand U2266 (N_2266,N_1789,N_1932);
nor U2267 (N_2267,N_1960,N_1946);
or U2268 (N_2268,N_1670,N_1561);
or U2269 (N_2269,N_1776,N_1698);
nor U2270 (N_2270,N_1596,N_1961);
nor U2271 (N_2271,N_1768,N_1793);
nand U2272 (N_2272,N_1871,N_1558);
and U2273 (N_2273,N_1855,N_1634);
xor U2274 (N_2274,N_1984,N_1677);
nor U2275 (N_2275,N_1995,N_1586);
or U2276 (N_2276,N_1678,N_1727);
or U2277 (N_2277,N_1854,N_1729);
nor U2278 (N_2278,N_1608,N_1915);
nand U2279 (N_2279,N_1893,N_1917);
xnor U2280 (N_2280,N_1740,N_1700);
nor U2281 (N_2281,N_1986,N_1825);
and U2282 (N_2282,N_1824,N_1899);
nand U2283 (N_2283,N_1526,N_1615);
xor U2284 (N_2284,N_1808,N_1761);
nand U2285 (N_2285,N_1803,N_1543);
nand U2286 (N_2286,N_1567,N_1766);
and U2287 (N_2287,N_1667,N_1663);
and U2288 (N_2288,N_1691,N_1561);
nand U2289 (N_2289,N_1634,N_1563);
and U2290 (N_2290,N_1706,N_1958);
and U2291 (N_2291,N_1606,N_1813);
nand U2292 (N_2292,N_1868,N_1893);
nor U2293 (N_2293,N_1741,N_1827);
nor U2294 (N_2294,N_1634,N_1939);
nor U2295 (N_2295,N_1975,N_1843);
and U2296 (N_2296,N_1668,N_1789);
or U2297 (N_2297,N_1869,N_1624);
nand U2298 (N_2298,N_1891,N_1876);
nand U2299 (N_2299,N_1971,N_1634);
nor U2300 (N_2300,N_1783,N_1650);
or U2301 (N_2301,N_1922,N_1605);
nand U2302 (N_2302,N_1606,N_1510);
xor U2303 (N_2303,N_1756,N_1909);
and U2304 (N_2304,N_1589,N_1533);
nand U2305 (N_2305,N_1715,N_1869);
or U2306 (N_2306,N_1637,N_1869);
nor U2307 (N_2307,N_1658,N_1678);
or U2308 (N_2308,N_1601,N_1660);
nor U2309 (N_2309,N_1715,N_1634);
and U2310 (N_2310,N_1822,N_1549);
xnor U2311 (N_2311,N_1901,N_1962);
or U2312 (N_2312,N_1530,N_1774);
and U2313 (N_2313,N_1619,N_1572);
or U2314 (N_2314,N_1518,N_1708);
xnor U2315 (N_2315,N_1748,N_1791);
nand U2316 (N_2316,N_1959,N_1620);
xor U2317 (N_2317,N_1944,N_1850);
nor U2318 (N_2318,N_1902,N_1965);
nand U2319 (N_2319,N_1923,N_1678);
or U2320 (N_2320,N_1531,N_1907);
nand U2321 (N_2321,N_1666,N_1618);
nor U2322 (N_2322,N_1941,N_1951);
and U2323 (N_2323,N_1644,N_1506);
and U2324 (N_2324,N_1678,N_1620);
nand U2325 (N_2325,N_1812,N_1612);
nand U2326 (N_2326,N_1795,N_1959);
and U2327 (N_2327,N_1522,N_1891);
nand U2328 (N_2328,N_1557,N_1589);
xnor U2329 (N_2329,N_1914,N_1647);
and U2330 (N_2330,N_1794,N_1933);
xor U2331 (N_2331,N_1669,N_1890);
and U2332 (N_2332,N_1774,N_1541);
xnor U2333 (N_2333,N_1769,N_1759);
or U2334 (N_2334,N_1758,N_1666);
or U2335 (N_2335,N_1845,N_1787);
and U2336 (N_2336,N_1937,N_1766);
nand U2337 (N_2337,N_1833,N_1555);
nor U2338 (N_2338,N_1804,N_1712);
and U2339 (N_2339,N_1757,N_1788);
nor U2340 (N_2340,N_1607,N_1777);
and U2341 (N_2341,N_1947,N_1977);
nand U2342 (N_2342,N_1797,N_1861);
nor U2343 (N_2343,N_1941,N_1922);
or U2344 (N_2344,N_1867,N_1700);
nor U2345 (N_2345,N_1527,N_1689);
nor U2346 (N_2346,N_1854,N_1594);
and U2347 (N_2347,N_1529,N_1772);
and U2348 (N_2348,N_1949,N_1961);
nor U2349 (N_2349,N_1886,N_1578);
nand U2350 (N_2350,N_1646,N_1848);
nor U2351 (N_2351,N_1990,N_1977);
or U2352 (N_2352,N_1947,N_1748);
and U2353 (N_2353,N_1606,N_1847);
xnor U2354 (N_2354,N_1642,N_1667);
xor U2355 (N_2355,N_1919,N_1509);
xor U2356 (N_2356,N_1899,N_1889);
nand U2357 (N_2357,N_1759,N_1680);
or U2358 (N_2358,N_1860,N_1958);
or U2359 (N_2359,N_1750,N_1877);
xnor U2360 (N_2360,N_1531,N_1751);
nand U2361 (N_2361,N_1547,N_1540);
and U2362 (N_2362,N_1646,N_1605);
xor U2363 (N_2363,N_1685,N_1986);
or U2364 (N_2364,N_1877,N_1679);
or U2365 (N_2365,N_1837,N_1654);
xor U2366 (N_2366,N_1615,N_1939);
and U2367 (N_2367,N_1812,N_1799);
nor U2368 (N_2368,N_1532,N_1628);
nor U2369 (N_2369,N_1706,N_1736);
xor U2370 (N_2370,N_1526,N_1753);
xnor U2371 (N_2371,N_1953,N_1970);
or U2372 (N_2372,N_1702,N_1632);
nor U2373 (N_2373,N_1514,N_1839);
nand U2374 (N_2374,N_1920,N_1760);
nor U2375 (N_2375,N_1646,N_1622);
nand U2376 (N_2376,N_1674,N_1847);
xor U2377 (N_2377,N_1519,N_1847);
xor U2378 (N_2378,N_1620,N_1658);
xnor U2379 (N_2379,N_1523,N_1976);
nand U2380 (N_2380,N_1551,N_1833);
xor U2381 (N_2381,N_1845,N_1943);
and U2382 (N_2382,N_1644,N_1503);
or U2383 (N_2383,N_1807,N_1825);
or U2384 (N_2384,N_1666,N_1961);
xnor U2385 (N_2385,N_1780,N_1902);
nand U2386 (N_2386,N_1805,N_1721);
nor U2387 (N_2387,N_1845,N_1660);
nor U2388 (N_2388,N_1973,N_1910);
or U2389 (N_2389,N_1648,N_1768);
nand U2390 (N_2390,N_1959,N_1772);
nand U2391 (N_2391,N_1961,N_1627);
or U2392 (N_2392,N_1517,N_1822);
nand U2393 (N_2393,N_1627,N_1645);
nand U2394 (N_2394,N_1617,N_1536);
nand U2395 (N_2395,N_1852,N_1801);
and U2396 (N_2396,N_1700,N_1732);
and U2397 (N_2397,N_1820,N_1838);
and U2398 (N_2398,N_1920,N_1834);
nor U2399 (N_2399,N_1802,N_1834);
nand U2400 (N_2400,N_1803,N_1999);
nor U2401 (N_2401,N_1571,N_1548);
xor U2402 (N_2402,N_1859,N_1876);
or U2403 (N_2403,N_1954,N_1712);
xor U2404 (N_2404,N_1765,N_1744);
nand U2405 (N_2405,N_1862,N_1780);
xor U2406 (N_2406,N_1540,N_1502);
and U2407 (N_2407,N_1724,N_1928);
nor U2408 (N_2408,N_1820,N_1640);
or U2409 (N_2409,N_1993,N_1919);
nor U2410 (N_2410,N_1642,N_1860);
nand U2411 (N_2411,N_1714,N_1516);
xor U2412 (N_2412,N_1942,N_1825);
nor U2413 (N_2413,N_1554,N_1947);
xnor U2414 (N_2414,N_1931,N_1662);
xor U2415 (N_2415,N_1525,N_1864);
or U2416 (N_2416,N_1547,N_1664);
nor U2417 (N_2417,N_1508,N_1664);
xnor U2418 (N_2418,N_1514,N_1772);
nand U2419 (N_2419,N_1656,N_1888);
nand U2420 (N_2420,N_1550,N_1519);
nand U2421 (N_2421,N_1797,N_1760);
xor U2422 (N_2422,N_1758,N_1849);
nor U2423 (N_2423,N_1786,N_1697);
nor U2424 (N_2424,N_1741,N_1684);
nand U2425 (N_2425,N_1560,N_1735);
nand U2426 (N_2426,N_1842,N_1527);
xnor U2427 (N_2427,N_1664,N_1818);
nand U2428 (N_2428,N_1922,N_1647);
and U2429 (N_2429,N_1851,N_1944);
nand U2430 (N_2430,N_1876,N_1825);
and U2431 (N_2431,N_1946,N_1631);
or U2432 (N_2432,N_1608,N_1647);
or U2433 (N_2433,N_1651,N_1978);
xor U2434 (N_2434,N_1522,N_1677);
and U2435 (N_2435,N_1970,N_1778);
and U2436 (N_2436,N_1776,N_1841);
nand U2437 (N_2437,N_1899,N_1582);
or U2438 (N_2438,N_1743,N_1672);
xor U2439 (N_2439,N_1780,N_1603);
and U2440 (N_2440,N_1957,N_1686);
nor U2441 (N_2441,N_1674,N_1592);
xnor U2442 (N_2442,N_1883,N_1570);
nor U2443 (N_2443,N_1832,N_1846);
nor U2444 (N_2444,N_1564,N_1848);
nor U2445 (N_2445,N_1761,N_1605);
nand U2446 (N_2446,N_1657,N_1619);
nor U2447 (N_2447,N_1800,N_1580);
and U2448 (N_2448,N_1855,N_1571);
or U2449 (N_2449,N_1873,N_1965);
or U2450 (N_2450,N_1901,N_1791);
xor U2451 (N_2451,N_1831,N_1643);
nand U2452 (N_2452,N_1940,N_1743);
nand U2453 (N_2453,N_1710,N_1612);
nand U2454 (N_2454,N_1735,N_1870);
or U2455 (N_2455,N_1731,N_1691);
or U2456 (N_2456,N_1947,N_1865);
xnor U2457 (N_2457,N_1733,N_1549);
and U2458 (N_2458,N_1603,N_1781);
and U2459 (N_2459,N_1686,N_1617);
nor U2460 (N_2460,N_1858,N_1743);
or U2461 (N_2461,N_1824,N_1825);
and U2462 (N_2462,N_1846,N_1807);
or U2463 (N_2463,N_1526,N_1650);
xor U2464 (N_2464,N_1738,N_1702);
nand U2465 (N_2465,N_1660,N_1922);
or U2466 (N_2466,N_1576,N_1686);
xor U2467 (N_2467,N_1762,N_1816);
xor U2468 (N_2468,N_1566,N_1597);
and U2469 (N_2469,N_1757,N_1824);
xor U2470 (N_2470,N_1945,N_1851);
xnor U2471 (N_2471,N_1567,N_1949);
or U2472 (N_2472,N_1920,N_1977);
xnor U2473 (N_2473,N_1519,N_1735);
and U2474 (N_2474,N_1975,N_1700);
xnor U2475 (N_2475,N_1531,N_1766);
nand U2476 (N_2476,N_1980,N_1603);
nor U2477 (N_2477,N_1918,N_1552);
nor U2478 (N_2478,N_1774,N_1965);
nand U2479 (N_2479,N_1910,N_1845);
and U2480 (N_2480,N_1691,N_1919);
xor U2481 (N_2481,N_1848,N_1648);
xnor U2482 (N_2482,N_1820,N_1586);
nor U2483 (N_2483,N_1526,N_1754);
nor U2484 (N_2484,N_1948,N_1713);
xor U2485 (N_2485,N_1794,N_1856);
nand U2486 (N_2486,N_1868,N_1751);
and U2487 (N_2487,N_1642,N_1976);
and U2488 (N_2488,N_1968,N_1741);
or U2489 (N_2489,N_1597,N_1813);
nand U2490 (N_2490,N_1627,N_1984);
and U2491 (N_2491,N_1534,N_1643);
nor U2492 (N_2492,N_1889,N_1581);
nand U2493 (N_2493,N_1961,N_1943);
xnor U2494 (N_2494,N_1777,N_1681);
or U2495 (N_2495,N_1625,N_1722);
nand U2496 (N_2496,N_1679,N_1644);
xor U2497 (N_2497,N_1908,N_1955);
nand U2498 (N_2498,N_1839,N_1835);
or U2499 (N_2499,N_1527,N_1912);
nand U2500 (N_2500,N_2296,N_2076);
xor U2501 (N_2501,N_2475,N_2041);
nor U2502 (N_2502,N_2034,N_2426);
and U2503 (N_2503,N_2406,N_2050);
nor U2504 (N_2504,N_2291,N_2047);
xor U2505 (N_2505,N_2381,N_2446);
nor U2506 (N_2506,N_2282,N_2256);
nand U2507 (N_2507,N_2244,N_2187);
and U2508 (N_2508,N_2167,N_2009);
or U2509 (N_2509,N_2103,N_2011);
xnor U2510 (N_2510,N_2361,N_2098);
and U2511 (N_2511,N_2124,N_2350);
xnor U2512 (N_2512,N_2452,N_2146);
nor U2513 (N_2513,N_2029,N_2169);
and U2514 (N_2514,N_2353,N_2100);
or U2515 (N_2515,N_2219,N_2437);
or U2516 (N_2516,N_2086,N_2273);
nand U2517 (N_2517,N_2195,N_2334);
and U2518 (N_2518,N_2237,N_2028);
nand U2519 (N_2519,N_2039,N_2003);
nor U2520 (N_2520,N_2374,N_2197);
nor U2521 (N_2521,N_2366,N_2078);
nor U2522 (N_2522,N_2059,N_2021);
xnor U2523 (N_2523,N_2307,N_2210);
nand U2524 (N_2524,N_2340,N_2153);
or U2525 (N_2525,N_2127,N_2403);
or U2526 (N_2526,N_2317,N_2405);
and U2527 (N_2527,N_2238,N_2480);
nand U2528 (N_2528,N_2170,N_2328);
and U2529 (N_2529,N_2033,N_2457);
xor U2530 (N_2530,N_2493,N_2278);
and U2531 (N_2531,N_2407,N_2188);
nor U2532 (N_2532,N_2433,N_2275);
and U2533 (N_2533,N_2201,N_2269);
or U2534 (N_2534,N_2134,N_2347);
nor U2535 (N_2535,N_2143,N_2126);
and U2536 (N_2536,N_2470,N_2140);
and U2537 (N_2537,N_2242,N_2408);
and U2538 (N_2538,N_2234,N_2357);
xor U2539 (N_2539,N_2318,N_2268);
and U2540 (N_2540,N_2451,N_2300);
and U2541 (N_2541,N_2031,N_2254);
and U2542 (N_2542,N_2016,N_2017);
or U2543 (N_2543,N_2399,N_2498);
and U2544 (N_2544,N_2092,N_2489);
and U2545 (N_2545,N_2469,N_2090);
and U2546 (N_2546,N_2232,N_2497);
nor U2547 (N_2547,N_2243,N_2066);
nor U2548 (N_2548,N_2428,N_2325);
or U2549 (N_2549,N_2385,N_2101);
xor U2550 (N_2550,N_2227,N_2330);
nor U2551 (N_2551,N_2258,N_2326);
or U2552 (N_2552,N_2311,N_2319);
nor U2553 (N_2553,N_2486,N_2211);
or U2554 (N_2554,N_2121,N_2024);
and U2555 (N_2555,N_2209,N_2056);
and U2556 (N_2556,N_2363,N_2423);
and U2557 (N_2557,N_2384,N_2231);
xnor U2558 (N_2558,N_2371,N_2065);
and U2559 (N_2559,N_2194,N_2249);
nor U2560 (N_2560,N_2485,N_2161);
nor U2561 (N_2561,N_2069,N_2320);
or U2562 (N_2562,N_2323,N_2099);
and U2563 (N_2563,N_2123,N_2263);
xor U2564 (N_2564,N_2159,N_2013);
and U2565 (N_2565,N_2149,N_2046);
xnor U2566 (N_2566,N_2255,N_2075);
and U2567 (N_2567,N_2151,N_2344);
and U2568 (N_2568,N_2040,N_2295);
nand U2569 (N_2569,N_2142,N_2080);
nand U2570 (N_2570,N_2487,N_2432);
or U2571 (N_2571,N_2310,N_2084);
and U2572 (N_2572,N_2496,N_2491);
and U2573 (N_2573,N_2358,N_2055);
nand U2574 (N_2574,N_2157,N_2276);
or U2575 (N_2575,N_2145,N_2365);
nand U2576 (N_2576,N_2203,N_2081);
nor U2577 (N_2577,N_2181,N_2175);
and U2578 (N_2578,N_2492,N_2035);
and U2579 (N_2579,N_2332,N_2252);
xor U2580 (N_2580,N_2349,N_2120);
xnor U2581 (N_2581,N_2147,N_2217);
nand U2582 (N_2582,N_2091,N_2345);
xnor U2583 (N_2583,N_2094,N_2410);
nand U2584 (N_2584,N_2096,N_2193);
or U2585 (N_2585,N_2038,N_2304);
nand U2586 (N_2586,N_2057,N_2464);
or U2587 (N_2587,N_2422,N_2052);
and U2588 (N_2588,N_2483,N_2383);
xnor U2589 (N_2589,N_2199,N_2324);
xor U2590 (N_2590,N_2179,N_2429);
or U2591 (N_2591,N_2401,N_2162);
nand U2592 (N_2592,N_2477,N_2436);
and U2593 (N_2593,N_2479,N_2434);
nor U2594 (N_2594,N_2155,N_2198);
xnor U2595 (N_2595,N_2236,N_2061);
xnor U2596 (N_2596,N_2286,N_2200);
and U2597 (N_2597,N_2251,N_2130);
nor U2598 (N_2598,N_2459,N_2224);
nand U2599 (N_2599,N_2182,N_2221);
nor U2600 (N_2600,N_2196,N_2490);
nand U2601 (N_2601,N_2277,N_2192);
or U2602 (N_2602,N_2413,N_2495);
nand U2603 (N_2603,N_2336,N_2455);
nor U2604 (N_2604,N_2095,N_2362);
and U2605 (N_2605,N_2002,N_2112);
nor U2606 (N_2606,N_2230,N_2085);
nor U2607 (N_2607,N_2245,N_2343);
or U2608 (N_2608,N_2253,N_2453);
and U2609 (N_2609,N_2132,N_2414);
nand U2610 (N_2610,N_2247,N_2032);
or U2611 (N_2611,N_2183,N_2229);
or U2612 (N_2612,N_2356,N_2222);
and U2613 (N_2613,N_2036,N_2398);
and U2614 (N_2614,N_2207,N_2087);
or U2615 (N_2615,N_2136,N_2404);
xor U2616 (N_2616,N_2113,N_2180);
nand U2617 (N_2617,N_2394,N_2215);
or U2618 (N_2618,N_2462,N_2083);
nor U2619 (N_2619,N_2139,N_2392);
nor U2620 (N_2620,N_2082,N_2054);
xor U2621 (N_2621,N_2156,N_2114);
xnor U2622 (N_2622,N_2122,N_2335);
nand U2623 (N_2623,N_2176,N_2264);
and U2624 (N_2624,N_2220,N_2128);
and U2625 (N_2625,N_2257,N_2388);
xor U2626 (N_2626,N_2416,N_2309);
nand U2627 (N_2627,N_2178,N_2014);
or U2628 (N_2628,N_2077,N_2369);
nor U2629 (N_2629,N_2418,N_2158);
nor U2630 (N_2630,N_2360,N_2088);
nand U2631 (N_2631,N_2216,N_2206);
and U2632 (N_2632,N_2163,N_2129);
and U2633 (N_2633,N_2386,N_2352);
or U2634 (N_2634,N_2270,N_2060);
or U2635 (N_2635,N_2051,N_2089);
or U2636 (N_2636,N_2005,N_2316);
or U2637 (N_2637,N_2261,N_2281);
nand U2638 (N_2638,N_2391,N_2331);
nand U2639 (N_2639,N_2072,N_2445);
nor U2640 (N_2640,N_2355,N_2043);
or U2641 (N_2641,N_2225,N_2321);
or U2642 (N_2642,N_2292,N_2107);
nand U2643 (N_2643,N_2400,N_2359);
nand U2644 (N_2644,N_2481,N_2454);
or U2645 (N_2645,N_2138,N_2303);
or U2646 (N_2646,N_2073,N_2189);
nand U2647 (N_2647,N_2015,N_2450);
nand U2648 (N_2648,N_2456,N_2287);
nor U2649 (N_2649,N_2327,N_2063);
and U2650 (N_2650,N_2144,N_2315);
xnor U2651 (N_2651,N_2379,N_2419);
xor U2652 (N_2652,N_2338,N_2233);
xnor U2653 (N_2653,N_2111,N_2045);
xor U2654 (N_2654,N_2299,N_2191);
or U2655 (N_2655,N_2164,N_2471);
or U2656 (N_2656,N_2466,N_2186);
or U2657 (N_2657,N_2006,N_2106);
and U2658 (N_2658,N_2427,N_2213);
or U2659 (N_2659,N_2415,N_2484);
nand U2660 (N_2660,N_2150,N_2067);
xnor U2661 (N_2661,N_2322,N_2118);
or U2662 (N_2662,N_2152,N_2007);
nand U2663 (N_2663,N_2022,N_2488);
or U2664 (N_2664,N_2341,N_2262);
xnor U2665 (N_2665,N_2026,N_2294);
and U2666 (N_2666,N_2053,N_2160);
and U2667 (N_2667,N_2302,N_2439);
and U2668 (N_2668,N_2494,N_2337);
nor U2669 (N_2669,N_2267,N_2214);
xor U2670 (N_2670,N_2444,N_2174);
xnor U2671 (N_2671,N_2468,N_2062);
nor U2672 (N_2672,N_2297,N_2125);
xnor U2673 (N_2673,N_2239,N_2283);
nor U2674 (N_2674,N_2478,N_2166);
or U2675 (N_2675,N_2027,N_2438);
nor U2676 (N_2676,N_2265,N_2367);
and U2677 (N_2677,N_2271,N_2393);
nor U2678 (N_2678,N_2012,N_2463);
xnor U2679 (N_2679,N_2260,N_2376);
or U2680 (N_2680,N_2373,N_2461);
nor U2681 (N_2681,N_2228,N_2131);
xor U2682 (N_2682,N_2389,N_2308);
nor U2683 (N_2683,N_2048,N_2259);
and U2684 (N_2684,N_2020,N_2467);
and U2685 (N_2685,N_2154,N_2448);
xor U2686 (N_2686,N_2458,N_2093);
and U2687 (N_2687,N_2285,N_2226);
xor U2688 (N_2688,N_2208,N_2148);
nor U2689 (N_2689,N_2411,N_2212);
xor U2690 (N_2690,N_2447,N_2290);
and U2691 (N_2691,N_2000,N_2313);
xnor U2692 (N_2692,N_2348,N_2049);
and U2693 (N_2693,N_2417,N_2339);
and U2694 (N_2694,N_2070,N_2312);
nand U2695 (N_2695,N_2284,N_2074);
xor U2696 (N_2696,N_2443,N_2010);
nand U2697 (N_2697,N_2442,N_2037);
xor U2698 (N_2698,N_2068,N_2171);
nand U2699 (N_2699,N_2117,N_2402);
xor U2700 (N_2700,N_2204,N_2165);
nand U2701 (N_2701,N_2190,N_2058);
nand U2702 (N_2702,N_2202,N_2205);
nand U2703 (N_2703,N_2272,N_2474);
nand U2704 (N_2704,N_2246,N_2421);
or U2705 (N_2705,N_2395,N_2440);
and U2706 (N_2706,N_2235,N_2449);
or U2707 (N_2707,N_2185,N_2172);
nand U2708 (N_2708,N_2223,N_2430);
and U2709 (N_2709,N_2079,N_2241);
nand U2710 (N_2710,N_2102,N_2168);
or U2711 (N_2711,N_2301,N_2266);
nand U2712 (N_2712,N_2333,N_2105);
xnor U2713 (N_2713,N_2119,N_2372);
or U2714 (N_2714,N_2298,N_2097);
nor U2715 (N_2715,N_2116,N_2364);
and U2716 (N_2716,N_2435,N_2173);
nand U2717 (N_2717,N_2064,N_2248);
nor U2718 (N_2718,N_2397,N_2293);
and U2719 (N_2719,N_2141,N_2004);
xor U2720 (N_2720,N_2375,N_2044);
nor U2721 (N_2721,N_2431,N_2377);
xor U2722 (N_2722,N_2314,N_2218);
nor U2723 (N_2723,N_2409,N_2329);
xor U2724 (N_2724,N_2424,N_2482);
and U2725 (N_2725,N_2071,N_2378);
and U2726 (N_2726,N_2380,N_2019);
xor U2727 (N_2727,N_2135,N_2025);
nor U2728 (N_2728,N_2250,N_2274);
xor U2729 (N_2729,N_2370,N_2354);
and U2730 (N_2730,N_2342,N_2109);
nand U2731 (N_2731,N_2008,N_2023);
nor U2732 (N_2732,N_2368,N_2288);
nand U2733 (N_2733,N_2240,N_2460);
xor U2734 (N_2734,N_2018,N_2441);
and U2735 (N_2735,N_2001,N_2279);
nand U2736 (N_2736,N_2306,N_2108);
or U2737 (N_2737,N_2425,N_2476);
and U2738 (N_2738,N_2104,N_2390);
nand U2739 (N_2739,N_2465,N_2387);
or U2740 (N_2740,N_2280,N_2412);
xor U2741 (N_2741,N_2030,N_2133);
xor U2742 (N_2742,N_2042,N_2137);
nor U2743 (N_2743,N_2420,N_2382);
xor U2744 (N_2744,N_2184,N_2346);
or U2745 (N_2745,N_2473,N_2177);
and U2746 (N_2746,N_2396,N_2115);
and U2747 (N_2747,N_2351,N_2289);
xnor U2748 (N_2748,N_2305,N_2499);
nor U2749 (N_2749,N_2110,N_2472);
and U2750 (N_2750,N_2060,N_2029);
or U2751 (N_2751,N_2392,N_2494);
xnor U2752 (N_2752,N_2266,N_2204);
nand U2753 (N_2753,N_2184,N_2357);
nor U2754 (N_2754,N_2150,N_2237);
nand U2755 (N_2755,N_2290,N_2332);
nand U2756 (N_2756,N_2232,N_2385);
xor U2757 (N_2757,N_2383,N_2306);
or U2758 (N_2758,N_2312,N_2181);
nor U2759 (N_2759,N_2330,N_2176);
nand U2760 (N_2760,N_2117,N_2175);
or U2761 (N_2761,N_2480,N_2376);
xnor U2762 (N_2762,N_2204,N_2227);
and U2763 (N_2763,N_2408,N_2156);
nand U2764 (N_2764,N_2492,N_2437);
xor U2765 (N_2765,N_2288,N_2007);
nand U2766 (N_2766,N_2269,N_2077);
xnor U2767 (N_2767,N_2213,N_2402);
nor U2768 (N_2768,N_2005,N_2039);
xor U2769 (N_2769,N_2139,N_2152);
nand U2770 (N_2770,N_2158,N_2431);
xor U2771 (N_2771,N_2321,N_2499);
and U2772 (N_2772,N_2021,N_2136);
and U2773 (N_2773,N_2373,N_2004);
nand U2774 (N_2774,N_2489,N_2237);
nor U2775 (N_2775,N_2204,N_2256);
or U2776 (N_2776,N_2266,N_2379);
and U2777 (N_2777,N_2289,N_2133);
xor U2778 (N_2778,N_2395,N_2047);
nor U2779 (N_2779,N_2165,N_2481);
or U2780 (N_2780,N_2245,N_2131);
and U2781 (N_2781,N_2068,N_2437);
nor U2782 (N_2782,N_2313,N_2451);
xor U2783 (N_2783,N_2351,N_2424);
nand U2784 (N_2784,N_2335,N_2044);
or U2785 (N_2785,N_2391,N_2250);
and U2786 (N_2786,N_2166,N_2366);
nand U2787 (N_2787,N_2258,N_2237);
xnor U2788 (N_2788,N_2349,N_2153);
nor U2789 (N_2789,N_2253,N_2422);
nand U2790 (N_2790,N_2175,N_2289);
xor U2791 (N_2791,N_2301,N_2453);
or U2792 (N_2792,N_2010,N_2362);
xor U2793 (N_2793,N_2379,N_2045);
or U2794 (N_2794,N_2175,N_2108);
or U2795 (N_2795,N_2326,N_2452);
xnor U2796 (N_2796,N_2268,N_2069);
xnor U2797 (N_2797,N_2443,N_2263);
and U2798 (N_2798,N_2276,N_2392);
and U2799 (N_2799,N_2320,N_2375);
or U2800 (N_2800,N_2172,N_2408);
nor U2801 (N_2801,N_2327,N_2440);
xor U2802 (N_2802,N_2490,N_2159);
and U2803 (N_2803,N_2244,N_2125);
and U2804 (N_2804,N_2123,N_2181);
xnor U2805 (N_2805,N_2356,N_2423);
nand U2806 (N_2806,N_2285,N_2190);
xnor U2807 (N_2807,N_2427,N_2120);
and U2808 (N_2808,N_2302,N_2070);
and U2809 (N_2809,N_2188,N_2377);
nand U2810 (N_2810,N_2470,N_2120);
and U2811 (N_2811,N_2034,N_2013);
xnor U2812 (N_2812,N_2014,N_2111);
and U2813 (N_2813,N_2445,N_2082);
xnor U2814 (N_2814,N_2413,N_2335);
xnor U2815 (N_2815,N_2269,N_2023);
nand U2816 (N_2816,N_2479,N_2129);
nand U2817 (N_2817,N_2424,N_2327);
or U2818 (N_2818,N_2005,N_2469);
xnor U2819 (N_2819,N_2470,N_2465);
xnor U2820 (N_2820,N_2129,N_2486);
or U2821 (N_2821,N_2121,N_2431);
or U2822 (N_2822,N_2468,N_2084);
and U2823 (N_2823,N_2415,N_2400);
or U2824 (N_2824,N_2205,N_2374);
nand U2825 (N_2825,N_2261,N_2210);
or U2826 (N_2826,N_2129,N_2153);
xnor U2827 (N_2827,N_2169,N_2105);
or U2828 (N_2828,N_2098,N_2177);
nor U2829 (N_2829,N_2424,N_2281);
or U2830 (N_2830,N_2351,N_2412);
nor U2831 (N_2831,N_2209,N_2300);
and U2832 (N_2832,N_2100,N_2231);
nor U2833 (N_2833,N_2447,N_2235);
or U2834 (N_2834,N_2224,N_2104);
xor U2835 (N_2835,N_2242,N_2311);
xor U2836 (N_2836,N_2228,N_2050);
or U2837 (N_2837,N_2401,N_2351);
nand U2838 (N_2838,N_2017,N_2141);
nand U2839 (N_2839,N_2249,N_2040);
and U2840 (N_2840,N_2479,N_2384);
or U2841 (N_2841,N_2235,N_2406);
and U2842 (N_2842,N_2112,N_2060);
nor U2843 (N_2843,N_2159,N_2473);
or U2844 (N_2844,N_2359,N_2236);
or U2845 (N_2845,N_2025,N_2298);
nor U2846 (N_2846,N_2071,N_2314);
or U2847 (N_2847,N_2404,N_2365);
nor U2848 (N_2848,N_2190,N_2478);
nor U2849 (N_2849,N_2447,N_2417);
or U2850 (N_2850,N_2405,N_2120);
and U2851 (N_2851,N_2199,N_2486);
xor U2852 (N_2852,N_2158,N_2443);
nor U2853 (N_2853,N_2454,N_2301);
and U2854 (N_2854,N_2262,N_2418);
xnor U2855 (N_2855,N_2240,N_2318);
nor U2856 (N_2856,N_2301,N_2494);
and U2857 (N_2857,N_2223,N_2468);
nor U2858 (N_2858,N_2442,N_2398);
or U2859 (N_2859,N_2422,N_2118);
nor U2860 (N_2860,N_2116,N_2496);
nand U2861 (N_2861,N_2474,N_2231);
and U2862 (N_2862,N_2316,N_2125);
and U2863 (N_2863,N_2285,N_2442);
xor U2864 (N_2864,N_2145,N_2322);
nor U2865 (N_2865,N_2086,N_2460);
nand U2866 (N_2866,N_2243,N_2428);
nand U2867 (N_2867,N_2227,N_2293);
and U2868 (N_2868,N_2290,N_2111);
xor U2869 (N_2869,N_2016,N_2498);
nor U2870 (N_2870,N_2152,N_2195);
and U2871 (N_2871,N_2156,N_2281);
xnor U2872 (N_2872,N_2441,N_2398);
or U2873 (N_2873,N_2496,N_2290);
or U2874 (N_2874,N_2164,N_2231);
and U2875 (N_2875,N_2152,N_2078);
and U2876 (N_2876,N_2429,N_2493);
nand U2877 (N_2877,N_2201,N_2274);
nand U2878 (N_2878,N_2365,N_2136);
nor U2879 (N_2879,N_2111,N_2300);
nor U2880 (N_2880,N_2193,N_2001);
nand U2881 (N_2881,N_2016,N_2247);
nand U2882 (N_2882,N_2394,N_2259);
or U2883 (N_2883,N_2176,N_2125);
nor U2884 (N_2884,N_2137,N_2465);
nor U2885 (N_2885,N_2472,N_2473);
nand U2886 (N_2886,N_2187,N_2195);
xor U2887 (N_2887,N_2161,N_2377);
and U2888 (N_2888,N_2135,N_2250);
or U2889 (N_2889,N_2497,N_2414);
xor U2890 (N_2890,N_2446,N_2412);
nor U2891 (N_2891,N_2206,N_2148);
or U2892 (N_2892,N_2434,N_2457);
or U2893 (N_2893,N_2281,N_2134);
and U2894 (N_2894,N_2209,N_2283);
nand U2895 (N_2895,N_2417,N_2085);
nand U2896 (N_2896,N_2329,N_2100);
xnor U2897 (N_2897,N_2061,N_2436);
nor U2898 (N_2898,N_2043,N_2234);
xnor U2899 (N_2899,N_2395,N_2005);
nand U2900 (N_2900,N_2487,N_2024);
or U2901 (N_2901,N_2082,N_2223);
and U2902 (N_2902,N_2485,N_2462);
and U2903 (N_2903,N_2370,N_2362);
or U2904 (N_2904,N_2039,N_2031);
xnor U2905 (N_2905,N_2480,N_2278);
or U2906 (N_2906,N_2466,N_2442);
xnor U2907 (N_2907,N_2275,N_2107);
or U2908 (N_2908,N_2033,N_2371);
and U2909 (N_2909,N_2469,N_2198);
nor U2910 (N_2910,N_2020,N_2216);
xor U2911 (N_2911,N_2111,N_2259);
and U2912 (N_2912,N_2390,N_2389);
xor U2913 (N_2913,N_2274,N_2026);
or U2914 (N_2914,N_2139,N_2478);
nand U2915 (N_2915,N_2463,N_2485);
or U2916 (N_2916,N_2313,N_2282);
or U2917 (N_2917,N_2047,N_2437);
nor U2918 (N_2918,N_2222,N_2247);
nor U2919 (N_2919,N_2393,N_2064);
nor U2920 (N_2920,N_2034,N_2331);
nand U2921 (N_2921,N_2116,N_2190);
nand U2922 (N_2922,N_2246,N_2255);
nand U2923 (N_2923,N_2317,N_2088);
nor U2924 (N_2924,N_2174,N_2282);
nand U2925 (N_2925,N_2120,N_2089);
or U2926 (N_2926,N_2022,N_2497);
or U2927 (N_2927,N_2484,N_2457);
nand U2928 (N_2928,N_2195,N_2233);
nand U2929 (N_2929,N_2047,N_2161);
nor U2930 (N_2930,N_2272,N_2349);
nor U2931 (N_2931,N_2256,N_2018);
nor U2932 (N_2932,N_2462,N_2155);
nand U2933 (N_2933,N_2215,N_2268);
or U2934 (N_2934,N_2096,N_2198);
nand U2935 (N_2935,N_2063,N_2318);
or U2936 (N_2936,N_2198,N_2135);
or U2937 (N_2937,N_2430,N_2380);
or U2938 (N_2938,N_2448,N_2002);
xnor U2939 (N_2939,N_2322,N_2015);
or U2940 (N_2940,N_2373,N_2106);
or U2941 (N_2941,N_2293,N_2325);
nand U2942 (N_2942,N_2116,N_2431);
nand U2943 (N_2943,N_2126,N_2316);
nand U2944 (N_2944,N_2093,N_2089);
nand U2945 (N_2945,N_2412,N_2237);
xnor U2946 (N_2946,N_2255,N_2058);
nand U2947 (N_2947,N_2098,N_2002);
xnor U2948 (N_2948,N_2130,N_2193);
nand U2949 (N_2949,N_2443,N_2217);
or U2950 (N_2950,N_2041,N_2115);
nand U2951 (N_2951,N_2058,N_2276);
nor U2952 (N_2952,N_2331,N_2231);
nand U2953 (N_2953,N_2080,N_2209);
and U2954 (N_2954,N_2172,N_2177);
nor U2955 (N_2955,N_2473,N_2105);
nand U2956 (N_2956,N_2403,N_2344);
xor U2957 (N_2957,N_2462,N_2084);
nor U2958 (N_2958,N_2286,N_2222);
nor U2959 (N_2959,N_2127,N_2281);
nand U2960 (N_2960,N_2200,N_2177);
nor U2961 (N_2961,N_2382,N_2159);
xor U2962 (N_2962,N_2001,N_2457);
or U2963 (N_2963,N_2440,N_2417);
or U2964 (N_2964,N_2067,N_2178);
or U2965 (N_2965,N_2291,N_2035);
and U2966 (N_2966,N_2261,N_2219);
nor U2967 (N_2967,N_2194,N_2351);
or U2968 (N_2968,N_2022,N_2464);
nor U2969 (N_2969,N_2168,N_2476);
or U2970 (N_2970,N_2147,N_2062);
nand U2971 (N_2971,N_2359,N_2300);
and U2972 (N_2972,N_2171,N_2432);
xor U2973 (N_2973,N_2349,N_2072);
nor U2974 (N_2974,N_2482,N_2309);
and U2975 (N_2975,N_2466,N_2091);
or U2976 (N_2976,N_2130,N_2116);
xor U2977 (N_2977,N_2055,N_2328);
xnor U2978 (N_2978,N_2316,N_2413);
and U2979 (N_2979,N_2168,N_2034);
nor U2980 (N_2980,N_2199,N_2275);
and U2981 (N_2981,N_2473,N_2321);
or U2982 (N_2982,N_2097,N_2145);
nor U2983 (N_2983,N_2447,N_2037);
nand U2984 (N_2984,N_2260,N_2215);
nand U2985 (N_2985,N_2377,N_2085);
nor U2986 (N_2986,N_2116,N_2456);
xor U2987 (N_2987,N_2107,N_2081);
nand U2988 (N_2988,N_2016,N_2064);
and U2989 (N_2989,N_2025,N_2305);
xnor U2990 (N_2990,N_2331,N_2078);
xor U2991 (N_2991,N_2397,N_2319);
nor U2992 (N_2992,N_2091,N_2299);
or U2993 (N_2993,N_2486,N_2000);
nand U2994 (N_2994,N_2290,N_2425);
nand U2995 (N_2995,N_2234,N_2203);
and U2996 (N_2996,N_2139,N_2233);
or U2997 (N_2997,N_2172,N_2080);
xnor U2998 (N_2998,N_2469,N_2246);
nor U2999 (N_2999,N_2103,N_2127);
nor U3000 (N_3000,N_2858,N_2595);
and U3001 (N_3001,N_2657,N_2952);
nand U3002 (N_3002,N_2544,N_2732);
and U3003 (N_3003,N_2670,N_2503);
or U3004 (N_3004,N_2794,N_2652);
xor U3005 (N_3005,N_2564,N_2869);
xor U3006 (N_3006,N_2863,N_2534);
nor U3007 (N_3007,N_2761,N_2658);
nand U3008 (N_3008,N_2524,N_2663);
or U3009 (N_3009,N_2728,N_2558);
nand U3010 (N_3010,N_2557,N_2973);
nor U3011 (N_3011,N_2923,N_2796);
nor U3012 (N_3012,N_2783,N_2946);
or U3013 (N_3013,N_2938,N_2601);
and U3014 (N_3014,N_2698,N_2539);
nor U3015 (N_3015,N_2874,N_2617);
and U3016 (N_3016,N_2905,N_2784);
xnor U3017 (N_3017,N_2561,N_2549);
or U3018 (N_3018,N_2958,N_2779);
nand U3019 (N_3019,N_2724,N_2582);
nor U3020 (N_3020,N_2580,N_2686);
or U3021 (N_3021,N_2845,N_2701);
xnor U3022 (N_3022,N_2739,N_2959);
and U3023 (N_3023,N_2883,N_2550);
nand U3024 (N_3024,N_2909,N_2989);
and U3025 (N_3025,N_2540,N_2639);
and U3026 (N_3026,N_2713,N_2554);
or U3027 (N_3027,N_2528,N_2625);
or U3028 (N_3028,N_2849,N_2994);
or U3029 (N_3029,N_2681,N_2894);
nor U3030 (N_3030,N_2945,N_2797);
nor U3031 (N_3031,N_2548,N_2935);
nor U3032 (N_3032,N_2815,N_2543);
and U3033 (N_3033,N_2943,N_2574);
or U3034 (N_3034,N_2819,N_2934);
and U3035 (N_3035,N_2611,N_2970);
nand U3036 (N_3036,N_2804,N_2850);
and U3037 (N_3037,N_2963,N_2978);
xor U3038 (N_3038,N_2756,N_2600);
and U3039 (N_3039,N_2620,N_2987);
and U3040 (N_3040,N_2829,N_2764);
or U3041 (N_3041,N_2769,N_2593);
xnor U3042 (N_3042,N_2594,N_2809);
or U3043 (N_3043,N_2862,N_2846);
nand U3044 (N_3044,N_2626,N_2805);
and U3045 (N_3045,N_2985,N_2810);
or U3046 (N_3046,N_2974,N_2720);
or U3047 (N_3047,N_2527,N_2953);
and U3048 (N_3048,N_2800,N_2906);
and U3049 (N_3049,N_2910,N_2705);
nand U3050 (N_3050,N_2834,N_2868);
and U3051 (N_3051,N_2791,N_2598);
or U3052 (N_3052,N_2696,N_2505);
xnor U3053 (N_3053,N_2758,N_2932);
xor U3054 (N_3054,N_2745,N_2526);
nor U3055 (N_3055,N_2838,N_2707);
xor U3056 (N_3056,N_2763,N_2591);
xor U3057 (N_3057,N_2744,N_2789);
xor U3058 (N_3058,N_2826,N_2637);
xor U3059 (N_3059,N_2683,N_2878);
nand U3060 (N_3060,N_2828,N_2772);
nand U3061 (N_3061,N_2913,N_2609);
xor U3062 (N_3062,N_2502,N_2866);
or U3063 (N_3063,N_2673,N_2518);
and U3064 (N_3064,N_2753,N_2969);
nand U3065 (N_3065,N_2513,N_2983);
nor U3066 (N_3066,N_2867,N_2900);
or U3067 (N_3067,N_2781,N_2991);
nand U3068 (N_3068,N_2577,N_2651);
xnor U3069 (N_3069,N_2602,N_2802);
or U3070 (N_3070,N_2795,N_2857);
xnor U3071 (N_3071,N_2852,N_2837);
nor U3072 (N_3072,N_2871,N_2759);
or U3073 (N_3073,N_2522,N_2552);
or U3074 (N_3074,N_2592,N_2741);
nor U3075 (N_3075,N_2608,N_2603);
nand U3076 (N_3076,N_2508,N_2955);
nor U3077 (N_3077,N_2699,N_2914);
xor U3078 (N_3078,N_2532,N_2619);
or U3079 (N_3079,N_2997,N_2790);
xor U3080 (N_3080,N_2965,N_2853);
or U3081 (N_3081,N_2954,N_2859);
nor U3082 (N_3082,N_2642,N_2578);
nand U3083 (N_3083,N_2632,N_2976);
and U3084 (N_3084,N_2519,N_2830);
and U3085 (N_3085,N_2629,N_2998);
or U3086 (N_3086,N_2604,N_2563);
nor U3087 (N_3087,N_2517,N_2562);
or U3088 (N_3088,N_2730,N_2674);
and U3089 (N_3089,N_2876,N_2892);
nor U3090 (N_3090,N_2507,N_2788);
xor U3091 (N_3091,N_2525,N_2638);
or U3092 (N_3092,N_2811,N_2556);
or U3093 (N_3093,N_2931,N_2654);
xnor U3094 (N_3094,N_2856,N_2835);
nand U3095 (N_3095,N_2623,N_2827);
nor U3096 (N_3096,N_2520,N_2715);
or U3097 (N_3097,N_2687,N_2731);
xor U3098 (N_3098,N_2723,N_2662);
nand U3099 (N_3099,N_2690,N_2590);
or U3100 (N_3100,N_2706,N_2545);
nand U3101 (N_3101,N_2907,N_2551);
and U3102 (N_3102,N_2566,N_2615);
nor U3103 (N_3103,N_2773,N_2812);
nor U3104 (N_3104,N_2521,N_2915);
and U3105 (N_3105,N_2610,N_2864);
xnor U3106 (N_3106,N_2599,N_2515);
or U3107 (N_3107,N_2684,N_2668);
xor U3108 (N_3108,N_2917,N_2921);
and U3109 (N_3109,N_2988,N_2823);
or U3110 (N_3110,N_2650,N_2672);
nor U3111 (N_3111,N_2660,N_2896);
nor U3112 (N_3112,N_2992,N_2588);
nand U3113 (N_3113,N_2714,N_2933);
nand U3114 (N_3114,N_2531,N_2614);
and U3115 (N_3115,N_2891,N_2725);
and U3116 (N_3116,N_2755,N_2721);
nand U3117 (N_3117,N_2606,N_2680);
and U3118 (N_3118,N_2555,N_2716);
nor U3119 (N_3119,N_2803,N_2972);
and U3120 (N_3120,N_2565,N_2695);
and U3121 (N_3121,N_2995,N_2785);
xnor U3122 (N_3122,N_2752,N_2685);
xor U3123 (N_3123,N_2799,N_2840);
xnor U3124 (N_3124,N_2579,N_2736);
nand U3125 (N_3125,N_2999,N_2816);
nand U3126 (N_3126,N_2635,N_2583);
nand U3127 (N_3127,N_2833,N_2726);
or U3128 (N_3128,N_2589,N_2990);
nor U3129 (N_3129,N_2627,N_2986);
xnor U3130 (N_3130,N_2806,N_2612);
xnor U3131 (N_3131,N_2500,N_2908);
and U3132 (N_3132,N_2960,N_2509);
and U3133 (N_3133,N_2581,N_2722);
or U3134 (N_3134,N_2746,N_2980);
or U3135 (N_3135,N_2655,N_2882);
and U3136 (N_3136,N_2872,N_2754);
and U3137 (N_3137,N_2586,N_2832);
nand U3138 (N_3138,N_2675,N_2679);
and U3139 (N_3139,N_2760,N_2899);
or U3140 (N_3140,N_2975,N_2911);
nand U3141 (N_3141,N_2870,N_2553);
or U3142 (N_3142,N_2622,N_2504);
nand U3143 (N_3143,N_2630,N_2982);
xnor U3144 (N_3144,N_2537,N_2648);
xnor U3145 (N_3145,N_2904,N_2571);
nor U3146 (N_3146,N_2559,N_2697);
nand U3147 (N_3147,N_2814,N_2645);
xnor U3148 (N_3148,N_2860,N_2700);
nor U3149 (N_3149,N_2942,N_2718);
nand U3150 (N_3150,N_2768,N_2708);
and U3151 (N_3151,N_2692,N_2538);
nand U3152 (N_3152,N_2664,N_2666);
and U3153 (N_3153,N_2893,N_2777);
xor U3154 (N_3154,N_2901,N_2780);
and U3155 (N_3155,N_2735,N_2895);
or U3156 (N_3156,N_2573,N_2847);
and U3157 (N_3157,N_2950,N_2861);
nor U3158 (N_3158,N_2966,N_2808);
xor U3159 (N_3159,N_2688,N_2511);
and U3160 (N_3160,N_2941,N_2616);
nand U3161 (N_3161,N_2854,N_2776);
or U3162 (N_3162,N_2875,N_2584);
or U3163 (N_3163,N_2964,N_2596);
or U3164 (N_3164,N_2743,N_2855);
nor U3165 (N_3165,N_2567,N_2618);
nand U3166 (N_3166,N_2902,N_2535);
xor U3167 (N_3167,N_2865,N_2766);
or U3168 (N_3168,N_2922,N_2512);
nand U3169 (N_3169,N_2897,N_2824);
xor U3170 (N_3170,N_2719,N_2798);
nand U3171 (N_3171,N_2689,N_2587);
nand U3172 (N_3172,N_2979,N_2903);
nand U3173 (N_3173,N_2993,N_2671);
or U3174 (N_3174,N_2649,N_2977);
nand U3175 (N_3175,N_2740,N_2782);
xor U3176 (N_3176,N_2920,N_2930);
xnor U3177 (N_3177,N_2928,N_2624);
or U3178 (N_3178,N_2501,N_2842);
or U3179 (N_3179,N_2844,N_2646);
xor U3180 (N_3180,N_2961,N_2962);
xor U3181 (N_3181,N_2676,N_2702);
and U3182 (N_3182,N_2542,N_2711);
or U3183 (N_3183,N_2704,N_2925);
or U3184 (N_3184,N_2929,N_2643);
xor U3185 (N_3185,N_2807,N_2641);
and U3186 (N_3186,N_2887,N_2510);
xor U3187 (N_3187,N_2981,N_2631);
or U3188 (N_3188,N_2748,N_2569);
and U3189 (N_3189,N_2628,N_2644);
or U3190 (N_3190,N_2541,N_2778);
xnor U3191 (N_3191,N_2613,N_2793);
nor U3192 (N_3192,N_2749,N_2792);
nand U3193 (N_3193,N_2712,N_2734);
nand U3194 (N_3194,N_2822,N_2747);
xnor U3195 (N_3195,N_2572,N_2813);
nor U3196 (N_3196,N_2762,N_2971);
or U3197 (N_3197,N_2786,N_2956);
and U3198 (N_3198,N_2787,N_2656);
or U3199 (N_3199,N_2729,N_2514);
or U3200 (N_3200,N_2968,N_2831);
xor U3201 (N_3201,N_2585,N_2516);
nor U3202 (N_3202,N_2733,N_2843);
xor U3203 (N_3203,N_2839,N_2546);
xnor U3204 (N_3204,N_2817,N_2948);
nand U3205 (N_3205,N_2633,N_2751);
nand U3206 (N_3206,N_2750,N_2890);
nand U3207 (N_3207,N_2881,N_2694);
xor U3208 (N_3208,N_2944,N_2774);
nand U3209 (N_3209,N_2703,N_2880);
nand U3210 (N_3210,N_2889,N_2560);
or U3211 (N_3211,N_2506,N_2940);
nor U3212 (N_3212,N_2825,N_2742);
or U3213 (N_3213,N_2529,N_2770);
nor U3214 (N_3214,N_2738,N_2710);
xnor U3215 (N_3215,N_2661,N_2669);
nor U3216 (N_3216,N_2667,N_2873);
nand U3217 (N_3217,N_2607,N_2659);
xor U3218 (N_3218,N_2775,N_2820);
nor U3219 (N_3219,N_2927,N_2924);
or U3220 (N_3220,N_2530,N_2523);
nor U3221 (N_3221,N_2682,N_2547);
nor U3222 (N_3222,N_2533,N_2898);
and U3223 (N_3223,N_2653,N_2918);
xnor U3224 (N_3224,N_2841,N_2767);
nand U3225 (N_3225,N_2919,N_2536);
xor U3226 (N_3226,N_2634,N_2568);
and U3227 (N_3227,N_2636,N_2771);
nor U3228 (N_3228,N_2709,N_2848);
and U3229 (N_3229,N_2818,N_2916);
or U3230 (N_3230,N_2621,N_2575);
and U3231 (N_3231,N_2647,N_2691);
nor U3232 (N_3232,N_2996,N_2877);
xnor U3233 (N_3233,N_2765,N_2576);
or U3234 (N_3234,N_2886,N_2757);
nand U3235 (N_3235,N_2836,N_2821);
nand U3236 (N_3236,N_2737,N_2693);
nand U3237 (N_3237,N_2851,N_2570);
xor U3238 (N_3238,N_2949,N_2884);
and U3239 (N_3239,N_2678,N_2937);
or U3240 (N_3240,N_2677,N_2879);
or U3241 (N_3241,N_2912,N_2947);
xnor U3242 (N_3242,N_2984,N_2951);
nor U3243 (N_3243,N_2640,N_2717);
xnor U3244 (N_3244,N_2888,N_2967);
or U3245 (N_3245,N_2605,N_2801);
nor U3246 (N_3246,N_2597,N_2936);
xor U3247 (N_3247,N_2957,N_2885);
nand U3248 (N_3248,N_2727,N_2926);
xnor U3249 (N_3249,N_2939,N_2665);
and U3250 (N_3250,N_2785,N_2747);
xor U3251 (N_3251,N_2825,N_2654);
or U3252 (N_3252,N_2740,N_2801);
nor U3253 (N_3253,N_2797,N_2724);
or U3254 (N_3254,N_2559,N_2610);
nor U3255 (N_3255,N_2994,N_2741);
and U3256 (N_3256,N_2672,N_2767);
and U3257 (N_3257,N_2738,N_2671);
and U3258 (N_3258,N_2856,N_2734);
nor U3259 (N_3259,N_2614,N_2863);
xor U3260 (N_3260,N_2502,N_2518);
nand U3261 (N_3261,N_2574,N_2720);
or U3262 (N_3262,N_2662,N_2944);
xnor U3263 (N_3263,N_2647,N_2670);
or U3264 (N_3264,N_2776,N_2747);
and U3265 (N_3265,N_2881,N_2985);
nor U3266 (N_3266,N_2671,N_2533);
nor U3267 (N_3267,N_2677,N_2814);
nand U3268 (N_3268,N_2686,N_2850);
nor U3269 (N_3269,N_2916,N_2906);
xor U3270 (N_3270,N_2699,N_2705);
nor U3271 (N_3271,N_2900,N_2931);
or U3272 (N_3272,N_2591,N_2883);
nor U3273 (N_3273,N_2589,N_2925);
and U3274 (N_3274,N_2829,N_2909);
nand U3275 (N_3275,N_2786,N_2890);
and U3276 (N_3276,N_2730,N_2760);
nor U3277 (N_3277,N_2522,N_2897);
xor U3278 (N_3278,N_2576,N_2648);
xor U3279 (N_3279,N_2950,N_2700);
or U3280 (N_3280,N_2781,N_2833);
xnor U3281 (N_3281,N_2705,N_2509);
nand U3282 (N_3282,N_2632,N_2762);
or U3283 (N_3283,N_2876,N_2874);
nor U3284 (N_3284,N_2748,N_2868);
nand U3285 (N_3285,N_2528,N_2957);
nor U3286 (N_3286,N_2982,N_2520);
or U3287 (N_3287,N_2903,N_2766);
or U3288 (N_3288,N_2612,N_2835);
nand U3289 (N_3289,N_2511,N_2651);
xnor U3290 (N_3290,N_2642,N_2713);
or U3291 (N_3291,N_2818,N_2924);
or U3292 (N_3292,N_2658,N_2782);
and U3293 (N_3293,N_2528,N_2688);
nor U3294 (N_3294,N_2515,N_2505);
nand U3295 (N_3295,N_2658,N_2600);
xor U3296 (N_3296,N_2864,N_2902);
xor U3297 (N_3297,N_2603,N_2861);
nor U3298 (N_3298,N_2764,N_2912);
nand U3299 (N_3299,N_2545,N_2753);
or U3300 (N_3300,N_2622,N_2993);
and U3301 (N_3301,N_2825,N_2973);
xor U3302 (N_3302,N_2897,N_2647);
nand U3303 (N_3303,N_2507,N_2886);
and U3304 (N_3304,N_2574,N_2839);
or U3305 (N_3305,N_2914,N_2757);
xnor U3306 (N_3306,N_2530,N_2579);
and U3307 (N_3307,N_2613,N_2680);
or U3308 (N_3308,N_2780,N_2552);
nand U3309 (N_3309,N_2992,N_2653);
xnor U3310 (N_3310,N_2887,N_2973);
nor U3311 (N_3311,N_2755,N_2839);
nand U3312 (N_3312,N_2598,N_2670);
xnor U3313 (N_3313,N_2865,N_2527);
or U3314 (N_3314,N_2946,N_2703);
and U3315 (N_3315,N_2680,N_2978);
xnor U3316 (N_3316,N_2934,N_2608);
xnor U3317 (N_3317,N_2833,N_2960);
and U3318 (N_3318,N_2944,N_2875);
or U3319 (N_3319,N_2571,N_2569);
nor U3320 (N_3320,N_2534,N_2508);
or U3321 (N_3321,N_2974,N_2882);
and U3322 (N_3322,N_2533,N_2731);
xor U3323 (N_3323,N_2924,N_2583);
xor U3324 (N_3324,N_2967,N_2835);
nand U3325 (N_3325,N_2652,N_2801);
nand U3326 (N_3326,N_2783,N_2554);
nand U3327 (N_3327,N_2662,N_2584);
and U3328 (N_3328,N_2779,N_2769);
and U3329 (N_3329,N_2827,N_2655);
nor U3330 (N_3330,N_2895,N_2778);
nor U3331 (N_3331,N_2672,N_2974);
or U3332 (N_3332,N_2774,N_2849);
nand U3333 (N_3333,N_2816,N_2512);
nor U3334 (N_3334,N_2886,N_2522);
xnor U3335 (N_3335,N_2831,N_2785);
nand U3336 (N_3336,N_2971,N_2844);
xor U3337 (N_3337,N_2562,N_2809);
nand U3338 (N_3338,N_2648,N_2970);
xor U3339 (N_3339,N_2786,N_2942);
xor U3340 (N_3340,N_2891,N_2756);
or U3341 (N_3341,N_2500,N_2787);
nand U3342 (N_3342,N_2985,N_2771);
and U3343 (N_3343,N_2687,N_2652);
nor U3344 (N_3344,N_2870,N_2841);
xnor U3345 (N_3345,N_2789,N_2855);
nor U3346 (N_3346,N_2616,N_2874);
xor U3347 (N_3347,N_2881,N_2512);
nand U3348 (N_3348,N_2540,N_2753);
nand U3349 (N_3349,N_2798,N_2897);
nor U3350 (N_3350,N_2697,N_2957);
and U3351 (N_3351,N_2736,N_2734);
xor U3352 (N_3352,N_2920,N_2942);
and U3353 (N_3353,N_2865,N_2722);
nor U3354 (N_3354,N_2994,N_2545);
xnor U3355 (N_3355,N_2805,N_2775);
or U3356 (N_3356,N_2528,N_2766);
xnor U3357 (N_3357,N_2882,N_2669);
and U3358 (N_3358,N_2574,N_2679);
nand U3359 (N_3359,N_2640,N_2548);
or U3360 (N_3360,N_2599,N_2868);
xnor U3361 (N_3361,N_2808,N_2674);
or U3362 (N_3362,N_2552,N_2830);
nand U3363 (N_3363,N_2577,N_2691);
nand U3364 (N_3364,N_2748,N_2682);
or U3365 (N_3365,N_2879,N_2635);
or U3366 (N_3366,N_2870,N_2534);
or U3367 (N_3367,N_2996,N_2636);
and U3368 (N_3368,N_2815,N_2888);
or U3369 (N_3369,N_2891,N_2969);
nor U3370 (N_3370,N_2706,N_2563);
and U3371 (N_3371,N_2993,N_2966);
xor U3372 (N_3372,N_2907,N_2571);
nand U3373 (N_3373,N_2513,N_2888);
xnor U3374 (N_3374,N_2637,N_2766);
or U3375 (N_3375,N_2832,N_2548);
xnor U3376 (N_3376,N_2962,N_2955);
xor U3377 (N_3377,N_2567,N_2796);
nor U3378 (N_3378,N_2598,N_2953);
xnor U3379 (N_3379,N_2829,N_2628);
and U3380 (N_3380,N_2556,N_2717);
xnor U3381 (N_3381,N_2839,N_2572);
xor U3382 (N_3382,N_2701,N_2797);
xnor U3383 (N_3383,N_2835,N_2947);
xnor U3384 (N_3384,N_2772,N_2881);
or U3385 (N_3385,N_2780,N_2571);
and U3386 (N_3386,N_2724,N_2888);
nand U3387 (N_3387,N_2770,N_2662);
nor U3388 (N_3388,N_2626,N_2896);
and U3389 (N_3389,N_2633,N_2670);
and U3390 (N_3390,N_2568,N_2713);
nor U3391 (N_3391,N_2801,N_2756);
xor U3392 (N_3392,N_2815,N_2685);
nor U3393 (N_3393,N_2508,N_2726);
nor U3394 (N_3394,N_2579,N_2801);
nor U3395 (N_3395,N_2797,N_2843);
or U3396 (N_3396,N_2757,N_2690);
nor U3397 (N_3397,N_2717,N_2907);
or U3398 (N_3398,N_2909,N_2957);
nand U3399 (N_3399,N_2951,N_2963);
or U3400 (N_3400,N_2563,N_2655);
nand U3401 (N_3401,N_2713,N_2739);
and U3402 (N_3402,N_2678,N_2842);
xor U3403 (N_3403,N_2723,N_2793);
nand U3404 (N_3404,N_2638,N_2732);
or U3405 (N_3405,N_2771,N_2608);
or U3406 (N_3406,N_2814,N_2684);
nor U3407 (N_3407,N_2622,N_2503);
nor U3408 (N_3408,N_2967,N_2523);
xor U3409 (N_3409,N_2508,N_2504);
nor U3410 (N_3410,N_2879,N_2841);
xor U3411 (N_3411,N_2662,N_2621);
nor U3412 (N_3412,N_2575,N_2755);
nand U3413 (N_3413,N_2633,N_2553);
xnor U3414 (N_3414,N_2604,N_2935);
or U3415 (N_3415,N_2931,N_2982);
xor U3416 (N_3416,N_2793,N_2770);
xnor U3417 (N_3417,N_2717,N_2637);
nor U3418 (N_3418,N_2645,N_2822);
or U3419 (N_3419,N_2642,N_2573);
or U3420 (N_3420,N_2909,N_2982);
xor U3421 (N_3421,N_2952,N_2634);
nand U3422 (N_3422,N_2906,N_2555);
xnor U3423 (N_3423,N_2840,N_2785);
xor U3424 (N_3424,N_2931,N_2700);
or U3425 (N_3425,N_2752,N_2583);
or U3426 (N_3426,N_2842,N_2690);
and U3427 (N_3427,N_2979,N_2642);
nand U3428 (N_3428,N_2927,N_2837);
xor U3429 (N_3429,N_2841,N_2617);
and U3430 (N_3430,N_2847,N_2978);
xor U3431 (N_3431,N_2529,N_2593);
and U3432 (N_3432,N_2821,N_2783);
nor U3433 (N_3433,N_2970,N_2512);
nand U3434 (N_3434,N_2559,N_2742);
and U3435 (N_3435,N_2887,N_2910);
and U3436 (N_3436,N_2972,N_2525);
xnor U3437 (N_3437,N_2676,N_2609);
or U3438 (N_3438,N_2930,N_2997);
xnor U3439 (N_3439,N_2985,N_2792);
xor U3440 (N_3440,N_2923,N_2647);
and U3441 (N_3441,N_2896,N_2980);
xor U3442 (N_3442,N_2999,N_2518);
and U3443 (N_3443,N_2563,N_2991);
and U3444 (N_3444,N_2605,N_2623);
nand U3445 (N_3445,N_2710,N_2816);
nand U3446 (N_3446,N_2689,N_2670);
xor U3447 (N_3447,N_2943,N_2600);
nor U3448 (N_3448,N_2576,N_2633);
or U3449 (N_3449,N_2631,N_2700);
and U3450 (N_3450,N_2551,N_2564);
and U3451 (N_3451,N_2739,N_2747);
xor U3452 (N_3452,N_2767,N_2725);
nor U3453 (N_3453,N_2963,N_2718);
xor U3454 (N_3454,N_2917,N_2575);
and U3455 (N_3455,N_2545,N_2848);
nor U3456 (N_3456,N_2600,N_2696);
nand U3457 (N_3457,N_2516,N_2697);
nand U3458 (N_3458,N_2808,N_2560);
nand U3459 (N_3459,N_2799,N_2542);
nor U3460 (N_3460,N_2990,N_2602);
and U3461 (N_3461,N_2758,N_2673);
xnor U3462 (N_3462,N_2804,N_2602);
and U3463 (N_3463,N_2848,N_2523);
nand U3464 (N_3464,N_2900,N_2724);
or U3465 (N_3465,N_2988,N_2837);
xnor U3466 (N_3466,N_2586,N_2566);
nor U3467 (N_3467,N_2954,N_2880);
or U3468 (N_3468,N_2524,N_2910);
and U3469 (N_3469,N_2719,N_2629);
and U3470 (N_3470,N_2624,N_2680);
and U3471 (N_3471,N_2804,N_2741);
nand U3472 (N_3472,N_2889,N_2814);
nor U3473 (N_3473,N_2997,N_2743);
xnor U3474 (N_3474,N_2867,N_2544);
or U3475 (N_3475,N_2622,N_2756);
xnor U3476 (N_3476,N_2637,N_2640);
xor U3477 (N_3477,N_2578,N_2751);
nand U3478 (N_3478,N_2634,N_2792);
xor U3479 (N_3479,N_2503,N_2762);
and U3480 (N_3480,N_2939,N_2546);
or U3481 (N_3481,N_2689,N_2677);
xnor U3482 (N_3482,N_2764,N_2751);
nor U3483 (N_3483,N_2624,N_2970);
and U3484 (N_3484,N_2502,N_2906);
xnor U3485 (N_3485,N_2559,N_2975);
nor U3486 (N_3486,N_2753,N_2924);
xnor U3487 (N_3487,N_2681,N_2932);
nand U3488 (N_3488,N_2925,N_2763);
or U3489 (N_3489,N_2832,N_2529);
or U3490 (N_3490,N_2906,N_2874);
or U3491 (N_3491,N_2760,N_2916);
nand U3492 (N_3492,N_2532,N_2790);
or U3493 (N_3493,N_2731,N_2893);
and U3494 (N_3494,N_2776,N_2861);
xor U3495 (N_3495,N_2669,N_2530);
xnor U3496 (N_3496,N_2550,N_2596);
nor U3497 (N_3497,N_2623,N_2631);
xor U3498 (N_3498,N_2603,N_2821);
nor U3499 (N_3499,N_2601,N_2766);
and U3500 (N_3500,N_3221,N_3444);
xnor U3501 (N_3501,N_3000,N_3181);
and U3502 (N_3502,N_3051,N_3114);
nand U3503 (N_3503,N_3091,N_3278);
xnor U3504 (N_3504,N_3293,N_3412);
nand U3505 (N_3505,N_3447,N_3156);
and U3506 (N_3506,N_3301,N_3405);
or U3507 (N_3507,N_3426,N_3282);
and U3508 (N_3508,N_3111,N_3003);
and U3509 (N_3509,N_3407,N_3090);
or U3510 (N_3510,N_3033,N_3038);
and U3511 (N_3511,N_3153,N_3427);
and U3512 (N_3512,N_3258,N_3267);
and U3513 (N_3513,N_3007,N_3312);
and U3514 (N_3514,N_3232,N_3175);
nand U3515 (N_3515,N_3057,N_3096);
nand U3516 (N_3516,N_3131,N_3120);
or U3517 (N_3517,N_3343,N_3435);
and U3518 (N_3518,N_3230,N_3471);
or U3519 (N_3519,N_3254,N_3121);
and U3520 (N_3520,N_3260,N_3197);
nand U3521 (N_3521,N_3452,N_3018);
and U3522 (N_3522,N_3355,N_3286);
nor U3523 (N_3523,N_3129,N_3315);
and U3524 (N_3524,N_3160,N_3306);
or U3525 (N_3525,N_3261,N_3478);
nor U3526 (N_3526,N_3037,N_3314);
and U3527 (N_3527,N_3028,N_3448);
nor U3528 (N_3528,N_3337,N_3087);
or U3529 (N_3529,N_3014,N_3185);
and U3530 (N_3530,N_3399,N_3487);
nand U3531 (N_3531,N_3458,N_3137);
or U3532 (N_3532,N_3468,N_3474);
nor U3533 (N_3533,N_3217,N_3348);
nand U3534 (N_3534,N_3250,N_3335);
and U3535 (N_3535,N_3070,N_3274);
xor U3536 (N_3536,N_3187,N_3079);
nor U3537 (N_3537,N_3415,N_3128);
xor U3538 (N_3538,N_3015,N_3193);
xor U3539 (N_3539,N_3398,N_3296);
and U3540 (N_3540,N_3159,N_3290);
nand U3541 (N_3541,N_3397,N_3103);
or U3542 (N_3542,N_3059,N_3430);
xor U3543 (N_3543,N_3225,N_3277);
xnor U3544 (N_3544,N_3017,N_3419);
xor U3545 (N_3545,N_3256,N_3326);
or U3546 (N_3546,N_3239,N_3052);
and U3547 (N_3547,N_3002,N_3288);
nor U3548 (N_3548,N_3494,N_3085);
xor U3549 (N_3549,N_3302,N_3171);
and U3550 (N_3550,N_3086,N_3388);
or U3551 (N_3551,N_3354,N_3307);
or U3552 (N_3552,N_3358,N_3176);
and U3553 (N_3553,N_3164,N_3350);
and U3554 (N_3554,N_3105,N_3019);
nand U3555 (N_3555,N_3270,N_3265);
nor U3556 (N_3556,N_3384,N_3034);
and U3557 (N_3557,N_3077,N_3402);
xor U3558 (N_3558,N_3414,N_3373);
nand U3559 (N_3559,N_3456,N_3489);
and U3560 (N_3560,N_3149,N_3110);
or U3561 (N_3561,N_3180,N_3395);
and U3562 (N_3562,N_3387,N_3362);
or U3563 (N_3563,N_3032,N_3202);
xor U3564 (N_3564,N_3392,N_3211);
and U3565 (N_3565,N_3163,N_3048);
and U3566 (N_3566,N_3054,N_3196);
or U3567 (N_3567,N_3006,N_3162);
and U3568 (N_3568,N_3024,N_3279);
nand U3569 (N_3569,N_3493,N_3453);
and U3570 (N_3570,N_3040,N_3372);
and U3571 (N_3571,N_3194,N_3416);
and U3572 (N_3572,N_3466,N_3467);
nand U3573 (N_3573,N_3207,N_3191);
nor U3574 (N_3574,N_3136,N_3375);
and U3575 (N_3575,N_3030,N_3368);
or U3576 (N_3576,N_3046,N_3049);
and U3577 (N_3577,N_3316,N_3262);
xor U3578 (N_3578,N_3023,N_3229);
and U3579 (N_3579,N_3205,N_3147);
or U3580 (N_3580,N_3055,N_3013);
nand U3581 (N_3581,N_3473,N_3309);
and U3582 (N_3582,N_3438,N_3390);
and U3583 (N_3583,N_3450,N_3039);
and U3584 (N_3584,N_3168,N_3319);
nand U3585 (N_3585,N_3124,N_3109);
and U3586 (N_3586,N_3078,N_3332);
xor U3587 (N_3587,N_3200,N_3341);
or U3588 (N_3588,N_3081,N_3008);
xnor U3589 (N_3589,N_3238,N_3165);
xnor U3590 (N_3590,N_3401,N_3280);
or U3591 (N_3591,N_3409,N_3069);
nand U3592 (N_3592,N_3071,N_3068);
or U3593 (N_3593,N_3490,N_3499);
and U3594 (N_3594,N_3248,N_3336);
or U3595 (N_3595,N_3252,N_3449);
nand U3596 (N_3596,N_3101,N_3233);
xnor U3597 (N_3597,N_3495,N_3463);
xnor U3598 (N_3598,N_3393,N_3255);
and U3599 (N_3599,N_3357,N_3031);
nor U3600 (N_3600,N_3310,N_3406);
and U3601 (N_3601,N_3488,N_3135);
or U3602 (N_3602,N_3376,N_3367);
nand U3603 (N_3603,N_3464,N_3421);
xor U3604 (N_3604,N_3143,N_3480);
nand U3605 (N_3605,N_3361,N_3083);
xor U3606 (N_3606,N_3383,N_3408);
or U3607 (N_3607,N_3273,N_3042);
xor U3608 (N_3608,N_3011,N_3351);
and U3609 (N_3609,N_3174,N_3064);
nand U3610 (N_3610,N_3269,N_3418);
or U3611 (N_3611,N_3422,N_3072);
or U3612 (N_3612,N_3027,N_3182);
xnor U3613 (N_3613,N_3423,N_3184);
nand U3614 (N_3614,N_3106,N_3304);
nand U3615 (N_3615,N_3366,N_3266);
nor U3616 (N_3616,N_3330,N_3016);
nor U3617 (N_3617,N_3303,N_3245);
xor U3618 (N_3618,N_3313,N_3243);
xnor U3619 (N_3619,N_3212,N_3118);
or U3620 (N_3620,N_3432,N_3022);
and U3621 (N_3621,N_3144,N_3317);
and U3622 (N_3622,N_3146,N_3094);
nor U3623 (N_3623,N_3138,N_3237);
xor U3624 (N_3624,N_3497,N_3206);
xnor U3625 (N_3625,N_3053,N_3108);
or U3626 (N_3626,N_3411,N_3479);
xnor U3627 (N_3627,N_3215,N_3065);
nor U3628 (N_3628,N_3344,N_3218);
and U3629 (N_3629,N_3287,N_3104);
or U3630 (N_3630,N_3271,N_3446);
nor U3631 (N_3631,N_3352,N_3477);
and U3632 (N_3632,N_3257,N_3043);
nand U3633 (N_3633,N_3154,N_3329);
or U3634 (N_3634,N_3155,N_3360);
xor U3635 (N_3635,N_3119,N_3169);
nor U3636 (N_3636,N_3268,N_3377);
nand U3637 (N_3637,N_3074,N_3454);
or U3638 (N_3638,N_3325,N_3457);
and U3639 (N_3639,N_3204,N_3199);
xor U3640 (N_3640,N_3323,N_3151);
xor U3641 (N_3641,N_3063,N_3130);
xnor U3642 (N_3642,N_3349,N_3484);
and U3643 (N_3643,N_3050,N_3095);
or U3644 (N_3644,N_3025,N_3084);
nand U3645 (N_3645,N_3076,N_3338);
nand U3646 (N_3646,N_3192,N_3213);
or U3647 (N_3647,N_3424,N_3334);
nand U3648 (N_3648,N_3041,N_3005);
xor U3649 (N_3649,N_3216,N_3141);
and U3650 (N_3650,N_3152,N_3189);
xnor U3651 (N_3651,N_3481,N_3067);
or U3652 (N_3652,N_3333,N_3492);
nor U3653 (N_3653,N_3431,N_3324);
xor U3654 (N_3654,N_3320,N_3080);
nor U3655 (N_3655,N_3442,N_3188);
nand U3656 (N_3656,N_3440,N_3382);
or U3657 (N_3657,N_3403,N_3223);
nand U3658 (N_3658,N_3133,N_3340);
xor U3659 (N_3659,N_3482,N_3483);
or U3660 (N_3660,N_3486,N_3391);
nor U3661 (N_3661,N_3020,N_3092);
and U3662 (N_3662,N_3246,N_3142);
or U3663 (N_3663,N_3170,N_3498);
and U3664 (N_3664,N_3396,N_3347);
xor U3665 (N_3665,N_3469,N_3369);
xor U3666 (N_3666,N_3236,N_3089);
nor U3667 (N_3667,N_3292,N_3112);
nand U3668 (N_3668,N_3394,N_3443);
and U3669 (N_3669,N_3179,N_3073);
nand U3670 (N_3670,N_3220,N_3161);
or U3671 (N_3671,N_3178,N_3385);
nor U3672 (N_3672,N_3044,N_3098);
and U3673 (N_3673,N_3115,N_3127);
xor U3674 (N_3674,N_3295,N_3364);
or U3675 (N_3675,N_3183,N_3201);
xor U3676 (N_3676,N_3420,N_3434);
xnor U3677 (N_3677,N_3433,N_3389);
xor U3678 (N_3678,N_3380,N_3088);
or U3679 (N_3679,N_3134,N_3308);
or U3680 (N_3680,N_3428,N_3470);
and U3681 (N_3681,N_3012,N_3026);
nor U3682 (N_3682,N_3125,N_3439);
or U3683 (N_3683,N_3462,N_3496);
nor U3684 (N_3684,N_3297,N_3036);
or U3685 (N_3685,N_3298,N_3208);
nand U3686 (N_3686,N_3167,N_3219);
and U3687 (N_3687,N_3253,N_3010);
or U3688 (N_3688,N_3413,N_3276);
xor U3689 (N_3689,N_3491,N_3173);
xnor U3690 (N_3690,N_3410,N_3441);
and U3691 (N_3691,N_3126,N_3460);
nand U3692 (N_3692,N_3242,N_3331);
xnor U3693 (N_3693,N_3417,N_3097);
xor U3694 (N_3694,N_3294,N_3107);
and U3695 (N_3695,N_3284,N_3321);
nand U3696 (N_3696,N_3139,N_3140);
or U3697 (N_3697,N_3061,N_3001);
nor U3698 (N_3698,N_3339,N_3475);
nand U3699 (N_3699,N_3035,N_3378);
or U3700 (N_3700,N_3285,N_3485);
nand U3701 (N_3701,N_3058,N_3150);
nor U3702 (N_3702,N_3045,N_3345);
nand U3703 (N_3703,N_3082,N_3198);
nand U3704 (N_3704,N_3356,N_3289);
nor U3705 (N_3705,N_3327,N_3209);
xnor U3706 (N_3706,N_3145,N_3465);
and U3707 (N_3707,N_3259,N_3459);
and U3708 (N_3708,N_3228,N_3060);
xnor U3709 (N_3709,N_3224,N_3056);
or U3710 (N_3710,N_3240,N_3300);
nand U3711 (N_3711,N_3190,N_3436);
nor U3712 (N_3712,N_3322,N_3203);
or U3713 (N_3713,N_3117,N_3047);
nand U3714 (N_3714,N_3177,N_3227);
or U3715 (N_3715,N_3123,N_3291);
nor U3716 (N_3716,N_3226,N_3359);
and U3717 (N_3717,N_3472,N_3158);
and U3718 (N_3718,N_3235,N_3029);
and U3719 (N_3719,N_3100,N_3099);
xor U3720 (N_3720,N_3381,N_3461);
nand U3721 (N_3721,N_3102,N_3122);
nand U3722 (N_3722,N_3342,N_3004);
and U3723 (N_3723,N_3275,N_3132);
nand U3724 (N_3724,N_3281,N_3263);
nor U3725 (N_3725,N_3210,N_3241);
nor U3726 (N_3726,N_3379,N_3374);
nand U3727 (N_3727,N_3249,N_3429);
nand U3728 (N_3728,N_3234,N_3264);
nor U3729 (N_3729,N_3445,N_3425);
or U3730 (N_3730,N_3311,N_3371);
or U3731 (N_3731,N_3476,N_3386);
nand U3732 (N_3732,N_3400,N_3305);
nor U3733 (N_3733,N_3093,N_3066);
xnor U3734 (N_3734,N_3272,N_3363);
nand U3735 (N_3735,N_3370,N_3247);
xor U3736 (N_3736,N_3113,N_3318);
and U3737 (N_3737,N_3346,N_3328);
nor U3738 (N_3738,N_3451,N_3244);
nor U3739 (N_3739,N_3404,N_3166);
xor U3740 (N_3740,N_3231,N_3222);
or U3741 (N_3741,N_3186,N_3075);
xor U3742 (N_3742,N_3009,N_3195);
xnor U3743 (N_3743,N_3455,N_3437);
nand U3744 (N_3744,N_3214,N_3148);
and U3745 (N_3745,N_3021,N_3251);
and U3746 (N_3746,N_3157,N_3062);
or U3747 (N_3747,N_3116,N_3365);
nand U3748 (N_3748,N_3353,N_3172);
xor U3749 (N_3749,N_3283,N_3299);
nor U3750 (N_3750,N_3230,N_3214);
xnor U3751 (N_3751,N_3157,N_3414);
xor U3752 (N_3752,N_3456,N_3186);
nand U3753 (N_3753,N_3495,N_3096);
and U3754 (N_3754,N_3010,N_3046);
xnor U3755 (N_3755,N_3171,N_3377);
and U3756 (N_3756,N_3104,N_3454);
nor U3757 (N_3757,N_3384,N_3254);
nor U3758 (N_3758,N_3419,N_3165);
nand U3759 (N_3759,N_3362,N_3140);
or U3760 (N_3760,N_3341,N_3347);
or U3761 (N_3761,N_3169,N_3006);
xor U3762 (N_3762,N_3083,N_3297);
nor U3763 (N_3763,N_3483,N_3122);
nand U3764 (N_3764,N_3130,N_3333);
nand U3765 (N_3765,N_3451,N_3288);
nand U3766 (N_3766,N_3317,N_3058);
nor U3767 (N_3767,N_3437,N_3079);
and U3768 (N_3768,N_3359,N_3142);
nand U3769 (N_3769,N_3127,N_3052);
nand U3770 (N_3770,N_3022,N_3305);
nand U3771 (N_3771,N_3403,N_3044);
or U3772 (N_3772,N_3368,N_3298);
and U3773 (N_3773,N_3295,N_3270);
xnor U3774 (N_3774,N_3012,N_3043);
nand U3775 (N_3775,N_3434,N_3040);
and U3776 (N_3776,N_3041,N_3132);
xor U3777 (N_3777,N_3334,N_3482);
nand U3778 (N_3778,N_3464,N_3148);
or U3779 (N_3779,N_3054,N_3443);
or U3780 (N_3780,N_3151,N_3393);
and U3781 (N_3781,N_3451,N_3233);
or U3782 (N_3782,N_3037,N_3034);
or U3783 (N_3783,N_3462,N_3372);
or U3784 (N_3784,N_3260,N_3203);
or U3785 (N_3785,N_3260,N_3487);
nand U3786 (N_3786,N_3032,N_3121);
nand U3787 (N_3787,N_3301,N_3357);
nand U3788 (N_3788,N_3076,N_3343);
nor U3789 (N_3789,N_3015,N_3201);
xnor U3790 (N_3790,N_3304,N_3343);
nor U3791 (N_3791,N_3182,N_3487);
and U3792 (N_3792,N_3140,N_3412);
xnor U3793 (N_3793,N_3074,N_3366);
and U3794 (N_3794,N_3085,N_3042);
and U3795 (N_3795,N_3307,N_3180);
nand U3796 (N_3796,N_3141,N_3328);
nand U3797 (N_3797,N_3332,N_3236);
nand U3798 (N_3798,N_3350,N_3292);
or U3799 (N_3799,N_3049,N_3415);
or U3800 (N_3800,N_3469,N_3161);
and U3801 (N_3801,N_3174,N_3379);
nand U3802 (N_3802,N_3330,N_3059);
and U3803 (N_3803,N_3095,N_3093);
or U3804 (N_3804,N_3304,N_3314);
xnor U3805 (N_3805,N_3329,N_3070);
xor U3806 (N_3806,N_3054,N_3365);
nand U3807 (N_3807,N_3210,N_3473);
xor U3808 (N_3808,N_3153,N_3362);
nand U3809 (N_3809,N_3301,N_3221);
xor U3810 (N_3810,N_3218,N_3325);
or U3811 (N_3811,N_3007,N_3359);
and U3812 (N_3812,N_3113,N_3022);
and U3813 (N_3813,N_3268,N_3398);
or U3814 (N_3814,N_3497,N_3122);
xnor U3815 (N_3815,N_3462,N_3419);
nor U3816 (N_3816,N_3262,N_3204);
or U3817 (N_3817,N_3103,N_3405);
or U3818 (N_3818,N_3168,N_3287);
xnor U3819 (N_3819,N_3377,N_3057);
or U3820 (N_3820,N_3299,N_3305);
nor U3821 (N_3821,N_3288,N_3390);
nor U3822 (N_3822,N_3356,N_3304);
or U3823 (N_3823,N_3317,N_3278);
xnor U3824 (N_3824,N_3107,N_3084);
nand U3825 (N_3825,N_3075,N_3407);
nor U3826 (N_3826,N_3171,N_3435);
nor U3827 (N_3827,N_3316,N_3435);
and U3828 (N_3828,N_3300,N_3214);
xor U3829 (N_3829,N_3261,N_3409);
or U3830 (N_3830,N_3000,N_3064);
nand U3831 (N_3831,N_3032,N_3465);
or U3832 (N_3832,N_3025,N_3127);
nor U3833 (N_3833,N_3464,N_3232);
xnor U3834 (N_3834,N_3071,N_3463);
xnor U3835 (N_3835,N_3062,N_3069);
xnor U3836 (N_3836,N_3013,N_3466);
or U3837 (N_3837,N_3472,N_3477);
nor U3838 (N_3838,N_3256,N_3282);
nand U3839 (N_3839,N_3488,N_3424);
or U3840 (N_3840,N_3320,N_3222);
or U3841 (N_3841,N_3302,N_3289);
and U3842 (N_3842,N_3433,N_3156);
nor U3843 (N_3843,N_3334,N_3104);
nand U3844 (N_3844,N_3174,N_3181);
nor U3845 (N_3845,N_3299,N_3071);
or U3846 (N_3846,N_3391,N_3219);
or U3847 (N_3847,N_3211,N_3255);
nand U3848 (N_3848,N_3402,N_3364);
xor U3849 (N_3849,N_3278,N_3057);
xnor U3850 (N_3850,N_3131,N_3017);
or U3851 (N_3851,N_3059,N_3338);
nor U3852 (N_3852,N_3189,N_3160);
and U3853 (N_3853,N_3254,N_3404);
xor U3854 (N_3854,N_3258,N_3463);
or U3855 (N_3855,N_3239,N_3202);
xor U3856 (N_3856,N_3208,N_3101);
nor U3857 (N_3857,N_3009,N_3035);
xor U3858 (N_3858,N_3414,N_3266);
nor U3859 (N_3859,N_3331,N_3199);
nor U3860 (N_3860,N_3019,N_3402);
or U3861 (N_3861,N_3392,N_3102);
nand U3862 (N_3862,N_3108,N_3106);
nor U3863 (N_3863,N_3446,N_3304);
or U3864 (N_3864,N_3192,N_3470);
nor U3865 (N_3865,N_3245,N_3233);
or U3866 (N_3866,N_3007,N_3468);
nor U3867 (N_3867,N_3102,N_3091);
nor U3868 (N_3868,N_3067,N_3463);
or U3869 (N_3869,N_3379,N_3419);
or U3870 (N_3870,N_3205,N_3332);
and U3871 (N_3871,N_3042,N_3416);
or U3872 (N_3872,N_3213,N_3470);
nand U3873 (N_3873,N_3123,N_3341);
nand U3874 (N_3874,N_3393,N_3057);
nor U3875 (N_3875,N_3377,N_3023);
xor U3876 (N_3876,N_3311,N_3219);
and U3877 (N_3877,N_3425,N_3186);
or U3878 (N_3878,N_3125,N_3462);
or U3879 (N_3879,N_3463,N_3129);
nand U3880 (N_3880,N_3396,N_3376);
nand U3881 (N_3881,N_3301,N_3447);
nand U3882 (N_3882,N_3089,N_3306);
or U3883 (N_3883,N_3436,N_3359);
xnor U3884 (N_3884,N_3029,N_3246);
nor U3885 (N_3885,N_3032,N_3016);
nor U3886 (N_3886,N_3427,N_3096);
and U3887 (N_3887,N_3376,N_3473);
xor U3888 (N_3888,N_3136,N_3196);
nand U3889 (N_3889,N_3197,N_3380);
nand U3890 (N_3890,N_3244,N_3441);
xnor U3891 (N_3891,N_3437,N_3258);
and U3892 (N_3892,N_3336,N_3328);
nand U3893 (N_3893,N_3087,N_3340);
or U3894 (N_3894,N_3372,N_3365);
or U3895 (N_3895,N_3322,N_3006);
nor U3896 (N_3896,N_3460,N_3310);
xor U3897 (N_3897,N_3239,N_3000);
nor U3898 (N_3898,N_3174,N_3176);
xnor U3899 (N_3899,N_3373,N_3076);
or U3900 (N_3900,N_3185,N_3465);
nor U3901 (N_3901,N_3325,N_3370);
nor U3902 (N_3902,N_3079,N_3236);
and U3903 (N_3903,N_3093,N_3479);
or U3904 (N_3904,N_3149,N_3395);
and U3905 (N_3905,N_3011,N_3029);
nor U3906 (N_3906,N_3412,N_3306);
nor U3907 (N_3907,N_3015,N_3398);
xor U3908 (N_3908,N_3479,N_3275);
and U3909 (N_3909,N_3403,N_3011);
nor U3910 (N_3910,N_3391,N_3287);
nor U3911 (N_3911,N_3351,N_3244);
or U3912 (N_3912,N_3117,N_3144);
and U3913 (N_3913,N_3143,N_3206);
or U3914 (N_3914,N_3007,N_3344);
xor U3915 (N_3915,N_3497,N_3463);
xnor U3916 (N_3916,N_3041,N_3456);
xnor U3917 (N_3917,N_3079,N_3348);
and U3918 (N_3918,N_3136,N_3011);
and U3919 (N_3919,N_3292,N_3186);
or U3920 (N_3920,N_3330,N_3216);
or U3921 (N_3921,N_3328,N_3168);
nand U3922 (N_3922,N_3024,N_3048);
or U3923 (N_3923,N_3190,N_3388);
or U3924 (N_3924,N_3014,N_3042);
or U3925 (N_3925,N_3428,N_3253);
xnor U3926 (N_3926,N_3056,N_3378);
nand U3927 (N_3927,N_3356,N_3402);
nor U3928 (N_3928,N_3037,N_3145);
xor U3929 (N_3929,N_3222,N_3446);
nor U3930 (N_3930,N_3116,N_3086);
nor U3931 (N_3931,N_3329,N_3306);
or U3932 (N_3932,N_3377,N_3160);
nor U3933 (N_3933,N_3081,N_3158);
or U3934 (N_3934,N_3413,N_3049);
and U3935 (N_3935,N_3489,N_3302);
or U3936 (N_3936,N_3268,N_3272);
xnor U3937 (N_3937,N_3108,N_3391);
nor U3938 (N_3938,N_3224,N_3436);
and U3939 (N_3939,N_3428,N_3257);
nand U3940 (N_3940,N_3383,N_3428);
nor U3941 (N_3941,N_3276,N_3269);
nand U3942 (N_3942,N_3011,N_3247);
or U3943 (N_3943,N_3061,N_3158);
or U3944 (N_3944,N_3116,N_3136);
xnor U3945 (N_3945,N_3175,N_3119);
and U3946 (N_3946,N_3182,N_3294);
or U3947 (N_3947,N_3183,N_3355);
xnor U3948 (N_3948,N_3205,N_3124);
and U3949 (N_3949,N_3278,N_3209);
or U3950 (N_3950,N_3334,N_3447);
nor U3951 (N_3951,N_3389,N_3341);
and U3952 (N_3952,N_3272,N_3442);
nor U3953 (N_3953,N_3219,N_3122);
nand U3954 (N_3954,N_3178,N_3279);
xor U3955 (N_3955,N_3442,N_3388);
nand U3956 (N_3956,N_3383,N_3455);
nor U3957 (N_3957,N_3337,N_3352);
nand U3958 (N_3958,N_3473,N_3275);
xor U3959 (N_3959,N_3336,N_3456);
and U3960 (N_3960,N_3395,N_3480);
nand U3961 (N_3961,N_3111,N_3184);
or U3962 (N_3962,N_3107,N_3372);
nor U3963 (N_3963,N_3361,N_3165);
nand U3964 (N_3964,N_3183,N_3454);
nand U3965 (N_3965,N_3307,N_3059);
xor U3966 (N_3966,N_3411,N_3494);
xnor U3967 (N_3967,N_3341,N_3104);
nor U3968 (N_3968,N_3177,N_3411);
or U3969 (N_3969,N_3256,N_3263);
xnor U3970 (N_3970,N_3162,N_3231);
nand U3971 (N_3971,N_3424,N_3218);
nand U3972 (N_3972,N_3200,N_3033);
nand U3973 (N_3973,N_3206,N_3129);
or U3974 (N_3974,N_3054,N_3244);
nand U3975 (N_3975,N_3385,N_3161);
xnor U3976 (N_3976,N_3052,N_3266);
and U3977 (N_3977,N_3370,N_3442);
or U3978 (N_3978,N_3113,N_3191);
and U3979 (N_3979,N_3008,N_3165);
nor U3980 (N_3980,N_3311,N_3487);
or U3981 (N_3981,N_3049,N_3068);
nand U3982 (N_3982,N_3045,N_3334);
nor U3983 (N_3983,N_3061,N_3028);
xor U3984 (N_3984,N_3101,N_3032);
nor U3985 (N_3985,N_3351,N_3328);
or U3986 (N_3986,N_3426,N_3409);
xor U3987 (N_3987,N_3252,N_3175);
or U3988 (N_3988,N_3263,N_3197);
xnor U3989 (N_3989,N_3305,N_3245);
nand U3990 (N_3990,N_3184,N_3419);
or U3991 (N_3991,N_3230,N_3211);
nand U3992 (N_3992,N_3175,N_3218);
or U3993 (N_3993,N_3301,N_3176);
nand U3994 (N_3994,N_3391,N_3091);
or U3995 (N_3995,N_3198,N_3142);
and U3996 (N_3996,N_3473,N_3050);
and U3997 (N_3997,N_3049,N_3064);
and U3998 (N_3998,N_3068,N_3359);
xor U3999 (N_3999,N_3279,N_3383);
or U4000 (N_4000,N_3925,N_3633);
or U4001 (N_4001,N_3806,N_3675);
nand U4002 (N_4002,N_3501,N_3653);
xor U4003 (N_4003,N_3708,N_3683);
nand U4004 (N_4004,N_3737,N_3640);
nor U4005 (N_4005,N_3868,N_3790);
nor U4006 (N_4006,N_3978,N_3884);
nor U4007 (N_4007,N_3687,N_3605);
xnor U4008 (N_4008,N_3814,N_3587);
nor U4009 (N_4009,N_3541,N_3982);
or U4010 (N_4010,N_3970,N_3942);
or U4011 (N_4011,N_3503,N_3515);
or U4012 (N_4012,N_3718,N_3817);
nor U4013 (N_4013,N_3983,N_3971);
nor U4014 (N_4014,N_3957,N_3592);
or U4015 (N_4015,N_3599,N_3873);
or U4016 (N_4016,N_3664,N_3616);
xor U4017 (N_4017,N_3972,N_3899);
nor U4018 (N_4018,N_3935,N_3560);
and U4019 (N_4019,N_3980,N_3837);
xnor U4020 (N_4020,N_3967,N_3938);
nor U4021 (N_4021,N_3870,N_3529);
nand U4022 (N_4022,N_3630,N_3584);
or U4023 (N_4023,N_3966,N_3569);
nor U4024 (N_4024,N_3857,N_3841);
or U4025 (N_4025,N_3830,N_3949);
nand U4026 (N_4026,N_3840,N_3694);
xor U4027 (N_4027,N_3792,N_3937);
xor U4028 (N_4028,N_3712,N_3676);
or U4029 (N_4029,N_3988,N_3845);
xor U4030 (N_4030,N_3717,N_3741);
and U4031 (N_4031,N_3991,N_3822);
and U4032 (N_4032,N_3839,N_3920);
xor U4033 (N_4033,N_3586,N_3593);
and U4034 (N_4034,N_3698,N_3934);
or U4035 (N_4035,N_3849,N_3753);
or U4036 (N_4036,N_3827,N_3521);
nand U4037 (N_4037,N_3953,N_3848);
nand U4038 (N_4038,N_3894,N_3582);
and U4039 (N_4039,N_3716,N_3754);
xnor U4040 (N_4040,N_3766,N_3581);
xnor U4041 (N_4041,N_3929,N_3546);
or U4042 (N_4042,N_3910,N_3617);
nand U4043 (N_4043,N_3629,N_3862);
xor U4044 (N_4044,N_3921,N_3940);
or U4045 (N_4045,N_3787,N_3877);
or U4046 (N_4046,N_3583,N_3656);
or U4047 (N_4047,N_3986,N_3740);
xor U4048 (N_4048,N_3665,N_3891);
or U4049 (N_4049,N_3504,N_3872);
nand U4050 (N_4050,N_3632,N_3644);
nor U4051 (N_4051,N_3707,N_3819);
nand U4052 (N_4052,N_3695,N_3906);
and U4053 (N_4053,N_3522,N_3526);
or U4054 (N_4054,N_3607,N_3936);
nand U4055 (N_4055,N_3709,N_3770);
or U4056 (N_4056,N_3506,N_3677);
nand U4057 (N_4057,N_3610,N_3693);
xnor U4058 (N_4058,N_3730,N_3543);
nand U4059 (N_4059,N_3844,N_3537);
nor U4060 (N_4060,N_3525,N_3650);
xor U4061 (N_4061,N_3674,N_3763);
nand U4062 (N_4062,N_3828,N_3671);
xor U4063 (N_4063,N_3829,N_3775);
or U4064 (N_4064,N_3811,N_3952);
nand U4065 (N_4065,N_3643,N_3851);
and U4066 (N_4066,N_3636,N_3500);
nor U4067 (N_4067,N_3897,N_3551);
nor U4068 (N_4068,N_3590,N_3803);
nor U4069 (N_4069,N_3502,N_3878);
or U4070 (N_4070,N_3977,N_3756);
or U4071 (N_4071,N_3946,N_3686);
xnor U4072 (N_4072,N_3659,N_3696);
or U4073 (N_4073,N_3947,N_3784);
nor U4074 (N_4074,N_3963,N_3507);
or U4075 (N_4075,N_3706,N_3669);
xor U4076 (N_4076,N_3945,N_3511);
nor U4077 (N_4077,N_3612,N_3679);
nand U4078 (N_4078,N_3725,N_3833);
nand U4079 (N_4079,N_3987,N_3818);
xor U4080 (N_4080,N_3777,N_3533);
or U4081 (N_4081,N_3520,N_3611);
or U4082 (N_4082,N_3514,N_3743);
xnor U4083 (N_4083,N_3700,N_3585);
nor U4084 (N_4084,N_3580,N_3747);
nand U4085 (N_4085,N_3749,N_3997);
nand U4086 (N_4086,N_3961,N_3875);
nor U4087 (N_4087,N_3524,N_3867);
and U4088 (N_4088,N_3703,N_3994);
or U4089 (N_4089,N_3579,N_3981);
nor U4090 (N_4090,N_3745,N_3542);
xnor U4091 (N_4091,N_3859,N_3668);
nand U4092 (N_4092,N_3536,N_3785);
nand U4093 (N_4093,N_3815,N_3689);
xor U4094 (N_4094,N_3655,N_3638);
or U4095 (N_4095,N_3760,N_3780);
xnor U4096 (N_4096,N_3768,N_3562);
nor U4097 (N_4097,N_3588,N_3911);
or U4098 (N_4098,N_3681,N_3869);
or U4099 (N_4099,N_3736,N_3879);
nand U4100 (N_4100,N_3534,N_3619);
nor U4101 (N_4101,N_3842,N_3765);
or U4102 (N_4102,N_3758,N_3606);
or U4103 (N_4103,N_3998,N_3751);
and U4104 (N_4104,N_3888,N_3850);
and U4105 (N_4105,N_3701,N_3820);
xnor U4106 (N_4106,N_3672,N_3527);
xnor U4107 (N_4107,N_3547,N_3923);
nand U4108 (N_4108,N_3578,N_3834);
xor U4109 (N_4109,N_3955,N_3532);
and U4110 (N_4110,N_3904,N_3623);
nor U4111 (N_4111,N_3889,N_3565);
or U4112 (N_4112,N_3575,N_3666);
xor U4113 (N_4113,N_3720,N_3864);
or U4114 (N_4114,N_3965,N_3908);
nor U4115 (N_4115,N_3791,N_3890);
nor U4116 (N_4116,N_3762,N_3809);
nand U4117 (N_4117,N_3715,N_3926);
or U4118 (N_4118,N_3558,N_3801);
nand U4119 (N_4119,N_3528,N_3846);
xnor U4120 (N_4120,N_3985,N_3727);
xor U4121 (N_4121,N_3723,N_3519);
or U4122 (N_4122,N_3613,N_3721);
or U4123 (N_4123,N_3789,N_3959);
nand U4124 (N_4124,N_3895,N_3928);
xnor U4125 (N_4125,N_3748,N_3788);
nand U4126 (N_4126,N_3932,N_3549);
nor U4127 (N_4127,N_3734,N_3711);
nand U4128 (N_4128,N_3648,N_3944);
xor U4129 (N_4129,N_3905,N_3861);
nand U4130 (N_4130,N_3692,N_3571);
and U4131 (N_4131,N_3847,N_3783);
or U4132 (N_4132,N_3962,N_3512);
or U4133 (N_4133,N_3603,N_3535);
nor U4134 (N_4134,N_3805,N_3728);
and U4135 (N_4135,N_3996,N_3724);
or U4136 (N_4136,N_3572,N_3950);
or U4137 (N_4137,N_3931,N_3639);
and U4138 (N_4138,N_3954,N_3979);
xor U4139 (N_4139,N_3568,N_3854);
and U4140 (N_4140,N_3880,N_3968);
xor U4141 (N_4141,N_3634,N_3913);
nand U4142 (N_4142,N_3812,N_3685);
nand U4143 (N_4143,N_3604,N_3750);
nand U4144 (N_4144,N_3976,N_3662);
nor U4145 (N_4145,N_3802,N_3807);
or U4146 (N_4146,N_3793,N_3800);
xor U4147 (N_4147,N_3622,N_3804);
nor U4148 (N_4148,N_3919,N_3600);
and U4149 (N_4149,N_3796,N_3596);
nand U4150 (N_4150,N_3999,N_3538);
or U4151 (N_4151,N_3559,N_3641);
and U4152 (N_4152,N_3898,N_3513);
and U4153 (N_4153,N_3903,N_3984);
nor U4154 (N_4154,N_3719,N_3699);
nand U4155 (N_4155,N_3948,N_3647);
nor U4156 (N_4156,N_3915,N_3651);
xnor U4157 (N_4157,N_3660,N_3798);
or U4158 (N_4158,N_3990,N_3794);
nor U4159 (N_4159,N_3530,N_3975);
xor U4160 (N_4160,N_3958,N_3769);
or U4161 (N_4161,N_3702,N_3732);
nand U4162 (N_4162,N_3539,N_3645);
nand U4163 (N_4163,N_3620,N_3658);
xnor U4164 (N_4164,N_3509,N_3757);
nand U4165 (N_4165,N_3821,N_3912);
or U4166 (N_4166,N_3667,N_3993);
or U4167 (N_4167,N_3924,N_3893);
nand U4168 (N_4168,N_3799,N_3939);
or U4169 (N_4169,N_3597,N_3782);
and U4170 (N_4170,N_3714,N_3518);
xnor U4171 (N_4171,N_3927,N_3823);
and U4172 (N_4172,N_3776,N_3544);
nor U4173 (N_4173,N_3508,N_3637);
and U4174 (N_4174,N_3900,N_3673);
and U4175 (N_4175,N_3505,N_3609);
and U4176 (N_4176,N_3855,N_3810);
nand U4177 (N_4177,N_3545,N_3726);
nand U4178 (N_4178,N_3836,N_3557);
nor U4179 (N_4179,N_3646,N_3523);
xnor U4180 (N_4180,N_3863,N_3556);
nor U4181 (N_4181,N_3914,N_3614);
and U4182 (N_4182,N_3853,N_3813);
nor U4183 (N_4183,N_3824,N_3601);
and U4184 (N_4184,N_3553,N_3767);
and U4185 (N_4185,N_3883,N_3866);
nand U4186 (N_4186,N_3941,N_3690);
xor U4187 (N_4187,N_3567,N_3627);
xnor U4188 (N_4188,N_3602,N_3826);
nor U4189 (N_4189,N_3995,N_3779);
or U4190 (N_4190,N_3552,N_3550);
and U4191 (N_4191,N_3577,N_3843);
nor U4192 (N_4192,N_3781,N_3680);
nand U4193 (N_4193,N_3704,N_3631);
xor U4194 (N_4194,N_3684,N_3901);
or U4195 (N_4195,N_3956,N_3852);
nor U4196 (N_4196,N_3682,N_3570);
and U4197 (N_4197,N_3598,N_3896);
or U4198 (N_4198,N_3835,N_3886);
xor U4199 (N_4199,N_3531,N_3710);
nand U4200 (N_4200,N_3739,N_3786);
xor U4201 (N_4201,N_3917,N_3621);
nand U4202 (N_4202,N_3759,N_3576);
nor U4203 (N_4203,N_3729,N_3831);
nor U4204 (N_4204,N_3755,N_3573);
and U4205 (N_4205,N_3738,N_3973);
nor U4206 (N_4206,N_3874,N_3772);
nor U4207 (N_4207,N_3635,N_3663);
or U4208 (N_4208,N_3858,N_3892);
xnor U4209 (N_4209,N_3881,N_3642);
xor U4210 (N_4210,N_3918,N_3554);
nor U4211 (N_4211,N_3774,N_3628);
xor U4212 (N_4212,N_3742,N_3566);
xor U4213 (N_4213,N_3618,N_3561);
and U4214 (N_4214,N_3649,N_3625);
nand U4215 (N_4215,N_3885,N_3691);
nor U4216 (N_4216,N_3902,N_3816);
xor U4217 (N_4217,N_3916,N_3865);
or U4218 (N_4218,N_3746,N_3555);
nor U4219 (N_4219,N_3797,N_3933);
or U4220 (N_4220,N_3960,N_3654);
or U4221 (N_4221,N_3517,N_3969);
nor U4222 (N_4222,N_3657,N_3697);
nor U4223 (N_4223,N_3856,N_3773);
nor U4224 (N_4224,N_3761,N_3992);
and U4225 (N_4225,N_3989,N_3907);
or U4226 (N_4226,N_3778,N_3615);
nand U4227 (N_4227,N_3882,N_3808);
xnor U4228 (N_4228,N_3733,N_3731);
nand U4229 (N_4229,N_3838,N_3832);
nand U4230 (N_4230,N_3930,N_3688);
or U4231 (N_4231,N_3964,N_3661);
or U4232 (N_4232,N_3510,N_3876);
and U4233 (N_4233,N_3670,N_3764);
nor U4234 (N_4234,N_3887,N_3744);
nor U4235 (N_4235,N_3735,N_3624);
nand U4236 (N_4236,N_3871,N_3860);
or U4237 (N_4237,N_3595,N_3795);
or U4238 (N_4238,N_3652,N_3722);
nand U4239 (N_4239,N_3563,N_3825);
nor U4240 (N_4240,N_3594,N_3574);
and U4241 (N_4241,N_3591,N_3922);
or U4242 (N_4242,N_3909,N_3974);
nand U4243 (N_4243,N_3705,N_3713);
xor U4244 (N_4244,N_3564,N_3608);
nand U4245 (N_4245,N_3752,N_3589);
or U4246 (N_4246,N_3678,N_3540);
nand U4247 (N_4247,N_3626,N_3943);
xor U4248 (N_4248,N_3548,N_3516);
and U4249 (N_4249,N_3951,N_3771);
nand U4250 (N_4250,N_3988,N_3980);
or U4251 (N_4251,N_3637,N_3530);
nor U4252 (N_4252,N_3923,N_3795);
nand U4253 (N_4253,N_3765,N_3739);
nand U4254 (N_4254,N_3648,N_3924);
xnor U4255 (N_4255,N_3534,N_3963);
and U4256 (N_4256,N_3566,N_3525);
or U4257 (N_4257,N_3839,N_3785);
xor U4258 (N_4258,N_3767,N_3514);
and U4259 (N_4259,N_3936,N_3729);
nor U4260 (N_4260,N_3982,N_3544);
nand U4261 (N_4261,N_3732,N_3917);
xnor U4262 (N_4262,N_3907,N_3942);
and U4263 (N_4263,N_3710,N_3553);
nor U4264 (N_4264,N_3748,N_3575);
xor U4265 (N_4265,N_3713,N_3992);
xnor U4266 (N_4266,N_3683,N_3841);
nand U4267 (N_4267,N_3846,N_3770);
or U4268 (N_4268,N_3899,N_3716);
and U4269 (N_4269,N_3890,N_3736);
nor U4270 (N_4270,N_3801,N_3886);
or U4271 (N_4271,N_3890,N_3899);
xnor U4272 (N_4272,N_3743,N_3814);
nand U4273 (N_4273,N_3500,N_3522);
and U4274 (N_4274,N_3858,N_3812);
xor U4275 (N_4275,N_3996,N_3515);
xor U4276 (N_4276,N_3576,N_3978);
xor U4277 (N_4277,N_3572,N_3600);
xor U4278 (N_4278,N_3631,N_3811);
xor U4279 (N_4279,N_3655,N_3833);
xor U4280 (N_4280,N_3615,N_3620);
or U4281 (N_4281,N_3502,N_3621);
nor U4282 (N_4282,N_3610,N_3935);
xor U4283 (N_4283,N_3539,N_3651);
xnor U4284 (N_4284,N_3623,N_3951);
and U4285 (N_4285,N_3672,N_3757);
and U4286 (N_4286,N_3524,N_3821);
nor U4287 (N_4287,N_3667,N_3890);
or U4288 (N_4288,N_3869,N_3745);
xor U4289 (N_4289,N_3983,N_3623);
and U4290 (N_4290,N_3856,N_3849);
and U4291 (N_4291,N_3960,N_3728);
and U4292 (N_4292,N_3559,N_3804);
or U4293 (N_4293,N_3929,N_3921);
xor U4294 (N_4294,N_3609,N_3860);
xor U4295 (N_4295,N_3935,N_3573);
and U4296 (N_4296,N_3984,N_3949);
xor U4297 (N_4297,N_3548,N_3500);
and U4298 (N_4298,N_3754,N_3747);
or U4299 (N_4299,N_3648,N_3900);
xor U4300 (N_4300,N_3818,N_3675);
or U4301 (N_4301,N_3879,N_3560);
and U4302 (N_4302,N_3511,N_3679);
xnor U4303 (N_4303,N_3572,N_3903);
nand U4304 (N_4304,N_3820,N_3731);
and U4305 (N_4305,N_3589,N_3559);
or U4306 (N_4306,N_3553,N_3802);
and U4307 (N_4307,N_3673,N_3988);
nor U4308 (N_4308,N_3889,N_3895);
nand U4309 (N_4309,N_3616,N_3827);
or U4310 (N_4310,N_3636,N_3503);
and U4311 (N_4311,N_3856,N_3682);
nand U4312 (N_4312,N_3985,N_3942);
xor U4313 (N_4313,N_3744,N_3627);
and U4314 (N_4314,N_3552,N_3991);
nor U4315 (N_4315,N_3905,N_3723);
and U4316 (N_4316,N_3884,N_3742);
and U4317 (N_4317,N_3617,N_3854);
nand U4318 (N_4318,N_3929,N_3979);
nor U4319 (N_4319,N_3887,N_3953);
nand U4320 (N_4320,N_3661,N_3688);
nor U4321 (N_4321,N_3660,N_3610);
or U4322 (N_4322,N_3889,N_3954);
xnor U4323 (N_4323,N_3878,N_3937);
and U4324 (N_4324,N_3891,N_3977);
nor U4325 (N_4325,N_3677,N_3562);
and U4326 (N_4326,N_3792,N_3715);
xnor U4327 (N_4327,N_3705,N_3967);
or U4328 (N_4328,N_3547,N_3571);
and U4329 (N_4329,N_3998,N_3609);
xnor U4330 (N_4330,N_3595,N_3701);
nor U4331 (N_4331,N_3503,N_3530);
nor U4332 (N_4332,N_3770,N_3509);
nor U4333 (N_4333,N_3746,N_3868);
nor U4334 (N_4334,N_3630,N_3912);
nor U4335 (N_4335,N_3929,N_3843);
and U4336 (N_4336,N_3562,N_3681);
and U4337 (N_4337,N_3555,N_3907);
and U4338 (N_4338,N_3791,N_3708);
or U4339 (N_4339,N_3916,N_3563);
xnor U4340 (N_4340,N_3900,N_3621);
nand U4341 (N_4341,N_3930,N_3876);
and U4342 (N_4342,N_3550,N_3780);
nor U4343 (N_4343,N_3673,N_3650);
or U4344 (N_4344,N_3857,N_3579);
nor U4345 (N_4345,N_3729,N_3797);
or U4346 (N_4346,N_3559,N_3604);
nor U4347 (N_4347,N_3799,N_3684);
or U4348 (N_4348,N_3631,N_3978);
and U4349 (N_4349,N_3856,N_3526);
nand U4350 (N_4350,N_3898,N_3878);
nand U4351 (N_4351,N_3969,N_3759);
xor U4352 (N_4352,N_3636,N_3596);
and U4353 (N_4353,N_3574,N_3645);
nand U4354 (N_4354,N_3802,N_3717);
nand U4355 (N_4355,N_3553,N_3772);
nand U4356 (N_4356,N_3828,N_3818);
nand U4357 (N_4357,N_3912,N_3504);
or U4358 (N_4358,N_3850,N_3953);
or U4359 (N_4359,N_3550,N_3791);
xnor U4360 (N_4360,N_3783,N_3952);
nand U4361 (N_4361,N_3875,N_3635);
and U4362 (N_4362,N_3819,N_3887);
or U4363 (N_4363,N_3686,N_3963);
xnor U4364 (N_4364,N_3601,N_3641);
nor U4365 (N_4365,N_3734,N_3760);
xnor U4366 (N_4366,N_3534,N_3958);
nor U4367 (N_4367,N_3775,N_3833);
or U4368 (N_4368,N_3983,N_3560);
or U4369 (N_4369,N_3957,N_3729);
xor U4370 (N_4370,N_3889,N_3662);
nand U4371 (N_4371,N_3883,N_3777);
or U4372 (N_4372,N_3714,N_3998);
nor U4373 (N_4373,N_3807,N_3626);
and U4374 (N_4374,N_3786,N_3827);
or U4375 (N_4375,N_3928,N_3824);
nor U4376 (N_4376,N_3982,N_3575);
xor U4377 (N_4377,N_3990,N_3869);
or U4378 (N_4378,N_3507,N_3785);
or U4379 (N_4379,N_3954,N_3851);
xor U4380 (N_4380,N_3751,N_3666);
nand U4381 (N_4381,N_3935,N_3899);
nor U4382 (N_4382,N_3553,N_3993);
or U4383 (N_4383,N_3524,N_3783);
and U4384 (N_4384,N_3965,N_3636);
or U4385 (N_4385,N_3888,N_3944);
xor U4386 (N_4386,N_3873,N_3552);
or U4387 (N_4387,N_3579,N_3826);
nand U4388 (N_4388,N_3728,N_3828);
or U4389 (N_4389,N_3700,N_3798);
or U4390 (N_4390,N_3621,N_3645);
nand U4391 (N_4391,N_3589,N_3688);
nand U4392 (N_4392,N_3770,N_3940);
or U4393 (N_4393,N_3766,N_3993);
nor U4394 (N_4394,N_3660,N_3716);
or U4395 (N_4395,N_3866,N_3570);
nor U4396 (N_4396,N_3939,N_3854);
or U4397 (N_4397,N_3924,N_3626);
nand U4398 (N_4398,N_3636,N_3910);
or U4399 (N_4399,N_3596,N_3917);
nor U4400 (N_4400,N_3500,N_3549);
or U4401 (N_4401,N_3560,N_3980);
and U4402 (N_4402,N_3818,N_3854);
nand U4403 (N_4403,N_3677,N_3652);
nor U4404 (N_4404,N_3927,N_3827);
nor U4405 (N_4405,N_3678,N_3727);
or U4406 (N_4406,N_3652,N_3736);
nor U4407 (N_4407,N_3907,N_3559);
and U4408 (N_4408,N_3986,N_3571);
xnor U4409 (N_4409,N_3994,N_3830);
nor U4410 (N_4410,N_3804,N_3915);
and U4411 (N_4411,N_3950,N_3671);
nand U4412 (N_4412,N_3557,N_3903);
nor U4413 (N_4413,N_3575,N_3532);
nand U4414 (N_4414,N_3798,N_3856);
nor U4415 (N_4415,N_3948,N_3705);
or U4416 (N_4416,N_3513,N_3673);
and U4417 (N_4417,N_3757,N_3514);
nor U4418 (N_4418,N_3675,N_3683);
xnor U4419 (N_4419,N_3795,N_3935);
nor U4420 (N_4420,N_3824,N_3916);
nor U4421 (N_4421,N_3609,N_3559);
xnor U4422 (N_4422,N_3663,N_3626);
nor U4423 (N_4423,N_3695,N_3615);
and U4424 (N_4424,N_3650,N_3644);
or U4425 (N_4425,N_3505,N_3784);
nand U4426 (N_4426,N_3568,N_3705);
nor U4427 (N_4427,N_3594,N_3912);
and U4428 (N_4428,N_3534,N_3648);
and U4429 (N_4429,N_3878,N_3523);
nand U4430 (N_4430,N_3996,N_3711);
nor U4431 (N_4431,N_3515,N_3944);
nor U4432 (N_4432,N_3737,N_3767);
and U4433 (N_4433,N_3619,N_3966);
nand U4434 (N_4434,N_3717,N_3911);
or U4435 (N_4435,N_3886,N_3981);
nand U4436 (N_4436,N_3811,N_3804);
xor U4437 (N_4437,N_3944,N_3694);
or U4438 (N_4438,N_3866,N_3943);
and U4439 (N_4439,N_3780,N_3772);
or U4440 (N_4440,N_3557,N_3780);
or U4441 (N_4441,N_3623,N_3716);
or U4442 (N_4442,N_3966,N_3961);
or U4443 (N_4443,N_3597,N_3910);
and U4444 (N_4444,N_3815,N_3804);
xor U4445 (N_4445,N_3750,N_3830);
nand U4446 (N_4446,N_3851,N_3805);
nand U4447 (N_4447,N_3645,N_3671);
or U4448 (N_4448,N_3799,N_3529);
nor U4449 (N_4449,N_3505,N_3686);
and U4450 (N_4450,N_3656,N_3635);
and U4451 (N_4451,N_3770,N_3564);
xnor U4452 (N_4452,N_3703,N_3554);
or U4453 (N_4453,N_3807,N_3625);
nand U4454 (N_4454,N_3785,N_3520);
xnor U4455 (N_4455,N_3551,N_3821);
xnor U4456 (N_4456,N_3999,N_3703);
nor U4457 (N_4457,N_3937,N_3916);
and U4458 (N_4458,N_3612,N_3873);
and U4459 (N_4459,N_3683,N_3818);
or U4460 (N_4460,N_3997,N_3580);
and U4461 (N_4461,N_3547,N_3740);
and U4462 (N_4462,N_3726,N_3877);
xnor U4463 (N_4463,N_3962,N_3718);
nand U4464 (N_4464,N_3980,N_3546);
nand U4465 (N_4465,N_3942,N_3662);
nor U4466 (N_4466,N_3516,N_3789);
nor U4467 (N_4467,N_3877,N_3987);
nand U4468 (N_4468,N_3556,N_3630);
or U4469 (N_4469,N_3901,N_3660);
xnor U4470 (N_4470,N_3937,N_3616);
or U4471 (N_4471,N_3696,N_3809);
nand U4472 (N_4472,N_3957,N_3876);
and U4473 (N_4473,N_3773,N_3913);
or U4474 (N_4474,N_3980,N_3825);
nor U4475 (N_4475,N_3998,N_3902);
nor U4476 (N_4476,N_3769,N_3722);
xor U4477 (N_4477,N_3605,N_3694);
nand U4478 (N_4478,N_3859,N_3878);
nand U4479 (N_4479,N_3873,N_3678);
or U4480 (N_4480,N_3551,N_3674);
xor U4481 (N_4481,N_3878,N_3672);
xor U4482 (N_4482,N_3603,N_3900);
or U4483 (N_4483,N_3745,N_3820);
nand U4484 (N_4484,N_3629,N_3520);
nor U4485 (N_4485,N_3543,N_3714);
nor U4486 (N_4486,N_3625,N_3835);
nor U4487 (N_4487,N_3700,N_3772);
or U4488 (N_4488,N_3563,N_3621);
nand U4489 (N_4489,N_3710,N_3573);
nor U4490 (N_4490,N_3582,N_3907);
nand U4491 (N_4491,N_3572,N_3987);
xnor U4492 (N_4492,N_3625,N_3720);
nor U4493 (N_4493,N_3638,N_3888);
xor U4494 (N_4494,N_3885,N_3593);
or U4495 (N_4495,N_3723,N_3729);
nor U4496 (N_4496,N_3828,N_3805);
nand U4497 (N_4497,N_3644,N_3717);
xor U4498 (N_4498,N_3987,N_3575);
nor U4499 (N_4499,N_3660,N_3872);
nand U4500 (N_4500,N_4474,N_4094);
or U4501 (N_4501,N_4318,N_4475);
nor U4502 (N_4502,N_4031,N_4007);
nor U4503 (N_4503,N_4411,N_4317);
nor U4504 (N_4504,N_4446,N_4419);
and U4505 (N_4505,N_4357,N_4280);
xnor U4506 (N_4506,N_4493,N_4195);
xnor U4507 (N_4507,N_4012,N_4454);
and U4508 (N_4508,N_4127,N_4128);
nor U4509 (N_4509,N_4371,N_4078);
or U4510 (N_4510,N_4131,N_4458);
nand U4511 (N_4511,N_4499,N_4162);
xor U4512 (N_4512,N_4457,N_4402);
or U4513 (N_4513,N_4145,N_4141);
or U4514 (N_4514,N_4441,N_4137);
and U4515 (N_4515,N_4027,N_4358);
nor U4516 (N_4516,N_4050,N_4235);
nand U4517 (N_4517,N_4146,N_4334);
and U4518 (N_4518,N_4498,N_4006);
or U4519 (N_4519,N_4108,N_4172);
nand U4520 (N_4520,N_4427,N_4183);
nor U4521 (N_4521,N_4226,N_4210);
and U4522 (N_4522,N_4477,N_4372);
xor U4523 (N_4523,N_4169,N_4250);
xnor U4524 (N_4524,N_4433,N_4016);
and U4525 (N_4525,N_4177,N_4439);
or U4526 (N_4526,N_4001,N_4236);
xor U4527 (N_4527,N_4018,N_4178);
and U4528 (N_4528,N_4289,N_4034);
nand U4529 (N_4529,N_4201,N_4174);
and U4530 (N_4530,N_4426,N_4438);
or U4531 (N_4531,N_4331,N_4167);
nor U4532 (N_4532,N_4377,N_4086);
nor U4533 (N_4533,N_4393,N_4030);
or U4534 (N_4534,N_4026,N_4211);
or U4535 (N_4535,N_4272,N_4179);
nand U4536 (N_4536,N_4436,N_4487);
or U4537 (N_4537,N_4380,N_4231);
nor U4538 (N_4538,N_4310,N_4148);
nand U4539 (N_4539,N_4081,N_4077);
nand U4540 (N_4540,N_4144,N_4326);
xor U4541 (N_4541,N_4413,N_4332);
nand U4542 (N_4542,N_4375,N_4353);
nor U4543 (N_4543,N_4218,N_4068);
nand U4544 (N_4544,N_4150,N_4472);
xor U4545 (N_4545,N_4107,N_4307);
nand U4546 (N_4546,N_4232,N_4469);
nor U4547 (N_4547,N_4437,N_4215);
nand U4548 (N_4548,N_4240,N_4140);
nor U4549 (N_4549,N_4257,N_4370);
and U4550 (N_4550,N_4204,N_4359);
xor U4551 (N_4551,N_4005,N_4062);
nand U4552 (N_4552,N_4020,N_4462);
nor U4553 (N_4553,N_4089,N_4406);
and U4554 (N_4554,N_4401,N_4299);
nor U4555 (N_4555,N_4302,N_4087);
nor U4556 (N_4556,N_4327,N_4329);
or U4557 (N_4557,N_4494,N_4361);
nand U4558 (N_4558,N_4263,N_4160);
xnor U4559 (N_4559,N_4058,N_4279);
nor U4560 (N_4560,N_4190,N_4194);
nor U4561 (N_4561,N_4425,N_4482);
and U4562 (N_4562,N_4287,N_4133);
or U4563 (N_4563,N_4364,N_4239);
and U4564 (N_4564,N_4398,N_4197);
nand U4565 (N_4565,N_4216,N_4149);
nor U4566 (N_4566,N_4467,N_4082);
nand U4567 (N_4567,N_4410,N_4092);
and U4568 (N_4568,N_4415,N_4230);
or U4569 (N_4569,N_4024,N_4112);
or U4570 (N_4570,N_4036,N_4013);
xnor U4571 (N_4571,N_4276,N_4188);
nor U4572 (N_4572,N_4391,N_4200);
xnor U4573 (N_4573,N_4032,N_4228);
xor U4574 (N_4574,N_4348,N_4165);
nand U4575 (N_4575,N_4176,N_4374);
or U4576 (N_4576,N_4470,N_4076);
and U4577 (N_4577,N_4392,N_4121);
nand U4578 (N_4578,N_4171,N_4155);
nand U4579 (N_4579,N_4489,N_4021);
xnor U4580 (N_4580,N_4111,N_4440);
or U4581 (N_4581,N_4252,N_4074);
or U4582 (N_4582,N_4124,N_4277);
nand U4583 (N_4583,N_4224,N_4382);
xor U4584 (N_4584,N_4497,N_4412);
and U4585 (N_4585,N_4429,N_4403);
or U4586 (N_4586,N_4066,N_4039);
nand U4587 (N_4587,N_4321,N_4262);
nand U4588 (N_4588,N_4091,N_4110);
nor U4589 (N_4589,N_4452,N_4009);
or U4590 (N_4590,N_4481,N_4322);
nand U4591 (N_4591,N_4266,N_4126);
and U4592 (N_4592,N_4022,N_4098);
xnor U4593 (N_4593,N_4465,N_4294);
nand U4594 (N_4594,N_4152,N_4147);
nand U4595 (N_4595,N_4135,N_4373);
and U4596 (N_4596,N_4023,N_4293);
and U4597 (N_4597,N_4453,N_4309);
or U4598 (N_4598,N_4113,N_4356);
or U4599 (N_4599,N_4456,N_4109);
nand U4600 (N_4600,N_4379,N_4255);
and U4601 (N_4601,N_4043,N_4350);
or U4602 (N_4602,N_4234,N_4435);
or U4603 (N_4603,N_4308,N_4442);
nand U4604 (N_4604,N_4344,N_4123);
and U4605 (N_4605,N_4000,N_4284);
and U4606 (N_4606,N_4296,N_4464);
xor U4607 (N_4607,N_4245,N_4455);
nor U4608 (N_4608,N_4256,N_4396);
xnor U4609 (N_4609,N_4431,N_4400);
or U4610 (N_4610,N_4288,N_4432);
nand U4611 (N_4611,N_4151,N_4241);
nand U4612 (N_4612,N_4217,N_4101);
or U4613 (N_4613,N_4227,N_4193);
nor U4614 (N_4614,N_4118,N_4164);
nand U4615 (N_4615,N_4461,N_4096);
nor U4616 (N_4616,N_4486,N_4315);
and U4617 (N_4617,N_4106,N_4019);
nand U4618 (N_4618,N_4029,N_4278);
nor U4619 (N_4619,N_4229,N_4251);
and U4620 (N_4620,N_4214,N_4285);
or U4621 (N_4621,N_4367,N_4341);
or U4622 (N_4622,N_4064,N_4430);
nor U4623 (N_4623,N_4421,N_4045);
nor U4624 (N_4624,N_4340,N_4170);
nand U4625 (N_4625,N_4207,N_4225);
or U4626 (N_4626,N_4328,N_4182);
or U4627 (N_4627,N_4354,N_4209);
and U4628 (N_4628,N_4304,N_4071);
nor U4629 (N_4629,N_4424,N_4002);
xor U4630 (N_4630,N_4420,N_4095);
and U4631 (N_4631,N_4423,N_4491);
nand U4632 (N_4632,N_4038,N_4208);
or U4633 (N_4633,N_4366,N_4417);
nand U4634 (N_4634,N_4386,N_4466);
nand U4635 (N_4635,N_4189,N_4254);
nand U4636 (N_4636,N_4345,N_4488);
and U4637 (N_4637,N_4363,N_4157);
xnor U4638 (N_4638,N_4319,N_4282);
nor U4639 (N_4639,N_4090,N_4159);
nor U4640 (N_4640,N_4409,N_4053);
xor U4641 (N_4641,N_4443,N_4173);
and U4642 (N_4642,N_4492,N_4362);
or U4643 (N_4643,N_4444,N_4185);
nand U4644 (N_4644,N_4388,N_4237);
xor U4645 (N_4645,N_4168,N_4048);
nand U4646 (N_4646,N_4125,N_4291);
xnor U4647 (N_4647,N_4450,N_4324);
xor U4648 (N_4648,N_4408,N_4273);
and U4649 (N_4649,N_4463,N_4342);
or U4650 (N_4650,N_4389,N_4191);
nand U4651 (N_4651,N_4479,N_4313);
and U4652 (N_4652,N_4259,N_4192);
and U4653 (N_4653,N_4346,N_4014);
nor U4654 (N_4654,N_4075,N_4360);
and U4655 (N_4655,N_4057,N_4290);
nor U4656 (N_4656,N_4221,N_4268);
xor U4657 (N_4657,N_4059,N_4283);
and U4658 (N_4658,N_4033,N_4447);
and U4659 (N_4659,N_4264,N_4368);
xor U4660 (N_4660,N_4478,N_4166);
or U4661 (N_4661,N_4369,N_4198);
nand U4662 (N_4662,N_4117,N_4246);
nand U4663 (N_4663,N_4343,N_4365);
nand U4664 (N_4664,N_4203,N_4010);
nor U4665 (N_4665,N_4314,N_4422);
nand U4666 (N_4666,N_4376,N_4267);
or U4667 (N_4667,N_4247,N_4434);
nand U4668 (N_4668,N_4325,N_4445);
nand U4669 (N_4669,N_4142,N_4054);
and U4670 (N_4670,N_4303,N_4473);
and U4671 (N_4671,N_4060,N_4122);
xor U4672 (N_4672,N_4281,N_4017);
xor U4673 (N_4673,N_4130,N_4115);
and U4674 (N_4674,N_4298,N_4330);
or U4675 (N_4675,N_4046,N_4015);
and U4676 (N_4676,N_4079,N_4301);
nand U4677 (N_4677,N_4085,N_4381);
or U4678 (N_4678,N_4187,N_4212);
and U4679 (N_4679,N_4352,N_4274);
or U4680 (N_4680,N_4116,N_4312);
nand U4681 (N_4681,N_4286,N_4485);
or U4682 (N_4682,N_4051,N_4037);
nor U4683 (N_4683,N_4163,N_4196);
and U4684 (N_4684,N_4333,N_4186);
and U4685 (N_4685,N_4483,N_4136);
nor U4686 (N_4686,N_4336,N_4297);
nor U4687 (N_4687,N_4011,N_4270);
or U4688 (N_4688,N_4099,N_4154);
xor U4689 (N_4689,N_4161,N_4100);
xnor U4690 (N_4690,N_4258,N_4223);
nor U4691 (N_4691,N_4260,N_4405);
xor U4692 (N_4692,N_4496,N_4047);
and U4693 (N_4693,N_4351,N_4175);
xor U4694 (N_4694,N_4056,N_4414);
xor U4695 (N_4695,N_4271,N_4004);
and U4696 (N_4696,N_4138,N_4253);
and U4697 (N_4697,N_4428,N_4338);
or U4698 (N_4698,N_4055,N_4202);
nor U4699 (N_4699,N_4003,N_4495);
and U4700 (N_4700,N_4384,N_4335);
and U4701 (N_4701,N_4311,N_4153);
or U4702 (N_4702,N_4156,N_4143);
and U4703 (N_4703,N_4480,N_4069);
or U4704 (N_4704,N_4184,N_4265);
nor U4705 (N_4705,N_4390,N_4088);
or U4706 (N_4706,N_4222,N_4093);
nor U4707 (N_4707,N_4134,N_4399);
nand U4708 (N_4708,N_4459,N_4451);
and U4709 (N_4709,N_4248,N_4083);
xnor U4710 (N_4710,N_4181,N_4180);
or U4711 (N_4711,N_4394,N_4061);
nand U4712 (N_4712,N_4008,N_4484);
xnor U4713 (N_4713,N_4490,N_4404);
and U4714 (N_4714,N_4213,N_4041);
nand U4715 (N_4715,N_4269,N_4387);
nand U4716 (N_4716,N_4418,N_4025);
nand U4717 (N_4717,N_4105,N_4097);
nor U4718 (N_4718,N_4220,N_4102);
or U4719 (N_4719,N_4040,N_4242);
xnor U4720 (N_4720,N_4244,N_4471);
nand U4721 (N_4721,N_4233,N_4070);
or U4722 (N_4722,N_4139,N_4292);
or U4723 (N_4723,N_4468,N_4249);
or U4724 (N_4724,N_4407,N_4114);
xnor U4725 (N_4725,N_4323,N_4383);
xor U4726 (N_4726,N_4120,N_4243);
nor U4727 (N_4727,N_4049,N_4044);
and U4728 (N_4728,N_4063,N_4349);
nor U4729 (N_4729,N_4199,N_4067);
nor U4730 (N_4730,N_4104,N_4084);
and U4731 (N_4731,N_4385,N_4378);
nor U4732 (N_4732,N_4072,N_4416);
or U4733 (N_4733,N_4460,N_4275);
nor U4734 (N_4734,N_4042,N_4080);
xnor U4735 (N_4735,N_4300,N_4448);
or U4736 (N_4736,N_4206,N_4119);
or U4737 (N_4737,N_4103,N_4132);
xor U4738 (N_4738,N_4129,N_4295);
or U4739 (N_4739,N_4305,N_4028);
nor U4740 (N_4740,N_4065,N_4397);
and U4741 (N_4741,N_4320,N_4158);
nand U4742 (N_4742,N_4238,N_4261);
nor U4743 (N_4743,N_4052,N_4347);
nand U4744 (N_4744,N_4395,N_4306);
nor U4745 (N_4745,N_4339,N_4355);
and U4746 (N_4746,N_4219,N_4205);
xor U4747 (N_4747,N_4035,N_4337);
nor U4748 (N_4748,N_4449,N_4316);
and U4749 (N_4749,N_4476,N_4073);
nand U4750 (N_4750,N_4287,N_4168);
nand U4751 (N_4751,N_4211,N_4152);
and U4752 (N_4752,N_4335,N_4454);
xnor U4753 (N_4753,N_4432,N_4453);
xnor U4754 (N_4754,N_4151,N_4439);
and U4755 (N_4755,N_4052,N_4172);
nand U4756 (N_4756,N_4061,N_4283);
and U4757 (N_4757,N_4001,N_4250);
nand U4758 (N_4758,N_4210,N_4020);
or U4759 (N_4759,N_4376,N_4335);
nor U4760 (N_4760,N_4148,N_4023);
or U4761 (N_4761,N_4329,N_4446);
and U4762 (N_4762,N_4077,N_4416);
nand U4763 (N_4763,N_4282,N_4234);
xor U4764 (N_4764,N_4369,N_4291);
or U4765 (N_4765,N_4304,N_4281);
nand U4766 (N_4766,N_4231,N_4324);
nor U4767 (N_4767,N_4074,N_4432);
or U4768 (N_4768,N_4169,N_4441);
and U4769 (N_4769,N_4331,N_4087);
xnor U4770 (N_4770,N_4455,N_4217);
xor U4771 (N_4771,N_4299,N_4429);
or U4772 (N_4772,N_4282,N_4217);
and U4773 (N_4773,N_4274,N_4231);
and U4774 (N_4774,N_4482,N_4088);
and U4775 (N_4775,N_4312,N_4314);
nand U4776 (N_4776,N_4177,N_4286);
nand U4777 (N_4777,N_4094,N_4209);
nand U4778 (N_4778,N_4060,N_4081);
nand U4779 (N_4779,N_4208,N_4002);
and U4780 (N_4780,N_4456,N_4135);
nor U4781 (N_4781,N_4070,N_4410);
nand U4782 (N_4782,N_4253,N_4407);
and U4783 (N_4783,N_4455,N_4025);
nand U4784 (N_4784,N_4469,N_4353);
xnor U4785 (N_4785,N_4435,N_4412);
nand U4786 (N_4786,N_4476,N_4394);
nand U4787 (N_4787,N_4494,N_4078);
nand U4788 (N_4788,N_4443,N_4480);
or U4789 (N_4789,N_4106,N_4371);
nand U4790 (N_4790,N_4064,N_4289);
xor U4791 (N_4791,N_4229,N_4226);
nand U4792 (N_4792,N_4347,N_4209);
xnor U4793 (N_4793,N_4189,N_4203);
nor U4794 (N_4794,N_4443,N_4316);
nor U4795 (N_4795,N_4133,N_4052);
nand U4796 (N_4796,N_4480,N_4285);
xor U4797 (N_4797,N_4418,N_4448);
and U4798 (N_4798,N_4082,N_4198);
xnor U4799 (N_4799,N_4317,N_4096);
nor U4800 (N_4800,N_4190,N_4007);
xnor U4801 (N_4801,N_4164,N_4314);
or U4802 (N_4802,N_4220,N_4318);
or U4803 (N_4803,N_4376,N_4427);
or U4804 (N_4804,N_4297,N_4173);
nor U4805 (N_4805,N_4282,N_4406);
and U4806 (N_4806,N_4013,N_4071);
nor U4807 (N_4807,N_4300,N_4071);
nor U4808 (N_4808,N_4452,N_4296);
and U4809 (N_4809,N_4316,N_4057);
nor U4810 (N_4810,N_4157,N_4103);
xor U4811 (N_4811,N_4171,N_4497);
nand U4812 (N_4812,N_4443,N_4252);
nor U4813 (N_4813,N_4148,N_4421);
nand U4814 (N_4814,N_4054,N_4304);
or U4815 (N_4815,N_4478,N_4304);
or U4816 (N_4816,N_4208,N_4270);
and U4817 (N_4817,N_4122,N_4446);
and U4818 (N_4818,N_4354,N_4125);
and U4819 (N_4819,N_4059,N_4090);
xnor U4820 (N_4820,N_4235,N_4448);
nor U4821 (N_4821,N_4217,N_4437);
xor U4822 (N_4822,N_4460,N_4403);
or U4823 (N_4823,N_4056,N_4238);
or U4824 (N_4824,N_4075,N_4298);
nand U4825 (N_4825,N_4059,N_4176);
nand U4826 (N_4826,N_4001,N_4346);
xor U4827 (N_4827,N_4059,N_4378);
nand U4828 (N_4828,N_4356,N_4242);
or U4829 (N_4829,N_4402,N_4455);
xnor U4830 (N_4830,N_4162,N_4122);
nand U4831 (N_4831,N_4441,N_4254);
and U4832 (N_4832,N_4162,N_4412);
nor U4833 (N_4833,N_4207,N_4003);
nand U4834 (N_4834,N_4253,N_4469);
and U4835 (N_4835,N_4298,N_4031);
nand U4836 (N_4836,N_4186,N_4052);
xor U4837 (N_4837,N_4414,N_4141);
and U4838 (N_4838,N_4447,N_4156);
xnor U4839 (N_4839,N_4043,N_4149);
xor U4840 (N_4840,N_4140,N_4225);
and U4841 (N_4841,N_4154,N_4305);
or U4842 (N_4842,N_4309,N_4359);
nand U4843 (N_4843,N_4277,N_4439);
nor U4844 (N_4844,N_4231,N_4480);
or U4845 (N_4845,N_4029,N_4079);
or U4846 (N_4846,N_4229,N_4345);
nor U4847 (N_4847,N_4372,N_4136);
and U4848 (N_4848,N_4432,N_4068);
or U4849 (N_4849,N_4015,N_4300);
nand U4850 (N_4850,N_4231,N_4282);
or U4851 (N_4851,N_4351,N_4159);
xnor U4852 (N_4852,N_4032,N_4286);
or U4853 (N_4853,N_4284,N_4165);
nand U4854 (N_4854,N_4043,N_4048);
nor U4855 (N_4855,N_4486,N_4169);
or U4856 (N_4856,N_4478,N_4032);
and U4857 (N_4857,N_4421,N_4269);
or U4858 (N_4858,N_4017,N_4026);
or U4859 (N_4859,N_4031,N_4179);
nor U4860 (N_4860,N_4481,N_4412);
nand U4861 (N_4861,N_4324,N_4283);
nand U4862 (N_4862,N_4435,N_4269);
or U4863 (N_4863,N_4398,N_4239);
nand U4864 (N_4864,N_4263,N_4486);
and U4865 (N_4865,N_4097,N_4167);
and U4866 (N_4866,N_4494,N_4028);
or U4867 (N_4867,N_4423,N_4086);
xnor U4868 (N_4868,N_4269,N_4343);
or U4869 (N_4869,N_4189,N_4176);
nand U4870 (N_4870,N_4198,N_4124);
or U4871 (N_4871,N_4115,N_4081);
or U4872 (N_4872,N_4038,N_4266);
nor U4873 (N_4873,N_4357,N_4470);
nand U4874 (N_4874,N_4256,N_4089);
xor U4875 (N_4875,N_4094,N_4365);
and U4876 (N_4876,N_4494,N_4274);
nor U4877 (N_4877,N_4434,N_4041);
nand U4878 (N_4878,N_4003,N_4262);
xnor U4879 (N_4879,N_4441,N_4419);
or U4880 (N_4880,N_4303,N_4499);
xor U4881 (N_4881,N_4396,N_4155);
and U4882 (N_4882,N_4480,N_4197);
or U4883 (N_4883,N_4302,N_4055);
and U4884 (N_4884,N_4196,N_4377);
and U4885 (N_4885,N_4298,N_4025);
nor U4886 (N_4886,N_4472,N_4230);
xnor U4887 (N_4887,N_4237,N_4432);
xnor U4888 (N_4888,N_4139,N_4185);
and U4889 (N_4889,N_4347,N_4004);
nor U4890 (N_4890,N_4127,N_4494);
and U4891 (N_4891,N_4298,N_4390);
nor U4892 (N_4892,N_4413,N_4025);
or U4893 (N_4893,N_4239,N_4120);
and U4894 (N_4894,N_4110,N_4320);
or U4895 (N_4895,N_4250,N_4115);
and U4896 (N_4896,N_4475,N_4451);
xor U4897 (N_4897,N_4334,N_4320);
xnor U4898 (N_4898,N_4421,N_4216);
nor U4899 (N_4899,N_4338,N_4157);
or U4900 (N_4900,N_4389,N_4245);
nand U4901 (N_4901,N_4001,N_4124);
nor U4902 (N_4902,N_4473,N_4437);
nand U4903 (N_4903,N_4414,N_4263);
xor U4904 (N_4904,N_4483,N_4261);
nor U4905 (N_4905,N_4394,N_4480);
nand U4906 (N_4906,N_4197,N_4293);
and U4907 (N_4907,N_4134,N_4088);
nand U4908 (N_4908,N_4025,N_4319);
xor U4909 (N_4909,N_4076,N_4343);
nand U4910 (N_4910,N_4340,N_4412);
and U4911 (N_4911,N_4156,N_4384);
or U4912 (N_4912,N_4164,N_4463);
or U4913 (N_4913,N_4248,N_4379);
nand U4914 (N_4914,N_4240,N_4303);
nor U4915 (N_4915,N_4362,N_4143);
and U4916 (N_4916,N_4071,N_4313);
xnor U4917 (N_4917,N_4020,N_4323);
nor U4918 (N_4918,N_4008,N_4227);
xnor U4919 (N_4919,N_4328,N_4219);
nor U4920 (N_4920,N_4215,N_4429);
nand U4921 (N_4921,N_4256,N_4028);
nand U4922 (N_4922,N_4429,N_4130);
nor U4923 (N_4923,N_4204,N_4043);
nand U4924 (N_4924,N_4298,N_4160);
nor U4925 (N_4925,N_4448,N_4055);
nor U4926 (N_4926,N_4171,N_4044);
nand U4927 (N_4927,N_4320,N_4472);
or U4928 (N_4928,N_4036,N_4260);
nand U4929 (N_4929,N_4008,N_4061);
or U4930 (N_4930,N_4185,N_4227);
nand U4931 (N_4931,N_4253,N_4097);
xor U4932 (N_4932,N_4032,N_4071);
and U4933 (N_4933,N_4123,N_4093);
or U4934 (N_4934,N_4192,N_4153);
nand U4935 (N_4935,N_4040,N_4443);
nor U4936 (N_4936,N_4105,N_4351);
or U4937 (N_4937,N_4124,N_4190);
and U4938 (N_4938,N_4036,N_4157);
nor U4939 (N_4939,N_4241,N_4314);
nand U4940 (N_4940,N_4436,N_4086);
xnor U4941 (N_4941,N_4443,N_4030);
and U4942 (N_4942,N_4074,N_4442);
nor U4943 (N_4943,N_4082,N_4234);
nor U4944 (N_4944,N_4041,N_4407);
or U4945 (N_4945,N_4083,N_4272);
or U4946 (N_4946,N_4266,N_4005);
nand U4947 (N_4947,N_4496,N_4144);
or U4948 (N_4948,N_4253,N_4312);
nand U4949 (N_4949,N_4476,N_4039);
and U4950 (N_4950,N_4326,N_4317);
xnor U4951 (N_4951,N_4352,N_4205);
and U4952 (N_4952,N_4088,N_4425);
nand U4953 (N_4953,N_4437,N_4180);
or U4954 (N_4954,N_4100,N_4021);
nor U4955 (N_4955,N_4245,N_4361);
nand U4956 (N_4956,N_4200,N_4212);
and U4957 (N_4957,N_4414,N_4304);
nand U4958 (N_4958,N_4020,N_4431);
xnor U4959 (N_4959,N_4218,N_4289);
nand U4960 (N_4960,N_4420,N_4497);
or U4961 (N_4961,N_4052,N_4005);
or U4962 (N_4962,N_4213,N_4218);
and U4963 (N_4963,N_4164,N_4101);
xor U4964 (N_4964,N_4308,N_4009);
xnor U4965 (N_4965,N_4230,N_4120);
and U4966 (N_4966,N_4347,N_4020);
xnor U4967 (N_4967,N_4472,N_4170);
or U4968 (N_4968,N_4339,N_4253);
xor U4969 (N_4969,N_4171,N_4097);
nor U4970 (N_4970,N_4124,N_4257);
or U4971 (N_4971,N_4258,N_4410);
and U4972 (N_4972,N_4014,N_4432);
nand U4973 (N_4973,N_4147,N_4348);
and U4974 (N_4974,N_4082,N_4029);
or U4975 (N_4975,N_4218,N_4150);
nand U4976 (N_4976,N_4163,N_4245);
nand U4977 (N_4977,N_4486,N_4165);
and U4978 (N_4978,N_4116,N_4019);
nor U4979 (N_4979,N_4043,N_4482);
and U4980 (N_4980,N_4187,N_4317);
and U4981 (N_4981,N_4343,N_4138);
or U4982 (N_4982,N_4442,N_4468);
and U4983 (N_4983,N_4152,N_4186);
or U4984 (N_4984,N_4384,N_4073);
xor U4985 (N_4985,N_4240,N_4067);
nand U4986 (N_4986,N_4437,N_4135);
and U4987 (N_4987,N_4403,N_4204);
nor U4988 (N_4988,N_4324,N_4078);
and U4989 (N_4989,N_4161,N_4399);
nand U4990 (N_4990,N_4468,N_4048);
nand U4991 (N_4991,N_4298,N_4180);
or U4992 (N_4992,N_4280,N_4043);
nor U4993 (N_4993,N_4135,N_4342);
and U4994 (N_4994,N_4038,N_4456);
or U4995 (N_4995,N_4171,N_4328);
or U4996 (N_4996,N_4383,N_4188);
nor U4997 (N_4997,N_4473,N_4194);
or U4998 (N_4998,N_4125,N_4132);
nand U4999 (N_4999,N_4337,N_4211);
and UO_0 (O_0,N_4766,N_4623);
and UO_1 (O_1,N_4721,N_4890);
nand UO_2 (O_2,N_4981,N_4765);
nor UO_3 (O_3,N_4661,N_4996);
or UO_4 (O_4,N_4643,N_4936);
or UO_5 (O_5,N_4690,N_4512);
and UO_6 (O_6,N_4944,N_4923);
and UO_7 (O_7,N_4859,N_4926);
nand UO_8 (O_8,N_4559,N_4578);
or UO_9 (O_9,N_4642,N_4939);
xnor UO_10 (O_10,N_4851,N_4845);
and UO_11 (O_11,N_4969,N_4551);
or UO_12 (O_12,N_4806,N_4786);
and UO_13 (O_13,N_4664,N_4889);
nand UO_14 (O_14,N_4897,N_4532);
or UO_15 (O_15,N_4997,N_4908);
xor UO_16 (O_16,N_4764,N_4612);
or UO_17 (O_17,N_4634,N_4757);
and UO_18 (O_18,N_4542,N_4910);
nor UO_19 (O_19,N_4956,N_4695);
and UO_20 (O_20,N_4892,N_4724);
xnor UO_21 (O_21,N_4694,N_4844);
nand UO_22 (O_22,N_4941,N_4976);
and UO_23 (O_23,N_4625,N_4887);
xor UO_24 (O_24,N_4907,N_4547);
and UO_25 (O_25,N_4648,N_4616);
and UO_26 (O_26,N_4769,N_4790);
and UO_27 (O_27,N_4539,N_4654);
xnor UO_28 (O_28,N_4633,N_4574);
nor UO_29 (O_29,N_4853,N_4776);
or UO_30 (O_30,N_4651,N_4788);
or UO_31 (O_31,N_4602,N_4508);
nand UO_32 (O_32,N_4506,N_4793);
or UO_33 (O_33,N_4550,N_4727);
and UO_34 (O_34,N_4999,N_4658);
nand UO_35 (O_35,N_4868,N_4697);
or UO_36 (O_36,N_4819,N_4528);
and UO_37 (O_37,N_4515,N_4884);
nor UO_38 (O_38,N_4977,N_4659);
nor UO_39 (O_39,N_4967,N_4987);
or UO_40 (O_40,N_4590,N_4605);
nor UO_41 (O_41,N_4781,N_4621);
nor UO_42 (O_42,N_4774,N_4826);
xor UO_43 (O_43,N_4900,N_4915);
or UO_44 (O_44,N_4829,N_4677);
nor UO_45 (O_45,N_4922,N_4873);
xor UO_46 (O_46,N_4912,N_4921);
nand UO_47 (O_47,N_4901,N_4975);
xnor UO_48 (O_48,N_4741,N_4593);
nand UO_49 (O_49,N_4720,N_4875);
nor UO_50 (O_50,N_4777,N_4636);
xnor UO_51 (O_51,N_4840,N_4945);
or UO_52 (O_52,N_4647,N_4738);
xor UO_53 (O_53,N_4750,N_4834);
and UO_54 (O_54,N_4606,N_4656);
and UO_55 (O_55,N_4570,N_4848);
and UO_56 (O_56,N_4548,N_4713);
and UO_57 (O_57,N_4615,N_4723);
or UO_58 (O_58,N_4828,N_4671);
xnor UO_59 (O_59,N_4913,N_4965);
nor UO_60 (O_60,N_4689,N_4505);
and UO_61 (O_61,N_4595,N_4983);
nor UO_62 (O_62,N_4718,N_4755);
nor UO_63 (O_63,N_4526,N_4904);
nand UO_64 (O_64,N_4843,N_4905);
nand UO_65 (O_65,N_4816,N_4730);
or UO_66 (O_66,N_4674,N_4745);
nor UO_67 (O_67,N_4847,N_4811);
nor UO_68 (O_68,N_4799,N_4955);
nor UO_69 (O_69,N_4672,N_4796);
or UO_70 (O_70,N_4657,N_4563);
xor UO_71 (O_71,N_4998,N_4837);
or UO_72 (O_72,N_4771,N_4763);
nand UO_73 (O_73,N_4702,N_4872);
nor UO_74 (O_74,N_4637,N_4917);
nand UO_75 (O_75,N_4778,N_4669);
and UO_76 (O_76,N_4557,N_4952);
and UO_77 (O_77,N_4833,N_4920);
xor UO_78 (O_78,N_4985,N_4747);
and UO_79 (O_79,N_4968,N_4589);
xnor UO_80 (O_80,N_4814,N_4725);
and UO_81 (O_81,N_4712,N_4553);
xnor UO_82 (O_82,N_4504,N_4959);
or UO_83 (O_83,N_4673,N_4680);
nand UO_84 (O_84,N_4536,N_4620);
nor UO_85 (O_85,N_4575,N_4916);
xor UO_86 (O_86,N_4783,N_4644);
and UO_87 (O_87,N_4839,N_4537);
or UO_88 (O_88,N_4626,N_4773);
xor UO_89 (O_89,N_4744,N_4991);
nor UO_90 (O_90,N_4514,N_4767);
nor UO_91 (O_91,N_4742,N_4632);
nand UO_92 (O_92,N_4792,N_4770);
xnor UO_93 (O_93,N_4813,N_4984);
nor UO_94 (O_94,N_4762,N_4972);
nand UO_95 (O_95,N_4911,N_4645);
nor UO_96 (O_96,N_4963,N_4544);
or UO_97 (O_97,N_4604,N_4679);
and UO_98 (O_98,N_4638,N_4520);
nand UO_99 (O_99,N_4925,N_4879);
or UO_100 (O_100,N_4617,N_4601);
and UO_101 (O_101,N_4698,N_4650);
xnor UO_102 (O_102,N_4599,N_4940);
or UO_103 (O_103,N_4893,N_4619);
xor UO_104 (O_104,N_4979,N_4622);
nand UO_105 (O_105,N_4501,N_4989);
xor UO_106 (O_106,N_4701,N_4753);
and UO_107 (O_107,N_4865,N_4596);
nand UO_108 (O_108,N_4871,N_4681);
and UO_109 (O_109,N_4630,N_4877);
xnor UO_110 (O_110,N_4800,N_4540);
nor UO_111 (O_111,N_4885,N_4947);
xor UO_112 (O_112,N_4715,N_4739);
nor UO_113 (O_113,N_4899,N_4541);
nand UO_114 (O_114,N_4565,N_4519);
or UO_115 (O_115,N_4988,N_4958);
and UO_116 (O_116,N_4962,N_4954);
and UO_117 (O_117,N_4631,N_4585);
and UO_118 (O_118,N_4618,N_4719);
nand UO_119 (O_119,N_4861,N_4543);
xor UO_120 (O_120,N_4749,N_4835);
nand UO_121 (O_121,N_4676,N_4867);
or UO_122 (O_122,N_4614,N_4737);
or UO_123 (O_123,N_4662,N_4818);
or UO_124 (O_124,N_4572,N_4948);
or UO_125 (O_125,N_4576,N_4990);
xnor UO_126 (O_126,N_4896,N_4588);
xnor UO_127 (O_127,N_4928,N_4971);
and UO_128 (O_128,N_4707,N_4660);
xor UO_129 (O_129,N_4743,N_4809);
nor UO_130 (O_130,N_4726,N_4561);
nor UO_131 (O_131,N_4521,N_4552);
nand UO_132 (O_132,N_4937,N_4670);
and UO_133 (O_133,N_4728,N_4652);
xnor UO_134 (O_134,N_4586,N_4663);
nand UO_135 (O_135,N_4748,N_4527);
xnor UO_136 (O_136,N_4869,N_4761);
or UO_137 (O_137,N_4609,N_4863);
or UO_138 (O_138,N_4525,N_4775);
xor UO_139 (O_139,N_4556,N_4667);
nand UO_140 (O_140,N_4927,N_4569);
nor UO_141 (O_141,N_4759,N_4898);
and UO_142 (O_142,N_4850,N_4894);
or UO_143 (O_143,N_4949,N_4534);
or UO_144 (O_144,N_4655,N_4597);
or UO_145 (O_145,N_4895,N_4964);
nor UO_146 (O_146,N_4772,N_4583);
and UO_147 (O_147,N_4627,N_4874);
or UO_148 (O_148,N_4524,N_4780);
xor UO_149 (O_149,N_4810,N_4919);
nor UO_150 (O_150,N_4629,N_4584);
nor UO_151 (O_151,N_4691,N_4932);
xnor UO_152 (O_152,N_4852,N_4994);
nand UO_153 (O_153,N_4831,N_4500);
xor UO_154 (O_154,N_4902,N_4815);
and UO_155 (O_155,N_4704,N_4933);
and UO_156 (O_156,N_4533,N_4705);
xnor UO_157 (O_157,N_4685,N_4560);
nand UO_158 (O_158,N_4870,N_4717);
nand UO_159 (O_159,N_4931,N_4581);
xnor UO_160 (O_160,N_4752,N_4960);
xnor UO_161 (O_161,N_4607,N_4817);
nand UO_162 (O_162,N_4836,N_4830);
and UO_163 (O_163,N_4562,N_4503);
nor UO_164 (O_164,N_4883,N_4710);
nor UO_165 (O_165,N_4608,N_4930);
or UO_166 (O_166,N_4974,N_4567);
or UO_167 (O_167,N_4687,N_4878);
or UO_168 (O_168,N_4522,N_4866);
nand UO_169 (O_169,N_4880,N_4882);
nor UO_170 (O_170,N_4758,N_4760);
nand UO_171 (O_171,N_4555,N_4846);
or UO_172 (O_172,N_4918,N_4973);
or UO_173 (O_173,N_4914,N_4785);
and UO_174 (O_174,N_4838,N_4798);
xnor UO_175 (O_175,N_4754,N_4807);
or UO_176 (O_176,N_4906,N_4805);
nand UO_177 (O_177,N_4832,N_4736);
and UO_178 (O_178,N_4703,N_4888);
nor UO_179 (O_179,N_4782,N_4688);
and UO_180 (O_180,N_4641,N_4531);
xnor UO_181 (O_181,N_4943,N_4876);
xor UO_182 (O_182,N_4862,N_4823);
and UO_183 (O_183,N_4518,N_4678);
nand UO_184 (O_184,N_4535,N_4530);
xnor UO_185 (O_185,N_4995,N_4509);
and UO_186 (O_186,N_4993,N_4957);
xor UO_187 (O_187,N_4558,N_4624);
xor UO_188 (O_188,N_4803,N_4529);
xnor UO_189 (O_189,N_4756,N_4966);
or UO_190 (O_190,N_4784,N_4566);
nand UO_191 (O_191,N_4942,N_4804);
or UO_192 (O_192,N_4857,N_4709);
and UO_193 (O_193,N_4716,N_4545);
or UO_194 (O_194,N_4986,N_4582);
nor UO_195 (O_195,N_4711,N_4683);
and UO_196 (O_196,N_4841,N_4502);
or UO_197 (O_197,N_4881,N_4646);
and UO_198 (O_198,N_4822,N_4682);
nor UO_199 (O_199,N_4577,N_4587);
and UO_200 (O_200,N_4980,N_4953);
and UO_201 (O_201,N_4668,N_4794);
or UO_202 (O_202,N_4801,N_4549);
nor UO_203 (O_203,N_4978,N_4789);
nor UO_204 (O_204,N_4538,N_4600);
xnor UO_205 (O_205,N_4787,N_4860);
and UO_206 (O_206,N_4797,N_4523);
nand UO_207 (O_207,N_4666,N_4729);
and UO_208 (O_208,N_4935,N_4579);
nor UO_209 (O_209,N_4517,N_4946);
nand UO_210 (O_210,N_4573,N_4929);
xnor UO_211 (O_211,N_4675,N_4849);
or UO_212 (O_212,N_4706,N_4610);
or UO_213 (O_213,N_4722,N_4580);
nand UO_214 (O_214,N_4568,N_4795);
nand UO_215 (O_215,N_4516,N_4603);
nor UO_216 (O_216,N_4571,N_4733);
xor UO_217 (O_217,N_4686,N_4891);
or UO_218 (O_218,N_4909,N_4858);
xor UO_219 (O_219,N_4700,N_4938);
nand UO_220 (O_220,N_4842,N_4692);
nor UO_221 (O_221,N_4653,N_4903);
and UO_222 (O_222,N_4820,N_4827);
or UO_223 (O_223,N_4513,N_4649);
or UO_224 (O_224,N_4684,N_4714);
or UO_225 (O_225,N_4731,N_4951);
nand UO_226 (O_226,N_4825,N_4591);
or UO_227 (O_227,N_4854,N_4779);
nand UO_228 (O_228,N_4734,N_4992);
nor UO_229 (O_229,N_4768,N_4511);
or UO_230 (O_230,N_4934,N_4924);
nand UO_231 (O_231,N_4802,N_4635);
or UO_232 (O_232,N_4639,N_4732);
xor UO_233 (O_233,N_4640,N_4665);
xor UO_234 (O_234,N_4824,N_4982);
nor UO_235 (O_235,N_4864,N_4546);
nor UO_236 (O_236,N_4696,N_4510);
nand UO_237 (O_237,N_4821,N_4611);
nand UO_238 (O_238,N_4886,N_4751);
nand UO_239 (O_239,N_4592,N_4746);
nand UO_240 (O_240,N_4708,N_4961);
nand UO_241 (O_241,N_4808,N_4856);
nor UO_242 (O_242,N_4970,N_4598);
or UO_243 (O_243,N_4554,N_4812);
or UO_244 (O_244,N_4735,N_4507);
and UO_245 (O_245,N_4855,N_4693);
and UO_246 (O_246,N_4564,N_4791);
or UO_247 (O_247,N_4740,N_4628);
nor UO_248 (O_248,N_4950,N_4594);
nor UO_249 (O_249,N_4699,N_4613);
xnor UO_250 (O_250,N_4661,N_4903);
and UO_251 (O_251,N_4980,N_4568);
nor UO_252 (O_252,N_4730,N_4970);
nor UO_253 (O_253,N_4975,N_4508);
xnor UO_254 (O_254,N_4929,N_4617);
xnor UO_255 (O_255,N_4989,N_4518);
and UO_256 (O_256,N_4904,N_4941);
and UO_257 (O_257,N_4784,N_4830);
nand UO_258 (O_258,N_4698,N_4908);
xor UO_259 (O_259,N_4989,N_4799);
nand UO_260 (O_260,N_4967,N_4639);
or UO_261 (O_261,N_4892,N_4804);
nor UO_262 (O_262,N_4698,N_4822);
nor UO_263 (O_263,N_4959,N_4647);
nand UO_264 (O_264,N_4500,N_4774);
nand UO_265 (O_265,N_4812,N_4908);
xnor UO_266 (O_266,N_4945,N_4806);
or UO_267 (O_267,N_4588,N_4586);
and UO_268 (O_268,N_4947,N_4710);
or UO_269 (O_269,N_4581,N_4599);
and UO_270 (O_270,N_4664,N_4882);
xnor UO_271 (O_271,N_4871,N_4928);
nand UO_272 (O_272,N_4902,N_4659);
nand UO_273 (O_273,N_4572,N_4533);
nor UO_274 (O_274,N_4581,N_4831);
nor UO_275 (O_275,N_4933,N_4565);
nor UO_276 (O_276,N_4733,N_4613);
nand UO_277 (O_277,N_4561,N_4940);
xnor UO_278 (O_278,N_4607,N_4914);
or UO_279 (O_279,N_4850,N_4769);
and UO_280 (O_280,N_4859,N_4692);
and UO_281 (O_281,N_4635,N_4733);
or UO_282 (O_282,N_4751,N_4827);
nor UO_283 (O_283,N_4828,N_4921);
nand UO_284 (O_284,N_4841,N_4892);
or UO_285 (O_285,N_4535,N_4572);
xnor UO_286 (O_286,N_4527,N_4861);
nand UO_287 (O_287,N_4793,N_4699);
and UO_288 (O_288,N_4942,N_4934);
or UO_289 (O_289,N_4532,N_4961);
nand UO_290 (O_290,N_4650,N_4992);
nand UO_291 (O_291,N_4963,N_4964);
and UO_292 (O_292,N_4884,N_4932);
nand UO_293 (O_293,N_4601,N_4814);
xor UO_294 (O_294,N_4587,N_4726);
or UO_295 (O_295,N_4691,N_4875);
and UO_296 (O_296,N_4964,N_4609);
and UO_297 (O_297,N_4964,N_4588);
xor UO_298 (O_298,N_4976,N_4583);
nor UO_299 (O_299,N_4747,N_4745);
xnor UO_300 (O_300,N_4676,N_4527);
and UO_301 (O_301,N_4663,N_4501);
nand UO_302 (O_302,N_4680,N_4665);
nor UO_303 (O_303,N_4944,N_4883);
and UO_304 (O_304,N_4518,N_4696);
xor UO_305 (O_305,N_4921,N_4965);
and UO_306 (O_306,N_4518,N_4802);
xor UO_307 (O_307,N_4569,N_4834);
or UO_308 (O_308,N_4756,N_4534);
nand UO_309 (O_309,N_4828,N_4973);
and UO_310 (O_310,N_4547,N_4984);
xnor UO_311 (O_311,N_4674,N_4930);
and UO_312 (O_312,N_4542,N_4719);
or UO_313 (O_313,N_4593,N_4525);
xor UO_314 (O_314,N_4711,N_4627);
nand UO_315 (O_315,N_4607,N_4715);
and UO_316 (O_316,N_4965,N_4864);
nand UO_317 (O_317,N_4507,N_4827);
xor UO_318 (O_318,N_4806,N_4661);
nand UO_319 (O_319,N_4784,N_4735);
and UO_320 (O_320,N_4520,N_4682);
nor UO_321 (O_321,N_4981,N_4734);
xor UO_322 (O_322,N_4898,N_4624);
xor UO_323 (O_323,N_4588,N_4534);
or UO_324 (O_324,N_4893,N_4923);
nor UO_325 (O_325,N_4830,N_4822);
nor UO_326 (O_326,N_4984,N_4688);
or UO_327 (O_327,N_4784,N_4738);
and UO_328 (O_328,N_4815,N_4771);
nor UO_329 (O_329,N_4568,N_4949);
or UO_330 (O_330,N_4621,N_4994);
or UO_331 (O_331,N_4795,N_4893);
nor UO_332 (O_332,N_4757,N_4533);
nor UO_333 (O_333,N_4990,N_4726);
and UO_334 (O_334,N_4616,N_4714);
and UO_335 (O_335,N_4759,N_4809);
xor UO_336 (O_336,N_4892,N_4590);
xnor UO_337 (O_337,N_4664,N_4972);
or UO_338 (O_338,N_4684,N_4737);
xnor UO_339 (O_339,N_4729,N_4595);
xor UO_340 (O_340,N_4846,N_4718);
and UO_341 (O_341,N_4941,N_4532);
nor UO_342 (O_342,N_4993,N_4576);
nand UO_343 (O_343,N_4795,N_4727);
xor UO_344 (O_344,N_4669,N_4854);
and UO_345 (O_345,N_4782,N_4557);
and UO_346 (O_346,N_4890,N_4832);
xor UO_347 (O_347,N_4594,N_4882);
nor UO_348 (O_348,N_4619,N_4559);
and UO_349 (O_349,N_4675,N_4602);
xor UO_350 (O_350,N_4870,N_4725);
xnor UO_351 (O_351,N_4977,N_4883);
and UO_352 (O_352,N_4776,N_4680);
or UO_353 (O_353,N_4932,N_4559);
and UO_354 (O_354,N_4836,N_4851);
nand UO_355 (O_355,N_4807,N_4953);
nand UO_356 (O_356,N_4838,N_4839);
or UO_357 (O_357,N_4771,N_4830);
and UO_358 (O_358,N_4789,N_4838);
or UO_359 (O_359,N_4897,N_4602);
nor UO_360 (O_360,N_4566,N_4579);
xor UO_361 (O_361,N_4932,N_4721);
or UO_362 (O_362,N_4659,N_4688);
or UO_363 (O_363,N_4993,N_4921);
xnor UO_364 (O_364,N_4520,N_4781);
nand UO_365 (O_365,N_4704,N_4586);
and UO_366 (O_366,N_4887,N_4546);
nor UO_367 (O_367,N_4857,N_4559);
and UO_368 (O_368,N_4842,N_4807);
or UO_369 (O_369,N_4707,N_4573);
nand UO_370 (O_370,N_4768,N_4713);
nand UO_371 (O_371,N_4646,N_4854);
and UO_372 (O_372,N_4689,N_4889);
nand UO_373 (O_373,N_4856,N_4724);
nand UO_374 (O_374,N_4758,N_4647);
nor UO_375 (O_375,N_4560,N_4759);
nor UO_376 (O_376,N_4881,N_4844);
or UO_377 (O_377,N_4644,N_4651);
nor UO_378 (O_378,N_4511,N_4632);
and UO_379 (O_379,N_4871,N_4770);
nor UO_380 (O_380,N_4997,N_4859);
nor UO_381 (O_381,N_4535,N_4952);
and UO_382 (O_382,N_4781,N_4810);
and UO_383 (O_383,N_4789,N_4641);
nor UO_384 (O_384,N_4599,N_4509);
xnor UO_385 (O_385,N_4506,N_4803);
nand UO_386 (O_386,N_4670,N_4950);
nor UO_387 (O_387,N_4773,N_4511);
nor UO_388 (O_388,N_4913,N_4954);
or UO_389 (O_389,N_4690,N_4520);
nand UO_390 (O_390,N_4645,N_4634);
xor UO_391 (O_391,N_4963,N_4980);
and UO_392 (O_392,N_4874,N_4659);
nand UO_393 (O_393,N_4985,N_4780);
or UO_394 (O_394,N_4832,N_4642);
xnor UO_395 (O_395,N_4657,N_4698);
or UO_396 (O_396,N_4558,N_4676);
nand UO_397 (O_397,N_4869,N_4923);
or UO_398 (O_398,N_4943,N_4851);
and UO_399 (O_399,N_4894,N_4962);
nand UO_400 (O_400,N_4685,N_4865);
nand UO_401 (O_401,N_4599,N_4554);
xor UO_402 (O_402,N_4740,N_4508);
and UO_403 (O_403,N_4845,N_4584);
or UO_404 (O_404,N_4983,N_4553);
and UO_405 (O_405,N_4530,N_4701);
xnor UO_406 (O_406,N_4820,N_4886);
nor UO_407 (O_407,N_4898,N_4732);
nor UO_408 (O_408,N_4520,N_4820);
and UO_409 (O_409,N_4549,N_4631);
nor UO_410 (O_410,N_4824,N_4609);
or UO_411 (O_411,N_4710,N_4510);
nand UO_412 (O_412,N_4981,N_4674);
nand UO_413 (O_413,N_4959,N_4598);
xor UO_414 (O_414,N_4692,N_4620);
and UO_415 (O_415,N_4602,N_4708);
nor UO_416 (O_416,N_4735,N_4768);
xnor UO_417 (O_417,N_4903,N_4592);
xor UO_418 (O_418,N_4893,N_4657);
nand UO_419 (O_419,N_4732,N_4775);
nor UO_420 (O_420,N_4868,N_4949);
nor UO_421 (O_421,N_4624,N_4924);
or UO_422 (O_422,N_4767,N_4889);
xor UO_423 (O_423,N_4500,N_4572);
and UO_424 (O_424,N_4768,N_4822);
nand UO_425 (O_425,N_4919,N_4931);
or UO_426 (O_426,N_4938,N_4701);
or UO_427 (O_427,N_4629,N_4684);
nand UO_428 (O_428,N_4954,N_4563);
nand UO_429 (O_429,N_4673,N_4968);
or UO_430 (O_430,N_4617,N_4680);
xor UO_431 (O_431,N_4645,N_4879);
nand UO_432 (O_432,N_4652,N_4593);
or UO_433 (O_433,N_4506,N_4584);
or UO_434 (O_434,N_4947,N_4565);
xor UO_435 (O_435,N_4931,N_4681);
or UO_436 (O_436,N_4545,N_4886);
or UO_437 (O_437,N_4828,N_4978);
nand UO_438 (O_438,N_4582,N_4642);
and UO_439 (O_439,N_4754,N_4589);
nand UO_440 (O_440,N_4527,N_4654);
nor UO_441 (O_441,N_4563,N_4835);
nor UO_442 (O_442,N_4862,N_4795);
and UO_443 (O_443,N_4728,N_4903);
nor UO_444 (O_444,N_4897,N_4629);
nor UO_445 (O_445,N_4584,N_4755);
and UO_446 (O_446,N_4753,N_4526);
xnor UO_447 (O_447,N_4803,N_4631);
nor UO_448 (O_448,N_4852,N_4669);
and UO_449 (O_449,N_4780,N_4543);
and UO_450 (O_450,N_4542,N_4690);
nand UO_451 (O_451,N_4692,N_4736);
or UO_452 (O_452,N_4942,N_4751);
and UO_453 (O_453,N_4892,N_4878);
or UO_454 (O_454,N_4557,N_4875);
nand UO_455 (O_455,N_4572,N_4686);
or UO_456 (O_456,N_4984,N_4740);
nor UO_457 (O_457,N_4830,N_4976);
nand UO_458 (O_458,N_4950,N_4687);
and UO_459 (O_459,N_4856,N_4892);
or UO_460 (O_460,N_4854,N_4974);
xor UO_461 (O_461,N_4711,N_4628);
or UO_462 (O_462,N_4862,N_4942);
and UO_463 (O_463,N_4765,N_4932);
or UO_464 (O_464,N_4801,N_4718);
nor UO_465 (O_465,N_4798,N_4546);
nand UO_466 (O_466,N_4755,N_4669);
nor UO_467 (O_467,N_4681,N_4519);
nor UO_468 (O_468,N_4574,N_4745);
and UO_469 (O_469,N_4877,N_4832);
and UO_470 (O_470,N_4636,N_4736);
or UO_471 (O_471,N_4909,N_4704);
or UO_472 (O_472,N_4680,N_4917);
or UO_473 (O_473,N_4688,N_4673);
xnor UO_474 (O_474,N_4668,N_4886);
and UO_475 (O_475,N_4940,N_4815);
xnor UO_476 (O_476,N_4983,N_4504);
or UO_477 (O_477,N_4910,N_4582);
or UO_478 (O_478,N_4755,N_4546);
nor UO_479 (O_479,N_4633,N_4556);
nand UO_480 (O_480,N_4692,N_4554);
or UO_481 (O_481,N_4935,N_4784);
nor UO_482 (O_482,N_4808,N_4738);
xnor UO_483 (O_483,N_4553,N_4623);
or UO_484 (O_484,N_4807,N_4933);
xor UO_485 (O_485,N_4664,N_4749);
and UO_486 (O_486,N_4695,N_4786);
nor UO_487 (O_487,N_4751,N_4732);
and UO_488 (O_488,N_4559,N_4538);
or UO_489 (O_489,N_4816,N_4974);
or UO_490 (O_490,N_4906,N_4890);
nand UO_491 (O_491,N_4691,N_4572);
and UO_492 (O_492,N_4949,N_4595);
nand UO_493 (O_493,N_4696,N_4565);
xor UO_494 (O_494,N_4817,N_4841);
nor UO_495 (O_495,N_4977,N_4707);
nand UO_496 (O_496,N_4733,N_4543);
and UO_497 (O_497,N_4770,N_4511);
nor UO_498 (O_498,N_4914,N_4850);
or UO_499 (O_499,N_4735,N_4825);
nor UO_500 (O_500,N_4941,N_4735);
nand UO_501 (O_501,N_4751,N_4762);
nor UO_502 (O_502,N_4537,N_4799);
xnor UO_503 (O_503,N_4634,N_4944);
or UO_504 (O_504,N_4856,N_4623);
nor UO_505 (O_505,N_4566,N_4584);
or UO_506 (O_506,N_4534,N_4507);
xor UO_507 (O_507,N_4639,N_4516);
or UO_508 (O_508,N_4524,N_4612);
nor UO_509 (O_509,N_4737,N_4799);
xnor UO_510 (O_510,N_4662,N_4871);
or UO_511 (O_511,N_4607,N_4870);
or UO_512 (O_512,N_4816,N_4805);
nand UO_513 (O_513,N_4666,N_4508);
or UO_514 (O_514,N_4767,N_4788);
nor UO_515 (O_515,N_4632,N_4524);
xnor UO_516 (O_516,N_4777,N_4723);
nor UO_517 (O_517,N_4880,N_4692);
xor UO_518 (O_518,N_4680,N_4952);
xnor UO_519 (O_519,N_4961,N_4825);
xnor UO_520 (O_520,N_4741,N_4874);
or UO_521 (O_521,N_4742,N_4972);
or UO_522 (O_522,N_4921,N_4930);
and UO_523 (O_523,N_4612,N_4631);
or UO_524 (O_524,N_4828,N_4529);
or UO_525 (O_525,N_4896,N_4853);
nor UO_526 (O_526,N_4887,N_4869);
xnor UO_527 (O_527,N_4830,N_4989);
nor UO_528 (O_528,N_4991,N_4980);
nor UO_529 (O_529,N_4951,N_4704);
nor UO_530 (O_530,N_4732,N_4616);
nor UO_531 (O_531,N_4888,N_4930);
and UO_532 (O_532,N_4947,N_4972);
or UO_533 (O_533,N_4934,N_4531);
and UO_534 (O_534,N_4500,N_4874);
nor UO_535 (O_535,N_4524,N_4746);
xnor UO_536 (O_536,N_4924,N_4871);
nand UO_537 (O_537,N_4663,N_4529);
nor UO_538 (O_538,N_4924,N_4568);
nor UO_539 (O_539,N_4943,N_4538);
nand UO_540 (O_540,N_4551,N_4852);
xor UO_541 (O_541,N_4983,N_4746);
nor UO_542 (O_542,N_4689,N_4631);
nor UO_543 (O_543,N_4602,N_4795);
and UO_544 (O_544,N_4591,N_4845);
xnor UO_545 (O_545,N_4580,N_4736);
nand UO_546 (O_546,N_4837,N_4878);
nand UO_547 (O_547,N_4831,N_4664);
and UO_548 (O_548,N_4533,N_4845);
nand UO_549 (O_549,N_4977,N_4856);
and UO_550 (O_550,N_4657,N_4606);
or UO_551 (O_551,N_4501,N_4512);
xnor UO_552 (O_552,N_4694,N_4800);
nor UO_553 (O_553,N_4677,N_4982);
xnor UO_554 (O_554,N_4531,N_4867);
nand UO_555 (O_555,N_4832,N_4552);
or UO_556 (O_556,N_4711,N_4764);
or UO_557 (O_557,N_4765,N_4875);
nand UO_558 (O_558,N_4880,N_4981);
nand UO_559 (O_559,N_4611,N_4662);
xor UO_560 (O_560,N_4851,N_4910);
nand UO_561 (O_561,N_4534,N_4761);
nor UO_562 (O_562,N_4782,N_4649);
or UO_563 (O_563,N_4688,N_4619);
nor UO_564 (O_564,N_4698,N_4708);
and UO_565 (O_565,N_4880,N_4568);
nor UO_566 (O_566,N_4722,N_4851);
nor UO_567 (O_567,N_4652,N_4806);
or UO_568 (O_568,N_4698,N_4669);
nand UO_569 (O_569,N_4749,N_4644);
nor UO_570 (O_570,N_4912,N_4685);
nand UO_571 (O_571,N_4795,N_4674);
xor UO_572 (O_572,N_4804,N_4903);
or UO_573 (O_573,N_4627,N_4825);
xnor UO_574 (O_574,N_4928,N_4686);
xor UO_575 (O_575,N_4554,N_4739);
nand UO_576 (O_576,N_4707,N_4544);
and UO_577 (O_577,N_4964,N_4653);
and UO_578 (O_578,N_4812,N_4716);
xor UO_579 (O_579,N_4568,N_4926);
or UO_580 (O_580,N_4751,N_4910);
nand UO_581 (O_581,N_4744,N_4518);
or UO_582 (O_582,N_4921,N_4771);
or UO_583 (O_583,N_4820,N_4854);
xnor UO_584 (O_584,N_4631,N_4998);
xnor UO_585 (O_585,N_4511,N_4855);
or UO_586 (O_586,N_4996,N_4782);
or UO_587 (O_587,N_4661,N_4731);
or UO_588 (O_588,N_4781,N_4706);
and UO_589 (O_589,N_4602,N_4739);
nand UO_590 (O_590,N_4590,N_4638);
and UO_591 (O_591,N_4820,N_4798);
nor UO_592 (O_592,N_4567,N_4797);
and UO_593 (O_593,N_4696,N_4591);
nand UO_594 (O_594,N_4757,N_4611);
or UO_595 (O_595,N_4660,N_4578);
or UO_596 (O_596,N_4856,N_4930);
or UO_597 (O_597,N_4823,N_4726);
xor UO_598 (O_598,N_4625,N_4967);
nand UO_599 (O_599,N_4542,N_4887);
nor UO_600 (O_600,N_4960,N_4764);
or UO_601 (O_601,N_4580,N_4981);
and UO_602 (O_602,N_4806,N_4859);
nor UO_603 (O_603,N_4712,N_4592);
nor UO_604 (O_604,N_4737,N_4872);
or UO_605 (O_605,N_4656,N_4668);
or UO_606 (O_606,N_4901,N_4822);
xnor UO_607 (O_607,N_4909,N_4768);
xnor UO_608 (O_608,N_4921,N_4728);
nand UO_609 (O_609,N_4965,N_4556);
xnor UO_610 (O_610,N_4636,N_4996);
nor UO_611 (O_611,N_4817,N_4771);
and UO_612 (O_612,N_4677,N_4564);
and UO_613 (O_613,N_4830,N_4973);
xor UO_614 (O_614,N_4670,N_4795);
or UO_615 (O_615,N_4942,N_4762);
nor UO_616 (O_616,N_4911,N_4574);
or UO_617 (O_617,N_4812,N_4539);
xnor UO_618 (O_618,N_4564,N_4559);
nand UO_619 (O_619,N_4615,N_4987);
or UO_620 (O_620,N_4886,N_4653);
nand UO_621 (O_621,N_4819,N_4755);
nand UO_622 (O_622,N_4976,N_4747);
nor UO_623 (O_623,N_4796,N_4932);
nand UO_624 (O_624,N_4549,N_4541);
nand UO_625 (O_625,N_4500,N_4628);
nand UO_626 (O_626,N_4784,N_4514);
and UO_627 (O_627,N_4596,N_4591);
nor UO_628 (O_628,N_4904,N_4890);
xor UO_629 (O_629,N_4997,N_4773);
xor UO_630 (O_630,N_4528,N_4731);
nor UO_631 (O_631,N_4799,N_4585);
nor UO_632 (O_632,N_4882,N_4723);
or UO_633 (O_633,N_4730,N_4814);
xor UO_634 (O_634,N_4550,N_4654);
and UO_635 (O_635,N_4927,N_4894);
nand UO_636 (O_636,N_4911,N_4710);
xnor UO_637 (O_637,N_4795,N_4649);
and UO_638 (O_638,N_4630,N_4572);
nor UO_639 (O_639,N_4593,N_4675);
or UO_640 (O_640,N_4843,N_4886);
and UO_641 (O_641,N_4691,N_4726);
and UO_642 (O_642,N_4560,N_4565);
or UO_643 (O_643,N_4824,N_4949);
and UO_644 (O_644,N_4597,N_4610);
or UO_645 (O_645,N_4946,N_4581);
nor UO_646 (O_646,N_4831,N_4772);
xnor UO_647 (O_647,N_4526,N_4819);
xor UO_648 (O_648,N_4603,N_4840);
or UO_649 (O_649,N_4898,N_4739);
xnor UO_650 (O_650,N_4650,N_4819);
nor UO_651 (O_651,N_4698,N_4573);
and UO_652 (O_652,N_4795,N_4929);
xnor UO_653 (O_653,N_4821,N_4699);
nor UO_654 (O_654,N_4705,N_4888);
nor UO_655 (O_655,N_4667,N_4999);
or UO_656 (O_656,N_4593,N_4824);
and UO_657 (O_657,N_4874,N_4993);
nor UO_658 (O_658,N_4957,N_4900);
nand UO_659 (O_659,N_4906,N_4753);
and UO_660 (O_660,N_4920,N_4670);
or UO_661 (O_661,N_4752,N_4852);
nor UO_662 (O_662,N_4621,N_4500);
nand UO_663 (O_663,N_4561,N_4807);
nor UO_664 (O_664,N_4803,N_4868);
nand UO_665 (O_665,N_4552,N_4871);
or UO_666 (O_666,N_4817,N_4557);
xor UO_667 (O_667,N_4528,N_4600);
nor UO_668 (O_668,N_4662,N_4542);
nand UO_669 (O_669,N_4629,N_4972);
nor UO_670 (O_670,N_4603,N_4745);
nor UO_671 (O_671,N_4517,N_4534);
nand UO_672 (O_672,N_4601,N_4834);
nand UO_673 (O_673,N_4554,N_4697);
and UO_674 (O_674,N_4594,N_4944);
and UO_675 (O_675,N_4825,N_4927);
and UO_676 (O_676,N_4967,N_4881);
and UO_677 (O_677,N_4827,N_4876);
xor UO_678 (O_678,N_4700,N_4528);
nand UO_679 (O_679,N_4775,N_4677);
nor UO_680 (O_680,N_4855,N_4954);
or UO_681 (O_681,N_4611,N_4793);
xor UO_682 (O_682,N_4982,N_4707);
nor UO_683 (O_683,N_4900,N_4577);
and UO_684 (O_684,N_4851,N_4867);
nand UO_685 (O_685,N_4905,N_4883);
or UO_686 (O_686,N_4854,N_4867);
nor UO_687 (O_687,N_4584,N_4706);
nor UO_688 (O_688,N_4610,N_4806);
nor UO_689 (O_689,N_4886,N_4749);
nand UO_690 (O_690,N_4838,N_4932);
and UO_691 (O_691,N_4724,N_4766);
and UO_692 (O_692,N_4629,N_4775);
nor UO_693 (O_693,N_4979,N_4926);
and UO_694 (O_694,N_4828,N_4766);
nor UO_695 (O_695,N_4802,N_4903);
nor UO_696 (O_696,N_4974,N_4575);
or UO_697 (O_697,N_4711,N_4606);
xor UO_698 (O_698,N_4915,N_4921);
or UO_699 (O_699,N_4713,N_4555);
xnor UO_700 (O_700,N_4735,N_4951);
nand UO_701 (O_701,N_4773,N_4951);
and UO_702 (O_702,N_4753,N_4796);
or UO_703 (O_703,N_4822,N_4585);
nor UO_704 (O_704,N_4639,N_4789);
and UO_705 (O_705,N_4686,N_4847);
and UO_706 (O_706,N_4615,N_4978);
nor UO_707 (O_707,N_4941,N_4658);
nand UO_708 (O_708,N_4819,N_4918);
nor UO_709 (O_709,N_4829,N_4760);
nor UO_710 (O_710,N_4897,N_4510);
nand UO_711 (O_711,N_4618,N_4737);
nand UO_712 (O_712,N_4805,N_4522);
nor UO_713 (O_713,N_4621,N_4840);
nor UO_714 (O_714,N_4689,N_4704);
and UO_715 (O_715,N_4665,N_4686);
and UO_716 (O_716,N_4934,N_4676);
nand UO_717 (O_717,N_4862,N_4819);
nand UO_718 (O_718,N_4959,N_4731);
nand UO_719 (O_719,N_4956,N_4537);
or UO_720 (O_720,N_4976,N_4703);
and UO_721 (O_721,N_4859,N_4550);
xnor UO_722 (O_722,N_4639,N_4592);
xor UO_723 (O_723,N_4939,N_4820);
nand UO_724 (O_724,N_4962,N_4981);
xor UO_725 (O_725,N_4784,N_4886);
nand UO_726 (O_726,N_4679,N_4634);
nand UO_727 (O_727,N_4854,N_4827);
nor UO_728 (O_728,N_4919,N_4975);
or UO_729 (O_729,N_4919,N_4507);
nor UO_730 (O_730,N_4865,N_4744);
and UO_731 (O_731,N_4879,N_4951);
nand UO_732 (O_732,N_4883,N_4592);
xor UO_733 (O_733,N_4906,N_4648);
or UO_734 (O_734,N_4813,N_4997);
or UO_735 (O_735,N_4896,N_4650);
nor UO_736 (O_736,N_4891,N_4869);
and UO_737 (O_737,N_4771,N_4828);
or UO_738 (O_738,N_4742,N_4926);
xnor UO_739 (O_739,N_4660,N_4524);
nor UO_740 (O_740,N_4831,N_4813);
xnor UO_741 (O_741,N_4571,N_4514);
xnor UO_742 (O_742,N_4951,N_4609);
and UO_743 (O_743,N_4758,N_4768);
and UO_744 (O_744,N_4889,N_4621);
or UO_745 (O_745,N_4712,N_4833);
and UO_746 (O_746,N_4591,N_4833);
and UO_747 (O_747,N_4703,N_4885);
xor UO_748 (O_748,N_4969,N_4824);
nor UO_749 (O_749,N_4521,N_4507);
and UO_750 (O_750,N_4547,N_4520);
or UO_751 (O_751,N_4857,N_4627);
xor UO_752 (O_752,N_4929,N_4931);
nor UO_753 (O_753,N_4574,N_4799);
and UO_754 (O_754,N_4873,N_4964);
nor UO_755 (O_755,N_4861,N_4540);
and UO_756 (O_756,N_4524,N_4676);
nor UO_757 (O_757,N_4841,N_4919);
nor UO_758 (O_758,N_4990,N_4786);
nor UO_759 (O_759,N_4943,N_4579);
or UO_760 (O_760,N_4626,N_4790);
nand UO_761 (O_761,N_4706,N_4707);
xnor UO_762 (O_762,N_4671,N_4718);
and UO_763 (O_763,N_4992,N_4698);
xnor UO_764 (O_764,N_4740,N_4969);
xor UO_765 (O_765,N_4810,N_4716);
nor UO_766 (O_766,N_4738,N_4765);
or UO_767 (O_767,N_4735,N_4762);
or UO_768 (O_768,N_4647,N_4918);
or UO_769 (O_769,N_4777,N_4653);
xnor UO_770 (O_770,N_4815,N_4833);
nor UO_771 (O_771,N_4680,N_4948);
and UO_772 (O_772,N_4936,N_4998);
nor UO_773 (O_773,N_4707,N_4753);
and UO_774 (O_774,N_4646,N_4737);
nand UO_775 (O_775,N_4753,N_4849);
xor UO_776 (O_776,N_4717,N_4898);
xnor UO_777 (O_777,N_4565,N_4735);
nor UO_778 (O_778,N_4867,N_4734);
and UO_779 (O_779,N_4544,N_4603);
or UO_780 (O_780,N_4740,N_4621);
xnor UO_781 (O_781,N_4765,N_4915);
xnor UO_782 (O_782,N_4880,N_4577);
or UO_783 (O_783,N_4834,N_4689);
nand UO_784 (O_784,N_4908,N_4501);
and UO_785 (O_785,N_4509,N_4971);
nor UO_786 (O_786,N_4680,N_4513);
xor UO_787 (O_787,N_4898,N_4674);
and UO_788 (O_788,N_4917,N_4624);
xnor UO_789 (O_789,N_4606,N_4544);
nor UO_790 (O_790,N_4607,N_4521);
xor UO_791 (O_791,N_4842,N_4781);
xor UO_792 (O_792,N_4583,N_4635);
nor UO_793 (O_793,N_4535,N_4772);
xnor UO_794 (O_794,N_4577,N_4603);
nor UO_795 (O_795,N_4661,N_4883);
or UO_796 (O_796,N_4851,N_4751);
xor UO_797 (O_797,N_4837,N_4682);
nor UO_798 (O_798,N_4694,N_4904);
nor UO_799 (O_799,N_4896,N_4935);
nand UO_800 (O_800,N_4534,N_4902);
xor UO_801 (O_801,N_4918,N_4930);
nand UO_802 (O_802,N_4772,N_4725);
and UO_803 (O_803,N_4753,N_4951);
and UO_804 (O_804,N_4784,N_4630);
or UO_805 (O_805,N_4667,N_4854);
and UO_806 (O_806,N_4748,N_4881);
or UO_807 (O_807,N_4524,N_4689);
and UO_808 (O_808,N_4504,N_4533);
or UO_809 (O_809,N_4868,N_4891);
or UO_810 (O_810,N_4861,N_4945);
xnor UO_811 (O_811,N_4944,N_4675);
or UO_812 (O_812,N_4614,N_4620);
nand UO_813 (O_813,N_4715,N_4537);
and UO_814 (O_814,N_4555,N_4924);
nand UO_815 (O_815,N_4666,N_4949);
nand UO_816 (O_816,N_4653,N_4563);
nor UO_817 (O_817,N_4863,N_4551);
nand UO_818 (O_818,N_4545,N_4879);
nand UO_819 (O_819,N_4782,N_4726);
nor UO_820 (O_820,N_4635,N_4970);
and UO_821 (O_821,N_4710,N_4928);
xor UO_822 (O_822,N_4689,N_4653);
or UO_823 (O_823,N_4927,N_4629);
nand UO_824 (O_824,N_4529,N_4732);
xnor UO_825 (O_825,N_4929,N_4885);
or UO_826 (O_826,N_4731,N_4750);
or UO_827 (O_827,N_4826,N_4894);
or UO_828 (O_828,N_4983,N_4980);
or UO_829 (O_829,N_4513,N_4759);
and UO_830 (O_830,N_4592,N_4783);
nor UO_831 (O_831,N_4565,N_4870);
nand UO_832 (O_832,N_4854,N_4763);
nand UO_833 (O_833,N_4604,N_4745);
nand UO_834 (O_834,N_4949,N_4665);
nor UO_835 (O_835,N_4560,N_4577);
or UO_836 (O_836,N_4619,N_4533);
or UO_837 (O_837,N_4723,N_4554);
or UO_838 (O_838,N_4566,N_4901);
nor UO_839 (O_839,N_4586,N_4988);
xor UO_840 (O_840,N_4527,N_4871);
nand UO_841 (O_841,N_4766,N_4596);
or UO_842 (O_842,N_4694,N_4637);
nor UO_843 (O_843,N_4585,N_4740);
xor UO_844 (O_844,N_4867,N_4933);
nand UO_845 (O_845,N_4772,N_4946);
xnor UO_846 (O_846,N_4504,N_4510);
and UO_847 (O_847,N_4825,N_4611);
or UO_848 (O_848,N_4836,N_4580);
nand UO_849 (O_849,N_4814,N_4783);
nor UO_850 (O_850,N_4651,N_4878);
nand UO_851 (O_851,N_4915,N_4767);
nor UO_852 (O_852,N_4768,N_4559);
and UO_853 (O_853,N_4510,N_4649);
xnor UO_854 (O_854,N_4661,N_4602);
or UO_855 (O_855,N_4677,N_4787);
nor UO_856 (O_856,N_4873,N_4846);
xnor UO_857 (O_857,N_4528,N_4779);
and UO_858 (O_858,N_4973,N_4742);
xnor UO_859 (O_859,N_4511,N_4891);
nor UO_860 (O_860,N_4722,N_4853);
nand UO_861 (O_861,N_4904,N_4701);
or UO_862 (O_862,N_4861,N_4582);
nand UO_863 (O_863,N_4935,N_4603);
and UO_864 (O_864,N_4918,N_4804);
xnor UO_865 (O_865,N_4810,N_4729);
xnor UO_866 (O_866,N_4942,N_4656);
and UO_867 (O_867,N_4816,N_4999);
nor UO_868 (O_868,N_4551,N_4950);
and UO_869 (O_869,N_4664,N_4613);
xor UO_870 (O_870,N_4764,N_4746);
nor UO_871 (O_871,N_4869,N_4979);
nand UO_872 (O_872,N_4517,N_4987);
xor UO_873 (O_873,N_4885,N_4854);
and UO_874 (O_874,N_4795,N_4524);
nand UO_875 (O_875,N_4592,N_4585);
xor UO_876 (O_876,N_4575,N_4524);
or UO_877 (O_877,N_4608,N_4805);
or UO_878 (O_878,N_4604,N_4675);
nor UO_879 (O_879,N_4594,N_4892);
xor UO_880 (O_880,N_4762,N_4641);
nand UO_881 (O_881,N_4658,N_4725);
xnor UO_882 (O_882,N_4929,N_4865);
xor UO_883 (O_883,N_4622,N_4844);
nor UO_884 (O_884,N_4969,N_4616);
nand UO_885 (O_885,N_4769,N_4682);
and UO_886 (O_886,N_4742,N_4557);
nand UO_887 (O_887,N_4802,N_4918);
or UO_888 (O_888,N_4775,N_4630);
nand UO_889 (O_889,N_4732,N_4543);
nor UO_890 (O_890,N_4577,N_4665);
and UO_891 (O_891,N_4839,N_4904);
or UO_892 (O_892,N_4601,N_4777);
and UO_893 (O_893,N_4683,N_4581);
nor UO_894 (O_894,N_4697,N_4941);
or UO_895 (O_895,N_4590,N_4729);
or UO_896 (O_896,N_4509,N_4805);
or UO_897 (O_897,N_4998,N_4771);
and UO_898 (O_898,N_4637,N_4581);
nor UO_899 (O_899,N_4995,N_4856);
nor UO_900 (O_900,N_4704,N_4800);
nand UO_901 (O_901,N_4590,N_4507);
xnor UO_902 (O_902,N_4897,N_4740);
or UO_903 (O_903,N_4819,N_4747);
and UO_904 (O_904,N_4578,N_4863);
nand UO_905 (O_905,N_4710,N_4662);
or UO_906 (O_906,N_4996,N_4900);
nor UO_907 (O_907,N_4638,N_4911);
or UO_908 (O_908,N_4850,N_4577);
nor UO_909 (O_909,N_4918,N_4831);
xnor UO_910 (O_910,N_4683,N_4783);
and UO_911 (O_911,N_4992,N_4621);
xnor UO_912 (O_912,N_4514,N_4541);
nand UO_913 (O_913,N_4668,N_4652);
or UO_914 (O_914,N_4841,N_4918);
nand UO_915 (O_915,N_4604,N_4641);
and UO_916 (O_916,N_4988,N_4609);
and UO_917 (O_917,N_4682,N_4990);
xor UO_918 (O_918,N_4932,N_4805);
and UO_919 (O_919,N_4928,N_4618);
xor UO_920 (O_920,N_4616,N_4548);
or UO_921 (O_921,N_4684,N_4915);
nor UO_922 (O_922,N_4571,N_4606);
nor UO_923 (O_923,N_4739,N_4588);
and UO_924 (O_924,N_4907,N_4641);
and UO_925 (O_925,N_4882,N_4686);
or UO_926 (O_926,N_4618,N_4930);
or UO_927 (O_927,N_4992,N_4980);
or UO_928 (O_928,N_4581,N_4580);
xnor UO_929 (O_929,N_4895,N_4947);
or UO_930 (O_930,N_4975,N_4887);
or UO_931 (O_931,N_4825,N_4671);
and UO_932 (O_932,N_4531,N_4514);
xnor UO_933 (O_933,N_4867,N_4732);
xor UO_934 (O_934,N_4914,N_4718);
nor UO_935 (O_935,N_4791,N_4755);
nor UO_936 (O_936,N_4953,N_4601);
and UO_937 (O_937,N_4506,N_4754);
xnor UO_938 (O_938,N_4891,N_4503);
and UO_939 (O_939,N_4504,N_4895);
xnor UO_940 (O_940,N_4736,N_4975);
xnor UO_941 (O_941,N_4953,N_4644);
and UO_942 (O_942,N_4523,N_4932);
xnor UO_943 (O_943,N_4726,N_4952);
and UO_944 (O_944,N_4769,N_4636);
or UO_945 (O_945,N_4973,N_4980);
nor UO_946 (O_946,N_4952,N_4851);
xor UO_947 (O_947,N_4871,N_4781);
or UO_948 (O_948,N_4755,N_4926);
or UO_949 (O_949,N_4885,N_4627);
or UO_950 (O_950,N_4630,N_4632);
and UO_951 (O_951,N_4885,N_4927);
nand UO_952 (O_952,N_4549,N_4782);
nor UO_953 (O_953,N_4948,N_4789);
and UO_954 (O_954,N_4757,N_4570);
nor UO_955 (O_955,N_4907,N_4593);
or UO_956 (O_956,N_4706,N_4822);
or UO_957 (O_957,N_4534,N_4982);
nand UO_958 (O_958,N_4754,N_4900);
nand UO_959 (O_959,N_4888,N_4838);
nor UO_960 (O_960,N_4813,N_4896);
nor UO_961 (O_961,N_4715,N_4991);
nand UO_962 (O_962,N_4656,N_4558);
nand UO_963 (O_963,N_4834,N_4842);
xnor UO_964 (O_964,N_4873,N_4603);
and UO_965 (O_965,N_4904,N_4769);
and UO_966 (O_966,N_4804,N_4598);
nor UO_967 (O_967,N_4941,N_4598);
nand UO_968 (O_968,N_4830,N_4600);
xnor UO_969 (O_969,N_4943,N_4679);
or UO_970 (O_970,N_4962,N_4546);
nor UO_971 (O_971,N_4885,N_4715);
xnor UO_972 (O_972,N_4953,N_4885);
nor UO_973 (O_973,N_4930,N_4512);
and UO_974 (O_974,N_4705,N_4586);
xor UO_975 (O_975,N_4989,N_4847);
xnor UO_976 (O_976,N_4702,N_4706);
or UO_977 (O_977,N_4961,N_4917);
or UO_978 (O_978,N_4887,N_4589);
and UO_979 (O_979,N_4683,N_4702);
nor UO_980 (O_980,N_4860,N_4516);
or UO_981 (O_981,N_4575,N_4729);
and UO_982 (O_982,N_4540,N_4787);
or UO_983 (O_983,N_4862,N_4700);
and UO_984 (O_984,N_4891,N_4674);
xnor UO_985 (O_985,N_4750,N_4714);
or UO_986 (O_986,N_4745,N_4902);
or UO_987 (O_987,N_4675,N_4712);
or UO_988 (O_988,N_4899,N_4813);
and UO_989 (O_989,N_4787,N_4510);
and UO_990 (O_990,N_4613,N_4905);
xnor UO_991 (O_991,N_4558,N_4614);
nand UO_992 (O_992,N_4725,N_4800);
or UO_993 (O_993,N_4540,N_4580);
xnor UO_994 (O_994,N_4964,N_4502);
or UO_995 (O_995,N_4847,N_4815);
and UO_996 (O_996,N_4853,N_4595);
nand UO_997 (O_997,N_4803,N_4622);
xnor UO_998 (O_998,N_4780,N_4849);
nor UO_999 (O_999,N_4692,N_4970);
endmodule