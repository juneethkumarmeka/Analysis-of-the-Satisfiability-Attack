module basic_2500_25000_3000_125_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1861,In_1163);
nor U1 (N_1,In_1245,In_847);
and U2 (N_2,In_823,In_2266);
xor U3 (N_3,In_424,In_372);
xnor U4 (N_4,In_1486,In_562);
or U5 (N_5,In_2452,In_831);
nand U6 (N_6,In_206,In_510);
xnor U7 (N_7,In_1986,In_1519);
nand U8 (N_8,In_2048,In_2391);
and U9 (N_9,In_1025,In_989);
and U10 (N_10,In_2028,In_1637);
or U11 (N_11,In_1941,In_2331);
and U12 (N_12,In_1318,In_878);
nor U13 (N_13,In_1068,In_2160);
nor U14 (N_14,In_1288,In_144);
and U15 (N_15,In_1146,In_876);
and U16 (N_16,In_2435,In_289);
and U17 (N_17,In_811,In_2095);
nor U18 (N_18,In_610,In_404);
xor U19 (N_19,In_646,In_330);
xor U20 (N_20,In_1174,In_1239);
nand U21 (N_21,In_292,In_1868);
and U22 (N_22,In_502,In_1278);
and U23 (N_23,In_664,In_1022);
nand U24 (N_24,In_1058,In_12);
nand U25 (N_25,In_1301,In_1969);
xor U26 (N_26,In_2078,In_740);
nand U27 (N_27,In_2478,In_1963);
or U28 (N_28,In_2499,In_1414);
xnor U29 (N_29,In_2246,In_1464);
or U30 (N_30,In_1212,In_84);
xor U31 (N_31,In_2370,In_1125);
and U32 (N_32,In_2051,In_544);
nor U33 (N_33,In_2193,In_1470);
or U34 (N_34,In_737,In_370);
or U35 (N_35,In_489,In_963);
or U36 (N_36,In_2100,In_909);
nand U37 (N_37,In_215,In_1865);
or U38 (N_38,In_301,In_739);
xnor U39 (N_39,In_1319,In_600);
xor U40 (N_40,In_1635,In_1315);
nor U41 (N_41,In_1777,In_478);
xor U42 (N_42,In_1972,In_1467);
and U43 (N_43,In_1221,In_1912);
nor U44 (N_44,In_1211,In_304);
or U45 (N_45,In_114,In_2018);
and U46 (N_46,In_157,In_1766);
and U47 (N_47,In_2173,In_408);
and U48 (N_48,In_2453,In_2205);
xor U49 (N_49,In_1048,In_1256);
nand U50 (N_50,In_198,In_830);
nor U51 (N_51,In_1393,In_2359);
and U52 (N_52,In_1989,In_894);
nand U53 (N_53,In_1131,In_2345);
or U54 (N_54,In_712,In_1592);
nand U55 (N_55,In_797,In_1415);
or U56 (N_56,In_2374,In_2069);
nor U57 (N_57,In_1075,In_1425);
and U58 (N_58,In_33,In_842);
nand U59 (N_59,In_1533,In_1725);
nand U60 (N_60,In_1540,In_619);
nand U61 (N_61,In_549,In_711);
or U62 (N_62,In_103,In_1517);
nor U63 (N_63,In_18,In_2439);
or U64 (N_64,In_1490,In_921);
and U65 (N_65,In_1126,In_1175);
or U66 (N_66,In_1437,In_349);
and U67 (N_67,In_61,In_1276);
and U68 (N_68,In_940,In_633);
and U69 (N_69,In_2420,In_2187);
nor U70 (N_70,In_280,In_327);
nand U71 (N_71,In_1796,In_2011);
nor U72 (N_72,In_997,In_283);
nor U73 (N_73,In_1653,In_1896);
nand U74 (N_74,In_635,In_800);
and U75 (N_75,In_1597,In_1583);
nand U76 (N_76,In_200,In_1182);
nand U77 (N_77,In_1111,In_1917);
nor U78 (N_78,In_550,In_1613);
nor U79 (N_79,In_2274,In_824);
or U80 (N_80,In_1447,In_240);
or U81 (N_81,In_1909,In_604);
nand U82 (N_82,In_360,In_66);
nor U83 (N_83,In_2176,In_90);
nand U84 (N_84,In_249,In_165);
nor U85 (N_85,In_1718,In_852);
and U86 (N_86,In_1419,In_538);
nor U87 (N_87,In_775,In_2200);
or U88 (N_88,In_2158,In_2035);
nor U89 (N_89,In_1118,In_925);
or U90 (N_90,In_701,In_1678);
or U91 (N_91,In_1047,In_1140);
nand U92 (N_92,In_893,In_1112);
and U93 (N_93,In_2194,In_1784);
nor U94 (N_94,In_273,In_976);
or U95 (N_95,In_728,In_906);
nor U96 (N_96,In_34,In_1474);
and U97 (N_97,In_1325,In_93);
xnor U98 (N_98,In_2023,In_1975);
nand U99 (N_99,In_1355,In_2254);
nand U100 (N_100,In_275,In_1538);
nand U101 (N_101,In_576,In_1940);
nor U102 (N_102,In_2057,In_2324);
xnor U103 (N_103,In_67,In_261);
nand U104 (N_104,In_1968,In_445);
xor U105 (N_105,In_693,In_465);
or U106 (N_106,In_325,In_1685);
nand U107 (N_107,In_92,In_2099);
xor U108 (N_108,In_1114,In_645);
xor U109 (N_109,In_761,In_2358);
or U110 (N_110,In_559,In_133);
xnor U111 (N_111,In_312,In_802);
xor U112 (N_112,In_1847,In_410);
and U113 (N_113,In_691,In_1805);
nor U114 (N_114,In_613,In_1743);
or U115 (N_115,In_1370,In_2446);
xor U116 (N_116,In_1273,In_1709);
nor U117 (N_117,In_1042,In_453);
and U118 (N_118,In_581,In_2288);
nor U119 (N_119,In_203,In_1200);
or U120 (N_120,In_2143,In_1618);
nand U121 (N_121,In_160,In_520);
nor U122 (N_122,In_1888,In_1807);
or U123 (N_123,In_417,In_1109);
xnor U124 (N_124,In_362,In_1057);
or U125 (N_125,In_1387,In_2076);
or U126 (N_126,In_1116,In_2091);
or U127 (N_127,In_85,In_405);
nor U128 (N_128,In_2214,In_2423);
xnor U129 (N_129,In_1851,In_1281);
and U130 (N_130,In_780,In_2189);
xor U131 (N_131,In_1491,In_1157);
xnor U132 (N_132,In_1894,In_773);
or U133 (N_133,In_2341,In_2226);
and U134 (N_134,In_1161,In_1552);
xnor U135 (N_135,In_853,In_1611);
nor U136 (N_136,In_384,In_742);
nand U137 (N_137,In_2025,In_1401);
or U138 (N_138,In_794,In_340);
nand U139 (N_139,In_173,In_1361);
xor U140 (N_140,In_1086,In_2298);
and U141 (N_141,In_1426,In_1332);
and U142 (N_142,In_40,In_426);
nand U143 (N_143,In_522,In_1293);
or U144 (N_144,In_716,In_1787);
nand U145 (N_145,In_1554,In_2291);
or U146 (N_146,In_1832,In_653);
and U147 (N_147,In_2191,In_1850);
nand U148 (N_148,In_890,In_607);
xnor U149 (N_149,In_837,In_952);
nand U150 (N_150,In_936,In_1765);
or U151 (N_151,In_2265,In_386);
nor U152 (N_152,In_2042,In_10);
and U153 (N_153,In_22,In_922);
or U154 (N_154,In_651,In_2348);
or U155 (N_155,In_1323,In_2400);
nor U156 (N_156,In_400,In_590);
xnor U157 (N_157,In_785,In_2333);
nor U158 (N_158,In_1779,In_594);
and U159 (N_159,In_1976,In_1988);
xnor U160 (N_160,In_1340,In_1740);
nor U161 (N_161,In_1270,In_1795);
xnor U162 (N_162,In_766,In_1162);
nand U163 (N_163,In_2202,In_1672);
nand U164 (N_164,In_1403,In_2123);
nor U165 (N_165,In_1671,In_2212);
xnor U166 (N_166,In_606,In_428);
nor U167 (N_167,In_1735,In_2043);
and U168 (N_168,In_191,In_756);
and U169 (N_169,In_390,In_927);
and U170 (N_170,In_436,In_1308);
or U171 (N_171,In_2014,In_551);
xnor U172 (N_172,In_1910,In_271);
nor U173 (N_173,In_1781,In_109);
nor U174 (N_174,In_1745,In_2149);
and U175 (N_175,In_174,In_2422);
nand U176 (N_176,In_2007,In_2454);
nor U177 (N_177,In_1700,In_298);
nand U178 (N_178,In_31,In_625);
or U179 (N_179,In_1197,In_1139);
and U180 (N_180,In_490,In_1764);
nor U181 (N_181,In_726,In_214);
or U182 (N_182,In_262,In_965);
nor U183 (N_183,In_648,In_1166);
nor U184 (N_184,In_611,In_582);
nor U185 (N_185,In_1037,In_1721);
nor U186 (N_186,In_1237,In_668);
or U187 (N_187,In_112,In_2162);
nand U188 (N_188,In_2350,In_2171);
and U189 (N_189,In_1626,In_1946);
xor U190 (N_190,In_820,In_1181);
or U191 (N_191,In_1374,In_375);
nor U192 (N_192,In_2383,In_1217);
xor U193 (N_193,In_1170,In_284);
nand U194 (N_194,In_928,In_2244);
or U195 (N_195,In_2090,In_844);
xnor U196 (N_196,In_2394,In_720);
and U197 (N_197,In_530,In_1826);
or U198 (N_198,In_419,In_2306);
or U199 (N_199,In_345,In_185);
nand U200 (N_200,In_1578,In_96);
or U201 (N_201,In_2113,In_224);
and U202 (N_202,In_964,In_2027);
or U203 (N_203,In_1665,In_1012);
or U204 (N_204,In_1982,In_2085);
or U205 (N_205,In_113,N_63);
or U206 (N_206,In_973,In_88);
nand U207 (N_207,In_1882,In_1966);
nand U208 (N_208,In_320,In_1974);
or U209 (N_209,In_2138,N_182);
nor U210 (N_210,In_1821,In_1459);
nand U211 (N_211,In_1886,In_1351);
xor U212 (N_212,In_2355,N_57);
and U213 (N_213,In_300,In_2468);
nand U214 (N_214,In_1999,In_131);
or U215 (N_215,In_1099,In_1532);
nand U216 (N_216,In_1590,In_334);
nor U217 (N_217,In_988,In_621);
and U218 (N_218,In_279,In_1349);
nand U219 (N_219,In_168,In_2197);
xnor U220 (N_220,In_220,N_79);
or U221 (N_221,In_555,In_2210);
nand U222 (N_222,In_1680,In_1366);
nand U223 (N_223,In_752,In_1291);
and U224 (N_224,In_2408,In_2281);
xor U225 (N_225,In_2242,N_11);
xnor U226 (N_226,In_1229,In_1000);
nor U227 (N_227,In_42,In_1327);
and U228 (N_228,In_667,In_1246);
nor U229 (N_229,N_110,In_238);
and U230 (N_230,In_1621,In_1727);
or U231 (N_231,In_1185,In_1376);
nand U232 (N_232,In_931,In_654);
and U233 (N_233,In_1268,In_1412);
nor U234 (N_234,In_950,In_2001);
nand U235 (N_235,In_946,In_727);
or U236 (N_236,In_1294,In_1046);
or U237 (N_237,In_1479,In_583);
nor U238 (N_238,In_76,In_601);
and U239 (N_239,In_1708,In_1925);
nand U240 (N_240,In_2260,In_1069);
nor U241 (N_241,N_111,In_122);
nor U242 (N_242,In_1601,In_515);
xor U243 (N_243,In_73,In_1544);
xnor U244 (N_244,In_2185,In_1669);
nand U245 (N_245,In_860,In_286);
nor U246 (N_246,In_916,In_573);
and U247 (N_247,N_133,In_7);
nor U248 (N_248,In_2311,In_873);
or U249 (N_249,In_2141,In_1926);
nand U250 (N_250,In_2473,In_926);
xor U251 (N_251,In_984,In_1386);
nor U252 (N_252,In_361,N_139);
nor U253 (N_253,In_542,In_764);
xnor U254 (N_254,In_702,In_1790);
nor U255 (N_255,In_485,In_242);
or U256 (N_256,In_1799,In_38);
nand U257 (N_257,In_705,N_174);
nand U258 (N_258,In_2296,In_1548);
and U259 (N_259,In_881,In_2406);
or U260 (N_260,In_1101,In_1560);
nand U261 (N_261,In_1205,In_1612);
and U262 (N_262,In_1244,In_2405);
nand U263 (N_263,In_1056,In_2065);
and U264 (N_264,In_1493,In_1622);
nor U265 (N_265,In_908,In_2012);
or U266 (N_266,In_1749,N_103);
nor U267 (N_267,In_1756,In_995);
or U268 (N_268,In_476,In_867);
nor U269 (N_269,In_1593,N_9);
nor U270 (N_270,In_817,N_104);
nor U271 (N_271,In_1924,In_2310);
or U272 (N_272,N_166,In_2230);
nor U273 (N_273,In_2371,In_1512);
or U274 (N_274,In_430,N_99);
or U275 (N_275,N_40,In_1417);
xor U276 (N_276,In_1520,In_1701);
or U277 (N_277,In_2132,In_1916);
or U278 (N_278,In_1305,In_2096);
xnor U279 (N_279,In_1528,N_50);
nor U280 (N_280,In_1202,In_673);
or U281 (N_281,In_1248,In_529);
nor U282 (N_282,In_420,In_368);
or U283 (N_283,In_321,In_1816);
nor U284 (N_284,In_1335,In_1130);
xnor U285 (N_285,In_83,In_987);
nor U286 (N_286,In_905,N_91);
nor U287 (N_287,In_1176,In_2407);
or U288 (N_288,In_2077,In_137);
or U289 (N_289,In_1364,In_1298);
or U290 (N_290,N_175,In_1951);
and U291 (N_291,In_1516,In_1629);
nor U292 (N_292,In_159,N_149);
nor U293 (N_293,In_1550,In_1215);
and U294 (N_294,In_725,In_557);
nor U295 (N_295,In_929,In_2481);
xnor U296 (N_296,N_130,In_1715);
xor U297 (N_297,In_1646,In_1326);
nor U298 (N_298,In_655,In_1257);
nor U299 (N_299,In_1218,N_10);
or U300 (N_300,In_291,N_115);
nor U301 (N_301,N_101,In_1150);
xnor U302 (N_302,In_541,In_2102);
nand U303 (N_303,In_599,In_111);
nand U304 (N_304,In_644,In_1275);
nor U305 (N_305,In_49,In_1853);
xnor U306 (N_306,N_29,In_247);
and U307 (N_307,In_211,In_98);
or U308 (N_308,In_2322,In_2021);
nand U309 (N_309,In_1014,In_1300);
xor U310 (N_310,In_227,In_841);
and U311 (N_311,In_866,In_153);
and U312 (N_312,In_650,In_1943);
and U313 (N_313,In_1103,In_1418);
nor U314 (N_314,In_996,In_1854);
nand U315 (N_315,In_1303,In_2235);
or U316 (N_316,N_77,N_45);
nor U317 (N_317,In_2493,In_2047);
xnor U318 (N_318,In_2236,In_1785);
nor U319 (N_319,In_2257,In_1945);
or U320 (N_320,In_1586,In_1591);
nor U321 (N_321,In_2425,In_307);
and U322 (N_322,In_1371,In_1707);
xor U323 (N_323,In_353,In_782);
and U324 (N_324,In_318,N_156);
nand U325 (N_325,In_388,In_1884);
xnor U326 (N_326,In_2232,In_754);
xnor U327 (N_327,N_122,In_1249);
xnor U328 (N_328,In_1522,In_57);
or U329 (N_329,In_1067,In_1953);
xnor U330 (N_330,In_907,In_1242);
xnor U331 (N_331,In_1171,In_641);
or U332 (N_332,In_1456,In_1135);
xnor U333 (N_333,In_212,In_432);
xor U334 (N_334,In_1050,In_868);
xor U335 (N_335,N_134,In_439);
nand U336 (N_336,In_1353,In_1889);
nor U337 (N_337,In_1158,In_993);
or U338 (N_338,In_942,N_25);
or U339 (N_339,In_2179,In_1993);
and U340 (N_340,In_851,In_1193);
xor U341 (N_341,N_38,In_1077);
nor U342 (N_342,In_254,In_865);
xor U343 (N_343,In_1453,In_642);
or U344 (N_344,In_2395,In_229);
nor U345 (N_345,In_1570,In_1584);
nand U346 (N_346,In_1084,N_148);
or U347 (N_347,In_2484,In_2492);
nor U348 (N_348,In_1450,In_1880);
nor U349 (N_349,In_1480,In_2362);
nand U350 (N_350,N_145,In_1020);
nor U351 (N_351,In_1521,In_1706);
nand U352 (N_352,N_5,In_1682);
nand U353 (N_353,N_167,In_1726);
and U354 (N_354,N_184,In_1392);
nor U355 (N_355,In_887,In_679);
xor U356 (N_356,In_2120,In_1814);
nand U357 (N_357,In_1524,In_1530);
or U358 (N_358,In_1119,In_2292);
or U359 (N_359,In_1639,In_2170);
nand U360 (N_360,In_1028,In_571);
nand U361 (N_361,In_431,In_1149);
nand U362 (N_362,In_1169,In_1192);
nor U363 (N_363,In_164,In_2442);
nor U364 (N_364,In_233,In_1264);
and U365 (N_365,In_2486,N_160);
xor U366 (N_366,In_1132,In_1489);
xnor U367 (N_367,In_1930,In_1809);
nor U368 (N_368,In_1866,In_466);
xnor U369 (N_369,In_1822,N_43);
or U370 (N_370,In_24,In_1863);
nor U371 (N_371,In_1858,In_1339);
nor U372 (N_372,In_2225,In_323);
nor U373 (N_373,In_401,In_978);
or U374 (N_374,In_309,In_106);
xnor U375 (N_375,In_1660,In_1043);
and U376 (N_376,In_2351,In_1724);
nor U377 (N_377,In_1053,In_116);
nand U378 (N_378,In_2088,In_1825);
or U379 (N_379,In_1473,In_953);
nor U380 (N_380,In_196,In_1472);
nand U381 (N_381,In_829,In_2201);
and U382 (N_382,In_687,In_523);
xor U383 (N_383,In_140,In_707);
nor U384 (N_384,In_1431,In_373);
or U385 (N_385,In_2360,In_107);
nand U386 (N_386,In_504,In_586);
or U387 (N_387,In_188,In_1977);
xnor U388 (N_388,In_158,In_1204);
xor U389 (N_389,In_1151,In_879);
nand U390 (N_390,In_669,In_2245);
or U391 (N_391,In_2004,In_343);
nand U392 (N_392,N_105,In_1890);
or U393 (N_393,In_17,In_564);
xor U394 (N_394,In_661,In_1352);
nand U395 (N_395,In_1311,In_2475);
xnor U396 (N_396,In_2316,In_2217);
xor U397 (N_397,In_1156,In_937);
or U398 (N_398,In_2066,In_2156);
or U399 (N_399,In_1867,In_2046);
or U400 (N_400,In_2136,In_966);
xnor U401 (N_401,In_578,In_1497);
nor U402 (N_402,In_891,In_1599);
nand U403 (N_403,In_1191,In_2495);
xor U404 (N_404,N_373,In_209);
or U405 (N_405,In_1840,In_1658);
xor U406 (N_406,N_270,In_2125);
or U407 (N_407,In_1575,In_949);
or U408 (N_408,In_1738,In_536);
or U409 (N_409,In_1808,In_1834);
xor U410 (N_410,In_2378,In_790);
xor U411 (N_411,In_2241,In_861);
and U412 (N_412,In_1398,N_326);
and U413 (N_413,N_348,In_743);
or U414 (N_414,In_864,In_1971);
and U415 (N_415,In_1771,In_1849);
nor U416 (N_416,In_2263,In_855);
and U417 (N_417,In_2134,In_2008);
and U418 (N_418,In_477,In_1457);
nor U419 (N_419,In_1870,In_2448);
or U420 (N_420,N_202,In_1608);
or U421 (N_421,In_569,In_281);
and U422 (N_422,In_871,In_1720);
or U423 (N_423,In_1979,In_2427);
and U424 (N_424,In_1160,In_1723);
and U425 (N_425,In_117,In_380);
nand U426 (N_426,In_1164,In_1741);
xnor U427 (N_427,In_2152,In_719);
xor U428 (N_428,N_395,In_2022);
and U429 (N_429,In_1247,In_1588);
xnor U430 (N_430,N_370,N_264);
and U431 (N_431,In_1793,N_204);
or U432 (N_432,N_261,In_1461);
nor U433 (N_433,In_244,In_454);
nor U434 (N_434,In_2343,N_216);
or U435 (N_435,In_458,In_1983);
xnor U436 (N_436,N_136,In_95);
or U437 (N_437,In_148,In_1717);
xnor U438 (N_438,In_892,In_514);
nand U439 (N_439,In_1616,In_1188);
or U440 (N_440,In_2053,N_168);
nand U441 (N_441,N_154,In_1839);
nand U442 (N_442,In_1243,In_1235);
nand U443 (N_443,N_173,N_333);
nand U444 (N_444,N_170,In_1619);
or U445 (N_445,In_2290,In_2213);
or U446 (N_446,N_14,In_1549);
and U447 (N_447,In_1498,In_1337);
or U448 (N_448,In_758,In_2054);
xnor U449 (N_449,In_1692,In_1641);
or U450 (N_450,In_1468,In_348);
nor U451 (N_451,In_108,In_524);
nor U452 (N_452,In_722,In_1987);
or U453 (N_453,N_245,In_903);
and U454 (N_454,N_65,In_21);
or U455 (N_455,In_74,In_2261);
or U456 (N_456,In_2002,In_195);
and U457 (N_457,In_2133,In_2497);
and U458 (N_458,N_263,In_1656);
xnor U459 (N_459,In_1859,In_20);
xnor U460 (N_460,In_1733,In_50);
or U461 (N_461,In_2349,In_1476);
xnor U462 (N_462,N_294,N_12);
and U463 (N_463,In_2303,In_19);
or U464 (N_464,In_1297,In_2376);
nand U465 (N_465,In_1104,In_1329);
and U466 (N_466,In_934,In_1312);
and U467 (N_467,In_838,In_1848);
and U468 (N_468,In_2412,In_1838);
nand U469 (N_469,In_877,In_293);
and U470 (N_470,In_45,In_2344);
or U471 (N_471,N_292,N_346);
nand U472 (N_472,In_367,In_341);
or U473 (N_473,In_1748,N_80);
nor U474 (N_474,N_23,In_1348);
and U475 (N_475,N_201,In_1155);
nand U476 (N_476,In_435,In_1595);
or U477 (N_477,In_589,In_263);
nor U478 (N_478,In_598,In_1695);
xnor U479 (N_479,In_313,N_24);
nor U480 (N_480,In_2036,N_384);
nor U481 (N_481,N_150,In_418);
nor U482 (N_482,In_1072,In_448);
nor U483 (N_483,In_2186,N_345);
and U484 (N_484,In_1295,In_377);
nand U485 (N_485,N_269,In_427);
and U486 (N_486,In_2323,In_913);
nand U487 (N_487,In_2372,In_2466);
and U488 (N_488,In_2233,In_1615);
and U489 (N_489,N_140,In_347);
xor U490 (N_490,In_379,In_1980);
and U491 (N_491,In_703,In_1906);
nand U492 (N_492,In_1096,In_981);
xor U493 (N_493,In_1026,In_626);
and U494 (N_494,In_1451,In_1985);
nor U495 (N_495,N_375,In_1555);
or U496 (N_496,In_447,N_192);
or U497 (N_497,In_732,In_1798);
nor U498 (N_498,In_2000,In_2037);
or U499 (N_499,In_1913,In_1003);
and U500 (N_500,In_1095,In_1427);
nand U501 (N_501,In_136,In_2388);
nand U502 (N_502,In_771,In_2061);
nand U503 (N_503,In_1198,In_2312);
xor U504 (N_504,In_875,N_385);
xnor U505 (N_505,N_285,In_2115);
nor U506 (N_506,In_1435,In_3);
xnor U507 (N_507,In_525,N_236);
xor U508 (N_508,N_178,In_221);
nand U509 (N_509,N_92,In_2227);
nand U510 (N_510,N_138,In_506);
nand U511 (N_511,N_266,In_1090);
and U512 (N_512,In_305,In_2443);
or U513 (N_513,In_982,In_415);
or U514 (N_514,In_1703,N_76);
nand U515 (N_515,In_912,In_1509);
nand U516 (N_516,In_1803,In_1356);
and U517 (N_517,In_1958,In_172);
nor U518 (N_518,N_276,In_1690);
and U519 (N_519,In_857,In_1526);
nand U520 (N_520,In_335,In_2135);
and U521 (N_521,In_336,In_2332);
nand U522 (N_522,N_34,In_2072);
nor U523 (N_523,N_62,In_1274);
nand U524 (N_524,In_299,In_126);
and U525 (N_525,In_608,N_324);
nor U526 (N_526,In_883,In_1460);
or U527 (N_527,N_313,In_6);
or U528 (N_528,In_290,In_217);
xnor U529 (N_529,In_1947,In_342);
nand U530 (N_530,In_438,In_311);
or U531 (N_531,In_1673,In_511);
xnor U532 (N_532,In_2122,In_2366);
xnor U533 (N_533,N_318,In_120);
xnor U534 (N_534,In_355,In_2346);
and U535 (N_535,In_1442,In_236);
nand U536 (N_536,In_1429,In_1681);
nor U537 (N_537,In_741,In_2256);
and U538 (N_538,In_54,In_1408);
or U539 (N_539,In_1167,N_176);
nor U540 (N_540,In_731,In_1216);
or U541 (N_541,In_1712,In_986);
nand U542 (N_542,In_1504,In_1362);
and U543 (N_543,In_182,In_2469);
and U544 (N_544,In_295,In_1677);
nand U545 (N_545,In_809,N_210);
nand U546 (N_546,N_95,In_888);
nor U547 (N_547,N_277,In_1607);
nand U548 (N_548,In_1675,In_787);
or U549 (N_549,In_1927,N_234);
xnor U550 (N_550,In_1499,N_354);
and U551 (N_551,In_1341,In_332);
nor U552 (N_552,In_1553,In_592);
xnor U553 (N_553,In_480,In_1711);
xor U554 (N_554,In_1462,In_1492);
xor U555 (N_555,In_1981,In_41);
nor U556 (N_556,In_2297,In_1023);
and U557 (N_557,In_836,In_1407);
nor U558 (N_558,In_591,In_898);
nor U559 (N_559,In_695,In_1455);
nand U560 (N_560,In_1051,In_1513);
or U561 (N_561,N_151,In_1812);
nand U562 (N_562,In_1333,In_132);
nor U563 (N_563,In_674,In_2490);
nor U564 (N_564,In_2377,In_2059);
and U565 (N_565,In_729,In_1923);
nor U566 (N_566,In_1369,In_889);
or U567 (N_567,In_1604,In_696);
nor U568 (N_568,In_821,In_2465);
xnor U569 (N_569,In_1769,In_991);
and U570 (N_570,In_1410,In_1236);
xnor U571 (N_571,In_177,In_2093);
xnor U572 (N_572,In_935,In_1287);
nor U573 (N_573,In_1285,In_1574);
and U574 (N_574,In_750,In_2041);
xnor U575 (N_575,In_2164,In_1226);
nor U576 (N_576,In_662,N_380);
or U577 (N_577,In_955,N_171);
xnor U578 (N_578,In_1871,In_1994);
nor U579 (N_579,In_1134,In_1159);
nand U580 (N_580,In_1815,In_127);
and U581 (N_581,In_56,In_518);
nand U582 (N_582,In_2174,In_2268);
nand U583 (N_583,In_1177,N_129);
and U584 (N_584,In_770,In_1344);
and U585 (N_585,In_13,In_660);
nand U586 (N_586,In_2049,In_207);
or U587 (N_587,In_1676,In_1033);
nand U588 (N_588,N_220,In_919);
or U589 (N_589,In_63,In_1213);
xor U590 (N_590,In_1019,In_1190);
and U591 (N_591,In_2300,In_1214);
and U592 (N_592,In_1091,In_411);
xnor U593 (N_593,In_266,In_2034);
or U594 (N_594,In_470,In_337);
nor U595 (N_595,In_951,In_2229);
or U596 (N_596,In_2052,In_1962);
xnor U597 (N_597,In_2352,In_1350);
and U598 (N_598,N_332,In_2258);
nor U599 (N_599,In_464,In_1280);
nand U600 (N_600,In_2472,In_1648);
and U601 (N_601,N_445,N_8);
nand U602 (N_602,N_421,In_2431);
nor U603 (N_603,N_303,In_239);
xor U604 (N_604,N_436,In_1388);
nand U605 (N_605,In_1321,In_948);
xor U606 (N_606,In_1224,In_187);
nor U607 (N_607,In_686,In_990);
nand U608 (N_608,In_2253,In_503);
or U609 (N_609,N_557,N_365);
and U610 (N_610,In_2325,In_1967);
nor U611 (N_611,N_224,In_450);
nand U612 (N_612,N_545,In_1488);
or U613 (N_613,In_267,N_117);
nand U614 (N_614,N_85,In_1857);
xnor U615 (N_615,In_1651,In_2243);
or U616 (N_616,In_832,In_2339);
nand U617 (N_617,In_2067,In_62);
xor U618 (N_618,N_474,N_312);
and U619 (N_619,In_223,In_99);
or U620 (N_620,In_2084,In_708);
nor U621 (N_621,In_793,N_473);
nor U622 (N_622,N_252,In_1922);
nor U623 (N_623,In_1773,In_885);
xor U624 (N_624,In_1921,N_209);
or U625 (N_625,N_334,In_2380);
nand U626 (N_626,In_1477,In_804);
or U627 (N_627,In_1860,In_152);
nor U628 (N_628,N_287,In_2286);
and U629 (N_629,N_451,In_1955);
or U630 (N_630,N_226,In_2159);
or U631 (N_631,N_587,N_141);
and U632 (N_632,N_344,In_2154);
or U633 (N_633,In_43,In_1115);
xnor U634 (N_634,In_1556,In_1573);
xor U635 (N_635,In_1503,In_2416);
nor U636 (N_636,In_1168,In_161);
xor U637 (N_637,In_1603,In_886);
and U638 (N_638,In_1081,N_90);
nor U639 (N_639,In_998,In_451);
nand U640 (N_640,In_1794,In_2015);
xor U641 (N_641,In_1518,In_680);
nor U642 (N_642,In_678,In_218);
or U643 (N_643,In_1758,In_2005);
xnor U644 (N_644,In_1029,N_368);
and U645 (N_645,N_388,N_584);
or U646 (N_646,In_858,In_1624);
xnor U647 (N_647,N_70,N_19);
xnor U648 (N_648,In_245,N_515);
nor U649 (N_649,N_308,In_816);
xor U650 (N_650,N_409,In_77);
or U651 (N_651,In_399,N_288);
nand U652 (N_652,In_1265,In_2114);
nand U653 (N_653,In_1038,In_2364);
nor U654 (N_654,In_2130,In_1713);
or U655 (N_655,In_371,In_1846);
xnor U656 (N_656,N_490,N_530);
and U657 (N_657,N_2,In_2347);
or U658 (N_658,In_2392,In_1523);
nor U659 (N_659,In_80,N_200);
nor U660 (N_660,In_697,In_146);
nand U661 (N_661,In_2285,N_526);
and U662 (N_662,In_1561,N_462);
and U663 (N_663,In_1083,N_48);
or U664 (N_664,In_1127,In_2299);
nor U665 (N_665,In_969,In_580);
nor U666 (N_666,In_496,N_7);
nand U667 (N_667,In_1430,In_1507);
nor U668 (N_668,N_489,In_1018);
and U669 (N_669,In_129,N_400);
nor U670 (N_670,N_243,In_915);
xnor U671 (N_671,In_369,In_2030);
nand U672 (N_672,In_143,In_528);
nand U673 (N_673,N_161,N_282);
nand U674 (N_674,In_1390,In_602);
or U675 (N_675,In_1978,N_21);
nor U676 (N_676,In_736,In_1031);
or U677 (N_677,N_163,In_593);
nand U678 (N_678,N_106,In_251);
or U679 (N_679,In_1172,N_597);
xor U680 (N_680,In_2121,N_228);
nor U681 (N_681,In_2188,In_2340);
nor U682 (N_682,In_65,In_256);
nor U683 (N_683,N_546,N_447);
xnor U684 (N_684,In_1220,N_507);
or U685 (N_685,In_213,In_2304);
or U686 (N_686,In_1324,In_1547);
nor U687 (N_687,N_271,In_1995);
or U688 (N_688,In_1436,In_1027);
or U689 (N_689,In_2020,In_1572);
or U690 (N_690,In_394,In_154);
nand U691 (N_691,In_730,In_856);
xor U692 (N_692,N_390,In_605);
nand U693 (N_693,In_778,N_519);
xnor U694 (N_694,In_1864,In_1120);
or U695 (N_695,In_398,N_69);
xnor U696 (N_696,N_569,In_615);
xor U697 (N_697,N_541,In_709);
xor U698 (N_698,In_2368,N_439);
or U699 (N_699,N_492,N_244);
or U700 (N_700,In_473,In_517);
nor U701 (N_701,In_2277,N_107);
or U702 (N_702,In_434,N_219);
xor U703 (N_703,In_482,In_962);
xor U704 (N_704,In_1005,In_363);
and U705 (N_705,In_765,In_2131);
nand U706 (N_706,In_1606,In_237);
and U707 (N_707,In_690,N_461);
or U708 (N_708,In_1032,In_1117);
nand U709 (N_709,In_258,In_1875);
xor U710 (N_710,In_2064,N_510);
xor U711 (N_711,N_254,N_521);
and U712 (N_712,In_180,In_91);
or U713 (N_713,In_306,In_5);
and U714 (N_714,In_1073,N_379);
or U715 (N_715,In_2181,In_805);
nor U716 (N_716,In_994,In_2451);
nor U717 (N_717,In_1469,In_1505);
and U718 (N_718,In_575,N_460);
nand U719 (N_719,N_181,N_137);
xor U720 (N_720,N_291,In_1757);
nor U721 (N_721,In_959,In_1950);
nand U722 (N_722,In_1813,In_971);
or U723 (N_723,In_1309,N_438);
xor U724 (N_724,N_249,In_643);
nand U725 (N_725,In_2354,In_1992);
nand U726 (N_726,N_306,In_579);
and U727 (N_727,In_2415,In_1304);
and U728 (N_728,In_970,In_2);
and U729 (N_729,N_102,N_112);
nand U730 (N_730,In_1404,N_478);
xor U731 (N_731,In_1045,In_2447);
xor U732 (N_732,In_1862,In_683);
xor U733 (N_733,In_1092,In_1939);
nand U734 (N_734,N_416,In_486);
nand U735 (N_735,N_585,In_1770);
xor U736 (N_736,In_1173,In_1918);
xnor U737 (N_737,In_94,In_82);
xor U738 (N_738,In_1527,In_2218);
nor U739 (N_739,N_212,In_278);
and U740 (N_740,In_2190,In_1823);
nand U741 (N_741,In_452,In_776);
and U742 (N_742,In_121,In_1719);
nor U743 (N_743,In_252,N_470);
or U744 (N_744,In_1438,In_631);
nor U745 (N_745,N_417,In_2273);
nand U746 (N_746,In_1458,In_1932);
nor U747 (N_747,N_52,In_1954);
xor U748 (N_748,In_1642,N_16);
and U749 (N_749,In_1078,In_1891);
nand U750 (N_750,In_250,N_20);
or U751 (N_751,In_512,N_469);
nor U752 (N_752,In_1314,In_322);
or U753 (N_753,In_1439,In_296);
and U754 (N_754,In_2117,N_466);
or U755 (N_755,In_2393,In_2479);
or U756 (N_756,N_128,In_918);
and U757 (N_757,In_1009,N_267);
and U758 (N_758,In_1564,In_1948);
and U759 (N_759,In_1670,In_1011);
nand U760 (N_760,N_402,In_387);
xnor U761 (N_761,In_2199,N_397);
or U762 (N_762,N_401,In_119);
nor U763 (N_763,In_1557,In_2270);
and U764 (N_764,In_509,In_1087);
xor U765 (N_765,In_1296,In_2250);
or U766 (N_766,In_27,In_1316);
nand U767 (N_767,In_64,In_125);
xnor U768 (N_768,In_1935,In_957);
or U769 (N_769,N_471,In_1569);
or U770 (N_770,N_17,In_23);
and U771 (N_771,In_1290,N_15);
and U772 (N_772,In_979,In_1097);
nor U773 (N_773,In_828,In_603);
or U774 (N_774,In_2016,N_423);
xor U775 (N_775,In_1911,In_947);
and U776 (N_776,In_1959,In_475);
nand U777 (N_777,In_1802,In_1887);
nand U778 (N_778,N_273,In_1421);
nor U779 (N_779,N_561,In_677);
or U780 (N_780,In_1767,In_2278);
nor U781 (N_781,In_1730,In_2003);
or U782 (N_782,In_210,N_410);
xnor U783 (N_783,In_123,In_2234);
nor U784 (N_784,In_1259,In_1138);
nor U785 (N_785,N_93,In_16);
or U786 (N_786,In_2328,N_487);
or U787 (N_787,N_22,In_1267);
nand U788 (N_788,In_1686,In_2168);
nand U789 (N_789,In_423,In_1144);
or U790 (N_790,In_226,In_791);
xor U791 (N_791,In_1933,In_440);
and U792 (N_792,In_2308,In_48);
xor U793 (N_793,In_437,N_341);
or U794 (N_794,In_1006,In_2038);
and U795 (N_795,In_1973,In_843);
or U796 (N_796,N_68,In_339);
nand U797 (N_797,In_2224,In_1819);
xnor U798 (N_798,In_2207,N_367);
and U799 (N_799,N_222,In_1542);
nand U800 (N_800,In_139,N_452);
and U801 (N_801,In_2175,In_145);
nand U802 (N_802,In_596,In_2413);
xor U803 (N_803,In_2073,In_1630);
nor U804 (N_804,N_493,In_1638);
nor U805 (N_805,In_2148,N_4);
nand U806 (N_806,In_422,In_1817);
or U807 (N_807,In_2462,In_1510);
nand U808 (N_808,N_735,N_576);
nand U809 (N_809,In_378,In_2240);
and U810 (N_810,In_1184,N_511);
xor U811 (N_811,In_2389,In_494);
and U812 (N_812,N_664,In_2279);
and U813 (N_813,In_1384,In_2428);
and U814 (N_814,In_2086,In_1128);
nor U815 (N_815,In_704,N_768);
and U816 (N_816,In_44,In_421);
and U817 (N_817,In_1187,N_578);
or U818 (N_818,In_706,N_225);
or U819 (N_819,N_672,In_632);
and U820 (N_820,In_1487,In_505);
xor U821 (N_821,In_1800,In_1582);
and U822 (N_822,In_308,In_2107);
nand U823 (N_823,N_311,In_1666);
and U824 (N_824,In_967,N_755);
xnor U825 (N_825,In_1568,N_527);
or U826 (N_826,In_2441,N_337);
xor U827 (N_827,In_356,In_1837);
or U828 (N_828,In_2161,In_2060);
nand U829 (N_829,In_1089,In_1434);
and U830 (N_830,N_330,In_652);
or U831 (N_831,In_30,In_1650);
or U832 (N_832,In_567,N_604);
and U833 (N_833,N_227,In_11);
nor U834 (N_834,N_667,In_474);
nand U835 (N_835,N_459,N_443);
and U836 (N_836,N_61,In_682);
and U837 (N_837,N_383,In_0);
nor U838 (N_838,N_771,N_751);
xnor U839 (N_839,In_1034,In_1736);
and U840 (N_840,In_2146,In_1180);
or U841 (N_841,In_1874,N_30);
nand U842 (N_842,N_538,In_923);
nand U843 (N_843,N_157,In_588);
nor U844 (N_844,N_476,N_31);
xnor U845 (N_845,N_536,In_2436);
or U846 (N_846,In_1124,In_1585);
or U847 (N_847,N_681,N_477);
and U848 (N_848,In_1411,N_339);
nor U849 (N_849,N_610,N_630);
and U850 (N_850,In_2055,In_2317);
and U851 (N_851,N_786,In_807);
nor U852 (N_852,In_762,In_2373);
or U853 (N_853,In_746,In_1251);
nand U854 (N_854,In_52,In_845);
nor U855 (N_855,In_328,In_1965);
or U856 (N_856,In_1559,N_598);
xnor U857 (N_857,N_422,In_1627);
and U858 (N_858,N_734,N_729);
and U859 (N_859,In_2401,N_378);
and U860 (N_860,In_1179,N_320);
xnor U861 (N_861,In_1804,In_630);
nor U862 (N_862,N_305,In_939);
xnor U863 (N_863,N_188,N_432);
or U864 (N_864,In_2399,N_123);
xor U865 (N_865,In_870,In_774);
nor U866 (N_866,In_246,In_2147);
and U867 (N_867,In_357,In_1877);
xnor U868 (N_868,In_1831,In_1021);
nor U869 (N_869,N_634,N_82);
and U870 (N_870,In_1262,N_429);
nand U871 (N_871,In_1908,N_725);
xor U872 (N_872,N_54,In_2092);
xnor U873 (N_873,In_69,N_353);
xnor U874 (N_874,In_97,In_2498);
or U875 (N_875,N_753,In_1998);
or U876 (N_876,In_1753,N_205);
or U877 (N_877,N_374,In_393);
and U878 (N_878,In_1232,N_503);
xor U879 (N_879,N_198,In_2385);
or U880 (N_880,In_255,In_1949);
and U881 (N_881,In_2017,In_2094);
xnor U882 (N_882,In_2402,N_377);
nor U883 (N_883,N_539,In_938);
nor U884 (N_884,N_403,N_325);
nor U885 (N_885,N_791,In_1137);
and U886 (N_886,In_1154,In_1007);
xnor U887 (N_887,In_1336,In_500);
nor U888 (N_888,In_956,N_127);
nand U889 (N_889,In_1317,In_1391);
xnor U890 (N_890,In_492,N_468);
nand U891 (N_891,In_2142,In_1338);
nand U892 (N_892,In_130,In_977);
or U893 (N_893,N_756,N_230);
xor U894 (N_894,In_783,N_758);
or U895 (N_895,N_547,N_535);
nand U896 (N_896,In_640,In_734);
nor U897 (N_897,N_635,In_324);
xnor U898 (N_898,In_222,N_720);
nand U899 (N_899,In_1231,In_1331);
xor U900 (N_900,In_2269,In_1074);
xor U901 (N_901,N_625,N_728);
xor U902 (N_902,N_639,N_185);
or U903 (N_903,In_2184,In_199);
xnor U904 (N_904,N_435,N_571);
or U905 (N_905,In_1620,N_696);
and U906 (N_906,N_120,In_1365);
and U907 (N_907,In_467,In_2183);
and U908 (N_908,In_899,In_723);
nand U909 (N_909,In_351,N_297);
and U910 (N_910,In_1791,In_658);
nor U911 (N_911,N_338,In_849);
and U912 (N_912,In_533,N_238);
nor U913 (N_913,In_2033,In_1566);
nor U914 (N_914,In_2144,In_1655);
and U915 (N_915,In_1199,N_714);
nor U916 (N_916,N_211,N_631);
nand U917 (N_917,N_357,In_1071);
nand U918 (N_918,N_399,N_628);
nor U919 (N_919,N_626,N_441);
xor U920 (N_920,In_2460,N_687);
xnor U921 (N_921,In_763,N_464);
and U922 (N_922,In_1885,N_274);
xor U923 (N_923,In_1206,In_1065);
nand U924 (N_924,In_2381,In_1737);
and U925 (N_925,In_1088,In_1783);
xnor U926 (N_926,In_902,In_493);
or U927 (N_927,In_1636,In_2083);
nand U928 (N_928,In_1485,In_1253);
and U929 (N_929,N_792,N_662);
xnor U930 (N_930,In_1699,In_350);
and U931 (N_931,In_616,N_609);
and U932 (N_932,In_835,N_501);
nand U933 (N_933,In_463,In_1238);
nand U934 (N_934,N_685,In_1143);
nor U935 (N_935,In_1152,In_681);
or U936 (N_936,In_35,In_1313);
or U937 (N_937,In_1563,N_229);
xor U938 (N_938,In_1739,N_300);
and U939 (N_939,In_1082,N_235);
or U940 (N_940,In_1662,In_738);
xnor U941 (N_941,N_789,N_552);
xor U942 (N_942,In_1661,In_767);
or U943 (N_943,N_71,In_1878);
xnor U944 (N_944,In_1189,N_81);
nand U945 (N_945,In_819,In_2112);
and U946 (N_946,In_1667,In_1360);
xor U947 (N_947,N_711,In_1359);
and U948 (N_948,In_1334,N_27);
or U949 (N_949,In_1,In_413);
xnor U950 (N_950,In_1539,In_1372);
xnor U951 (N_951,In_1907,In_1729);
nor U952 (N_952,In_1484,In_1545);
and U953 (N_953,In_676,N_310);
nor U954 (N_954,In_595,In_799);
nor U955 (N_955,In_772,In_1571);
or U956 (N_956,In_796,In_231);
nand U957 (N_957,In_346,N_525);
and U958 (N_958,N_607,In_1389);
nand U959 (N_959,In_171,N_475);
xnor U960 (N_960,In_638,In_1433);
nor U961 (N_961,In_1322,N_376);
nand U962 (N_962,N_94,N_565);
nor U963 (N_963,In_287,N_795);
and U964 (N_964,In_1017,In_2215);
or U965 (N_965,In_2421,N_159);
nor U966 (N_966,N_679,In_519);
xnor U967 (N_967,In_1380,In_552);
or U968 (N_968,N_514,In_376);
nor U969 (N_969,In_374,In_1869);
and U970 (N_970,In_1587,N_158);
and U971 (N_971,In_1024,N_352);
nor U972 (N_972,In_265,N_648);
or U973 (N_973,In_1625,In_980);
and U974 (N_974,In_1508,N_619);
or U975 (N_975,N_573,N_321);
and U976 (N_976,In_118,N_649);
nand U977 (N_977,In_721,In_537);
or U978 (N_978,In_2262,In_1919);
nor U979 (N_979,In_2104,In_1742);
nand U980 (N_980,In_1110,In_896);
xor U981 (N_981,N_796,In_319);
xor U982 (N_982,N_66,In_135);
or U983 (N_983,In_1683,In_479);
nor U984 (N_984,In_412,In_710);
or U985 (N_985,N_559,In_1899);
or U986 (N_986,N_361,In_397);
nand U987 (N_987,In_1643,In_2456);
and U988 (N_988,In_1842,N_207);
xnor U989 (N_989,In_197,In_2319);
or U990 (N_990,In_194,In_1424);
nor U991 (N_991,In_1030,In_1961);
or U992 (N_992,N_671,N_767);
and U993 (N_993,N_437,N_440);
nor U994 (N_994,N_710,In_2153);
nor U995 (N_995,N_750,In_656);
nor U996 (N_996,In_688,N_516);
xnor U997 (N_997,In_1382,In_86);
nand U998 (N_998,In_2111,In_622);
and U999 (N_999,N_433,In_2150);
xnor U1000 (N_1000,N_716,In_2097);
nor U1001 (N_1001,N_355,In_1856);
or U1002 (N_1002,In_2081,N_591);
or U1003 (N_1003,N_988,N_144);
xnor U1004 (N_1004,In_2198,In_795);
nor U1005 (N_1005,In_620,In_260);
and U1006 (N_1006,N_763,N_759);
or U1007 (N_1007,N_363,In_2068);
xnor U1008 (N_1008,In_2496,In_1535);
nand U1009 (N_1009,In_364,In_2009);
and U1010 (N_1010,In_850,N_520);
nor U1011 (N_1011,In_1600,N_299);
nand U1012 (N_1012,N_785,In_316);
xnor U1013 (N_1013,In_487,In_484);
nor U1014 (N_1014,N_971,In_840);
or U1015 (N_1015,N_396,N_994);
nor U1016 (N_1016,In_1299,In_1631);
and U1017 (N_1017,N_83,In_2467);
or U1018 (N_1018,In_532,N_430);
and U1019 (N_1019,In_2169,In_1482);
nor U1020 (N_1020,In_72,In_2455);
nand U1021 (N_1021,In_2124,In_1210);
xor U1022 (N_1022,N_779,N_119);
nor U1023 (N_1023,In_1876,In_1035);
nand U1024 (N_1024,In_253,N_579);
nand U1025 (N_1025,In_1984,In_815);
xnor U1026 (N_1026,N_617,N_739);
nand U1027 (N_1027,N_614,In_170);
xor U1028 (N_1028,In_1441,N_843);
or U1029 (N_1029,N_766,N_703);
and U1030 (N_1030,N_665,N_948);
xor U1031 (N_1031,N_389,N_603);
nor U1032 (N_1032,In_2307,N_816);
and U1033 (N_1033,In_1446,N_688);
xnor U1034 (N_1034,N_424,In_2474);
and U1035 (N_1035,In_2165,N_776);
xnor U1036 (N_1036,N_653,In_2251);
xor U1037 (N_1037,N_772,N_706);
or U1038 (N_1038,In_71,N_543);
nor U1039 (N_1039,In_2167,In_933);
nor U1040 (N_1040,In_402,N_636);
or U1041 (N_1041,In_1059,N_595);
and U1042 (N_1042,In_1534,N_787);
and U1043 (N_1043,In_1691,In_156);
nand U1044 (N_1044,N_985,In_425);
and U1045 (N_1045,In_585,N_512);
nor U1046 (N_1046,In_617,N_821);
xor U1047 (N_1047,In_2284,N_335);
nand U1048 (N_1048,In_1346,In_1002);
nor U1049 (N_1049,In_1064,N_100);
nand U1050 (N_1050,N_442,N_788);
and U1051 (N_1051,N_544,N_661);
or U1052 (N_1052,N_713,N_842);
nand U1053 (N_1053,In_2206,N_97);
or U1054 (N_1054,N_656,N_600);
nor U1055 (N_1055,In_166,N_752);
nand U1056 (N_1056,N_496,N_912);
xnor U1057 (N_1057,In_1780,In_2477);
and U1058 (N_1058,In_974,In_1502);
or U1059 (N_1059,N_472,In_627);
and U1060 (N_1060,In_2071,N_582);
nand U1061 (N_1061,In_1422,In_540);
nor U1062 (N_1062,N_208,N_916);
xnor U1063 (N_1063,N_960,In_190);
nand U1064 (N_1064,In_1697,In_1385);
nand U1065 (N_1065,N_537,In_1302);
and U1066 (N_1066,In_527,N_386);
xor U1067 (N_1067,In_1223,In_769);
or U1068 (N_1068,In_46,In_1944);
or U1069 (N_1069,In_1755,In_2480);
xor U1070 (N_1070,In_1307,N_331);
xor U1071 (N_1071,N_898,In_572);
xor U1072 (N_1072,N_840,In_917);
and U1073 (N_1073,N_193,In_1623);
and U1074 (N_1074,N_701,In_2032);
xnor U1075 (N_1075,In_1036,N_990);
and U1076 (N_1076,In_1123,N_237);
nor U1077 (N_1077,In_941,N_957);
nand U1078 (N_1078,N_939,N_837);
and U1079 (N_1079,In_872,N_406);
and U1080 (N_1080,N_784,N_206);
and U1081 (N_1081,N_563,N_890);
nor U1082 (N_1082,In_2157,N_455);
nand U1083 (N_1083,N_265,In_2166);
or U1084 (N_1084,In_563,In_1640);
nand U1085 (N_1085,In_14,In_1957);
xor U1086 (N_1086,In_1960,N_412);
or U1087 (N_1087,N_709,N_343);
xnor U1088 (N_1088,In_2126,N_580);
nor U1089 (N_1089,In_58,N_947);
nand U1090 (N_1090,In_51,In_1443);
and U1091 (N_1091,In_225,In_79);
nor U1092 (N_1092,In_649,N_949);
and U1093 (N_1093,In_1230,N_824);
nand U1094 (N_1094,In_105,In_1827);
and U1095 (N_1095,N_84,N_859);
nor U1096 (N_1096,N_221,N_302);
nor U1097 (N_1097,In_2464,N_644);
or U1098 (N_1098,N_232,In_1879);
or U1099 (N_1099,N_450,In_55);
nor U1100 (N_1100,In_2417,N_844);
nor U1101 (N_1101,In_636,In_1872);
or U1102 (N_1102,In_1201,In_854);
nand U1103 (N_1103,In_2365,In_2128);
or U1104 (N_1104,In_547,N_913);
and U1105 (N_1105,In_2450,In_460);
nor U1106 (N_1106,In_1357,N_748);
nor U1107 (N_1107,In_2482,In_822);
nor U1108 (N_1108,N_983,In_178);
or U1109 (N_1109,N_504,In_268);
nor U1110 (N_1110,N_964,N_444);
or U1111 (N_1111,N_463,In_958);
nand U1112 (N_1112,In_1905,In_1277);
and U1113 (N_1113,N_765,N_637);
nor U1114 (N_1114,In_577,In_2209);
nor U1115 (N_1115,In_2387,N_855);
nand U1116 (N_1116,In_2327,In_39);
nand U1117 (N_1117,In_768,In_786);
xnor U1118 (N_1118,In_1183,N_131);
or U1119 (N_1119,In_333,In_1076);
xnor U1120 (N_1120,In_516,N_744);
and U1121 (N_1121,In_2182,N_620);
nand U1122 (N_1122,In_352,In_433);
nor U1123 (N_1123,N_246,In_1165);
xor U1124 (N_1124,In_2379,N_611);
nor U1125 (N_1125,N_839,In_1747);
nand U1126 (N_1126,N_899,In_1207);
and U1127 (N_1127,N_599,In_2432);
nand U1128 (N_1128,N_36,In_2228);
and U1129 (N_1129,In_1060,In_1252);
and U1130 (N_1130,N_568,In_205);
and U1131 (N_1131,In_1810,N_927);
nor U1132 (N_1132,In_230,N_831);
xnor U1133 (N_1133,In_1506,N_973);
nand U1134 (N_1134,N_78,N_730);
nand U1135 (N_1135,In_961,In_779);
or U1136 (N_1136,In_1762,N_351);
or U1137 (N_1137,In_1746,In_788);
xnor U1138 (N_1138,In_1496,In_2219);
nor U1139 (N_1139,N_629,N_56);
nor U1140 (N_1140,In_163,N_926);
nor U1141 (N_1141,N_88,N_3);
or U1142 (N_1142,In_565,In_1551);
nor U1143 (N_1143,In_2382,N_799);
nor U1144 (N_1144,In_798,N_956);
and U1145 (N_1145,N_555,In_2192);
or U1146 (N_1146,In_1208,N_862);
xnor U1147 (N_1147,N_359,N_0);
or U1148 (N_1148,In_1511,In_930);
or U1149 (N_1149,N_858,N_28);
nor U1150 (N_1150,In_2044,In_1824);
xnor U1151 (N_1151,N_109,In_1400);
nor U1152 (N_1152,In_449,N_283);
xnor U1153 (N_1153,N_18,In_1843);
and U1154 (N_1154,N_801,In_1610);
nor U1155 (N_1155,In_614,In_526);
nand U1156 (N_1156,N_608,In_59);
xnor U1157 (N_1157,N_372,In_469);
xnor U1158 (N_1158,In_612,In_1416);
and U1159 (N_1159,In_1241,In_498);
or U1160 (N_1160,In_1420,N_651);
nand U1161 (N_1161,N_708,In_2283);
xor U1162 (N_1162,In_179,N_413);
nor U1163 (N_1163,In_1501,N_307);
xnor U1164 (N_1164,N_700,In_1647);
nand U1165 (N_1165,In_2129,In_1841);
or U1166 (N_1166,In_2276,In_2029);
nand U1167 (N_1167,N_114,In_2414);
xor U1168 (N_1168,In_232,In_1565);
nand U1169 (N_1169,N_534,N_669);
nand U1170 (N_1170,N_407,In_2329);
xor U1171 (N_1171,In_444,N_6);
xnor U1172 (N_1172,N_847,N_548);
xnor U1173 (N_1173,In_1991,In_663);
nand U1174 (N_1174,N_645,In_1674);
or U1175 (N_1175,N_73,In_36);
or U1176 (N_1176,In_624,N_747);
nor U1177 (N_1177,In_2208,In_792);
nand U1178 (N_1178,N_732,N_121);
and U1179 (N_1179,In_1066,N_769);
xnor U1180 (N_1180,In_457,N_126);
xor U1181 (N_1181,In_1774,In_943);
xor U1182 (N_1182,N_195,In_2485);
nand U1183 (N_1183,In_2211,N_418);
nor U1184 (N_1184,In_189,In_748);
xor U1185 (N_1185,N_683,N_951);
or U1186 (N_1186,N_258,In_2437);
xor U1187 (N_1187,N_993,N_362);
and U1188 (N_1188,N_624,N_910);
or U1189 (N_1189,N_60,N_113);
or U1190 (N_1190,In_1728,In_1664);
nor U1191 (N_1191,In_481,In_2127);
nor U1192 (N_1192,N_857,N_39);
and U1193 (N_1193,N_911,N_189);
nor U1194 (N_1194,N_593,In_1964);
nand U1195 (N_1195,In_2040,In_2116);
nand U1196 (N_1196,N_482,N_867);
and U1197 (N_1197,N_419,N_909);
or U1198 (N_1198,In_747,N_762);
or U1199 (N_1199,N_53,In_2403);
nor U1200 (N_1200,N_715,N_1099);
nand U1201 (N_1201,In_1378,In_2282);
nor U1202 (N_1202,In_2398,N_1114);
nand U1203 (N_1203,N_1076,In_169);
nand U1204 (N_1204,N_1127,In_1562);
or U1205 (N_1205,N_1179,N_1141);
nand U1206 (N_1206,In_2063,In_2287);
and U1207 (N_1207,N_1185,N_827);
or U1208 (N_1208,N_922,In_1343);
and U1209 (N_1209,In_568,N_1064);
nand U1210 (N_1210,N_533,In_1070);
nor U1211 (N_1211,N_797,In_2386);
and U1212 (N_1212,N_1031,In_269);
nand U1213 (N_1213,N_1164,N_508);
or U1214 (N_1214,N_340,In_60);
nor U1215 (N_1215,In_2252,In_1644);
xnor U1216 (N_1216,In_1694,N_689);
and U1217 (N_1217,In_1054,In_2220);
nand U1218 (N_1218,N_32,In_2330);
xor U1219 (N_1219,In_972,In_1363);
xor U1220 (N_1220,N_945,In_302);
nand U1221 (N_1221,N_284,In_147);
nor U1222 (N_1222,N_690,N_781);
xnor U1223 (N_1223,In_2155,In_1970);
xnor U1224 (N_1224,In_383,In_104);
nor U1225 (N_1225,N_513,N_1125);
or U1226 (N_1226,N_1174,In_1413);
nand U1227 (N_1227,N_1104,In_1039);
and U1228 (N_1228,N_124,N_165);
nor U1229 (N_1229,In_1100,In_1567);
nor U1230 (N_1230,N_815,In_874);
and U1231 (N_1231,In_1732,In_1016);
xnor U1232 (N_1232,N_995,In_2494);
nand U1233 (N_1233,N_794,N_870);
nor U1234 (N_1234,In_698,N_465);
and U1235 (N_1235,In_359,In_219);
xnor U1236 (N_1236,In_1465,N_532);
nor U1237 (N_1237,N_290,In_1129);
xnor U1238 (N_1238,In_2026,N_1196);
or U1239 (N_1239,N_393,In_910);
and U1240 (N_1240,In_87,In_745);
or U1241 (N_1241,In_1537,N_722);
nand U1242 (N_1242,N_1103,In_1255);
nand U1243 (N_1243,In_1094,N_1154);
nor U1244 (N_1244,In_70,In_2488);
and U1245 (N_1245,In_2313,N_55);
nand U1246 (N_1246,In_128,N_968);
nor U1247 (N_1247,In_999,N_1106);
or U1248 (N_1248,In_2137,N_572);
or U1249 (N_1249,N_1181,In_992);
nor U1250 (N_1250,In_718,In_2105);
and U1251 (N_1251,In_1354,N_1015);
nor U1252 (N_1252,N_986,N_1117);
nor U1253 (N_1253,In_1536,In_288);
or U1254 (N_1254,In_749,N_1165);
nor U1255 (N_1255,In_1576,In_1778);
nand U1256 (N_1256,N_642,In_102);
and U1257 (N_1257,In_1085,N_304);
xnor U1258 (N_1258,In_2367,N_731);
xor U1259 (N_1259,In_2259,In_1900);
nand U1260 (N_1260,N_262,N_832);
nand U1261 (N_1261,In_869,N_887);
nand U1262 (N_1262,N_932,N_1017);
nor U1263 (N_1263,N_125,In_1759);
and U1264 (N_1264,N_382,N_1075);
nand U1265 (N_1265,N_349,In_545);
nor U1266 (N_1266,N_1091,In_344);
nand U1267 (N_1267,In_1605,N_239);
xor U1268 (N_1268,In_1010,In_1145);
xor U1269 (N_1269,N_871,In_385);
and U1270 (N_1270,N_41,In_2326);
xnor U1271 (N_1271,N_601,N_872);
or U1272 (N_1272,N_854,In_1633);
nor U1273 (N_1273,In_1062,In_784);
xnor U1274 (N_1274,In_1495,In_2140);
and U1275 (N_1275,N_885,N_1063);
xor U1276 (N_1276,In_1776,In_1990);
and U1277 (N_1277,N_893,N_1011);
or U1278 (N_1278,In_495,N_364);
nor U1279 (N_1279,In_1689,N_849);
and U1280 (N_1280,N_118,In_717);
or U1281 (N_1281,N_657,In_25);
and U1282 (N_1282,N_878,In_584);
or U1283 (N_1283,N_509,N_558);
and U1284 (N_1284,N_398,In_2079);
and U1285 (N_1285,N_967,N_240);
and U1286 (N_1286,In_167,N_805);
nor U1287 (N_1287,In_2396,In_1153);
xor U1288 (N_1288,N_775,In_277);
or U1289 (N_1289,In_15,N_1149);
and U1290 (N_1290,In_414,In_1782);
or U1291 (N_1291,In_141,N_499);
xnor U1292 (N_1292,In_781,N_660);
xor U1293 (N_1293,In_954,In_2180);
nor U1294 (N_1294,In_1952,N_908);
xor U1295 (N_1295,In_468,N_415);
and U1296 (N_1296,In_1688,In_639);
and U1297 (N_1297,N_567,N_1043);
nand U1298 (N_1298,In_895,In_1225);
and U1299 (N_1299,In_2293,In_694);
xnor U1300 (N_1300,N_745,In_806);
or U1301 (N_1301,N_963,N_680);
nor U1302 (N_1302,N_1096,N_1081);
or U1303 (N_1303,N_1172,In_1892);
xnor U1304 (N_1304,In_2445,N_404);
nand U1305 (N_1305,In_395,In_409);
nand U1306 (N_1306,N_1193,N_247);
xnor U1307 (N_1307,N_467,N_1121);
nand U1308 (N_1308,In_2459,In_1716);
or U1309 (N_1309,N_1183,In_521);
nor U1310 (N_1310,N_1086,N_670);
nand U1311 (N_1311,In_2424,N_941);
or U1312 (N_1312,N_860,N_1022);
xnor U1313 (N_1313,In_1044,N_1138);
nand U1314 (N_1314,N_592,In_184);
nor U1315 (N_1315,N_75,N_49);
xor U1316 (N_1316,In_834,N_605);
and U1317 (N_1317,N_655,N_197);
nand U1318 (N_1318,In_396,N_322);
and U1319 (N_1319,In_2271,N_869);
xor U1320 (N_1320,N_1173,In_1898);
or U1321 (N_1321,N_1059,N_977);
or U1322 (N_1322,N_663,In_1928);
or U1323 (N_1323,N_790,N_934);
nand U1324 (N_1324,In_150,N_214);
or U1325 (N_1325,N_1052,N_296);
and U1326 (N_1326,N_740,In_1121);
nand U1327 (N_1327,N_749,In_2483);
nand U1328 (N_1328,N_549,N_1048);
and U1329 (N_1329,In_235,In_570);
and U1330 (N_1330,N_773,N_1078);
and U1331 (N_1331,N_846,N_921);
and U1332 (N_1332,In_1649,N_259);
and U1333 (N_1333,In_2418,In_2336);
nor U1334 (N_1334,In_2139,N_13);
nor U1335 (N_1335,In_1761,N_1194);
or U1336 (N_1336,In_1367,N_806);
nand U1337 (N_1337,N_724,N_281);
nor U1338 (N_1338,In_1531,N_982);
nor U1339 (N_1339,N_336,N_169);
nor U1340 (N_1340,In_441,N_976);
or U1341 (N_1341,N_589,N_901);
and U1342 (N_1342,N_761,In_1525);
nor U1343 (N_1343,In_282,In_1543);
xor U1344 (N_1344,N_1192,In_1792);
nand U1345 (N_1345,N_1197,In_416);
or U1346 (N_1346,N_807,N_251);
nand U1347 (N_1347,In_1195,N_1042);
or U1348 (N_1348,N_1009,In_208);
nor U1349 (N_1349,N_754,In_2223);
or U1350 (N_1350,In_2216,In_960);
nor U1351 (N_1351,N_1016,In_216);
nand U1352 (N_1352,N_943,N_551);
or U1353 (N_1353,N_356,In_968);
nor U1354 (N_1354,In_2045,In_1915);
or U1355 (N_1355,N_978,In_812);
nor U1356 (N_1356,N_1093,In_2353);
nor U1357 (N_1357,N_659,N_256);
or U1358 (N_1358,N_961,N_155);
nand U1359 (N_1359,In_1250,N_638);
and U1360 (N_1360,In_2318,In_1228);
nand U1361 (N_1361,In_68,N_704);
and U1362 (N_1362,N_1045,N_712);
or U1363 (N_1363,In_1004,N_814);
nand U1364 (N_1364,N_879,In_507);
nand U1365 (N_1365,N_851,In_2429);
nand U1366 (N_1366,N_1195,N_575);
or U1367 (N_1367,In_1931,In_618);
nor U1368 (N_1368,In_124,N_707);
nor U1369 (N_1369,In_558,In_1598);
xor U1370 (N_1370,N_612,N_1080);
and U1371 (N_1371,In_1282,In_1614);
or U1372 (N_1372,In_310,N_458);
and U1373 (N_1373,N_590,N_918);
and U1374 (N_1374,In_381,In_1263);
or U1375 (N_1375,N_581,In_270);
or U1376 (N_1376,N_387,In_461);
nand U1377 (N_1377,In_2309,N_783);
nand U1378 (N_1378,In_1829,N_881);
nand U1379 (N_1379,In_2178,N_895);
or U1380 (N_1380,In_1828,In_1914);
nand U1381 (N_1381,In_1041,In_491);
nor U1382 (N_1382,N_992,N_833);
nand U1383 (N_1383,In_1687,N_564);
nand U1384 (N_1384,In_1102,N_64);
and U1385 (N_1385,In_2440,N_272);
xnor U1386 (N_1386,In_2369,N_804);
and U1387 (N_1387,N_1156,In_685);
xor U1388 (N_1388,In_1122,In_932);
xor U1389 (N_1389,N_556,In_2444);
xor U1390 (N_1390,In_193,In_671);
nand U1391 (N_1391,In_2103,N_1163);
xnor U1392 (N_1392,N_652,N_523);
nor U1393 (N_1393,N_1056,N_135);
or U1394 (N_1394,In_241,N_1090);
nor U1395 (N_1395,In_2101,N_485);
nand U1396 (N_1396,In_202,N_1068);
or U1397 (N_1397,N_917,N_866);
nand U1398 (N_1398,N_677,N_162);
nand U1399 (N_1399,In_1063,N_778);
nor U1400 (N_1400,N_142,In_2315);
or U1401 (N_1401,N_823,N_673);
nand U1402 (N_1402,N_329,In_1577);
nor U1403 (N_1403,N_1143,N_698);
and U1404 (N_1404,In_1789,In_1113);
xnor U1405 (N_1405,N_891,N_1280);
nor U1406 (N_1406,In_1801,N_705);
or U1407 (N_1407,N_1111,N_774);
xor U1408 (N_1408,In_2449,In_839);
xnor U1409 (N_1409,N_1242,In_1448);
nor U1410 (N_1410,In_2361,N_1360);
and U1411 (N_1411,N_1014,In_175);
nand U1412 (N_1412,In_1772,N_825);
and U1413 (N_1413,In_365,In_1483);
and U1414 (N_1414,N_1003,N_1237);
or U1415 (N_1415,N_613,In_833);
nor U1416 (N_1416,N_658,In_2087);
nand U1417 (N_1417,In_2119,In_89);
or U1418 (N_1418,N_1115,N_1110);
and U1419 (N_1419,In_2342,In_534);
nor U1420 (N_1420,N_1182,N_89);
xnor U1421 (N_1421,In_1209,N_1211);
and U1422 (N_1422,In_714,In_100);
nand U1423 (N_1423,N_902,N_1279);
nor U1424 (N_1424,In_1405,In_1375);
nand U1425 (N_1425,N_743,N_1293);
nor U1426 (N_1426,N_892,N_1220);
or U1427 (N_1427,N_1051,N_1105);
and U1428 (N_1428,N_1077,N_1155);
xor U1429 (N_1429,N_1199,In_2275);
or U1430 (N_1430,N_1392,N_760);
xnor U1431 (N_1431,N_1036,N_47);
or U1432 (N_1432,N_1302,N_1222);
or U1433 (N_1433,N_279,N_434);
nor U1434 (N_1434,In_548,In_1852);
xnor U1435 (N_1435,In_862,N_1292);
and U1436 (N_1436,In_1529,N_1316);
or U1437 (N_1437,N_877,N_1166);
or U1438 (N_1438,In_1541,In_1079);
and U1439 (N_1439,N_26,In_566);
xnor U1440 (N_1440,In_975,N_1053);
or U1441 (N_1441,In_1432,In_155);
xnor U1442 (N_1442,In_264,In_274);
xnor U1443 (N_1443,N_938,In_2487);
nand U1444 (N_1444,N_484,In_2302);
nor U1445 (N_1445,N_1284,N_448);
xor U1446 (N_1446,In_1463,N_1359);
nand U1447 (N_1447,N_1334,N_199);
nand U1448 (N_1448,In_2163,N_935);
and U1449 (N_1449,In_28,In_1602);
and U1450 (N_1450,N_1132,In_715);
nor U1451 (N_1451,In_276,N_358);
nand U1452 (N_1452,N_640,N_1116);
nor U1453 (N_1453,In_1452,N_1087);
or U1454 (N_1454,In_825,In_1652);
xor U1455 (N_1455,N_116,In_1881);
or U1456 (N_1456,N_1343,N_67);
or U1457 (N_1457,In_2106,N_1073);
nor U1458 (N_1458,N_1210,N_275);
and U1459 (N_1459,N_187,N_633);
and U1460 (N_1460,N_733,In_827);
nor U1461 (N_1461,N_1365,N_215);
and U1462 (N_1462,N_1004,N_1300);
nor U1463 (N_1463,In_382,In_2357);
nor U1464 (N_1464,N_1329,In_1679);
nand U1465 (N_1465,N_742,In_560);
nand U1466 (N_1466,N_1204,N_1285);
xnor U1467 (N_1467,In_8,N_1037);
nand U1468 (N_1468,In_561,N_528);
or U1469 (N_1469,In_1654,In_884);
xor U1470 (N_1470,N_1289,N_1386);
and U1471 (N_1471,N_1295,N_900);
or U1472 (N_1472,In_472,N_1035);
nand U1473 (N_1473,N_1350,N_980);
and U1474 (N_1474,N_622,In_459);
nor U1475 (N_1475,N_480,N_940);
or U1476 (N_1476,N_1061,N_1107);
nand U1477 (N_1477,In_2335,N_1393);
xor U1478 (N_1478,In_1788,In_814);
and U1479 (N_1479,N_323,N_1189);
xnor U1480 (N_1480,N_1349,In_1234);
or U1481 (N_1481,In_1731,N_1123);
nand U1482 (N_1482,In_110,N_1066);
or U1483 (N_1483,N_1338,In_1310);
nor U1484 (N_1484,N_621,N_1023);
nor U1485 (N_1485,N_553,N_813);
nor U1486 (N_1486,N_317,In_1500);
nand U1487 (N_1487,N_518,N_371);
xor U1488 (N_1488,In_1320,In_724);
xnor U1489 (N_1489,N_1232,N_868);
xnor U1490 (N_1490,N_1062,In_735);
or U1491 (N_1491,N_641,N_882);
nand U1492 (N_1492,N_1335,In_1396);
nand U1493 (N_1493,N_1323,N_1005);
or U1494 (N_1494,N_72,N_1021);
nand U1495 (N_1495,In_1833,N_172);
nand U1496 (N_1496,N_820,In_647);
and U1497 (N_1497,N_1018,N_1264);
nor U1498 (N_1498,N_1221,In_1893);
xor U1499 (N_1499,N_920,In_1196);
and U1500 (N_1500,N_1235,N_856);
nand U1501 (N_1501,N_1092,N_817);
nand U1502 (N_1502,In_2356,N_1270);
nand U1503 (N_1503,In_863,In_243);
and U1504 (N_1504,N_1345,In_29);
and U1505 (N_1505,N_194,N_1124);
xor U1506 (N_1506,N_1147,N_979);
xor U1507 (N_1507,N_491,N_1382);
nor U1508 (N_1508,In_257,N_616);
or U1509 (N_1509,N_812,N_1207);
nand U1510 (N_1510,N_1158,N_1347);
nor U1511 (N_1511,N_1344,In_900);
and U1512 (N_1512,N_1160,N_888);
and U1513 (N_1513,N_666,In_699);
or U1514 (N_1514,N_164,In_744);
or U1515 (N_1515,In_2056,In_442);
or U1516 (N_1516,N_826,In_546);
or U1517 (N_1517,In_272,In_2384);
nand U1518 (N_1518,N_479,N_1340);
and U1519 (N_1519,N_1304,N_524);
xnor U1520 (N_1520,N_1102,In_2247);
nor U1521 (N_1521,In_1286,N_446);
nor U1522 (N_1522,N_1231,In_407);
nor U1523 (N_1523,N_566,In_1705);
nand U1524 (N_1524,In_1558,In_1580);
nor U1525 (N_1525,N_1381,N_1252);
xnor U1526 (N_1526,In_1996,In_985);
and U1527 (N_1527,In_609,N_782);
nor U1528 (N_1528,In_880,N_1161);
nor U1529 (N_1529,In_1383,N_506);
nor U1530 (N_1530,N_676,N_1112);
nand U1531 (N_1531,N_495,In_897);
and U1532 (N_1532,N_1256,In_700);
and U1533 (N_1533,N_74,In_2231);
xnor U1534 (N_1534,N_391,N_1187);
or U1535 (N_1535,In_1133,N_1008);
and U1536 (N_1536,N_830,N_965);
xor U1537 (N_1537,In_2075,N_1229);
nand U1538 (N_1538,In_499,N_1305);
or U1539 (N_1539,N_1390,N_1299);
or U1540 (N_1540,N_1362,N_1303);
nor U1541 (N_1541,N_904,N_570);
nand U1542 (N_1542,N_1396,N_1040);
or U1543 (N_1543,In_1768,N_1169);
and U1544 (N_1544,N_906,N_1227);
nor U1545 (N_1545,N_803,In_2434);
nand U1546 (N_1546,N_1,N_1247);
or U1547 (N_1547,N_1170,In_1284);
and U1548 (N_1548,N_1258,N_408);
nand U1549 (N_1549,N_502,In_314);
and U1550 (N_1550,N_1209,N_241);
nor U1551 (N_1551,N_819,N_231);
xor U1552 (N_1552,In_803,N_1376);
xor U1553 (N_1553,N_1157,In_1763);
nor U1554 (N_1554,N_577,In_1760);
and U1555 (N_1555,N_1244,In_1751);
or U1556 (N_1556,N_1339,In_446);
xor U1557 (N_1557,N_1034,N_1233);
nor U1558 (N_1558,N_1355,In_1830);
and U1559 (N_1559,N_924,N_738);
xnor U1560 (N_1560,N_695,N_1089);
xnor U1561 (N_1561,In_1750,N_684);
nand U1562 (N_1562,N_1135,In_1106);
nor U1563 (N_1563,In_1358,N_809);
and U1564 (N_1564,N_87,N_697);
or U1565 (N_1565,In_366,N_987);
and U1566 (N_1566,In_1734,N_1375);
and U1567 (N_1567,N_876,In_1806);
xor U1568 (N_1568,N_991,In_2363);
or U1569 (N_1569,N_650,N_315);
or U1570 (N_1570,N_864,In_1883);
xnor U1571 (N_1571,In_1402,N_946);
or U1572 (N_1572,N_1322,In_911);
nor U1573 (N_1573,N_1281,In_2098);
and U1574 (N_1574,N_289,N_996);
xnor U1575 (N_1575,N_694,N_770);
nand U1576 (N_1576,N_841,In_1330);
and U1577 (N_1577,N_147,N_1071);
or U1578 (N_1578,N_1241,N_1083);
xor U1579 (N_1579,In_2222,In_1632);
or U1580 (N_1580,N_1228,In_1055);
nand U1581 (N_1581,In_81,N_360);
nor U1582 (N_1582,N_1041,N_915);
xor U1583 (N_1583,In_759,N_1245);
and U1584 (N_1584,N_223,N_981);
and U1585 (N_1585,N_540,In_37);
or U1586 (N_1586,In_1449,In_1901);
and U1587 (N_1587,N_44,In_1657);
nor U1588 (N_1588,N_1319,N_1290);
and U1589 (N_1589,N_560,N_298);
and U1590 (N_1590,N_838,In_1466);
nor U1591 (N_1591,N_835,N_975);
nand U1592 (N_1592,N_1318,N_350);
xor U1593 (N_1593,N_1332,N_999);
and U1594 (N_1594,In_2108,N_1159);
and U1595 (N_1595,N_1200,N_606);
nor U1596 (N_1596,N_1101,N_966);
and U1597 (N_1597,In_285,N_1088);
nor U1598 (N_1598,N_405,N_1108);
nor U1599 (N_1599,N_802,N_798);
xnor U1600 (N_1600,N_1460,In_1306);
and U1601 (N_1601,N_746,N_517);
xor U1602 (N_1602,In_392,In_901);
and U1603 (N_1603,In_665,In_659);
or U1604 (N_1604,In_2239,In_443);
xor U1605 (N_1605,N_1033,In_554);
or U1606 (N_1606,N_1129,In_2110);
xor U1607 (N_1607,In_2249,In_1579);
xnor U1608 (N_1608,N_852,N_1487);
and U1609 (N_1609,N_1324,N_1405);
and U1610 (N_1610,N_1351,N_414);
or U1611 (N_1611,In_2314,N_1213);
xnor U1612 (N_1612,N_453,N_1069);
nand U1613 (N_1613,N_691,N_741);
nor U1614 (N_1614,In_1008,In_1835);
xor U1615 (N_1615,In_1904,N_1579);
nor U1616 (N_1616,N_1180,In_1186);
nor U1617 (N_1617,In_1902,N_1561);
nor U1618 (N_1618,N_1341,In_1920);
nor U1619 (N_1619,In_2006,N_1388);
nand U1620 (N_1620,In_1395,In_1581);
nand U1621 (N_1621,In_403,N_692);
nor U1622 (N_1622,N_1568,N_1145);
nand U1623 (N_1623,N_278,N_1348);
or U1624 (N_1624,In_1379,In_1141);
nor U1625 (N_1625,In_2295,N_529);
xor U1626 (N_1626,N_1070,N_280);
and U1627 (N_1627,N_944,In_2195);
or U1628 (N_1628,N_1234,N_1587);
nand U1629 (N_1629,N_1067,In_637);
xor U1630 (N_1630,N_1595,In_138);
or U1631 (N_1631,N_1515,N_1248);
nor U1632 (N_1632,N_886,N_1424);
and U1633 (N_1633,N_1269,N_1459);
and U1634 (N_1634,N_1511,In_1997);
or U1635 (N_1635,N_42,N_1468);
xnor U1636 (N_1636,In_1342,N_143);
nand U1637 (N_1637,In_1328,N_1380);
xnor U1638 (N_1638,In_818,N_1488);
and U1639 (N_1639,N_449,N_1261);
nor U1640 (N_1640,N_1588,In_1240);
nor U1641 (N_1641,In_1628,In_2438);
nand U1642 (N_1642,In_553,In_429);
and U1643 (N_1643,N_33,N_1584);
or U1644 (N_1644,N_1259,N_998);
nor U1645 (N_1645,N_108,N_1030);
and U1646 (N_1646,N_1591,N_1451);
xnor U1647 (N_1647,N_845,In_1873);
and U1648 (N_1648,N_896,N_1581);
nand U1649 (N_1649,N_1342,N_301);
nor U1650 (N_1650,N_903,In_2082);
nand U1651 (N_1651,N_955,In_1820);
and U1652 (N_1652,In_2410,In_2289);
or U1653 (N_1653,N_1486,In_859);
or U1654 (N_1654,N_1217,N_1208);
nand U1655 (N_1655,N_1567,In_2031);
nand U1656 (N_1656,In_810,N_1462);
nor U1657 (N_1657,In_2221,N_1437);
nand U1658 (N_1658,In_53,N_800);
nor U1659 (N_1659,In_456,N_952);
and U1660 (N_1660,N_1007,N_255);
xor U1661 (N_1661,In_259,N_1407);
and U1662 (N_1662,In_983,In_914);
nand U1663 (N_1663,N_1253,N_250);
nor U1664 (N_1664,In_1478,N_1573);
or U1665 (N_1665,N_1570,N_1397);
xor U1666 (N_1666,N_1309,In_1698);
nand U1667 (N_1667,N_1024,N_1466);
and U1668 (N_1668,N_1128,In_1546);
xor U1669 (N_1669,N_1419,N_1496);
or U1670 (N_1670,N_1139,N_213);
or U1671 (N_1671,In_1219,N_1406);
or U1672 (N_1672,In_848,In_543);
or U1673 (N_1673,N_1225,In_1107);
or U1674 (N_1674,N_836,N_853);
or U1675 (N_1675,In_1744,N_488);
and U1676 (N_1676,N_1119,N_1593);
or U1677 (N_1677,In_2109,N_1134);
and U1678 (N_1678,In_1481,In_1254);
and U1679 (N_1679,In_1494,N_1074);
nor U1680 (N_1680,N_1491,N_1449);
or U1681 (N_1681,In_1609,N_1448);
or U1682 (N_1682,N_483,In_149);
nand U1683 (N_1683,In_2238,N_486);
and U1684 (N_1684,In_2463,In_338);
nand U1685 (N_1685,N_1524,N_1500);
nand U1686 (N_1686,N_1485,N_1477);
nand U1687 (N_1687,N_1465,In_944);
xor U1688 (N_1688,N_1438,N_719);
nor U1689 (N_1689,N_1404,N_1391);
and U1690 (N_1690,N_233,N_1427);
and U1691 (N_1691,N_1576,In_760);
or U1692 (N_1692,N_1368,N_1379);
or U1693 (N_1693,N_929,N_1373);
and U1694 (N_1694,N_1522,N_153);
or U1695 (N_1695,N_183,In_597);
nand U1696 (N_1696,In_675,In_1203);
nand U1697 (N_1697,N_1494,N_1146);
xor U1698 (N_1698,N_1513,In_1260);
nor U1699 (N_1699,In_1283,N_1095);
and U1700 (N_1700,N_627,N_1317);
nand U1701 (N_1701,In_1895,In_1754);
nor U1702 (N_1702,N_1554,N_257);
xor U1703 (N_1703,N_248,In_315);
nor U1704 (N_1704,N_1471,N_780);
xor U1705 (N_1705,N_931,In_162);
nand U1706 (N_1706,In_101,N_1403);
xnor U1707 (N_1707,N_1493,N_588);
nor U1708 (N_1708,N_1444,N_1268);
nand U1709 (N_1709,N_562,N_1428);
and U1710 (N_1710,N_457,N_1599);
or U1711 (N_1711,N_1336,In_201);
nor U1712 (N_1712,In_508,In_2433);
nand U1713 (N_1713,In_151,In_183);
and U1714 (N_1714,N_1226,N_1238);
nand U1715 (N_1715,N_632,N_1236);
nand U1716 (N_1716,N_1519,N_1473);
xor U1717 (N_1717,N_1333,N_1387);
nand U1718 (N_1718,N_1202,N_425);
nand U1719 (N_1719,In_2321,In_115);
or U1720 (N_1720,N_1130,In_1406);
or U1721 (N_1721,N_1505,N_1306);
nor U1722 (N_1722,N_1489,In_1080);
nand U1723 (N_1723,N_1543,In_1147);
nand U1724 (N_1724,In_2320,N_1520);
nor U1725 (N_1725,N_850,N_953);
or U1726 (N_1726,N_1480,N_427);
nand U1727 (N_1727,In_2409,N_1058);
nand U1728 (N_1728,N_454,N_1418);
xnor U1729 (N_1729,N_1508,N_1498);
and U1730 (N_1730,N_1082,N_1378);
xnor U1731 (N_1731,N_874,N_1298);
nand U1732 (N_1732,In_689,N_1562);
nor U1733 (N_1733,N_1408,N_1133);
nand U1734 (N_1734,N_905,In_2426);
and U1735 (N_1735,N_1212,N_1100);
xnor U1736 (N_1736,In_1098,N_481);
nand U1737 (N_1737,N_721,In_692);
xor U1738 (N_1738,In_1702,N_1510);
nor U1739 (N_1739,In_2305,In_2204);
or U1740 (N_1740,In_142,N_1286);
or U1741 (N_1741,N_1367,N_668);
nand U1742 (N_1742,N_1412,N_328);
and U1743 (N_1743,N_1525,In_326);
nand U1744 (N_1744,N_1144,N_829);
nand U1745 (N_1745,N_1594,N_1541);
and U1746 (N_1746,N_777,N_293);
xor U1747 (N_1747,N_505,N_1422);
xnor U1748 (N_1748,N_594,N_1571);
or U1749 (N_1749,N_191,N_186);
nor U1750 (N_1750,N_1538,N_1283);
nand U1751 (N_1751,In_1693,N_1553);
nor U1752 (N_1752,N_818,In_2267);
or U1753 (N_1753,N_1126,N_1085);
nand U1754 (N_1754,In_1818,N_1531);
nand U1755 (N_1755,N_1527,In_176);
and U1756 (N_1756,In_192,N_1416);
nor U1757 (N_1757,N_327,N_146);
nand U1758 (N_1758,In_204,N_1363);
and U1759 (N_1759,N_1190,In_808);
and U1760 (N_1760,In_2457,In_2390);
nand U1761 (N_1761,N_1297,N_554);
xor U1762 (N_1762,N_1440,N_1084);
xor U1763 (N_1763,In_1233,In_1929);
or U1764 (N_1764,In_1786,In_2471);
nor U1765 (N_1765,N_431,N_933);
nand U1766 (N_1766,N_1148,N_1389);
xor U1767 (N_1767,In_2089,In_1594);
xnor U1768 (N_1768,In_789,In_2151);
or U1769 (N_1769,N_1557,N_1507);
or U1770 (N_1770,N_1575,N_1203);
nand U1771 (N_1771,N_1267,N_1002);
xnor U1772 (N_1772,N_1251,In_1454);
xor U1773 (N_1773,In_1936,N_699);
and U1774 (N_1774,N_808,In_1897);
and U1775 (N_1775,N_997,N_1540);
nor U1776 (N_1776,In_1001,N_1530);
or U1777 (N_1777,N_1120,N_880);
or U1778 (N_1778,In_462,N_531);
or U1779 (N_1779,N_1239,N_623);
and U1780 (N_1780,In_587,N_1255);
and U1781 (N_1781,N_1257,In_26);
nand U1782 (N_1782,In_2338,N_1533);
or U1783 (N_1783,In_1289,In_1704);
nand U1784 (N_1784,N_1046,N_950);
nand U1785 (N_1785,In_1440,N_522);
nor U1786 (N_1786,N_1219,N_217);
nor U1787 (N_1787,N_764,N_1361);
or U1788 (N_1788,N_1596,N_1354);
or U1789 (N_1789,N_1331,N_1597);
nand U1790 (N_1790,N_1314,In_1345);
or U1791 (N_1791,N_494,In_9);
or U1792 (N_1792,In_1634,N_1327);
xnor U1793 (N_1793,N_1564,In_1266);
and U1794 (N_1794,N_1495,In_2489);
xor U1795 (N_1795,In_513,In_1589);
and U1796 (N_1796,N_420,N_1469);
or U1797 (N_1797,In_1409,In_1714);
or U1798 (N_1798,In_1428,N_1434);
and U1799 (N_1799,In_1272,N_1463);
xor U1800 (N_1800,N_1243,In_1397);
or U1801 (N_1801,N_1028,N_1682);
or U1802 (N_1802,N_1788,In_2337);
xnor U1803 (N_1803,N_1660,N_1565);
and U1804 (N_1804,N_1246,In_134);
nand U1805 (N_1805,N_1750,N_1600);
and U1806 (N_1806,N_1723,N_793);
or U1807 (N_1807,N_1551,In_488);
xnor U1808 (N_1808,N_51,N_1746);
xor U1809 (N_1809,In_2419,N_1577);
and U1810 (N_1810,In_497,N_426);
nand U1811 (N_1811,In_882,N_1648);
or U1812 (N_1812,In_354,N_1328);
nor U1813 (N_1813,N_1136,N_1415);
and U1814 (N_1814,N_1006,N_1782);
or U1815 (N_1815,N_1206,N_411);
nor U1816 (N_1816,N_394,N_1622);
and U1817 (N_1817,N_1372,In_2039);
xnor U1818 (N_1818,N_1686,N_1250);
nor U1819 (N_1819,N_675,N_1697);
or U1820 (N_1820,In_2458,N_1649);
and U1821 (N_1821,In_904,N_1693);
nor U1822 (N_1822,N_1443,N_1502);
or U1823 (N_1823,In_1013,N_1094);
and U1824 (N_1824,N_702,N_1162);
nor U1825 (N_1825,N_1675,N_1775);
or U1826 (N_1826,N_1188,N_1751);
xnor U1827 (N_1827,N_1658,N_1400);
or U1828 (N_1828,N_1696,N_1714);
and U1829 (N_1829,N_1641,N_1065);
or U1830 (N_1830,N_1484,N_268);
or U1831 (N_1831,N_1274,N_1249);
and U1832 (N_1832,N_1254,N_1504);
and U1833 (N_1833,N_1497,N_1445);
nor U1834 (N_1834,N_1635,In_1844);
and U1835 (N_1835,In_1052,N_1626);
nand U1836 (N_1836,N_1785,N_1770);
nand U1837 (N_1837,N_1296,N_1547);
or U1838 (N_1838,N_1650,In_234);
xor U1839 (N_1839,N_1178,N_574);
or U1840 (N_1840,N_1109,In_1258);
nand U1841 (N_1841,N_428,N_1621);
or U1842 (N_1842,N_1759,N_1032);
or U1843 (N_1843,In_666,N_1262);
or U1844 (N_1844,N_1442,N_1783);
or U1845 (N_1845,In_1347,N_1688);
nor U1846 (N_1846,N_1205,N_37);
or U1847 (N_1847,N_1768,N_1457);
or U1848 (N_1848,N_1453,In_1956);
or U1849 (N_1849,N_1464,N_1433);
or U1850 (N_1850,N_1754,In_1811);
nor U1851 (N_1851,In_2080,In_2058);
nand U1852 (N_1852,In_1148,N_1312);
nor U1853 (N_1853,In_455,N_1287);
nor U1854 (N_1854,N_1214,N_98);
nor U1855 (N_1855,N_1215,N_1690);
nor U1856 (N_1856,N_1369,N_1608);
nor U1857 (N_1857,N_1447,In_2470);
or U1858 (N_1858,In_2070,N_1478);
or U1859 (N_1859,In_1049,N_811);
or U1860 (N_1860,In_1108,N_1798);
nor U1861 (N_1861,N_1748,In_2196);
and U1862 (N_1862,N_810,N_928);
and U1863 (N_1863,N_1607,In_2264);
and U1864 (N_1864,N_693,N_1590);
nor U1865 (N_1865,N_1047,N_1401);
and U1866 (N_1866,N_1580,In_751);
nor U1867 (N_1867,N_1614,N_392);
xor U1868 (N_1868,In_1663,N_1727);
nor U1869 (N_1869,In_181,In_1142);
xor U1870 (N_1870,In_628,N_1606);
nand U1871 (N_1871,N_1644,N_1153);
or U1872 (N_1872,N_319,N_1672);
and U1873 (N_1873,In_539,N_1698);
xor U1874 (N_1874,N_1402,N_1534);
xnor U1875 (N_1875,N_1725,N_96);
or U1876 (N_1876,N_1628,N_1744);
xnor U1877 (N_1877,N_1712,N_1454);
nand U1878 (N_1878,N_1001,N_602);
nand U1879 (N_1879,N_1772,In_1696);
or U1880 (N_1880,N_1201,In_2334);
xor U1881 (N_1881,N_1734,N_1479);
and U1882 (N_1882,In_1659,N_1038);
xnor U1883 (N_1883,N_1481,N_497);
nor U1884 (N_1884,N_1313,N_1055);
nor U1885 (N_1885,N_1532,N_897);
nand U1886 (N_1886,N_1586,N_1787);
nor U1887 (N_1887,N_865,N_1634);
or U1888 (N_1888,N_1019,N_1223);
or U1889 (N_1889,N_1681,N_618);
and U1890 (N_1890,N_1475,In_331);
and U1891 (N_1891,In_2172,N_1394);
or U1892 (N_1892,N_1556,N_1630);
nor U1893 (N_1893,N_1411,N_46);
or U1894 (N_1894,N_1265,In_2074);
nand U1895 (N_1895,N_1781,In_1752);
or U1896 (N_1896,In_574,N_286);
and U1897 (N_1897,N_1760,In_1937);
and U1898 (N_1898,N_1715,N_1240);
xor U1899 (N_1899,N_1456,N_757);
nor U1900 (N_1900,N_1057,N_1724);
and U1901 (N_1901,N_1773,N_1079);
nand U1902 (N_1902,In_1710,N_1618);
and U1903 (N_1903,In_78,N_1692);
nand U1904 (N_1904,N_1545,N_1769);
xnor U1905 (N_1905,N_1663,N_1535);
nand U1906 (N_1906,N_1779,N_1151);
nor U1907 (N_1907,N_1582,N_1755);
or U1908 (N_1908,N_1054,N_1701);
and U1909 (N_1909,N_1012,N_1358);
or U1910 (N_1910,N_1273,N_586);
and U1911 (N_1911,In_2024,N_1000);
or U1912 (N_1912,N_366,In_2397);
xnor U1913 (N_1913,In_1093,N_1492);
xor U1914 (N_1914,N_1027,N_1414);
and U1915 (N_1915,N_1604,N_1677);
or U1916 (N_1916,N_1730,N_1738);
or U1917 (N_1917,N_972,N_1664);
or U1918 (N_1918,N_1429,N_1652);
and U1919 (N_1919,N_1446,N_1620);
and U1920 (N_1920,In_684,N_253);
or U1921 (N_1921,N_1421,N_1684);
xnor U1922 (N_1922,In_1934,N_894);
nand U1923 (N_1923,N_1320,N_1177);
nand U1924 (N_1924,In_1381,In_483);
nor U1925 (N_1925,N_1757,N_1683);
and U1926 (N_1926,N_1645,N_962);
nor U1927 (N_1927,In_753,N_1516);
nor U1928 (N_1928,N_1559,In_1645);
nor U1929 (N_1929,In_1775,N_1611);
nor U1930 (N_1930,In_1515,In_733);
nor U1931 (N_1931,N_152,N_1731);
or U1932 (N_1932,N_1741,N_1585);
or U1933 (N_1933,N_1653,N_1514);
nand U1934 (N_1934,N_1722,N_727);
or U1935 (N_1935,In_1903,N_1137);
nor U1936 (N_1936,N_1602,N_678);
or U1937 (N_1937,N_1631,N_1609);
nand U1938 (N_1938,N_1616,N_1353);
and U1939 (N_1939,N_1025,In_2050);
and U1940 (N_1940,In_1423,N_1168);
and U1941 (N_1941,N_937,N_542);
nor U1942 (N_1942,N_347,In_391);
nand U1943 (N_1943,N_1745,In_1942);
xnor U1944 (N_1944,N_1311,N_1713);
or U1945 (N_1945,N_1666,In_623);
xnor U1946 (N_1946,N_1558,N_1795);
nand U1947 (N_1947,In_1136,N_1572);
or U1948 (N_1948,N_1771,In_672);
and U1949 (N_1949,N_1122,N_1689);
nor U1950 (N_1950,N_1420,N_1776);
nor U1951 (N_1951,N_1700,N_1385);
nand U1952 (N_1952,N_177,N_1321);
or U1953 (N_1953,N_1762,N_1710);
nor U1954 (N_1954,N_1704,N_1529);
xor U1955 (N_1955,N_1374,N_1499);
or U1956 (N_1956,In_358,N_1753);
nand U1957 (N_1957,N_884,N_1799);
and U1958 (N_1958,N_1426,N_1797);
or U1959 (N_1959,N_1482,In_2013);
nand U1960 (N_1960,N_1560,N_1509);
nor U1961 (N_1961,In_2404,N_1764);
or U1962 (N_1962,N_369,N_1013);
xnor U1963 (N_1963,N_583,N_959);
nor U1964 (N_1964,In_1105,N_1439);
nand U1965 (N_1965,N_1703,N_1060);
nand U1966 (N_1966,N_936,In_2491);
nor U1967 (N_1967,N_717,N_1739);
xnor U1968 (N_1968,N_1260,N_1694);
nand U1969 (N_1969,N_1625,In_846);
and U1970 (N_1970,N_889,N_1330);
nand U1971 (N_1971,N_1566,In_1836);
and U1972 (N_1972,N_1702,In_1269);
and U1973 (N_1973,N_1517,N_615);
or U1974 (N_1974,In_47,N_1536);
nor U1975 (N_1975,N_1230,N_1638);
nor U1976 (N_1976,In_1227,In_1722);
nand U1977 (N_1977,N_1679,N_863);
and U1978 (N_1978,In_1373,N_550);
and U1979 (N_1979,N_1337,N_1578);
nor U1980 (N_1980,N_1432,In_186);
nor U1981 (N_1981,N_196,N_1659);
xnor U1982 (N_1982,N_1673,In_2461);
nand U1983 (N_1983,In_329,N_942);
xor U1984 (N_1984,In_713,N_1733);
nand U1985 (N_1985,N_1461,N_1793);
and U1986 (N_1986,N_1266,N_1026);
or U1987 (N_1987,In_1399,N_1118);
nand U1988 (N_1988,In_1394,N_1352);
xnor U1989 (N_1989,N_1191,N_1646);
nand U1990 (N_1990,N_86,In_32);
nor U1991 (N_1991,In_294,N_1624);
nor U1992 (N_1992,N_1550,In_389);
nand U1993 (N_1993,N_1637,N_1728);
xnor U1994 (N_1994,N_1669,N_1472);
nand U1995 (N_1995,N_58,N_218);
nand U1996 (N_1996,In_556,N_1467);
nor U1997 (N_1997,N_736,N_1470);
or U1998 (N_1998,N_1356,N_1794);
nor U1999 (N_1999,N_1544,N_1647);
and U2000 (N_2000,N_1810,N_1841);
xor U2001 (N_2001,In_248,N_1676);
nor U2002 (N_2002,N_1989,N_1828);
and U2003 (N_2003,In_75,N_1357);
nor U2004 (N_2004,N_1831,N_1097);
or U2005 (N_2005,In_2255,N_1603);
and U2006 (N_2006,N_1537,N_1718);
or U2007 (N_2007,N_1435,N_1417);
xnor U2008 (N_2008,N_1833,In_2010);
nand U2009 (N_2009,N_822,N_1506);
nor U2010 (N_2010,N_1835,N_1996);
nor U2011 (N_2011,In_317,N_1997);
xnor U2012 (N_2012,N_1827,N_1784);
and U2013 (N_2013,N_861,N_1821);
or U2014 (N_2014,N_1820,N_1049);
xnor U2015 (N_2015,N_1632,N_1801);
nor U2016 (N_2016,N_737,N_1263);
or U2017 (N_2017,N_1546,N_1623);
nor U2018 (N_2018,N_1490,In_2177);
and U2019 (N_2019,N_1992,N_1869);
nor U2020 (N_2020,N_1512,N_1911);
and U2021 (N_2021,N_1592,N_1927);
and U2022 (N_2022,N_1924,N_1526);
or U2023 (N_2023,In_2237,N_1474);
or U2024 (N_2024,N_1789,N_1371);
nand U2025 (N_2025,N_1855,N_1982);
and U2026 (N_2026,N_834,N_1098);
nor U2027 (N_2027,N_1922,N_1583);
xor U2028 (N_2028,N_1131,N_295);
nand U2029 (N_2029,N_1892,N_1847);
nand U2030 (N_2030,N_1929,N_1796);
or U2031 (N_2031,In_1475,N_1802);
nor U2032 (N_2032,N_309,N_1747);
nand U2033 (N_2033,N_1807,In_1684);
xnor U2034 (N_2034,N_1072,N_1955);
xor U2035 (N_2035,N_1627,N_1961);
and U2036 (N_2036,N_1655,N_1990);
and U2037 (N_2037,N_1729,N_1716);
and U2038 (N_2038,N_1930,N_1995);
nor U2039 (N_2039,N_1778,N_1891);
and U2040 (N_2040,N_1708,N_1914);
and U2041 (N_2041,In_1471,N_1978);
and U2042 (N_2042,N_1601,N_1843);
nor U2043 (N_2043,N_1410,N_1503);
xnor U2044 (N_2044,N_1431,In_1040);
xor U2045 (N_2045,N_1822,N_1938);
or U2046 (N_2046,N_1605,N_1947);
nand U2047 (N_2047,N_1680,N_1574);
and U2048 (N_2048,N_1931,N_1935);
and U2049 (N_2049,N_1780,N_1839);
or U2050 (N_2050,N_1423,N_1845);
nor U2051 (N_2051,In_228,N_1176);
or U2052 (N_2052,N_1804,N_1920);
nor U2053 (N_2053,N_1736,N_1792);
xor U2054 (N_2054,In_1377,N_875);
nor U2055 (N_2055,N_1950,N_1050);
and U2056 (N_2056,N_35,N_974);
and U2057 (N_2057,In_1279,N_1981);
xor U2058 (N_2058,N_1848,N_907);
nand U2059 (N_2059,N_1844,N_1818);
or U2060 (N_2060,N_1902,N_1612);
nand U2061 (N_2061,N_1842,N_1942);
nand U2062 (N_2062,N_1834,N_1949);
nor U2063 (N_2063,N_1271,N_1853);
and U2064 (N_2064,N_1812,N_1867);
nand U2065 (N_2065,N_1786,N_1983);
and U2066 (N_2066,In_2476,N_1939);
or U2067 (N_2067,N_1377,In_2019);
nor U2068 (N_2068,N_1216,N_1846);
or U2069 (N_2069,N_1963,N_1752);
and U2070 (N_2070,In_920,In_634);
or U2071 (N_2071,N_1829,N_1458);
nand U2072 (N_2072,N_342,N_1965);
xor U2073 (N_2073,N_1826,N_1901);
xor U2074 (N_2074,In_1061,N_1282);
or U2075 (N_2075,N_1817,N_1657);
nand U2076 (N_2076,N_1113,N_1824);
xnor U2077 (N_2077,N_726,In_2411);
xor U2078 (N_2078,N_1671,N_1039);
or U2079 (N_2079,In_1178,N_1917);
xor U2080 (N_2080,In_1617,N_1291);
and U2081 (N_2081,N_1275,In_657);
xnor U2082 (N_2082,N_1858,N_1919);
and U2083 (N_2083,N_1825,In_1596);
or U2084 (N_2084,N_1364,N_1384);
xnor U2085 (N_2085,In_1292,N_1928);
nand U2086 (N_2086,N_674,In_1855);
or U2087 (N_2087,N_1732,N_1370);
or U2088 (N_2088,N_1661,N_1926);
nand U2089 (N_2089,N_1020,N_1813);
or U2090 (N_2090,N_1866,N_1569);
xor U2091 (N_2091,N_1937,N_1876);
nand U2092 (N_2092,In_2294,N_1870);
nand U2093 (N_2093,N_1140,N_1999);
or U2094 (N_2094,N_1811,In_1271);
nor U2095 (N_2095,N_1875,N_1720);
nor U2096 (N_2096,N_923,N_59);
or U2097 (N_2097,N_1975,N_1932);
nor U2098 (N_2098,N_1310,N_1184);
or U2099 (N_2099,N_925,N_1974);
or U2100 (N_2100,N_1643,N_1629);
and U2101 (N_2101,N_1667,In_1368);
nor U2102 (N_2102,N_500,N_1977);
xor U2103 (N_2103,N_1906,N_1346);
nor U2104 (N_2104,N_1678,N_919);
nor U2105 (N_2105,N_1815,N_1819);
or U2106 (N_2106,N_1152,N_1954);
or U2107 (N_2107,In_2280,N_1742);
and U2108 (N_2108,In_2062,N_1921);
or U2109 (N_2109,N_1198,N_1994);
xnor U2110 (N_2110,N_1908,N_1959);
and U2111 (N_2111,N_1873,In_1668);
nand U2112 (N_2112,N_1964,N_1903);
nand U2113 (N_2113,N_1395,N_1883);
nand U2114 (N_2114,N_1836,N_1957);
and U2115 (N_2115,N_643,N_456);
xnor U2116 (N_2116,In_2118,N_1288);
nor U2117 (N_2117,N_1943,N_718);
xor U2118 (N_2118,N_1985,N_1980);
xor U2119 (N_2119,N_1973,N_873);
nand U2120 (N_2120,N_984,N_1868);
and U2121 (N_2121,In_2145,N_1806);
and U2122 (N_2122,N_1010,N_260);
nor U2123 (N_2123,N_1849,N_1850);
nor U2124 (N_2124,N_1325,N_1735);
xnor U2125 (N_2125,N_1528,N_1665);
xor U2126 (N_2126,N_1864,In_501);
or U2127 (N_2127,N_1619,N_1907);
and U2128 (N_2128,N_1615,N_1889);
nand U2129 (N_2129,N_1640,N_1719);
xor U2130 (N_2130,N_1707,N_1610);
and U2131 (N_2131,N_1308,In_1261);
xor U2132 (N_2132,N_1774,N_1948);
and U2133 (N_2133,N_1878,In_826);
xnor U2134 (N_2134,N_242,N_1272);
or U2135 (N_2135,N_1967,In_777);
or U2136 (N_2136,In_2272,N_1383);
or U2137 (N_2137,N_1915,N_180);
or U2138 (N_2138,In_303,In_1194);
and U2139 (N_2139,N_1809,N_1709);
nand U2140 (N_2140,N_1186,N_1862);
or U2141 (N_2141,N_1986,N_1450);
and U2142 (N_2142,In_2248,N_1856);
nor U2143 (N_2143,N_1946,N_1276);
nor U2144 (N_2144,N_1852,N_1940);
nand U2145 (N_2145,In_629,In_4);
or U2146 (N_2146,N_1636,N_1887);
and U2147 (N_2147,N_1670,In_471);
and U2148 (N_2148,N_958,N_1366);
and U2149 (N_2149,N_1175,In_531);
nor U2150 (N_2150,N_1971,N_1881);
nand U2151 (N_2151,N_1224,N_1910);
nand U2152 (N_2152,In_1445,N_1029);
xor U2153 (N_2153,N_1904,N_1711);
and U2154 (N_2154,N_1895,In_670);
xnor U2155 (N_2155,N_647,N_1639);
or U2156 (N_2156,N_314,N_1307);
nand U2157 (N_2157,N_1518,N_1944);
or U2158 (N_2158,N_1838,N_1687);
or U2159 (N_2159,N_1871,N_1523);
or U2160 (N_2160,N_1945,In_757);
and U2161 (N_2161,N_1717,N_1326);
nor U2162 (N_2162,N_1278,N_1549);
or U2163 (N_2163,N_190,N_1913);
nor U2164 (N_2164,N_1790,N_1765);
nor U2165 (N_2165,N_1898,N_1617);
nor U2166 (N_2166,N_1777,N_1167);
nand U2167 (N_2167,N_1589,N_1918);
xor U2168 (N_2168,N_930,N_1991);
and U2169 (N_2169,N_1984,N_1800);
nand U2170 (N_2170,N_203,N_1315);
and U2171 (N_2171,In_1938,N_1642);
or U2172 (N_2172,In_535,N_1613);
and U2173 (N_2173,In_801,N_970);
or U2174 (N_2174,N_1976,N_1882);
nand U2175 (N_2175,N_132,In_945);
and U2176 (N_2176,N_1695,N_1941);
xnor U2177 (N_2177,In_1444,N_1872);
nand U2178 (N_2178,N_1662,N_1483);
and U2179 (N_2179,N_1888,N_1656);
xor U2180 (N_2180,In_2375,N_1805);
nor U2181 (N_2181,N_1936,N_1791);
xor U2182 (N_2182,N_1425,In_924);
nor U2183 (N_2183,N_1668,In_1015);
or U2184 (N_2184,N_1044,N_1501);
or U2185 (N_2185,N_1968,N_1555);
nand U2186 (N_2186,In_755,N_1896);
nand U2187 (N_2187,N_1706,N_1563);
nor U2188 (N_2188,N_1987,N_1756);
nand U2189 (N_2189,N_1934,In_1514);
and U2190 (N_2190,N_1960,N_914);
and U2191 (N_2191,N_1476,N_1830);
xor U2192 (N_2192,N_1884,N_828);
nor U2193 (N_2193,N_498,N_1874);
xor U2194 (N_2194,N_1823,N_646);
xnor U2195 (N_2195,N_1758,In_1797);
and U2196 (N_2196,In_1845,N_1674);
nand U2197 (N_2197,N_1851,N_1880);
nor U2198 (N_2198,N_1933,N_1988);
or U2199 (N_2199,N_723,N_1860);
or U2200 (N_2200,N_2160,N_2079);
nor U2201 (N_2201,N_2197,N_2154);
xor U2202 (N_2202,N_2168,N_1865);
xor U2203 (N_2203,N_1816,N_2081);
and U2204 (N_2204,N_2130,N_2111);
xnor U2205 (N_2205,N_2019,N_1150);
nor U2206 (N_2206,N_2125,N_2186);
xnor U2207 (N_2207,N_2088,N_1861);
and U2208 (N_2208,N_2006,N_2162);
and U2209 (N_2209,N_2076,N_2029);
and U2210 (N_2210,In_2430,N_1294);
nor U2211 (N_2211,N_2196,N_2185);
nand U2212 (N_2212,N_2126,In_1222);
nand U2213 (N_2213,N_1277,N_1958);
and U2214 (N_2214,N_316,N_1521);
or U2215 (N_2215,N_2108,N_2097);
and U2216 (N_2216,N_2098,N_2116);
nor U2217 (N_2217,N_2017,N_2123);
xnor U2218 (N_2218,N_2177,N_1142);
or U2219 (N_2219,N_1436,N_2000);
nand U2220 (N_2220,N_2052,N_2134);
nand U2221 (N_2221,N_1916,N_2004);
or U2222 (N_2222,N_1969,N_1301);
or U2223 (N_2223,N_1726,N_2021);
nand U2224 (N_2224,N_2109,N_1399);
and U2225 (N_2225,N_2064,N_1863);
or U2226 (N_2226,N_848,N_1743);
xnor U2227 (N_2227,N_2033,N_2054);
nand U2228 (N_2228,N_2137,N_2166);
nor U2229 (N_2229,N_1740,In_813);
or U2230 (N_2230,N_2003,N_2188);
or U2231 (N_2231,N_2025,N_989);
nor U2232 (N_2232,N_2141,N_2193);
xnor U2233 (N_2233,N_1837,N_2107);
or U2234 (N_2234,N_1909,N_1552);
nor U2235 (N_2235,N_2032,N_2057);
nand U2236 (N_2236,N_2192,N_2173);
xor U2237 (N_2237,N_1766,N_2093);
nor U2238 (N_2238,N_2143,N_2152);
nand U2239 (N_2239,N_2059,N_1899);
nor U2240 (N_2240,N_2198,N_1685);
nand U2241 (N_2241,N_2014,N_2051);
or U2242 (N_2242,N_2191,N_2018);
or U2243 (N_2243,N_1998,N_2073);
nand U2244 (N_2244,N_2066,N_2176);
nand U2245 (N_2245,N_1699,N_2078);
nand U2246 (N_2246,N_1542,N_2169);
and U2247 (N_2247,N_2011,N_2138);
nor U2248 (N_2248,N_2187,N_2090);
and U2249 (N_2249,N_2070,N_1885);
or U2250 (N_2250,N_2053,N_2135);
nor U2251 (N_2251,N_954,N_2119);
nand U2252 (N_2252,N_2139,N_2157);
or U2253 (N_2253,N_1832,N_2085);
nor U2254 (N_2254,N_1721,N_2012);
xnor U2255 (N_2255,N_1897,N_2039);
nor U2256 (N_2256,N_1633,N_2048);
nor U2257 (N_2257,N_1452,N_2023);
and U2258 (N_2258,N_1972,N_2175);
nor U2259 (N_2259,N_2043,N_1970);
and U2260 (N_2260,N_2159,N_2071);
and U2261 (N_2261,N_2007,N_2199);
or U2262 (N_2262,N_1705,N_2100);
nand U2263 (N_2263,N_1413,N_2083);
nand U2264 (N_2264,N_2028,N_2163);
xor U2265 (N_2265,N_1761,N_2102);
or U2266 (N_2266,N_2115,N_2178);
nor U2267 (N_2267,N_2036,N_2158);
nand U2268 (N_2268,N_2183,N_2072);
nand U2269 (N_2269,N_2184,N_2118);
and U2270 (N_2270,N_2084,N_1651);
nor U2271 (N_2271,N_1900,N_2190);
and U2272 (N_2272,N_1430,N_2031);
or U2273 (N_2273,N_1905,N_2156);
nand U2274 (N_2274,N_2106,N_1952);
nand U2275 (N_2275,N_2124,N_2131);
xor U2276 (N_2276,N_2174,N_2127);
or U2277 (N_2277,N_1979,N_1814);
and U2278 (N_2278,N_1923,N_179);
nor U2279 (N_2279,In_2203,N_2182);
nand U2280 (N_2280,N_1859,N_2140);
xor U2281 (N_2281,N_1398,N_1539);
and U2282 (N_2282,N_2005,N_2150);
nor U2283 (N_2283,N_1966,N_2091);
nor U2284 (N_2284,N_2050,N_2008);
nor U2285 (N_2285,N_2049,N_2001);
or U2286 (N_2286,N_2009,N_2145);
or U2287 (N_2287,N_654,N_2171);
and U2288 (N_2288,N_2080,N_2027);
and U2289 (N_2289,N_1912,N_2110);
or U2290 (N_2290,N_2002,N_596);
or U2291 (N_2291,N_2170,N_2040);
and U2292 (N_2292,N_2112,N_2015);
and U2293 (N_2293,N_2058,N_1893);
or U2294 (N_2294,N_2055,N_2086);
or U2295 (N_2295,N_1409,N_1441);
nand U2296 (N_2296,N_2077,N_883);
and U2297 (N_2297,In_2301,N_2153);
nor U2298 (N_2298,N_2069,N_1749);
and U2299 (N_2299,N_2136,N_2092);
nand U2300 (N_2300,N_2041,N_2151);
nor U2301 (N_2301,N_2120,N_2128);
nor U2302 (N_2302,N_1886,N_2105);
nand U2303 (N_2303,N_2044,N_2172);
nand U2304 (N_2304,N_2065,N_2094);
or U2305 (N_2305,N_2056,N_2089);
xor U2306 (N_2306,N_2034,N_2148);
nand U2307 (N_2307,N_2195,N_2181);
and U2308 (N_2308,N_2167,N_2010);
and U2309 (N_2309,N_2061,N_2063);
nor U2310 (N_2310,N_2149,N_2165);
nor U2311 (N_2311,N_2122,N_1808);
nand U2312 (N_2312,N_686,N_2062);
xor U2313 (N_2313,N_2035,N_1218);
nor U2314 (N_2314,N_1548,N_2045);
nand U2315 (N_2315,N_2096,N_1877);
or U2316 (N_2316,N_2060,N_2024);
nand U2317 (N_2317,N_2104,N_2030);
and U2318 (N_2318,N_2114,N_1879);
xor U2319 (N_2319,N_2082,N_2038);
or U2320 (N_2320,N_2132,N_1654);
or U2321 (N_2321,N_1455,N_2087);
nand U2322 (N_2322,N_2142,N_1763);
nand U2323 (N_2323,N_2103,N_2164);
and U2324 (N_2324,N_682,N_2022);
and U2325 (N_2325,N_1854,N_2037);
xnor U2326 (N_2326,N_2067,N_2180);
nand U2327 (N_2327,N_2042,N_2113);
xnor U2328 (N_2328,N_2179,N_969);
and U2329 (N_2329,N_1691,N_2129);
nor U2330 (N_2330,N_2161,N_2068);
xnor U2331 (N_2331,N_2189,N_381);
nor U2332 (N_2332,N_2194,N_2155);
nor U2333 (N_2333,N_2020,N_1737);
nor U2334 (N_2334,N_1890,N_2013);
or U2335 (N_2335,N_1598,N_2046);
xnor U2336 (N_2336,N_2133,N_2117);
nor U2337 (N_2337,N_1803,N_1894);
nor U2338 (N_2338,N_1840,N_2121);
nand U2339 (N_2339,N_1767,N_2075);
nand U2340 (N_2340,In_406,N_2147);
or U2341 (N_2341,N_2146,N_1171);
nand U2342 (N_2342,N_2095,N_1953);
nand U2343 (N_2343,N_2074,N_2101);
or U2344 (N_2344,N_1951,N_1993);
nand U2345 (N_2345,N_1956,N_2047);
or U2346 (N_2346,N_1962,N_2144);
and U2347 (N_2347,N_1925,In_297);
nand U2348 (N_2348,N_2099,N_2026);
nand U2349 (N_2349,N_2016,N_1857);
xnor U2350 (N_2350,N_2184,N_2172);
or U2351 (N_2351,N_2092,N_2091);
nand U2352 (N_2352,N_2022,N_2026);
nor U2353 (N_2353,N_2038,N_1766);
nand U2354 (N_2354,N_1277,N_2044);
nand U2355 (N_2355,N_2006,N_2036);
or U2356 (N_2356,N_2058,N_2168);
nand U2357 (N_2357,N_1413,N_2055);
nor U2358 (N_2358,N_989,N_1993);
nand U2359 (N_2359,N_2023,N_1894);
and U2360 (N_2360,N_2198,N_2180);
xor U2361 (N_2361,N_2009,N_2061);
and U2362 (N_2362,N_2022,N_2126);
and U2363 (N_2363,N_1969,N_2060);
nor U2364 (N_2364,N_2089,N_1890);
xnor U2365 (N_2365,N_2103,N_2197);
or U2366 (N_2366,N_1857,N_2091);
nor U2367 (N_2367,N_1455,N_654);
or U2368 (N_2368,N_2172,N_2018);
nand U2369 (N_2369,N_2134,N_2031);
xnor U2370 (N_2370,N_2003,N_2028);
and U2371 (N_2371,N_2145,N_1916);
xor U2372 (N_2372,N_2192,N_1885);
nand U2373 (N_2373,N_2130,N_2033);
and U2374 (N_2374,N_2123,N_2066);
xnor U2375 (N_2375,N_2110,N_2128);
and U2376 (N_2376,N_2096,N_954);
nor U2377 (N_2377,N_1409,N_2011);
xnor U2378 (N_2378,N_2146,N_2160);
xor U2379 (N_2379,N_1691,N_1969);
or U2380 (N_2380,N_2030,N_2152);
or U2381 (N_2381,N_2003,N_2043);
xor U2382 (N_2382,N_2177,N_2024);
nor U2383 (N_2383,N_1413,N_2046);
and U2384 (N_2384,N_2049,N_2141);
and U2385 (N_2385,N_1816,N_2064);
nor U2386 (N_2386,N_1766,N_2193);
or U2387 (N_2387,N_2180,N_1962);
nand U2388 (N_2388,N_2095,N_2192);
nor U2389 (N_2389,N_1899,N_2145);
xor U2390 (N_2390,N_1767,In_2430);
xor U2391 (N_2391,N_2032,N_2068);
and U2392 (N_2392,N_2140,N_2127);
and U2393 (N_2393,N_2199,N_1763);
and U2394 (N_2394,N_2131,N_2083);
nand U2395 (N_2395,N_2102,N_1743);
nor U2396 (N_2396,N_1972,N_2060);
and U2397 (N_2397,N_1399,N_2113);
nand U2398 (N_2398,N_2039,N_2161);
nor U2399 (N_2399,N_2179,N_1409);
xnor U2400 (N_2400,N_2202,N_2380);
nand U2401 (N_2401,N_2264,N_2326);
nor U2402 (N_2402,N_2330,N_2274);
and U2403 (N_2403,N_2339,N_2341);
and U2404 (N_2404,N_2310,N_2304);
or U2405 (N_2405,N_2324,N_2381);
xnor U2406 (N_2406,N_2217,N_2207);
xor U2407 (N_2407,N_2303,N_2225);
nor U2408 (N_2408,N_2375,N_2231);
xor U2409 (N_2409,N_2353,N_2219);
xnor U2410 (N_2410,N_2329,N_2284);
nor U2411 (N_2411,N_2328,N_2226);
or U2412 (N_2412,N_2223,N_2277);
xnor U2413 (N_2413,N_2216,N_2359);
and U2414 (N_2414,N_2252,N_2369);
and U2415 (N_2415,N_2384,N_2221);
xnor U2416 (N_2416,N_2286,N_2292);
or U2417 (N_2417,N_2336,N_2230);
xnor U2418 (N_2418,N_2287,N_2334);
nand U2419 (N_2419,N_2398,N_2364);
or U2420 (N_2420,N_2262,N_2229);
nand U2421 (N_2421,N_2257,N_2352);
and U2422 (N_2422,N_2206,N_2245);
nand U2423 (N_2423,N_2210,N_2305);
xnor U2424 (N_2424,N_2315,N_2382);
and U2425 (N_2425,N_2360,N_2344);
nor U2426 (N_2426,N_2272,N_2255);
xnor U2427 (N_2427,N_2296,N_2233);
nand U2428 (N_2428,N_2201,N_2263);
xor U2429 (N_2429,N_2214,N_2378);
and U2430 (N_2430,N_2276,N_2337);
nor U2431 (N_2431,N_2271,N_2351);
or U2432 (N_2432,N_2390,N_2213);
and U2433 (N_2433,N_2312,N_2387);
xor U2434 (N_2434,N_2393,N_2388);
nor U2435 (N_2435,N_2363,N_2383);
nor U2436 (N_2436,N_2294,N_2306);
xnor U2437 (N_2437,N_2325,N_2280);
or U2438 (N_2438,N_2224,N_2307);
and U2439 (N_2439,N_2301,N_2237);
xor U2440 (N_2440,N_2204,N_2249);
nor U2441 (N_2441,N_2370,N_2343);
nand U2442 (N_2442,N_2205,N_2374);
nor U2443 (N_2443,N_2327,N_2289);
nand U2444 (N_2444,N_2253,N_2385);
xor U2445 (N_2445,N_2338,N_2357);
and U2446 (N_2446,N_2300,N_2349);
or U2447 (N_2447,N_2258,N_2200);
xor U2448 (N_2448,N_2317,N_2358);
xor U2449 (N_2449,N_2283,N_2256);
nand U2450 (N_2450,N_2278,N_2267);
and U2451 (N_2451,N_2270,N_2345);
xnor U2452 (N_2452,N_2247,N_2285);
and U2453 (N_2453,N_2319,N_2275);
and U2454 (N_2454,N_2346,N_2293);
nand U2455 (N_2455,N_2260,N_2361);
nand U2456 (N_2456,N_2318,N_2281);
xnor U2457 (N_2457,N_2279,N_2331);
or U2458 (N_2458,N_2391,N_2355);
and U2459 (N_2459,N_2362,N_2282);
xnor U2460 (N_2460,N_2323,N_2250);
or U2461 (N_2461,N_2392,N_2313);
or U2462 (N_2462,N_2308,N_2377);
xnor U2463 (N_2463,N_2350,N_2322);
or U2464 (N_2464,N_2290,N_2373);
nor U2465 (N_2465,N_2246,N_2269);
or U2466 (N_2466,N_2342,N_2297);
and U2467 (N_2467,N_2397,N_2356);
and U2468 (N_2468,N_2395,N_2396);
nor U2469 (N_2469,N_2365,N_2220);
nand U2470 (N_2470,N_2309,N_2288);
nand U2471 (N_2471,N_2242,N_2212);
xnor U2472 (N_2472,N_2248,N_2321);
xor U2473 (N_2473,N_2209,N_2314);
nand U2474 (N_2474,N_2228,N_2218);
and U2475 (N_2475,N_2244,N_2211);
nor U2476 (N_2476,N_2251,N_2273);
nand U2477 (N_2477,N_2239,N_2232);
and U2478 (N_2478,N_2203,N_2215);
nand U2479 (N_2479,N_2299,N_2222);
xor U2480 (N_2480,N_2302,N_2295);
nor U2481 (N_2481,N_2268,N_2261);
or U2482 (N_2482,N_2236,N_2311);
or U2483 (N_2483,N_2347,N_2234);
nand U2484 (N_2484,N_2320,N_2386);
or U2485 (N_2485,N_2265,N_2389);
and U2486 (N_2486,N_2376,N_2316);
and U2487 (N_2487,N_2394,N_2266);
xnor U2488 (N_2488,N_2259,N_2333);
or U2489 (N_2489,N_2298,N_2332);
nand U2490 (N_2490,N_2399,N_2354);
and U2491 (N_2491,N_2367,N_2379);
xor U2492 (N_2492,N_2208,N_2335);
and U2493 (N_2493,N_2240,N_2366);
or U2494 (N_2494,N_2243,N_2371);
nand U2495 (N_2495,N_2368,N_2291);
nand U2496 (N_2496,N_2348,N_2227);
nand U2497 (N_2497,N_2238,N_2241);
and U2498 (N_2498,N_2254,N_2372);
nor U2499 (N_2499,N_2235,N_2340);
nor U2500 (N_2500,N_2224,N_2376);
xnor U2501 (N_2501,N_2378,N_2258);
xor U2502 (N_2502,N_2323,N_2264);
nand U2503 (N_2503,N_2352,N_2268);
and U2504 (N_2504,N_2378,N_2219);
nor U2505 (N_2505,N_2245,N_2311);
xor U2506 (N_2506,N_2368,N_2308);
nor U2507 (N_2507,N_2397,N_2286);
xor U2508 (N_2508,N_2375,N_2311);
or U2509 (N_2509,N_2382,N_2233);
or U2510 (N_2510,N_2342,N_2299);
xnor U2511 (N_2511,N_2291,N_2344);
or U2512 (N_2512,N_2269,N_2227);
and U2513 (N_2513,N_2224,N_2275);
nand U2514 (N_2514,N_2213,N_2345);
nand U2515 (N_2515,N_2322,N_2327);
nor U2516 (N_2516,N_2224,N_2255);
or U2517 (N_2517,N_2266,N_2253);
nand U2518 (N_2518,N_2315,N_2345);
nor U2519 (N_2519,N_2326,N_2274);
or U2520 (N_2520,N_2225,N_2252);
and U2521 (N_2521,N_2212,N_2368);
or U2522 (N_2522,N_2311,N_2348);
and U2523 (N_2523,N_2386,N_2200);
xor U2524 (N_2524,N_2251,N_2293);
or U2525 (N_2525,N_2398,N_2205);
nand U2526 (N_2526,N_2255,N_2308);
nor U2527 (N_2527,N_2372,N_2241);
and U2528 (N_2528,N_2299,N_2311);
or U2529 (N_2529,N_2315,N_2284);
and U2530 (N_2530,N_2338,N_2237);
or U2531 (N_2531,N_2281,N_2370);
nor U2532 (N_2532,N_2324,N_2268);
or U2533 (N_2533,N_2332,N_2227);
or U2534 (N_2534,N_2330,N_2270);
nor U2535 (N_2535,N_2326,N_2233);
nand U2536 (N_2536,N_2234,N_2292);
xor U2537 (N_2537,N_2381,N_2203);
or U2538 (N_2538,N_2374,N_2381);
and U2539 (N_2539,N_2372,N_2341);
and U2540 (N_2540,N_2279,N_2219);
nand U2541 (N_2541,N_2268,N_2344);
and U2542 (N_2542,N_2368,N_2363);
and U2543 (N_2543,N_2295,N_2318);
xnor U2544 (N_2544,N_2230,N_2253);
nand U2545 (N_2545,N_2312,N_2356);
xnor U2546 (N_2546,N_2399,N_2319);
nor U2547 (N_2547,N_2386,N_2398);
nand U2548 (N_2548,N_2287,N_2376);
or U2549 (N_2549,N_2385,N_2252);
nand U2550 (N_2550,N_2214,N_2227);
or U2551 (N_2551,N_2321,N_2358);
xnor U2552 (N_2552,N_2206,N_2335);
or U2553 (N_2553,N_2309,N_2287);
nor U2554 (N_2554,N_2230,N_2339);
nand U2555 (N_2555,N_2333,N_2203);
nor U2556 (N_2556,N_2217,N_2250);
or U2557 (N_2557,N_2240,N_2283);
xnor U2558 (N_2558,N_2267,N_2240);
xor U2559 (N_2559,N_2250,N_2366);
or U2560 (N_2560,N_2227,N_2365);
nor U2561 (N_2561,N_2210,N_2231);
xor U2562 (N_2562,N_2379,N_2227);
and U2563 (N_2563,N_2382,N_2275);
nand U2564 (N_2564,N_2287,N_2250);
and U2565 (N_2565,N_2209,N_2386);
and U2566 (N_2566,N_2370,N_2232);
nor U2567 (N_2567,N_2380,N_2266);
nand U2568 (N_2568,N_2330,N_2314);
and U2569 (N_2569,N_2336,N_2329);
nand U2570 (N_2570,N_2385,N_2257);
nor U2571 (N_2571,N_2239,N_2389);
nand U2572 (N_2572,N_2311,N_2281);
nand U2573 (N_2573,N_2399,N_2340);
nand U2574 (N_2574,N_2208,N_2386);
nand U2575 (N_2575,N_2226,N_2377);
nand U2576 (N_2576,N_2356,N_2379);
xor U2577 (N_2577,N_2351,N_2203);
xnor U2578 (N_2578,N_2345,N_2282);
xnor U2579 (N_2579,N_2326,N_2372);
or U2580 (N_2580,N_2380,N_2273);
nand U2581 (N_2581,N_2225,N_2361);
and U2582 (N_2582,N_2363,N_2394);
nor U2583 (N_2583,N_2289,N_2244);
nor U2584 (N_2584,N_2259,N_2377);
or U2585 (N_2585,N_2221,N_2367);
xnor U2586 (N_2586,N_2374,N_2208);
and U2587 (N_2587,N_2319,N_2282);
xnor U2588 (N_2588,N_2296,N_2306);
nand U2589 (N_2589,N_2334,N_2363);
xnor U2590 (N_2590,N_2306,N_2313);
nor U2591 (N_2591,N_2330,N_2399);
nor U2592 (N_2592,N_2269,N_2385);
nand U2593 (N_2593,N_2399,N_2227);
nand U2594 (N_2594,N_2276,N_2236);
and U2595 (N_2595,N_2382,N_2296);
and U2596 (N_2596,N_2396,N_2324);
xor U2597 (N_2597,N_2371,N_2233);
nor U2598 (N_2598,N_2230,N_2211);
and U2599 (N_2599,N_2282,N_2276);
xnor U2600 (N_2600,N_2480,N_2477);
xnor U2601 (N_2601,N_2431,N_2555);
nand U2602 (N_2602,N_2509,N_2452);
nor U2603 (N_2603,N_2444,N_2508);
xnor U2604 (N_2604,N_2557,N_2550);
xnor U2605 (N_2605,N_2455,N_2473);
or U2606 (N_2606,N_2464,N_2450);
or U2607 (N_2607,N_2461,N_2564);
xnor U2608 (N_2608,N_2467,N_2499);
nand U2609 (N_2609,N_2527,N_2439);
xor U2610 (N_2610,N_2515,N_2534);
nor U2611 (N_2611,N_2574,N_2541);
xor U2612 (N_2612,N_2549,N_2538);
nand U2613 (N_2613,N_2490,N_2438);
or U2614 (N_2614,N_2456,N_2587);
nor U2615 (N_2615,N_2405,N_2568);
or U2616 (N_2616,N_2585,N_2488);
xnor U2617 (N_2617,N_2521,N_2453);
nor U2618 (N_2618,N_2487,N_2579);
nand U2619 (N_2619,N_2446,N_2544);
or U2620 (N_2620,N_2553,N_2573);
and U2621 (N_2621,N_2526,N_2594);
or U2622 (N_2622,N_2443,N_2502);
and U2623 (N_2623,N_2423,N_2427);
and U2624 (N_2624,N_2517,N_2460);
nand U2625 (N_2625,N_2503,N_2409);
or U2626 (N_2626,N_2507,N_2483);
nand U2627 (N_2627,N_2432,N_2414);
nand U2628 (N_2628,N_2430,N_2468);
nor U2629 (N_2629,N_2598,N_2422);
nand U2630 (N_2630,N_2403,N_2525);
and U2631 (N_2631,N_2451,N_2583);
and U2632 (N_2632,N_2472,N_2402);
nor U2633 (N_2633,N_2532,N_2537);
nor U2634 (N_2634,N_2479,N_2514);
nand U2635 (N_2635,N_2556,N_2596);
nand U2636 (N_2636,N_2400,N_2533);
nand U2637 (N_2637,N_2447,N_2463);
xor U2638 (N_2638,N_2582,N_2481);
nand U2639 (N_2639,N_2494,N_2572);
or U2640 (N_2640,N_2559,N_2591);
and U2641 (N_2641,N_2424,N_2548);
or U2642 (N_2642,N_2566,N_2558);
and U2643 (N_2643,N_2571,N_2492);
or U2644 (N_2644,N_2415,N_2419);
nand U2645 (N_2645,N_2576,N_2457);
xnor U2646 (N_2646,N_2404,N_2454);
and U2647 (N_2647,N_2426,N_2563);
xnor U2648 (N_2648,N_2408,N_2484);
xnor U2649 (N_2649,N_2540,N_2510);
nand U2650 (N_2650,N_2554,N_2471);
xor U2651 (N_2651,N_2441,N_2567);
or U2652 (N_2652,N_2428,N_2475);
nand U2653 (N_2653,N_2493,N_2506);
xor U2654 (N_2654,N_2575,N_2401);
and U2655 (N_2655,N_2466,N_2500);
nand U2656 (N_2656,N_2412,N_2599);
or U2657 (N_2657,N_2518,N_2542);
or U2658 (N_2658,N_2470,N_2562);
or U2659 (N_2659,N_2551,N_2501);
or U2660 (N_2660,N_2592,N_2411);
nand U2661 (N_2661,N_2436,N_2417);
nand U2662 (N_2662,N_2442,N_2445);
or U2663 (N_2663,N_2569,N_2420);
nor U2664 (N_2664,N_2440,N_2528);
nand U2665 (N_2665,N_2584,N_2529);
xor U2666 (N_2666,N_2519,N_2565);
nor U2667 (N_2667,N_2505,N_2590);
xnor U2668 (N_2668,N_2546,N_2407);
and U2669 (N_2669,N_2429,N_2469);
or U2670 (N_2670,N_2421,N_2513);
or U2671 (N_2671,N_2496,N_2416);
nand U2672 (N_2672,N_2560,N_2543);
xnor U2673 (N_2673,N_2504,N_2462);
xor U2674 (N_2674,N_2561,N_2433);
and U2675 (N_2675,N_2465,N_2570);
nor U2676 (N_2676,N_2448,N_2498);
nor U2677 (N_2677,N_2516,N_2523);
nor U2678 (N_2678,N_2578,N_2520);
and U2679 (N_2679,N_2459,N_2586);
nor U2680 (N_2680,N_2418,N_2530);
nor U2681 (N_2681,N_2485,N_2476);
xnor U2682 (N_2682,N_2536,N_2588);
nor U2683 (N_2683,N_2581,N_2486);
or U2684 (N_2684,N_2437,N_2434);
nor U2685 (N_2685,N_2413,N_2474);
or U2686 (N_2686,N_2597,N_2497);
nor U2687 (N_2687,N_2593,N_2449);
and U2688 (N_2688,N_2552,N_2495);
nor U2689 (N_2689,N_2435,N_2478);
nand U2690 (N_2690,N_2589,N_2489);
or U2691 (N_2691,N_2410,N_2425);
nand U2692 (N_2692,N_2482,N_2522);
xnor U2693 (N_2693,N_2595,N_2547);
or U2694 (N_2694,N_2512,N_2458);
xor U2695 (N_2695,N_2539,N_2535);
xor U2696 (N_2696,N_2511,N_2531);
nor U2697 (N_2697,N_2524,N_2580);
or U2698 (N_2698,N_2491,N_2406);
xor U2699 (N_2699,N_2577,N_2545);
or U2700 (N_2700,N_2474,N_2467);
nor U2701 (N_2701,N_2562,N_2539);
or U2702 (N_2702,N_2540,N_2509);
nor U2703 (N_2703,N_2534,N_2492);
nor U2704 (N_2704,N_2580,N_2528);
xor U2705 (N_2705,N_2438,N_2500);
nor U2706 (N_2706,N_2438,N_2477);
nand U2707 (N_2707,N_2442,N_2514);
and U2708 (N_2708,N_2466,N_2402);
nand U2709 (N_2709,N_2569,N_2408);
nor U2710 (N_2710,N_2421,N_2599);
nand U2711 (N_2711,N_2562,N_2442);
or U2712 (N_2712,N_2466,N_2509);
nand U2713 (N_2713,N_2531,N_2419);
xor U2714 (N_2714,N_2567,N_2456);
and U2715 (N_2715,N_2496,N_2434);
nor U2716 (N_2716,N_2428,N_2571);
xnor U2717 (N_2717,N_2589,N_2415);
or U2718 (N_2718,N_2495,N_2458);
nor U2719 (N_2719,N_2431,N_2423);
nand U2720 (N_2720,N_2478,N_2576);
nand U2721 (N_2721,N_2462,N_2577);
xnor U2722 (N_2722,N_2416,N_2584);
xor U2723 (N_2723,N_2555,N_2482);
or U2724 (N_2724,N_2443,N_2511);
or U2725 (N_2725,N_2416,N_2514);
or U2726 (N_2726,N_2440,N_2457);
and U2727 (N_2727,N_2492,N_2532);
xnor U2728 (N_2728,N_2583,N_2449);
nor U2729 (N_2729,N_2512,N_2436);
and U2730 (N_2730,N_2422,N_2520);
and U2731 (N_2731,N_2539,N_2525);
and U2732 (N_2732,N_2528,N_2497);
and U2733 (N_2733,N_2535,N_2452);
nand U2734 (N_2734,N_2543,N_2506);
xor U2735 (N_2735,N_2592,N_2453);
nand U2736 (N_2736,N_2489,N_2543);
or U2737 (N_2737,N_2526,N_2452);
nor U2738 (N_2738,N_2512,N_2504);
or U2739 (N_2739,N_2498,N_2442);
and U2740 (N_2740,N_2502,N_2446);
and U2741 (N_2741,N_2474,N_2545);
nand U2742 (N_2742,N_2582,N_2560);
xnor U2743 (N_2743,N_2443,N_2499);
nand U2744 (N_2744,N_2442,N_2444);
or U2745 (N_2745,N_2502,N_2561);
or U2746 (N_2746,N_2460,N_2435);
xnor U2747 (N_2747,N_2586,N_2465);
xor U2748 (N_2748,N_2404,N_2597);
nor U2749 (N_2749,N_2584,N_2576);
and U2750 (N_2750,N_2539,N_2522);
xor U2751 (N_2751,N_2434,N_2451);
or U2752 (N_2752,N_2470,N_2477);
and U2753 (N_2753,N_2447,N_2581);
or U2754 (N_2754,N_2544,N_2455);
or U2755 (N_2755,N_2407,N_2427);
nand U2756 (N_2756,N_2555,N_2450);
nor U2757 (N_2757,N_2554,N_2580);
or U2758 (N_2758,N_2599,N_2561);
and U2759 (N_2759,N_2537,N_2560);
xnor U2760 (N_2760,N_2418,N_2536);
nor U2761 (N_2761,N_2405,N_2549);
or U2762 (N_2762,N_2573,N_2591);
xnor U2763 (N_2763,N_2499,N_2464);
or U2764 (N_2764,N_2465,N_2495);
nand U2765 (N_2765,N_2474,N_2425);
nor U2766 (N_2766,N_2544,N_2514);
nor U2767 (N_2767,N_2422,N_2414);
nor U2768 (N_2768,N_2514,N_2597);
or U2769 (N_2769,N_2512,N_2412);
nand U2770 (N_2770,N_2450,N_2519);
nand U2771 (N_2771,N_2516,N_2501);
nor U2772 (N_2772,N_2529,N_2477);
nor U2773 (N_2773,N_2489,N_2412);
and U2774 (N_2774,N_2447,N_2507);
and U2775 (N_2775,N_2483,N_2414);
or U2776 (N_2776,N_2515,N_2596);
nand U2777 (N_2777,N_2431,N_2465);
and U2778 (N_2778,N_2512,N_2511);
and U2779 (N_2779,N_2589,N_2554);
and U2780 (N_2780,N_2451,N_2597);
xnor U2781 (N_2781,N_2499,N_2404);
or U2782 (N_2782,N_2513,N_2473);
or U2783 (N_2783,N_2562,N_2479);
or U2784 (N_2784,N_2423,N_2487);
and U2785 (N_2785,N_2438,N_2483);
nor U2786 (N_2786,N_2450,N_2588);
xnor U2787 (N_2787,N_2570,N_2423);
nor U2788 (N_2788,N_2517,N_2599);
nor U2789 (N_2789,N_2560,N_2478);
nor U2790 (N_2790,N_2571,N_2558);
nor U2791 (N_2791,N_2540,N_2497);
and U2792 (N_2792,N_2558,N_2514);
nand U2793 (N_2793,N_2577,N_2472);
and U2794 (N_2794,N_2474,N_2412);
xor U2795 (N_2795,N_2573,N_2465);
nor U2796 (N_2796,N_2556,N_2564);
xor U2797 (N_2797,N_2456,N_2434);
and U2798 (N_2798,N_2520,N_2511);
and U2799 (N_2799,N_2447,N_2579);
and U2800 (N_2800,N_2765,N_2661);
nand U2801 (N_2801,N_2601,N_2774);
nor U2802 (N_2802,N_2666,N_2669);
xnor U2803 (N_2803,N_2638,N_2751);
xor U2804 (N_2804,N_2759,N_2622);
or U2805 (N_2805,N_2673,N_2725);
nand U2806 (N_2806,N_2752,N_2743);
or U2807 (N_2807,N_2635,N_2675);
nand U2808 (N_2808,N_2772,N_2619);
and U2809 (N_2809,N_2604,N_2611);
xor U2810 (N_2810,N_2794,N_2625);
or U2811 (N_2811,N_2776,N_2670);
nand U2812 (N_2812,N_2730,N_2705);
or U2813 (N_2813,N_2798,N_2680);
xnor U2814 (N_2814,N_2754,N_2607);
nand U2815 (N_2815,N_2709,N_2783);
xor U2816 (N_2816,N_2746,N_2664);
and U2817 (N_2817,N_2779,N_2636);
nor U2818 (N_2818,N_2640,N_2642);
and U2819 (N_2819,N_2782,N_2793);
nor U2820 (N_2820,N_2718,N_2722);
xor U2821 (N_2821,N_2733,N_2608);
and U2822 (N_2822,N_2708,N_2656);
or U2823 (N_2823,N_2755,N_2602);
nor U2824 (N_2824,N_2788,N_2684);
and U2825 (N_2825,N_2749,N_2614);
or U2826 (N_2826,N_2643,N_2671);
xor U2827 (N_2827,N_2653,N_2775);
xor U2828 (N_2828,N_2711,N_2726);
or U2829 (N_2829,N_2649,N_2677);
nor U2830 (N_2830,N_2645,N_2744);
nand U2831 (N_2831,N_2663,N_2689);
xnor U2832 (N_2832,N_2715,N_2764);
or U2833 (N_2833,N_2791,N_2650);
nand U2834 (N_2834,N_2735,N_2693);
nor U2835 (N_2835,N_2658,N_2695);
nor U2836 (N_2836,N_2617,N_2696);
nor U2837 (N_2837,N_2787,N_2641);
and U2838 (N_2838,N_2699,N_2603);
xnor U2839 (N_2839,N_2648,N_2609);
nand U2840 (N_2840,N_2701,N_2651);
nor U2841 (N_2841,N_2685,N_2766);
nand U2842 (N_2842,N_2734,N_2769);
or U2843 (N_2843,N_2700,N_2728);
and U2844 (N_2844,N_2691,N_2703);
or U2845 (N_2845,N_2687,N_2729);
xor U2846 (N_2846,N_2646,N_2731);
and U2847 (N_2847,N_2799,N_2613);
and U2848 (N_2848,N_2668,N_2698);
or U2849 (N_2849,N_2786,N_2750);
nand U2850 (N_2850,N_2652,N_2763);
nor U2851 (N_2851,N_2720,N_2632);
or U2852 (N_2852,N_2626,N_2678);
and U2853 (N_2853,N_2712,N_2740);
xnor U2854 (N_2854,N_2785,N_2756);
nor U2855 (N_2855,N_2736,N_2686);
nand U2856 (N_2856,N_2615,N_2630);
nand U2857 (N_2857,N_2723,N_2706);
or U2858 (N_2858,N_2761,N_2717);
or U2859 (N_2859,N_2713,N_2672);
or U2860 (N_2860,N_2721,N_2781);
and U2861 (N_2861,N_2727,N_2753);
and U2862 (N_2862,N_2644,N_2605);
or U2863 (N_2863,N_2748,N_2679);
or U2864 (N_2864,N_2758,N_2612);
and U2865 (N_2865,N_2667,N_2771);
nor U2866 (N_2866,N_2704,N_2694);
nand U2867 (N_2867,N_2628,N_2631);
or U2868 (N_2868,N_2692,N_2747);
or U2869 (N_2869,N_2738,N_2657);
nor U2870 (N_2870,N_2610,N_2681);
nand U2871 (N_2871,N_2737,N_2623);
or U2872 (N_2872,N_2716,N_2778);
nor U2873 (N_2873,N_2707,N_2757);
xnor U2874 (N_2874,N_2784,N_2789);
nor U2875 (N_2875,N_2624,N_2768);
or U2876 (N_2876,N_2647,N_2659);
and U2877 (N_2877,N_2676,N_2741);
nor U2878 (N_2878,N_2682,N_2620);
and U2879 (N_2879,N_2618,N_2792);
and U2880 (N_2880,N_2780,N_2621);
nor U2881 (N_2881,N_2683,N_2742);
and U2882 (N_2882,N_2665,N_2777);
xnor U2883 (N_2883,N_2655,N_2633);
nand U2884 (N_2884,N_2627,N_2688);
nor U2885 (N_2885,N_2762,N_2674);
nand U2886 (N_2886,N_2662,N_2660);
xor U2887 (N_2887,N_2654,N_2739);
nor U2888 (N_2888,N_2629,N_2697);
xor U2889 (N_2889,N_2790,N_2796);
and U2890 (N_2890,N_2710,N_2634);
or U2891 (N_2891,N_2795,N_2637);
nor U2892 (N_2892,N_2616,N_2745);
nand U2893 (N_2893,N_2760,N_2732);
or U2894 (N_2894,N_2714,N_2702);
nor U2895 (N_2895,N_2600,N_2797);
nand U2896 (N_2896,N_2639,N_2719);
nor U2897 (N_2897,N_2690,N_2724);
and U2898 (N_2898,N_2767,N_2770);
xor U2899 (N_2899,N_2773,N_2606);
xnor U2900 (N_2900,N_2748,N_2734);
or U2901 (N_2901,N_2741,N_2618);
xnor U2902 (N_2902,N_2664,N_2748);
nor U2903 (N_2903,N_2766,N_2650);
and U2904 (N_2904,N_2721,N_2604);
and U2905 (N_2905,N_2651,N_2720);
nor U2906 (N_2906,N_2726,N_2704);
nor U2907 (N_2907,N_2785,N_2633);
xor U2908 (N_2908,N_2620,N_2656);
and U2909 (N_2909,N_2701,N_2716);
or U2910 (N_2910,N_2798,N_2742);
nor U2911 (N_2911,N_2612,N_2630);
nand U2912 (N_2912,N_2762,N_2692);
or U2913 (N_2913,N_2664,N_2722);
nand U2914 (N_2914,N_2682,N_2699);
or U2915 (N_2915,N_2700,N_2779);
nor U2916 (N_2916,N_2738,N_2733);
nand U2917 (N_2917,N_2650,N_2726);
and U2918 (N_2918,N_2600,N_2663);
and U2919 (N_2919,N_2681,N_2763);
xnor U2920 (N_2920,N_2797,N_2675);
nand U2921 (N_2921,N_2665,N_2608);
and U2922 (N_2922,N_2687,N_2619);
nand U2923 (N_2923,N_2782,N_2704);
nor U2924 (N_2924,N_2609,N_2785);
nand U2925 (N_2925,N_2799,N_2607);
and U2926 (N_2926,N_2709,N_2753);
nor U2927 (N_2927,N_2679,N_2729);
and U2928 (N_2928,N_2686,N_2619);
and U2929 (N_2929,N_2645,N_2746);
nand U2930 (N_2930,N_2608,N_2640);
xor U2931 (N_2931,N_2752,N_2723);
nand U2932 (N_2932,N_2602,N_2699);
and U2933 (N_2933,N_2715,N_2657);
or U2934 (N_2934,N_2648,N_2753);
nor U2935 (N_2935,N_2719,N_2792);
nand U2936 (N_2936,N_2745,N_2649);
and U2937 (N_2937,N_2737,N_2747);
or U2938 (N_2938,N_2796,N_2736);
nand U2939 (N_2939,N_2618,N_2636);
and U2940 (N_2940,N_2645,N_2616);
or U2941 (N_2941,N_2723,N_2624);
and U2942 (N_2942,N_2637,N_2732);
nor U2943 (N_2943,N_2733,N_2656);
xnor U2944 (N_2944,N_2709,N_2767);
nor U2945 (N_2945,N_2742,N_2676);
xor U2946 (N_2946,N_2693,N_2780);
xnor U2947 (N_2947,N_2640,N_2668);
nor U2948 (N_2948,N_2760,N_2685);
nand U2949 (N_2949,N_2648,N_2721);
xor U2950 (N_2950,N_2618,N_2746);
xor U2951 (N_2951,N_2604,N_2798);
nand U2952 (N_2952,N_2611,N_2792);
nor U2953 (N_2953,N_2665,N_2678);
nor U2954 (N_2954,N_2770,N_2772);
and U2955 (N_2955,N_2673,N_2678);
xor U2956 (N_2956,N_2773,N_2685);
and U2957 (N_2957,N_2701,N_2791);
xnor U2958 (N_2958,N_2646,N_2791);
and U2959 (N_2959,N_2665,N_2794);
or U2960 (N_2960,N_2659,N_2605);
xnor U2961 (N_2961,N_2748,N_2789);
xnor U2962 (N_2962,N_2751,N_2677);
xor U2963 (N_2963,N_2674,N_2744);
nand U2964 (N_2964,N_2601,N_2712);
xor U2965 (N_2965,N_2721,N_2710);
nand U2966 (N_2966,N_2782,N_2623);
or U2967 (N_2967,N_2720,N_2704);
nand U2968 (N_2968,N_2745,N_2789);
xor U2969 (N_2969,N_2703,N_2716);
nor U2970 (N_2970,N_2745,N_2613);
nor U2971 (N_2971,N_2757,N_2635);
xor U2972 (N_2972,N_2621,N_2604);
or U2973 (N_2973,N_2733,N_2622);
xor U2974 (N_2974,N_2755,N_2732);
xnor U2975 (N_2975,N_2692,N_2774);
xnor U2976 (N_2976,N_2785,N_2796);
or U2977 (N_2977,N_2652,N_2625);
xnor U2978 (N_2978,N_2601,N_2698);
nor U2979 (N_2979,N_2737,N_2735);
nor U2980 (N_2980,N_2679,N_2677);
and U2981 (N_2981,N_2783,N_2796);
or U2982 (N_2982,N_2670,N_2676);
or U2983 (N_2983,N_2742,N_2668);
and U2984 (N_2984,N_2681,N_2700);
nand U2985 (N_2985,N_2635,N_2605);
and U2986 (N_2986,N_2632,N_2673);
xor U2987 (N_2987,N_2761,N_2737);
and U2988 (N_2988,N_2631,N_2652);
nand U2989 (N_2989,N_2714,N_2758);
xor U2990 (N_2990,N_2703,N_2603);
or U2991 (N_2991,N_2675,N_2776);
nor U2992 (N_2992,N_2735,N_2776);
or U2993 (N_2993,N_2606,N_2644);
nor U2994 (N_2994,N_2789,N_2733);
nand U2995 (N_2995,N_2795,N_2615);
and U2996 (N_2996,N_2629,N_2632);
or U2997 (N_2997,N_2723,N_2748);
xnor U2998 (N_2998,N_2749,N_2703);
xnor U2999 (N_2999,N_2780,N_2776);
nand U3000 (N_3000,N_2911,N_2870);
xor U3001 (N_3001,N_2878,N_2932);
and U3002 (N_3002,N_2965,N_2836);
or U3003 (N_3003,N_2921,N_2951);
nor U3004 (N_3004,N_2944,N_2988);
nor U3005 (N_3005,N_2947,N_2991);
and U3006 (N_3006,N_2957,N_2939);
nor U3007 (N_3007,N_2928,N_2848);
nor U3008 (N_3008,N_2842,N_2905);
and U3009 (N_3009,N_2845,N_2854);
nor U3010 (N_3010,N_2973,N_2974);
nand U3011 (N_3011,N_2882,N_2889);
and U3012 (N_3012,N_2999,N_2995);
nand U3013 (N_3013,N_2879,N_2948);
or U3014 (N_3014,N_2952,N_2981);
and U3015 (N_3015,N_2880,N_2916);
xor U3016 (N_3016,N_2843,N_2942);
nor U3017 (N_3017,N_2908,N_2833);
and U3018 (N_3018,N_2868,N_2931);
xor U3019 (N_3019,N_2816,N_2962);
nor U3020 (N_3020,N_2919,N_2813);
or U3021 (N_3021,N_2881,N_2820);
nand U3022 (N_3022,N_2960,N_2976);
nand U3023 (N_3023,N_2896,N_2886);
xor U3024 (N_3024,N_2834,N_2998);
or U3025 (N_3025,N_2819,N_2923);
nand U3026 (N_3026,N_2968,N_2945);
or U3027 (N_3027,N_2828,N_2824);
and U3028 (N_3028,N_2812,N_2910);
nand U3029 (N_3029,N_2810,N_2993);
nand U3030 (N_3030,N_2985,N_2907);
nand U3031 (N_3031,N_2914,N_2953);
or U3032 (N_3032,N_2927,N_2829);
nand U3033 (N_3033,N_2863,N_2804);
and U3034 (N_3034,N_2969,N_2915);
xnor U3035 (N_3035,N_2891,N_2967);
nand U3036 (N_3036,N_2901,N_2857);
or U3037 (N_3037,N_2972,N_2899);
and U3038 (N_3038,N_2975,N_2887);
nor U3039 (N_3039,N_2809,N_2937);
nand U3040 (N_3040,N_2821,N_2984);
nor U3041 (N_3041,N_2992,N_2902);
or U3042 (N_3042,N_2971,N_2946);
xor U3043 (N_3043,N_2940,N_2979);
or U3044 (N_3044,N_2936,N_2963);
xor U3045 (N_3045,N_2823,N_2888);
nand U3046 (N_3046,N_2906,N_2930);
and U3047 (N_3047,N_2933,N_2996);
xnor U3048 (N_3048,N_2801,N_2935);
or U3049 (N_3049,N_2808,N_2943);
or U3050 (N_3050,N_2852,N_2966);
nand U3051 (N_3051,N_2990,N_2876);
or U3052 (N_3052,N_2949,N_2997);
xor U3053 (N_3053,N_2830,N_2856);
nand U3054 (N_3054,N_2818,N_2892);
xnor U3055 (N_3055,N_2982,N_2897);
xnor U3056 (N_3056,N_2867,N_2866);
and U3057 (N_3057,N_2929,N_2978);
nor U3058 (N_3058,N_2822,N_2846);
xnor U3059 (N_3059,N_2850,N_2826);
nand U3060 (N_3060,N_2954,N_2893);
nor U3061 (N_3061,N_2900,N_2851);
nand U3062 (N_3062,N_2865,N_2875);
and U3063 (N_3063,N_2844,N_2924);
and U3064 (N_3064,N_2917,N_2959);
xnor U3065 (N_3065,N_2849,N_2811);
nor U3066 (N_3066,N_2994,N_2904);
nor U3067 (N_3067,N_2847,N_2890);
and U3068 (N_3068,N_2831,N_2873);
xnor U3069 (N_3069,N_2869,N_2802);
or U3070 (N_3070,N_2970,N_2920);
or U3071 (N_3071,N_2961,N_2853);
or U3072 (N_3072,N_2835,N_2898);
xnor U3073 (N_3073,N_2977,N_2922);
xor U3074 (N_3074,N_2839,N_2909);
nor U3075 (N_3075,N_2837,N_2862);
nor U3076 (N_3076,N_2926,N_2964);
xor U3077 (N_3077,N_2934,N_2913);
and U3078 (N_3078,N_2912,N_2980);
xnor U3079 (N_3079,N_2827,N_2884);
or U3080 (N_3080,N_2817,N_2885);
and U3081 (N_3081,N_2983,N_2986);
nand U3082 (N_3082,N_2858,N_2941);
xor U3083 (N_3083,N_2958,N_2956);
nor U3084 (N_3084,N_2859,N_2832);
and U3085 (N_3085,N_2806,N_2894);
nor U3086 (N_3086,N_2838,N_2841);
xnor U3087 (N_3087,N_2825,N_2872);
nor U3088 (N_3088,N_2903,N_2815);
xor U3089 (N_3089,N_2938,N_2860);
nor U3090 (N_3090,N_2805,N_2883);
or U3091 (N_3091,N_2925,N_2871);
and U3092 (N_3092,N_2874,N_2989);
and U3093 (N_3093,N_2807,N_2803);
and U3094 (N_3094,N_2877,N_2987);
or U3095 (N_3095,N_2855,N_2861);
and U3096 (N_3096,N_2918,N_2800);
nand U3097 (N_3097,N_2840,N_2955);
xnor U3098 (N_3098,N_2814,N_2864);
nand U3099 (N_3099,N_2895,N_2950);
and U3100 (N_3100,N_2881,N_2848);
nand U3101 (N_3101,N_2849,N_2960);
nand U3102 (N_3102,N_2834,N_2851);
xor U3103 (N_3103,N_2958,N_2921);
or U3104 (N_3104,N_2873,N_2878);
or U3105 (N_3105,N_2871,N_2894);
nor U3106 (N_3106,N_2879,N_2904);
nand U3107 (N_3107,N_2972,N_2997);
and U3108 (N_3108,N_2950,N_2923);
nor U3109 (N_3109,N_2815,N_2897);
or U3110 (N_3110,N_2843,N_2934);
nand U3111 (N_3111,N_2930,N_2817);
nor U3112 (N_3112,N_2821,N_2994);
and U3113 (N_3113,N_2851,N_2961);
or U3114 (N_3114,N_2923,N_2852);
nand U3115 (N_3115,N_2865,N_2810);
xor U3116 (N_3116,N_2930,N_2849);
nor U3117 (N_3117,N_2982,N_2926);
nor U3118 (N_3118,N_2969,N_2815);
and U3119 (N_3119,N_2873,N_2815);
xnor U3120 (N_3120,N_2891,N_2965);
nor U3121 (N_3121,N_2951,N_2961);
xnor U3122 (N_3122,N_2900,N_2895);
and U3123 (N_3123,N_2882,N_2858);
nor U3124 (N_3124,N_2948,N_2870);
xnor U3125 (N_3125,N_2878,N_2946);
nor U3126 (N_3126,N_2961,N_2859);
nand U3127 (N_3127,N_2889,N_2897);
nand U3128 (N_3128,N_2941,N_2817);
or U3129 (N_3129,N_2846,N_2813);
nor U3130 (N_3130,N_2981,N_2830);
xnor U3131 (N_3131,N_2898,N_2858);
and U3132 (N_3132,N_2815,N_2994);
nand U3133 (N_3133,N_2823,N_2954);
and U3134 (N_3134,N_2828,N_2915);
xnor U3135 (N_3135,N_2854,N_2800);
or U3136 (N_3136,N_2866,N_2970);
nor U3137 (N_3137,N_2880,N_2831);
xnor U3138 (N_3138,N_2919,N_2958);
nand U3139 (N_3139,N_2802,N_2888);
xor U3140 (N_3140,N_2801,N_2941);
xnor U3141 (N_3141,N_2990,N_2994);
xnor U3142 (N_3142,N_2962,N_2922);
nand U3143 (N_3143,N_2819,N_2920);
nand U3144 (N_3144,N_2861,N_2929);
nand U3145 (N_3145,N_2992,N_2858);
nand U3146 (N_3146,N_2930,N_2816);
xnor U3147 (N_3147,N_2911,N_2890);
or U3148 (N_3148,N_2812,N_2894);
or U3149 (N_3149,N_2870,N_2986);
or U3150 (N_3150,N_2953,N_2980);
xnor U3151 (N_3151,N_2809,N_2846);
nand U3152 (N_3152,N_2835,N_2843);
nor U3153 (N_3153,N_2901,N_2989);
nand U3154 (N_3154,N_2848,N_2921);
nor U3155 (N_3155,N_2912,N_2868);
nor U3156 (N_3156,N_2877,N_2840);
nand U3157 (N_3157,N_2895,N_2859);
or U3158 (N_3158,N_2965,N_2809);
xor U3159 (N_3159,N_2867,N_2811);
nand U3160 (N_3160,N_2840,N_2957);
xor U3161 (N_3161,N_2909,N_2940);
and U3162 (N_3162,N_2911,N_2897);
nand U3163 (N_3163,N_2904,N_2927);
nand U3164 (N_3164,N_2973,N_2894);
nand U3165 (N_3165,N_2862,N_2920);
xnor U3166 (N_3166,N_2926,N_2920);
and U3167 (N_3167,N_2945,N_2875);
xnor U3168 (N_3168,N_2802,N_2818);
nor U3169 (N_3169,N_2915,N_2938);
nand U3170 (N_3170,N_2815,N_2872);
and U3171 (N_3171,N_2998,N_2890);
nor U3172 (N_3172,N_2857,N_2970);
or U3173 (N_3173,N_2824,N_2946);
or U3174 (N_3174,N_2946,N_2821);
xor U3175 (N_3175,N_2917,N_2906);
xor U3176 (N_3176,N_2944,N_2870);
xnor U3177 (N_3177,N_2883,N_2907);
or U3178 (N_3178,N_2837,N_2890);
nand U3179 (N_3179,N_2971,N_2817);
xor U3180 (N_3180,N_2918,N_2877);
nor U3181 (N_3181,N_2980,N_2844);
nand U3182 (N_3182,N_2948,N_2992);
and U3183 (N_3183,N_2923,N_2874);
nand U3184 (N_3184,N_2936,N_2916);
or U3185 (N_3185,N_2941,N_2940);
nand U3186 (N_3186,N_2871,N_2943);
or U3187 (N_3187,N_2859,N_2976);
or U3188 (N_3188,N_2812,N_2834);
nor U3189 (N_3189,N_2869,N_2815);
and U3190 (N_3190,N_2869,N_2922);
nand U3191 (N_3191,N_2980,N_2816);
nand U3192 (N_3192,N_2875,N_2877);
nand U3193 (N_3193,N_2963,N_2938);
or U3194 (N_3194,N_2920,N_2932);
and U3195 (N_3195,N_2851,N_2989);
nor U3196 (N_3196,N_2800,N_2801);
nor U3197 (N_3197,N_2823,N_2880);
nor U3198 (N_3198,N_2998,N_2824);
or U3199 (N_3199,N_2807,N_2892);
and U3200 (N_3200,N_3151,N_3196);
or U3201 (N_3201,N_3084,N_3003);
nor U3202 (N_3202,N_3125,N_3090);
nor U3203 (N_3203,N_3194,N_3122);
and U3204 (N_3204,N_3012,N_3145);
and U3205 (N_3205,N_3193,N_3011);
nand U3206 (N_3206,N_3126,N_3070);
xor U3207 (N_3207,N_3015,N_3035);
xor U3208 (N_3208,N_3078,N_3014);
nand U3209 (N_3209,N_3179,N_3008);
xnor U3210 (N_3210,N_3163,N_3173);
nor U3211 (N_3211,N_3152,N_3018);
or U3212 (N_3212,N_3186,N_3185);
nand U3213 (N_3213,N_3105,N_3057);
or U3214 (N_3214,N_3104,N_3007);
nand U3215 (N_3215,N_3089,N_3146);
nand U3216 (N_3216,N_3025,N_3170);
nand U3217 (N_3217,N_3140,N_3062);
nand U3218 (N_3218,N_3021,N_3165);
nor U3219 (N_3219,N_3156,N_3024);
nor U3220 (N_3220,N_3136,N_3027);
nand U3221 (N_3221,N_3181,N_3020);
and U3222 (N_3222,N_3046,N_3036);
nor U3223 (N_3223,N_3047,N_3132);
nor U3224 (N_3224,N_3041,N_3162);
nand U3225 (N_3225,N_3175,N_3115);
or U3226 (N_3226,N_3028,N_3100);
or U3227 (N_3227,N_3017,N_3191);
xor U3228 (N_3228,N_3139,N_3172);
or U3229 (N_3229,N_3000,N_3013);
nor U3230 (N_3230,N_3153,N_3135);
nor U3231 (N_3231,N_3096,N_3009);
nand U3232 (N_3232,N_3095,N_3155);
and U3233 (N_3233,N_3030,N_3079);
and U3234 (N_3234,N_3189,N_3032);
nor U3235 (N_3235,N_3004,N_3174);
nand U3236 (N_3236,N_3187,N_3177);
and U3237 (N_3237,N_3171,N_3023);
or U3238 (N_3238,N_3103,N_3001);
nand U3239 (N_3239,N_3161,N_3199);
nand U3240 (N_3240,N_3006,N_3048);
xor U3241 (N_3241,N_3108,N_3054);
xnor U3242 (N_3242,N_3167,N_3040);
xnor U3243 (N_3243,N_3160,N_3169);
nand U3244 (N_3244,N_3124,N_3183);
nand U3245 (N_3245,N_3073,N_3102);
and U3246 (N_3246,N_3086,N_3076);
or U3247 (N_3247,N_3097,N_3166);
and U3248 (N_3248,N_3168,N_3067);
nand U3249 (N_3249,N_3064,N_3099);
nand U3250 (N_3250,N_3195,N_3154);
and U3251 (N_3251,N_3019,N_3092);
and U3252 (N_3252,N_3144,N_3128);
nor U3253 (N_3253,N_3138,N_3134);
nor U3254 (N_3254,N_3112,N_3060);
nor U3255 (N_3255,N_3055,N_3031);
nor U3256 (N_3256,N_3029,N_3198);
nand U3257 (N_3257,N_3044,N_3053);
nand U3258 (N_3258,N_3045,N_3150);
or U3259 (N_3259,N_3093,N_3052);
nor U3260 (N_3260,N_3081,N_3065);
or U3261 (N_3261,N_3056,N_3120);
xnor U3262 (N_3262,N_3111,N_3075);
xor U3263 (N_3263,N_3107,N_3026);
nand U3264 (N_3264,N_3085,N_3087);
xnor U3265 (N_3265,N_3133,N_3016);
nor U3266 (N_3266,N_3159,N_3037);
xnor U3267 (N_3267,N_3157,N_3116);
xor U3268 (N_3268,N_3130,N_3106);
or U3269 (N_3269,N_3190,N_3119);
xor U3270 (N_3270,N_3083,N_3158);
xor U3271 (N_3271,N_3137,N_3034);
xor U3272 (N_3272,N_3042,N_3077);
nand U3273 (N_3273,N_3101,N_3066);
nor U3274 (N_3274,N_3039,N_3074);
or U3275 (N_3275,N_3082,N_3184);
and U3276 (N_3276,N_3188,N_3149);
nor U3277 (N_3277,N_3131,N_3002);
and U3278 (N_3278,N_3022,N_3061);
or U3279 (N_3279,N_3010,N_3118);
nor U3280 (N_3280,N_3114,N_3094);
and U3281 (N_3281,N_3141,N_3043);
nor U3282 (N_3282,N_3080,N_3091);
nand U3283 (N_3283,N_3197,N_3110);
or U3284 (N_3284,N_3143,N_3063);
or U3285 (N_3285,N_3038,N_3098);
nor U3286 (N_3286,N_3129,N_3072);
or U3287 (N_3287,N_3049,N_3180);
nor U3288 (N_3288,N_3109,N_3058);
nor U3289 (N_3289,N_3117,N_3068);
xnor U3290 (N_3290,N_3050,N_3182);
nor U3291 (N_3291,N_3176,N_3164);
xnor U3292 (N_3292,N_3121,N_3051);
or U3293 (N_3293,N_3071,N_3005);
and U3294 (N_3294,N_3088,N_3142);
and U3295 (N_3295,N_3192,N_3069);
nand U3296 (N_3296,N_3148,N_3059);
and U3297 (N_3297,N_3178,N_3123);
nor U3298 (N_3298,N_3033,N_3127);
nand U3299 (N_3299,N_3147,N_3113);
or U3300 (N_3300,N_3058,N_3007);
nor U3301 (N_3301,N_3111,N_3078);
or U3302 (N_3302,N_3016,N_3184);
and U3303 (N_3303,N_3191,N_3106);
nor U3304 (N_3304,N_3100,N_3030);
or U3305 (N_3305,N_3004,N_3021);
and U3306 (N_3306,N_3069,N_3091);
xor U3307 (N_3307,N_3046,N_3039);
nand U3308 (N_3308,N_3126,N_3119);
xor U3309 (N_3309,N_3059,N_3041);
nand U3310 (N_3310,N_3005,N_3004);
nor U3311 (N_3311,N_3008,N_3035);
xnor U3312 (N_3312,N_3024,N_3047);
or U3313 (N_3313,N_3036,N_3150);
xor U3314 (N_3314,N_3025,N_3100);
nor U3315 (N_3315,N_3030,N_3009);
and U3316 (N_3316,N_3174,N_3014);
or U3317 (N_3317,N_3062,N_3094);
and U3318 (N_3318,N_3032,N_3187);
or U3319 (N_3319,N_3036,N_3114);
xnor U3320 (N_3320,N_3181,N_3123);
xor U3321 (N_3321,N_3196,N_3072);
or U3322 (N_3322,N_3020,N_3067);
nor U3323 (N_3323,N_3001,N_3163);
or U3324 (N_3324,N_3127,N_3119);
nand U3325 (N_3325,N_3155,N_3041);
and U3326 (N_3326,N_3197,N_3006);
or U3327 (N_3327,N_3168,N_3060);
nand U3328 (N_3328,N_3119,N_3146);
xnor U3329 (N_3329,N_3069,N_3096);
nand U3330 (N_3330,N_3003,N_3119);
nand U3331 (N_3331,N_3177,N_3070);
nor U3332 (N_3332,N_3055,N_3136);
xor U3333 (N_3333,N_3082,N_3153);
and U3334 (N_3334,N_3172,N_3111);
nand U3335 (N_3335,N_3112,N_3023);
nor U3336 (N_3336,N_3060,N_3125);
nand U3337 (N_3337,N_3004,N_3009);
or U3338 (N_3338,N_3041,N_3176);
xor U3339 (N_3339,N_3035,N_3187);
nand U3340 (N_3340,N_3055,N_3048);
nor U3341 (N_3341,N_3083,N_3032);
nand U3342 (N_3342,N_3175,N_3010);
nor U3343 (N_3343,N_3096,N_3049);
nand U3344 (N_3344,N_3071,N_3042);
or U3345 (N_3345,N_3064,N_3151);
nand U3346 (N_3346,N_3001,N_3026);
or U3347 (N_3347,N_3151,N_3121);
nor U3348 (N_3348,N_3110,N_3181);
xnor U3349 (N_3349,N_3040,N_3021);
nor U3350 (N_3350,N_3033,N_3164);
nand U3351 (N_3351,N_3110,N_3139);
nand U3352 (N_3352,N_3011,N_3099);
or U3353 (N_3353,N_3135,N_3172);
and U3354 (N_3354,N_3028,N_3025);
or U3355 (N_3355,N_3181,N_3192);
and U3356 (N_3356,N_3078,N_3019);
and U3357 (N_3357,N_3171,N_3129);
xor U3358 (N_3358,N_3124,N_3111);
and U3359 (N_3359,N_3025,N_3064);
nand U3360 (N_3360,N_3188,N_3192);
nor U3361 (N_3361,N_3121,N_3196);
nor U3362 (N_3362,N_3029,N_3156);
nand U3363 (N_3363,N_3092,N_3196);
xnor U3364 (N_3364,N_3083,N_3065);
xor U3365 (N_3365,N_3138,N_3153);
xor U3366 (N_3366,N_3022,N_3118);
nor U3367 (N_3367,N_3130,N_3190);
or U3368 (N_3368,N_3022,N_3038);
nor U3369 (N_3369,N_3021,N_3057);
and U3370 (N_3370,N_3064,N_3080);
and U3371 (N_3371,N_3068,N_3039);
xor U3372 (N_3372,N_3150,N_3048);
or U3373 (N_3373,N_3109,N_3175);
nor U3374 (N_3374,N_3093,N_3066);
xnor U3375 (N_3375,N_3091,N_3184);
nand U3376 (N_3376,N_3072,N_3043);
and U3377 (N_3377,N_3084,N_3035);
xnor U3378 (N_3378,N_3196,N_3063);
nor U3379 (N_3379,N_3040,N_3051);
nor U3380 (N_3380,N_3112,N_3032);
or U3381 (N_3381,N_3014,N_3118);
nand U3382 (N_3382,N_3030,N_3190);
nor U3383 (N_3383,N_3191,N_3004);
or U3384 (N_3384,N_3136,N_3124);
and U3385 (N_3385,N_3197,N_3020);
and U3386 (N_3386,N_3180,N_3085);
nand U3387 (N_3387,N_3034,N_3058);
xnor U3388 (N_3388,N_3076,N_3075);
or U3389 (N_3389,N_3113,N_3061);
and U3390 (N_3390,N_3110,N_3054);
nor U3391 (N_3391,N_3098,N_3198);
nand U3392 (N_3392,N_3010,N_3176);
and U3393 (N_3393,N_3037,N_3183);
xnor U3394 (N_3394,N_3196,N_3068);
nand U3395 (N_3395,N_3147,N_3001);
and U3396 (N_3396,N_3152,N_3190);
and U3397 (N_3397,N_3140,N_3065);
nand U3398 (N_3398,N_3015,N_3014);
xnor U3399 (N_3399,N_3041,N_3064);
and U3400 (N_3400,N_3359,N_3267);
and U3401 (N_3401,N_3351,N_3385);
or U3402 (N_3402,N_3274,N_3275);
nand U3403 (N_3403,N_3379,N_3352);
or U3404 (N_3404,N_3280,N_3399);
or U3405 (N_3405,N_3337,N_3384);
or U3406 (N_3406,N_3374,N_3396);
and U3407 (N_3407,N_3207,N_3202);
xor U3408 (N_3408,N_3369,N_3398);
and U3409 (N_3409,N_3229,N_3317);
nor U3410 (N_3410,N_3355,N_3278);
or U3411 (N_3411,N_3247,N_3250);
and U3412 (N_3412,N_3201,N_3332);
xor U3413 (N_3413,N_3321,N_3233);
nand U3414 (N_3414,N_3328,N_3309);
or U3415 (N_3415,N_3272,N_3345);
or U3416 (N_3416,N_3387,N_3306);
nor U3417 (N_3417,N_3238,N_3331);
or U3418 (N_3418,N_3239,N_3393);
or U3419 (N_3419,N_3262,N_3269);
nand U3420 (N_3420,N_3375,N_3290);
and U3421 (N_3421,N_3282,N_3367);
and U3422 (N_3422,N_3397,N_3324);
nand U3423 (N_3423,N_3383,N_3330);
xor U3424 (N_3424,N_3211,N_3386);
nor U3425 (N_3425,N_3333,N_3329);
or U3426 (N_3426,N_3344,N_3235);
xor U3427 (N_3427,N_3214,N_3241);
nor U3428 (N_3428,N_3311,N_3292);
and U3429 (N_3429,N_3221,N_3303);
or U3430 (N_3430,N_3289,N_3276);
nor U3431 (N_3431,N_3213,N_3318);
nor U3432 (N_3432,N_3368,N_3360);
xnor U3433 (N_3433,N_3343,N_3300);
or U3434 (N_3434,N_3243,N_3200);
nand U3435 (N_3435,N_3381,N_3362);
xnor U3436 (N_3436,N_3316,N_3258);
nor U3437 (N_3437,N_3223,N_3224);
or U3438 (N_3438,N_3227,N_3312);
nand U3439 (N_3439,N_3287,N_3323);
and U3440 (N_3440,N_3257,N_3256);
nand U3441 (N_3441,N_3335,N_3288);
or U3442 (N_3442,N_3237,N_3326);
nand U3443 (N_3443,N_3391,N_3392);
nor U3444 (N_3444,N_3314,N_3325);
xnor U3445 (N_3445,N_3307,N_3281);
nand U3446 (N_3446,N_3242,N_3286);
xor U3447 (N_3447,N_3268,N_3259);
nor U3448 (N_3448,N_3266,N_3372);
nand U3449 (N_3449,N_3255,N_3219);
or U3450 (N_3450,N_3390,N_3327);
xor U3451 (N_3451,N_3299,N_3206);
or U3452 (N_3452,N_3231,N_3340);
or U3453 (N_3453,N_3226,N_3252);
xor U3454 (N_3454,N_3365,N_3203);
or U3455 (N_3455,N_3349,N_3320);
and U3456 (N_3456,N_3222,N_3310);
xor U3457 (N_3457,N_3382,N_3217);
and U3458 (N_3458,N_3277,N_3234);
nand U3459 (N_3459,N_3338,N_3302);
xnor U3460 (N_3460,N_3270,N_3295);
and U3461 (N_3461,N_3263,N_3251);
xor U3462 (N_3462,N_3209,N_3232);
or U3463 (N_3463,N_3357,N_3388);
and U3464 (N_3464,N_3236,N_3245);
xnor U3465 (N_3465,N_3293,N_3230);
nor U3466 (N_3466,N_3339,N_3377);
and U3467 (N_3467,N_3212,N_3348);
xnor U3468 (N_3468,N_3342,N_3366);
nand U3469 (N_3469,N_3294,N_3389);
xor U3470 (N_3470,N_3297,N_3248);
nand U3471 (N_3471,N_3341,N_3216);
or U3472 (N_3472,N_3336,N_3334);
nand U3473 (N_3473,N_3370,N_3395);
nand U3474 (N_3474,N_3308,N_3347);
nor U3475 (N_3475,N_3380,N_3264);
xnor U3476 (N_3476,N_3305,N_3271);
and U3477 (N_3477,N_3253,N_3204);
nor U3478 (N_3478,N_3225,N_3261);
xor U3479 (N_3479,N_3285,N_3353);
or U3480 (N_3480,N_3208,N_3358);
or U3481 (N_3481,N_3291,N_3298);
xor U3482 (N_3482,N_3220,N_3246);
xor U3483 (N_3483,N_3371,N_3356);
nor U3484 (N_3484,N_3364,N_3354);
nor U3485 (N_3485,N_3376,N_3254);
or U3486 (N_3486,N_3228,N_3249);
xnor U3487 (N_3487,N_3322,N_3273);
or U3488 (N_3488,N_3296,N_3361);
or U3489 (N_3489,N_3284,N_3279);
and U3490 (N_3490,N_3240,N_3301);
nand U3491 (N_3491,N_3218,N_3210);
nor U3492 (N_3492,N_3215,N_3315);
and U3493 (N_3493,N_3373,N_3304);
nand U3494 (N_3494,N_3319,N_3260);
nor U3495 (N_3495,N_3350,N_3265);
or U3496 (N_3496,N_3313,N_3244);
or U3497 (N_3497,N_3363,N_3346);
xor U3498 (N_3498,N_3378,N_3394);
nor U3499 (N_3499,N_3205,N_3283);
xor U3500 (N_3500,N_3290,N_3373);
nor U3501 (N_3501,N_3272,N_3356);
xor U3502 (N_3502,N_3326,N_3273);
nor U3503 (N_3503,N_3291,N_3201);
and U3504 (N_3504,N_3212,N_3270);
nor U3505 (N_3505,N_3253,N_3250);
nor U3506 (N_3506,N_3267,N_3275);
or U3507 (N_3507,N_3358,N_3246);
nor U3508 (N_3508,N_3255,N_3319);
and U3509 (N_3509,N_3350,N_3234);
nand U3510 (N_3510,N_3218,N_3219);
or U3511 (N_3511,N_3209,N_3349);
nand U3512 (N_3512,N_3368,N_3295);
nor U3513 (N_3513,N_3269,N_3246);
nand U3514 (N_3514,N_3312,N_3361);
nand U3515 (N_3515,N_3307,N_3386);
nand U3516 (N_3516,N_3258,N_3346);
or U3517 (N_3517,N_3262,N_3361);
xnor U3518 (N_3518,N_3326,N_3385);
xor U3519 (N_3519,N_3312,N_3360);
xnor U3520 (N_3520,N_3355,N_3228);
xor U3521 (N_3521,N_3203,N_3307);
or U3522 (N_3522,N_3208,N_3357);
nor U3523 (N_3523,N_3305,N_3241);
or U3524 (N_3524,N_3370,N_3270);
nand U3525 (N_3525,N_3352,N_3351);
nor U3526 (N_3526,N_3395,N_3332);
nand U3527 (N_3527,N_3278,N_3345);
or U3528 (N_3528,N_3216,N_3259);
nor U3529 (N_3529,N_3303,N_3236);
nor U3530 (N_3530,N_3225,N_3256);
nand U3531 (N_3531,N_3359,N_3384);
and U3532 (N_3532,N_3233,N_3313);
or U3533 (N_3533,N_3308,N_3279);
nor U3534 (N_3534,N_3378,N_3396);
xor U3535 (N_3535,N_3224,N_3236);
nor U3536 (N_3536,N_3289,N_3375);
or U3537 (N_3537,N_3234,N_3209);
nand U3538 (N_3538,N_3231,N_3302);
nor U3539 (N_3539,N_3365,N_3348);
nand U3540 (N_3540,N_3314,N_3273);
xor U3541 (N_3541,N_3248,N_3200);
or U3542 (N_3542,N_3292,N_3231);
xor U3543 (N_3543,N_3243,N_3222);
nand U3544 (N_3544,N_3278,N_3391);
xnor U3545 (N_3545,N_3365,N_3210);
nor U3546 (N_3546,N_3322,N_3225);
and U3547 (N_3547,N_3294,N_3398);
or U3548 (N_3548,N_3279,N_3324);
or U3549 (N_3549,N_3269,N_3397);
xor U3550 (N_3550,N_3203,N_3284);
nor U3551 (N_3551,N_3220,N_3366);
nor U3552 (N_3552,N_3201,N_3377);
nand U3553 (N_3553,N_3317,N_3293);
xnor U3554 (N_3554,N_3357,N_3344);
or U3555 (N_3555,N_3394,N_3383);
and U3556 (N_3556,N_3301,N_3243);
and U3557 (N_3557,N_3309,N_3233);
or U3558 (N_3558,N_3389,N_3366);
nand U3559 (N_3559,N_3374,N_3359);
and U3560 (N_3560,N_3267,N_3265);
nor U3561 (N_3561,N_3207,N_3257);
nor U3562 (N_3562,N_3340,N_3209);
xnor U3563 (N_3563,N_3230,N_3321);
nand U3564 (N_3564,N_3284,N_3212);
xnor U3565 (N_3565,N_3355,N_3354);
and U3566 (N_3566,N_3373,N_3354);
nor U3567 (N_3567,N_3238,N_3224);
and U3568 (N_3568,N_3241,N_3345);
or U3569 (N_3569,N_3344,N_3200);
nor U3570 (N_3570,N_3386,N_3215);
nand U3571 (N_3571,N_3362,N_3250);
xnor U3572 (N_3572,N_3377,N_3321);
nor U3573 (N_3573,N_3222,N_3225);
xnor U3574 (N_3574,N_3215,N_3242);
nand U3575 (N_3575,N_3260,N_3386);
nor U3576 (N_3576,N_3245,N_3232);
and U3577 (N_3577,N_3327,N_3370);
xnor U3578 (N_3578,N_3293,N_3390);
or U3579 (N_3579,N_3324,N_3204);
and U3580 (N_3580,N_3216,N_3387);
nor U3581 (N_3581,N_3257,N_3375);
nor U3582 (N_3582,N_3379,N_3209);
nor U3583 (N_3583,N_3340,N_3395);
and U3584 (N_3584,N_3202,N_3339);
nor U3585 (N_3585,N_3305,N_3312);
or U3586 (N_3586,N_3348,N_3242);
nand U3587 (N_3587,N_3396,N_3296);
or U3588 (N_3588,N_3262,N_3250);
and U3589 (N_3589,N_3332,N_3251);
or U3590 (N_3590,N_3232,N_3258);
and U3591 (N_3591,N_3231,N_3290);
nor U3592 (N_3592,N_3221,N_3288);
nand U3593 (N_3593,N_3276,N_3312);
nand U3594 (N_3594,N_3399,N_3213);
xnor U3595 (N_3595,N_3285,N_3220);
nand U3596 (N_3596,N_3390,N_3224);
nor U3597 (N_3597,N_3388,N_3271);
xnor U3598 (N_3598,N_3272,N_3228);
nand U3599 (N_3599,N_3256,N_3341);
nor U3600 (N_3600,N_3594,N_3593);
and U3601 (N_3601,N_3450,N_3424);
or U3602 (N_3602,N_3412,N_3568);
and U3603 (N_3603,N_3542,N_3487);
or U3604 (N_3604,N_3585,N_3565);
and U3605 (N_3605,N_3489,N_3414);
or U3606 (N_3606,N_3590,N_3512);
and U3607 (N_3607,N_3537,N_3519);
and U3608 (N_3608,N_3571,N_3488);
nor U3609 (N_3609,N_3456,N_3469);
or U3610 (N_3610,N_3422,N_3561);
nand U3611 (N_3611,N_3458,N_3452);
or U3612 (N_3612,N_3494,N_3521);
and U3613 (N_3613,N_3545,N_3535);
or U3614 (N_3614,N_3431,N_3549);
and U3615 (N_3615,N_3502,N_3510);
nand U3616 (N_3616,N_3598,N_3455);
nand U3617 (N_3617,N_3576,N_3527);
and U3618 (N_3618,N_3581,N_3485);
or U3619 (N_3619,N_3518,N_3575);
and U3620 (N_3620,N_3573,N_3532);
nor U3621 (N_3621,N_3451,N_3477);
nor U3622 (N_3622,N_3597,N_3484);
nor U3623 (N_3623,N_3459,N_3462);
nand U3624 (N_3624,N_3437,N_3470);
or U3625 (N_3625,N_3404,N_3479);
or U3626 (N_3626,N_3547,N_3531);
xor U3627 (N_3627,N_3413,N_3574);
or U3628 (N_3628,N_3406,N_3490);
nand U3629 (N_3629,N_3592,N_3583);
nor U3630 (N_3630,N_3523,N_3405);
nand U3631 (N_3631,N_3554,N_3541);
or U3632 (N_3632,N_3587,N_3460);
and U3633 (N_3633,N_3421,N_3572);
or U3634 (N_3634,N_3411,N_3441);
and U3635 (N_3635,N_3492,N_3520);
nor U3636 (N_3636,N_3553,N_3584);
nand U3637 (N_3637,N_3439,N_3524);
or U3638 (N_3638,N_3444,N_3534);
nand U3639 (N_3639,N_3430,N_3496);
and U3640 (N_3640,N_3434,N_3570);
nor U3641 (N_3641,N_3402,N_3419);
or U3642 (N_3642,N_3569,N_3528);
nand U3643 (N_3643,N_3500,N_3515);
xor U3644 (N_3644,N_3420,N_3445);
nand U3645 (N_3645,N_3408,N_3499);
and U3646 (N_3646,N_3474,N_3464);
or U3647 (N_3647,N_3539,N_3591);
and U3648 (N_3648,N_3476,N_3415);
and U3649 (N_3649,N_3461,N_3511);
nor U3650 (N_3650,N_3482,N_3557);
or U3651 (N_3651,N_3427,N_3416);
xnor U3652 (N_3652,N_3471,N_3401);
xor U3653 (N_3653,N_3447,N_3564);
and U3654 (N_3654,N_3507,N_3425);
or U3655 (N_3655,N_3446,N_3409);
xor U3656 (N_3656,N_3467,N_3544);
nor U3657 (N_3657,N_3580,N_3483);
or U3658 (N_3658,N_3448,N_3454);
xor U3659 (N_3659,N_3486,N_3522);
or U3660 (N_3660,N_3555,N_3400);
nor U3661 (N_3661,N_3589,N_3418);
and U3662 (N_3662,N_3509,N_3508);
nor U3663 (N_3663,N_3442,N_3440);
or U3664 (N_3664,N_3438,N_3540);
xor U3665 (N_3665,N_3497,N_3559);
and U3666 (N_3666,N_3503,N_3546);
or U3667 (N_3667,N_3588,N_3526);
nor U3668 (N_3668,N_3472,N_3428);
nor U3669 (N_3669,N_3562,N_3543);
and U3670 (N_3670,N_3533,N_3426);
xor U3671 (N_3671,N_3403,N_3566);
nand U3672 (N_3672,N_3468,N_3481);
and U3673 (N_3673,N_3505,N_3501);
xnor U3674 (N_3674,N_3465,N_3407);
xnor U3675 (N_3675,N_3550,N_3548);
xnor U3676 (N_3676,N_3586,N_3453);
nand U3677 (N_3677,N_3552,N_3560);
or U3678 (N_3678,N_3530,N_3595);
and U3679 (N_3679,N_3417,N_3516);
or U3680 (N_3680,N_3498,N_3475);
nand U3681 (N_3681,N_3457,N_3567);
or U3682 (N_3682,N_3579,N_3582);
and U3683 (N_3683,N_3563,N_3473);
nor U3684 (N_3684,N_3578,N_3551);
nor U3685 (N_3685,N_3599,N_3556);
or U3686 (N_3686,N_3495,N_3429);
xor U3687 (N_3687,N_3538,N_3436);
and U3688 (N_3688,N_3491,N_3536);
and U3689 (N_3689,N_3449,N_3517);
and U3690 (N_3690,N_3433,N_3577);
nand U3691 (N_3691,N_3410,N_3435);
nand U3692 (N_3692,N_3466,N_3432);
and U3693 (N_3693,N_3514,N_3529);
and U3694 (N_3694,N_3558,N_3596);
nor U3695 (N_3695,N_3463,N_3525);
nor U3696 (N_3696,N_3480,N_3443);
or U3697 (N_3697,N_3493,N_3504);
nand U3698 (N_3698,N_3513,N_3506);
xor U3699 (N_3699,N_3423,N_3478);
nand U3700 (N_3700,N_3524,N_3523);
and U3701 (N_3701,N_3482,N_3577);
nor U3702 (N_3702,N_3412,N_3401);
or U3703 (N_3703,N_3537,N_3584);
xnor U3704 (N_3704,N_3571,N_3474);
or U3705 (N_3705,N_3403,N_3569);
nand U3706 (N_3706,N_3522,N_3573);
xor U3707 (N_3707,N_3407,N_3405);
and U3708 (N_3708,N_3475,N_3559);
or U3709 (N_3709,N_3589,N_3492);
and U3710 (N_3710,N_3531,N_3420);
or U3711 (N_3711,N_3538,N_3461);
xor U3712 (N_3712,N_3502,N_3432);
and U3713 (N_3713,N_3527,N_3520);
and U3714 (N_3714,N_3590,N_3419);
and U3715 (N_3715,N_3572,N_3579);
and U3716 (N_3716,N_3586,N_3558);
nor U3717 (N_3717,N_3489,N_3548);
or U3718 (N_3718,N_3463,N_3472);
or U3719 (N_3719,N_3543,N_3510);
and U3720 (N_3720,N_3569,N_3482);
nand U3721 (N_3721,N_3420,N_3438);
or U3722 (N_3722,N_3555,N_3464);
nor U3723 (N_3723,N_3591,N_3455);
nand U3724 (N_3724,N_3503,N_3404);
xor U3725 (N_3725,N_3446,N_3532);
and U3726 (N_3726,N_3524,N_3513);
xor U3727 (N_3727,N_3504,N_3561);
and U3728 (N_3728,N_3418,N_3401);
nor U3729 (N_3729,N_3540,N_3441);
nand U3730 (N_3730,N_3563,N_3451);
xnor U3731 (N_3731,N_3543,N_3433);
nor U3732 (N_3732,N_3562,N_3424);
xor U3733 (N_3733,N_3423,N_3565);
nor U3734 (N_3734,N_3581,N_3594);
or U3735 (N_3735,N_3502,N_3462);
xor U3736 (N_3736,N_3429,N_3422);
xnor U3737 (N_3737,N_3494,N_3463);
or U3738 (N_3738,N_3435,N_3401);
xnor U3739 (N_3739,N_3537,N_3593);
nor U3740 (N_3740,N_3482,N_3565);
and U3741 (N_3741,N_3456,N_3526);
or U3742 (N_3742,N_3544,N_3586);
nand U3743 (N_3743,N_3583,N_3549);
and U3744 (N_3744,N_3452,N_3559);
or U3745 (N_3745,N_3591,N_3541);
nor U3746 (N_3746,N_3547,N_3566);
nand U3747 (N_3747,N_3449,N_3572);
xnor U3748 (N_3748,N_3402,N_3488);
and U3749 (N_3749,N_3511,N_3446);
or U3750 (N_3750,N_3424,N_3455);
nor U3751 (N_3751,N_3458,N_3415);
nand U3752 (N_3752,N_3590,N_3591);
and U3753 (N_3753,N_3482,N_3469);
xnor U3754 (N_3754,N_3525,N_3420);
nand U3755 (N_3755,N_3431,N_3519);
xor U3756 (N_3756,N_3579,N_3490);
nand U3757 (N_3757,N_3418,N_3470);
and U3758 (N_3758,N_3499,N_3467);
nand U3759 (N_3759,N_3454,N_3428);
xnor U3760 (N_3760,N_3451,N_3499);
nand U3761 (N_3761,N_3411,N_3536);
xor U3762 (N_3762,N_3473,N_3421);
or U3763 (N_3763,N_3507,N_3584);
nand U3764 (N_3764,N_3515,N_3430);
nor U3765 (N_3765,N_3502,N_3561);
xnor U3766 (N_3766,N_3494,N_3409);
nor U3767 (N_3767,N_3558,N_3597);
xor U3768 (N_3768,N_3483,N_3515);
nand U3769 (N_3769,N_3513,N_3515);
or U3770 (N_3770,N_3532,N_3445);
nand U3771 (N_3771,N_3467,N_3410);
and U3772 (N_3772,N_3411,N_3555);
and U3773 (N_3773,N_3401,N_3474);
xnor U3774 (N_3774,N_3434,N_3523);
and U3775 (N_3775,N_3451,N_3462);
or U3776 (N_3776,N_3448,N_3437);
xor U3777 (N_3777,N_3472,N_3412);
or U3778 (N_3778,N_3494,N_3588);
nand U3779 (N_3779,N_3445,N_3524);
nor U3780 (N_3780,N_3585,N_3577);
xor U3781 (N_3781,N_3557,N_3475);
xnor U3782 (N_3782,N_3494,N_3482);
nor U3783 (N_3783,N_3502,N_3451);
nand U3784 (N_3784,N_3470,N_3494);
nand U3785 (N_3785,N_3481,N_3560);
nand U3786 (N_3786,N_3578,N_3459);
or U3787 (N_3787,N_3477,N_3553);
xnor U3788 (N_3788,N_3459,N_3499);
nand U3789 (N_3789,N_3440,N_3569);
or U3790 (N_3790,N_3562,N_3514);
nand U3791 (N_3791,N_3501,N_3568);
nand U3792 (N_3792,N_3587,N_3443);
nand U3793 (N_3793,N_3416,N_3464);
nand U3794 (N_3794,N_3533,N_3505);
xnor U3795 (N_3795,N_3411,N_3494);
and U3796 (N_3796,N_3593,N_3522);
nor U3797 (N_3797,N_3417,N_3485);
and U3798 (N_3798,N_3549,N_3416);
xor U3799 (N_3799,N_3514,N_3465);
xnor U3800 (N_3800,N_3768,N_3726);
and U3801 (N_3801,N_3646,N_3612);
and U3802 (N_3802,N_3769,N_3622);
nand U3803 (N_3803,N_3642,N_3670);
nor U3804 (N_3804,N_3641,N_3770);
xor U3805 (N_3805,N_3674,N_3725);
xnor U3806 (N_3806,N_3693,N_3650);
nor U3807 (N_3807,N_3613,N_3796);
nand U3808 (N_3808,N_3748,N_3645);
xor U3809 (N_3809,N_3694,N_3719);
and U3810 (N_3810,N_3656,N_3679);
xnor U3811 (N_3811,N_3620,N_3604);
xnor U3812 (N_3812,N_3640,N_3734);
or U3813 (N_3813,N_3720,N_3696);
nor U3814 (N_3814,N_3706,N_3601);
nor U3815 (N_3815,N_3736,N_3795);
nand U3816 (N_3816,N_3794,N_3686);
or U3817 (N_3817,N_3799,N_3715);
nor U3818 (N_3818,N_3667,N_3684);
xor U3819 (N_3819,N_3784,N_3761);
nor U3820 (N_3820,N_3669,N_3786);
or U3821 (N_3821,N_3609,N_3659);
or U3822 (N_3822,N_3774,N_3658);
or U3823 (N_3823,N_3685,N_3618);
xor U3824 (N_3824,N_3742,N_3629);
and U3825 (N_3825,N_3729,N_3633);
and U3826 (N_3826,N_3712,N_3619);
xor U3827 (N_3827,N_3749,N_3792);
and U3828 (N_3828,N_3789,N_3615);
nor U3829 (N_3829,N_3625,N_3728);
or U3830 (N_3830,N_3771,N_3760);
nand U3831 (N_3831,N_3678,N_3772);
nor U3832 (N_3832,N_3745,N_3762);
xor U3833 (N_3833,N_3709,N_3705);
xnor U3834 (N_3834,N_3649,N_3727);
or U3835 (N_3835,N_3710,N_3775);
xnor U3836 (N_3836,N_3682,N_3702);
nand U3837 (N_3837,N_3605,N_3753);
nor U3838 (N_3838,N_3689,N_3765);
nor U3839 (N_3839,N_3647,N_3756);
or U3840 (N_3840,N_3747,N_3733);
nand U3841 (N_3841,N_3634,N_3636);
nand U3842 (N_3842,N_3781,N_3721);
xor U3843 (N_3843,N_3673,N_3758);
nand U3844 (N_3844,N_3637,N_3610);
or U3845 (N_3845,N_3611,N_3699);
and U3846 (N_3846,N_3780,N_3688);
or U3847 (N_3847,N_3690,N_3773);
or U3848 (N_3848,N_3737,N_3671);
xor U3849 (N_3849,N_3757,N_3664);
nor U3850 (N_3850,N_3677,N_3676);
xnor U3851 (N_3851,N_3707,N_3687);
nand U3852 (N_3852,N_3652,N_3793);
and U3853 (N_3853,N_3714,N_3730);
xnor U3854 (N_3854,N_3644,N_3738);
and U3855 (N_3855,N_3603,N_3695);
or U3856 (N_3856,N_3648,N_3788);
and U3857 (N_3857,N_3638,N_3732);
xor U3858 (N_3858,N_3755,N_3767);
or U3859 (N_3859,N_3751,N_3666);
xnor U3860 (N_3860,N_3627,N_3791);
and U3861 (N_3861,N_3750,N_3763);
nor U3862 (N_3862,N_3662,N_3731);
xor U3863 (N_3863,N_3766,N_3681);
nand U3864 (N_3864,N_3740,N_3779);
and U3865 (N_3865,N_3777,N_3717);
and U3866 (N_3866,N_3798,N_3746);
nor U3867 (N_3867,N_3692,N_3718);
xor U3868 (N_3868,N_3764,N_3680);
nand U3869 (N_3869,N_3660,N_3600);
nand U3870 (N_3870,N_3703,N_3653);
xor U3871 (N_3871,N_3602,N_3631);
nand U3872 (N_3872,N_3630,N_3708);
xor U3873 (N_3873,N_3744,N_3661);
xor U3874 (N_3874,N_3739,N_3655);
xor U3875 (N_3875,N_3635,N_3778);
or U3876 (N_3876,N_3665,N_3668);
nand U3877 (N_3877,N_3722,N_3621);
or U3878 (N_3878,N_3754,N_3785);
nand U3879 (N_3879,N_3651,N_3614);
and U3880 (N_3880,N_3790,N_3675);
or U3881 (N_3881,N_3628,N_3663);
nor U3882 (N_3882,N_3623,N_3741);
xnor U3883 (N_3883,N_3743,N_3697);
and U3884 (N_3884,N_3711,N_3643);
nor U3885 (N_3885,N_3776,N_3701);
nand U3886 (N_3886,N_3735,N_3783);
nand U3887 (N_3887,N_3626,N_3698);
nand U3888 (N_3888,N_3632,N_3608);
nor U3889 (N_3889,N_3759,N_3713);
xor U3890 (N_3890,N_3657,N_3716);
xnor U3891 (N_3891,N_3654,N_3672);
or U3892 (N_3892,N_3724,N_3606);
nor U3893 (N_3893,N_3639,N_3797);
nand U3894 (N_3894,N_3616,N_3617);
or U3895 (N_3895,N_3752,N_3723);
or U3896 (N_3896,N_3691,N_3700);
and U3897 (N_3897,N_3624,N_3787);
or U3898 (N_3898,N_3782,N_3683);
or U3899 (N_3899,N_3607,N_3704);
xor U3900 (N_3900,N_3679,N_3603);
nand U3901 (N_3901,N_3619,N_3784);
nor U3902 (N_3902,N_3762,N_3765);
and U3903 (N_3903,N_3660,N_3776);
nor U3904 (N_3904,N_3721,N_3614);
nand U3905 (N_3905,N_3736,N_3708);
and U3906 (N_3906,N_3795,N_3600);
xor U3907 (N_3907,N_3704,N_3738);
xor U3908 (N_3908,N_3619,N_3660);
nand U3909 (N_3909,N_3663,N_3600);
xor U3910 (N_3910,N_3702,N_3755);
and U3911 (N_3911,N_3687,N_3647);
nor U3912 (N_3912,N_3707,N_3665);
xnor U3913 (N_3913,N_3673,N_3698);
nand U3914 (N_3914,N_3600,N_3746);
or U3915 (N_3915,N_3611,N_3651);
or U3916 (N_3916,N_3607,N_3725);
and U3917 (N_3917,N_3745,N_3732);
and U3918 (N_3918,N_3640,N_3786);
or U3919 (N_3919,N_3761,N_3627);
and U3920 (N_3920,N_3613,N_3749);
and U3921 (N_3921,N_3703,N_3657);
xor U3922 (N_3922,N_3653,N_3758);
or U3923 (N_3923,N_3657,N_3766);
xnor U3924 (N_3924,N_3678,N_3716);
nor U3925 (N_3925,N_3762,N_3775);
or U3926 (N_3926,N_3708,N_3744);
and U3927 (N_3927,N_3795,N_3623);
xor U3928 (N_3928,N_3696,N_3728);
or U3929 (N_3929,N_3683,N_3775);
xor U3930 (N_3930,N_3699,N_3752);
and U3931 (N_3931,N_3757,N_3654);
nor U3932 (N_3932,N_3768,N_3715);
or U3933 (N_3933,N_3603,N_3669);
nand U3934 (N_3934,N_3705,N_3648);
nand U3935 (N_3935,N_3735,N_3682);
nor U3936 (N_3936,N_3722,N_3671);
nor U3937 (N_3937,N_3681,N_3684);
nand U3938 (N_3938,N_3740,N_3605);
or U3939 (N_3939,N_3701,N_3661);
nand U3940 (N_3940,N_3660,N_3652);
nand U3941 (N_3941,N_3685,N_3668);
nand U3942 (N_3942,N_3713,N_3676);
and U3943 (N_3943,N_3661,N_3763);
nand U3944 (N_3944,N_3789,N_3645);
or U3945 (N_3945,N_3701,N_3731);
xnor U3946 (N_3946,N_3618,N_3798);
and U3947 (N_3947,N_3723,N_3706);
or U3948 (N_3948,N_3767,N_3750);
or U3949 (N_3949,N_3769,N_3654);
nor U3950 (N_3950,N_3649,N_3750);
nor U3951 (N_3951,N_3613,N_3732);
nand U3952 (N_3952,N_3689,N_3690);
xor U3953 (N_3953,N_3713,N_3666);
xnor U3954 (N_3954,N_3769,N_3689);
xor U3955 (N_3955,N_3710,N_3767);
nor U3956 (N_3956,N_3708,N_3793);
or U3957 (N_3957,N_3791,N_3605);
xor U3958 (N_3958,N_3738,N_3634);
or U3959 (N_3959,N_3799,N_3733);
nor U3960 (N_3960,N_3656,N_3722);
nand U3961 (N_3961,N_3742,N_3604);
xor U3962 (N_3962,N_3740,N_3741);
nand U3963 (N_3963,N_3687,N_3723);
or U3964 (N_3964,N_3737,N_3749);
and U3965 (N_3965,N_3644,N_3736);
and U3966 (N_3966,N_3668,N_3731);
or U3967 (N_3967,N_3778,N_3797);
nand U3968 (N_3968,N_3608,N_3797);
nand U3969 (N_3969,N_3746,N_3622);
or U3970 (N_3970,N_3608,N_3743);
nor U3971 (N_3971,N_3777,N_3657);
xor U3972 (N_3972,N_3792,N_3623);
or U3973 (N_3973,N_3662,N_3717);
and U3974 (N_3974,N_3669,N_3691);
nor U3975 (N_3975,N_3700,N_3646);
nand U3976 (N_3976,N_3664,N_3710);
and U3977 (N_3977,N_3775,N_3647);
nor U3978 (N_3978,N_3776,N_3740);
xor U3979 (N_3979,N_3725,N_3644);
nand U3980 (N_3980,N_3746,N_3720);
or U3981 (N_3981,N_3789,N_3713);
or U3982 (N_3982,N_3750,N_3694);
nand U3983 (N_3983,N_3649,N_3661);
and U3984 (N_3984,N_3602,N_3709);
and U3985 (N_3985,N_3662,N_3752);
nor U3986 (N_3986,N_3651,N_3635);
or U3987 (N_3987,N_3797,N_3640);
nor U3988 (N_3988,N_3733,N_3646);
and U3989 (N_3989,N_3767,N_3681);
or U3990 (N_3990,N_3694,N_3767);
or U3991 (N_3991,N_3616,N_3742);
or U3992 (N_3992,N_3745,N_3707);
nand U3993 (N_3993,N_3643,N_3765);
xor U3994 (N_3994,N_3603,N_3683);
nand U3995 (N_3995,N_3766,N_3747);
nor U3996 (N_3996,N_3723,N_3635);
and U3997 (N_3997,N_3606,N_3754);
nor U3998 (N_3998,N_3722,N_3793);
nor U3999 (N_3999,N_3600,N_3778);
nor U4000 (N_4000,N_3852,N_3831);
xnor U4001 (N_4001,N_3921,N_3855);
nor U4002 (N_4002,N_3899,N_3830);
nor U4003 (N_4003,N_3835,N_3932);
xor U4004 (N_4004,N_3959,N_3860);
and U4005 (N_4005,N_3821,N_3867);
or U4006 (N_4006,N_3935,N_3968);
and U4007 (N_4007,N_3942,N_3979);
nand U4008 (N_4008,N_3995,N_3965);
nand U4009 (N_4009,N_3953,N_3863);
nor U4010 (N_4010,N_3895,N_3917);
or U4011 (N_4011,N_3927,N_3873);
nor U4012 (N_4012,N_3814,N_3924);
nor U4013 (N_4013,N_3950,N_3897);
nor U4014 (N_4014,N_3914,N_3809);
and U4015 (N_4015,N_3988,N_3816);
nor U4016 (N_4016,N_3994,N_3818);
xor U4017 (N_4017,N_3902,N_3874);
nor U4018 (N_4018,N_3956,N_3944);
or U4019 (N_4019,N_3938,N_3947);
and U4020 (N_4020,N_3879,N_3972);
nand U4021 (N_4021,N_3900,N_3910);
and U4022 (N_4022,N_3827,N_3990);
nand U4023 (N_4023,N_3850,N_3892);
or U4024 (N_4024,N_3909,N_3933);
and U4025 (N_4025,N_3847,N_3941);
xor U4026 (N_4026,N_3976,N_3851);
and U4027 (N_4027,N_3811,N_3802);
nand U4028 (N_4028,N_3999,N_3951);
nand U4029 (N_4029,N_3810,N_3896);
and U4030 (N_4030,N_3870,N_3982);
nor U4031 (N_4031,N_3925,N_3853);
or U4032 (N_4032,N_3964,N_3840);
xnor U4033 (N_4033,N_3930,N_3886);
and U4034 (N_4034,N_3916,N_3807);
and U4035 (N_4035,N_3829,N_3820);
nor U4036 (N_4036,N_3985,N_3884);
nand U4037 (N_4037,N_3923,N_3974);
xor U4038 (N_4038,N_3989,N_3839);
nand U4039 (N_4039,N_3905,N_3828);
or U4040 (N_4040,N_3971,N_3966);
nor U4041 (N_4041,N_3864,N_3987);
xnor U4042 (N_4042,N_3997,N_3889);
nand U4043 (N_4043,N_3911,N_3890);
nor U4044 (N_4044,N_3806,N_3996);
or U4045 (N_4045,N_3882,N_3913);
xnor U4046 (N_4046,N_3969,N_3862);
or U4047 (N_4047,N_3844,N_3826);
nand U4048 (N_4048,N_3919,N_3977);
nor U4049 (N_4049,N_3893,N_3812);
or U4050 (N_4050,N_3878,N_3825);
and U4051 (N_4051,N_3868,N_3984);
nor U4052 (N_4052,N_3904,N_3958);
xnor U4053 (N_4053,N_3842,N_3813);
and U4054 (N_4054,N_3936,N_3940);
and U4055 (N_4055,N_3957,N_3838);
and U4056 (N_4056,N_3801,N_3954);
nand U4057 (N_4057,N_3937,N_3960);
or U4058 (N_4058,N_3943,N_3967);
nand U4059 (N_4059,N_3948,N_3912);
or U4060 (N_4060,N_3887,N_3877);
nor U4061 (N_4061,N_3993,N_3849);
xnor U4062 (N_4062,N_3983,N_3992);
and U4063 (N_4063,N_3980,N_3856);
nor U4064 (N_4064,N_3804,N_3875);
nor U4065 (N_4065,N_3832,N_3836);
nor U4066 (N_4066,N_3837,N_3815);
xnor U4067 (N_4067,N_3834,N_3833);
and U4068 (N_4068,N_3822,N_3888);
nor U4069 (N_4069,N_3908,N_3929);
nand U4070 (N_4070,N_3991,N_3843);
xor U4071 (N_4071,N_3846,N_3934);
xor U4072 (N_4072,N_3926,N_3885);
or U4073 (N_4073,N_3891,N_3803);
xor U4074 (N_4074,N_3883,N_3961);
xor U4075 (N_4075,N_3939,N_3848);
nand U4076 (N_4076,N_3872,N_3808);
nand U4077 (N_4077,N_3978,N_3903);
or U4078 (N_4078,N_3922,N_3817);
and U4079 (N_4079,N_3845,N_3894);
and U4080 (N_4080,N_3920,N_3963);
xor U4081 (N_4081,N_3861,N_3970);
or U4082 (N_4082,N_3823,N_3949);
nor U4083 (N_4083,N_3975,N_3865);
and U4084 (N_4084,N_3881,N_3854);
or U4085 (N_4085,N_3876,N_3841);
or U4086 (N_4086,N_3928,N_3986);
nor U4087 (N_4087,N_3955,N_3857);
or U4088 (N_4088,N_3859,N_3907);
xor U4089 (N_4089,N_3981,N_3880);
and U4090 (N_4090,N_3866,N_3819);
or U4091 (N_4091,N_3898,N_3952);
nand U4092 (N_4092,N_3962,N_3858);
nor U4093 (N_4093,N_3946,N_3800);
nor U4094 (N_4094,N_3901,N_3869);
and U4095 (N_4095,N_3998,N_3973);
nand U4096 (N_4096,N_3945,N_3906);
nor U4097 (N_4097,N_3824,N_3918);
xor U4098 (N_4098,N_3871,N_3931);
xor U4099 (N_4099,N_3805,N_3915);
nand U4100 (N_4100,N_3969,N_3856);
xor U4101 (N_4101,N_3983,N_3938);
xor U4102 (N_4102,N_3835,N_3974);
xor U4103 (N_4103,N_3926,N_3863);
or U4104 (N_4104,N_3968,N_3815);
nand U4105 (N_4105,N_3829,N_3994);
nand U4106 (N_4106,N_3868,N_3966);
and U4107 (N_4107,N_3911,N_3878);
xnor U4108 (N_4108,N_3841,N_3941);
nor U4109 (N_4109,N_3834,N_3861);
or U4110 (N_4110,N_3822,N_3840);
nor U4111 (N_4111,N_3850,N_3825);
xor U4112 (N_4112,N_3944,N_3804);
nor U4113 (N_4113,N_3917,N_3910);
and U4114 (N_4114,N_3909,N_3977);
xor U4115 (N_4115,N_3977,N_3964);
and U4116 (N_4116,N_3992,N_3883);
nor U4117 (N_4117,N_3800,N_3844);
nor U4118 (N_4118,N_3998,N_3932);
nor U4119 (N_4119,N_3963,N_3859);
nor U4120 (N_4120,N_3939,N_3941);
nand U4121 (N_4121,N_3937,N_3884);
nand U4122 (N_4122,N_3960,N_3806);
or U4123 (N_4123,N_3895,N_3957);
nand U4124 (N_4124,N_3962,N_3882);
or U4125 (N_4125,N_3952,N_3843);
or U4126 (N_4126,N_3977,N_3988);
or U4127 (N_4127,N_3822,N_3904);
nand U4128 (N_4128,N_3830,N_3874);
nor U4129 (N_4129,N_3926,N_3803);
nand U4130 (N_4130,N_3848,N_3871);
xnor U4131 (N_4131,N_3934,N_3893);
or U4132 (N_4132,N_3910,N_3981);
or U4133 (N_4133,N_3941,N_3950);
nor U4134 (N_4134,N_3869,N_3848);
nand U4135 (N_4135,N_3974,N_3884);
xnor U4136 (N_4136,N_3803,N_3968);
nand U4137 (N_4137,N_3923,N_3882);
nor U4138 (N_4138,N_3908,N_3914);
xnor U4139 (N_4139,N_3998,N_3963);
nand U4140 (N_4140,N_3910,N_3993);
and U4141 (N_4141,N_3809,N_3858);
nand U4142 (N_4142,N_3985,N_3860);
xor U4143 (N_4143,N_3818,N_3981);
and U4144 (N_4144,N_3982,N_3887);
xor U4145 (N_4145,N_3970,N_3941);
or U4146 (N_4146,N_3948,N_3884);
nor U4147 (N_4147,N_3827,N_3885);
and U4148 (N_4148,N_3802,N_3880);
xnor U4149 (N_4149,N_3974,N_3801);
or U4150 (N_4150,N_3841,N_3972);
nor U4151 (N_4151,N_3848,N_3842);
nand U4152 (N_4152,N_3803,N_3979);
or U4153 (N_4153,N_3956,N_3971);
nor U4154 (N_4154,N_3855,N_3876);
and U4155 (N_4155,N_3813,N_3877);
or U4156 (N_4156,N_3916,N_3931);
or U4157 (N_4157,N_3990,N_3861);
and U4158 (N_4158,N_3882,N_3918);
nand U4159 (N_4159,N_3982,N_3873);
and U4160 (N_4160,N_3880,N_3873);
and U4161 (N_4161,N_3862,N_3815);
xor U4162 (N_4162,N_3906,N_3884);
or U4163 (N_4163,N_3963,N_3994);
xor U4164 (N_4164,N_3940,N_3951);
nand U4165 (N_4165,N_3960,N_3938);
nor U4166 (N_4166,N_3885,N_3841);
and U4167 (N_4167,N_3863,N_3908);
nand U4168 (N_4168,N_3895,N_3900);
nand U4169 (N_4169,N_3914,N_3916);
or U4170 (N_4170,N_3871,N_3830);
or U4171 (N_4171,N_3930,N_3895);
or U4172 (N_4172,N_3956,N_3947);
or U4173 (N_4173,N_3970,N_3995);
xor U4174 (N_4174,N_3813,N_3892);
xnor U4175 (N_4175,N_3925,N_3856);
and U4176 (N_4176,N_3944,N_3803);
nor U4177 (N_4177,N_3877,N_3853);
nand U4178 (N_4178,N_3898,N_3986);
nand U4179 (N_4179,N_3880,N_3899);
nor U4180 (N_4180,N_3947,N_3802);
or U4181 (N_4181,N_3999,N_3970);
or U4182 (N_4182,N_3992,N_3808);
or U4183 (N_4183,N_3856,N_3916);
and U4184 (N_4184,N_3867,N_3981);
nor U4185 (N_4185,N_3956,N_3916);
and U4186 (N_4186,N_3903,N_3865);
nand U4187 (N_4187,N_3869,N_3879);
xnor U4188 (N_4188,N_3802,N_3978);
or U4189 (N_4189,N_3934,N_3914);
or U4190 (N_4190,N_3916,N_3949);
nor U4191 (N_4191,N_3818,N_3843);
xor U4192 (N_4192,N_3974,N_3894);
xnor U4193 (N_4193,N_3889,N_3860);
nand U4194 (N_4194,N_3804,N_3918);
nor U4195 (N_4195,N_3972,N_3865);
nor U4196 (N_4196,N_3964,N_3914);
or U4197 (N_4197,N_3942,N_3883);
or U4198 (N_4198,N_3985,N_3853);
and U4199 (N_4199,N_3827,N_3936);
nand U4200 (N_4200,N_4157,N_4104);
nor U4201 (N_4201,N_4042,N_4162);
xnor U4202 (N_4202,N_4122,N_4166);
nand U4203 (N_4203,N_4126,N_4101);
xnor U4204 (N_4204,N_4083,N_4021);
or U4205 (N_4205,N_4170,N_4185);
xnor U4206 (N_4206,N_4048,N_4159);
and U4207 (N_4207,N_4179,N_4191);
xor U4208 (N_4208,N_4198,N_4006);
and U4209 (N_4209,N_4168,N_4046);
xor U4210 (N_4210,N_4149,N_4105);
and U4211 (N_4211,N_4011,N_4091);
or U4212 (N_4212,N_4161,N_4040);
nor U4213 (N_4213,N_4100,N_4088);
and U4214 (N_4214,N_4036,N_4098);
nand U4215 (N_4215,N_4132,N_4069);
nand U4216 (N_4216,N_4033,N_4073);
nand U4217 (N_4217,N_4052,N_4173);
nor U4218 (N_4218,N_4188,N_4026);
or U4219 (N_4219,N_4136,N_4193);
nor U4220 (N_4220,N_4063,N_4038);
xnor U4221 (N_4221,N_4109,N_4153);
nand U4222 (N_4222,N_4181,N_4107);
nand U4223 (N_4223,N_4061,N_4123);
or U4224 (N_4224,N_4054,N_4145);
nand U4225 (N_4225,N_4001,N_4096);
or U4226 (N_4226,N_4084,N_4090);
xor U4227 (N_4227,N_4092,N_4043);
nor U4228 (N_4228,N_4014,N_4031);
nor U4229 (N_4229,N_4089,N_4189);
or U4230 (N_4230,N_4039,N_4174);
or U4231 (N_4231,N_4087,N_4066);
nor U4232 (N_4232,N_4195,N_4130);
or U4233 (N_4233,N_4121,N_4051);
and U4234 (N_4234,N_4057,N_4065);
xor U4235 (N_4235,N_4028,N_4172);
nor U4236 (N_4236,N_4080,N_4111);
or U4237 (N_4237,N_4183,N_4150);
nand U4238 (N_4238,N_4176,N_4147);
nand U4239 (N_4239,N_4072,N_4005);
or U4240 (N_4240,N_4064,N_4029);
nor U4241 (N_4241,N_4143,N_4023);
or U4242 (N_4242,N_4171,N_4099);
nor U4243 (N_4243,N_4124,N_4160);
xnor U4244 (N_4244,N_4140,N_4118);
nor U4245 (N_4245,N_4192,N_4058);
or U4246 (N_4246,N_4075,N_4167);
or U4247 (N_4247,N_4041,N_4044);
xnor U4248 (N_4248,N_4017,N_4196);
nand U4249 (N_4249,N_4102,N_4094);
nand U4250 (N_4250,N_4128,N_4116);
nand U4251 (N_4251,N_4151,N_4027);
nand U4252 (N_4252,N_4154,N_4049);
xnor U4253 (N_4253,N_4097,N_4178);
or U4254 (N_4254,N_4060,N_4067);
or U4255 (N_4255,N_4062,N_4025);
nand U4256 (N_4256,N_4139,N_4035);
or U4257 (N_4257,N_4169,N_4165);
and U4258 (N_4258,N_4115,N_4022);
xor U4259 (N_4259,N_4095,N_4037);
or U4260 (N_4260,N_4148,N_4138);
xor U4261 (N_4261,N_4079,N_4155);
xor U4262 (N_4262,N_4158,N_4110);
and U4263 (N_4263,N_4137,N_4142);
xnor U4264 (N_4264,N_4125,N_4177);
nand U4265 (N_4265,N_4004,N_4070);
xnor U4266 (N_4266,N_4010,N_4112);
or U4267 (N_4267,N_4059,N_4019);
nand U4268 (N_4268,N_4009,N_4103);
nand U4269 (N_4269,N_4032,N_4146);
or U4270 (N_4270,N_4013,N_4068);
nor U4271 (N_4271,N_4002,N_4175);
nand U4272 (N_4272,N_4093,N_4141);
nor U4273 (N_4273,N_4082,N_4199);
nor U4274 (N_4274,N_4020,N_4197);
xnor U4275 (N_4275,N_4108,N_4056);
nand U4276 (N_4276,N_4007,N_4074);
or U4277 (N_4277,N_4053,N_4047);
or U4278 (N_4278,N_4078,N_4045);
nor U4279 (N_4279,N_4106,N_4120);
or U4280 (N_4280,N_4113,N_4024);
nor U4281 (N_4281,N_4144,N_4184);
and U4282 (N_4282,N_4050,N_4071);
or U4283 (N_4283,N_4076,N_4163);
or U4284 (N_4284,N_4012,N_4086);
and U4285 (N_4285,N_4187,N_4134);
xnor U4286 (N_4286,N_4085,N_4030);
and U4287 (N_4287,N_4129,N_4034);
nand U4288 (N_4288,N_4081,N_4117);
nor U4289 (N_4289,N_4164,N_4055);
or U4290 (N_4290,N_4152,N_4018);
and U4291 (N_4291,N_4190,N_4194);
nor U4292 (N_4292,N_4077,N_4135);
xnor U4293 (N_4293,N_4015,N_4156);
xnor U4294 (N_4294,N_4008,N_4182);
xnor U4295 (N_4295,N_4003,N_4133);
nand U4296 (N_4296,N_4114,N_4186);
nand U4297 (N_4297,N_4127,N_4180);
or U4298 (N_4298,N_4131,N_4016);
and U4299 (N_4299,N_4119,N_4000);
nand U4300 (N_4300,N_4181,N_4160);
or U4301 (N_4301,N_4099,N_4165);
nand U4302 (N_4302,N_4166,N_4180);
xnor U4303 (N_4303,N_4045,N_4185);
or U4304 (N_4304,N_4176,N_4180);
and U4305 (N_4305,N_4148,N_4018);
and U4306 (N_4306,N_4192,N_4129);
xor U4307 (N_4307,N_4116,N_4042);
or U4308 (N_4308,N_4153,N_4017);
and U4309 (N_4309,N_4117,N_4089);
and U4310 (N_4310,N_4082,N_4012);
nor U4311 (N_4311,N_4149,N_4136);
and U4312 (N_4312,N_4038,N_4183);
and U4313 (N_4313,N_4186,N_4086);
and U4314 (N_4314,N_4055,N_4096);
nand U4315 (N_4315,N_4006,N_4079);
nand U4316 (N_4316,N_4016,N_4113);
and U4317 (N_4317,N_4038,N_4022);
nor U4318 (N_4318,N_4137,N_4116);
or U4319 (N_4319,N_4128,N_4143);
nand U4320 (N_4320,N_4052,N_4191);
or U4321 (N_4321,N_4065,N_4177);
nand U4322 (N_4322,N_4003,N_4022);
xnor U4323 (N_4323,N_4036,N_4190);
nor U4324 (N_4324,N_4076,N_4142);
nor U4325 (N_4325,N_4057,N_4177);
and U4326 (N_4326,N_4053,N_4168);
xor U4327 (N_4327,N_4127,N_4116);
nand U4328 (N_4328,N_4009,N_4020);
nand U4329 (N_4329,N_4100,N_4058);
nand U4330 (N_4330,N_4064,N_4036);
or U4331 (N_4331,N_4119,N_4026);
or U4332 (N_4332,N_4007,N_4066);
nand U4333 (N_4333,N_4091,N_4128);
nor U4334 (N_4334,N_4083,N_4126);
xor U4335 (N_4335,N_4162,N_4002);
and U4336 (N_4336,N_4124,N_4189);
nor U4337 (N_4337,N_4103,N_4045);
xor U4338 (N_4338,N_4047,N_4151);
or U4339 (N_4339,N_4093,N_4138);
or U4340 (N_4340,N_4154,N_4176);
nor U4341 (N_4341,N_4080,N_4130);
and U4342 (N_4342,N_4125,N_4192);
nor U4343 (N_4343,N_4078,N_4122);
nand U4344 (N_4344,N_4028,N_4072);
and U4345 (N_4345,N_4125,N_4158);
nor U4346 (N_4346,N_4162,N_4096);
nand U4347 (N_4347,N_4123,N_4039);
nor U4348 (N_4348,N_4007,N_4055);
or U4349 (N_4349,N_4197,N_4090);
or U4350 (N_4350,N_4030,N_4116);
nor U4351 (N_4351,N_4118,N_4008);
nand U4352 (N_4352,N_4078,N_4161);
and U4353 (N_4353,N_4087,N_4038);
xnor U4354 (N_4354,N_4184,N_4084);
nor U4355 (N_4355,N_4012,N_4087);
nand U4356 (N_4356,N_4131,N_4155);
or U4357 (N_4357,N_4000,N_4187);
and U4358 (N_4358,N_4034,N_4080);
nand U4359 (N_4359,N_4109,N_4106);
nor U4360 (N_4360,N_4160,N_4025);
or U4361 (N_4361,N_4113,N_4151);
xnor U4362 (N_4362,N_4165,N_4189);
nor U4363 (N_4363,N_4042,N_4092);
nor U4364 (N_4364,N_4133,N_4005);
nand U4365 (N_4365,N_4051,N_4027);
nand U4366 (N_4366,N_4081,N_4138);
nand U4367 (N_4367,N_4179,N_4145);
nor U4368 (N_4368,N_4178,N_4080);
nand U4369 (N_4369,N_4091,N_4025);
nor U4370 (N_4370,N_4067,N_4098);
and U4371 (N_4371,N_4081,N_4055);
nand U4372 (N_4372,N_4121,N_4029);
nand U4373 (N_4373,N_4027,N_4168);
xor U4374 (N_4374,N_4069,N_4160);
and U4375 (N_4375,N_4110,N_4186);
nand U4376 (N_4376,N_4084,N_4083);
and U4377 (N_4377,N_4187,N_4072);
and U4378 (N_4378,N_4020,N_4110);
xnor U4379 (N_4379,N_4021,N_4192);
or U4380 (N_4380,N_4014,N_4102);
or U4381 (N_4381,N_4050,N_4034);
and U4382 (N_4382,N_4016,N_4023);
or U4383 (N_4383,N_4142,N_4010);
and U4384 (N_4384,N_4122,N_4127);
nand U4385 (N_4385,N_4099,N_4121);
nand U4386 (N_4386,N_4186,N_4004);
and U4387 (N_4387,N_4032,N_4137);
or U4388 (N_4388,N_4098,N_4081);
nand U4389 (N_4389,N_4028,N_4070);
nand U4390 (N_4390,N_4006,N_4152);
or U4391 (N_4391,N_4044,N_4084);
xnor U4392 (N_4392,N_4030,N_4026);
nor U4393 (N_4393,N_4127,N_4111);
nand U4394 (N_4394,N_4138,N_4120);
xnor U4395 (N_4395,N_4074,N_4081);
xnor U4396 (N_4396,N_4198,N_4017);
nand U4397 (N_4397,N_4006,N_4054);
and U4398 (N_4398,N_4076,N_4049);
and U4399 (N_4399,N_4024,N_4192);
nand U4400 (N_4400,N_4204,N_4374);
or U4401 (N_4401,N_4371,N_4269);
nand U4402 (N_4402,N_4211,N_4238);
or U4403 (N_4403,N_4214,N_4376);
xor U4404 (N_4404,N_4347,N_4283);
or U4405 (N_4405,N_4206,N_4277);
and U4406 (N_4406,N_4393,N_4242);
xnor U4407 (N_4407,N_4378,N_4304);
xor U4408 (N_4408,N_4240,N_4261);
nand U4409 (N_4409,N_4249,N_4330);
or U4410 (N_4410,N_4389,N_4341);
xnor U4411 (N_4411,N_4383,N_4245);
or U4412 (N_4412,N_4287,N_4220);
xor U4413 (N_4413,N_4346,N_4243);
xnor U4414 (N_4414,N_4273,N_4201);
nor U4415 (N_4415,N_4328,N_4307);
and U4416 (N_4416,N_4316,N_4230);
nor U4417 (N_4417,N_4372,N_4293);
and U4418 (N_4418,N_4280,N_4298);
and U4419 (N_4419,N_4381,N_4260);
nor U4420 (N_4420,N_4311,N_4396);
and U4421 (N_4421,N_4315,N_4336);
xor U4422 (N_4422,N_4392,N_4387);
nand U4423 (N_4423,N_4366,N_4213);
and U4424 (N_4424,N_4369,N_4275);
and U4425 (N_4425,N_4340,N_4297);
xor U4426 (N_4426,N_4253,N_4377);
xnor U4427 (N_4427,N_4251,N_4332);
and U4428 (N_4428,N_4241,N_4278);
nand U4429 (N_4429,N_4239,N_4248);
xnor U4430 (N_4430,N_4270,N_4344);
or U4431 (N_4431,N_4385,N_4256);
nor U4432 (N_4432,N_4319,N_4320);
and U4433 (N_4433,N_4360,N_4382);
nand U4434 (N_4434,N_4244,N_4294);
nor U4435 (N_4435,N_4342,N_4227);
xnor U4436 (N_4436,N_4345,N_4365);
or U4437 (N_4437,N_4289,N_4303);
or U4438 (N_4438,N_4209,N_4208);
nor U4439 (N_4439,N_4339,N_4224);
nand U4440 (N_4440,N_4218,N_4234);
and U4441 (N_4441,N_4397,N_4312);
and U4442 (N_4442,N_4321,N_4355);
xor U4443 (N_4443,N_4246,N_4284);
xor U4444 (N_4444,N_4394,N_4237);
nand U4445 (N_4445,N_4325,N_4235);
xor U4446 (N_4446,N_4354,N_4301);
or U4447 (N_4447,N_4221,N_4254);
nor U4448 (N_4448,N_4228,N_4250);
and U4449 (N_4449,N_4216,N_4231);
xnor U4450 (N_4450,N_4290,N_4252);
or U4451 (N_4451,N_4317,N_4322);
nor U4452 (N_4452,N_4257,N_4205);
and U4453 (N_4453,N_4375,N_4306);
or U4454 (N_4454,N_4364,N_4262);
nand U4455 (N_4455,N_4236,N_4274);
xor U4456 (N_4456,N_4357,N_4348);
nor U4457 (N_4457,N_4281,N_4395);
nand U4458 (N_4458,N_4329,N_4265);
or U4459 (N_4459,N_4258,N_4313);
nand U4460 (N_4460,N_4279,N_4217);
or U4461 (N_4461,N_4398,N_4334);
nand U4462 (N_4462,N_4222,N_4386);
nor U4463 (N_4463,N_4215,N_4314);
or U4464 (N_4464,N_4363,N_4350);
and U4465 (N_4465,N_4362,N_4223);
nand U4466 (N_4466,N_4384,N_4391);
nand U4467 (N_4467,N_4296,N_4352);
nor U4468 (N_4468,N_4361,N_4351);
nand U4469 (N_4469,N_4202,N_4327);
or U4470 (N_4470,N_4318,N_4232);
or U4471 (N_4471,N_4309,N_4367);
and U4472 (N_4472,N_4305,N_4247);
and U4473 (N_4473,N_4299,N_4388);
nor U4474 (N_4474,N_4380,N_4292);
and U4475 (N_4475,N_4356,N_4308);
nor U4476 (N_4476,N_4337,N_4358);
and U4477 (N_4477,N_4291,N_4268);
nand U4478 (N_4478,N_4379,N_4255);
or U4479 (N_4479,N_4333,N_4370);
and U4480 (N_4480,N_4288,N_4263);
nand U4481 (N_4481,N_4302,N_4267);
nor U4482 (N_4482,N_4353,N_4200);
nand U4483 (N_4483,N_4259,N_4207);
xnor U4484 (N_4484,N_4285,N_4368);
xnor U4485 (N_4485,N_4272,N_4295);
nand U4486 (N_4486,N_4399,N_4226);
nor U4487 (N_4487,N_4359,N_4324);
xnor U4488 (N_4488,N_4271,N_4210);
xor U4489 (N_4489,N_4323,N_4310);
and U4490 (N_4490,N_4373,N_4331);
and U4491 (N_4491,N_4343,N_4349);
nand U4492 (N_4492,N_4282,N_4286);
nor U4493 (N_4493,N_4203,N_4264);
nand U4494 (N_4494,N_4233,N_4338);
or U4495 (N_4495,N_4335,N_4219);
nand U4496 (N_4496,N_4326,N_4390);
xor U4497 (N_4497,N_4229,N_4276);
nor U4498 (N_4498,N_4212,N_4266);
nand U4499 (N_4499,N_4300,N_4225);
nor U4500 (N_4500,N_4282,N_4212);
nand U4501 (N_4501,N_4329,N_4268);
or U4502 (N_4502,N_4380,N_4253);
nand U4503 (N_4503,N_4298,N_4371);
nor U4504 (N_4504,N_4384,N_4286);
xor U4505 (N_4505,N_4384,N_4228);
or U4506 (N_4506,N_4277,N_4224);
and U4507 (N_4507,N_4326,N_4302);
nor U4508 (N_4508,N_4319,N_4310);
or U4509 (N_4509,N_4302,N_4276);
or U4510 (N_4510,N_4328,N_4324);
nand U4511 (N_4511,N_4380,N_4398);
nor U4512 (N_4512,N_4263,N_4206);
nand U4513 (N_4513,N_4232,N_4361);
nand U4514 (N_4514,N_4244,N_4371);
nand U4515 (N_4515,N_4271,N_4253);
nor U4516 (N_4516,N_4205,N_4277);
xnor U4517 (N_4517,N_4395,N_4264);
or U4518 (N_4518,N_4289,N_4360);
nor U4519 (N_4519,N_4298,N_4337);
or U4520 (N_4520,N_4329,N_4394);
or U4521 (N_4521,N_4268,N_4373);
xnor U4522 (N_4522,N_4236,N_4243);
and U4523 (N_4523,N_4352,N_4353);
or U4524 (N_4524,N_4274,N_4220);
xnor U4525 (N_4525,N_4321,N_4264);
and U4526 (N_4526,N_4286,N_4222);
nand U4527 (N_4527,N_4240,N_4200);
xnor U4528 (N_4528,N_4397,N_4265);
and U4529 (N_4529,N_4256,N_4311);
and U4530 (N_4530,N_4224,N_4266);
or U4531 (N_4531,N_4246,N_4268);
or U4532 (N_4532,N_4313,N_4242);
and U4533 (N_4533,N_4247,N_4263);
xnor U4534 (N_4534,N_4368,N_4372);
nand U4535 (N_4535,N_4248,N_4398);
xor U4536 (N_4536,N_4347,N_4256);
xnor U4537 (N_4537,N_4249,N_4338);
and U4538 (N_4538,N_4262,N_4287);
xor U4539 (N_4539,N_4361,N_4315);
or U4540 (N_4540,N_4238,N_4294);
nor U4541 (N_4541,N_4349,N_4345);
or U4542 (N_4542,N_4236,N_4213);
xor U4543 (N_4543,N_4387,N_4398);
and U4544 (N_4544,N_4378,N_4288);
or U4545 (N_4545,N_4370,N_4248);
or U4546 (N_4546,N_4329,N_4335);
xor U4547 (N_4547,N_4357,N_4235);
nor U4548 (N_4548,N_4334,N_4307);
nand U4549 (N_4549,N_4311,N_4341);
xnor U4550 (N_4550,N_4320,N_4395);
and U4551 (N_4551,N_4303,N_4377);
xnor U4552 (N_4552,N_4213,N_4389);
or U4553 (N_4553,N_4397,N_4227);
xnor U4554 (N_4554,N_4228,N_4262);
and U4555 (N_4555,N_4350,N_4344);
nor U4556 (N_4556,N_4375,N_4385);
nor U4557 (N_4557,N_4346,N_4307);
and U4558 (N_4558,N_4399,N_4287);
nor U4559 (N_4559,N_4218,N_4225);
nand U4560 (N_4560,N_4294,N_4395);
or U4561 (N_4561,N_4331,N_4223);
or U4562 (N_4562,N_4323,N_4226);
nand U4563 (N_4563,N_4238,N_4295);
or U4564 (N_4564,N_4321,N_4317);
or U4565 (N_4565,N_4385,N_4287);
or U4566 (N_4566,N_4389,N_4279);
nor U4567 (N_4567,N_4251,N_4208);
nor U4568 (N_4568,N_4330,N_4244);
nor U4569 (N_4569,N_4203,N_4229);
and U4570 (N_4570,N_4379,N_4238);
xor U4571 (N_4571,N_4280,N_4259);
nor U4572 (N_4572,N_4312,N_4236);
nand U4573 (N_4573,N_4399,N_4368);
or U4574 (N_4574,N_4305,N_4309);
nor U4575 (N_4575,N_4387,N_4281);
or U4576 (N_4576,N_4210,N_4200);
and U4577 (N_4577,N_4273,N_4369);
nand U4578 (N_4578,N_4270,N_4226);
or U4579 (N_4579,N_4383,N_4311);
or U4580 (N_4580,N_4215,N_4226);
or U4581 (N_4581,N_4378,N_4351);
nand U4582 (N_4582,N_4364,N_4357);
or U4583 (N_4583,N_4392,N_4361);
and U4584 (N_4584,N_4392,N_4267);
nor U4585 (N_4585,N_4209,N_4250);
and U4586 (N_4586,N_4226,N_4207);
and U4587 (N_4587,N_4263,N_4323);
xor U4588 (N_4588,N_4370,N_4200);
and U4589 (N_4589,N_4289,N_4333);
nand U4590 (N_4590,N_4364,N_4278);
nor U4591 (N_4591,N_4339,N_4217);
nand U4592 (N_4592,N_4302,N_4215);
nand U4593 (N_4593,N_4216,N_4214);
nand U4594 (N_4594,N_4315,N_4256);
or U4595 (N_4595,N_4297,N_4310);
and U4596 (N_4596,N_4228,N_4311);
nand U4597 (N_4597,N_4334,N_4316);
nand U4598 (N_4598,N_4214,N_4255);
nand U4599 (N_4599,N_4374,N_4369);
nor U4600 (N_4600,N_4427,N_4468);
nor U4601 (N_4601,N_4437,N_4584);
and U4602 (N_4602,N_4500,N_4570);
nand U4603 (N_4603,N_4535,N_4475);
xnor U4604 (N_4604,N_4477,N_4435);
xor U4605 (N_4605,N_4483,N_4403);
xnor U4606 (N_4606,N_4506,N_4471);
and U4607 (N_4607,N_4556,N_4514);
and U4608 (N_4608,N_4488,N_4561);
nand U4609 (N_4609,N_4515,N_4452);
or U4610 (N_4610,N_4441,N_4461);
or U4611 (N_4611,N_4557,N_4428);
xor U4612 (N_4612,N_4594,N_4432);
or U4613 (N_4613,N_4577,N_4495);
nand U4614 (N_4614,N_4578,N_4402);
nor U4615 (N_4615,N_4543,N_4559);
or U4616 (N_4616,N_4558,N_4498);
nor U4617 (N_4617,N_4569,N_4587);
nor U4618 (N_4618,N_4502,N_4491);
nand U4619 (N_4619,N_4479,N_4534);
and U4620 (N_4620,N_4512,N_4451);
nand U4621 (N_4621,N_4473,N_4522);
nor U4622 (N_4622,N_4467,N_4472);
xor U4623 (N_4623,N_4423,N_4519);
or U4624 (N_4624,N_4419,N_4417);
or U4625 (N_4625,N_4484,N_4444);
and U4626 (N_4626,N_4540,N_4576);
and U4627 (N_4627,N_4497,N_4562);
xnor U4628 (N_4628,N_4529,N_4548);
nand U4629 (N_4629,N_4518,N_4593);
xnor U4630 (N_4630,N_4538,N_4589);
or U4631 (N_4631,N_4412,N_4455);
xnor U4632 (N_4632,N_4517,N_4406);
xnor U4633 (N_4633,N_4436,N_4504);
xnor U4634 (N_4634,N_4575,N_4418);
or U4635 (N_4635,N_4501,N_4553);
nor U4636 (N_4636,N_4521,N_4454);
or U4637 (N_4637,N_4499,N_4541);
nand U4638 (N_4638,N_4401,N_4446);
nor U4639 (N_4639,N_4460,N_4490);
or U4640 (N_4640,N_4598,N_4542);
or U4641 (N_4641,N_4592,N_4431);
or U4642 (N_4642,N_4516,N_4456);
or U4643 (N_4643,N_4599,N_4448);
or U4644 (N_4644,N_4554,N_4469);
or U4645 (N_4645,N_4486,N_4413);
nor U4646 (N_4646,N_4574,N_4595);
nor U4647 (N_4647,N_4466,N_4430);
nor U4648 (N_4648,N_4583,N_4416);
and U4649 (N_4649,N_4474,N_4462);
nor U4650 (N_4650,N_4410,N_4588);
nor U4651 (N_4651,N_4533,N_4513);
xnor U4652 (N_4652,N_4508,N_4586);
or U4653 (N_4653,N_4404,N_4450);
nand U4654 (N_4654,N_4503,N_4581);
and U4655 (N_4655,N_4480,N_4414);
nand U4656 (N_4656,N_4549,N_4447);
xnor U4657 (N_4657,N_4492,N_4550);
or U4658 (N_4658,N_4568,N_4579);
xnor U4659 (N_4659,N_4596,N_4457);
nand U4660 (N_4660,N_4470,N_4573);
nand U4661 (N_4661,N_4482,N_4433);
nand U4662 (N_4662,N_4421,N_4453);
and U4663 (N_4663,N_4571,N_4537);
nor U4664 (N_4664,N_4458,N_4425);
nand U4665 (N_4665,N_4563,N_4439);
or U4666 (N_4666,N_4411,N_4400);
and U4667 (N_4667,N_4478,N_4438);
xor U4668 (N_4668,N_4539,N_4551);
nor U4669 (N_4669,N_4509,N_4565);
nand U4670 (N_4670,N_4405,N_4505);
or U4671 (N_4671,N_4572,N_4426);
and U4672 (N_4672,N_4567,N_4552);
and U4673 (N_4673,N_4532,N_4442);
xnor U4674 (N_4674,N_4528,N_4481);
xor U4675 (N_4675,N_4546,N_4485);
or U4676 (N_4676,N_4429,N_4424);
xnor U4677 (N_4677,N_4564,N_4531);
and U4678 (N_4678,N_4524,N_4510);
or U4679 (N_4679,N_4597,N_4489);
xor U4680 (N_4680,N_4465,N_4523);
nor U4681 (N_4681,N_4525,N_4590);
xnor U4682 (N_4682,N_4544,N_4487);
xor U4683 (N_4683,N_4494,N_4420);
nor U4684 (N_4684,N_4496,N_4422);
or U4685 (N_4685,N_4507,N_4415);
xor U4686 (N_4686,N_4555,N_4545);
nor U4687 (N_4687,N_4511,N_4434);
and U4688 (N_4688,N_4407,N_4526);
and U4689 (N_4689,N_4530,N_4520);
nand U4690 (N_4690,N_4585,N_4443);
nor U4691 (N_4691,N_4591,N_4409);
and U4692 (N_4692,N_4560,N_4445);
nor U4693 (N_4693,N_4440,N_4527);
nand U4694 (N_4694,N_4463,N_4476);
or U4695 (N_4695,N_4580,N_4464);
and U4696 (N_4696,N_4408,N_4459);
xnor U4697 (N_4697,N_4493,N_4582);
and U4698 (N_4698,N_4547,N_4449);
and U4699 (N_4699,N_4566,N_4536);
nor U4700 (N_4700,N_4471,N_4584);
and U4701 (N_4701,N_4481,N_4521);
or U4702 (N_4702,N_4574,N_4535);
nor U4703 (N_4703,N_4402,N_4500);
nor U4704 (N_4704,N_4486,N_4592);
nor U4705 (N_4705,N_4595,N_4493);
nor U4706 (N_4706,N_4533,N_4553);
nor U4707 (N_4707,N_4496,N_4411);
or U4708 (N_4708,N_4595,N_4413);
nand U4709 (N_4709,N_4431,N_4415);
xnor U4710 (N_4710,N_4558,N_4593);
xnor U4711 (N_4711,N_4407,N_4460);
nor U4712 (N_4712,N_4594,N_4444);
or U4713 (N_4713,N_4403,N_4444);
nand U4714 (N_4714,N_4536,N_4563);
nor U4715 (N_4715,N_4462,N_4421);
xor U4716 (N_4716,N_4557,N_4497);
nand U4717 (N_4717,N_4518,N_4538);
nor U4718 (N_4718,N_4556,N_4418);
nand U4719 (N_4719,N_4500,N_4579);
nor U4720 (N_4720,N_4405,N_4490);
nor U4721 (N_4721,N_4502,N_4549);
and U4722 (N_4722,N_4587,N_4526);
nor U4723 (N_4723,N_4518,N_4498);
xor U4724 (N_4724,N_4418,N_4480);
nor U4725 (N_4725,N_4486,N_4577);
xor U4726 (N_4726,N_4427,N_4470);
and U4727 (N_4727,N_4480,N_4478);
or U4728 (N_4728,N_4432,N_4409);
xor U4729 (N_4729,N_4484,N_4434);
nand U4730 (N_4730,N_4408,N_4516);
nand U4731 (N_4731,N_4572,N_4424);
xor U4732 (N_4732,N_4501,N_4492);
xnor U4733 (N_4733,N_4539,N_4544);
xor U4734 (N_4734,N_4527,N_4505);
xnor U4735 (N_4735,N_4543,N_4466);
nand U4736 (N_4736,N_4437,N_4450);
xor U4737 (N_4737,N_4538,N_4411);
nor U4738 (N_4738,N_4419,N_4422);
xor U4739 (N_4739,N_4580,N_4417);
or U4740 (N_4740,N_4435,N_4594);
xor U4741 (N_4741,N_4453,N_4435);
nand U4742 (N_4742,N_4430,N_4483);
nor U4743 (N_4743,N_4468,N_4481);
or U4744 (N_4744,N_4473,N_4402);
or U4745 (N_4745,N_4473,N_4536);
xor U4746 (N_4746,N_4475,N_4492);
xor U4747 (N_4747,N_4490,N_4543);
xor U4748 (N_4748,N_4567,N_4556);
or U4749 (N_4749,N_4586,N_4472);
xor U4750 (N_4750,N_4400,N_4440);
xor U4751 (N_4751,N_4542,N_4574);
or U4752 (N_4752,N_4523,N_4409);
nand U4753 (N_4753,N_4403,N_4493);
nand U4754 (N_4754,N_4577,N_4557);
or U4755 (N_4755,N_4540,N_4429);
or U4756 (N_4756,N_4486,N_4456);
xnor U4757 (N_4757,N_4584,N_4549);
xnor U4758 (N_4758,N_4499,N_4496);
xnor U4759 (N_4759,N_4494,N_4568);
or U4760 (N_4760,N_4498,N_4505);
xnor U4761 (N_4761,N_4513,N_4503);
nand U4762 (N_4762,N_4470,N_4489);
and U4763 (N_4763,N_4550,N_4499);
or U4764 (N_4764,N_4465,N_4437);
nand U4765 (N_4765,N_4573,N_4575);
xor U4766 (N_4766,N_4554,N_4485);
or U4767 (N_4767,N_4451,N_4476);
and U4768 (N_4768,N_4555,N_4513);
or U4769 (N_4769,N_4477,N_4453);
xnor U4770 (N_4770,N_4455,N_4449);
nand U4771 (N_4771,N_4454,N_4485);
and U4772 (N_4772,N_4531,N_4442);
xnor U4773 (N_4773,N_4440,N_4572);
nand U4774 (N_4774,N_4500,N_4530);
and U4775 (N_4775,N_4569,N_4596);
nor U4776 (N_4776,N_4596,N_4495);
xnor U4777 (N_4777,N_4495,N_4581);
and U4778 (N_4778,N_4552,N_4442);
nor U4779 (N_4779,N_4524,N_4420);
or U4780 (N_4780,N_4457,N_4506);
xnor U4781 (N_4781,N_4579,N_4484);
xnor U4782 (N_4782,N_4473,N_4476);
or U4783 (N_4783,N_4415,N_4564);
and U4784 (N_4784,N_4545,N_4548);
or U4785 (N_4785,N_4497,N_4445);
nand U4786 (N_4786,N_4535,N_4569);
nor U4787 (N_4787,N_4418,N_4403);
or U4788 (N_4788,N_4482,N_4468);
and U4789 (N_4789,N_4564,N_4409);
and U4790 (N_4790,N_4430,N_4477);
xor U4791 (N_4791,N_4506,N_4591);
nand U4792 (N_4792,N_4489,N_4419);
nand U4793 (N_4793,N_4408,N_4513);
and U4794 (N_4794,N_4437,N_4579);
xnor U4795 (N_4795,N_4597,N_4487);
or U4796 (N_4796,N_4465,N_4438);
nand U4797 (N_4797,N_4458,N_4555);
nor U4798 (N_4798,N_4441,N_4447);
or U4799 (N_4799,N_4487,N_4480);
nand U4800 (N_4800,N_4692,N_4757);
nor U4801 (N_4801,N_4751,N_4752);
and U4802 (N_4802,N_4766,N_4618);
nand U4803 (N_4803,N_4672,N_4638);
xnor U4804 (N_4804,N_4755,N_4625);
and U4805 (N_4805,N_4743,N_4785);
xor U4806 (N_4806,N_4714,N_4771);
nand U4807 (N_4807,N_4654,N_4601);
or U4808 (N_4808,N_4607,N_4648);
nand U4809 (N_4809,N_4762,N_4649);
nand U4810 (N_4810,N_4687,N_4790);
nand U4811 (N_4811,N_4716,N_4722);
nand U4812 (N_4812,N_4622,N_4665);
or U4813 (N_4813,N_4764,N_4663);
and U4814 (N_4814,N_4783,N_4781);
nor U4815 (N_4815,N_4754,N_4736);
xor U4816 (N_4816,N_4688,N_4697);
xnor U4817 (N_4817,N_4698,N_4765);
nor U4818 (N_4818,N_4702,N_4711);
xor U4819 (N_4819,N_4720,N_4729);
or U4820 (N_4820,N_4763,N_4701);
and U4821 (N_4821,N_4627,N_4675);
or U4822 (N_4822,N_4680,N_4749);
and U4823 (N_4823,N_4619,N_4655);
nand U4824 (N_4824,N_4776,N_4778);
or U4825 (N_4825,N_4700,N_4636);
nor U4826 (N_4826,N_4773,N_4658);
or U4827 (N_4827,N_4794,N_4769);
nor U4828 (N_4828,N_4721,N_4617);
nand U4829 (N_4829,N_4793,N_4728);
xor U4830 (N_4830,N_4632,N_4661);
or U4831 (N_4831,N_4774,N_4691);
nand U4832 (N_4832,N_4685,N_4624);
or U4833 (N_4833,N_4727,N_4719);
nor U4834 (N_4834,N_4657,N_4696);
xnor U4835 (N_4835,N_4730,N_4626);
and U4836 (N_4836,N_4643,N_4713);
xor U4837 (N_4837,N_4671,N_4613);
xnor U4838 (N_4838,N_4640,N_4786);
or U4839 (N_4839,N_4628,N_4637);
or U4840 (N_4840,N_4792,N_4726);
xnor U4841 (N_4841,N_4686,N_4784);
or U4842 (N_4842,N_4779,N_4789);
nor U4843 (N_4843,N_4760,N_4767);
nor U4844 (N_4844,N_4695,N_4735);
xnor U4845 (N_4845,N_4642,N_4761);
xor U4846 (N_4846,N_4746,N_4740);
nor U4847 (N_4847,N_4758,N_4679);
or U4848 (N_4848,N_4709,N_4724);
or U4849 (N_4849,N_4768,N_4739);
xor U4850 (N_4850,N_4662,N_4699);
and U4851 (N_4851,N_4689,N_4667);
xor U4852 (N_4852,N_4704,N_4731);
or U4853 (N_4853,N_4710,N_4602);
or U4854 (N_4854,N_4775,N_4707);
nand U4855 (N_4855,N_4718,N_4635);
or U4856 (N_4856,N_4623,N_4693);
or U4857 (N_4857,N_4703,N_4633);
nor U4858 (N_4858,N_4742,N_4690);
nor U4859 (N_4859,N_4741,N_4608);
nor U4860 (N_4860,N_4644,N_4777);
xor U4861 (N_4861,N_4631,N_4606);
xor U4862 (N_4862,N_4629,N_4744);
and U4863 (N_4863,N_4603,N_4694);
nor U4864 (N_4864,N_4734,N_4634);
nand U4865 (N_4865,N_4674,N_4616);
xnor U4866 (N_4866,N_4670,N_4610);
nor U4867 (N_4867,N_4798,N_4600);
or U4868 (N_4868,N_4673,N_4782);
xor U4869 (N_4869,N_4615,N_4770);
xor U4870 (N_4870,N_4641,N_4723);
nand U4871 (N_4871,N_4605,N_4630);
or U4872 (N_4872,N_4659,N_4677);
xnor U4873 (N_4873,N_4604,N_4668);
or U4874 (N_4874,N_4780,N_4748);
or U4875 (N_4875,N_4791,N_4614);
nor U4876 (N_4876,N_4708,N_4620);
nor U4877 (N_4877,N_4797,N_4650);
xnor U4878 (N_4878,N_4664,N_4611);
nand U4879 (N_4879,N_4609,N_4717);
nand U4880 (N_4880,N_4795,N_4621);
nor U4881 (N_4881,N_4759,N_4646);
nor U4882 (N_4882,N_4683,N_4682);
nand U4883 (N_4883,N_4725,N_4750);
xnor U4884 (N_4884,N_4753,N_4684);
nor U4885 (N_4885,N_4737,N_4660);
nand U4886 (N_4886,N_4732,N_4656);
or U4887 (N_4887,N_4799,N_4681);
or U4888 (N_4888,N_4676,N_4666);
or U4889 (N_4889,N_4745,N_4645);
xnor U4890 (N_4890,N_4738,N_4706);
nand U4891 (N_4891,N_4712,N_4678);
xnor U4892 (N_4892,N_4639,N_4669);
nand U4893 (N_4893,N_4788,N_4652);
xnor U4894 (N_4894,N_4733,N_4653);
xnor U4895 (N_4895,N_4756,N_4796);
nor U4896 (N_4896,N_4705,N_4747);
or U4897 (N_4897,N_4612,N_4715);
xnor U4898 (N_4898,N_4651,N_4787);
xor U4899 (N_4899,N_4647,N_4772);
xor U4900 (N_4900,N_4720,N_4690);
nor U4901 (N_4901,N_4727,N_4765);
xor U4902 (N_4902,N_4784,N_4705);
nand U4903 (N_4903,N_4655,N_4763);
and U4904 (N_4904,N_4633,N_4731);
and U4905 (N_4905,N_4695,N_4716);
nand U4906 (N_4906,N_4671,N_4742);
or U4907 (N_4907,N_4690,N_4670);
xor U4908 (N_4908,N_4776,N_4642);
nand U4909 (N_4909,N_4643,N_4690);
or U4910 (N_4910,N_4780,N_4659);
nor U4911 (N_4911,N_4661,N_4693);
or U4912 (N_4912,N_4768,N_4623);
nand U4913 (N_4913,N_4648,N_4720);
nand U4914 (N_4914,N_4621,N_4796);
and U4915 (N_4915,N_4792,N_4676);
nand U4916 (N_4916,N_4753,N_4762);
and U4917 (N_4917,N_4782,N_4768);
and U4918 (N_4918,N_4681,N_4780);
xnor U4919 (N_4919,N_4610,N_4674);
or U4920 (N_4920,N_4733,N_4766);
and U4921 (N_4921,N_4600,N_4728);
xor U4922 (N_4922,N_4773,N_4662);
and U4923 (N_4923,N_4753,N_4621);
nand U4924 (N_4924,N_4674,N_4765);
and U4925 (N_4925,N_4791,N_4714);
nand U4926 (N_4926,N_4796,N_4777);
xnor U4927 (N_4927,N_4712,N_4720);
and U4928 (N_4928,N_4778,N_4720);
xnor U4929 (N_4929,N_4767,N_4623);
or U4930 (N_4930,N_4791,N_4744);
or U4931 (N_4931,N_4659,N_4799);
nand U4932 (N_4932,N_4650,N_4649);
nor U4933 (N_4933,N_4662,N_4665);
or U4934 (N_4934,N_4777,N_4760);
nand U4935 (N_4935,N_4650,N_4700);
and U4936 (N_4936,N_4620,N_4784);
and U4937 (N_4937,N_4695,N_4606);
xor U4938 (N_4938,N_4775,N_4692);
xor U4939 (N_4939,N_4641,N_4785);
nand U4940 (N_4940,N_4683,N_4693);
xor U4941 (N_4941,N_4781,N_4727);
nor U4942 (N_4942,N_4619,N_4688);
xor U4943 (N_4943,N_4753,N_4635);
or U4944 (N_4944,N_4754,N_4620);
or U4945 (N_4945,N_4757,N_4689);
and U4946 (N_4946,N_4685,N_4661);
nand U4947 (N_4947,N_4764,N_4667);
and U4948 (N_4948,N_4660,N_4673);
xnor U4949 (N_4949,N_4737,N_4717);
or U4950 (N_4950,N_4779,N_4755);
nand U4951 (N_4951,N_4677,N_4692);
nor U4952 (N_4952,N_4618,N_4643);
and U4953 (N_4953,N_4698,N_4734);
and U4954 (N_4954,N_4785,N_4616);
nand U4955 (N_4955,N_4731,N_4700);
xor U4956 (N_4956,N_4777,N_4665);
or U4957 (N_4957,N_4746,N_4669);
nor U4958 (N_4958,N_4614,N_4792);
nor U4959 (N_4959,N_4603,N_4645);
nor U4960 (N_4960,N_4708,N_4601);
or U4961 (N_4961,N_4649,N_4774);
or U4962 (N_4962,N_4751,N_4633);
nor U4963 (N_4963,N_4708,N_4656);
nand U4964 (N_4964,N_4759,N_4631);
xnor U4965 (N_4965,N_4691,N_4658);
nor U4966 (N_4966,N_4735,N_4711);
or U4967 (N_4967,N_4760,N_4757);
and U4968 (N_4968,N_4684,N_4728);
nor U4969 (N_4969,N_4654,N_4628);
nor U4970 (N_4970,N_4707,N_4778);
nand U4971 (N_4971,N_4680,N_4691);
or U4972 (N_4972,N_4783,N_4754);
nor U4973 (N_4973,N_4790,N_4724);
nand U4974 (N_4974,N_4739,N_4725);
nor U4975 (N_4975,N_4783,N_4740);
or U4976 (N_4976,N_4721,N_4717);
and U4977 (N_4977,N_4692,N_4750);
xor U4978 (N_4978,N_4607,N_4741);
nand U4979 (N_4979,N_4620,N_4647);
nor U4980 (N_4980,N_4657,N_4787);
nor U4981 (N_4981,N_4737,N_4606);
nor U4982 (N_4982,N_4629,N_4797);
xnor U4983 (N_4983,N_4788,N_4734);
xnor U4984 (N_4984,N_4654,N_4744);
xnor U4985 (N_4985,N_4651,N_4762);
or U4986 (N_4986,N_4755,N_4639);
and U4987 (N_4987,N_4625,N_4739);
nand U4988 (N_4988,N_4705,N_4778);
and U4989 (N_4989,N_4757,N_4627);
nor U4990 (N_4990,N_4619,N_4778);
xnor U4991 (N_4991,N_4637,N_4653);
nand U4992 (N_4992,N_4605,N_4793);
xnor U4993 (N_4993,N_4612,N_4797);
and U4994 (N_4994,N_4795,N_4604);
nor U4995 (N_4995,N_4669,N_4742);
nand U4996 (N_4996,N_4669,N_4726);
xor U4997 (N_4997,N_4664,N_4701);
xor U4998 (N_4998,N_4710,N_4631);
xor U4999 (N_4999,N_4708,N_4751);
or U5000 (N_5000,N_4821,N_4915);
nand U5001 (N_5001,N_4833,N_4902);
nand U5002 (N_5002,N_4993,N_4802);
and U5003 (N_5003,N_4886,N_4817);
and U5004 (N_5004,N_4986,N_4848);
or U5005 (N_5005,N_4871,N_4892);
nand U5006 (N_5006,N_4983,N_4859);
or U5007 (N_5007,N_4942,N_4846);
nor U5008 (N_5008,N_4836,N_4861);
xor U5009 (N_5009,N_4988,N_4815);
and U5010 (N_5010,N_4837,N_4864);
or U5011 (N_5011,N_4933,N_4858);
nor U5012 (N_5012,N_4998,N_4877);
and U5013 (N_5013,N_4956,N_4926);
nor U5014 (N_5014,N_4995,N_4894);
and U5015 (N_5015,N_4854,N_4899);
and U5016 (N_5016,N_4873,N_4925);
or U5017 (N_5017,N_4984,N_4826);
or U5018 (N_5018,N_4967,N_4876);
or U5019 (N_5019,N_4945,N_4985);
xnor U5020 (N_5020,N_4830,N_4870);
and U5021 (N_5021,N_4869,N_4906);
xor U5022 (N_5022,N_4808,N_4816);
nand U5023 (N_5023,N_4843,N_4951);
nor U5024 (N_5024,N_4818,N_4936);
and U5025 (N_5025,N_4874,N_4857);
nor U5026 (N_5026,N_4934,N_4944);
or U5027 (N_5027,N_4928,N_4914);
xnor U5028 (N_5028,N_4987,N_4883);
and U5029 (N_5029,N_4992,N_4994);
and U5030 (N_5030,N_4810,N_4852);
nand U5031 (N_5031,N_4980,N_4800);
or U5032 (N_5032,N_4975,N_4989);
nand U5033 (N_5033,N_4882,N_4964);
or U5034 (N_5034,N_4913,N_4943);
nor U5035 (N_5035,N_4901,N_4827);
nand U5036 (N_5036,N_4890,N_4960);
or U5037 (N_5037,N_4841,N_4898);
nor U5038 (N_5038,N_4904,N_4855);
nand U5039 (N_5039,N_4820,N_4955);
or U5040 (N_5040,N_4961,N_4813);
nor U5041 (N_5041,N_4842,N_4863);
or U5042 (N_5042,N_4805,N_4812);
and U5043 (N_5043,N_4916,N_4949);
and U5044 (N_5044,N_4979,N_4959);
and U5045 (N_5045,N_4946,N_4909);
nor U5046 (N_5046,N_4968,N_4974);
nor U5047 (N_5047,N_4811,N_4908);
and U5048 (N_5048,N_4911,N_4977);
or U5049 (N_5049,N_4875,N_4880);
and U5050 (N_5050,N_4862,N_4912);
or U5051 (N_5051,N_4895,N_4900);
and U5052 (N_5052,N_4844,N_4929);
nand U5053 (N_5053,N_4840,N_4803);
nand U5054 (N_5054,N_4860,N_4825);
or U5055 (N_5055,N_4918,N_4937);
and U5056 (N_5056,N_4990,N_4919);
nor U5057 (N_5057,N_4966,N_4930);
and U5058 (N_5058,N_4982,N_4896);
nand U5059 (N_5059,N_4927,N_4973);
and U5060 (N_5060,N_4903,N_4872);
xor U5061 (N_5061,N_4976,N_4828);
xor U5062 (N_5062,N_4958,N_4878);
nor U5063 (N_5063,N_4981,N_4935);
nand U5064 (N_5064,N_4962,N_4822);
nand U5065 (N_5065,N_4807,N_4887);
nand U5066 (N_5066,N_4856,N_4917);
xnor U5067 (N_5067,N_4845,N_4885);
nand U5068 (N_5068,N_4865,N_4963);
nor U5069 (N_5069,N_4868,N_4835);
or U5070 (N_5070,N_4851,N_4938);
nor U5071 (N_5071,N_4997,N_4867);
and U5072 (N_5072,N_4965,N_4823);
nor U5073 (N_5073,N_4970,N_4999);
xor U5074 (N_5074,N_4931,N_4957);
or U5075 (N_5075,N_4923,N_4953);
or U5076 (N_5076,N_4801,N_4839);
xnor U5077 (N_5077,N_4847,N_4806);
or U5078 (N_5078,N_4905,N_4850);
or U5079 (N_5079,N_4907,N_4971);
nand U5080 (N_5080,N_4996,N_4814);
nand U5081 (N_5081,N_4950,N_4952);
or U5082 (N_5082,N_4881,N_4819);
nand U5083 (N_5083,N_4978,N_4804);
or U5084 (N_5084,N_4866,N_4884);
or U5085 (N_5085,N_4891,N_4939);
and U5086 (N_5086,N_4829,N_4991);
or U5087 (N_5087,N_4897,N_4954);
nor U5088 (N_5088,N_4889,N_4910);
xnor U5089 (N_5089,N_4969,N_4853);
nor U5090 (N_5090,N_4893,N_4831);
nor U5091 (N_5091,N_4824,N_4924);
or U5092 (N_5092,N_4948,N_4832);
or U5093 (N_5093,N_4940,N_4972);
nor U5094 (N_5094,N_4879,N_4922);
xnor U5095 (N_5095,N_4834,N_4941);
nor U5096 (N_5096,N_4920,N_4849);
nor U5097 (N_5097,N_4947,N_4932);
and U5098 (N_5098,N_4838,N_4888);
xor U5099 (N_5099,N_4809,N_4921);
and U5100 (N_5100,N_4917,N_4830);
and U5101 (N_5101,N_4815,N_4957);
or U5102 (N_5102,N_4907,N_4963);
or U5103 (N_5103,N_4917,N_4958);
nand U5104 (N_5104,N_4926,N_4886);
xor U5105 (N_5105,N_4909,N_4824);
and U5106 (N_5106,N_4900,N_4832);
nand U5107 (N_5107,N_4983,N_4951);
xor U5108 (N_5108,N_4822,N_4835);
or U5109 (N_5109,N_4939,N_4937);
xnor U5110 (N_5110,N_4947,N_4981);
xnor U5111 (N_5111,N_4903,N_4917);
or U5112 (N_5112,N_4990,N_4822);
nor U5113 (N_5113,N_4916,N_4994);
and U5114 (N_5114,N_4983,N_4936);
nand U5115 (N_5115,N_4812,N_4866);
or U5116 (N_5116,N_4827,N_4967);
nand U5117 (N_5117,N_4853,N_4985);
nor U5118 (N_5118,N_4954,N_4964);
nand U5119 (N_5119,N_4972,N_4816);
and U5120 (N_5120,N_4856,N_4887);
or U5121 (N_5121,N_4970,N_4943);
nor U5122 (N_5122,N_4801,N_4906);
nor U5123 (N_5123,N_4834,N_4821);
nor U5124 (N_5124,N_4875,N_4824);
xnor U5125 (N_5125,N_4939,N_4916);
and U5126 (N_5126,N_4957,N_4928);
nand U5127 (N_5127,N_4886,N_4965);
nand U5128 (N_5128,N_4810,N_4927);
xnor U5129 (N_5129,N_4988,N_4808);
nand U5130 (N_5130,N_4829,N_4971);
and U5131 (N_5131,N_4938,N_4976);
nand U5132 (N_5132,N_4801,N_4916);
or U5133 (N_5133,N_4945,N_4907);
xor U5134 (N_5134,N_4804,N_4861);
nor U5135 (N_5135,N_4943,N_4954);
and U5136 (N_5136,N_4890,N_4958);
nand U5137 (N_5137,N_4830,N_4915);
nand U5138 (N_5138,N_4861,N_4823);
and U5139 (N_5139,N_4868,N_4914);
xor U5140 (N_5140,N_4901,N_4974);
nand U5141 (N_5141,N_4992,N_4941);
and U5142 (N_5142,N_4909,N_4901);
nand U5143 (N_5143,N_4886,N_4854);
nor U5144 (N_5144,N_4940,N_4907);
xor U5145 (N_5145,N_4860,N_4940);
and U5146 (N_5146,N_4900,N_4874);
or U5147 (N_5147,N_4940,N_4920);
nand U5148 (N_5148,N_4991,N_4930);
and U5149 (N_5149,N_4951,N_4852);
nor U5150 (N_5150,N_4941,N_4866);
nand U5151 (N_5151,N_4853,N_4875);
nand U5152 (N_5152,N_4929,N_4927);
nor U5153 (N_5153,N_4800,N_4904);
or U5154 (N_5154,N_4926,N_4998);
and U5155 (N_5155,N_4898,N_4804);
or U5156 (N_5156,N_4824,N_4853);
or U5157 (N_5157,N_4910,N_4848);
xor U5158 (N_5158,N_4965,N_4928);
nor U5159 (N_5159,N_4888,N_4935);
and U5160 (N_5160,N_4812,N_4995);
or U5161 (N_5161,N_4940,N_4976);
nand U5162 (N_5162,N_4988,N_4990);
and U5163 (N_5163,N_4816,N_4958);
nor U5164 (N_5164,N_4989,N_4822);
nor U5165 (N_5165,N_4960,N_4822);
and U5166 (N_5166,N_4830,N_4901);
and U5167 (N_5167,N_4827,N_4896);
xor U5168 (N_5168,N_4855,N_4997);
xor U5169 (N_5169,N_4900,N_4932);
nor U5170 (N_5170,N_4932,N_4890);
nor U5171 (N_5171,N_4883,N_4864);
xor U5172 (N_5172,N_4860,N_4927);
xnor U5173 (N_5173,N_4953,N_4909);
and U5174 (N_5174,N_4992,N_4816);
xnor U5175 (N_5175,N_4862,N_4857);
or U5176 (N_5176,N_4930,N_4879);
nand U5177 (N_5177,N_4803,N_4873);
and U5178 (N_5178,N_4881,N_4814);
or U5179 (N_5179,N_4939,N_4887);
xor U5180 (N_5180,N_4973,N_4801);
nand U5181 (N_5181,N_4938,N_4982);
nor U5182 (N_5182,N_4902,N_4940);
nand U5183 (N_5183,N_4949,N_4863);
nor U5184 (N_5184,N_4991,N_4843);
or U5185 (N_5185,N_4858,N_4916);
and U5186 (N_5186,N_4927,N_4855);
nor U5187 (N_5187,N_4814,N_4902);
or U5188 (N_5188,N_4950,N_4921);
nor U5189 (N_5189,N_4994,N_4883);
nor U5190 (N_5190,N_4818,N_4885);
or U5191 (N_5191,N_4891,N_4999);
nor U5192 (N_5192,N_4962,N_4914);
nand U5193 (N_5193,N_4981,N_4843);
or U5194 (N_5194,N_4812,N_4903);
and U5195 (N_5195,N_4929,N_4945);
nor U5196 (N_5196,N_4936,N_4829);
and U5197 (N_5197,N_4900,N_4965);
nor U5198 (N_5198,N_4960,N_4895);
or U5199 (N_5199,N_4901,N_4863);
or U5200 (N_5200,N_5150,N_5081);
and U5201 (N_5201,N_5030,N_5161);
and U5202 (N_5202,N_5134,N_5051);
nor U5203 (N_5203,N_5073,N_5152);
nand U5204 (N_5204,N_5164,N_5076);
and U5205 (N_5205,N_5101,N_5086);
nand U5206 (N_5206,N_5003,N_5070);
xnor U5207 (N_5207,N_5050,N_5144);
xnor U5208 (N_5208,N_5140,N_5084);
xnor U5209 (N_5209,N_5099,N_5016);
and U5210 (N_5210,N_5177,N_5008);
nand U5211 (N_5211,N_5172,N_5056);
or U5212 (N_5212,N_5168,N_5021);
nor U5213 (N_5213,N_5107,N_5041);
nand U5214 (N_5214,N_5156,N_5124);
xor U5215 (N_5215,N_5106,N_5136);
or U5216 (N_5216,N_5162,N_5186);
nand U5217 (N_5217,N_5032,N_5179);
and U5218 (N_5218,N_5159,N_5147);
and U5219 (N_5219,N_5115,N_5171);
xor U5220 (N_5220,N_5046,N_5091);
or U5221 (N_5221,N_5113,N_5079);
xor U5222 (N_5222,N_5135,N_5038);
and U5223 (N_5223,N_5065,N_5018);
and U5224 (N_5224,N_5157,N_5042);
nor U5225 (N_5225,N_5154,N_5092);
nor U5226 (N_5226,N_5044,N_5185);
xor U5227 (N_5227,N_5094,N_5075);
or U5228 (N_5228,N_5039,N_5170);
xor U5229 (N_5229,N_5108,N_5000);
and U5230 (N_5230,N_5082,N_5196);
xor U5231 (N_5231,N_5037,N_5045);
nor U5232 (N_5232,N_5035,N_5173);
nand U5233 (N_5233,N_5145,N_5143);
or U5234 (N_5234,N_5013,N_5034);
or U5235 (N_5235,N_5095,N_5176);
and U5236 (N_5236,N_5178,N_5067);
nand U5237 (N_5237,N_5012,N_5011);
or U5238 (N_5238,N_5193,N_5119);
nand U5239 (N_5239,N_5146,N_5111);
nor U5240 (N_5240,N_5175,N_5017);
nor U5241 (N_5241,N_5121,N_5031);
nand U5242 (N_5242,N_5199,N_5110);
and U5243 (N_5243,N_5188,N_5088);
or U5244 (N_5244,N_5160,N_5190);
nand U5245 (N_5245,N_5104,N_5052);
nor U5246 (N_5246,N_5063,N_5090);
xor U5247 (N_5247,N_5112,N_5189);
and U5248 (N_5248,N_5139,N_5182);
xnor U5249 (N_5249,N_5040,N_5049);
nand U5250 (N_5250,N_5130,N_5026);
or U5251 (N_5251,N_5165,N_5151);
nand U5252 (N_5252,N_5006,N_5127);
nor U5253 (N_5253,N_5187,N_5169);
xnor U5254 (N_5254,N_5117,N_5093);
nor U5255 (N_5255,N_5133,N_5128);
nor U5256 (N_5256,N_5005,N_5053);
xor U5257 (N_5257,N_5123,N_5077);
xor U5258 (N_5258,N_5072,N_5071);
nor U5259 (N_5259,N_5001,N_5184);
nand U5260 (N_5260,N_5043,N_5036);
nor U5261 (N_5261,N_5138,N_5033);
or U5262 (N_5262,N_5142,N_5014);
or U5263 (N_5263,N_5167,N_5129);
and U5264 (N_5264,N_5102,N_5183);
and U5265 (N_5265,N_5059,N_5197);
nor U5266 (N_5266,N_5023,N_5089);
xnor U5267 (N_5267,N_5058,N_5149);
or U5268 (N_5268,N_5148,N_5061);
and U5269 (N_5269,N_5181,N_5166);
nand U5270 (N_5270,N_5062,N_5024);
or U5271 (N_5271,N_5007,N_5029);
nand U5272 (N_5272,N_5010,N_5191);
nand U5273 (N_5273,N_5098,N_5192);
nor U5274 (N_5274,N_5158,N_5195);
or U5275 (N_5275,N_5020,N_5132);
and U5276 (N_5276,N_5131,N_5125);
nand U5277 (N_5277,N_5048,N_5153);
nor U5278 (N_5278,N_5120,N_5137);
and U5279 (N_5279,N_5141,N_5078);
and U5280 (N_5280,N_5105,N_5155);
xor U5281 (N_5281,N_5025,N_5163);
or U5282 (N_5282,N_5109,N_5015);
nor U5283 (N_5283,N_5114,N_5097);
and U5284 (N_5284,N_5019,N_5002);
nor U5285 (N_5285,N_5055,N_5080);
and U5286 (N_5286,N_5180,N_5118);
nand U5287 (N_5287,N_5064,N_5004);
or U5288 (N_5288,N_5122,N_5009);
or U5289 (N_5289,N_5022,N_5198);
nor U5290 (N_5290,N_5066,N_5103);
xnor U5291 (N_5291,N_5096,N_5060);
nor U5292 (N_5292,N_5057,N_5100);
or U5293 (N_5293,N_5074,N_5068);
nor U5294 (N_5294,N_5069,N_5028);
nand U5295 (N_5295,N_5116,N_5085);
xnor U5296 (N_5296,N_5174,N_5083);
xor U5297 (N_5297,N_5054,N_5126);
nor U5298 (N_5298,N_5027,N_5047);
or U5299 (N_5299,N_5194,N_5087);
nand U5300 (N_5300,N_5105,N_5089);
or U5301 (N_5301,N_5013,N_5007);
nor U5302 (N_5302,N_5151,N_5021);
nor U5303 (N_5303,N_5199,N_5160);
nor U5304 (N_5304,N_5082,N_5006);
nor U5305 (N_5305,N_5010,N_5007);
nor U5306 (N_5306,N_5131,N_5026);
or U5307 (N_5307,N_5168,N_5135);
nor U5308 (N_5308,N_5081,N_5037);
xor U5309 (N_5309,N_5191,N_5069);
and U5310 (N_5310,N_5166,N_5021);
or U5311 (N_5311,N_5057,N_5058);
or U5312 (N_5312,N_5196,N_5181);
nor U5313 (N_5313,N_5138,N_5113);
xnor U5314 (N_5314,N_5076,N_5132);
nor U5315 (N_5315,N_5092,N_5104);
nor U5316 (N_5316,N_5075,N_5033);
nand U5317 (N_5317,N_5137,N_5076);
nand U5318 (N_5318,N_5108,N_5014);
xor U5319 (N_5319,N_5132,N_5042);
and U5320 (N_5320,N_5053,N_5039);
and U5321 (N_5321,N_5028,N_5040);
nand U5322 (N_5322,N_5176,N_5166);
nand U5323 (N_5323,N_5097,N_5042);
nor U5324 (N_5324,N_5044,N_5151);
xnor U5325 (N_5325,N_5007,N_5111);
or U5326 (N_5326,N_5118,N_5067);
xnor U5327 (N_5327,N_5057,N_5117);
and U5328 (N_5328,N_5010,N_5092);
nand U5329 (N_5329,N_5155,N_5180);
nand U5330 (N_5330,N_5171,N_5070);
xor U5331 (N_5331,N_5008,N_5191);
xor U5332 (N_5332,N_5019,N_5065);
xor U5333 (N_5333,N_5136,N_5041);
and U5334 (N_5334,N_5077,N_5160);
nand U5335 (N_5335,N_5098,N_5022);
nand U5336 (N_5336,N_5147,N_5146);
nand U5337 (N_5337,N_5117,N_5052);
nor U5338 (N_5338,N_5109,N_5007);
and U5339 (N_5339,N_5174,N_5165);
xor U5340 (N_5340,N_5187,N_5194);
nand U5341 (N_5341,N_5186,N_5138);
and U5342 (N_5342,N_5126,N_5067);
or U5343 (N_5343,N_5036,N_5153);
and U5344 (N_5344,N_5185,N_5147);
nor U5345 (N_5345,N_5028,N_5141);
xnor U5346 (N_5346,N_5116,N_5047);
xnor U5347 (N_5347,N_5046,N_5116);
or U5348 (N_5348,N_5087,N_5075);
nor U5349 (N_5349,N_5058,N_5025);
nor U5350 (N_5350,N_5181,N_5077);
and U5351 (N_5351,N_5112,N_5013);
nand U5352 (N_5352,N_5161,N_5087);
nor U5353 (N_5353,N_5037,N_5006);
xor U5354 (N_5354,N_5123,N_5149);
nand U5355 (N_5355,N_5026,N_5019);
nor U5356 (N_5356,N_5098,N_5057);
nor U5357 (N_5357,N_5044,N_5031);
or U5358 (N_5358,N_5121,N_5127);
or U5359 (N_5359,N_5053,N_5022);
and U5360 (N_5360,N_5090,N_5060);
and U5361 (N_5361,N_5081,N_5146);
and U5362 (N_5362,N_5144,N_5124);
and U5363 (N_5363,N_5099,N_5062);
and U5364 (N_5364,N_5091,N_5170);
nand U5365 (N_5365,N_5033,N_5179);
nand U5366 (N_5366,N_5123,N_5006);
and U5367 (N_5367,N_5190,N_5185);
nor U5368 (N_5368,N_5141,N_5066);
and U5369 (N_5369,N_5048,N_5005);
nor U5370 (N_5370,N_5152,N_5090);
nor U5371 (N_5371,N_5044,N_5072);
xnor U5372 (N_5372,N_5191,N_5054);
nand U5373 (N_5373,N_5019,N_5044);
nor U5374 (N_5374,N_5116,N_5011);
xnor U5375 (N_5375,N_5124,N_5152);
or U5376 (N_5376,N_5138,N_5129);
nor U5377 (N_5377,N_5192,N_5169);
nor U5378 (N_5378,N_5189,N_5046);
nor U5379 (N_5379,N_5182,N_5025);
and U5380 (N_5380,N_5096,N_5145);
and U5381 (N_5381,N_5011,N_5110);
xnor U5382 (N_5382,N_5097,N_5190);
xnor U5383 (N_5383,N_5020,N_5130);
nor U5384 (N_5384,N_5110,N_5196);
and U5385 (N_5385,N_5070,N_5063);
nand U5386 (N_5386,N_5160,N_5043);
xnor U5387 (N_5387,N_5040,N_5133);
nand U5388 (N_5388,N_5043,N_5181);
nand U5389 (N_5389,N_5096,N_5135);
and U5390 (N_5390,N_5028,N_5068);
or U5391 (N_5391,N_5027,N_5105);
nor U5392 (N_5392,N_5180,N_5191);
xnor U5393 (N_5393,N_5074,N_5080);
or U5394 (N_5394,N_5112,N_5180);
xnor U5395 (N_5395,N_5124,N_5130);
and U5396 (N_5396,N_5093,N_5171);
nor U5397 (N_5397,N_5040,N_5138);
or U5398 (N_5398,N_5009,N_5110);
nand U5399 (N_5399,N_5071,N_5000);
nand U5400 (N_5400,N_5332,N_5212);
or U5401 (N_5401,N_5257,N_5364);
nor U5402 (N_5402,N_5256,N_5301);
or U5403 (N_5403,N_5297,N_5389);
nand U5404 (N_5404,N_5219,N_5233);
nand U5405 (N_5405,N_5320,N_5341);
xnor U5406 (N_5406,N_5308,N_5342);
xor U5407 (N_5407,N_5246,N_5281);
nor U5408 (N_5408,N_5296,N_5350);
nor U5409 (N_5409,N_5238,N_5226);
nand U5410 (N_5410,N_5357,N_5244);
and U5411 (N_5411,N_5227,N_5280);
and U5412 (N_5412,N_5351,N_5339);
xnor U5413 (N_5413,N_5265,N_5326);
xnor U5414 (N_5414,N_5269,N_5287);
xor U5415 (N_5415,N_5385,N_5220);
xor U5416 (N_5416,N_5217,N_5271);
or U5417 (N_5417,N_5239,N_5295);
nor U5418 (N_5418,N_5333,N_5231);
nor U5419 (N_5419,N_5316,N_5282);
and U5420 (N_5420,N_5209,N_5312);
xnor U5421 (N_5421,N_5254,N_5381);
xor U5422 (N_5422,N_5386,N_5262);
or U5423 (N_5423,N_5223,N_5345);
nand U5424 (N_5424,N_5234,N_5362);
nand U5425 (N_5425,N_5348,N_5236);
nor U5426 (N_5426,N_5277,N_5328);
xnor U5427 (N_5427,N_5336,N_5298);
and U5428 (N_5428,N_5398,N_5330);
nand U5429 (N_5429,N_5285,N_5208);
nor U5430 (N_5430,N_5365,N_5360);
nand U5431 (N_5431,N_5371,N_5384);
or U5432 (N_5432,N_5275,N_5214);
nand U5433 (N_5433,N_5396,N_5253);
or U5434 (N_5434,N_5374,N_5379);
xor U5435 (N_5435,N_5200,N_5340);
nand U5436 (N_5436,N_5225,N_5318);
or U5437 (N_5437,N_5211,N_5272);
xor U5438 (N_5438,N_5321,N_5358);
and U5439 (N_5439,N_5395,N_5367);
xnor U5440 (N_5440,N_5309,N_5354);
nand U5441 (N_5441,N_5329,N_5268);
or U5442 (N_5442,N_5240,N_5352);
or U5443 (N_5443,N_5390,N_5278);
or U5444 (N_5444,N_5222,N_5324);
nor U5445 (N_5445,N_5288,N_5243);
nor U5446 (N_5446,N_5270,N_5274);
nor U5447 (N_5447,N_5286,N_5300);
xor U5448 (N_5448,N_5224,N_5302);
xnor U5449 (N_5449,N_5306,N_5313);
and U5450 (N_5450,N_5393,N_5292);
or U5451 (N_5451,N_5303,N_5361);
or U5452 (N_5452,N_5215,N_5378);
xnor U5453 (N_5453,N_5338,N_5279);
nand U5454 (N_5454,N_5264,N_5369);
xnor U5455 (N_5455,N_5377,N_5237);
xor U5456 (N_5456,N_5334,N_5387);
nor U5457 (N_5457,N_5251,N_5353);
nor U5458 (N_5458,N_5213,N_5346);
or U5459 (N_5459,N_5310,N_5261);
xor U5460 (N_5460,N_5299,N_5291);
or U5461 (N_5461,N_5383,N_5229);
nor U5462 (N_5462,N_5373,N_5221);
nor U5463 (N_5463,N_5397,N_5245);
nand U5464 (N_5464,N_5356,N_5266);
xor U5465 (N_5465,N_5355,N_5205);
nor U5466 (N_5466,N_5323,N_5230);
and U5467 (N_5467,N_5289,N_5210);
nand U5468 (N_5468,N_5325,N_5366);
nor U5469 (N_5469,N_5276,N_5207);
xnor U5470 (N_5470,N_5392,N_5347);
xnor U5471 (N_5471,N_5283,N_5273);
nor U5472 (N_5472,N_5370,N_5304);
and U5473 (N_5473,N_5327,N_5203);
nor U5474 (N_5474,N_5259,N_5248);
or U5475 (N_5475,N_5368,N_5228);
and U5476 (N_5476,N_5344,N_5263);
or U5477 (N_5477,N_5250,N_5252);
nand U5478 (N_5478,N_5260,N_5391);
or U5479 (N_5479,N_5319,N_5202);
nor U5480 (N_5480,N_5305,N_5314);
nor U5481 (N_5481,N_5307,N_5242);
and U5482 (N_5482,N_5255,N_5241);
nor U5483 (N_5483,N_5399,N_5218);
and U5484 (N_5484,N_5363,N_5394);
or U5485 (N_5485,N_5315,N_5337);
and U5486 (N_5486,N_5201,N_5331);
or U5487 (N_5487,N_5343,N_5258);
or U5488 (N_5488,N_5216,N_5376);
and U5489 (N_5489,N_5293,N_5317);
nor U5490 (N_5490,N_5247,N_5232);
and U5491 (N_5491,N_5335,N_5206);
xor U5492 (N_5492,N_5311,N_5267);
or U5493 (N_5493,N_5235,N_5349);
nor U5494 (N_5494,N_5375,N_5284);
and U5495 (N_5495,N_5372,N_5294);
or U5496 (N_5496,N_5290,N_5382);
and U5497 (N_5497,N_5388,N_5204);
xor U5498 (N_5498,N_5359,N_5380);
nor U5499 (N_5499,N_5249,N_5322);
nor U5500 (N_5500,N_5229,N_5319);
or U5501 (N_5501,N_5358,N_5347);
and U5502 (N_5502,N_5320,N_5382);
nand U5503 (N_5503,N_5339,N_5237);
nor U5504 (N_5504,N_5293,N_5394);
nor U5505 (N_5505,N_5348,N_5272);
nor U5506 (N_5506,N_5315,N_5210);
nor U5507 (N_5507,N_5367,N_5366);
xnor U5508 (N_5508,N_5378,N_5351);
or U5509 (N_5509,N_5342,N_5330);
nand U5510 (N_5510,N_5364,N_5343);
xnor U5511 (N_5511,N_5336,N_5207);
xor U5512 (N_5512,N_5275,N_5345);
xor U5513 (N_5513,N_5209,N_5289);
or U5514 (N_5514,N_5361,N_5202);
xnor U5515 (N_5515,N_5322,N_5373);
or U5516 (N_5516,N_5211,N_5314);
and U5517 (N_5517,N_5351,N_5261);
xnor U5518 (N_5518,N_5335,N_5300);
nor U5519 (N_5519,N_5210,N_5280);
and U5520 (N_5520,N_5227,N_5223);
nor U5521 (N_5521,N_5255,N_5336);
nor U5522 (N_5522,N_5342,N_5373);
xor U5523 (N_5523,N_5295,N_5365);
xnor U5524 (N_5524,N_5265,N_5347);
xor U5525 (N_5525,N_5308,N_5284);
or U5526 (N_5526,N_5312,N_5357);
or U5527 (N_5527,N_5350,N_5231);
and U5528 (N_5528,N_5361,N_5394);
xnor U5529 (N_5529,N_5301,N_5295);
xnor U5530 (N_5530,N_5327,N_5396);
nor U5531 (N_5531,N_5262,N_5228);
and U5532 (N_5532,N_5350,N_5337);
and U5533 (N_5533,N_5200,N_5249);
xnor U5534 (N_5534,N_5332,N_5301);
and U5535 (N_5535,N_5297,N_5233);
and U5536 (N_5536,N_5361,N_5246);
xnor U5537 (N_5537,N_5225,N_5270);
nand U5538 (N_5538,N_5253,N_5299);
xor U5539 (N_5539,N_5368,N_5394);
and U5540 (N_5540,N_5225,N_5327);
nor U5541 (N_5541,N_5357,N_5246);
or U5542 (N_5542,N_5242,N_5253);
nor U5543 (N_5543,N_5387,N_5300);
nor U5544 (N_5544,N_5335,N_5220);
xor U5545 (N_5545,N_5325,N_5230);
nor U5546 (N_5546,N_5228,N_5315);
xnor U5547 (N_5547,N_5361,N_5278);
and U5548 (N_5548,N_5224,N_5383);
or U5549 (N_5549,N_5361,N_5357);
and U5550 (N_5550,N_5218,N_5271);
nor U5551 (N_5551,N_5340,N_5227);
xor U5552 (N_5552,N_5270,N_5276);
or U5553 (N_5553,N_5293,N_5224);
nor U5554 (N_5554,N_5216,N_5385);
xor U5555 (N_5555,N_5369,N_5284);
or U5556 (N_5556,N_5283,N_5328);
xnor U5557 (N_5557,N_5395,N_5302);
nor U5558 (N_5558,N_5314,N_5363);
nor U5559 (N_5559,N_5234,N_5278);
xnor U5560 (N_5560,N_5372,N_5371);
and U5561 (N_5561,N_5265,N_5314);
and U5562 (N_5562,N_5230,N_5250);
nand U5563 (N_5563,N_5361,N_5304);
xnor U5564 (N_5564,N_5397,N_5262);
xnor U5565 (N_5565,N_5299,N_5329);
or U5566 (N_5566,N_5266,N_5265);
or U5567 (N_5567,N_5234,N_5296);
nor U5568 (N_5568,N_5371,N_5277);
nor U5569 (N_5569,N_5223,N_5217);
nor U5570 (N_5570,N_5263,N_5275);
nand U5571 (N_5571,N_5346,N_5221);
nand U5572 (N_5572,N_5386,N_5322);
and U5573 (N_5573,N_5236,N_5353);
nand U5574 (N_5574,N_5302,N_5290);
nand U5575 (N_5575,N_5365,N_5302);
nand U5576 (N_5576,N_5247,N_5293);
nor U5577 (N_5577,N_5344,N_5387);
xor U5578 (N_5578,N_5290,N_5235);
xnor U5579 (N_5579,N_5205,N_5226);
and U5580 (N_5580,N_5275,N_5386);
nor U5581 (N_5581,N_5306,N_5234);
xor U5582 (N_5582,N_5355,N_5254);
and U5583 (N_5583,N_5354,N_5347);
and U5584 (N_5584,N_5301,N_5286);
or U5585 (N_5585,N_5374,N_5297);
xor U5586 (N_5586,N_5247,N_5222);
or U5587 (N_5587,N_5334,N_5312);
nand U5588 (N_5588,N_5222,N_5266);
xnor U5589 (N_5589,N_5248,N_5262);
xnor U5590 (N_5590,N_5377,N_5246);
nand U5591 (N_5591,N_5204,N_5226);
nand U5592 (N_5592,N_5398,N_5322);
or U5593 (N_5593,N_5253,N_5391);
or U5594 (N_5594,N_5261,N_5302);
or U5595 (N_5595,N_5354,N_5398);
nor U5596 (N_5596,N_5301,N_5267);
nand U5597 (N_5597,N_5259,N_5384);
or U5598 (N_5598,N_5330,N_5346);
nand U5599 (N_5599,N_5376,N_5353);
nor U5600 (N_5600,N_5465,N_5570);
and U5601 (N_5601,N_5501,N_5464);
and U5602 (N_5602,N_5406,N_5585);
nand U5603 (N_5603,N_5451,N_5595);
and U5604 (N_5604,N_5514,N_5461);
xor U5605 (N_5605,N_5591,N_5490);
or U5606 (N_5606,N_5547,N_5411);
nor U5607 (N_5607,N_5432,N_5594);
nand U5608 (N_5608,N_5436,N_5450);
or U5609 (N_5609,N_5418,N_5565);
nor U5610 (N_5610,N_5520,N_5409);
nand U5611 (N_5611,N_5425,N_5471);
and U5612 (N_5612,N_5574,N_5573);
and U5613 (N_5613,N_5568,N_5588);
nor U5614 (N_5614,N_5477,N_5423);
or U5615 (N_5615,N_5576,N_5557);
and U5616 (N_5616,N_5597,N_5463);
nor U5617 (N_5617,N_5455,N_5422);
and U5618 (N_5618,N_5518,N_5527);
nor U5619 (N_5619,N_5428,N_5505);
or U5620 (N_5620,N_5442,N_5545);
xor U5621 (N_5621,N_5507,N_5458);
and U5622 (N_5622,N_5402,N_5410);
and U5623 (N_5623,N_5445,N_5486);
xnor U5624 (N_5624,N_5586,N_5504);
or U5625 (N_5625,N_5438,N_5531);
or U5626 (N_5626,N_5589,N_5524);
xnor U5627 (N_5627,N_5408,N_5511);
nand U5628 (N_5628,N_5434,N_5500);
and U5629 (N_5629,N_5554,N_5599);
nand U5630 (N_5630,N_5489,N_5476);
xor U5631 (N_5631,N_5405,N_5470);
or U5632 (N_5632,N_5467,N_5496);
xor U5633 (N_5633,N_5466,N_5530);
or U5634 (N_5634,N_5572,N_5487);
nand U5635 (N_5635,N_5479,N_5493);
nor U5636 (N_5636,N_5532,N_5549);
nand U5637 (N_5637,N_5447,N_5564);
or U5638 (N_5638,N_5429,N_5566);
or U5639 (N_5639,N_5499,N_5481);
nand U5640 (N_5640,N_5494,N_5508);
or U5641 (N_5641,N_5483,N_5578);
xnor U5642 (N_5642,N_5400,N_5412);
and U5643 (N_5643,N_5468,N_5517);
nor U5644 (N_5644,N_5421,N_5540);
xnor U5645 (N_5645,N_5430,N_5569);
or U5646 (N_5646,N_5401,N_5521);
nand U5647 (N_5647,N_5431,N_5435);
nand U5648 (N_5648,N_5415,N_5516);
and U5649 (N_5649,N_5509,N_5528);
xnor U5650 (N_5650,N_5541,N_5482);
nor U5651 (N_5651,N_5539,N_5506);
xor U5652 (N_5652,N_5502,N_5550);
xnor U5653 (N_5653,N_5439,N_5558);
nand U5654 (N_5654,N_5498,N_5403);
nor U5655 (N_5655,N_5491,N_5598);
and U5656 (N_5656,N_5556,N_5592);
xnor U5657 (N_5657,N_5561,N_5581);
and U5658 (N_5658,N_5596,N_5536);
xnor U5659 (N_5659,N_5407,N_5563);
nor U5660 (N_5660,N_5462,N_5551);
nor U5661 (N_5661,N_5460,N_5575);
nand U5662 (N_5662,N_5484,N_5526);
or U5663 (N_5663,N_5478,N_5522);
xnor U5664 (N_5664,N_5559,N_5452);
and U5665 (N_5665,N_5542,N_5454);
and U5666 (N_5666,N_5453,N_5579);
nand U5667 (N_5667,N_5417,N_5587);
or U5668 (N_5668,N_5593,N_5525);
xor U5669 (N_5669,N_5529,N_5571);
and U5670 (N_5670,N_5426,N_5538);
or U5671 (N_5671,N_5583,N_5475);
nor U5672 (N_5672,N_5562,N_5441);
or U5673 (N_5673,N_5495,N_5444);
or U5674 (N_5674,N_5537,N_5420);
xor U5675 (N_5675,N_5419,N_5437);
nand U5676 (N_5676,N_5560,N_5533);
xnor U5677 (N_5677,N_5546,N_5473);
or U5678 (N_5678,N_5427,N_5446);
xnor U5679 (N_5679,N_5535,N_5469);
xnor U5680 (N_5680,N_5433,N_5552);
xnor U5681 (N_5681,N_5456,N_5416);
xor U5682 (N_5682,N_5414,N_5480);
nand U5683 (N_5683,N_5584,N_5510);
nor U5684 (N_5684,N_5497,N_5503);
xnor U5685 (N_5685,N_5488,N_5448);
nor U5686 (N_5686,N_5443,N_5534);
or U5687 (N_5687,N_5440,N_5543);
xor U5688 (N_5688,N_5459,N_5449);
xnor U5689 (N_5689,N_5512,N_5580);
and U5690 (N_5690,N_5523,N_5577);
nor U5691 (N_5691,N_5472,N_5555);
and U5692 (N_5692,N_5553,N_5548);
nor U5693 (N_5693,N_5457,N_5544);
nor U5694 (N_5694,N_5413,N_5590);
nor U5695 (N_5695,N_5513,N_5404);
xor U5696 (N_5696,N_5515,N_5519);
or U5697 (N_5697,N_5485,N_5492);
and U5698 (N_5698,N_5582,N_5424);
xor U5699 (N_5699,N_5567,N_5474);
or U5700 (N_5700,N_5419,N_5481);
xor U5701 (N_5701,N_5540,N_5576);
or U5702 (N_5702,N_5468,N_5507);
nor U5703 (N_5703,N_5445,N_5416);
nor U5704 (N_5704,N_5484,N_5550);
xnor U5705 (N_5705,N_5472,N_5431);
or U5706 (N_5706,N_5552,N_5508);
or U5707 (N_5707,N_5504,N_5591);
and U5708 (N_5708,N_5532,N_5513);
nor U5709 (N_5709,N_5490,N_5470);
and U5710 (N_5710,N_5506,N_5419);
nor U5711 (N_5711,N_5454,N_5405);
nand U5712 (N_5712,N_5583,N_5411);
xnor U5713 (N_5713,N_5455,N_5460);
nor U5714 (N_5714,N_5570,N_5407);
nor U5715 (N_5715,N_5477,N_5597);
nor U5716 (N_5716,N_5502,N_5419);
and U5717 (N_5717,N_5486,N_5433);
xor U5718 (N_5718,N_5424,N_5554);
xnor U5719 (N_5719,N_5534,N_5553);
nor U5720 (N_5720,N_5572,N_5599);
or U5721 (N_5721,N_5589,N_5575);
and U5722 (N_5722,N_5438,N_5488);
xor U5723 (N_5723,N_5439,N_5539);
nand U5724 (N_5724,N_5544,N_5552);
nand U5725 (N_5725,N_5452,N_5533);
nor U5726 (N_5726,N_5597,N_5411);
xnor U5727 (N_5727,N_5497,N_5448);
and U5728 (N_5728,N_5445,N_5429);
xnor U5729 (N_5729,N_5477,N_5518);
nor U5730 (N_5730,N_5560,N_5497);
nor U5731 (N_5731,N_5425,N_5595);
nand U5732 (N_5732,N_5511,N_5433);
and U5733 (N_5733,N_5559,N_5440);
and U5734 (N_5734,N_5493,N_5414);
and U5735 (N_5735,N_5409,N_5580);
nor U5736 (N_5736,N_5439,N_5540);
nand U5737 (N_5737,N_5582,N_5566);
or U5738 (N_5738,N_5428,N_5481);
nor U5739 (N_5739,N_5519,N_5580);
or U5740 (N_5740,N_5460,N_5431);
and U5741 (N_5741,N_5491,N_5489);
and U5742 (N_5742,N_5421,N_5425);
nand U5743 (N_5743,N_5525,N_5599);
or U5744 (N_5744,N_5434,N_5453);
and U5745 (N_5745,N_5481,N_5449);
nor U5746 (N_5746,N_5437,N_5405);
xor U5747 (N_5747,N_5441,N_5444);
or U5748 (N_5748,N_5561,N_5482);
nand U5749 (N_5749,N_5457,N_5594);
and U5750 (N_5750,N_5478,N_5553);
nor U5751 (N_5751,N_5583,N_5419);
or U5752 (N_5752,N_5592,N_5576);
and U5753 (N_5753,N_5487,N_5512);
nand U5754 (N_5754,N_5431,N_5458);
and U5755 (N_5755,N_5597,N_5407);
and U5756 (N_5756,N_5522,N_5567);
and U5757 (N_5757,N_5593,N_5464);
and U5758 (N_5758,N_5459,N_5485);
or U5759 (N_5759,N_5555,N_5479);
nand U5760 (N_5760,N_5456,N_5468);
xor U5761 (N_5761,N_5428,N_5578);
xnor U5762 (N_5762,N_5415,N_5547);
or U5763 (N_5763,N_5420,N_5548);
nand U5764 (N_5764,N_5455,N_5503);
and U5765 (N_5765,N_5461,N_5486);
nor U5766 (N_5766,N_5429,N_5541);
or U5767 (N_5767,N_5523,N_5405);
nor U5768 (N_5768,N_5504,N_5492);
nand U5769 (N_5769,N_5599,N_5485);
or U5770 (N_5770,N_5505,N_5478);
and U5771 (N_5771,N_5576,N_5453);
nand U5772 (N_5772,N_5492,N_5542);
xnor U5773 (N_5773,N_5565,N_5442);
and U5774 (N_5774,N_5594,N_5550);
xnor U5775 (N_5775,N_5435,N_5422);
or U5776 (N_5776,N_5563,N_5491);
and U5777 (N_5777,N_5412,N_5524);
or U5778 (N_5778,N_5476,N_5588);
xor U5779 (N_5779,N_5473,N_5460);
and U5780 (N_5780,N_5472,N_5575);
and U5781 (N_5781,N_5580,N_5578);
nor U5782 (N_5782,N_5466,N_5476);
or U5783 (N_5783,N_5550,N_5406);
and U5784 (N_5784,N_5442,N_5483);
nor U5785 (N_5785,N_5440,N_5507);
xor U5786 (N_5786,N_5572,N_5440);
nand U5787 (N_5787,N_5496,N_5454);
nand U5788 (N_5788,N_5529,N_5405);
xor U5789 (N_5789,N_5414,N_5423);
nand U5790 (N_5790,N_5561,N_5511);
xnor U5791 (N_5791,N_5529,N_5502);
nand U5792 (N_5792,N_5436,N_5513);
nand U5793 (N_5793,N_5561,N_5452);
and U5794 (N_5794,N_5464,N_5566);
or U5795 (N_5795,N_5406,N_5567);
nand U5796 (N_5796,N_5478,N_5508);
and U5797 (N_5797,N_5403,N_5503);
nand U5798 (N_5798,N_5522,N_5420);
and U5799 (N_5799,N_5500,N_5519);
nor U5800 (N_5800,N_5671,N_5736);
and U5801 (N_5801,N_5642,N_5639);
nor U5802 (N_5802,N_5614,N_5740);
and U5803 (N_5803,N_5654,N_5660);
and U5804 (N_5804,N_5719,N_5612);
nor U5805 (N_5805,N_5763,N_5703);
or U5806 (N_5806,N_5688,N_5712);
xnor U5807 (N_5807,N_5794,N_5786);
nor U5808 (N_5808,N_5638,N_5622);
nand U5809 (N_5809,N_5726,N_5760);
or U5810 (N_5810,N_5635,N_5680);
xor U5811 (N_5811,N_5697,N_5686);
nor U5812 (N_5812,N_5776,N_5746);
or U5813 (N_5813,N_5675,N_5669);
xnor U5814 (N_5814,N_5792,N_5771);
nand U5815 (N_5815,N_5750,N_5618);
nand U5816 (N_5816,N_5742,N_5714);
or U5817 (N_5817,N_5748,N_5749);
xnor U5818 (N_5818,N_5640,N_5615);
nor U5819 (N_5819,N_5787,N_5788);
and U5820 (N_5820,N_5708,N_5772);
and U5821 (N_5821,N_5646,N_5626);
and U5822 (N_5822,N_5758,N_5636);
and U5823 (N_5823,N_5713,N_5670);
nand U5824 (N_5824,N_5665,N_5644);
nor U5825 (N_5825,N_5661,N_5616);
nand U5826 (N_5826,N_5667,N_5691);
xor U5827 (N_5827,N_5751,N_5798);
nand U5828 (N_5828,N_5630,N_5651);
xnor U5829 (N_5829,N_5756,N_5725);
and U5830 (N_5830,N_5657,N_5608);
nor U5831 (N_5831,N_5732,N_5699);
and U5832 (N_5832,N_5782,N_5747);
nor U5833 (N_5833,N_5655,N_5765);
xnor U5834 (N_5834,N_5621,N_5648);
nor U5835 (N_5835,N_5724,N_5768);
or U5836 (N_5836,N_5679,N_5643);
xnor U5837 (N_5837,N_5650,N_5779);
nor U5838 (N_5838,N_5666,N_5743);
and U5839 (N_5839,N_5609,N_5777);
or U5840 (N_5840,N_5753,N_5637);
and U5841 (N_5841,N_5767,N_5668);
or U5842 (N_5842,N_5656,N_5766);
nand U5843 (N_5843,N_5705,N_5775);
nand U5844 (N_5844,N_5603,N_5602);
nor U5845 (N_5845,N_5789,N_5662);
or U5846 (N_5846,N_5625,N_5600);
nor U5847 (N_5847,N_5659,N_5623);
nand U5848 (N_5848,N_5734,N_5702);
or U5849 (N_5849,N_5704,N_5664);
and U5850 (N_5850,N_5658,N_5723);
nor U5851 (N_5851,N_5678,N_5715);
nor U5852 (N_5852,N_5793,N_5663);
nor U5853 (N_5853,N_5716,N_5711);
nand U5854 (N_5854,N_5687,N_5709);
or U5855 (N_5855,N_5795,N_5721);
nand U5856 (N_5856,N_5677,N_5604);
and U5857 (N_5857,N_5647,N_5718);
and U5858 (N_5858,N_5729,N_5745);
xnor U5859 (N_5859,N_5733,N_5674);
xnor U5860 (N_5860,N_5601,N_5755);
and U5861 (N_5861,N_5681,N_5693);
nor U5862 (N_5862,N_5683,N_5762);
or U5863 (N_5863,N_5744,N_5629);
or U5864 (N_5864,N_5781,N_5757);
or U5865 (N_5865,N_5796,N_5627);
and U5866 (N_5866,N_5738,N_5791);
and U5867 (N_5867,N_5631,N_5619);
nor U5868 (N_5868,N_5720,N_5672);
or U5869 (N_5869,N_5695,N_5613);
nand U5870 (N_5870,N_5628,N_5790);
or U5871 (N_5871,N_5717,N_5676);
or U5872 (N_5872,N_5769,N_5690);
nor U5873 (N_5873,N_5710,N_5694);
and U5874 (N_5874,N_5764,N_5739);
or U5875 (N_5875,N_5701,N_5700);
nand U5876 (N_5876,N_5652,N_5780);
or U5877 (N_5877,N_5761,N_5606);
nor U5878 (N_5878,N_5607,N_5797);
nand U5879 (N_5879,N_5706,N_5633);
xnor U5880 (N_5880,N_5774,N_5785);
xnor U5881 (N_5881,N_5684,N_5645);
and U5882 (N_5882,N_5673,N_5741);
or U5883 (N_5883,N_5641,N_5752);
nor U5884 (N_5884,N_5611,N_5692);
and U5885 (N_5885,N_5682,N_5634);
or U5886 (N_5886,N_5783,N_5685);
and U5887 (N_5887,N_5624,N_5784);
nand U5888 (N_5888,N_5722,N_5735);
or U5889 (N_5889,N_5778,N_5728);
and U5890 (N_5890,N_5617,N_5698);
nand U5891 (N_5891,N_5773,N_5770);
or U5892 (N_5892,N_5759,N_5610);
nor U5893 (N_5893,N_5754,N_5731);
xor U5894 (N_5894,N_5653,N_5605);
and U5895 (N_5895,N_5737,N_5707);
or U5896 (N_5896,N_5689,N_5799);
and U5897 (N_5897,N_5632,N_5696);
or U5898 (N_5898,N_5727,N_5649);
nor U5899 (N_5899,N_5620,N_5730);
nor U5900 (N_5900,N_5762,N_5724);
or U5901 (N_5901,N_5737,N_5799);
and U5902 (N_5902,N_5732,N_5703);
nand U5903 (N_5903,N_5692,N_5764);
xnor U5904 (N_5904,N_5680,N_5643);
xnor U5905 (N_5905,N_5647,N_5672);
nor U5906 (N_5906,N_5787,N_5647);
and U5907 (N_5907,N_5610,N_5794);
or U5908 (N_5908,N_5679,N_5793);
or U5909 (N_5909,N_5712,N_5686);
or U5910 (N_5910,N_5661,N_5774);
and U5911 (N_5911,N_5798,N_5647);
and U5912 (N_5912,N_5610,N_5699);
nand U5913 (N_5913,N_5737,N_5792);
and U5914 (N_5914,N_5674,N_5665);
or U5915 (N_5915,N_5696,N_5644);
and U5916 (N_5916,N_5753,N_5724);
nand U5917 (N_5917,N_5746,N_5690);
or U5918 (N_5918,N_5605,N_5652);
xnor U5919 (N_5919,N_5611,N_5630);
nor U5920 (N_5920,N_5683,N_5627);
and U5921 (N_5921,N_5779,N_5697);
nor U5922 (N_5922,N_5682,N_5728);
and U5923 (N_5923,N_5729,N_5753);
nand U5924 (N_5924,N_5633,N_5781);
xnor U5925 (N_5925,N_5748,N_5797);
nand U5926 (N_5926,N_5657,N_5722);
or U5927 (N_5927,N_5718,N_5738);
nand U5928 (N_5928,N_5767,N_5714);
xnor U5929 (N_5929,N_5741,N_5779);
and U5930 (N_5930,N_5648,N_5729);
xnor U5931 (N_5931,N_5725,N_5601);
or U5932 (N_5932,N_5694,N_5767);
or U5933 (N_5933,N_5782,N_5633);
xor U5934 (N_5934,N_5750,N_5772);
xor U5935 (N_5935,N_5634,N_5666);
xor U5936 (N_5936,N_5620,N_5790);
or U5937 (N_5937,N_5711,N_5670);
and U5938 (N_5938,N_5723,N_5669);
or U5939 (N_5939,N_5798,N_5715);
and U5940 (N_5940,N_5617,N_5667);
nor U5941 (N_5941,N_5747,N_5665);
nand U5942 (N_5942,N_5783,N_5749);
nor U5943 (N_5943,N_5759,N_5635);
and U5944 (N_5944,N_5717,N_5765);
and U5945 (N_5945,N_5664,N_5779);
or U5946 (N_5946,N_5600,N_5784);
and U5947 (N_5947,N_5656,N_5726);
nand U5948 (N_5948,N_5696,N_5737);
or U5949 (N_5949,N_5602,N_5659);
nor U5950 (N_5950,N_5618,N_5617);
and U5951 (N_5951,N_5624,N_5609);
and U5952 (N_5952,N_5737,N_5642);
xor U5953 (N_5953,N_5673,N_5776);
or U5954 (N_5954,N_5724,N_5774);
nor U5955 (N_5955,N_5782,N_5780);
nor U5956 (N_5956,N_5764,N_5763);
nor U5957 (N_5957,N_5614,N_5668);
and U5958 (N_5958,N_5787,N_5702);
nor U5959 (N_5959,N_5745,N_5775);
xnor U5960 (N_5960,N_5655,N_5604);
or U5961 (N_5961,N_5623,N_5712);
nand U5962 (N_5962,N_5797,N_5781);
xnor U5963 (N_5963,N_5769,N_5660);
and U5964 (N_5964,N_5683,N_5759);
or U5965 (N_5965,N_5678,N_5786);
nand U5966 (N_5966,N_5788,N_5615);
xnor U5967 (N_5967,N_5776,N_5709);
and U5968 (N_5968,N_5645,N_5679);
xor U5969 (N_5969,N_5709,N_5615);
nor U5970 (N_5970,N_5776,N_5603);
or U5971 (N_5971,N_5744,N_5689);
nor U5972 (N_5972,N_5758,N_5713);
and U5973 (N_5973,N_5728,N_5788);
and U5974 (N_5974,N_5661,N_5600);
and U5975 (N_5975,N_5670,N_5766);
and U5976 (N_5976,N_5756,N_5692);
xnor U5977 (N_5977,N_5759,N_5675);
and U5978 (N_5978,N_5767,N_5775);
and U5979 (N_5979,N_5715,N_5680);
nor U5980 (N_5980,N_5747,N_5741);
nor U5981 (N_5981,N_5676,N_5674);
xor U5982 (N_5982,N_5745,N_5632);
or U5983 (N_5983,N_5726,N_5663);
nor U5984 (N_5984,N_5666,N_5720);
nor U5985 (N_5985,N_5749,N_5670);
or U5986 (N_5986,N_5704,N_5720);
or U5987 (N_5987,N_5748,N_5631);
xnor U5988 (N_5988,N_5760,N_5660);
nand U5989 (N_5989,N_5767,N_5713);
or U5990 (N_5990,N_5691,N_5710);
nor U5991 (N_5991,N_5753,N_5623);
nor U5992 (N_5992,N_5690,N_5667);
nor U5993 (N_5993,N_5619,N_5616);
and U5994 (N_5994,N_5724,N_5685);
xnor U5995 (N_5995,N_5620,N_5795);
xor U5996 (N_5996,N_5767,N_5739);
nand U5997 (N_5997,N_5685,N_5777);
nand U5998 (N_5998,N_5721,N_5690);
nand U5999 (N_5999,N_5634,N_5600);
nand U6000 (N_6000,N_5817,N_5837);
nor U6001 (N_6001,N_5944,N_5862);
nand U6002 (N_6002,N_5877,N_5997);
nand U6003 (N_6003,N_5946,N_5863);
nand U6004 (N_6004,N_5925,N_5991);
nor U6005 (N_6005,N_5869,N_5822);
xnor U6006 (N_6006,N_5897,N_5834);
nand U6007 (N_6007,N_5823,N_5998);
xor U6008 (N_6008,N_5811,N_5835);
or U6009 (N_6009,N_5990,N_5814);
nand U6010 (N_6010,N_5865,N_5892);
and U6011 (N_6011,N_5910,N_5994);
nor U6012 (N_6012,N_5971,N_5839);
nand U6013 (N_6013,N_5833,N_5856);
or U6014 (N_6014,N_5953,N_5969);
xnor U6015 (N_6015,N_5857,N_5900);
and U6016 (N_6016,N_5840,N_5975);
nand U6017 (N_6017,N_5887,N_5976);
or U6018 (N_6018,N_5884,N_5945);
or U6019 (N_6019,N_5813,N_5851);
and U6020 (N_6020,N_5893,N_5977);
xnor U6021 (N_6021,N_5861,N_5988);
nand U6022 (N_6022,N_5939,N_5923);
nand U6023 (N_6023,N_5830,N_5885);
nor U6024 (N_6024,N_5993,N_5938);
or U6025 (N_6025,N_5846,N_5956);
and U6026 (N_6026,N_5906,N_5920);
and U6027 (N_6027,N_5806,N_5951);
and U6028 (N_6028,N_5888,N_5917);
xnor U6029 (N_6029,N_5864,N_5911);
nor U6030 (N_6030,N_5809,N_5886);
nand U6031 (N_6031,N_5881,N_5967);
nand U6032 (N_6032,N_5899,N_5876);
nand U6033 (N_6033,N_5818,N_5890);
or U6034 (N_6034,N_5859,N_5875);
nand U6035 (N_6035,N_5867,N_5970);
or U6036 (N_6036,N_5921,N_5836);
xnor U6037 (N_6037,N_5803,N_5821);
nor U6038 (N_6038,N_5807,N_5812);
and U6039 (N_6039,N_5802,N_5962);
nor U6040 (N_6040,N_5826,N_5941);
nor U6041 (N_6041,N_5901,N_5903);
or U6042 (N_6042,N_5905,N_5908);
nor U6043 (N_6043,N_5928,N_5879);
and U6044 (N_6044,N_5842,N_5847);
xnor U6045 (N_6045,N_5954,N_5889);
or U6046 (N_6046,N_5963,N_5855);
nand U6047 (N_6047,N_5979,N_5950);
or U6048 (N_6048,N_5932,N_5915);
xor U6049 (N_6049,N_5853,N_5808);
xor U6050 (N_6050,N_5849,N_5828);
nand U6051 (N_6051,N_5987,N_5918);
or U6052 (N_6052,N_5843,N_5919);
nor U6053 (N_6053,N_5986,N_5931);
nand U6054 (N_6054,N_5972,N_5958);
or U6055 (N_6055,N_5978,N_5848);
nor U6056 (N_6056,N_5858,N_5914);
or U6057 (N_6057,N_5937,N_5955);
nor U6058 (N_6058,N_5926,N_5819);
nand U6059 (N_6059,N_5841,N_5996);
xor U6060 (N_6060,N_5952,N_5912);
nand U6061 (N_6061,N_5825,N_5973);
and U6062 (N_6062,N_5820,N_5999);
or U6063 (N_6063,N_5844,N_5829);
and U6064 (N_6064,N_5966,N_5929);
or U6065 (N_6065,N_5816,N_5949);
xnor U6066 (N_6066,N_5805,N_5930);
or U6067 (N_6067,N_5832,N_5831);
xor U6068 (N_6068,N_5810,N_5981);
nand U6069 (N_6069,N_5922,N_5804);
and U6070 (N_6070,N_5873,N_5870);
nor U6071 (N_6071,N_5924,N_5852);
nor U6072 (N_6072,N_5800,N_5933);
xnor U6073 (N_6073,N_5936,N_5868);
nand U6074 (N_6074,N_5882,N_5801);
and U6075 (N_6075,N_5824,N_5947);
and U6076 (N_6076,N_5974,N_5913);
xor U6077 (N_6077,N_5907,N_5943);
nand U6078 (N_6078,N_5959,N_5904);
nor U6079 (N_6079,N_5935,N_5902);
xor U6080 (N_6080,N_5992,N_5850);
nand U6081 (N_6081,N_5815,N_5965);
or U6082 (N_6082,N_5895,N_5871);
and U6083 (N_6083,N_5934,N_5898);
and U6084 (N_6084,N_5909,N_5891);
nor U6085 (N_6085,N_5872,N_5916);
and U6086 (N_6086,N_5957,N_5982);
nor U6087 (N_6087,N_5860,N_5854);
or U6088 (N_6088,N_5942,N_5961);
nor U6089 (N_6089,N_5985,N_5980);
nor U6090 (N_6090,N_5984,N_5995);
and U6091 (N_6091,N_5968,N_5927);
nor U6092 (N_6092,N_5878,N_5838);
xor U6093 (N_6093,N_5827,N_5874);
nor U6094 (N_6094,N_5894,N_5960);
nand U6095 (N_6095,N_5964,N_5983);
nor U6096 (N_6096,N_5880,N_5845);
nand U6097 (N_6097,N_5989,N_5948);
nand U6098 (N_6098,N_5866,N_5940);
and U6099 (N_6099,N_5896,N_5883);
nand U6100 (N_6100,N_5889,N_5812);
or U6101 (N_6101,N_5910,N_5894);
xor U6102 (N_6102,N_5885,N_5946);
or U6103 (N_6103,N_5808,N_5928);
nand U6104 (N_6104,N_5967,N_5908);
and U6105 (N_6105,N_5964,N_5875);
and U6106 (N_6106,N_5962,N_5876);
nand U6107 (N_6107,N_5939,N_5806);
xnor U6108 (N_6108,N_5981,N_5953);
or U6109 (N_6109,N_5992,N_5986);
nor U6110 (N_6110,N_5895,N_5909);
nand U6111 (N_6111,N_5883,N_5890);
and U6112 (N_6112,N_5805,N_5851);
nor U6113 (N_6113,N_5938,N_5870);
or U6114 (N_6114,N_5986,N_5899);
or U6115 (N_6115,N_5870,N_5968);
or U6116 (N_6116,N_5833,N_5835);
xor U6117 (N_6117,N_5974,N_5959);
and U6118 (N_6118,N_5981,N_5808);
nand U6119 (N_6119,N_5872,N_5905);
nand U6120 (N_6120,N_5874,N_5993);
and U6121 (N_6121,N_5886,N_5993);
xnor U6122 (N_6122,N_5926,N_5896);
or U6123 (N_6123,N_5983,N_5895);
and U6124 (N_6124,N_5803,N_5834);
nand U6125 (N_6125,N_5888,N_5894);
nor U6126 (N_6126,N_5889,N_5823);
nor U6127 (N_6127,N_5841,N_5818);
xnor U6128 (N_6128,N_5867,N_5949);
and U6129 (N_6129,N_5980,N_5802);
and U6130 (N_6130,N_5837,N_5881);
or U6131 (N_6131,N_5823,N_5824);
or U6132 (N_6132,N_5911,N_5983);
or U6133 (N_6133,N_5821,N_5869);
or U6134 (N_6134,N_5908,N_5808);
nor U6135 (N_6135,N_5855,N_5837);
xnor U6136 (N_6136,N_5915,N_5806);
xnor U6137 (N_6137,N_5960,N_5904);
or U6138 (N_6138,N_5957,N_5973);
and U6139 (N_6139,N_5818,N_5907);
xor U6140 (N_6140,N_5828,N_5946);
xor U6141 (N_6141,N_5892,N_5897);
nor U6142 (N_6142,N_5877,N_5940);
and U6143 (N_6143,N_5829,N_5920);
and U6144 (N_6144,N_5988,N_5981);
nor U6145 (N_6145,N_5986,N_5967);
nand U6146 (N_6146,N_5971,N_5997);
or U6147 (N_6147,N_5863,N_5841);
and U6148 (N_6148,N_5988,N_5870);
nor U6149 (N_6149,N_5948,N_5886);
and U6150 (N_6150,N_5958,N_5971);
and U6151 (N_6151,N_5854,N_5905);
xor U6152 (N_6152,N_5928,N_5913);
and U6153 (N_6153,N_5987,N_5833);
nand U6154 (N_6154,N_5820,N_5900);
or U6155 (N_6155,N_5917,N_5916);
and U6156 (N_6156,N_5973,N_5853);
nand U6157 (N_6157,N_5924,N_5947);
nor U6158 (N_6158,N_5847,N_5809);
nor U6159 (N_6159,N_5868,N_5946);
xor U6160 (N_6160,N_5913,N_5812);
nand U6161 (N_6161,N_5883,N_5914);
nor U6162 (N_6162,N_5976,N_5978);
and U6163 (N_6163,N_5850,N_5890);
xor U6164 (N_6164,N_5955,N_5811);
nor U6165 (N_6165,N_5921,N_5972);
xor U6166 (N_6166,N_5820,N_5906);
xnor U6167 (N_6167,N_5932,N_5867);
nand U6168 (N_6168,N_5955,N_5849);
nand U6169 (N_6169,N_5934,N_5991);
nor U6170 (N_6170,N_5817,N_5984);
nand U6171 (N_6171,N_5942,N_5966);
xnor U6172 (N_6172,N_5987,N_5893);
or U6173 (N_6173,N_5862,N_5904);
and U6174 (N_6174,N_5876,N_5879);
nor U6175 (N_6175,N_5844,N_5996);
and U6176 (N_6176,N_5913,N_5811);
nor U6177 (N_6177,N_5967,N_5809);
nor U6178 (N_6178,N_5812,N_5820);
nand U6179 (N_6179,N_5953,N_5838);
and U6180 (N_6180,N_5860,N_5859);
nand U6181 (N_6181,N_5870,N_5939);
xnor U6182 (N_6182,N_5998,N_5973);
or U6183 (N_6183,N_5895,N_5917);
nand U6184 (N_6184,N_5918,N_5911);
or U6185 (N_6185,N_5822,N_5975);
xnor U6186 (N_6186,N_5931,N_5827);
and U6187 (N_6187,N_5816,N_5907);
and U6188 (N_6188,N_5890,N_5941);
nor U6189 (N_6189,N_5982,N_5910);
nand U6190 (N_6190,N_5848,N_5874);
xor U6191 (N_6191,N_5974,N_5810);
nor U6192 (N_6192,N_5890,N_5822);
xor U6193 (N_6193,N_5818,N_5941);
nor U6194 (N_6194,N_5911,N_5950);
nand U6195 (N_6195,N_5828,N_5916);
or U6196 (N_6196,N_5845,N_5905);
nor U6197 (N_6197,N_5981,N_5850);
and U6198 (N_6198,N_5879,N_5918);
nand U6199 (N_6199,N_5955,N_5933);
and U6200 (N_6200,N_6139,N_6101);
nor U6201 (N_6201,N_6035,N_6104);
and U6202 (N_6202,N_6148,N_6002);
or U6203 (N_6203,N_6106,N_6188);
nor U6204 (N_6204,N_6156,N_6066);
xnor U6205 (N_6205,N_6013,N_6081);
xor U6206 (N_6206,N_6029,N_6086);
nand U6207 (N_6207,N_6087,N_6033);
or U6208 (N_6208,N_6090,N_6126);
or U6209 (N_6209,N_6059,N_6018);
xnor U6210 (N_6210,N_6099,N_6129);
nand U6211 (N_6211,N_6187,N_6116);
or U6212 (N_6212,N_6056,N_6068);
and U6213 (N_6213,N_6162,N_6118);
xnor U6214 (N_6214,N_6113,N_6042);
nand U6215 (N_6215,N_6149,N_6171);
xor U6216 (N_6216,N_6192,N_6055);
or U6217 (N_6217,N_6112,N_6084);
or U6218 (N_6218,N_6095,N_6091);
and U6219 (N_6219,N_6021,N_6164);
and U6220 (N_6220,N_6000,N_6168);
xnor U6221 (N_6221,N_6170,N_6058);
or U6222 (N_6222,N_6130,N_6184);
nand U6223 (N_6223,N_6123,N_6011);
nor U6224 (N_6224,N_6193,N_6017);
nand U6225 (N_6225,N_6077,N_6098);
or U6226 (N_6226,N_6159,N_6031);
xor U6227 (N_6227,N_6146,N_6134);
and U6228 (N_6228,N_6092,N_6183);
nand U6229 (N_6229,N_6069,N_6097);
nor U6230 (N_6230,N_6132,N_6120);
nand U6231 (N_6231,N_6030,N_6065);
xor U6232 (N_6232,N_6199,N_6075);
nand U6233 (N_6233,N_6125,N_6073);
xor U6234 (N_6234,N_6180,N_6052);
or U6235 (N_6235,N_6185,N_6102);
and U6236 (N_6236,N_6107,N_6043);
nor U6237 (N_6237,N_6103,N_6181);
or U6238 (N_6238,N_6145,N_6191);
xnor U6239 (N_6239,N_6001,N_6061);
nor U6240 (N_6240,N_6062,N_6039);
and U6241 (N_6241,N_6195,N_6140);
or U6242 (N_6242,N_6023,N_6109);
or U6243 (N_6243,N_6009,N_6105);
nor U6244 (N_6244,N_6190,N_6147);
or U6245 (N_6245,N_6122,N_6079);
nand U6246 (N_6246,N_6198,N_6182);
or U6247 (N_6247,N_6005,N_6111);
nor U6248 (N_6248,N_6119,N_6114);
nor U6249 (N_6249,N_6027,N_6110);
nand U6250 (N_6250,N_6142,N_6025);
xor U6251 (N_6251,N_6089,N_6050);
and U6252 (N_6252,N_6172,N_6071);
nand U6253 (N_6253,N_6076,N_6007);
nor U6254 (N_6254,N_6006,N_6128);
or U6255 (N_6255,N_6177,N_6088);
or U6256 (N_6256,N_6173,N_6040);
xor U6257 (N_6257,N_6044,N_6083);
and U6258 (N_6258,N_6048,N_6014);
and U6259 (N_6259,N_6189,N_6060);
nor U6260 (N_6260,N_6136,N_6019);
and U6261 (N_6261,N_6127,N_6155);
and U6262 (N_6262,N_6037,N_6175);
nor U6263 (N_6263,N_6135,N_6020);
xnor U6264 (N_6264,N_6161,N_6022);
xnor U6265 (N_6265,N_6012,N_6196);
xnor U6266 (N_6266,N_6047,N_6057);
nor U6267 (N_6267,N_6024,N_6165);
xnor U6268 (N_6268,N_6169,N_6094);
nor U6269 (N_6269,N_6036,N_6072);
or U6270 (N_6270,N_6045,N_6074);
and U6271 (N_6271,N_6131,N_6034);
and U6272 (N_6272,N_6160,N_6016);
xnor U6273 (N_6273,N_6176,N_6115);
nand U6274 (N_6274,N_6153,N_6008);
xnor U6275 (N_6275,N_6166,N_6194);
xor U6276 (N_6276,N_6124,N_6054);
nand U6277 (N_6277,N_6137,N_6151);
xor U6278 (N_6278,N_6041,N_6004);
and U6279 (N_6279,N_6138,N_6010);
or U6280 (N_6280,N_6051,N_6152);
nand U6281 (N_6281,N_6157,N_6108);
or U6282 (N_6282,N_6064,N_6144);
nor U6283 (N_6283,N_6067,N_6178);
or U6284 (N_6284,N_6143,N_6049);
nor U6285 (N_6285,N_6085,N_6082);
xnor U6286 (N_6286,N_6121,N_6078);
nor U6287 (N_6287,N_6133,N_6015);
nand U6288 (N_6288,N_6026,N_6032);
nor U6289 (N_6289,N_6154,N_6038);
nor U6290 (N_6290,N_6046,N_6100);
and U6291 (N_6291,N_6163,N_6028);
nor U6292 (N_6292,N_6158,N_6197);
and U6293 (N_6293,N_6117,N_6167);
nor U6294 (N_6294,N_6096,N_6070);
nand U6295 (N_6295,N_6063,N_6093);
nand U6296 (N_6296,N_6003,N_6141);
xnor U6297 (N_6297,N_6080,N_6186);
nand U6298 (N_6298,N_6174,N_6150);
xor U6299 (N_6299,N_6053,N_6179);
nand U6300 (N_6300,N_6057,N_6197);
nand U6301 (N_6301,N_6085,N_6095);
or U6302 (N_6302,N_6035,N_6012);
xor U6303 (N_6303,N_6091,N_6006);
xnor U6304 (N_6304,N_6066,N_6178);
xor U6305 (N_6305,N_6045,N_6164);
and U6306 (N_6306,N_6105,N_6074);
nor U6307 (N_6307,N_6084,N_6198);
and U6308 (N_6308,N_6122,N_6185);
nand U6309 (N_6309,N_6123,N_6158);
nor U6310 (N_6310,N_6065,N_6076);
nand U6311 (N_6311,N_6006,N_6008);
or U6312 (N_6312,N_6041,N_6076);
xnor U6313 (N_6313,N_6143,N_6041);
xnor U6314 (N_6314,N_6061,N_6064);
nor U6315 (N_6315,N_6152,N_6042);
nand U6316 (N_6316,N_6112,N_6182);
nor U6317 (N_6317,N_6020,N_6163);
and U6318 (N_6318,N_6065,N_6109);
or U6319 (N_6319,N_6059,N_6110);
or U6320 (N_6320,N_6165,N_6152);
xnor U6321 (N_6321,N_6110,N_6053);
nand U6322 (N_6322,N_6027,N_6083);
nand U6323 (N_6323,N_6181,N_6182);
nor U6324 (N_6324,N_6048,N_6166);
nand U6325 (N_6325,N_6042,N_6053);
xnor U6326 (N_6326,N_6068,N_6172);
xor U6327 (N_6327,N_6159,N_6059);
and U6328 (N_6328,N_6153,N_6093);
xnor U6329 (N_6329,N_6103,N_6037);
nand U6330 (N_6330,N_6160,N_6010);
nor U6331 (N_6331,N_6056,N_6014);
nand U6332 (N_6332,N_6199,N_6168);
and U6333 (N_6333,N_6095,N_6142);
or U6334 (N_6334,N_6145,N_6123);
xnor U6335 (N_6335,N_6098,N_6178);
nand U6336 (N_6336,N_6093,N_6075);
xnor U6337 (N_6337,N_6064,N_6146);
nor U6338 (N_6338,N_6120,N_6149);
or U6339 (N_6339,N_6144,N_6100);
xnor U6340 (N_6340,N_6018,N_6014);
nand U6341 (N_6341,N_6199,N_6066);
or U6342 (N_6342,N_6152,N_6159);
and U6343 (N_6343,N_6149,N_6027);
and U6344 (N_6344,N_6151,N_6008);
xnor U6345 (N_6345,N_6161,N_6016);
and U6346 (N_6346,N_6131,N_6009);
and U6347 (N_6347,N_6130,N_6138);
nor U6348 (N_6348,N_6057,N_6117);
and U6349 (N_6349,N_6094,N_6173);
nor U6350 (N_6350,N_6023,N_6056);
or U6351 (N_6351,N_6028,N_6142);
nand U6352 (N_6352,N_6185,N_6116);
and U6353 (N_6353,N_6022,N_6112);
nand U6354 (N_6354,N_6134,N_6039);
nor U6355 (N_6355,N_6055,N_6085);
nor U6356 (N_6356,N_6031,N_6172);
xor U6357 (N_6357,N_6050,N_6162);
xnor U6358 (N_6358,N_6164,N_6012);
and U6359 (N_6359,N_6120,N_6091);
and U6360 (N_6360,N_6018,N_6171);
nand U6361 (N_6361,N_6022,N_6013);
or U6362 (N_6362,N_6134,N_6119);
and U6363 (N_6363,N_6149,N_6089);
or U6364 (N_6364,N_6012,N_6059);
nor U6365 (N_6365,N_6069,N_6096);
nand U6366 (N_6366,N_6159,N_6182);
nor U6367 (N_6367,N_6088,N_6190);
xnor U6368 (N_6368,N_6114,N_6144);
xnor U6369 (N_6369,N_6179,N_6001);
or U6370 (N_6370,N_6106,N_6078);
xor U6371 (N_6371,N_6055,N_6127);
xnor U6372 (N_6372,N_6002,N_6127);
xor U6373 (N_6373,N_6194,N_6173);
nor U6374 (N_6374,N_6185,N_6015);
nand U6375 (N_6375,N_6059,N_6086);
or U6376 (N_6376,N_6005,N_6195);
and U6377 (N_6377,N_6184,N_6106);
nand U6378 (N_6378,N_6146,N_6099);
xnor U6379 (N_6379,N_6135,N_6084);
nand U6380 (N_6380,N_6099,N_6049);
xnor U6381 (N_6381,N_6127,N_6029);
nand U6382 (N_6382,N_6062,N_6040);
xor U6383 (N_6383,N_6160,N_6098);
nor U6384 (N_6384,N_6013,N_6143);
nor U6385 (N_6385,N_6138,N_6035);
and U6386 (N_6386,N_6115,N_6096);
nor U6387 (N_6387,N_6035,N_6097);
or U6388 (N_6388,N_6152,N_6049);
or U6389 (N_6389,N_6176,N_6120);
nand U6390 (N_6390,N_6113,N_6024);
or U6391 (N_6391,N_6066,N_6105);
nand U6392 (N_6392,N_6144,N_6148);
nand U6393 (N_6393,N_6019,N_6114);
and U6394 (N_6394,N_6047,N_6157);
and U6395 (N_6395,N_6152,N_6154);
nor U6396 (N_6396,N_6124,N_6163);
and U6397 (N_6397,N_6088,N_6093);
xnor U6398 (N_6398,N_6062,N_6198);
xnor U6399 (N_6399,N_6120,N_6114);
nor U6400 (N_6400,N_6385,N_6298);
nor U6401 (N_6401,N_6367,N_6350);
xor U6402 (N_6402,N_6299,N_6259);
or U6403 (N_6403,N_6279,N_6226);
nor U6404 (N_6404,N_6366,N_6258);
nand U6405 (N_6405,N_6390,N_6257);
and U6406 (N_6406,N_6239,N_6396);
xor U6407 (N_6407,N_6382,N_6281);
nor U6408 (N_6408,N_6236,N_6254);
nand U6409 (N_6409,N_6305,N_6381);
nor U6410 (N_6410,N_6276,N_6204);
and U6411 (N_6411,N_6373,N_6261);
nand U6412 (N_6412,N_6380,N_6317);
nand U6413 (N_6413,N_6384,N_6231);
nor U6414 (N_6414,N_6219,N_6272);
nand U6415 (N_6415,N_6289,N_6245);
nand U6416 (N_6416,N_6343,N_6216);
nor U6417 (N_6417,N_6293,N_6395);
or U6418 (N_6418,N_6360,N_6229);
or U6419 (N_6419,N_6277,N_6206);
xnor U6420 (N_6420,N_6205,N_6364);
or U6421 (N_6421,N_6394,N_6342);
and U6422 (N_6422,N_6301,N_6324);
nor U6423 (N_6423,N_6307,N_6212);
xor U6424 (N_6424,N_6297,N_6320);
nor U6425 (N_6425,N_6203,N_6354);
xnor U6426 (N_6426,N_6339,N_6311);
nor U6427 (N_6427,N_6250,N_6291);
and U6428 (N_6428,N_6295,N_6252);
or U6429 (N_6429,N_6282,N_6287);
or U6430 (N_6430,N_6338,N_6334);
nand U6431 (N_6431,N_6238,N_6316);
or U6432 (N_6432,N_6363,N_6294);
and U6433 (N_6433,N_6312,N_6327);
and U6434 (N_6434,N_6228,N_6248);
xor U6435 (N_6435,N_6217,N_6362);
nand U6436 (N_6436,N_6268,N_6233);
nand U6437 (N_6437,N_6335,N_6329);
and U6438 (N_6438,N_6377,N_6345);
xor U6439 (N_6439,N_6242,N_6237);
xor U6440 (N_6440,N_6256,N_6370);
xor U6441 (N_6441,N_6280,N_6222);
and U6442 (N_6442,N_6368,N_6365);
xnor U6443 (N_6443,N_6274,N_6220);
and U6444 (N_6444,N_6292,N_6232);
or U6445 (N_6445,N_6314,N_6375);
and U6446 (N_6446,N_6319,N_6318);
nor U6447 (N_6447,N_6397,N_6322);
xnor U6448 (N_6448,N_6234,N_6313);
and U6449 (N_6449,N_6208,N_6266);
and U6450 (N_6450,N_6227,N_6218);
and U6451 (N_6451,N_6347,N_6315);
nor U6452 (N_6452,N_6388,N_6358);
and U6453 (N_6453,N_6340,N_6378);
nand U6454 (N_6454,N_6303,N_6399);
or U6455 (N_6455,N_6356,N_6223);
nand U6456 (N_6456,N_6249,N_6288);
and U6457 (N_6457,N_6207,N_6210);
and U6458 (N_6458,N_6202,N_6251);
nand U6459 (N_6459,N_6309,N_6283);
nand U6460 (N_6460,N_6213,N_6304);
nand U6461 (N_6461,N_6284,N_6392);
or U6462 (N_6462,N_6214,N_6391);
xnor U6463 (N_6463,N_6271,N_6326);
or U6464 (N_6464,N_6243,N_6225);
and U6465 (N_6465,N_6308,N_6336);
nand U6466 (N_6466,N_6383,N_6247);
or U6467 (N_6467,N_6264,N_6328);
nand U6468 (N_6468,N_6331,N_6371);
nor U6469 (N_6469,N_6349,N_6270);
xnor U6470 (N_6470,N_6260,N_6398);
nor U6471 (N_6471,N_6201,N_6269);
nor U6472 (N_6472,N_6300,N_6348);
nor U6473 (N_6473,N_6351,N_6337);
nand U6474 (N_6474,N_6273,N_6372);
nor U6475 (N_6475,N_6253,N_6389);
xor U6476 (N_6476,N_6346,N_6355);
nor U6477 (N_6477,N_6359,N_6369);
nand U6478 (N_6478,N_6296,N_6341);
and U6479 (N_6479,N_6200,N_6306);
and U6480 (N_6480,N_6262,N_6265);
xor U6481 (N_6481,N_6230,N_6330);
or U6482 (N_6482,N_6255,N_6333);
xnor U6483 (N_6483,N_6224,N_6332);
nand U6484 (N_6484,N_6321,N_6290);
or U6485 (N_6485,N_6310,N_6386);
and U6486 (N_6486,N_6374,N_6357);
nand U6487 (N_6487,N_6235,N_6376);
xnor U6488 (N_6488,N_6221,N_6275);
nand U6489 (N_6489,N_6393,N_6286);
nor U6490 (N_6490,N_6240,N_6352);
xor U6491 (N_6491,N_6267,N_6353);
and U6492 (N_6492,N_6244,N_6344);
or U6493 (N_6493,N_6215,N_6323);
nand U6494 (N_6494,N_6278,N_6246);
and U6495 (N_6495,N_6387,N_6241);
and U6496 (N_6496,N_6211,N_6263);
and U6497 (N_6497,N_6285,N_6325);
or U6498 (N_6498,N_6361,N_6302);
nand U6499 (N_6499,N_6379,N_6209);
and U6500 (N_6500,N_6304,N_6234);
nor U6501 (N_6501,N_6358,N_6287);
nor U6502 (N_6502,N_6325,N_6349);
nand U6503 (N_6503,N_6327,N_6226);
and U6504 (N_6504,N_6267,N_6236);
and U6505 (N_6505,N_6388,N_6332);
and U6506 (N_6506,N_6330,N_6246);
or U6507 (N_6507,N_6263,N_6371);
xor U6508 (N_6508,N_6254,N_6290);
xor U6509 (N_6509,N_6375,N_6239);
and U6510 (N_6510,N_6382,N_6338);
or U6511 (N_6511,N_6238,N_6317);
or U6512 (N_6512,N_6238,N_6379);
nand U6513 (N_6513,N_6291,N_6201);
nor U6514 (N_6514,N_6360,N_6240);
and U6515 (N_6515,N_6344,N_6307);
or U6516 (N_6516,N_6302,N_6272);
or U6517 (N_6517,N_6233,N_6235);
nand U6518 (N_6518,N_6204,N_6237);
nor U6519 (N_6519,N_6278,N_6234);
xnor U6520 (N_6520,N_6215,N_6234);
and U6521 (N_6521,N_6365,N_6318);
and U6522 (N_6522,N_6243,N_6323);
nand U6523 (N_6523,N_6334,N_6308);
and U6524 (N_6524,N_6392,N_6311);
nor U6525 (N_6525,N_6380,N_6385);
and U6526 (N_6526,N_6310,N_6214);
nand U6527 (N_6527,N_6366,N_6281);
nor U6528 (N_6528,N_6308,N_6388);
nand U6529 (N_6529,N_6278,N_6218);
nor U6530 (N_6530,N_6239,N_6213);
nor U6531 (N_6531,N_6213,N_6298);
and U6532 (N_6532,N_6335,N_6206);
nand U6533 (N_6533,N_6228,N_6249);
or U6534 (N_6534,N_6277,N_6204);
and U6535 (N_6535,N_6209,N_6351);
or U6536 (N_6536,N_6353,N_6248);
nor U6537 (N_6537,N_6382,N_6300);
nand U6538 (N_6538,N_6230,N_6336);
xor U6539 (N_6539,N_6378,N_6365);
xor U6540 (N_6540,N_6286,N_6389);
or U6541 (N_6541,N_6230,N_6267);
xor U6542 (N_6542,N_6273,N_6308);
nor U6543 (N_6543,N_6311,N_6332);
and U6544 (N_6544,N_6229,N_6345);
nand U6545 (N_6545,N_6350,N_6351);
or U6546 (N_6546,N_6350,N_6323);
nor U6547 (N_6547,N_6305,N_6236);
nand U6548 (N_6548,N_6306,N_6359);
nor U6549 (N_6549,N_6375,N_6380);
and U6550 (N_6550,N_6289,N_6237);
or U6551 (N_6551,N_6353,N_6250);
xor U6552 (N_6552,N_6346,N_6303);
or U6553 (N_6553,N_6282,N_6333);
and U6554 (N_6554,N_6232,N_6268);
nand U6555 (N_6555,N_6319,N_6389);
xnor U6556 (N_6556,N_6264,N_6324);
or U6557 (N_6557,N_6266,N_6259);
nand U6558 (N_6558,N_6376,N_6216);
and U6559 (N_6559,N_6220,N_6295);
nor U6560 (N_6560,N_6221,N_6397);
nor U6561 (N_6561,N_6391,N_6357);
nor U6562 (N_6562,N_6298,N_6345);
nand U6563 (N_6563,N_6302,N_6345);
or U6564 (N_6564,N_6395,N_6210);
nand U6565 (N_6565,N_6232,N_6389);
nor U6566 (N_6566,N_6332,N_6322);
nand U6567 (N_6567,N_6371,N_6306);
or U6568 (N_6568,N_6379,N_6297);
xnor U6569 (N_6569,N_6308,N_6319);
nand U6570 (N_6570,N_6314,N_6344);
or U6571 (N_6571,N_6320,N_6273);
nand U6572 (N_6572,N_6236,N_6218);
or U6573 (N_6573,N_6297,N_6216);
or U6574 (N_6574,N_6220,N_6372);
nand U6575 (N_6575,N_6221,N_6354);
and U6576 (N_6576,N_6350,N_6211);
nor U6577 (N_6577,N_6372,N_6333);
nand U6578 (N_6578,N_6322,N_6276);
nor U6579 (N_6579,N_6250,N_6294);
or U6580 (N_6580,N_6388,N_6362);
xnor U6581 (N_6581,N_6206,N_6399);
nor U6582 (N_6582,N_6274,N_6393);
and U6583 (N_6583,N_6248,N_6264);
xnor U6584 (N_6584,N_6336,N_6365);
or U6585 (N_6585,N_6211,N_6348);
nand U6586 (N_6586,N_6354,N_6251);
xor U6587 (N_6587,N_6378,N_6200);
nand U6588 (N_6588,N_6280,N_6317);
or U6589 (N_6589,N_6257,N_6283);
and U6590 (N_6590,N_6292,N_6275);
xor U6591 (N_6591,N_6336,N_6223);
xnor U6592 (N_6592,N_6349,N_6374);
or U6593 (N_6593,N_6282,N_6219);
xor U6594 (N_6594,N_6235,N_6255);
and U6595 (N_6595,N_6351,N_6360);
nand U6596 (N_6596,N_6217,N_6213);
or U6597 (N_6597,N_6336,N_6261);
or U6598 (N_6598,N_6383,N_6208);
or U6599 (N_6599,N_6329,N_6233);
nor U6600 (N_6600,N_6590,N_6526);
xor U6601 (N_6601,N_6456,N_6572);
and U6602 (N_6602,N_6549,N_6569);
xor U6603 (N_6603,N_6540,N_6525);
nand U6604 (N_6604,N_6518,N_6424);
or U6605 (N_6605,N_6442,N_6584);
or U6606 (N_6606,N_6560,N_6508);
and U6607 (N_6607,N_6513,N_6479);
xor U6608 (N_6608,N_6585,N_6514);
nand U6609 (N_6609,N_6594,N_6598);
nor U6610 (N_6610,N_6457,N_6470);
nand U6611 (N_6611,N_6480,N_6539);
xnor U6612 (N_6612,N_6472,N_6478);
nand U6613 (N_6613,N_6505,N_6571);
and U6614 (N_6614,N_6555,N_6524);
xnor U6615 (N_6615,N_6429,N_6586);
nand U6616 (N_6616,N_6577,N_6495);
nor U6617 (N_6617,N_6527,N_6402);
xor U6618 (N_6618,N_6499,N_6529);
and U6619 (N_6619,N_6484,N_6553);
and U6620 (N_6620,N_6474,N_6599);
xor U6621 (N_6621,N_6477,N_6556);
nor U6622 (N_6622,N_6522,N_6412);
and U6623 (N_6623,N_6596,N_6436);
nand U6624 (N_6624,N_6546,N_6548);
nor U6625 (N_6625,N_6578,N_6419);
xnor U6626 (N_6626,N_6515,N_6426);
or U6627 (N_6627,N_6592,N_6496);
nor U6628 (N_6628,N_6545,N_6587);
and U6629 (N_6629,N_6417,N_6427);
and U6630 (N_6630,N_6489,N_6543);
xnor U6631 (N_6631,N_6531,N_6454);
nand U6632 (N_6632,N_6512,N_6469);
or U6633 (N_6633,N_6400,N_6408);
xnor U6634 (N_6634,N_6475,N_6589);
nor U6635 (N_6635,N_6453,N_6583);
xnor U6636 (N_6636,N_6404,N_6523);
nor U6637 (N_6637,N_6559,N_6581);
xnor U6638 (N_6638,N_6554,N_6441);
or U6639 (N_6639,N_6542,N_6416);
or U6640 (N_6640,N_6401,N_6538);
nor U6641 (N_6641,N_6562,N_6503);
and U6642 (N_6642,N_6588,N_6485);
xor U6643 (N_6643,N_6593,N_6422);
nor U6644 (N_6644,N_6493,N_6445);
xor U6645 (N_6645,N_6551,N_6415);
xor U6646 (N_6646,N_6406,N_6520);
and U6647 (N_6647,N_6506,N_6434);
xor U6648 (N_6648,N_6521,N_6534);
xnor U6649 (N_6649,N_6440,N_6439);
and U6650 (N_6650,N_6530,N_6491);
xnor U6651 (N_6651,N_6411,N_6544);
nand U6652 (N_6652,N_6570,N_6430);
nand U6653 (N_6653,N_6482,N_6438);
nor U6654 (N_6654,N_6459,N_6446);
nand U6655 (N_6655,N_6494,N_6565);
xnor U6656 (N_6656,N_6533,N_6464);
nor U6657 (N_6657,N_6418,N_6580);
xor U6658 (N_6658,N_6448,N_6579);
xor U6659 (N_6659,N_6471,N_6490);
or U6660 (N_6660,N_6407,N_6447);
and U6661 (N_6661,N_6409,N_6547);
or U6662 (N_6662,N_6483,N_6425);
nor U6663 (N_6663,N_6516,N_6476);
or U6664 (N_6664,N_6443,N_6423);
nor U6665 (N_6665,N_6450,N_6566);
nor U6666 (N_6666,N_6458,N_6557);
and U6667 (N_6667,N_6486,N_6481);
or U6668 (N_6668,N_6410,N_6414);
nand U6669 (N_6669,N_6502,N_6455);
nand U6670 (N_6670,N_6403,N_6449);
nand U6671 (N_6671,N_6468,N_6509);
nand U6672 (N_6672,N_6552,N_6561);
xor U6673 (N_6673,N_6528,N_6519);
xor U6674 (N_6674,N_6517,N_6507);
or U6675 (N_6675,N_6487,N_6591);
nand U6676 (N_6676,N_6451,N_6510);
xnor U6677 (N_6677,N_6435,N_6421);
and U6678 (N_6678,N_6575,N_6597);
nand U6679 (N_6679,N_6563,N_6431);
or U6680 (N_6680,N_6500,N_6467);
nand U6681 (N_6681,N_6413,N_6576);
nor U6682 (N_6682,N_6504,N_6473);
xor U6683 (N_6683,N_6463,N_6574);
nor U6684 (N_6684,N_6537,N_6460);
nor U6685 (N_6685,N_6541,N_6432);
xnor U6686 (N_6686,N_6466,N_6452);
nor U6687 (N_6687,N_6535,N_6465);
xnor U6688 (N_6688,N_6564,N_6511);
and U6689 (N_6689,N_6444,N_6582);
nor U6690 (N_6690,N_6498,N_6492);
or U6691 (N_6691,N_6405,N_6573);
xnor U6692 (N_6692,N_6462,N_6532);
and U6693 (N_6693,N_6420,N_6550);
nand U6694 (N_6694,N_6461,N_6433);
xor U6695 (N_6695,N_6567,N_6497);
and U6696 (N_6696,N_6568,N_6428);
nor U6697 (N_6697,N_6595,N_6437);
and U6698 (N_6698,N_6501,N_6536);
or U6699 (N_6699,N_6558,N_6488);
xor U6700 (N_6700,N_6487,N_6496);
and U6701 (N_6701,N_6536,N_6496);
or U6702 (N_6702,N_6525,N_6517);
or U6703 (N_6703,N_6532,N_6565);
xnor U6704 (N_6704,N_6414,N_6545);
xor U6705 (N_6705,N_6587,N_6540);
nand U6706 (N_6706,N_6510,N_6558);
and U6707 (N_6707,N_6427,N_6591);
or U6708 (N_6708,N_6545,N_6494);
xor U6709 (N_6709,N_6501,N_6586);
and U6710 (N_6710,N_6548,N_6550);
xor U6711 (N_6711,N_6513,N_6549);
or U6712 (N_6712,N_6494,N_6551);
nand U6713 (N_6713,N_6487,N_6431);
or U6714 (N_6714,N_6556,N_6500);
and U6715 (N_6715,N_6475,N_6546);
or U6716 (N_6716,N_6463,N_6408);
nor U6717 (N_6717,N_6440,N_6562);
and U6718 (N_6718,N_6450,N_6507);
and U6719 (N_6719,N_6562,N_6495);
nand U6720 (N_6720,N_6432,N_6504);
xnor U6721 (N_6721,N_6580,N_6546);
nor U6722 (N_6722,N_6412,N_6537);
nor U6723 (N_6723,N_6521,N_6550);
nor U6724 (N_6724,N_6447,N_6558);
or U6725 (N_6725,N_6517,N_6595);
nor U6726 (N_6726,N_6417,N_6597);
nand U6727 (N_6727,N_6421,N_6520);
and U6728 (N_6728,N_6487,N_6517);
nand U6729 (N_6729,N_6577,N_6538);
or U6730 (N_6730,N_6494,N_6574);
xor U6731 (N_6731,N_6586,N_6492);
xnor U6732 (N_6732,N_6432,N_6585);
nor U6733 (N_6733,N_6557,N_6573);
nand U6734 (N_6734,N_6583,N_6566);
nand U6735 (N_6735,N_6484,N_6400);
and U6736 (N_6736,N_6466,N_6416);
xor U6737 (N_6737,N_6432,N_6426);
nand U6738 (N_6738,N_6407,N_6488);
xnor U6739 (N_6739,N_6558,N_6554);
or U6740 (N_6740,N_6467,N_6503);
nand U6741 (N_6741,N_6456,N_6581);
nor U6742 (N_6742,N_6546,N_6559);
xnor U6743 (N_6743,N_6579,N_6572);
nand U6744 (N_6744,N_6474,N_6492);
or U6745 (N_6745,N_6522,N_6535);
nand U6746 (N_6746,N_6453,N_6486);
or U6747 (N_6747,N_6530,N_6410);
nor U6748 (N_6748,N_6413,N_6482);
xor U6749 (N_6749,N_6499,N_6434);
nor U6750 (N_6750,N_6594,N_6578);
and U6751 (N_6751,N_6488,N_6579);
nand U6752 (N_6752,N_6504,N_6518);
and U6753 (N_6753,N_6439,N_6507);
nor U6754 (N_6754,N_6526,N_6507);
or U6755 (N_6755,N_6599,N_6463);
and U6756 (N_6756,N_6465,N_6436);
nand U6757 (N_6757,N_6587,N_6549);
and U6758 (N_6758,N_6454,N_6446);
nor U6759 (N_6759,N_6527,N_6517);
nor U6760 (N_6760,N_6463,N_6539);
nand U6761 (N_6761,N_6557,N_6553);
xnor U6762 (N_6762,N_6446,N_6447);
and U6763 (N_6763,N_6500,N_6434);
nand U6764 (N_6764,N_6591,N_6540);
nand U6765 (N_6765,N_6460,N_6583);
xnor U6766 (N_6766,N_6594,N_6421);
or U6767 (N_6767,N_6571,N_6526);
xnor U6768 (N_6768,N_6573,N_6451);
nand U6769 (N_6769,N_6535,N_6411);
or U6770 (N_6770,N_6415,N_6424);
or U6771 (N_6771,N_6467,N_6577);
and U6772 (N_6772,N_6437,N_6429);
or U6773 (N_6773,N_6599,N_6548);
or U6774 (N_6774,N_6406,N_6474);
nand U6775 (N_6775,N_6442,N_6525);
nor U6776 (N_6776,N_6517,N_6446);
and U6777 (N_6777,N_6461,N_6597);
and U6778 (N_6778,N_6454,N_6594);
or U6779 (N_6779,N_6516,N_6547);
and U6780 (N_6780,N_6419,N_6538);
xor U6781 (N_6781,N_6475,N_6441);
nor U6782 (N_6782,N_6593,N_6457);
xnor U6783 (N_6783,N_6466,N_6585);
and U6784 (N_6784,N_6432,N_6495);
nor U6785 (N_6785,N_6519,N_6490);
and U6786 (N_6786,N_6449,N_6407);
nor U6787 (N_6787,N_6501,N_6485);
and U6788 (N_6788,N_6433,N_6457);
nor U6789 (N_6789,N_6495,N_6493);
nand U6790 (N_6790,N_6442,N_6435);
nand U6791 (N_6791,N_6517,N_6510);
nand U6792 (N_6792,N_6480,N_6579);
and U6793 (N_6793,N_6558,N_6420);
or U6794 (N_6794,N_6409,N_6426);
or U6795 (N_6795,N_6541,N_6576);
nand U6796 (N_6796,N_6436,N_6416);
or U6797 (N_6797,N_6485,N_6410);
and U6798 (N_6798,N_6410,N_6446);
and U6799 (N_6799,N_6410,N_6451);
or U6800 (N_6800,N_6662,N_6650);
and U6801 (N_6801,N_6749,N_6648);
and U6802 (N_6802,N_6631,N_6776);
or U6803 (N_6803,N_6767,N_6728);
nand U6804 (N_6804,N_6654,N_6768);
nand U6805 (N_6805,N_6640,N_6669);
xnor U6806 (N_6806,N_6794,N_6651);
nor U6807 (N_6807,N_6684,N_6762);
and U6808 (N_6808,N_6618,N_6619);
xor U6809 (N_6809,N_6686,N_6740);
xor U6810 (N_6810,N_6642,N_6629);
nand U6811 (N_6811,N_6663,N_6770);
nor U6812 (N_6812,N_6699,N_6710);
nand U6813 (N_6813,N_6692,N_6688);
and U6814 (N_6814,N_6636,N_6644);
nand U6815 (N_6815,N_6639,N_6726);
and U6816 (N_6816,N_6681,N_6622);
xor U6817 (N_6817,N_6623,N_6687);
nand U6818 (N_6818,N_6665,N_6779);
or U6819 (N_6819,N_6750,N_6709);
nor U6820 (N_6820,N_6700,N_6691);
xnor U6821 (N_6821,N_6731,N_6707);
or U6822 (N_6822,N_6689,N_6675);
and U6823 (N_6823,N_6628,N_6753);
nand U6824 (N_6824,N_6676,N_6652);
nand U6825 (N_6825,N_6733,N_6714);
or U6826 (N_6826,N_6789,N_6765);
or U6827 (N_6827,N_6715,N_6772);
nor U6828 (N_6828,N_6778,N_6633);
and U6829 (N_6829,N_6612,N_6730);
nand U6830 (N_6830,N_6664,N_6655);
and U6831 (N_6831,N_6603,N_6696);
and U6832 (N_6832,N_6754,N_6683);
nand U6833 (N_6833,N_6751,N_6799);
or U6834 (N_6834,N_6725,N_6624);
or U6835 (N_6835,N_6713,N_6634);
nor U6836 (N_6836,N_6656,N_6620);
xor U6837 (N_6837,N_6744,N_6784);
and U6838 (N_6838,N_6788,N_6600);
xnor U6839 (N_6839,N_6758,N_6705);
or U6840 (N_6840,N_6679,N_6658);
and U6841 (N_6841,N_6660,N_6748);
nor U6842 (N_6842,N_6601,N_6611);
nand U6843 (N_6843,N_6605,N_6617);
nor U6844 (N_6844,N_6697,N_6775);
nor U6845 (N_6845,N_6674,N_6785);
nand U6846 (N_6846,N_6786,N_6614);
and U6847 (N_6847,N_6649,N_6616);
nand U6848 (N_6848,N_6659,N_6630);
or U6849 (N_6849,N_6791,N_6737);
and U6850 (N_6850,N_6701,N_6635);
nor U6851 (N_6851,N_6613,N_6747);
nand U6852 (N_6852,N_6643,N_6678);
xnor U6853 (N_6853,N_6717,N_6718);
nor U6854 (N_6854,N_6780,N_6706);
or U6855 (N_6855,N_6766,N_6774);
or U6856 (N_6856,N_6720,N_6698);
xor U6857 (N_6857,N_6761,N_6738);
or U6858 (N_6858,N_6690,N_6797);
or U6859 (N_6859,N_6657,N_6661);
or U6860 (N_6860,N_6702,N_6615);
and U6861 (N_6861,N_6756,N_6742);
and U6862 (N_6862,N_6666,N_6653);
xnor U6863 (N_6863,N_6695,N_6741);
xnor U6864 (N_6864,N_6637,N_6783);
and U6865 (N_6865,N_6781,N_6773);
nor U6866 (N_6866,N_6608,N_6757);
xor U6867 (N_6867,N_6682,N_6743);
nor U6868 (N_6868,N_6724,N_6793);
nor U6869 (N_6869,N_6712,N_6673);
nor U6870 (N_6870,N_6752,N_6764);
nand U6871 (N_6871,N_6711,N_6645);
and U6872 (N_6872,N_6693,N_6703);
or U6873 (N_6873,N_6668,N_6771);
and U6874 (N_6874,N_6796,N_6722);
nand U6875 (N_6875,N_6739,N_6708);
and U6876 (N_6876,N_6604,N_6647);
and U6877 (N_6877,N_6646,N_6723);
and U6878 (N_6878,N_6680,N_6719);
or U6879 (N_6879,N_6759,N_6625);
nor U6880 (N_6880,N_6704,N_6798);
xor U6881 (N_6881,N_6609,N_6736);
and U6882 (N_6882,N_6792,N_6777);
nor U6883 (N_6883,N_6602,N_6626);
nor U6884 (N_6884,N_6760,N_6621);
nor U6885 (N_6885,N_6746,N_6694);
or U6886 (N_6886,N_6721,N_6732);
nand U6887 (N_6887,N_6638,N_6641);
nor U6888 (N_6888,N_6769,N_6734);
or U6889 (N_6889,N_6677,N_6672);
nand U6890 (N_6890,N_6716,N_6727);
nor U6891 (N_6891,N_6607,N_6632);
xor U6892 (N_6892,N_6610,N_6627);
and U6893 (N_6893,N_6729,N_6671);
or U6894 (N_6894,N_6735,N_6787);
and U6895 (N_6895,N_6667,N_6745);
nand U6896 (N_6896,N_6670,N_6685);
nand U6897 (N_6897,N_6755,N_6790);
and U6898 (N_6898,N_6795,N_6606);
nand U6899 (N_6899,N_6782,N_6763);
and U6900 (N_6900,N_6715,N_6624);
nor U6901 (N_6901,N_6702,N_6614);
nand U6902 (N_6902,N_6718,N_6796);
nor U6903 (N_6903,N_6703,N_6782);
or U6904 (N_6904,N_6733,N_6682);
nor U6905 (N_6905,N_6657,N_6668);
or U6906 (N_6906,N_6686,N_6610);
or U6907 (N_6907,N_6763,N_6691);
xor U6908 (N_6908,N_6630,N_6744);
nor U6909 (N_6909,N_6780,N_6674);
or U6910 (N_6910,N_6674,N_6765);
nor U6911 (N_6911,N_6657,N_6788);
and U6912 (N_6912,N_6683,N_6715);
nand U6913 (N_6913,N_6781,N_6672);
xnor U6914 (N_6914,N_6681,N_6728);
or U6915 (N_6915,N_6661,N_6603);
and U6916 (N_6916,N_6717,N_6728);
and U6917 (N_6917,N_6650,N_6750);
or U6918 (N_6918,N_6715,N_6734);
nor U6919 (N_6919,N_6652,N_6626);
or U6920 (N_6920,N_6700,N_6704);
and U6921 (N_6921,N_6675,N_6789);
nor U6922 (N_6922,N_6601,N_6767);
xnor U6923 (N_6923,N_6666,N_6792);
nor U6924 (N_6924,N_6660,N_6635);
or U6925 (N_6925,N_6679,N_6716);
nand U6926 (N_6926,N_6745,N_6743);
nor U6927 (N_6927,N_6709,N_6684);
xnor U6928 (N_6928,N_6650,N_6693);
nand U6929 (N_6929,N_6693,N_6750);
or U6930 (N_6930,N_6716,N_6628);
nor U6931 (N_6931,N_6617,N_6731);
nand U6932 (N_6932,N_6705,N_6794);
or U6933 (N_6933,N_6722,N_6621);
nor U6934 (N_6934,N_6756,N_6738);
and U6935 (N_6935,N_6780,N_6622);
xor U6936 (N_6936,N_6611,N_6658);
nand U6937 (N_6937,N_6666,N_6721);
or U6938 (N_6938,N_6721,N_6761);
xnor U6939 (N_6939,N_6719,N_6778);
or U6940 (N_6940,N_6679,N_6687);
nor U6941 (N_6941,N_6795,N_6778);
nor U6942 (N_6942,N_6628,N_6608);
or U6943 (N_6943,N_6794,N_6623);
and U6944 (N_6944,N_6696,N_6702);
or U6945 (N_6945,N_6719,N_6692);
or U6946 (N_6946,N_6772,N_6729);
or U6947 (N_6947,N_6793,N_6645);
nand U6948 (N_6948,N_6783,N_6625);
nand U6949 (N_6949,N_6715,N_6774);
nor U6950 (N_6950,N_6770,N_6660);
nand U6951 (N_6951,N_6748,N_6753);
or U6952 (N_6952,N_6689,N_6768);
nand U6953 (N_6953,N_6653,N_6649);
or U6954 (N_6954,N_6788,N_6753);
or U6955 (N_6955,N_6665,N_6731);
nor U6956 (N_6956,N_6778,N_6792);
xor U6957 (N_6957,N_6702,N_6706);
or U6958 (N_6958,N_6668,N_6610);
nand U6959 (N_6959,N_6662,N_6788);
and U6960 (N_6960,N_6715,N_6746);
or U6961 (N_6961,N_6662,N_6698);
or U6962 (N_6962,N_6616,N_6735);
or U6963 (N_6963,N_6771,N_6696);
nor U6964 (N_6964,N_6760,N_6734);
nor U6965 (N_6965,N_6651,N_6786);
nand U6966 (N_6966,N_6738,N_6791);
xor U6967 (N_6967,N_6799,N_6691);
nand U6968 (N_6968,N_6744,N_6785);
nor U6969 (N_6969,N_6614,N_6608);
xnor U6970 (N_6970,N_6712,N_6720);
nor U6971 (N_6971,N_6749,N_6798);
nand U6972 (N_6972,N_6769,N_6650);
nor U6973 (N_6973,N_6767,N_6632);
and U6974 (N_6974,N_6740,N_6667);
nand U6975 (N_6975,N_6601,N_6770);
and U6976 (N_6976,N_6664,N_6687);
xor U6977 (N_6977,N_6698,N_6763);
nand U6978 (N_6978,N_6636,N_6681);
nand U6979 (N_6979,N_6689,N_6766);
or U6980 (N_6980,N_6647,N_6665);
nor U6981 (N_6981,N_6640,N_6644);
and U6982 (N_6982,N_6602,N_6631);
or U6983 (N_6983,N_6720,N_6605);
xor U6984 (N_6984,N_6752,N_6667);
nand U6985 (N_6985,N_6700,N_6612);
nor U6986 (N_6986,N_6703,N_6709);
nor U6987 (N_6987,N_6665,N_6727);
nor U6988 (N_6988,N_6729,N_6789);
xnor U6989 (N_6989,N_6779,N_6602);
and U6990 (N_6990,N_6687,N_6772);
nand U6991 (N_6991,N_6710,N_6649);
and U6992 (N_6992,N_6663,N_6772);
nand U6993 (N_6993,N_6683,N_6684);
xnor U6994 (N_6994,N_6755,N_6627);
or U6995 (N_6995,N_6786,N_6668);
nor U6996 (N_6996,N_6680,N_6710);
xnor U6997 (N_6997,N_6772,N_6601);
nor U6998 (N_6998,N_6622,N_6753);
or U6999 (N_6999,N_6718,N_6741);
and U7000 (N_7000,N_6907,N_6963);
and U7001 (N_7001,N_6829,N_6837);
nor U7002 (N_7002,N_6964,N_6816);
xnor U7003 (N_7003,N_6913,N_6947);
and U7004 (N_7004,N_6958,N_6950);
or U7005 (N_7005,N_6868,N_6967);
nand U7006 (N_7006,N_6831,N_6838);
nor U7007 (N_7007,N_6874,N_6921);
or U7008 (N_7008,N_6880,N_6915);
or U7009 (N_7009,N_6849,N_6995);
nand U7010 (N_7010,N_6982,N_6832);
xor U7011 (N_7011,N_6997,N_6961);
and U7012 (N_7012,N_6936,N_6830);
or U7013 (N_7013,N_6973,N_6949);
nand U7014 (N_7014,N_6979,N_6955);
nand U7015 (N_7015,N_6905,N_6891);
nor U7016 (N_7016,N_6910,N_6878);
xnor U7017 (N_7017,N_6861,N_6933);
and U7018 (N_7018,N_6909,N_6962);
xnor U7019 (N_7019,N_6946,N_6866);
nor U7020 (N_7020,N_6920,N_6990);
nand U7021 (N_7021,N_6869,N_6810);
xor U7022 (N_7022,N_6820,N_6917);
nor U7023 (N_7023,N_6835,N_6833);
or U7024 (N_7024,N_6911,N_6846);
nor U7025 (N_7025,N_6806,N_6983);
and U7026 (N_7026,N_6894,N_6814);
or U7027 (N_7027,N_6988,N_6822);
or U7028 (N_7028,N_6970,N_6914);
nor U7029 (N_7029,N_6938,N_6918);
xor U7030 (N_7030,N_6904,N_6931);
and U7031 (N_7031,N_6934,N_6939);
xnor U7032 (N_7032,N_6898,N_6848);
xnor U7033 (N_7033,N_6850,N_6986);
and U7034 (N_7034,N_6900,N_6875);
or U7035 (N_7035,N_6935,N_6926);
nand U7036 (N_7036,N_6801,N_6828);
and U7037 (N_7037,N_6940,N_6937);
xor U7038 (N_7038,N_6867,N_6860);
and U7039 (N_7039,N_6877,N_6932);
xnor U7040 (N_7040,N_6889,N_6927);
or U7041 (N_7041,N_6890,N_6992);
nor U7042 (N_7042,N_6865,N_6882);
xnor U7043 (N_7043,N_6976,N_6808);
or U7044 (N_7044,N_6859,N_6948);
nor U7045 (N_7045,N_6841,N_6923);
xor U7046 (N_7046,N_6998,N_6968);
or U7047 (N_7047,N_6811,N_6944);
or U7048 (N_7048,N_6842,N_6881);
xnor U7049 (N_7049,N_6834,N_6888);
nor U7050 (N_7050,N_6984,N_6978);
nor U7051 (N_7051,N_6928,N_6972);
nor U7052 (N_7052,N_6942,N_6980);
nand U7053 (N_7053,N_6912,N_6953);
nand U7054 (N_7054,N_6965,N_6817);
and U7055 (N_7055,N_6922,N_6969);
nand U7056 (N_7056,N_6993,N_6805);
nand U7057 (N_7057,N_6886,N_6899);
and U7058 (N_7058,N_6892,N_6809);
nand U7059 (N_7059,N_6908,N_6919);
nand U7060 (N_7060,N_6873,N_6857);
nand U7061 (N_7061,N_6959,N_6893);
and U7062 (N_7062,N_6956,N_6856);
xnor U7063 (N_7063,N_6844,N_6903);
or U7064 (N_7064,N_6839,N_6852);
nor U7065 (N_7065,N_6952,N_6924);
nor U7066 (N_7066,N_6800,N_6826);
xnor U7067 (N_7067,N_6985,N_6804);
xnor U7068 (N_7068,N_6854,N_6960);
nor U7069 (N_7069,N_6845,N_6925);
nand U7070 (N_7070,N_6971,N_6836);
nor U7071 (N_7071,N_6819,N_6902);
xor U7072 (N_7072,N_6858,N_6813);
or U7073 (N_7073,N_6863,N_6807);
or U7074 (N_7074,N_6876,N_6929);
nand U7075 (N_7075,N_6840,N_6855);
or U7076 (N_7076,N_6824,N_6974);
or U7077 (N_7077,N_6941,N_6930);
nand U7078 (N_7078,N_6870,N_6885);
and U7079 (N_7079,N_6987,N_6847);
nand U7080 (N_7080,N_6887,N_6943);
xor U7081 (N_7081,N_6966,N_6871);
nand U7082 (N_7082,N_6879,N_6851);
and U7083 (N_7083,N_6981,N_6872);
and U7084 (N_7084,N_6954,N_6975);
nor U7085 (N_7085,N_6901,N_6812);
xor U7086 (N_7086,N_6916,N_6883);
nor U7087 (N_7087,N_6864,N_6996);
and U7088 (N_7088,N_6821,N_6827);
and U7089 (N_7089,N_6957,N_6991);
nor U7090 (N_7090,N_6977,N_6825);
and U7091 (N_7091,N_6802,N_6896);
nand U7092 (N_7092,N_6897,N_6823);
nand U7093 (N_7093,N_6853,N_6999);
or U7094 (N_7094,N_6906,N_6818);
and U7095 (N_7095,N_6815,N_6994);
xor U7096 (N_7096,N_6884,N_6951);
and U7097 (N_7097,N_6895,N_6989);
nor U7098 (N_7098,N_6803,N_6843);
nor U7099 (N_7099,N_6945,N_6862);
or U7100 (N_7100,N_6871,N_6987);
or U7101 (N_7101,N_6900,N_6865);
xnor U7102 (N_7102,N_6893,N_6904);
and U7103 (N_7103,N_6876,N_6968);
nand U7104 (N_7104,N_6860,N_6838);
and U7105 (N_7105,N_6813,N_6931);
nand U7106 (N_7106,N_6832,N_6949);
nand U7107 (N_7107,N_6852,N_6812);
nand U7108 (N_7108,N_6962,N_6964);
nor U7109 (N_7109,N_6839,N_6895);
or U7110 (N_7110,N_6955,N_6885);
and U7111 (N_7111,N_6913,N_6849);
nand U7112 (N_7112,N_6905,N_6973);
nand U7113 (N_7113,N_6998,N_6990);
and U7114 (N_7114,N_6869,N_6974);
xor U7115 (N_7115,N_6872,N_6862);
and U7116 (N_7116,N_6918,N_6923);
nor U7117 (N_7117,N_6976,N_6912);
and U7118 (N_7118,N_6829,N_6832);
nand U7119 (N_7119,N_6840,N_6971);
or U7120 (N_7120,N_6970,N_6903);
and U7121 (N_7121,N_6950,N_6875);
and U7122 (N_7122,N_6945,N_6936);
or U7123 (N_7123,N_6962,N_6818);
nand U7124 (N_7124,N_6840,N_6984);
xor U7125 (N_7125,N_6981,N_6890);
or U7126 (N_7126,N_6936,N_6813);
and U7127 (N_7127,N_6908,N_6977);
or U7128 (N_7128,N_6983,N_6940);
and U7129 (N_7129,N_6849,N_6923);
xnor U7130 (N_7130,N_6859,N_6804);
nor U7131 (N_7131,N_6829,N_6850);
nand U7132 (N_7132,N_6873,N_6865);
xor U7133 (N_7133,N_6806,N_6859);
nor U7134 (N_7134,N_6867,N_6885);
nand U7135 (N_7135,N_6843,N_6991);
or U7136 (N_7136,N_6990,N_6914);
xnor U7137 (N_7137,N_6867,N_6953);
nand U7138 (N_7138,N_6817,N_6826);
xor U7139 (N_7139,N_6949,N_6970);
and U7140 (N_7140,N_6968,N_6882);
nand U7141 (N_7141,N_6826,N_6845);
nand U7142 (N_7142,N_6842,N_6920);
or U7143 (N_7143,N_6984,N_6887);
nand U7144 (N_7144,N_6957,N_6859);
xnor U7145 (N_7145,N_6962,N_6922);
nor U7146 (N_7146,N_6891,N_6902);
nor U7147 (N_7147,N_6848,N_6977);
nand U7148 (N_7148,N_6931,N_6932);
nand U7149 (N_7149,N_6904,N_6838);
nor U7150 (N_7150,N_6878,N_6889);
nor U7151 (N_7151,N_6930,N_6954);
and U7152 (N_7152,N_6802,N_6994);
and U7153 (N_7153,N_6930,N_6851);
or U7154 (N_7154,N_6939,N_6827);
and U7155 (N_7155,N_6836,N_6976);
xor U7156 (N_7156,N_6841,N_6965);
nand U7157 (N_7157,N_6921,N_6907);
nor U7158 (N_7158,N_6836,N_6904);
and U7159 (N_7159,N_6970,N_6895);
nor U7160 (N_7160,N_6911,N_6913);
and U7161 (N_7161,N_6865,N_6953);
xor U7162 (N_7162,N_6820,N_6900);
nand U7163 (N_7163,N_6811,N_6806);
nand U7164 (N_7164,N_6893,N_6883);
xnor U7165 (N_7165,N_6918,N_6877);
and U7166 (N_7166,N_6828,N_6833);
and U7167 (N_7167,N_6885,N_6903);
xor U7168 (N_7168,N_6883,N_6873);
and U7169 (N_7169,N_6820,N_6868);
xor U7170 (N_7170,N_6981,N_6883);
xor U7171 (N_7171,N_6945,N_6930);
or U7172 (N_7172,N_6948,N_6856);
nand U7173 (N_7173,N_6845,N_6879);
nor U7174 (N_7174,N_6812,N_6998);
and U7175 (N_7175,N_6821,N_6894);
and U7176 (N_7176,N_6828,N_6848);
nand U7177 (N_7177,N_6848,N_6976);
and U7178 (N_7178,N_6855,N_6941);
or U7179 (N_7179,N_6908,N_6867);
nor U7180 (N_7180,N_6858,N_6817);
nand U7181 (N_7181,N_6808,N_6856);
nor U7182 (N_7182,N_6984,N_6820);
xnor U7183 (N_7183,N_6833,N_6930);
and U7184 (N_7184,N_6820,N_6931);
or U7185 (N_7185,N_6962,N_6899);
nand U7186 (N_7186,N_6814,N_6925);
nor U7187 (N_7187,N_6881,N_6894);
nand U7188 (N_7188,N_6935,N_6937);
or U7189 (N_7189,N_6810,N_6879);
and U7190 (N_7190,N_6864,N_6987);
xnor U7191 (N_7191,N_6883,N_6823);
nand U7192 (N_7192,N_6909,N_6841);
xnor U7193 (N_7193,N_6937,N_6894);
and U7194 (N_7194,N_6802,N_6853);
xnor U7195 (N_7195,N_6899,N_6918);
or U7196 (N_7196,N_6910,N_6960);
and U7197 (N_7197,N_6909,N_6842);
xnor U7198 (N_7198,N_6930,N_6986);
and U7199 (N_7199,N_6992,N_6833);
xor U7200 (N_7200,N_7012,N_7180);
and U7201 (N_7201,N_7147,N_7135);
nor U7202 (N_7202,N_7165,N_7081);
nand U7203 (N_7203,N_7150,N_7108);
or U7204 (N_7204,N_7064,N_7030);
and U7205 (N_7205,N_7092,N_7152);
nor U7206 (N_7206,N_7025,N_7063);
or U7207 (N_7207,N_7134,N_7123);
or U7208 (N_7208,N_7074,N_7115);
and U7209 (N_7209,N_7102,N_7166);
xor U7210 (N_7210,N_7097,N_7111);
and U7211 (N_7211,N_7083,N_7021);
nor U7212 (N_7212,N_7154,N_7181);
nand U7213 (N_7213,N_7185,N_7119);
xnor U7214 (N_7214,N_7141,N_7007);
nor U7215 (N_7215,N_7172,N_7036);
or U7216 (N_7216,N_7197,N_7067);
nand U7217 (N_7217,N_7171,N_7062);
and U7218 (N_7218,N_7029,N_7056);
or U7219 (N_7219,N_7043,N_7051);
xor U7220 (N_7220,N_7184,N_7131);
nand U7221 (N_7221,N_7148,N_7018);
xnor U7222 (N_7222,N_7168,N_7075);
nand U7223 (N_7223,N_7140,N_7109);
xnor U7224 (N_7224,N_7085,N_7035);
nand U7225 (N_7225,N_7122,N_7020);
xor U7226 (N_7226,N_7041,N_7077);
and U7227 (N_7227,N_7189,N_7159);
and U7228 (N_7228,N_7026,N_7016);
xnor U7229 (N_7229,N_7090,N_7101);
xor U7230 (N_7230,N_7130,N_7065);
xor U7231 (N_7231,N_7046,N_7044);
nand U7232 (N_7232,N_7006,N_7014);
or U7233 (N_7233,N_7151,N_7017);
nand U7234 (N_7234,N_7124,N_7003);
nand U7235 (N_7235,N_7001,N_7023);
or U7236 (N_7236,N_7005,N_7186);
nor U7237 (N_7237,N_7175,N_7027);
and U7238 (N_7238,N_7053,N_7091);
nand U7239 (N_7239,N_7069,N_7072);
nand U7240 (N_7240,N_7137,N_7049);
and U7241 (N_7241,N_7022,N_7133);
nor U7242 (N_7242,N_7191,N_7011);
xnor U7243 (N_7243,N_7161,N_7073);
or U7244 (N_7244,N_7132,N_7104);
xnor U7245 (N_7245,N_7088,N_7037);
nand U7246 (N_7246,N_7176,N_7099);
nand U7247 (N_7247,N_7169,N_7028);
and U7248 (N_7248,N_7008,N_7094);
nand U7249 (N_7249,N_7079,N_7173);
nand U7250 (N_7250,N_7183,N_7127);
or U7251 (N_7251,N_7125,N_7019);
nand U7252 (N_7252,N_7149,N_7103);
or U7253 (N_7253,N_7004,N_7162);
nand U7254 (N_7254,N_7057,N_7178);
xnor U7255 (N_7255,N_7114,N_7084);
or U7256 (N_7256,N_7070,N_7059);
nor U7257 (N_7257,N_7066,N_7199);
nand U7258 (N_7258,N_7117,N_7187);
or U7259 (N_7259,N_7071,N_7100);
and U7260 (N_7260,N_7047,N_7060);
xor U7261 (N_7261,N_7136,N_7196);
nand U7262 (N_7262,N_7156,N_7188);
nand U7263 (N_7263,N_7034,N_7120);
and U7264 (N_7264,N_7153,N_7086);
and U7265 (N_7265,N_7042,N_7095);
or U7266 (N_7266,N_7009,N_7192);
nand U7267 (N_7267,N_7048,N_7055);
nor U7268 (N_7268,N_7015,N_7010);
nand U7269 (N_7269,N_7128,N_7198);
xnor U7270 (N_7270,N_7052,N_7000);
or U7271 (N_7271,N_7076,N_7082);
xnor U7272 (N_7272,N_7157,N_7058);
xor U7273 (N_7273,N_7144,N_7142);
or U7274 (N_7274,N_7174,N_7045);
and U7275 (N_7275,N_7096,N_7129);
nand U7276 (N_7276,N_7032,N_7080);
xnor U7277 (N_7277,N_7105,N_7013);
nor U7278 (N_7278,N_7039,N_7160);
and U7279 (N_7279,N_7164,N_7163);
and U7280 (N_7280,N_7106,N_7054);
or U7281 (N_7281,N_7033,N_7193);
xor U7282 (N_7282,N_7118,N_7050);
xor U7283 (N_7283,N_7113,N_7170);
nor U7284 (N_7284,N_7107,N_7112);
xor U7285 (N_7285,N_7061,N_7182);
nor U7286 (N_7286,N_7143,N_7126);
xor U7287 (N_7287,N_7040,N_7089);
or U7288 (N_7288,N_7179,N_7098);
nand U7289 (N_7289,N_7146,N_7110);
xnor U7290 (N_7290,N_7155,N_7068);
xnor U7291 (N_7291,N_7002,N_7190);
and U7292 (N_7292,N_7078,N_7145);
nor U7293 (N_7293,N_7195,N_7167);
or U7294 (N_7294,N_7194,N_7093);
and U7295 (N_7295,N_7177,N_7158);
and U7296 (N_7296,N_7087,N_7121);
and U7297 (N_7297,N_7139,N_7138);
nand U7298 (N_7298,N_7031,N_7038);
nor U7299 (N_7299,N_7024,N_7116);
xnor U7300 (N_7300,N_7183,N_7085);
or U7301 (N_7301,N_7023,N_7098);
and U7302 (N_7302,N_7070,N_7026);
and U7303 (N_7303,N_7147,N_7098);
nand U7304 (N_7304,N_7095,N_7002);
xnor U7305 (N_7305,N_7147,N_7118);
xor U7306 (N_7306,N_7134,N_7055);
or U7307 (N_7307,N_7103,N_7189);
nand U7308 (N_7308,N_7194,N_7010);
nand U7309 (N_7309,N_7006,N_7143);
nand U7310 (N_7310,N_7097,N_7038);
xnor U7311 (N_7311,N_7139,N_7116);
nor U7312 (N_7312,N_7022,N_7053);
and U7313 (N_7313,N_7115,N_7083);
nor U7314 (N_7314,N_7021,N_7075);
or U7315 (N_7315,N_7015,N_7114);
and U7316 (N_7316,N_7060,N_7044);
and U7317 (N_7317,N_7178,N_7068);
or U7318 (N_7318,N_7030,N_7087);
nand U7319 (N_7319,N_7117,N_7100);
xnor U7320 (N_7320,N_7016,N_7192);
nand U7321 (N_7321,N_7169,N_7156);
xor U7322 (N_7322,N_7093,N_7196);
nor U7323 (N_7323,N_7088,N_7177);
or U7324 (N_7324,N_7145,N_7002);
nand U7325 (N_7325,N_7155,N_7038);
nor U7326 (N_7326,N_7181,N_7170);
nor U7327 (N_7327,N_7037,N_7047);
and U7328 (N_7328,N_7198,N_7163);
xor U7329 (N_7329,N_7085,N_7093);
nor U7330 (N_7330,N_7114,N_7180);
and U7331 (N_7331,N_7128,N_7186);
or U7332 (N_7332,N_7193,N_7121);
nor U7333 (N_7333,N_7047,N_7140);
xor U7334 (N_7334,N_7022,N_7109);
or U7335 (N_7335,N_7173,N_7192);
and U7336 (N_7336,N_7012,N_7011);
or U7337 (N_7337,N_7014,N_7178);
nand U7338 (N_7338,N_7021,N_7073);
xnor U7339 (N_7339,N_7108,N_7173);
xor U7340 (N_7340,N_7104,N_7180);
or U7341 (N_7341,N_7129,N_7080);
nand U7342 (N_7342,N_7182,N_7149);
and U7343 (N_7343,N_7004,N_7040);
and U7344 (N_7344,N_7011,N_7136);
and U7345 (N_7345,N_7084,N_7163);
nor U7346 (N_7346,N_7118,N_7047);
nand U7347 (N_7347,N_7026,N_7006);
nand U7348 (N_7348,N_7170,N_7107);
xor U7349 (N_7349,N_7147,N_7164);
xor U7350 (N_7350,N_7166,N_7176);
or U7351 (N_7351,N_7153,N_7063);
or U7352 (N_7352,N_7160,N_7101);
or U7353 (N_7353,N_7114,N_7199);
nor U7354 (N_7354,N_7109,N_7095);
and U7355 (N_7355,N_7019,N_7151);
xor U7356 (N_7356,N_7195,N_7099);
or U7357 (N_7357,N_7146,N_7024);
nor U7358 (N_7358,N_7148,N_7095);
nor U7359 (N_7359,N_7011,N_7088);
and U7360 (N_7360,N_7042,N_7046);
xnor U7361 (N_7361,N_7055,N_7179);
nor U7362 (N_7362,N_7090,N_7084);
or U7363 (N_7363,N_7010,N_7196);
or U7364 (N_7364,N_7158,N_7121);
and U7365 (N_7365,N_7182,N_7125);
nand U7366 (N_7366,N_7077,N_7074);
xor U7367 (N_7367,N_7018,N_7015);
or U7368 (N_7368,N_7002,N_7114);
and U7369 (N_7369,N_7114,N_7097);
or U7370 (N_7370,N_7127,N_7125);
nor U7371 (N_7371,N_7191,N_7022);
or U7372 (N_7372,N_7021,N_7051);
or U7373 (N_7373,N_7066,N_7132);
or U7374 (N_7374,N_7071,N_7199);
nor U7375 (N_7375,N_7091,N_7142);
nor U7376 (N_7376,N_7181,N_7137);
xor U7377 (N_7377,N_7139,N_7124);
and U7378 (N_7378,N_7003,N_7041);
nor U7379 (N_7379,N_7007,N_7055);
xnor U7380 (N_7380,N_7026,N_7077);
nor U7381 (N_7381,N_7028,N_7145);
nor U7382 (N_7382,N_7147,N_7179);
or U7383 (N_7383,N_7160,N_7137);
or U7384 (N_7384,N_7166,N_7153);
and U7385 (N_7385,N_7161,N_7104);
nor U7386 (N_7386,N_7007,N_7107);
or U7387 (N_7387,N_7092,N_7062);
nand U7388 (N_7388,N_7050,N_7091);
nor U7389 (N_7389,N_7047,N_7061);
nor U7390 (N_7390,N_7169,N_7117);
xnor U7391 (N_7391,N_7026,N_7192);
or U7392 (N_7392,N_7041,N_7139);
nand U7393 (N_7393,N_7035,N_7089);
nor U7394 (N_7394,N_7012,N_7120);
or U7395 (N_7395,N_7064,N_7021);
and U7396 (N_7396,N_7182,N_7126);
xnor U7397 (N_7397,N_7119,N_7002);
and U7398 (N_7398,N_7055,N_7001);
nand U7399 (N_7399,N_7180,N_7165);
and U7400 (N_7400,N_7210,N_7365);
xor U7401 (N_7401,N_7315,N_7352);
or U7402 (N_7402,N_7230,N_7289);
and U7403 (N_7403,N_7380,N_7209);
nand U7404 (N_7404,N_7261,N_7207);
or U7405 (N_7405,N_7258,N_7346);
and U7406 (N_7406,N_7322,N_7313);
xnor U7407 (N_7407,N_7341,N_7375);
xnor U7408 (N_7408,N_7343,N_7299);
or U7409 (N_7409,N_7269,N_7392);
or U7410 (N_7410,N_7281,N_7353);
nor U7411 (N_7411,N_7287,N_7300);
or U7412 (N_7412,N_7381,N_7387);
xnor U7413 (N_7413,N_7208,N_7275);
or U7414 (N_7414,N_7271,N_7323);
nand U7415 (N_7415,N_7327,N_7285);
xor U7416 (N_7416,N_7237,N_7391);
xor U7417 (N_7417,N_7232,N_7386);
nor U7418 (N_7418,N_7309,N_7222);
nor U7419 (N_7419,N_7373,N_7350);
xnor U7420 (N_7420,N_7340,N_7349);
and U7421 (N_7421,N_7253,N_7204);
nand U7422 (N_7422,N_7297,N_7329);
or U7423 (N_7423,N_7214,N_7263);
and U7424 (N_7424,N_7211,N_7276);
and U7425 (N_7425,N_7267,N_7235);
nor U7426 (N_7426,N_7213,N_7254);
or U7427 (N_7427,N_7382,N_7308);
or U7428 (N_7428,N_7264,N_7390);
nor U7429 (N_7429,N_7282,N_7370);
nor U7430 (N_7430,N_7371,N_7226);
and U7431 (N_7431,N_7348,N_7311);
nor U7432 (N_7432,N_7330,N_7272);
xnor U7433 (N_7433,N_7295,N_7333);
or U7434 (N_7434,N_7314,N_7312);
or U7435 (N_7435,N_7274,N_7292);
nor U7436 (N_7436,N_7307,N_7376);
or U7437 (N_7437,N_7302,N_7336);
nand U7438 (N_7438,N_7339,N_7369);
nor U7439 (N_7439,N_7225,N_7286);
nor U7440 (N_7440,N_7310,N_7257);
nor U7441 (N_7441,N_7294,N_7378);
and U7442 (N_7442,N_7236,N_7316);
nor U7443 (N_7443,N_7344,N_7277);
nand U7444 (N_7444,N_7227,N_7249);
or U7445 (N_7445,N_7372,N_7219);
nor U7446 (N_7446,N_7288,N_7298);
or U7447 (N_7447,N_7319,N_7255);
nor U7448 (N_7448,N_7395,N_7328);
nand U7449 (N_7449,N_7355,N_7345);
and U7450 (N_7450,N_7205,N_7363);
nor U7451 (N_7451,N_7359,N_7266);
nand U7452 (N_7452,N_7342,N_7325);
or U7453 (N_7453,N_7293,N_7379);
xor U7454 (N_7454,N_7393,N_7366);
nor U7455 (N_7455,N_7399,N_7241);
nor U7456 (N_7456,N_7384,N_7245);
nor U7457 (N_7457,N_7335,N_7332);
nand U7458 (N_7458,N_7200,N_7221);
nor U7459 (N_7459,N_7396,N_7223);
and U7460 (N_7460,N_7290,N_7270);
or U7461 (N_7461,N_7216,N_7240);
xor U7462 (N_7462,N_7242,N_7231);
nand U7463 (N_7463,N_7278,N_7306);
xnor U7464 (N_7464,N_7217,N_7303);
and U7465 (N_7465,N_7234,N_7351);
xor U7466 (N_7466,N_7320,N_7291);
xnor U7467 (N_7467,N_7244,N_7260);
and U7468 (N_7468,N_7229,N_7367);
nand U7469 (N_7469,N_7388,N_7394);
xor U7470 (N_7470,N_7360,N_7364);
xor U7471 (N_7471,N_7251,N_7279);
and U7472 (N_7472,N_7233,N_7321);
xnor U7473 (N_7473,N_7358,N_7338);
xor U7474 (N_7474,N_7383,N_7228);
xor U7475 (N_7475,N_7215,N_7324);
nor U7476 (N_7476,N_7354,N_7374);
nor U7477 (N_7477,N_7283,N_7398);
nor U7478 (N_7478,N_7304,N_7318);
xnor U7479 (N_7479,N_7334,N_7385);
and U7480 (N_7480,N_7347,N_7284);
or U7481 (N_7481,N_7224,N_7326);
nand U7482 (N_7482,N_7361,N_7252);
nor U7483 (N_7483,N_7201,N_7265);
nor U7484 (N_7484,N_7239,N_7305);
nor U7485 (N_7485,N_7220,N_7317);
xnor U7486 (N_7486,N_7256,N_7357);
nor U7487 (N_7487,N_7218,N_7203);
nand U7488 (N_7488,N_7243,N_7268);
nand U7489 (N_7489,N_7362,N_7206);
or U7490 (N_7490,N_7202,N_7356);
or U7491 (N_7491,N_7246,N_7250);
and U7492 (N_7492,N_7273,N_7331);
and U7493 (N_7493,N_7296,N_7247);
or U7494 (N_7494,N_7337,N_7212);
xor U7495 (N_7495,N_7389,N_7280);
xnor U7496 (N_7496,N_7259,N_7248);
nand U7497 (N_7497,N_7397,N_7262);
xor U7498 (N_7498,N_7301,N_7368);
nand U7499 (N_7499,N_7238,N_7377);
or U7500 (N_7500,N_7205,N_7271);
xor U7501 (N_7501,N_7283,N_7376);
and U7502 (N_7502,N_7281,N_7204);
xnor U7503 (N_7503,N_7280,N_7367);
xor U7504 (N_7504,N_7330,N_7349);
or U7505 (N_7505,N_7306,N_7201);
nor U7506 (N_7506,N_7395,N_7382);
nor U7507 (N_7507,N_7207,N_7355);
and U7508 (N_7508,N_7361,N_7238);
nand U7509 (N_7509,N_7263,N_7291);
nand U7510 (N_7510,N_7322,N_7259);
nand U7511 (N_7511,N_7342,N_7250);
and U7512 (N_7512,N_7234,N_7254);
or U7513 (N_7513,N_7346,N_7353);
nor U7514 (N_7514,N_7334,N_7375);
xor U7515 (N_7515,N_7230,N_7281);
and U7516 (N_7516,N_7324,N_7267);
or U7517 (N_7517,N_7297,N_7203);
nand U7518 (N_7518,N_7331,N_7298);
xnor U7519 (N_7519,N_7384,N_7210);
nor U7520 (N_7520,N_7213,N_7306);
nand U7521 (N_7521,N_7214,N_7371);
nor U7522 (N_7522,N_7381,N_7392);
and U7523 (N_7523,N_7319,N_7242);
or U7524 (N_7524,N_7355,N_7363);
and U7525 (N_7525,N_7324,N_7269);
and U7526 (N_7526,N_7391,N_7229);
xnor U7527 (N_7527,N_7379,N_7333);
nand U7528 (N_7528,N_7355,N_7291);
nand U7529 (N_7529,N_7381,N_7212);
xnor U7530 (N_7530,N_7371,N_7263);
xor U7531 (N_7531,N_7234,N_7248);
xnor U7532 (N_7532,N_7366,N_7362);
or U7533 (N_7533,N_7251,N_7389);
nand U7534 (N_7534,N_7264,N_7319);
nor U7535 (N_7535,N_7344,N_7253);
and U7536 (N_7536,N_7229,N_7216);
xnor U7537 (N_7537,N_7346,N_7367);
and U7538 (N_7538,N_7216,N_7389);
or U7539 (N_7539,N_7354,N_7370);
nand U7540 (N_7540,N_7347,N_7279);
xor U7541 (N_7541,N_7336,N_7291);
or U7542 (N_7542,N_7218,N_7375);
xor U7543 (N_7543,N_7397,N_7242);
nor U7544 (N_7544,N_7385,N_7237);
and U7545 (N_7545,N_7259,N_7218);
nor U7546 (N_7546,N_7332,N_7272);
nand U7547 (N_7547,N_7261,N_7235);
nand U7548 (N_7548,N_7360,N_7298);
nor U7549 (N_7549,N_7212,N_7267);
nor U7550 (N_7550,N_7277,N_7221);
nand U7551 (N_7551,N_7239,N_7235);
nand U7552 (N_7552,N_7356,N_7271);
nor U7553 (N_7553,N_7374,N_7340);
and U7554 (N_7554,N_7266,N_7271);
nor U7555 (N_7555,N_7268,N_7302);
nand U7556 (N_7556,N_7245,N_7315);
nand U7557 (N_7557,N_7237,N_7281);
or U7558 (N_7558,N_7332,N_7239);
nand U7559 (N_7559,N_7365,N_7256);
xnor U7560 (N_7560,N_7328,N_7240);
nor U7561 (N_7561,N_7344,N_7260);
nor U7562 (N_7562,N_7222,N_7349);
nand U7563 (N_7563,N_7390,N_7272);
or U7564 (N_7564,N_7377,N_7211);
or U7565 (N_7565,N_7269,N_7328);
xor U7566 (N_7566,N_7213,N_7203);
nor U7567 (N_7567,N_7231,N_7311);
nor U7568 (N_7568,N_7212,N_7376);
nand U7569 (N_7569,N_7350,N_7244);
or U7570 (N_7570,N_7323,N_7373);
and U7571 (N_7571,N_7248,N_7227);
nand U7572 (N_7572,N_7386,N_7227);
xnor U7573 (N_7573,N_7313,N_7221);
and U7574 (N_7574,N_7227,N_7230);
nand U7575 (N_7575,N_7393,N_7361);
or U7576 (N_7576,N_7337,N_7237);
nor U7577 (N_7577,N_7243,N_7205);
nand U7578 (N_7578,N_7382,N_7231);
nand U7579 (N_7579,N_7256,N_7213);
nand U7580 (N_7580,N_7398,N_7362);
and U7581 (N_7581,N_7389,N_7281);
and U7582 (N_7582,N_7226,N_7225);
nor U7583 (N_7583,N_7214,N_7305);
and U7584 (N_7584,N_7363,N_7310);
or U7585 (N_7585,N_7311,N_7270);
nand U7586 (N_7586,N_7340,N_7222);
nand U7587 (N_7587,N_7223,N_7392);
xor U7588 (N_7588,N_7371,N_7278);
nand U7589 (N_7589,N_7232,N_7205);
xor U7590 (N_7590,N_7333,N_7375);
or U7591 (N_7591,N_7330,N_7295);
nand U7592 (N_7592,N_7329,N_7282);
nor U7593 (N_7593,N_7328,N_7387);
nor U7594 (N_7594,N_7306,N_7328);
xnor U7595 (N_7595,N_7304,N_7373);
nand U7596 (N_7596,N_7229,N_7308);
or U7597 (N_7597,N_7364,N_7399);
nor U7598 (N_7598,N_7224,N_7328);
or U7599 (N_7599,N_7287,N_7387);
xnor U7600 (N_7600,N_7452,N_7492);
nand U7601 (N_7601,N_7483,N_7453);
xnor U7602 (N_7602,N_7523,N_7418);
and U7603 (N_7603,N_7551,N_7474);
xnor U7604 (N_7604,N_7577,N_7574);
and U7605 (N_7605,N_7567,N_7414);
nor U7606 (N_7606,N_7588,N_7438);
and U7607 (N_7607,N_7511,N_7444);
and U7608 (N_7608,N_7466,N_7491);
xnor U7609 (N_7609,N_7400,N_7548);
and U7610 (N_7610,N_7473,N_7500);
and U7611 (N_7611,N_7533,N_7544);
and U7612 (N_7612,N_7572,N_7421);
xnor U7613 (N_7613,N_7516,N_7481);
xnor U7614 (N_7614,N_7527,N_7519);
xor U7615 (N_7615,N_7543,N_7476);
nor U7616 (N_7616,N_7431,N_7554);
xor U7617 (N_7617,N_7568,N_7484);
and U7618 (N_7618,N_7560,N_7424);
and U7619 (N_7619,N_7573,N_7512);
nor U7620 (N_7620,N_7461,N_7417);
xor U7621 (N_7621,N_7435,N_7443);
and U7622 (N_7622,N_7545,N_7487);
nand U7623 (N_7623,N_7427,N_7455);
nand U7624 (N_7624,N_7482,N_7475);
nand U7625 (N_7625,N_7445,N_7426);
xor U7626 (N_7626,N_7490,N_7555);
xnor U7627 (N_7627,N_7441,N_7458);
nor U7628 (N_7628,N_7460,N_7501);
and U7629 (N_7629,N_7580,N_7563);
or U7630 (N_7630,N_7522,N_7409);
and U7631 (N_7631,N_7447,N_7457);
or U7632 (N_7632,N_7589,N_7517);
nand U7633 (N_7633,N_7469,N_7585);
nand U7634 (N_7634,N_7436,N_7597);
xor U7635 (N_7635,N_7599,N_7536);
xnor U7636 (N_7636,N_7525,N_7496);
and U7637 (N_7637,N_7413,N_7472);
and U7638 (N_7638,N_7402,N_7539);
nor U7639 (N_7639,N_7564,N_7468);
xor U7640 (N_7640,N_7583,N_7538);
nand U7641 (N_7641,N_7587,N_7448);
nand U7642 (N_7642,N_7486,N_7579);
nand U7643 (N_7643,N_7419,N_7465);
or U7644 (N_7644,N_7526,N_7510);
nand U7645 (N_7645,N_7578,N_7429);
and U7646 (N_7646,N_7456,N_7464);
and U7647 (N_7647,N_7423,N_7401);
or U7648 (N_7648,N_7590,N_7432);
or U7649 (N_7649,N_7422,N_7557);
or U7650 (N_7650,N_7416,N_7594);
nor U7651 (N_7651,N_7528,N_7477);
xnor U7652 (N_7652,N_7479,N_7504);
nor U7653 (N_7653,N_7521,N_7471);
and U7654 (N_7654,N_7547,N_7485);
and U7655 (N_7655,N_7440,N_7459);
xor U7656 (N_7656,N_7462,N_7507);
xor U7657 (N_7657,N_7550,N_7582);
and U7658 (N_7658,N_7598,N_7463);
nor U7659 (N_7659,N_7561,N_7509);
and U7660 (N_7660,N_7513,N_7530);
nor U7661 (N_7661,N_7532,N_7565);
xnor U7662 (N_7662,N_7451,N_7531);
and U7663 (N_7663,N_7407,N_7470);
and U7664 (N_7664,N_7576,N_7595);
or U7665 (N_7665,N_7450,N_7406);
or U7666 (N_7666,N_7570,N_7446);
nand U7667 (N_7667,N_7425,N_7562);
and U7668 (N_7668,N_7495,N_7437);
and U7669 (N_7669,N_7442,N_7434);
and U7670 (N_7670,N_7410,N_7494);
and U7671 (N_7671,N_7404,N_7535);
or U7672 (N_7672,N_7596,N_7489);
or U7673 (N_7673,N_7415,N_7581);
nor U7674 (N_7674,N_7439,N_7454);
xor U7675 (N_7675,N_7488,N_7499);
and U7676 (N_7676,N_7575,N_7433);
nand U7677 (N_7677,N_7497,N_7503);
xnor U7678 (N_7678,N_7549,N_7514);
xnor U7679 (N_7679,N_7558,N_7569);
xor U7680 (N_7680,N_7518,N_7559);
xnor U7681 (N_7681,N_7498,N_7546);
and U7682 (N_7682,N_7540,N_7430);
nand U7683 (N_7683,N_7542,N_7480);
and U7684 (N_7684,N_7524,N_7553);
xnor U7685 (N_7685,N_7571,N_7403);
nand U7686 (N_7686,N_7541,N_7449);
xor U7687 (N_7687,N_7534,N_7515);
or U7688 (N_7688,N_7467,N_7506);
xnor U7689 (N_7689,N_7493,N_7502);
or U7690 (N_7690,N_7537,N_7584);
nand U7691 (N_7691,N_7592,N_7508);
xor U7692 (N_7692,N_7505,N_7420);
xnor U7693 (N_7693,N_7586,N_7556);
or U7694 (N_7694,N_7552,N_7408);
or U7695 (N_7695,N_7529,N_7591);
nor U7696 (N_7696,N_7428,N_7405);
or U7697 (N_7697,N_7593,N_7478);
and U7698 (N_7698,N_7412,N_7520);
and U7699 (N_7699,N_7411,N_7566);
nor U7700 (N_7700,N_7442,N_7533);
xor U7701 (N_7701,N_7527,N_7447);
nor U7702 (N_7702,N_7561,N_7554);
or U7703 (N_7703,N_7432,N_7573);
nor U7704 (N_7704,N_7522,N_7405);
xor U7705 (N_7705,N_7557,N_7584);
xor U7706 (N_7706,N_7560,N_7432);
nand U7707 (N_7707,N_7436,N_7485);
nor U7708 (N_7708,N_7417,N_7561);
nor U7709 (N_7709,N_7527,N_7481);
nor U7710 (N_7710,N_7420,N_7448);
or U7711 (N_7711,N_7406,N_7487);
xor U7712 (N_7712,N_7407,N_7490);
xnor U7713 (N_7713,N_7515,N_7425);
nor U7714 (N_7714,N_7584,N_7411);
nand U7715 (N_7715,N_7425,N_7506);
xnor U7716 (N_7716,N_7414,N_7504);
xor U7717 (N_7717,N_7489,N_7550);
nor U7718 (N_7718,N_7588,N_7506);
and U7719 (N_7719,N_7468,N_7512);
nor U7720 (N_7720,N_7559,N_7423);
nand U7721 (N_7721,N_7422,N_7532);
nor U7722 (N_7722,N_7505,N_7452);
nor U7723 (N_7723,N_7547,N_7534);
or U7724 (N_7724,N_7450,N_7483);
nor U7725 (N_7725,N_7476,N_7584);
xor U7726 (N_7726,N_7530,N_7522);
and U7727 (N_7727,N_7504,N_7526);
nand U7728 (N_7728,N_7547,N_7430);
nor U7729 (N_7729,N_7443,N_7535);
nand U7730 (N_7730,N_7436,N_7554);
xor U7731 (N_7731,N_7579,N_7447);
xnor U7732 (N_7732,N_7591,N_7436);
and U7733 (N_7733,N_7413,N_7533);
nand U7734 (N_7734,N_7422,N_7590);
nor U7735 (N_7735,N_7436,N_7475);
xor U7736 (N_7736,N_7404,N_7505);
nand U7737 (N_7737,N_7516,N_7454);
or U7738 (N_7738,N_7453,N_7449);
nor U7739 (N_7739,N_7528,N_7422);
and U7740 (N_7740,N_7549,N_7554);
nand U7741 (N_7741,N_7470,N_7587);
or U7742 (N_7742,N_7580,N_7401);
xor U7743 (N_7743,N_7445,N_7583);
xnor U7744 (N_7744,N_7575,N_7545);
nor U7745 (N_7745,N_7592,N_7578);
nor U7746 (N_7746,N_7551,N_7446);
xnor U7747 (N_7747,N_7435,N_7476);
xnor U7748 (N_7748,N_7564,N_7471);
nor U7749 (N_7749,N_7418,N_7405);
and U7750 (N_7750,N_7583,N_7423);
or U7751 (N_7751,N_7481,N_7559);
nand U7752 (N_7752,N_7439,N_7539);
and U7753 (N_7753,N_7464,N_7453);
nor U7754 (N_7754,N_7584,N_7409);
xor U7755 (N_7755,N_7510,N_7527);
or U7756 (N_7756,N_7414,N_7419);
xor U7757 (N_7757,N_7588,N_7490);
or U7758 (N_7758,N_7519,N_7409);
or U7759 (N_7759,N_7477,N_7479);
xnor U7760 (N_7760,N_7402,N_7449);
xnor U7761 (N_7761,N_7473,N_7594);
nor U7762 (N_7762,N_7588,N_7453);
or U7763 (N_7763,N_7421,N_7569);
or U7764 (N_7764,N_7541,N_7482);
nor U7765 (N_7765,N_7519,N_7400);
and U7766 (N_7766,N_7489,N_7587);
xnor U7767 (N_7767,N_7438,N_7465);
or U7768 (N_7768,N_7536,N_7504);
or U7769 (N_7769,N_7462,N_7405);
and U7770 (N_7770,N_7590,N_7529);
nor U7771 (N_7771,N_7593,N_7442);
or U7772 (N_7772,N_7406,N_7529);
xor U7773 (N_7773,N_7595,N_7563);
and U7774 (N_7774,N_7587,N_7530);
or U7775 (N_7775,N_7570,N_7552);
and U7776 (N_7776,N_7468,N_7529);
nand U7777 (N_7777,N_7548,N_7599);
or U7778 (N_7778,N_7441,N_7509);
xor U7779 (N_7779,N_7448,N_7476);
nor U7780 (N_7780,N_7422,N_7594);
and U7781 (N_7781,N_7509,N_7485);
and U7782 (N_7782,N_7464,N_7587);
and U7783 (N_7783,N_7577,N_7465);
and U7784 (N_7784,N_7523,N_7424);
xnor U7785 (N_7785,N_7559,N_7420);
nand U7786 (N_7786,N_7433,N_7441);
xor U7787 (N_7787,N_7537,N_7576);
and U7788 (N_7788,N_7561,N_7588);
xnor U7789 (N_7789,N_7434,N_7531);
and U7790 (N_7790,N_7456,N_7459);
nor U7791 (N_7791,N_7478,N_7587);
xor U7792 (N_7792,N_7504,N_7506);
xor U7793 (N_7793,N_7413,N_7495);
nor U7794 (N_7794,N_7468,N_7590);
and U7795 (N_7795,N_7581,N_7450);
xor U7796 (N_7796,N_7575,N_7597);
nand U7797 (N_7797,N_7484,N_7574);
and U7798 (N_7798,N_7510,N_7568);
and U7799 (N_7799,N_7513,N_7415);
xor U7800 (N_7800,N_7669,N_7769);
xor U7801 (N_7801,N_7699,N_7690);
nand U7802 (N_7802,N_7675,N_7752);
and U7803 (N_7803,N_7634,N_7641);
nor U7804 (N_7804,N_7784,N_7651);
or U7805 (N_7805,N_7781,N_7731);
xnor U7806 (N_7806,N_7629,N_7631);
xor U7807 (N_7807,N_7665,N_7645);
nor U7808 (N_7808,N_7745,N_7661);
or U7809 (N_7809,N_7799,N_7642);
xor U7810 (N_7810,N_7736,N_7617);
nand U7811 (N_7811,N_7622,N_7720);
and U7812 (N_7812,N_7635,N_7709);
nor U7813 (N_7813,N_7742,N_7630);
xnor U7814 (N_7814,N_7793,N_7671);
nor U7815 (N_7815,N_7673,N_7640);
xnor U7816 (N_7816,N_7703,N_7654);
and U7817 (N_7817,N_7646,N_7653);
xor U7818 (N_7818,N_7691,N_7750);
or U7819 (N_7819,N_7636,N_7607);
xnor U7820 (N_7820,N_7765,N_7763);
and U7821 (N_7821,N_7624,N_7776);
and U7822 (N_7822,N_7606,N_7710);
or U7823 (N_7823,N_7743,N_7678);
or U7824 (N_7824,N_7663,N_7701);
nor U7825 (N_7825,N_7726,N_7647);
nor U7826 (N_7826,N_7615,N_7774);
nand U7827 (N_7827,N_7733,N_7603);
xnor U7828 (N_7828,N_7626,N_7608);
nor U7829 (N_7829,N_7753,N_7785);
xor U7830 (N_7830,N_7715,N_7760);
nor U7831 (N_7831,N_7604,N_7689);
or U7832 (N_7832,N_7755,N_7790);
and U7833 (N_7833,N_7712,N_7702);
or U7834 (N_7834,N_7734,N_7660);
nor U7835 (N_7835,N_7637,N_7724);
or U7836 (N_7836,N_7766,N_7789);
or U7837 (N_7837,N_7794,N_7714);
nor U7838 (N_7838,N_7609,N_7782);
and U7839 (N_7839,N_7713,N_7666);
nor U7840 (N_7840,N_7659,N_7718);
nor U7841 (N_7841,N_7758,N_7674);
nor U7842 (N_7842,N_7686,N_7610);
nand U7843 (N_7843,N_7795,N_7627);
xnor U7844 (N_7844,N_7680,N_7762);
xor U7845 (N_7845,N_7600,N_7735);
nand U7846 (N_7846,N_7677,N_7652);
nor U7847 (N_7847,N_7768,N_7706);
nor U7848 (N_7848,N_7728,N_7643);
xor U7849 (N_7849,N_7664,N_7614);
xor U7850 (N_7850,N_7616,N_7620);
xnor U7851 (N_7851,N_7773,N_7628);
xor U7852 (N_7852,N_7685,N_7775);
nor U7853 (N_7853,N_7757,N_7751);
or U7854 (N_7854,N_7679,N_7612);
nor U7855 (N_7855,N_7700,N_7696);
xor U7856 (N_7856,N_7780,N_7602);
or U7857 (N_7857,N_7681,N_7698);
or U7858 (N_7858,N_7633,N_7601);
nand U7859 (N_7859,N_7730,N_7704);
xor U7860 (N_7860,N_7725,N_7740);
xor U7861 (N_7861,N_7632,N_7759);
xnor U7862 (N_7862,N_7747,N_7741);
nor U7863 (N_7863,N_7694,N_7721);
and U7864 (N_7864,N_7738,N_7746);
xor U7865 (N_7865,N_7771,N_7798);
and U7866 (N_7866,N_7623,N_7707);
and U7867 (N_7867,N_7796,N_7711);
or U7868 (N_7868,N_7717,N_7770);
nor U7869 (N_7869,N_7772,N_7658);
nand U7870 (N_7870,N_7719,N_7619);
nor U7871 (N_7871,N_7697,N_7670);
and U7872 (N_7872,N_7687,N_7754);
nor U7873 (N_7873,N_7749,N_7656);
xnor U7874 (N_7874,N_7767,N_7723);
and U7875 (N_7875,N_7621,N_7737);
nor U7876 (N_7876,N_7639,N_7748);
nor U7877 (N_7877,N_7618,N_7787);
or U7878 (N_7878,N_7613,N_7682);
nor U7879 (N_7879,N_7777,N_7744);
nor U7880 (N_7880,N_7655,N_7792);
nand U7881 (N_7881,N_7708,N_7722);
or U7882 (N_7882,N_7644,N_7791);
xnor U7883 (N_7883,N_7657,N_7739);
nor U7884 (N_7884,N_7778,N_7625);
xnor U7885 (N_7885,N_7684,N_7732);
nand U7886 (N_7886,N_7638,N_7756);
or U7887 (N_7887,N_7783,N_7662);
or U7888 (N_7888,N_7695,N_7667);
nor U7889 (N_7889,N_7705,N_7716);
nor U7890 (N_7890,N_7764,N_7761);
xnor U7891 (N_7891,N_7683,N_7692);
nand U7892 (N_7892,N_7788,N_7605);
or U7893 (N_7893,N_7688,N_7649);
nor U7894 (N_7894,N_7729,N_7797);
and U7895 (N_7895,N_7648,N_7676);
nor U7896 (N_7896,N_7668,N_7779);
and U7897 (N_7897,N_7611,N_7786);
xnor U7898 (N_7898,N_7693,N_7672);
nor U7899 (N_7899,N_7650,N_7727);
nand U7900 (N_7900,N_7789,N_7673);
and U7901 (N_7901,N_7726,N_7633);
xor U7902 (N_7902,N_7767,N_7661);
nand U7903 (N_7903,N_7782,N_7769);
nand U7904 (N_7904,N_7628,N_7734);
and U7905 (N_7905,N_7665,N_7674);
xor U7906 (N_7906,N_7687,N_7645);
and U7907 (N_7907,N_7686,N_7760);
nand U7908 (N_7908,N_7733,N_7756);
and U7909 (N_7909,N_7620,N_7767);
nand U7910 (N_7910,N_7685,N_7713);
nand U7911 (N_7911,N_7692,N_7600);
and U7912 (N_7912,N_7794,N_7668);
nor U7913 (N_7913,N_7788,N_7677);
or U7914 (N_7914,N_7744,N_7698);
or U7915 (N_7915,N_7685,N_7601);
xor U7916 (N_7916,N_7624,N_7643);
xor U7917 (N_7917,N_7774,N_7689);
xnor U7918 (N_7918,N_7631,N_7608);
or U7919 (N_7919,N_7723,N_7638);
nand U7920 (N_7920,N_7644,N_7694);
xnor U7921 (N_7921,N_7657,N_7702);
and U7922 (N_7922,N_7683,N_7656);
or U7923 (N_7923,N_7667,N_7645);
xnor U7924 (N_7924,N_7795,N_7744);
nand U7925 (N_7925,N_7640,N_7705);
nor U7926 (N_7926,N_7784,N_7654);
and U7927 (N_7927,N_7644,N_7781);
nand U7928 (N_7928,N_7708,N_7786);
and U7929 (N_7929,N_7749,N_7675);
and U7930 (N_7930,N_7717,N_7704);
and U7931 (N_7931,N_7625,N_7796);
and U7932 (N_7932,N_7780,N_7693);
or U7933 (N_7933,N_7739,N_7694);
xor U7934 (N_7934,N_7676,N_7755);
xor U7935 (N_7935,N_7650,N_7732);
nor U7936 (N_7936,N_7610,N_7756);
xnor U7937 (N_7937,N_7669,N_7697);
nor U7938 (N_7938,N_7686,N_7728);
and U7939 (N_7939,N_7620,N_7758);
and U7940 (N_7940,N_7739,N_7637);
nand U7941 (N_7941,N_7693,N_7759);
nor U7942 (N_7942,N_7627,N_7726);
or U7943 (N_7943,N_7648,N_7633);
nand U7944 (N_7944,N_7663,N_7630);
nand U7945 (N_7945,N_7621,N_7660);
nor U7946 (N_7946,N_7710,N_7718);
and U7947 (N_7947,N_7724,N_7615);
nand U7948 (N_7948,N_7705,N_7699);
and U7949 (N_7949,N_7774,N_7621);
xor U7950 (N_7950,N_7705,N_7780);
nor U7951 (N_7951,N_7601,N_7651);
nor U7952 (N_7952,N_7739,N_7667);
nor U7953 (N_7953,N_7681,N_7683);
nor U7954 (N_7954,N_7714,N_7708);
nand U7955 (N_7955,N_7748,N_7672);
nor U7956 (N_7956,N_7618,N_7780);
xnor U7957 (N_7957,N_7760,N_7662);
and U7958 (N_7958,N_7760,N_7601);
xnor U7959 (N_7959,N_7604,N_7750);
nor U7960 (N_7960,N_7681,N_7669);
nand U7961 (N_7961,N_7797,N_7785);
or U7962 (N_7962,N_7668,N_7762);
nand U7963 (N_7963,N_7714,N_7726);
nand U7964 (N_7964,N_7651,N_7782);
nor U7965 (N_7965,N_7714,N_7680);
nand U7966 (N_7966,N_7625,N_7708);
nor U7967 (N_7967,N_7697,N_7663);
and U7968 (N_7968,N_7655,N_7766);
or U7969 (N_7969,N_7734,N_7608);
nor U7970 (N_7970,N_7724,N_7667);
xor U7971 (N_7971,N_7607,N_7792);
and U7972 (N_7972,N_7730,N_7619);
or U7973 (N_7973,N_7717,N_7675);
and U7974 (N_7974,N_7746,N_7719);
xor U7975 (N_7975,N_7681,N_7790);
or U7976 (N_7976,N_7755,N_7668);
or U7977 (N_7977,N_7680,N_7756);
or U7978 (N_7978,N_7793,N_7667);
nor U7979 (N_7979,N_7719,N_7791);
nand U7980 (N_7980,N_7719,N_7724);
and U7981 (N_7981,N_7662,N_7665);
and U7982 (N_7982,N_7784,N_7680);
or U7983 (N_7983,N_7649,N_7643);
nand U7984 (N_7984,N_7698,N_7779);
or U7985 (N_7985,N_7755,N_7694);
and U7986 (N_7986,N_7693,N_7652);
nor U7987 (N_7987,N_7652,N_7699);
nor U7988 (N_7988,N_7763,N_7625);
xor U7989 (N_7989,N_7761,N_7614);
xor U7990 (N_7990,N_7658,N_7741);
or U7991 (N_7991,N_7758,N_7628);
xor U7992 (N_7992,N_7747,N_7736);
xnor U7993 (N_7993,N_7631,N_7733);
nand U7994 (N_7994,N_7676,N_7643);
nor U7995 (N_7995,N_7704,N_7783);
nand U7996 (N_7996,N_7658,N_7639);
or U7997 (N_7997,N_7637,N_7750);
or U7998 (N_7998,N_7640,N_7679);
nand U7999 (N_7999,N_7673,N_7647);
nor U8000 (N_8000,N_7835,N_7922);
nand U8001 (N_8001,N_7936,N_7844);
nand U8002 (N_8002,N_7809,N_7807);
or U8003 (N_8003,N_7894,N_7893);
nor U8004 (N_8004,N_7943,N_7965);
or U8005 (N_8005,N_7947,N_7886);
xnor U8006 (N_8006,N_7828,N_7854);
and U8007 (N_8007,N_7957,N_7982);
nor U8008 (N_8008,N_7910,N_7892);
and U8009 (N_8009,N_7932,N_7956);
or U8010 (N_8010,N_7913,N_7950);
nor U8011 (N_8011,N_7816,N_7827);
or U8012 (N_8012,N_7852,N_7900);
and U8013 (N_8013,N_7916,N_7838);
or U8014 (N_8014,N_7963,N_7880);
nand U8015 (N_8015,N_7981,N_7918);
nand U8016 (N_8016,N_7866,N_7818);
nand U8017 (N_8017,N_7912,N_7977);
nor U8018 (N_8018,N_7917,N_7871);
nor U8019 (N_8019,N_7858,N_7948);
xor U8020 (N_8020,N_7878,N_7914);
nand U8021 (N_8021,N_7840,N_7968);
xnor U8022 (N_8022,N_7883,N_7890);
nor U8023 (N_8023,N_7806,N_7974);
or U8024 (N_8024,N_7868,N_7902);
xnor U8025 (N_8025,N_7908,N_7915);
nor U8026 (N_8026,N_7990,N_7966);
and U8027 (N_8027,N_7933,N_7837);
and U8028 (N_8028,N_7939,N_7879);
nor U8029 (N_8029,N_7951,N_7821);
nor U8030 (N_8030,N_7802,N_7920);
nand U8031 (N_8031,N_7823,N_7889);
and U8032 (N_8032,N_7847,N_7833);
or U8033 (N_8033,N_7994,N_7831);
and U8034 (N_8034,N_7969,N_7953);
nor U8035 (N_8035,N_7906,N_7986);
or U8036 (N_8036,N_7876,N_7848);
or U8037 (N_8037,N_7928,N_7949);
and U8038 (N_8038,N_7870,N_7984);
nor U8039 (N_8039,N_7874,N_7832);
and U8040 (N_8040,N_7921,N_7972);
or U8041 (N_8041,N_7891,N_7971);
xor U8042 (N_8042,N_7896,N_7810);
or U8043 (N_8043,N_7851,N_7803);
nand U8044 (N_8044,N_7997,N_7938);
and U8045 (N_8045,N_7985,N_7903);
or U8046 (N_8046,N_7826,N_7814);
and U8047 (N_8047,N_7907,N_7877);
nand U8048 (N_8048,N_7875,N_7905);
nor U8049 (N_8049,N_7887,N_7813);
nor U8050 (N_8050,N_7993,N_7929);
nand U8051 (N_8051,N_7960,N_7859);
nand U8052 (N_8052,N_7869,N_7873);
nand U8053 (N_8053,N_7857,N_7976);
nand U8054 (N_8054,N_7961,N_7849);
and U8055 (N_8055,N_7995,N_7925);
xor U8056 (N_8056,N_7808,N_7860);
xor U8057 (N_8057,N_7867,N_7935);
and U8058 (N_8058,N_7952,N_7946);
nor U8059 (N_8059,N_7964,N_7805);
nand U8060 (N_8060,N_7884,N_7864);
nand U8061 (N_8061,N_7830,N_7872);
and U8062 (N_8062,N_7979,N_7861);
nor U8063 (N_8063,N_7944,N_7958);
and U8064 (N_8064,N_7845,N_7801);
nor U8065 (N_8065,N_7962,N_7853);
nand U8066 (N_8066,N_7811,N_7911);
and U8067 (N_8067,N_7897,N_7834);
nand U8068 (N_8068,N_7885,N_7898);
and U8069 (N_8069,N_7980,N_7927);
xor U8070 (N_8070,N_7800,N_7988);
or U8071 (N_8071,N_7919,N_7846);
nor U8072 (N_8072,N_7973,N_7959);
nand U8073 (N_8073,N_7954,N_7978);
nor U8074 (N_8074,N_7862,N_7940);
nor U8075 (N_8075,N_7999,N_7817);
nand U8076 (N_8076,N_7812,N_7839);
or U8077 (N_8077,N_7895,N_7829);
nor U8078 (N_8078,N_7942,N_7924);
nand U8079 (N_8079,N_7820,N_7882);
and U8080 (N_8080,N_7987,N_7926);
nor U8081 (N_8081,N_7819,N_7855);
xor U8082 (N_8082,N_7991,N_7930);
or U8083 (N_8083,N_7881,N_7804);
or U8084 (N_8084,N_7989,N_7909);
or U8085 (N_8085,N_7822,N_7975);
nor U8086 (N_8086,N_7983,N_7923);
and U8087 (N_8087,N_7941,N_7931);
xor U8088 (N_8088,N_7825,N_7934);
nand U8089 (N_8089,N_7901,N_7996);
xnor U8090 (N_8090,N_7937,N_7945);
or U8091 (N_8091,N_7850,N_7970);
or U8092 (N_8092,N_7955,N_7836);
or U8093 (N_8093,N_7815,N_7865);
xor U8094 (N_8094,N_7863,N_7841);
and U8095 (N_8095,N_7856,N_7998);
nor U8096 (N_8096,N_7967,N_7904);
xor U8097 (N_8097,N_7824,N_7843);
nand U8098 (N_8098,N_7842,N_7899);
nor U8099 (N_8099,N_7888,N_7992);
nand U8100 (N_8100,N_7903,N_7999);
nor U8101 (N_8101,N_7966,N_7803);
and U8102 (N_8102,N_7927,N_7990);
nor U8103 (N_8103,N_7970,N_7816);
xor U8104 (N_8104,N_7943,N_7823);
or U8105 (N_8105,N_7925,N_7983);
and U8106 (N_8106,N_7876,N_7952);
and U8107 (N_8107,N_7835,N_7825);
or U8108 (N_8108,N_7923,N_7971);
xnor U8109 (N_8109,N_7875,N_7988);
and U8110 (N_8110,N_7911,N_7845);
or U8111 (N_8111,N_7840,N_7909);
nor U8112 (N_8112,N_7859,N_7928);
or U8113 (N_8113,N_7964,N_7947);
and U8114 (N_8114,N_7805,N_7892);
nor U8115 (N_8115,N_7933,N_7897);
xnor U8116 (N_8116,N_7938,N_7975);
or U8117 (N_8117,N_7852,N_7813);
nand U8118 (N_8118,N_7990,N_7941);
xor U8119 (N_8119,N_7930,N_7824);
nor U8120 (N_8120,N_7822,N_7876);
and U8121 (N_8121,N_7990,N_7893);
and U8122 (N_8122,N_7814,N_7842);
or U8123 (N_8123,N_7924,N_7982);
or U8124 (N_8124,N_7813,N_7871);
or U8125 (N_8125,N_7804,N_7859);
nor U8126 (N_8126,N_7913,N_7874);
xnor U8127 (N_8127,N_7860,N_7914);
xor U8128 (N_8128,N_7977,N_7803);
nor U8129 (N_8129,N_7962,N_7808);
nand U8130 (N_8130,N_7807,N_7915);
or U8131 (N_8131,N_7803,N_7937);
or U8132 (N_8132,N_7940,N_7939);
or U8133 (N_8133,N_7930,N_7967);
and U8134 (N_8134,N_7913,N_7864);
nand U8135 (N_8135,N_7826,N_7978);
nor U8136 (N_8136,N_7878,N_7815);
nor U8137 (N_8137,N_7923,N_7991);
nor U8138 (N_8138,N_7964,N_7905);
or U8139 (N_8139,N_7909,N_7823);
nor U8140 (N_8140,N_7803,N_7945);
and U8141 (N_8141,N_7995,N_7861);
or U8142 (N_8142,N_7928,N_7852);
xor U8143 (N_8143,N_7824,N_7886);
or U8144 (N_8144,N_7939,N_7846);
nand U8145 (N_8145,N_7985,N_7846);
or U8146 (N_8146,N_7949,N_7802);
nor U8147 (N_8147,N_7913,N_7988);
nor U8148 (N_8148,N_7814,N_7866);
nand U8149 (N_8149,N_7986,N_7952);
xnor U8150 (N_8150,N_7999,N_7875);
nor U8151 (N_8151,N_7892,N_7963);
or U8152 (N_8152,N_7820,N_7992);
nor U8153 (N_8153,N_7825,N_7838);
xnor U8154 (N_8154,N_7815,N_7841);
xnor U8155 (N_8155,N_7819,N_7832);
or U8156 (N_8156,N_7995,N_7951);
nor U8157 (N_8157,N_7944,N_7930);
and U8158 (N_8158,N_7844,N_7836);
xor U8159 (N_8159,N_7979,N_7899);
nand U8160 (N_8160,N_7851,N_7975);
and U8161 (N_8161,N_7837,N_7842);
nand U8162 (N_8162,N_7930,N_7862);
and U8163 (N_8163,N_7886,N_7975);
nand U8164 (N_8164,N_7937,N_7864);
or U8165 (N_8165,N_7996,N_7812);
nand U8166 (N_8166,N_7989,N_7947);
or U8167 (N_8167,N_7898,N_7820);
nand U8168 (N_8168,N_7996,N_7914);
or U8169 (N_8169,N_7868,N_7828);
nand U8170 (N_8170,N_7973,N_7902);
nand U8171 (N_8171,N_7819,N_7956);
and U8172 (N_8172,N_7950,N_7876);
xnor U8173 (N_8173,N_7829,N_7980);
nor U8174 (N_8174,N_7855,N_7875);
and U8175 (N_8175,N_7903,N_7963);
and U8176 (N_8176,N_7955,N_7943);
and U8177 (N_8177,N_7943,N_7803);
nor U8178 (N_8178,N_7930,N_7804);
xnor U8179 (N_8179,N_7938,N_7821);
or U8180 (N_8180,N_7875,N_7921);
and U8181 (N_8181,N_7902,N_7965);
nand U8182 (N_8182,N_7808,N_7964);
or U8183 (N_8183,N_7815,N_7885);
or U8184 (N_8184,N_7947,N_7978);
xor U8185 (N_8185,N_7861,N_7905);
nand U8186 (N_8186,N_7836,N_7866);
and U8187 (N_8187,N_7976,N_7841);
nand U8188 (N_8188,N_7845,N_7841);
nand U8189 (N_8189,N_7951,N_7987);
nand U8190 (N_8190,N_7874,N_7894);
and U8191 (N_8191,N_7980,N_7917);
nand U8192 (N_8192,N_7853,N_7928);
xor U8193 (N_8193,N_7831,N_7987);
and U8194 (N_8194,N_7941,N_7812);
nand U8195 (N_8195,N_7989,N_7889);
or U8196 (N_8196,N_7976,N_7991);
xor U8197 (N_8197,N_7931,N_7899);
nor U8198 (N_8198,N_7907,N_7930);
nand U8199 (N_8199,N_7824,N_7862);
or U8200 (N_8200,N_8017,N_8125);
and U8201 (N_8201,N_8123,N_8075);
or U8202 (N_8202,N_8196,N_8081);
or U8203 (N_8203,N_8035,N_8004);
or U8204 (N_8204,N_8107,N_8157);
nand U8205 (N_8205,N_8134,N_8188);
xor U8206 (N_8206,N_8176,N_8066);
nor U8207 (N_8207,N_8161,N_8088);
and U8208 (N_8208,N_8077,N_8085);
xor U8209 (N_8209,N_8136,N_8140);
xor U8210 (N_8210,N_8187,N_8053);
xnor U8211 (N_8211,N_8034,N_8014);
xnor U8212 (N_8212,N_8122,N_8104);
or U8213 (N_8213,N_8058,N_8128);
and U8214 (N_8214,N_8048,N_8180);
xnor U8215 (N_8215,N_8001,N_8159);
or U8216 (N_8216,N_8111,N_8160);
xor U8217 (N_8217,N_8072,N_8163);
xnor U8218 (N_8218,N_8026,N_8002);
or U8219 (N_8219,N_8194,N_8198);
xor U8220 (N_8220,N_8091,N_8158);
xor U8221 (N_8221,N_8031,N_8155);
or U8222 (N_8222,N_8129,N_8065);
and U8223 (N_8223,N_8106,N_8010);
and U8224 (N_8224,N_8033,N_8191);
nor U8225 (N_8225,N_8108,N_8015);
or U8226 (N_8226,N_8118,N_8131);
and U8227 (N_8227,N_8071,N_8126);
xnor U8228 (N_8228,N_8069,N_8102);
nor U8229 (N_8229,N_8051,N_8199);
nand U8230 (N_8230,N_8164,N_8184);
and U8231 (N_8231,N_8092,N_8132);
xnor U8232 (N_8232,N_8074,N_8055);
or U8233 (N_8233,N_8142,N_8008);
nor U8234 (N_8234,N_8078,N_8062);
nor U8235 (N_8235,N_8024,N_8137);
or U8236 (N_8236,N_8165,N_8090);
nor U8237 (N_8237,N_8154,N_8022);
nand U8238 (N_8238,N_8143,N_8027);
or U8239 (N_8239,N_8120,N_8037);
and U8240 (N_8240,N_8113,N_8135);
nor U8241 (N_8241,N_8086,N_8080);
xnor U8242 (N_8242,N_8149,N_8192);
nor U8243 (N_8243,N_8119,N_8012);
nor U8244 (N_8244,N_8049,N_8133);
nand U8245 (N_8245,N_8045,N_8067);
nor U8246 (N_8246,N_8029,N_8038);
or U8247 (N_8247,N_8181,N_8153);
xor U8248 (N_8248,N_8173,N_8032);
nor U8249 (N_8249,N_8121,N_8050);
nor U8250 (N_8250,N_8046,N_8185);
and U8251 (N_8251,N_8167,N_8193);
nor U8252 (N_8252,N_8079,N_8094);
nand U8253 (N_8253,N_8190,N_8098);
nand U8254 (N_8254,N_8114,N_8101);
xor U8255 (N_8255,N_8082,N_8087);
or U8256 (N_8256,N_8171,N_8068);
xor U8257 (N_8257,N_8182,N_8179);
and U8258 (N_8258,N_8039,N_8020);
nor U8259 (N_8259,N_8152,N_8097);
nor U8260 (N_8260,N_8197,N_8059);
xnor U8261 (N_8261,N_8052,N_8150);
xnor U8262 (N_8262,N_8073,N_8186);
or U8263 (N_8263,N_8195,N_8041);
and U8264 (N_8264,N_8175,N_8007);
and U8265 (N_8265,N_8021,N_8183);
nor U8266 (N_8266,N_8138,N_8060);
nor U8267 (N_8267,N_8044,N_8156);
nand U8268 (N_8268,N_8043,N_8109);
nand U8269 (N_8269,N_8141,N_8169);
xor U8270 (N_8270,N_8124,N_8168);
and U8271 (N_8271,N_8189,N_8009);
nor U8272 (N_8272,N_8095,N_8030);
or U8273 (N_8273,N_8145,N_8130);
nand U8274 (N_8274,N_8025,N_8047);
or U8275 (N_8275,N_8076,N_8054);
nand U8276 (N_8276,N_8070,N_8110);
and U8277 (N_8277,N_8170,N_8172);
nor U8278 (N_8278,N_8013,N_8042);
and U8279 (N_8279,N_8064,N_8174);
and U8280 (N_8280,N_8083,N_8117);
or U8281 (N_8281,N_8127,N_8018);
xor U8282 (N_8282,N_8016,N_8139);
and U8283 (N_8283,N_8177,N_8112);
nor U8284 (N_8284,N_8144,N_8178);
and U8285 (N_8285,N_8096,N_8148);
nor U8286 (N_8286,N_8011,N_8061);
nor U8287 (N_8287,N_8162,N_8146);
xnor U8288 (N_8288,N_8093,N_8105);
xnor U8289 (N_8289,N_8040,N_8057);
nand U8290 (N_8290,N_8056,N_8019);
or U8291 (N_8291,N_8006,N_8151);
and U8292 (N_8292,N_8003,N_8115);
nand U8293 (N_8293,N_8116,N_8028);
and U8294 (N_8294,N_8023,N_8063);
and U8295 (N_8295,N_8036,N_8166);
nand U8296 (N_8296,N_8099,N_8103);
or U8297 (N_8297,N_8005,N_8147);
nor U8298 (N_8298,N_8084,N_8089);
xnor U8299 (N_8299,N_8000,N_8100);
or U8300 (N_8300,N_8009,N_8071);
xor U8301 (N_8301,N_8161,N_8042);
xor U8302 (N_8302,N_8070,N_8111);
nor U8303 (N_8303,N_8186,N_8066);
nor U8304 (N_8304,N_8130,N_8027);
and U8305 (N_8305,N_8160,N_8179);
nor U8306 (N_8306,N_8180,N_8095);
xnor U8307 (N_8307,N_8100,N_8141);
and U8308 (N_8308,N_8045,N_8129);
and U8309 (N_8309,N_8111,N_8028);
nor U8310 (N_8310,N_8078,N_8091);
or U8311 (N_8311,N_8088,N_8092);
and U8312 (N_8312,N_8164,N_8053);
nor U8313 (N_8313,N_8156,N_8102);
and U8314 (N_8314,N_8013,N_8104);
nor U8315 (N_8315,N_8090,N_8053);
nand U8316 (N_8316,N_8130,N_8046);
nor U8317 (N_8317,N_8140,N_8160);
and U8318 (N_8318,N_8095,N_8129);
xnor U8319 (N_8319,N_8110,N_8030);
nor U8320 (N_8320,N_8105,N_8097);
nand U8321 (N_8321,N_8051,N_8107);
xnor U8322 (N_8322,N_8090,N_8196);
nor U8323 (N_8323,N_8127,N_8133);
xor U8324 (N_8324,N_8144,N_8039);
or U8325 (N_8325,N_8010,N_8030);
nor U8326 (N_8326,N_8071,N_8198);
and U8327 (N_8327,N_8114,N_8123);
nor U8328 (N_8328,N_8172,N_8114);
or U8329 (N_8329,N_8183,N_8072);
or U8330 (N_8330,N_8076,N_8185);
or U8331 (N_8331,N_8173,N_8170);
nand U8332 (N_8332,N_8156,N_8035);
nor U8333 (N_8333,N_8084,N_8146);
nand U8334 (N_8334,N_8076,N_8178);
nand U8335 (N_8335,N_8153,N_8169);
nand U8336 (N_8336,N_8145,N_8044);
xor U8337 (N_8337,N_8196,N_8114);
xor U8338 (N_8338,N_8110,N_8123);
nand U8339 (N_8339,N_8019,N_8196);
xnor U8340 (N_8340,N_8190,N_8151);
nand U8341 (N_8341,N_8190,N_8122);
nand U8342 (N_8342,N_8013,N_8037);
nor U8343 (N_8343,N_8024,N_8136);
or U8344 (N_8344,N_8110,N_8135);
xor U8345 (N_8345,N_8046,N_8039);
and U8346 (N_8346,N_8175,N_8126);
nand U8347 (N_8347,N_8141,N_8067);
or U8348 (N_8348,N_8096,N_8074);
nor U8349 (N_8349,N_8164,N_8069);
or U8350 (N_8350,N_8182,N_8159);
nor U8351 (N_8351,N_8115,N_8140);
or U8352 (N_8352,N_8096,N_8000);
nor U8353 (N_8353,N_8139,N_8121);
nor U8354 (N_8354,N_8022,N_8166);
nand U8355 (N_8355,N_8158,N_8174);
or U8356 (N_8356,N_8016,N_8015);
nand U8357 (N_8357,N_8096,N_8187);
nor U8358 (N_8358,N_8066,N_8168);
nand U8359 (N_8359,N_8112,N_8024);
or U8360 (N_8360,N_8124,N_8191);
or U8361 (N_8361,N_8007,N_8199);
nand U8362 (N_8362,N_8066,N_8170);
nand U8363 (N_8363,N_8119,N_8191);
nand U8364 (N_8364,N_8110,N_8196);
nand U8365 (N_8365,N_8063,N_8189);
or U8366 (N_8366,N_8048,N_8181);
or U8367 (N_8367,N_8093,N_8011);
xor U8368 (N_8368,N_8131,N_8045);
nor U8369 (N_8369,N_8114,N_8086);
and U8370 (N_8370,N_8079,N_8051);
or U8371 (N_8371,N_8093,N_8171);
and U8372 (N_8372,N_8192,N_8067);
nor U8373 (N_8373,N_8132,N_8043);
nand U8374 (N_8374,N_8084,N_8067);
or U8375 (N_8375,N_8011,N_8106);
xnor U8376 (N_8376,N_8114,N_8173);
or U8377 (N_8377,N_8136,N_8121);
xnor U8378 (N_8378,N_8180,N_8125);
nor U8379 (N_8379,N_8025,N_8166);
and U8380 (N_8380,N_8109,N_8120);
or U8381 (N_8381,N_8016,N_8035);
or U8382 (N_8382,N_8015,N_8027);
nand U8383 (N_8383,N_8155,N_8064);
or U8384 (N_8384,N_8070,N_8180);
xor U8385 (N_8385,N_8115,N_8038);
and U8386 (N_8386,N_8184,N_8181);
nand U8387 (N_8387,N_8073,N_8191);
and U8388 (N_8388,N_8042,N_8059);
and U8389 (N_8389,N_8020,N_8135);
xor U8390 (N_8390,N_8164,N_8051);
and U8391 (N_8391,N_8163,N_8011);
xnor U8392 (N_8392,N_8081,N_8030);
nor U8393 (N_8393,N_8146,N_8060);
or U8394 (N_8394,N_8199,N_8166);
xor U8395 (N_8395,N_8057,N_8034);
nor U8396 (N_8396,N_8007,N_8002);
nor U8397 (N_8397,N_8156,N_8031);
xor U8398 (N_8398,N_8056,N_8062);
and U8399 (N_8399,N_8140,N_8125);
nand U8400 (N_8400,N_8278,N_8310);
xor U8401 (N_8401,N_8263,N_8358);
nand U8402 (N_8402,N_8339,N_8221);
xnor U8403 (N_8403,N_8350,N_8335);
nand U8404 (N_8404,N_8276,N_8302);
nand U8405 (N_8405,N_8215,N_8385);
xor U8406 (N_8406,N_8298,N_8395);
xnor U8407 (N_8407,N_8295,N_8355);
nor U8408 (N_8408,N_8280,N_8206);
and U8409 (N_8409,N_8284,N_8379);
nor U8410 (N_8410,N_8290,N_8325);
or U8411 (N_8411,N_8315,N_8270);
or U8412 (N_8412,N_8305,N_8308);
xor U8413 (N_8413,N_8397,N_8340);
nand U8414 (N_8414,N_8238,N_8234);
nor U8415 (N_8415,N_8211,N_8345);
xnor U8416 (N_8416,N_8248,N_8329);
or U8417 (N_8417,N_8218,N_8285);
xnor U8418 (N_8418,N_8202,N_8399);
and U8419 (N_8419,N_8387,N_8247);
nor U8420 (N_8420,N_8275,N_8341);
nor U8421 (N_8421,N_8360,N_8256);
and U8422 (N_8422,N_8378,N_8210);
and U8423 (N_8423,N_8237,N_8220);
nand U8424 (N_8424,N_8363,N_8351);
nor U8425 (N_8425,N_8318,N_8229);
and U8426 (N_8426,N_8313,N_8373);
xnor U8427 (N_8427,N_8370,N_8236);
and U8428 (N_8428,N_8224,N_8286);
nand U8429 (N_8429,N_8376,N_8214);
and U8430 (N_8430,N_8266,N_8309);
nand U8431 (N_8431,N_8249,N_8391);
nor U8432 (N_8432,N_8364,N_8265);
xor U8433 (N_8433,N_8288,N_8388);
xnor U8434 (N_8434,N_8314,N_8246);
nor U8435 (N_8435,N_8216,N_8271);
nor U8436 (N_8436,N_8316,N_8269);
nor U8437 (N_8437,N_8257,N_8333);
xnor U8438 (N_8438,N_8344,N_8337);
xor U8439 (N_8439,N_8287,N_8331);
nand U8440 (N_8440,N_8203,N_8207);
or U8441 (N_8441,N_8384,N_8368);
xor U8442 (N_8442,N_8289,N_8264);
and U8443 (N_8443,N_8381,N_8226);
nand U8444 (N_8444,N_8204,N_8267);
and U8445 (N_8445,N_8208,N_8394);
nor U8446 (N_8446,N_8235,N_8241);
or U8447 (N_8447,N_8253,N_8297);
nor U8448 (N_8448,N_8259,N_8365);
nand U8449 (N_8449,N_8361,N_8382);
nor U8450 (N_8450,N_8239,N_8349);
and U8451 (N_8451,N_8294,N_8390);
xor U8452 (N_8452,N_8342,N_8304);
nor U8453 (N_8453,N_8320,N_8225);
xor U8454 (N_8454,N_8354,N_8213);
nand U8455 (N_8455,N_8396,N_8352);
nor U8456 (N_8456,N_8343,N_8217);
or U8457 (N_8457,N_8332,N_8347);
and U8458 (N_8458,N_8219,N_8367);
and U8459 (N_8459,N_8323,N_8380);
nor U8460 (N_8460,N_8303,N_8353);
or U8461 (N_8461,N_8228,N_8283);
or U8462 (N_8462,N_8362,N_8356);
or U8463 (N_8463,N_8282,N_8261);
nor U8464 (N_8464,N_8330,N_8324);
and U8465 (N_8465,N_8301,N_8231);
and U8466 (N_8466,N_8205,N_8312);
or U8467 (N_8467,N_8321,N_8245);
or U8468 (N_8468,N_8383,N_8268);
xnor U8469 (N_8469,N_8311,N_8292);
nand U8470 (N_8470,N_8334,N_8291);
or U8471 (N_8471,N_8306,N_8232);
xor U8472 (N_8472,N_8338,N_8209);
and U8473 (N_8473,N_8242,N_8262);
nand U8474 (N_8474,N_8227,N_8375);
nor U8475 (N_8475,N_8348,N_8369);
nand U8476 (N_8476,N_8389,N_8326);
xnor U8477 (N_8477,N_8366,N_8374);
and U8478 (N_8478,N_8371,N_8300);
or U8479 (N_8479,N_8254,N_8252);
or U8480 (N_8480,N_8346,N_8222);
xnor U8481 (N_8481,N_8317,N_8307);
nand U8482 (N_8482,N_8277,N_8274);
and U8483 (N_8483,N_8250,N_8319);
xor U8484 (N_8484,N_8377,N_8279);
nor U8485 (N_8485,N_8392,N_8273);
and U8486 (N_8486,N_8244,N_8255);
or U8487 (N_8487,N_8359,N_8299);
nor U8488 (N_8488,N_8293,N_8243);
nand U8489 (N_8489,N_8233,N_8296);
nand U8490 (N_8490,N_8336,N_8328);
or U8491 (N_8491,N_8398,N_8357);
nand U8492 (N_8492,N_8258,N_8322);
nand U8493 (N_8493,N_8281,N_8201);
and U8494 (N_8494,N_8230,N_8212);
nand U8495 (N_8495,N_8372,N_8272);
xor U8496 (N_8496,N_8240,N_8260);
or U8497 (N_8497,N_8251,N_8393);
nor U8498 (N_8498,N_8386,N_8327);
nand U8499 (N_8499,N_8223,N_8200);
xor U8500 (N_8500,N_8292,N_8245);
or U8501 (N_8501,N_8330,N_8263);
or U8502 (N_8502,N_8244,N_8257);
nand U8503 (N_8503,N_8239,N_8283);
xnor U8504 (N_8504,N_8225,N_8202);
and U8505 (N_8505,N_8284,N_8249);
nand U8506 (N_8506,N_8254,N_8220);
xor U8507 (N_8507,N_8227,N_8215);
nor U8508 (N_8508,N_8363,N_8366);
nor U8509 (N_8509,N_8305,N_8346);
or U8510 (N_8510,N_8391,N_8330);
and U8511 (N_8511,N_8286,N_8207);
and U8512 (N_8512,N_8356,N_8305);
and U8513 (N_8513,N_8308,N_8302);
nand U8514 (N_8514,N_8374,N_8352);
and U8515 (N_8515,N_8374,N_8264);
and U8516 (N_8516,N_8344,N_8252);
nand U8517 (N_8517,N_8331,N_8380);
and U8518 (N_8518,N_8331,N_8279);
nand U8519 (N_8519,N_8309,N_8318);
and U8520 (N_8520,N_8224,N_8335);
xor U8521 (N_8521,N_8320,N_8341);
and U8522 (N_8522,N_8337,N_8347);
or U8523 (N_8523,N_8361,N_8383);
xnor U8524 (N_8524,N_8236,N_8392);
xnor U8525 (N_8525,N_8287,N_8257);
or U8526 (N_8526,N_8223,N_8267);
or U8527 (N_8527,N_8229,N_8210);
and U8528 (N_8528,N_8206,N_8371);
and U8529 (N_8529,N_8341,N_8342);
nand U8530 (N_8530,N_8203,N_8242);
nor U8531 (N_8531,N_8344,N_8207);
xnor U8532 (N_8532,N_8375,N_8216);
nand U8533 (N_8533,N_8397,N_8389);
xnor U8534 (N_8534,N_8397,N_8279);
nand U8535 (N_8535,N_8341,N_8356);
nor U8536 (N_8536,N_8223,N_8224);
xnor U8537 (N_8537,N_8373,N_8266);
xnor U8538 (N_8538,N_8386,N_8231);
nand U8539 (N_8539,N_8379,N_8246);
and U8540 (N_8540,N_8259,N_8358);
nand U8541 (N_8541,N_8367,N_8299);
xor U8542 (N_8542,N_8212,N_8213);
xnor U8543 (N_8543,N_8335,N_8359);
nor U8544 (N_8544,N_8209,N_8327);
nand U8545 (N_8545,N_8227,N_8397);
nand U8546 (N_8546,N_8323,N_8272);
nor U8547 (N_8547,N_8296,N_8300);
or U8548 (N_8548,N_8218,N_8250);
and U8549 (N_8549,N_8266,N_8221);
and U8550 (N_8550,N_8355,N_8337);
xnor U8551 (N_8551,N_8393,N_8318);
nor U8552 (N_8552,N_8239,N_8371);
or U8553 (N_8553,N_8213,N_8252);
or U8554 (N_8554,N_8206,N_8286);
nor U8555 (N_8555,N_8332,N_8302);
nand U8556 (N_8556,N_8387,N_8222);
or U8557 (N_8557,N_8202,N_8307);
nand U8558 (N_8558,N_8374,N_8377);
xnor U8559 (N_8559,N_8220,N_8399);
nand U8560 (N_8560,N_8370,N_8246);
xnor U8561 (N_8561,N_8202,N_8299);
nand U8562 (N_8562,N_8358,N_8326);
nand U8563 (N_8563,N_8207,N_8224);
xor U8564 (N_8564,N_8233,N_8270);
nor U8565 (N_8565,N_8324,N_8316);
xnor U8566 (N_8566,N_8380,N_8282);
or U8567 (N_8567,N_8383,N_8351);
nand U8568 (N_8568,N_8347,N_8328);
nor U8569 (N_8569,N_8242,N_8327);
nand U8570 (N_8570,N_8381,N_8245);
xor U8571 (N_8571,N_8318,N_8314);
xnor U8572 (N_8572,N_8214,N_8324);
and U8573 (N_8573,N_8296,N_8379);
or U8574 (N_8574,N_8252,N_8383);
xnor U8575 (N_8575,N_8382,N_8283);
nor U8576 (N_8576,N_8234,N_8226);
and U8577 (N_8577,N_8332,N_8272);
xnor U8578 (N_8578,N_8320,N_8265);
xor U8579 (N_8579,N_8230,N_8367);
or U8580 (N_8580,N_8363,N_8247);
xor U8581 (N_8581,N_8369,N_8284);
xor U8582 (N_8582,N_8326,N_8288);
and U8583 (N_8583,N_8334,N_8364);
xnor U8584 (N_8584,N_8255,N_8344);
xor U8585 (N_8585,N_8295,N_8351);
or U8586 (N_8586,N_8235,N_8370);
and U8587 (N_8587,N_8325,N_8246);
and U8588 (N_8588,N_8300,N_8270);
or U8589 (N_8589,N_8316,N_8386);
nand U8590 (N_8590,N_8256,N_8343);
nor U8591 (N_8591,N_8223,N_8227);
and U8592 (N_8592,N_8352,N_8391);
and U8593 (N_8593,N_8260,N_8359);
nand U8594 (N_8594,N_8317,N_8251);
xnor U8595 (N_8595,N_8335,N_8373);
or U8596 (N_8596,N_8273,N_8281);
or U8597 (N_8597,N_8290,N_8318);
nand U8598 (N_8598,N_8353,N_8203);
xor U8599 (N_8599,N_8232,N_8317);
or U8600 (N_8600,N_8439,N_8478);
and U8601 (N_8601,N_8510,N_8537);
xnor U8602 (N_8602,N_8539,N_8425);
nor U8603 (N_8603,N_8444,N_8528);
or U8604 (N_8604,N_8483,N_8450);
nand U8605 (N_8605,N_8496,N_8462);
nor U8606 (N_8606,N_8431,N_8557);
nor U8607 (N_8607,N_8429,N_8564);
or U8608 (N_8608,N_8403,N_8596);
xor U8609 (N_8609,N_8445,N_8466);
or U8610 (N_8610,N_8476,N_8477);
and U8611 (N_8611,N_8416,N_8409);
nor U8612 (N_8612,N_8480,N_8518);
and U8613 (N_8613,N_8583,N_8411);
nor U8614 (N_8614,N_8491,N_8458);
nand U8615 (N_8615,N_8543,N_8446);
nand U8616 (N_8616,N_8532,N_8547);
nand U8617 (N_8617,N_8418,N_8512);
nor U8618 (N_8618,N_8567,N_8407);
nand U8619 (N_8619,N_8570,N_8436);
nor U8620 (N_8620,N_8501,N_8454);
or U8621 (N_8621,N_8402,N_8420);
nand U8622 (N_8622,N_8516,N_8423);
nand U8623 (N_8623,N_8560,N_8461);
and U8624 (N_8624,N_8593,N_8424);
nand U8625 (N_8625,N_8542,N_8574);
xnor U8626 (N_8626,N_8434,N_8495);
and U8627 (N_8627,N_8492,N_8555);
nand U8628 (N_8628,N_8587,N_8522);
xor U8629 (N_8629,N_8440,N_8410);
or U8630 (N_8630,N_8447,N_8486);
nor U8631 (N_8631,N_8548,N_8408);
and U8632 (N_8632,N_8580,N_8400);
and U8633 (N_8633,N_8500,N_8467);
and U8634 (N_8634,N_8471,N_8432);
and U8635 (N_8635,N_8511,N_8590);
nor U8636 (N_8636,N_8465,N_8459);
nor U8637 (N_8637,N_8561,N_8493);
and U8638 (N_8638,N_8562,N_8479);
nand U8639 (N_8639,N_8468,N_8517);
nor U8640 (N_8640,N_8415,N_8552);
or U8641 (N_8641,N_8503,N_8451);
xor U8642 (N_8642,N_8598,N_8558);
nand U8643 (N_8643,N_8426,N_8581);
nor U8644 (N_8644,N_8448,N_8455);
or U8645 (N_8645,N_8419,N_8414);
xor U8646 (N_8646,N_8482,N_8531);
or U8647 (N_8647,N_8499,N_8497);
nor U8648 (N_8648,N_8422,N_8515);
and U8649 (N_8649,N_8487,N_8549);
nand U8650 (N_8650,N_8508,N_8591);
nor U8651 (N_8651,N_8433,N_8441);
xor U8652 (N_8652,N_8504,N_8401);
nor U8653 (N_8653,N_8505,N_8437);
nor U8654 (N_8654,N_8563,N_8592);
and U8655 (N_8655,N_8582,N_8442);
xor U8656 (N_8656,N_8559,N_8575);
or U8657 (N_8657,N_8586,N_8525);
nand U8658 (N_8658,N_8453,N_8464);
xnor U8659 (N_8659,N_8481,N_8530);
nor U8660 (N_8660,N_8597,N_8594);
nand U8661 (N_8661,N_8494,N_8578);
xnor U8662 (N_8662,N_8551,N_8488);
xor U8663 (N_8663,N_8460,N_8438);
or U8664 (N_8664,N_8473,N_8584);
or U8665 (N_8665,N_8435,N_8421);
and U8666 (N_8666,N_8538,N_8474);
and U8667 (N_8667,N_8472,N_8475);
and U8668 (N_8668,N_8571,N_8521);
nand U8669 (N_8669,N_8585,N_8577);
or U8670 (N_8670,N_8456,N_8404);
nor U8671 (N_8671,N_8556,N_8536);
or U8672 (N_8672,N_8541,N_8470);
nand U8673 (N_8673,N_8553,N_8509);
nor U8674 (N_8674,N_8507,N_8520);
xor U8675 (N_8675,N_8519,N_8412);
or U8676 (N_8676,N_8430,N_8463);
xnor U8677 (N_8677,N_8514,N_8406);
nand U8678 (N_8678,N_8573,N_8566);
and U8679 (N_8679,N_8545,N_8427);
and U8680 (N_8680,N_8535,N_8534);
nor U8681 (N_8681,N_8449,N_8405);
or U8682 (N_8682,N_8529,N_8452);
nor U8683 (N_8683,N_8569,N_8544);
xor U8684 (N_8684,N_8498,N_8417);
nor U8685 (N_8685,N_8469,N_8579);
nor U8686 (N_8686,N_8485,N_8546);
and U8687 (N_8687,N_8489,N_8589);
xor U8688 (N_8688,N_8484,N_8565);
nor U8689 (N_8689,N_8550,N_8540);
or U8690 (N_8690,N_8490,N_8413);
xnor U8691 (N_8691,N_8554,N_8576);
nor U8692 (N_8692,N_8568,N_8443);
and U8693 (N_8693,N_8526,N_8588);
and U8694 (N_8694,N_8428,N_8513);
nand U8695 (N_8695,N_8457,N_8506);
xor U8696 (N_8696,N_8524,N_8599);
xor U8697 (N_8697,N_8527,N_8533);
xnor U8698 (N_8698,N_8572,N_8523);
nor U8699 (N_8699,N_8502,N_8595);
xnor U8700 (N_8700,N_8572,N_8577);
nor U8701 (N_8701,N_8581,N_8480);
xor U8702 (N_8702,N_8540,N_8590);
and U8703 (N_8703,N_8567,N_8547);
nand U8704 (N_8704,N_8421,N_8507);
nand U8705 (N_8705,N_8593,N_8425);
xor U8706 (N_8706,N_8445,N_8494);
nand U8707 (N_8707,N_8584,N_8427);
or U8708 (N_8708,N_8457,N_8522);
and U8709 (N_8709,N_8484,N_8587);
xor U8710 (N_8710,N_8575,N_8491);
xor U8711 (N_8711,N_8529,N_8585);
nand U8712 (N_8712,N_8585,N_8454);
xor U8713 (N_8713,N_8469,N_8568);
and U8714 (N_8714,N_8585,N_8515);
xnor U8715 (N_8715,N_8412,N_8469);
and U8716 (N_8716,N_8518,N_8532);
nand U8717 (N_8717,N_8458,N_8483);
and U8718 (N_8718,N_8478,N_8485);
xnor U8719 (N_8719,N_8478,N_8490);
nor U8720 (N_8720,N_8594,N_8570);
nor U8721 (N_8721,N_8476,N_8510);
nor U8722 (N_8722,N_8490,N_8439);
nand U8723 (N_8723,N_8466,N_8591);
nand U8724 (N_8724,N_8442,N_8423);
nor U8725 (N_8725,N_8533,N_8555);
nor U8726 (N_8726,N_8412,N_8516);
xnor U8727 (N_8727,N_8401,N_8499);
nor U8728 (N_8728,N_8544,N_8454);
nor U8729 (N_8729,N_8450,N_8599);
nor U8730 (N_8730,N_8456,N_8434);
and U8731 (N_8731,N_8424,N_8470);
nor U8732 (N_8732,N_8411,N_8504);
and U8733 (N_8733,N_8481,N_8497);
or U8734 (N_8734,N_8406,N_8529);
nand U8735 (N_8735,N_8492,N_8548);
and U8736 (N_8736,N_8470,N_8579);
xnor U8737 (N_8737,N_8460,N_8498);
xor U8738 (N_8738,N_8519,N_8599);
or U8739 (N_8739,N_8489,N_8440);
or U8740 (N_8740,N_8493,N_8590);
nand U8741 (N_8741,N_8515,N_8572);
xor U8742 (N_8742,N_8501,N_8510);
or U8743 (N_8743,N_8564,N_8430);
xor U8744 (N_8744,N_8501,N_8410);
nand U8745 (N_8745,N_8496,N_8427);
or U8746 (N_8746,N_8558,N_8458);
or U8747 (N_8747,N_8460,N_8455);
or U8748 (N_8748,N_8521,N_8589);
or U8749 (N_8749,N_8594,N_8471);
nor U8750 (N_8750,N_8519,N_8507);
and U8751 (N_8751,N_8454,N_8404);
or U8752 (N_8752,N_8471,N_8517);
xnor U8753 (N_8753,N_8492,N_8404);
or U8754 (N_8754,N_8516,N_8488);
and U8755 (N_8755,N_8537,N_8449);
or U8756 (N_8756,N_8582,N_8591);
nand U8757 (N_8757,N_8542,N_8451);
nor U8758 (N_8758,N_8506,N_8478);
or U8759 (N_8759,N_8586,N_8441);
nand U8760 (N_8760,N_8449,N_8585);
xnor U8761 (N_8761,N_8597,N_8551);
and U8762 (N_8762,N_8548,N_8437);
nand U8763 (N_8763,N_8400,N_8538);
xor U8764 (N_8764,N_8582,N_8416);
and U8765 (N_8765,N_8465,N_8452);
and U8766 (N_8766,N_8411,N_8452);
xnor U8767 (N_8767,N_8578,N_8466);
nor U8768 (N_8768,N_8432,N_8439);
and U8769 (N_8769,N_8445,N_8533);
and U8770 (N_8770,N_8524,N_8595);
xnor U8771 (N_8771,N_8455,N_8430);
or U8772 (N_8772,N_8457,N_8477);
xnor U8773 (N_8773,N_8595,N_8594);
nand U8774 (N_8774,N_8455,N_8596);
or U8775 (N_8775,N_8411,N_8473);
and U8776 (N_8776,N_8529,N_8552);
or U8777 (N_8777,N_8571,N_8543);
and U8778 (N_8778,N_8581,N_8569);
and U8779 (N_8779,N_8519,N_8487);
xnor U8780 (N_8780,N_8482,N_8541);
nor U8781 (N_8781,N_8435,N_8438);
nor U8782 (N_8782,N_8553,N_8410);
or U8783 (N_8783,N_8547,N_8477);
nor U8784 (N_8784,N_8515,N_8581);
or U8785 (N_8785,N_8583,N_8400);
or U8786 (N_8786,N_8460,N_8427);
nor U8787 (N_8787,N_8486,N_8549);
xor U8788 (N_8788,N_8515,N_8598);
and U8789 (N_8789,N_8597,N_8459);
nor U8790 (N_8790,N_8471,N_8458);
nand U8791 (N_8791,N_8468,N_8485);
and U8792 (N_8792,N_8413,N_8504);
nor U8793 (N_8793,N_8428,N_8569);
nor U8794 (N_8794,N_8511,N_8410);
and U8795 (N_8795,N_8501,N_8584);
nand U8796 (N_8796,N_8405,N_8522);
nand U8797 (N_8797,N_8503,N_8556);
and U8798 (N_8798,N_8529,N_8493);
nand U8799 (N_8799,N_8434,N_8571);
or U8800 (N_8800,N_8612,N_8752);
and U8801 (N_8801,N_8670,N_8601);
nand U8802 (N_8802,N_8683,N_8781);
or U8803 (N_8803,N_8637,N_8716);
xnor U8804 (N_8804,N_8724,N_8749);
and U8805 (N_8805,N_8650,N_8793);
nand U8806 (N_8806,N_8698,N_8773);
nand U8807 (N_8807,N_8762,N_8770);
nor U8808 (N_8808,N_8606,N_8731);
xnor U8809 (N_8809,N_8639,N_8715);
nand U8810 (N_8810,N_8766,N_8680);
xor U8811 (N_8811,N_8662,N_8779);
nand U8812 (N_8812,N_8772,N_8693);
xor U8813 (N_8813,N_8735,N_8712);
and U8814 (N_8814,N_8767,N_8722);
or U8815 (N_8815,N_8728,N_8732);
and U8816 (N_8816,N_8621,N_8763);
and U8817 (N_8817,N_8685,N_8797);
and U8818 (N_8818,N_8681,N_8765);
nor U8819 (N_8819,N_8696,N_8653);
xor U8820 (N_8820,N_8784,N_8655);
or U8821 (N_8821,N_8613,N_8713);
or U8822 (N_8822,N_8786,N_8726);
and U8823 (N_8823,N_8764,N_8631);
nand U8824 (N_8824,N_8633,N_8751);
nand U8825 (N_8825,N_8791,N_8618);
nor U8826 (N_8826,N_8660,N_8743);
nand U8827 (N_8827,N_8604,N_8672);
nor U8828 (N_8828,N_8665,N_8753);
nand U8829 (N_8829,N_8607,N_8795);
xnor U8830 (N_8830,N_8748,N_8616);
nor U8831 (N_8831,N_8656,N_8688);
or U8832 (N_8832,N_8649,N_8630);
nor U8833 (N_8833,N_8709,N_8706);
and U8834 (N_8834,N_8674,N_8792);
nand U8835 (N_8835,N_8669,N_8700);
xor U8836 (N_8836,N_8730,N_8617);
or U8837 (N_8837,N_8744,N_8647);
xnor U8838 (N_8838,N_8788,N_8707);
or U8839 (N_8839,N_8760,N_8652);
and U8840 (N_8840,N_8657,N_8636);
nand U8841 (N_8841,N_8678,N_8739);
or U8842 (N_8842,N_8611,N_8798);
xor U8843 (N_8843,N_8737,N_8721);
nand U8844 (N_8844,N_8704,N_8796);
xor U8845 (N_8845,N_8780,N_8708);
nor U8846 (N_8846,N_8710,N_8648);
and U8847 (N_8847,N_8741,N_8635);
nand U8848 (N_8848,N_8776,N_8642);
nor U8849 (N_8849,N_8646,N_8734);
xnor U8850 (N_8850,N_8628,N_8625);
and U8851 (N_8851,N_8641,N_8783);
nor U8852 (N_8852,N_8690,N_8692);
and U8853 (N_8853,N_8658,N_8759);
or U8854 (N_8854,N_8755,N_8727);
nand U8855 (N_8855,N_8677,N_8640);
or U8856 (N_8856,N_8729,N_8673);
and U8857 (N_8857,N_8758,N_8719);
nor U8858 (N_8858,N_8761,N_8736);
nor U8859 (N_8859,N_8733,N_8750);
nand U8860 (N_8860,N_8620,N_8745);
nand U8861 (N_8861,N_8624,N_8651);
nand U8862 (N_8862,N_8754,N_8775);
nand U8863 (N_8863,N_8723,N_8659);
nor U8864 (N_8864,N_8643,N_8747);
and U8865 (N_8865,N_8768,N_8771);
nor U8866 (N_8866,N_8600,N_8725);
xnor U8867 (N_8867,N_8605,N_8695);
xor U8868 (N_8868,N_8691,N_8711);
nor U8869 (N_8869,N_8663,N_8703);
or U8870 (N_8870,N_8738,N_8623);
nor U8871 (N_8871,N_8668,N_8769);
nand U8872 (N_8872,N_8684,N_8603);
nor U8873 (N_8873,N_8697,N_8757);
nor U8874 (N_8874,N_8644,N_8676);
nor U8875 (N_8875,N_8667,N_8756);
and U8876 (N_8876,N_8789,N_8790);
or U8877 (N_8877,N_8610,N_8627);
or U8878 (N_8878,N_8686,N_8666);
or U8879 (N_8879,N_8785,N_8702);
nand U8880 (N_8880,N_8634,N_8602);
and U8881 (N_8881,N_8687,N_8777);
and U8882 (N_8882,N_8619,N_8664);
xor U8883 (N_8883,N_8632,N_8682);
nand U8884 (N_8884,N_8626,N_8675);
or U8885 (N_8885,N_8614,N_8689);
and U8886 (N_8886,N_8718,N_8699);
and U8887 (N_8887,N_8701,N_8705);
and U8888 (N_8888,N_8720,N_8740);
xnor U8889 (N_8889,N_8794,N_8661);
nand U8890 (N_8890,N_8782,N_8645);
and U8891 (N_8891,N_8638,N_8609);
or U8892 (N_8892,N_8629,N_8615);
xnor U8893 (N_8893,N_8714,N_8746);
and U8894 (N_8894,N_8694,N_8622);
nand U8895 (N_8895,N_8717,N_8671);
and U8896 (N_8896,N_8654,N_8774);
nor U8897 (N_8897,N_8608,N_8778);
nor U8898 (N_8898,N_8679,N_8742);
and U8899 (N_8899,N_8799,N_8787);
or U8900 (N_8900,N_8698,N_8772);
nand U8901 (N_8901,N_8641,N_8705);
and U8902 (N_8902,N_8657,N_8758);
nor U8903 (N_8903,N_8604,N_8748);
nand U8904 (N_8904,N_8631,N_8632);
and U8905 (N_8905,N_8747,N_8796);
nor U8906 (N_8906,N_8782,N_8643);
or U8907 (N_8907,N_8667,N_8703);
nand U8908 (N_8908,N_8798,N_8645);
and U8909 (N_8909,N_8661,N_8778);
xor U8910 (N_8910,N_8649,N_8754);
xnor U8911 (N_8911,N_8625,N_8751);
and U8912 (N_8912,N_8770,N_8791);
nor U8913 (N_8913,N_8753,N_8738);
nor U8914 (N_8914,N_8625,N_8785);
or U8915 (N_8915,N_8636,N_8651);
nor U8916 (N_8916,N_8654,N_8611);
nand U8917 (N_8917,N_8684,N_8672);
nand U8918 (N_8918,N_8623,N_8639);
or U8919 (N_8919,N_8710,N_8722);
nand U8920 (N_8920,N_8786,N_8760);
nor U8921 (N_8921,N_8606,N_8727);
and U8922 (N_8922,N_8716,N_8788);
nor U8923 (N_8923,N_8725,N_8611);
or U8924 (N_8924,N_8735,N_8688);
or U8925 (N_8925,N_8693,N_8717);
or U8926 (N_8926,N_8613,N_8770);
and U8927 (N_8927,N_8693,N_8719);
and U8928 (N_8928,N_8758,N_8641);
xor U8929 (N_8929,N_8749,N_8690);
and U8930 (N_8930,N_8630,N_8776);
xor U8931 (N_8931,N_8718,N_8693);
xor U8932 (N_8932,N_8744,N_8769);
xor U8933 (N_8933,N_8749,N_8682);
and U8934 (N_8934,N_8630,N_8673);
and U8935 (N_8935,N_8737,N_8667);
xnor U8936 (N_8936,N_8757,N_8734);
or U8937 (N_8937,N_8666,N_8715);
nand U8938 (N_8938,N_8706,N_8748);
xor U8939 (N_8939,N_8784,N_8723);
and U8940 (N_8940,N_8771,N_8639);
nor U8941 (N_8941,N_8625,N_8775);
nand U8942 (N_8942,N_8751,N_8754);
or U8943 (N_8943,N_8698,N_8646);
xor U8944 (N_8944,N_8703,N_8625);
nor U8945 (N_8945,N_8635,N_8711);
xor U8946 (N_8946,N_8763,N_8777);
nor U8947 (N_8947,N_8642,N_8654);
or U8948 (N_8948,N_8755,N_8716);
xor U8949 (N_8949,N_8744,N_8610);
or U8950 (N_8950,N_8684,N_8653);
xor U8951 (N_8951,N_8713,N_8628);
or U8952 (N_8952,N_8716,N_8776);
nor U8953 (N_8953,N_8743,N_8747);
nor U8954 (N_8954,N_8740,N_8778);
or U8955 (N_8955,N_8633,N_8707);
xor U8956 (N_8956,N_8646,N_8609);
xnor U8957 (N_8957,N_8696,N_8708);
or U8958 (N_8958,N_8614,N_8769);
nand U8959 (N_8959,N_8665,N_8760);
or U8960 (N_8960,N_8606,N_8677);
or U8961 (N_8961,N_8717,N_8728);
nor U8962 (N_8962,N_8799,N_8754);
or U8963 (N_8963,N_8667,N_8788);
nor U8964 (N_8964,N_8720,N_8759);
and U8965 (N_8965,N_8753,N_8636);
nor U8966 (N_8966,N_8799,N_8790);
and U8967 (N_8967,N_8671,N_8629);
nand U8968 (N_8968,N_8748,N_8605);
and U8969 (N_8969,N_8728,N_8796);
or U8970 (N_8970,N_8672,N_8696);
xor U8971 (N_8971,N_8774,N_8773);
and U8972 (N_8972,N_8710,N_8729);
and U8973 (N_8973,N_8677,N_8666);
nand U8974 (N_8974,N_8619,N_8732);
xnor U8975 (N_8975,N_8616,N_8679);
xor U8976 (N_8976,N_8774,N_8768);
nand U8977 (N_8977,N_8793,N_8761);
and U8978 (N_8978,N_8618,N_8765);
or U8979 (N_8979,N_8607,N_8659);
and U8980 (N_8980,N_8734,N_8695);
and U8981 (N_8981,N_8792,N_8624);
or U8982 (N_8982,N_8765,N_8677);
nand U8983 (N_8983,N_8604,N_8729);
or U8984 (N_8984,N_8774,N_8737);
nand U8985 (N_8985,N_8786,N_8658);
nand U8986 (N_8986,N_8749,N_8600);
nor U8987 (N_8987,N_8617,N_8731);
nor U8988 (N_8988,N_8728,N_8781);
nand U8989 (N_8989,N_8726,N_8784);
nand U8990 (N_8990,N_8766,N_8794);
nand U8991 (N_8991,N_8763,N_8738);
or U8992 (N_8992,N_8734,N_8711);
or U8993 (N_8993,N_8751,N_8755);
or U8994 (N_8994,N_8673,N_8791);
nand U8995 (N_8995,N_8690,N_8728);
or U8996 (N_8996,N_8733,N_8789);
nor U8997 (N_8997,N_8673,N_8617);
nand U8998 (N_8998,N_8763,N_8686);
nor U8999 (N_8999,N_8671,N_8669);
and U9000 (N_9000,N_8881,N_8899);
nor U9001 (N_9001,N_8994,N_8954);
or U9002 (N_9002,N_8979,N_8876);
or U9003 (N_9003,N_8803,N_8961);
xnor U9004 (N_9004,N_8978,N_8897);
nand U9005 (N_9005,N_8810,N_8862);
xor U9006 (N_9006,N_8868,N_8925);
and U9007 (N_9007,N_8814,N_8828);
or U9008 (N_9008,N_8912,N_8920);
and U9009 (N_9009,N_8929,N_8984);
xor U9010 (N_9010,N_8879,N_8940);
nand U9011 (N_9011,N_8817,N_8932);
xnor U9012 (N_9012,N_8953,N_8809);
and U9013 (N_9013,N_8964,N_8894);
nor U9014 (N_9014,N_8808,N_8943);
nor U9015 (N_9015,N_8819,N_8844);
nor U9016 (N_9016,N_8823,N_8873);
or U9017 (N_9017,N_8865,N_8833);
nor U9018 (N_9018,N_8826,N_8860);
nor U9019 (N_9019,N_8805,N_8927);
and U9020 (N_9020,N_8992,N_8822);
nor U9021 (N_9021,N_8840,N_8812);
nand U9022 (N_9022,N_8866,N_8852);
xor U9023 (N_9023,N_8883,N_8821);
and U9024 (N_9024,N_8903,N_8854);
nand U9025 (N_9025,N_8869,N_8872);
nand U9026 (N_9026,N_8995,N_8913);
or U9027 (N_9027,N_8993,N_8848);
nor U9028 (N_9028,N_8838,N_8857);
nor U9029 (N_9029,N_8981,N_8951);
nand U9030 (N_9030,N_8813,N_8829);
nand U9031 (N_9031,N_8858,N_8917);
or U9032 (N_9032,N_8924,N_8971);
nor U9033 (N_9033,N_8907,N_8905);
nand U9034 (N_9034,N_8959,N_8856);
xnor U9035 (N_9035,N_8950,N_8855);
or U9036 (N_9036,N_8887,N_8898);
nor U9037 (N_9037,N_8958,N_8891);
or U9038 (N_9038,N_8987,N_8885);
xnor U9039 (N_9039,N_8933,N_8921);
xor U9040 (N_9040,N_8801,N_8847);
nand U9041 (N_9041,N_8834,N_8939);
or U9042 (N_9042,N_8874,N_8945);
nand U9043 (N_9043,N_8835,N_8928);
nand U9044 (N_9044,N_8851,N_8831);
and U9045 (N_9045,N_8909,N_8991);
xnor U9046 (N_9046,N_8982,N_8989);
nand U9047 (N_9047,N_8906,N_8916);
or U9048 (N_9048,N_8919,N_8893);
or U9049 (N_9049,N_8861,N_8842);
or U9050 (N_9050,N_8941,N_8948);
nor U9051 (N_9051,N_8955,N_8990);
nand U9052 (N_9052,N_8841,N_8914);
nor U9053 (N_9053,N_8931,N_8867);
or U9054 (N_9054,N_8832,N_8870);
or U9055 (N_9055,N_8966,N_8807);
and U9056 (N_9056,N_8902,N_8996);
nand U9057 (N_9057,N_8871,N_8952);
or U9058 (N_9058,N_8908,N_8888);
or U9059 (N_9059,N_8837,N_8944);
nand U9060 (N_9060,N_8864,N_8830);
nor U9061 (N_9061,N_8930,N_8910);
and U9062 (N_9062,N_8892,N_8849);
nand U9063 (N_9063,N_8949,N_8877);
nand U9064 (N_9064,N_8882,N_8886);
nor U9065 (N_9065,N_8922,N_8999);
xor U9066 (N_9066,N_8973,N_8839);
xnor U9067 (N_9067,N_8968,N_8947);
or U9068 (N_9068,N_8977,N_8975);
or U9069 (N_9069,N_8974,N_8880);
nor U9070 (N_9070,N_8818,N_8878);
and U9071 (N_9071,N_8926,N_8998);
nand U9072 (N_9072,N_8859,N_8825);
or U9073 (N_9073,N_8889,N_8976);
and U9074 (N_9074,N_8936,N_8904);
and U9075 (N_9075,N_8875,N_8804);
and U9076 (N_9076,N_8850,N_8923);
or U9077 (N_9077,N_8863,N_8960);
and U9078 (N_9078,N_8970,N_8937);
and U9079 (N_9079,N_8985,N_8853);
xnor U9080 (N_9080,N_8911,N_8988);
nand U9081 (N_9081,N_8935,N_8980);
and U9082 (N_9082,N_8845,N_8956);
or U9083 (N_9083,N_8983,N_8827);
nand U9084 (N_9084,N_8806,N_8972);
or U9085 (N_9085,N_8946,N_8800);
nand U9086 (N_9086,N_8811,N_8836);
nor U9087 (N_9087,N_8890,N_8901);
and U9088 (N_9088,N_8997,N_8938);
or U9089 (N_9089,N_8934,N_8942);
nor U9090 (N_9090,N_8957,N_8884);
xor U9091 (N_9091,N_8802,N_8895);
or U9092 (N_9092,N_8824,N_8986);
or U9093 (N_9093,N_8846,N_8962);
xnor U9094 (N_9094,N_8965,N_8900);
nor U9095 (N_9095,N_8815,N_8915);
nand U9096 (N_9096,N_8967,N_8918);
xnor U9097 (N_9097,N_8969,N_8843);
nor U9098 (N_9098,N_8963,N_8820);
xor U9099 (N_9099,N_8816,N_8896);
or U9100 (N_9100,N_8976,N_8959);
and U9101 (N_9101,N_8856,N_8937);
xor U9102 (N_9102,N_8969,N_8915);
nor U9103 (N_9103,N_8934,N_8896);
or U9104 (N_9104,N_8984,N_8931);
nand U9105 (N_9105,N_8907,N_8820);
nand U9106 (N_9106,N_8864,N_8979);
or U9107 (N_9107,N_8898,N_8891);
nand U9108 (N_9108,N_8837,N_8981);
nand U9109 (N_9109,N_8846,N_8957);
nand U9110 (N_9110,N_8816,N_8853);
or U9111 (N_9111,N_8859,N_8895);
nand U9112 (N_9112,N_8806,N_8829);
and U9113 (N_9113,N_8927,N_8825);
nand U9114 (N_9114,N_8982,N_8907);
nand U9115 (N_9115,N_8823,N_8894);
nand U9116 (N_9116,N_8972,N_8904);
xnor U9117 (N_9117,N_8830,N_8841);
nand U9118 (N_9118,N_8926,N_8848);
and U9119 (N_9119,N_8948,N_8960);
and U9120 (N_9120,N_8867,N_8855);
or U9121 (N_9121,N_8942,N_8961);
and U9122 (N_9122,N_8845,N_8959);
xor U9123 (N_9123,N_8850,N_8946);
xnor U9124 (N_9124,N_8903,N_8848);
xnor U9125 (N_9125,N_8867,N_8822);
and U9126 (N_9126,N_8971,N_8846);
or U9127 (N_9127,N_8857,N_8803);
nand U9128 (N_9128,N_8869,N_8880);
nand U9129 (N_9129,N_8933,N_8854);
xor U9130 (N_9130,N_8948,N_8890);
or U9131 (N_9131,N_8912,N_8810);
nand U9132 (N_9132,N_8868,N_8949);
nor U9133 (N_9133,N_8819,N_8971);
nor U9134 (N_9134,N_8823,N_8985);
and U9135 (N_9135,N_8862,N_8899);
and U9136 (N_9136,N_8964,N_8919);
or U9137 (N_9137,N_8926,N_8874);
and U9138 (N_9138,N_8819,N_8959);
or U9139 (N_9139,N_8904,N_8814);
nand U9140 (N_9140,N_8898,N_8856);
nor U9141 (N_9141,N_8839,N_8979);
and U9142 (N_9142,N_8987,N_8858);
and U9143 (N_9143,N_8916,N_8977);
and U9144 (N_9144,N_8924,N_8862);
and U9145 (N_9145,N_8874,N_8907);
nand U9146 (N_9146,N_8880,N_8923);
or U9147 (N_9147,N_8974,N_8879);
nand U9148 (N_9148,N_8994,N_8819);
or U9149 (N_9149,N_8973,N_8858);
nor U9150 (N_9150,N_8952,N_8935);
or U9151 (N_9151,N_8837,N_8984);
nor U9152 (N_9152,N_8857,N_8831);
and U9153 (N_9153,N_8898,N_8877);
and U9154 (N_9154,N_8818,N_8877);
and U9155 (N_9155,N_8942,N_8966);
nor U9156 (N_9156,N_8861,N_8943);
and U9157 (N_9157,N_8903,N_8820);
or U9158 (N_9158,N_8828,N_8838);
and U9159 (N_9159,N_8801,N_8966);
and U9160 (N_9160,N_8975,N_8899);
and U9161 (N_9161,N_8802,N_8890);
and U9162 (N_9162,N_8873,N_8872);
xnor U9163 (N_9163,N_8991,N_8813);
xnor U9164 (N_9164,N_8816,N_8843);
or U9165 (N_9165,N_8984,N_8961);
or U9166 (N_9166,N_8855,N_8981);
nor U9167 (N_9167,N_8840,N_8801);
nor U9168 (N_9168,N_8951,N_8942);
or U9169 (N_9169,N_8943,N_8934);
xor U9170 (N_9170,N_8813,N_8980);
nand U9171 (N_9171,N_8991,N_8944);
and U9172 (N_9172,N_8828,N_8887);
xor U9173 (N_9173,N_8904,N_8885);
nor U9174 (N_9174,N_8808,N_8854);
and U9175 (N_9175,N_8981,N_8917);
xor U9176 (N_9176,N_8867,N_8832);
and U9177 (N_9177,N_8867,N_8996);
xor U9178 (N_9178,N_8983,N_8867);
or U9179 (N_9179,N_8927,N_8972);
or U9180 (N_9180,N_8929,N_8864);
xor U9181 (N_9181,N_8879,N_8898);
nand U9182 (N_9182,N_8888,N_8852);
nand U9183 (N_9183,N_8842,N_8962);
nand U9184 (N_9184,N_8845,N_8881);
xnor U9185 (N_9185,N_8826,N_8831);
xnor U9186 (N_9186,N_8971,N_8831);
nand U9187 (N_9187,N_8919,N_8896);
xor U9188 (N_9188,N_8992,N_8818);
nor U9189 (N_9189,N_8949,N_8954);
and U9190 (N_9190,N_8951,N_8993);
xor U9191 (N_9191,N_8993,N_8871);
xor U9192 (N_9192,N_8836,N_8953);
or U9193 (N_9193,N_8847,N_8992);
nor U9194 (N_9194,N_8985,N_8844);
xor U9195 (N_9195,N_8891,N_8802);
and U9196 (N_9196,N_8886,N_8832);
xor U9197 (N_9197,N_8913,N_8999);
nand U9198 (N_9198,N_8971,N_8870);
nor U9199 (N_9199,N_8943,N_8896);
and U9200 (N_9200,N_9163,N_9122);
and U9201 (N_9201,N_9028,N_9164);
or U9202 (N_9202,N_9167,N_9171);
nand U9203 (N_9203,N_9121,N_9099);
and U9204 (N_9204,N_9187,N_9084);
or U9205 (N_9205,N_9117,N_9166);
and U9206 (N_9206,N_9114,N_9052);
and U9207 (N_9207,N_9103,N_9046);
nor U9208 (N_9208,N_9079,N_9105);
nor U9209 (N_9209,N_9081,N_9075);
nor U9210 (N_9210,N_9051,N_9186);
nand U9211 (N_9211,N_9199,N_9038);
xnor U9212 (N_9212,N_9024,N_9080);
nor U9213 (N_9213,N_9193,N_9062);
and U9214 (N_9214,N_9009,N_9030);
or U9215 (N_9215,N_9053,N_9148);
or U9216 (N_9216,N_9029,N_9093);
nand U9217 (N_9217,N_9017,N_9184);
and U9218 (N_9218,N_9194,N_9014);
nor U9219 (N_9219,N_9133,N_9174);
nor U9220 (N_9220,N_9144,N_9097);
and U9221 (N_9221,N_9137,N_9160);
xor U9222 (N_9222,N_9073,N_9043);
and U9223 (N_9223,N_9092,N_9027);
or U9224 (N_9224,N_9112,N_9107);
or U9225 (N_9225,N_9153,N_9087);
or U9226 (N_9226,N_9070,N_9151);
and U9227 (N_9227,N_9188,N_9002);
or U9228 (N_9228,N_9124,N_9150);
or U9229 (N_9229,N_9086,N_9198);
nand U9230 (N_9230,N_9060,N_9101);
and U9231 (N_9231,N_9031,N_9104);
xor U9232 (N_9232,N_9021,N_9015);
xnor U9233 (N_9233,N_9000,N_9077);
xnor U9234 (N_9234,N_9019,N_9094);
or U9235 (N_9235,N_9130,N_9047);
nor U9236 (N_9236,N_9149,N_9018);
or U9237 (N_9237,N_9197,N_9040);
nand U9238 (N_9238,N_9145,N_9135);
or U9239 (N_9239,N_9126,N_9066);
and U9240 (N_9240,N_9123,N_9162);
or U9241 (N_9241,N_9158,N_9057);
and U9242 (N_9242,N_9128,N_9055);
or U9243 (N_9243,N_9134,N_9168);
or U9244 (N_9244,N_9006,N_9192);
and U9245 (N_9245,N_9195,N_9156);
nor U9246 (N_9246,N_9049,N_9115);
nand U9247 (N_9247,N_9143,N_9102);
and U9248 (N_9248,N_9147,N_9089);
nand U9249 (N_9249,N_9085,N_9118);
or U9250 (N_9250,N_9146,N_9165);
xnor U9251 (N_9251,N_9191,N_9106);
xor U9252 (N_9252,N_9025,N_9007);
xnor U9253 (N_9253,N_9076,N_9068);
or U9254 (N_9254,N_9119,N_9056);
and U9255 (N_9255,N_9120,N_9152);
or U9256 (N_9256,N_9141,N_9196);
xor U9257 (N_9257,N_9010,N_9178);
or U9258 (N_9258,N_9078,N_9035);
and U9259 (N_9259,N_9059,N_9058);
and U9260 (N_9260,N_9169,N_9176);
nor U9261 (N_9261,N_9067,N_9100);
xnor U9262 (N_9262,N_9142,N_9065);
or U9263 (N_9263,N_9033,N_9008);
nor U9264 (N_9264,N_9136,N_9154);
xnor U9265 (N_9265,N_9177,N_9189);
and U9266 (N_9266,N_9175,N_9044);
nand U9267 (N_9267,N_9036,N_9069);
or U9268 (N_9268,N_9039,N_9096);
nor U9269 (N_9269,N_9042,N_9155);
and U9270 (N_9270,N_9173,N_9083);
and U9271 (N_9271,N_9125,N_9071);
xnor U9272 (N_9272,N_9001,N_9016);
xor U9273 (N_9273,N_9063,N_9020);
or U9274 (N_9274,N_9127,N_9034);
nand U9275 (N_9275,N_9109,N_9111);
or U9276 (N_9276,N_9098,N_9183);
and U9277 (N_9277,N_9032,N_9091);
and U9278 (N_9278,N_9140,N_9090);
or U9279 (N_9279,N_9180,N_9190);
nand U9280 (N_9280,N_9045,N_9061);
nor U9281 (N_9281,N_9023,N_9082);
or U9282 (N_9282,N_9108,N_9132);
nand U9283 (N_9283,N_9074,N_9159);
nor U9284 (N_9284,N_9138,N_9003);
xnor U9285 (N_9285,N_9185,N_9026);
or U9286 (N_9286,N_9041,N_9095);
or U9287 (N_9287,N_9110,N_9157);
and U9288 (N_9288,N_9139,N_9012);
nor U9289 (N_9289,N_9022,N_9131);
nor U9290 (N_9290,N_9161,N_9072);
nor U9291 (N_9291,N_9048,N_9172);
xor U9292 (N_9292,N_9181,N_9054);
xnor U9293 (N_9293,N_9004,N_9011);
xnor U9294 (N_9294,N_9170,N_9013);
and U9295 (N_9295,N_9005,N_9037);
nor U9296 (N_9296,N_9129,N_9088);
nand U9297 (N_9297,N_9113,N_9179);
xnor U9298 (N_9298,N_9182,N_9050);
or U9299 (N_9299,N_9064,N_9116);
nand U9300 (N_9300,N_9192,N_9161);
xnor U9301 (N_9301,N_9048,N_9182);
nor U9302 (N_9302,N_9111,N_9194);
or U9303 (N_9303,N_9119,N_9023);
nor U9304 (N_9304,N_9034,N_9063);
and U9305 (N_9305,N_9095,N_9154);
nand U9306 (N_9306,N_9082,N_9078);
or U9307 (N_9307,N_9027,N_9127);
and U9308 (N_9308,N_9026,N_9028);
nor U9309 (N_9309,N_9137,N_9197);
nand U9310 (N_9310,N_9100,N_9089);
or U9311 (N_9311,N_9003,N_9040);
nand U9312 (N_9312,N_9170,N_9008);
and U9313 (N_9313,N_9036,N_9088);
and U9314 (N_9314,N_9087,N_9187);
nor U9315 (N_9315,N_9114,N_9122);
and U9316 (N_9316,N_9179,N_9056);
nor U9317 (N_9317,N_9029,N_9128);
xor U9318 (N_9318,N_9103,N_9194);
and U9319 (N_9319,N_9116,N_9031);
xnor U9320 (N_9320,N_9131,N_9121);
and U9321 (N_9321,N_9160,N_9199);
or U9322 (N_9322,N_9017,N_9116);
nand U9323 (N_9323,N_9034,N_9169);
or U9324 (N_9324,N_9077,N_9143);
nand U9325 (N_9325,N_9028,N_9146);
nand U9326 (N_9326,N_9103,N_9136);
and U9327 (N_9327,N_9166,N_9077);
nand U9328 (N_9328,N_9097,N_9000);
nand U9329 (N_9329,N_9073,N_9171);
nor U9330 (N_9330,N_9076,N_9009);
nor U9331 (N_9331,N_9014,N_9106);
nor U9332 (N_9332,N_9149,N_9038);
and U9333 (N_9333,N_9170,N_9074);
nor U9334 (N_9334,N_9191,N_9152);
nor U9335 (N_9335,N_9119,N_9163);
or U9336 (N_9336,N_9141,N_9013);
nand U9337 (N_9337,N_9157,N_9070);
xor U9338 (N_9338,N_9121,N_9178);
nor U9339 (N_9339,N_9137,N_9039);
nor U9340 (N_9340,N_9162,N_9157);
nand U9341 (N_9341,N_9170,N_9105);
or U9342 (N_9342,N_9070,N_9180);
xor U9343 (N_9343,N_9061,N_9170);
xnor U9344 (N_9344,N_9183,N_9061);
xnor U9345 (N_9345,N_9160,N_9133);
nand U9346 (N_9346,N_9090,N_9072);
nor U9347 (N_9347,N_9012,N_9143);
or U9348 (N_9348,N_9001,N_9174);
or U9349 (N_9349,N_9040,N_9002);
xor U9350 (N_9350,N_9188,N_9013);
xnor U9351 (N_9351,N_9124,N_9033);
nor U9352 (N_9352,N_9150,N_9059);
nor U9353 (N_9353,N_9119,N_9039);
nor U9354 (N_9354,N_9113,N_9125);
nand U9355 (N_9355,N_9129,N_9174);
nand U9356 (N_9356,N_9066,N_9016);
nand U9357 (N_9357,N_9084,N_9077);
and U9358 (N_9358,N_9152,N_9012);
or U9359 (N_9359,N_9032,N_9073);
nor U9360 (N_9360,N_9159,N_9011);
nor U9361 (N_9361,N_9100,N_9025);
or U9362 (N_9362,N_9190,N_9005);
or U9363 (N_9363,N_9173,N_9023);
nand U9364 (N_9364,N_9001,N_9045);
nand U9365 (N_9365,N_9107,N_9196);
or U9366 (N_9366,N_9103,N_9002);
xnor U9367 (N_9367,N_9090,N_9165);
nand U9368 (N_9368,N_9067,N_9082);
xor U9369 (N_9369,N_9009,N_9080);
nor U9370 (N_9370,N_9058,N_9087);
nand U9371 (N_9371,N_9159,N_9180);
nor U9372 (N_9372,N_9093,N_9089);
nor U9373 (N_9373,N_9037,N_9051);
nand U9374 (N_9374,N_9132,N_9119);
and U9375 (N_9375,N_9038,N_9138);
nor U9376 (N_9376,N_9110,N_9069);
xor U9377 (N_9377,N_9025,N_9094);
nand U9378 (N_9378,N_9050,N_9046);
and U9379 (N_9379,N_9032,N_9189);
and U9380 (N_9380,N_9033,N_9045);
nor U9381 (N_9381,N_9112,N_9097);
nor U9382 (N_9382,N_9113,N_9199);
or U9383 (N_9383,N_9140,N_9129);
or U9384 (N_9384,N_9037,N_9077);
and U9385 (N_9385,N_9065,N_9166);
nand U9386 (N_9386,N_9153,N_9040);
and U9387 (N_9387,N_9031,N_9049);
xor U9388 (N_9388,N_9042,N_9166);
nor U9389 (N_9389,N_9003,N_9080);
or U9390 (N_9390,N_9040,N_9041);
nor U9391 (N_9391,N_9121,N_9110);
or U9392 (N_9392,N_9123,N_9049);
xor U9393 (N_9393,N_9001,N_9017);
and U9394 (N_9394,N_9141,N_9026);
or U9395 (N_9395,N_9094,N_9065);
nand U9396 (N_9396,N_9047,N_9078);
and U9397 (N_9397,N_9155,N_9128);
or U9398 (N_9398,N_9102,N_9100);
xor U9399 (N_9399,N_9058,N_9083);
nand U9400 (N_9400,N_9382,N_9238);
xnor U9401 (N_9401,N_9322,N_9266);
nor U9402 (N_9402,N_9388,N_9327);
nor U9403 (N_9403,N_9334,N_9253);
and U9404 (N_9404,N_9227,N_9330);
and U9405 (N_9405,N_9301,N_9352);
nand U9406 (N_9406,N_9343,N_9347);
and U9407 (N_9407,N_9201,N_9296);
nor U9408 (N_9408,N_9243,N_9284);
and U9409 (N_9409,N_9306,N_9293);
nor U9410 (N_9410,N_9254,N_9361);
and U9411 (N_9411,N_9211,N_9289);
or U9412 (N_9412,N_9267,N_9274);
nand U9413 (N_9413,N_9256,N_9329);
nand U9414 (N_9414,N_9335,N_9323);
nand U9415 (N_9415,N_9321,N_9264);
nor U9416 (N_9416,N_9362,N_9351);
nor U9417 (N_9417,N_9360,N_9369);
nand U9418 (N_9418,N_9390,N_9270);
or U9419 (N_9419,N_9288,N_9255);
or U9420 (N_9420,N_9358,N_9318);
and U9421 (N_9421,N_9367,N_9282);
nor U9422 (N_9422,N_9204,N_9278);
and U9423 (N_9423,N_9275,N_9345);
nor U9424 (N_9424,N_9313,N_9210);
and U9425 (N_9425,N_9220,N_9355);
and U9426 (N_9426,N_9200,N_9228);
nand U9427 (N_9427,N_9315,N_9260);
nor U9428 (N_9428,N_9257,N_9385);
or U9429 (N_9429,N_9250,N_9280);
xor U9430 (N_9430,N_9205,N_9237);
xnor U9431 (N_9431,N_9249,N_9374);
xor U9432 (N_9432,N_9309,N_9396);
nand U9433 (N_9433,N_9217,N_9319);
and U9434 (N_9434,N_9245,N_9341);
and U9435 (N_9435,N_9252,N_9276);
nand U9436 (N_9436,N_9261,N_9379);
or U9437 (N_9437,N_9285,N_9277);
xor U9438 (N_9438,N_9308,N_9348);
nand U9439 (N_9439,N_9234,N_9221);
nor U9440 (N_9440,N_9356,N_9246);
and U9441 (N_9441,N_9392,N_9202);
or U9442 (N_9442,N_9224,N_9225);
nor U9443 (N_9443,N_9300,N_9279);
xnor U9444 (N_9444,N_9287,N_9337);
nor U9445 (N_9445,N_9258,N_9214);
nor U9446 (N_9446,N_9320,N_9305);
xnor U9447 (N_9447,N_9378,N_9357);
nor U9448 (N_9448,N_9286,N_9241);
and U9449 (N_9449,N_9375,N_9219);
xnor U9450 (N_9450,N_9304,N_9230);
xnor U9451 (N_9451,N_9244,N_9283);
nor U9452 (N_9452,N_9317,N_9368);
and U9453 (N_9453,N_9251,N_9353);
or U9454 (N_9454,N_9269,N_9248);
xor U9455 (N_9455,N_9271,N_9370);
xnor U9456 (N_9456,N_9222,N_9294);
xor U9457 (N_9457,N_9399,N_9218);
xor U9458 (N_9458,N_9298,N_9311);
and U9459 (N_9459,N_9207,N_9310);
or U9460 (N_9460,N_9312,N_9339);
and U9461 (N_9461,N_9340,N_9397);
xor U9462 (N_9462,N_9328,N_9366);
xnor U9463 (N_9463,N_9203,N_9232);
and U9464 (N_9464,N_9235,N_9297);
and U9465 (N_9465,N_9342,N_9216);
nor U9466 (N_9466,N_9262,N_9391);
nand U9467 (N_9467,N_9331,N_9354);
and U9468 (N_9468,N_9336,N_9389);
nor U9469 (N_9469,N_9380,N_9333);
and U9470 (N_9470,N_9363,N_9398);
and U9471 (N_9471,N_9299,N_9387);
nand U9472 (N_9472,N_9303,N_9229);
xor U9473 (N_9473,N_9359,N_9212);
nor U9474 (N_9474,N_9349,N_9247);
nand U9475 (N_9475,N_9236,N_9281);
and U9476 (N_9476,N_9307,N_9302);
and U9477 (N_9477,N_9215,N_9364);
and U9478 (N_9478,N_9332,N_9242);
and U9479 (N_9479,N_9263,N_9223);
or U9480 (N_9480,N_9372,N_9384);
and U9481 (N_9481,N_9316,N_9314);
xor U9482 (N_9482,N_9239,N_9259);
nand U9483 (N_9483,N_9394,N_9213);
xor U9484 (N_9484,N_9324,N_9383);
nor U9485 (N_9485,N_9338,N_9209);
xnor U9486 (N_9486,N_9240,N_9265);
nand U9487 (N_9487,N_9344,N_9233);
or U9488 (N_9488,N_9325,N_9371);
nor U9489 (N_9489,N_9377,N_9346);
xor U9490 (N_9490,N_9231,N_9273);
nand U9491 (N_9491,N_9206,N_9272);
and U9492 (N_9492,N_9226,N_9373);
or U9493 (N_9493,N_9268,N_9295);
and U9494 (N_9494,N_9365,N_9291);
or U9495 (N_9495,N_9393,N_9395);
nor U9496 (N_9496,N_9326,N_9386);
xnor U9497 (N_9497,N_9376,N_9381);
or U9498 (N_9498,N_9208,N_9290);
xor U9499 (N_9499,N_9292,N_9350);
and U9500 (N_9500,N_9293,N_9353);
or U9501 (N_9501,N_9202,N_9204);
nor U9502 (N_9502,N_9354,N_9386);
nand U9503 (N_9503,N_9351,N_9251);
and U9504 (N_9504,N_9272,N_9254);
or U9505 (N_9505,N_9379,N_9268);
xor U9506 (N_9506,N_9324,N_9209);
xor U9507 (N_9507,N_9224,N_9239);
nor U9508 (N_9508,N_9282,N_9349);
and U9509 (N_9509,N_9273,N_9283);
and U9510 (N_9510,N_9302,N_9265);
xor U9511 (N_9511,N_9272,N_9292);
or U9512 (N_9512,N_9325,N_9261);
xor U9513 (N_9513,N_9310,N_9274);
and U9514 (N_9514,N_9289,N_9318);
or U9515 (N_9515,N_9384,N_9326);
or U9516 (N_9516,N_9337,N_9327);
xnor U9517 (N_9517,N_9216,N_9204);
and U9518 (N_9518,N_9378,N_9338);
nand U9519 (N_9519,N_9393,N_9203);
nor U9520 (N_9520,N_9203,N_9240);
nand U9521 (N_9521,N_9335,N_9291);
nor U9522 (N_9522,N_9293,N_9375);
nor U9523 (N_9523,N_9396,N_9327);
and U9524 (N_9524,N_9280,N_9347);
xor U9525 (N_9525,N_9399,N_9282);
or U9526 (N_9526,N_9357,N_9306);
nand U9527 (N_9527,N_9276,N_9234);
and U9528 (N_9528,N_9285,N_9302);
and U9529 (N_9529,N_9255,N_9390);
xnor U9530 (N_9530,N_9346,N_9233);
xor U9531 (N_9531,N_9328,N_9397);
and U9532 (N_9532,N_9251,N_9382);
xor U9533 (N_9533,N_9346,N_9245);
nor U9534 (N_9534,N_9353,N_9267);
nand U9535 (N_9535,N_9274,N_9297);
nor U9536 (N_9536,N_9208,N_9203);
or U9537 (N_9537,N_9250,N_9323);
and U9538 (N_9538,N_9353,N_9225);
nor U9539 (N_9539,N_9292,N_9255);
and U9540 (N_9540,N_9266,N_9367);
or U9541 (N_9541,N_9267,N_9384);
or U9542 (N_9542,N_9342,N_9371);
xor U9543 (N_9543,N_9314,N_9395);
nand U9544 (N_9544,N_9358,N_9201);
nor U9545 (N_9545,N_9217,N_9309);
nor U9546 (N_9546,N_9245,N_9372);
xnor U9547 (N_9547,N_9219,N_9254);
nor U9548 (N_9548,N_9315,N_9324);
and U9549 (N_9549,N_9266,N_9274);
xnor U9550 (N_9550,N_9325,N_9250);
nor U9551 (N_9551,N_9389,N_9365);
or U9552 (N_9552,N_9352,N_9222);
nand U9553 (N_9553,N_9267,N_9359);
xor U9554 (N_9554,N_9397,N_9233);
or U9555 (N_9555,N_9222,N_9231);
nor U9556 (N_9556,N_9252,N_9235);
or U9557 (N_9557,N_9239,N_9312);
xor U9558 (N_9558,N_9253,N_9277);
nor U9559 (N_9559,N_9338,N_9248);
and U9560 (N_9560,N_9241,N_9217);
nor U9561 (N_9561,N_9295,N_9292);
nor U9562 (N_9562,N_9359,N_9376);
or U9563 (N_9563,N_9365,N_9293);
nand U9564 (N_9564,N_9301,N_9333);
or U9565 (N_9565,N_9313,N_9256);
nand U9566 (N_9566,N_9304,N_9327);
nand U9567 (N_9567,N_9259,N_9383);
nor U9568 (N_9568,N_9363,N_9302);
nor U9569 (N_9569,N_9210,N_9227);
nand U9570 (N_9570,N_9386,N_9315);
xor U9571 (N_9571,N_9244,N_9267);
and U9572 (N_9572,N_9255,N_9242);
nor U9573 (N_9573,N_9316,N_9215);
nor U9574 (N_9574,N_9244,N_9307);
nor U9575 (N_9575,N_9269,N_9300);
nand U9576 (N_9576,N_9315,N_9290);
and U9577 (N_9577,N_9227,N_9247);
xnor U9578 (N_9578,N_9378,N_9278);
or U9579 (N_9579,N_9255,N_9391);
xnor U9580 (N_9580,N_9392,N_9245);
xor U9581 (N_9581,N_9399,N_9333);
and U9582 (N_9582,N_9297,N_9383);
or U9583 (N_9583,N_9372,N_9391);
nor U9584 (N_9584,N_9245,N_9248);
nand U9585 (N_9585,N_9370,N_9263);
and U9586 (N_9586,N_9303,N_9258);
nand U9587 (N_9587,N_9355,N_9380);
xnor U9588 (N_9588,N_9378,N_9242);
xnor U9589 (N_9589,N_9285,N_9267);
and U9590 (N_9590,N_9200,N_9325);
xor U9591 (N_9591,N_9328,N_9294);
or U9592 (N_9592,N_9374,N_9327);
nand U9593 (N_9593,N_9318,N_9228);
and U9594 (N_9594,N_9357,N_9350);
xnor U9595 (N_9595,N_9220,N_9311);
or U9596 (N_9596,N_9324,N_9393);
and U9597 (N_9597,N_9284,N_9299);
or U9598 (N_9598,N_9341,N_9321);
or U9599 (N_9599,N_9341,N_9232);
nand U9600 (N_9600,N_9556,N_9534);
and U9601 (N_9601,N_9525,N_9417);
or U9602 (N_9602,N_9549,N_9467);
nor U9603 (N_9603,N_9518,N_9486);
xor U9604 (N_9604,N_9506,N_9435);
nor U9605 (N_9605,N_9434,N_9451);
nor U9606 (N_9606,N_9481,N_9414);
nor U9607 (N_9607,N_9421,N_9497);
and U9608 (N_9608,N_9543,N_9589);
nand U9609 (N_9609,N_9469,N_9483);
or U9610 (N_9610,N_9429,N_9465);
and U9611 (N_9611,N_9541,N_9564);
and U9612 (N_9612,N_9427,N_9570);
or U9613 (N_9613,N_9586,N_9412);
nand U9614 (N_9614,N_9575,N_9544);
and U9615 (N_9615,N_9474,N_9471);
nor U9616 (N_9616,N_9598,N_9425);
or U9617 (N_9617,N_9475,N_9487);
xor U9618 (N_9618,N_9515,N_9576);
xnor U9619 (N_9619,N_9594,N_9583);
and U9620 (N_9620,N_9446,N_9500);
nand U9621 (N_9621,N_9561,N_9512);
xor U9622 (N_9622,N_9519,N_9579);
nor U9623 (N_9623,N_9513,N_9522);
nand U9624 (N_9624,N_9562,N_9504);
and U9625 (N_9625,N_9418,N_9565);
and U9626 (N_9626,N_9533,N_9440);
xnor U9627 (N_9627,N_9479,N_9490);
nor U9628 (N_9628,N_9404,N_9463);
or U9629 (N_9629,N_9529,N_9585);
and U9630 (N_9630,N_9595,N_9431);
nand U9631 (N_9631,N_9577,N_9539);
xor U9632 (N_9632,N_9596,N_9400);
or U9633 (N_9633,N_9457,N_9540);
or U9634 (N_9634,N_9447,N_9532);
nand U9635 (N_9635,N_9423,N_9547);
nor U9636 (N_9636,N_9505,N_9593);
nand U9637 (N_9637,N_9439,N_9563);
and U9638 (N_9638,N_9426,N_9551);
or U9639 (N_9639,N_9507,N_9436);
or U9640 (N_9640,N_9550,N_9492);
nand U9641 (N_9641,N_9413,N_9588);
xnor U9642 (N_9642,N_9542,N_9408);
or U9643 (N_9643,N_9578,N_9458);
nand U9644 (N_9644,N_9514,N_9555);
nand U9645 (N_9645,N_9489,N_9557);
xnor U9646 (N_9646,N_9510,N_9537);
nand U9647 (N_9647,N_9580,N_9437);
nor U9648 (N_9648,N_9493,N_9597);
or U9649 (N_9649,N_9432,N_9528);
nand U9650 (N_9650,N_9511,N_9484);
xor U9651 (N_9651,N_9503,N_9464);
nand U9652 (N_9652,N_9480,N_9590);
and U9653 (N_9653,N_9476,N_9462);
nand U9654 (N_9654,N_9402,N_9401);
xor U9655 (N_9655,N_9523,N_9571);
xor U9656 (N_9656,N_9526,N_9407);
xor U9657 (N_9657,N_9461,N_9494);
or U9658 (N_9658,N_9456,N_9430);
or U9659 (N_9659,N_9478,N_9442);
and U9660 (N_9660,N_9454,N_9568);
or U9661 (N_9661,N_9419,N_9449);
or U9662 (N_9662,N_9524,N_9485);
nand U9663 (N_9663,N_9411,N_9569);
and U9664 (N_9664,N_9517,N_9482);
and U9665 (N_9665,N_9501,N_9558);
nand U9666 (N_9666,N_9520,N_9488);
nand U9667 (N_9667,N_9591,N_9582);
nor U9668 (N_9668,N_9498,N_9448);
or U9669 (N_9669,N_9445,N_9516);
and U9670 (N_9670,N_9466,N_9502);
or U9671 (N_9671,N_9574,N_9468);
nand U9672 (N_9672,N_9415,N_9496);
and U9673 (N_9673,N_9592,N_9554);
xor U9674 (N_9674,N_9530,N_9455);
nand U9675 (N_9675,N_9531,N_9420);
nand U9676 (N_9676,N_9409,N_9491);
and U9677 (N_9677,N_9403,N_9473);
xnor U9678 (N_9678,N_9422,N_9552);
and U9679 (N_9679,N_9416,N_9460);
and U9680 (N_9680,N_9548,N_9560);
or U9681 (N_9681,N_9584,N_9453);
nand U9682 (N_9682,N_9545,N_9566);
and U9683 (N_9683,N_9450,N_9438);
nand U9684 (N_9684,N_9567,N_9509);
or U9685 (N_9685,N_9599,N_9433);
nor U9686 (N_9686,N_9581,N_9572);
xnor U9687 (N_9687,N_9546,N_9535);
nor U9688 (N_9688,N_9527,N_9521);
and U9689 (N_9689,N_9508,N_9452);
and U9690 (N_9690,N_9573,N_9405);
nand U9691 (N_9691,N_9587,N_9470);
nor U9692 (N_9692,N_9553,N_9424);
or U9693 (N_9693,N_9444,N_9472);
nor U9694 (N_9694,N_9443,N_9459);
or U9695 (N_9695,N_9559,N_9477);
nand U9696 (N_9696,N_9410,N_9536);
or U9697 (N_9697,N_9538,N_9428);
nand U9698 (N_9698,N_9495,N_9441);
and U9699 (N_9699,N_9406,N_9499);
and U9700 (N_9700,N_9455,N_9583);
nor U9701 (N_9701,N_9461,N_9591);
nor U9702 (N_9702,N_9496,N_9587);
nand U9703 (N_9703,N_9408,N_9426);
xnor U9704 (N_9704,N_9516,N_9404);
nand U9705 (N_9705,N_9445,N_9405);
xor U9706 (N_9706,N_9483,N_9548);
and U9707 (N_9707,N_9560,N_9578);
and U9708 (N_9708,N_9516,N_9518);
or U9709 (N_9709,N_9474,N_9592);
xor U9710 (N_9710,N_9452,N_9593);
xnor U9711 (N_9711,N_9416,N_9507);
nand U9712 (N_9712,N_9408,N_9576);
and U9713 (N_9713,N_9504,N_9447);
nand U9714 (N_9714,N_9408,N_9593);
nor U9715 (N_9715,N_9474,N_9562);
and U9716 (N_9716,N_9542,N_9498);
or U9717 (N_9717,N_9511,N_9492);
nor U9718 (N_9718,N_9511,N_9579);
nand U9719 (N_9719,N_9599,N_9494);
nand U9720 (N_9720,N_9586,N_9419);
and U9721 (N_9721,N_9483,N_9506);
and U9722 (N_9722,N_9512,N_9524);
and U9723 (N_9723,N_9469,N_9564);
nand U9724 (N_9724,N_9421,N_9431);
nand U9725 (N_9725,N_9447,N_9405);
or U9726 (N_9726,N_9456,N_9572);
or U9727 (N_9727,N_9472,N_9510);
or U9728 (N_9728,N_9475,N_9498);
or U9729 (N_9729,N_9546,N_9533);
nand U9730 (N_9730,N_9418,N_9578);
nor U9731 (N_9731,N_9455,N_9515);
nor U9732 (N_9732,N_9439,N_9407);
nor U9733 (N_9733,N_9545,N_9583);
nand U9734 (N_9734,N_9529,N_9443);
nor U9735 (N_9735,N_9502,N_9483);
nor U9736 (N_9736,N_9436,N_9448);
and U9737 (N_9737,N_9432,N_9422);
xnor U9738 (N_9738,N_9525,N_9428);
nand U9739 (N_9739,N_9474,N_9582);
or U9740 (N_9740,N_9415,N_9510);
nor U9741 (N_9741,N_9564,N_9411);
xor U9742 (N_9742,N_9583,N_9522);
nor U9743 (N_9743,N_9440,N_9569);
nand U9744 (N_9744,N_9451,N_9531);
xnor U9745 (N_9745,N_9531,N_9564);
xor U9746 (N_9746,N_9512,N_9427);
xor U9747 (N_9747,N_9405,N_9463);
nand U9748 (N_9748,N_9581,N_9571);
and U9749 (N_9749,N_9524,N_9461);
xor U9750 (N_9750,N_9470,N_9495);
nand U9751 (N_9751,N_9505,N_9455);
or U9752 (N_9752,N_9468,N_9446);
xnor U9753 (N_9753,N_9459,N_9532);
or U9754 (N_9754,N_9548,N_9590);
and U9755 (N_9755,N_9571,N_9556);
and U9756 (N_9756,N_9476,N_9403);
and U9757 (N_9757,N_9480,N_9550);
nand U9758 (N_9758,N_9492,N_9565);
nand U9759 (N_9759,N_9414,N_9436);
and U9760 (N_9760,N_9432,N_9524);
and U9761 (N_9761,N_9457,N_9488);
nor U9762 (N_9762,N_9498,N_9470);
nor U9763 (N_9763,N_9587,N_9510);
and U9764 (N_9764,N_9442,N_9546);
nor U9765 (N_9765,N_9414,N_9411);
and U9766 (N_9766,N_9401,N_9546);
or U9767 (N_9767,N_9574,N_9481);
and U9768 (N_9768,N_9575,N_9500);
nor U9769 (N_9769,N_9503,N_9523);
nand U9770 (N_9770,N_9455,N_9504);
xnor U9771 (N_9771,N_9581,N_9521);
xor U9772 (N_9772,N_9575,N_9437);
and U9773 (N_9773,N_9458,N_9508);
and U9774 (N_9774,N_9408,N_9578);
or U9775 (N_9775,N_9461,N_9427);
nor U9776 (N_9776,N_9567,N_9435);
xnor U9777 (N_9777,N_9423,N_9561);
or U9778 (N_9778,N_9454,N_9535);
and U9779 (N_9779,N_9464,N_9508);
nand U9780 (N_9780,N_9414,N_9549);
nand U9781 (N_9781,N_9444,N_9544);
nor U9782 (N_9782,N_9505,N_9500);
nor U9783 (N_9783,N_9561,N_9469);
and U9784 (N_9784,N_9480,N_9564);
or U9785 (N_9785,N_9482,N_9515);
nor U9786 (N_9786,N_9437,N_9483);
nand U9787 (N_9787,N_9416,N_9497);
or U9788 (N_9788,N_9448,N_9517);
xnor U9789 (N_9789,N_9414,N_9555);
or U9790 (N_9790,N_9526,N_9577);
xor U9791 (N_9791,N_9486,N_9434);
xnor U9792 (N_9792,N_9544,N_9472);
nand U9793 (N_9793,N_9484,N_9431);
xor U9794 (N_9794,N_9436,N_9519);
nor U9795 (N_9795,N_9545,N_9594);
nor U9796 (N_9796,N_9584,N_9592);
or U9797 (N_9797,N_9530,N_9450);
or U9798 (N_9798,N_9441,N_9426);
nand U9799 (N_9799,N_9437,N_9468);
nor U9800 (N_9800,N_9653,N_9796);
nand U9801 (N_9801,N_9618,N_9761);
or U9802 (N_9802,N_9671,N_9692);
nor U9803 (N_9803,N_9737,N_9745);
nor U9804 (N_9804,N_9783,N_9749);
nor U9805 (N_9805,N_9655,N_9756);
and U9806 (N_9806,N_9657,N_9685);
xor U9807 (N_9807,N_9677,N_9682);
and U9808 (N_9808,N_9781,N_9722);
nand U9809 (N_9809,N_9689,N_9673);
nor U9810 (N_9810,N_9617,N_9752);
nor U9811 (N_9811,N_9795,N_9674);
or U9812 (N_9812,N_9764,N_9770);
xnor U9813 (N_9813,N_9612,N_9747);
or U9814 (N_9814,N_9684,N_9630);
and U9815 (N_9815,N_9734,N_9777);
or U9816 (N_9816,N_9654,N_9710);
nor U9817 (N_9817,N_9751,N_9721);
nand U9818 (N_9818,N_9631,N_9714);
and U9819 (N_9819,N_9735,N_9759);
or U9820 (N_9820,N_9648,N_9715);
and U9821 (N_9821,N_9793,N_9750);
or U9822 (N_9822,N_9744,N_9627);
nand U9823 (N_9823,N_9628,N_9738);
and U9824 (N_9824,N_9665,N_9773);
and U9825 (N_9825,N_9691,N_9700);
nand U9826 (N_9826,N_9694,N_9603);
xnor U9827 (N_9827,N_9688,N_9767);
xnor U9828 (N_9828,N_9778,N_9669);
nor U9829 (N_9829,N_9789,N_9658);
and U9830 (N_9830,N_9664,N_9797);
nand U9831 (N_9831,N_9641,N_9794);
or U9832 (N_9832,N_9733,N_9642);
or U9833 (N_9833,N_9727,N_9718);
nor U9834 (N_9834,N_9629,N_9766);
nand U9835 (N_9835,N_9632,N_9662);
or U9836 (N_9836,N_9698,N_9765);
and U9837 (N_9837,N_9755,N_9625);
xnor U9838 (N_9838,N_9731,N_9670);
nand U9839 (N_9839,N_9711,N_9659);
and U9840 (N_9840,N_9637,N_9743);
nand U9841 (N_9841,N_9701,N_9678);
nand U9842 (N_9842,N_9696,N_9713);
or U9843 (N_9843,N_9712,N_9640);
xor U9844 (N_9844,N_9620,N_9788);
xnor U9845 (N_9845,N_9667,N_9616);
nor U9846 (N_9846,N_9697,N_9621);
and U9847 (N_9847,N_9719,N_9791);
nand U9848 (N_9848,N_9675,N_9754);
nand U9849 (N_9849,N_9619,N_9638);
or U9850 (N_9850,N_9650,N_9652);
xor U9851 (N_9851,N_9763,N_9699);
or U9852 (N_9852,N_9775,N_9720);
nand U9853 (N_9853,N_9646,N_9615);
xnor U9854 (N_9854,N_9706,N_9739);
nor U9855 (N_9855,N_9798,N_9626);
or U9856 (N_9856,N_9790,N_9774);
and U9857 (N_9857,N_9622,N_9786);
and U9858 (N_9858,N_9611,N_9708);
and U9859 (N_9859,N_9600,N_9610);
nand U9860 (N_9860,N_9676,N_9633);
nor U9861 (N_9861,N_9776,N_9787);
nand U9862 (N_9862,N_9746,N_9748);
nand U9863 (N_9863,N_9649,N_9680);
or U9864 (N_9864,N_9753,N_9799);
nand U9865 (N_9865,N_9782,N_9686);
and U9866 (N_9866,N_9607,N_9762);
and U9867 (N_9867,N_9608,N_9771);
nand U9868 (N_9868,N_9651,N_9703);
or U9869 (N_9869,N_9660,N_9726);
and U9870 (N_9870,N_9757,N_9644);
nand U9871 (N_9871,N_9687,N_9647);
or U9872 (N_9872,N_9602,N_9679);
nor U9873 (N_9873,N_9717,N_9732);
or U9874 (N_9874,N_9663,N_9709);
xor U9875 (N_9875,N_9690,N_9636);
and U9876 (N_9876,N_9639,N_9601);
xor U9877 (N_9877,N_9723,N_9695);
nor U9878 (N_9878,N_9736,N_9772);
nand U9879 (N_9879,N_9693,N_9728);
nor U9880 (N_9880,N_9742,N_9606);
xor U9881 (N_9881,N_9784,N_9704);
nand U9882 (N_9882,N_9741,N_9779);
nor U9883 (N_9883,N_9707,N_9716);
xnor U9884 (N_9884,N_9656,N_9792);
nor U9885 (N_9885,N_9635,N_9661);
and U9886 (N_9886,N_9724,N_9702);
nor U9887 (N_9887,N_9769,N_9683);
and U9888 (N_9888,N_9740,N_9725);
nor U9889 (N_9889,N_9681,N_9604);
and U9890 (N_9890,N_9760,N_9785);
xor U9891 (N_9891,N_9614,N_9729);
and U9892 (N_9892,N_9645,N_9623);
and U9893 (N_9893,N_9624,N_9780);
and U9894 (N_9894,N_9672,N_9730);
or U9895 (N_9895,N_9634,N_9613);
and U9896 (N_9896,N_9705,N_9668);
nand U9897 (N_9897,N_9768,N_9605);
xnor U9898 (N_9898,N_9758,N_9666);
nand U9899 (N_9899,N_9643,N_9609);
nand U9900 (N_9900,N_9700,N_9628);
nand U9901 (N_9901,N_9685,N_9696);
nor U9902 (N_9902,N_9772,N_9713);
or U9903 (N_9903,N_9755,N_9670);
xor U9904 (N_9904,N_9727,N_9782);
and U9905 (N_9905,N_9623,N_9705);
xor U9906 (N_9906,N_9780,N_9672);
and U9907 (N_9907,N_9719,N_9699);
xor U9908 (N_9908,N_9790,N_9634);
xnor U9909 (N_9909,N_9716,N_9709);
or U9910 (N_9910,N_9780,N_9617);
xnor U9911 (N_9911,N_9794,N_9602);
or U9912 (N_9912,N_9741,N_9697);
xnor U9913 (N_9913,N_9637,N_9645);
and U9914 (N_9914,N_9665,N_9743);
nand U9915 (N_9915,N_9731,N_9671);
nand U9916 (N_9916,N_9675,N_9657);
or U9917 (N_9917,N_9680,N_9759);
nor U9918 (N_9918,N_9748,N_9718);
and U9919 (N_9919,N_9625,N_9759);
nor U9920 (N_9920,N_9784,N_9657);
nor U9921 (N_9921,N_9657,N_9793);
or U9922 (N_9922,N_9600,N_9643);
nand U9923 (N_9923,N_9659,N_9649);
xnor U9924 (N_9924,N_9722,N_9741);
and U9925 (N_9925,N_9773,N_9721);
nor U9926 (N_9926,N_9604,N_9762);
nand U9927 (N_9927,N_9745,N_9631);
and U9928 (N_9928,N_9670,N_9794);
and U9929 (N_9929,N_9614,N_9646);
nor U9930 (N_9930,N_9764,N_9681);
nand U9931 (N_9931,N_9619,N_9710);
nand U9932 (N_9932,N_9656,N_9709);
or U9933 (N_9933,N_9799,N_9711);
and U9934 (N_9934,N_9683,N_9640);
nor U9935 (N_9935,N_9664,N_9621);
and U9936 (N_9936,N_9604,N_9650);
nor U9937 (N_9937,N_9685,N_9673);
nand U9938 (N_9938,N_9743,N_9705);
and U9939 (N_9939,N_9612,N_9614);
xnor U9940 (N_9940,N_9736,N_9755);
and U9941 (N_9941,N_9725,N_9762);
or U9942 (N_9942,N_9721,N_9698);
nor U9943 (N_9943,N_9695,N_9742);
nor U9944 (N_9944,N_9759,N_9622);
and U9945 (N_9945,N_9728,N_9765);
and U9946 (N_9946,N_9692,N_9786);
or U9947 (N_9947,N_9753,N_9681);
nand U9948 (N_9948,N_9618,N_9672);
nand U9949 (N_9949,N_9729,N_9675);
or U9950 (N_9950,N_9759,N_9756);
nand U9951 (N_9951,N_9660,N_9797);
xnor U9952 (N_9952,N_9655,N_9644);
nand U9953 (N_9953,N_9706,N_9781);
or U9954 (N_9954,N_9681,N_9631);
nor U9955 (N_9955,N_9608,N_9677);
nand U9956 (N_9956,N_9600,N_9609);
nor U9957 (N_9957,N_9732,N_9697);
or U9958 (N_9958,N_9692,N_9722);
nor U9959 (N_9959,N_9728,N_9789);
nand U9960 (N_9960,N_9752,N_9715);
xnor U9961 (N_9961,N_9709,N_9646);
and U9962 (N_9962,N_9702,N_9620);
nand U9963 (N_9963,N_9638,N_9794);
nor U9964 (N_9964,N_9793,N_9624);
xnor U9965 (N_9965,N_9631,N_9684);
nand U9966 (N_9966,N_9793,N_9716);
nand U9967 (N_9967,N_9617,N_9629);
nor U9968 (N_9968,N_9720,N_9602);
and U9969 (N_9969,N_9754,N_9681);
xnor U9970 (N_9970,N_9628,N_9720);
xor U9971 (N_9971,N_9745,N_9771);
or U9972 (N_9972,N_9644,N_9700);
and U9973 (N_9973,N_9695,N_9604);
or U9974 (N_9974,N_9663,N_9777);
xnor U9975 (N_9975,N_9703,N_9627);
nand U9976 (N_9976,N_9729,N_9703);
xnor U9977 (N_9977,N_9635,N_9756);
nor U9978 (N_9978,N_9691,N_9751);
and U9979 (N_9979,N_9691,N_9759);
nand U9980 (N_9980,N_9600,N_9680);
or U9981 (N_9981,N_9662,N_9770);
or U9982 (N_9982,N_9612,N_9746);
nand U9983 (N_9983,N_9617,N_9636);
and U9984 (N_9984,N_9628,N_9609);
or U9985 (N_9985,N_9614,N_9763);
and U9986 (N_9986,N_9696,N_9755);
nor U9987 (N_9987,N_9760,N_9652);
nand U9988 (N_9988,N_9658,N_9627);
and U9989 (N_9989,N_9621,N_9754);
or U9990 (N_9990,N_9710,N_9615);
nand U9991 (N_9991,N_9667,N_9796);
or U9992 (N_9992,N_9605,N_9627);
nand U9993 (N_9993,N_9635,N_9649);
xnor U9994 (N_9994,N_9618,N_9762);
and U9995 (N_9995,N_9744,N_9686);
xnor U9996 (N_9996,N_9610,N_9687);
and U9997 (N_9997,N_9703,N_9767);
nand U9998 (N_9998,N_9667,N_9651);
nor U9999 (N_9999,N_9682,N_9722);
xnor U10000 (N_10000,N_9951,N_9832);
and U10001 (N_10001,N_9812,N_9807);
or U10002 (N_10002,N_9937,N_9920);
nor U10003 (N_10003,N_9903,N_9908);
xor U10004 (N_10004,N_9823,N_9995);
or U10005 (N_10005,N_9929,N_9916);
xor U10006 (N_10006,N_9860,N_9848);
nor U10007 (N_10007,N_9969,N_9905);
nand U10008 (N_10008,N_9983,N_9829);
nand U10009 (N_10009,N_9888,N_9869);
xor U10010 (N_10010,N_9846,N_9843);
xnor U10011 (N_10011,N_9965,N_9982);
nand U10012 (N_10012,N_9894,N_9868);
and U10013 (N_10013,N_9815,N_9874);
nand U10014 (N_10014,N_9956,N_9914);
xnor U10015 (N_10015,N_9990,N_9886);
xor U10016 (N_10016,N_9981,N_9917);
nor U10017 (N_10017,N_9810,N_9871);
xor U10018 (N_10018,N_9882,N_9827);
xnor U10019 (N_10019,N_9831,N_9986);
and U10020 (N_10020,N_9800,N_9849);
or U10021 (N_10021,N_9936,N_9852);
or U10022 (N_10022,N_9850,N_9893);
nand U10023 (N_10023,N_9892,N_9944);
or U10024 (N_10024,N_9862,N_9952);
xor U10025 (N_10025,N_9875,N_9977);
or U10026 (N_10026,N_9974,N_9996);
xnor U10027 (N_10027,N_9992,N_9988);
xor U10028 (N_10028,N_9961,N_9873);
xor U10029 (N_10029,N_9805,N_9941);
nor U10030 (N_10030,N_9939,N_9863);
nor U10031 (N_10031,N_9925,N_9821);
and U10032 (N_10032,N_9809,N_9844);
xnor U10033 (N_10033,N_9975,N_9879);
and U10034 (N_10034,N_9858,N_9979);
xnor U10035 (N_10035,N_9887,N_9891);
nand U10036 (N_10036,N_9976,N_9930);
xnor U10037 (N_10037,N_9987,N_9942);
or U10038 (N_10038,N_9839,N_9813);
and U10039 (N_10039,N_9907,N_9998);
nor U10040 (N_10040,N_9880,N_9932);
nor U10041 (N_10041,N_9803,N_9993);
nor U10042 (N_10042,N_9808,N_9816);
or U10043 (N_10043,N_9881,N_9851);
xnor U10044 (N_10044,N_9898,N_9943);
nor U10045 (N_10045,N_9968,N_9811);
xnor U10046 (N_10046,N_9924,N_9854);
nand U10047 (N_10047,N_9949,N_9984);
nor U10048 (N_10048,N_9994,N_9927);
nand U10049 (N_10049,N_9955,N_9902);
or U10050 (N_10050,N_9847,N_9818);
nor U10051 (N_10051,N_9856,N_9814);
nand U10052 (N_10052,N_9897,N_9820);
or U10053 (N_10053,N_9973,N_9940);
nand U10054 (N_10054,N_9928,N_9801);
xor U10055 (N_10055,N_9910,N_9890);
and U10056 (N_10056,N_9855,N_9953);
nor U10057 (N_10057,N_9950,N_9835);
or U10058 (N_10058,N_9954,N_9833);
nand U10059 (N_10059,N_9918,N_9980);
nor U10060 (N_10060,N_9933,N_9967);
or U10061 (N_10061,N_9870,N_9876);
and U10062 (N_10062,N_9828,N_9997);
xor U10063 (N_10063,N_9958,N_9913);
nor U10064 (N_10064,N_9957,N_9853);
or U10065 (N_10065,N_9819,N_9904);
xor U10066 (N_10066,N_9841,N_9945);
xor U10067 (N_10067,N_9878,N_9883);
nor U10068 (N_10068,N_9836,N_9865);
nand U10069 (N_10069,N_9861,N_9838);
and U10070 (N_10070,N_9921,N_9830);
xor U10071 (N_10071,N_9926,N_9912);
or U10072 (N_10072,N_9989,N_9962);
nor U10073 (N_10073,N_9889,N_9806);
nor U10074 (N_10074,N_9971,N_9872);
and U10075 (N_10075,N_9947,N_9959);
nor U10076 (N_10076,N_9946,N_9964);
nor U10077 (N_10077,N_9931,N_9885);
nand U10078 (N_10078,N_9970,N_9804);
xnor U10079 (N_10079,N_9859,N_9867);
nor U10080 (N_10080,N_9906,N_9909);
or U10081 (N_10081,N_9985,N_9923);
and U10082 (N_10082,N_9837,N_9948);
nor U10083 (N_10083,N_9922,N_9817);
or U10084 (N_10084,N_9960,N_9900);
and U10085 (N_10085,N_9866,N_9919);
xor U10086 (N_10086,N_9845,N_9895);
xnor U10087 (N_10087,N_9935,N_9915);
xnor U10088 (N_10088,N_9824,N_9899);
or U10089 (N_10089,N_9864,N_9825);
nand U10090 (N_10090,N_9857,N_9911);
nor U10091 (N_10091,N_9822,N_9877);
nor U10092 (N_10092,N_9842,N_9901);
and U10093 (N_10093,N_9963,N_9826);
nand U10094 (N_10094,N_9834,N_9934);
nor U10095 (N_10095,N_9991,N_9884);
xor U10096 (N_10096,N_9938,N_9840);
nor U10097 (N_10097,N_9978,N_9966);
or U10098 (N_10098,N_9896,N_9972);
or U10099 (N_10099,N_9999,N_9802);
xor U10100 (N_10100,N_9958,N_9902);
nor U10101 (N_10101,N_9911,N_9960);
or U10102 (N_10102,N_9808,N_9954);
or U10103 (N_10103,N_9819,N_9961);
nand U10104 (N_10104,N_9968,N_9994);
and U10105 (N_10105,N_9808,N_9926);
and U10106 (N_10106,N_9816,N_9856);
and U10107 (N_10107,N_9940,N_9963);
nor U10108 (N_10108,N_9991,N_9895);
and U10109 (N_10109,N_9918,N_9860);
xor U10110 (N_10110,N_9905,N_9874);
or U10111 (N_10111,N_9893,N_9830);
nor U10112 (N_10112,N_9938,N_9894);
nor U10113 (N_10113,N_9833,N_9936);
or U10114 (N_10114,N_9992,N_9814);
and U10115 (N_10115,N_9992,N_9804);
nand U10116 (N_10116,N_9923,N_9860);
or U10117 (N_10117,N_9974,N_9819);
or U10118 (N_10118,N_9897,N_9810);
and U10119 (N_10119,N_9899,N_9852);
nor U10120 (N_10120,N_9983,N_9827);
nand U10121 (N_10121,N_9851,N_9819);
xnor U10122 (N_10122,N_9802,N_9983);
nor U10123 (N_10123,N_9990,N_9864);
or U10124 (N_10124,N_9898,N_9867);
nand U10125 (N_10125,N_9978,N_9861);
nand U10126 (N_10126,N_9813,N_9881);
or U10127 (N_10127,N_9920,N_9908);
xnor U10128 (N_10128,N_9956,N_9951);
or U10129 (N_10129,N_9838,N_9869);
nand U10130 (N_10130,N_9912,N_9805);
xor U10131 (N_10131,N_9871,N_9977);
nor U10132 (N_10132,N_9871,N_9812);
and U10133 (N_10133,N_9915,N_9872);
nand U10134 (N_10134,N_9919,N_9918);
and U10135 (N_10135,N_9906,N_9925);
nand U10136 (N_10136,N_9835,N_9986);
nor U10137 (N_10137,N_9840,N_9875);
and U10138 (N_10138,N_9993,N_9968);
xnor U10139 (N_10139,N_9827,N_9837);
xor U10140 (N_10140,N_9820,N_9855);
or U10141 (N_10141,N_9963,N_9930);
xnor U10142 (N_10142,N_9831,N_9801);
and U10143 (N_10143,N_9978,N_9972);
nor U10144 (N_10144,N_9895,N_9928);
xnor U10145 (N_10145,N_9907,N_9942);
nor U10146 (N_10146,N_9949,N_9808);
xnor U10147 (N_10147,N_9946,N_9825);
or U10148 (N_10148,N_9905,N_9955);
nand U10149 (N_10149,N_9930,N_9874);
and U10150 (N_10150,N_9825,N_9920);
nor U10151 (N_10151,N_9997,N_9878);
nand U10152 (N_10152,N_9999,N_9922);
nor U10153 (N_10153,N_9867,N_9945);
nor U10154 (N_10154,N_9904,N_9887);
or U10155 (N_10155,N_9995,N_9942);
nor U10156 (N_10156,N_9986,N_9846);
nor U10157 (N_10157,N_9888,N_9816);
nand U10158 (N_10158,N_9977,N_9886);
or U10159 (N_10159,N_9803,N_9849);
or U10160 (N_10160,N_9836,N_9980);
or U10161 (N_10161,N_9991,N_9818);
or U10162 (N_10162,N_9938,N_9807);
nor U10163 (N_10163,N_9885,N_9982);
xor U10164 (N_10164,N_9839,N_9887);
nand U10165 (N_10165,N_9895,N_9880);
and U10166 (N_10166,N_9910,N_9883);
nor U10167 (N_10167,N_9918,N_9926);
or U10168 (N_10168,N_9988,N_9880);
xor U10169 (N_10169,N_9955,N_9971);
xor U10170 (N_10170,N_9841,N_9974);
and U10171 (N_10171,N_9808,N_9838);
and U10172 (N_10172,N_9893,N_9997);
nand U10173 (N_10173,N_9915,N_9941);
xnor U10174 (N_10174,N_9902,N_9982);
nor U10175 (N_10175,N_9857,N_9854);
nand U10176 (N_10176,N_9819,N_9945);
and U10177 (N_10177,N_9805,N_9896);
xnor U10178 (N_10178,N_9937,N_9803);
and U10179 (N_10179,N_9951,N_9998);
xor U10180 (N_10180,N_9855,N_9932);
nor U10181 (N_10181,N_9934,N_9933);
nand U10182 (N_10182,N_9983,N_9864);
and U10183 (N_10183,N_9954,N_9905);
and U10184 (N_10184,N_9881,N_9945);
or U10185 (N_10185,N_9866,N_9898);
nand U10186 (N_10186,N_9848,N_9889);
nor U10187 (N_10187,N_9964,N_9979);
nand U10188 (N_10188,N_9804,N_9848);
and U10189 (N_10189,N_9936,N_9828);
nor U10190 (N_10190,N_9995,N_9814);
or U10191 (N_10191,N_9959,N_9830);
nand U10192 (N_10192,N_9948,N_9899);
nand U10193 (N_10193,N_9913,N_9845);
and U10194 (N_10194,N_9871,N_9933);
or U10195 (N_10195,N_9969,N_9888);
or U10196 (N_10196,N_9882,N_9862);
or U10197 (N_10197,N_9907,N_9912);
xor U10198 (N_10198,N_9902,N_9893);
nor U10199 (N_10199,N_9824,N_9818);
and U10200 (N_10200,N_10145,N_10185);
nand U10201 (N_10201,N_10127,N_10189);
or U10202 (N_10202,N_10161,N_10162);
or U10203 (N_10203,N_10053,N_10181);
or U10204 (N_10204,N_10019,N_10095);
and U10205 (N_10205,N_10134,N_10013);
nand U10206 (N_10206,N_10198,N_10186);
nand U10207 (N_10207,N_10111,N_10089);
nor U10208 (N_10208,N_10141,N_10098);
xnor U10209 (N_10209,N_10178,N_10085);
xor U10210 (N_10210,N_10149,N_10122);
and U10211 (N_10211,N_10135,N_10124);
nor U10212 (N_10212,N_10087,N_10103);
and U10213 (N_10213,N_10064,N_10176);
nor U10214 (N_10214,N_10160,N_10070);
nand U10215 (N_10215,N_10068,N_10012);
xor U10216 (N_10216,N_10180,N_10056);
xor U10217 (N_10217,N_10038,N_10071);
or U10218 (N_10218,N_10049,N_10173);
or U10219 (N_10219,N_10061,N_10036);
and U10220 (N_10220,N_10073,N_10129);
and U10221 (N_10221,N_10104,N_10072);
and U10222 (N_10222,N_10051,N_10066);
nor U10223 (N_10223,N_10065,N_10022);
xor U10224 (N_10224,N_10188,N_10110);
and U10225 (N_10225,N_10034,N_10037);
or U10226 (N_10226,N_10083,N_10184);
nand U10227 (N_10227,N_10004,N_10168);
nand U10228 (N_10228,N_10047,N_10005);
and U10229 (N_10229,N_10133,N_10120);
and U10230 (N_10230,N_10170,N_10128);
nor U10231 (N_10231,N_10026,N_10076);
and U10232 (N_10232,N_10190,N_10101);
and U10233 (N_10233,N_10165,N_10094);
xor U10234 (N_10234,N_10194,N_10041);
nor U10235 (N_10235,N_10016,N_10107);
and U10236 (N_10236,N_10154,N_10179);
and U10237 (N_10237,N_10130,N_10069);
or U10238 (N_10238,N_10132,N_10057);
nor U10239 (N_10239,N_10100,N_10027);
nor U10240 (N_10240,N_10082,N_10075);
and U10241 (N_10241,N_10096,N_10192);
nor U10242 (N_10242,N_10153,N_10163);
nand U10243 (N_10243,N_10108,N_10003);
and U10244 (N_10244,N_10114,N_10102);
or U10245 (N_10245,N_10099,N_10055);
or U10246 (N_10246,N_10164,N_10024);
nor U10247 (N_10247,N_10028,N_10147);
nand U10248 (N_10248,N_10182,N_10140);
and U10249 (N_10249,N_10007,N_10001);
xnor U10250 (N_10250,N_10009,N_10126);
nor U10251 (N_10251,N_10044,N_10115);
xnor U10252 (N_10252,N_10052,N_10000);
nor U10253 (N_10253,N_10172,N_10146);
nor U10254 (N_10254,N_10008,N_10105);
xnor U10255 (N_10255,N_10020,N_10035);
and U10256 (N_10256,N_10029,N_10112);
nand U10257 (N_10257,N_10050,N_10091);
nor U10258 (N_10258,N_10086,N_10011);
and U10259 (N_10259,N_10117,N_10199);
nor U10260 (N_10260,N_10157,N_10155);
nor U10261 (N_10261,N_10023,N_10006);
or U10262 (N_10262,N_10002,N_10018);
nand U10263 (N_10263,N_10142,N_10097);
and U10264 (N_10264,N_10040,N_10088);
or U10265 (N_10265,N_10197,N_10067);
or U10266 (N_10266,N_10166,N_10191);
xnor U10267 (N_10267,N_10169,N_10109);
or U10268 (N_10268,N_10148,N_10042);
or U10269 (N_10269,N_10046,N_10017);
and U10270 (N_10270,N_10113,N_10062);
and U10271 (N_10271,N_10144,N_10021);
nand U10272 (N_10272,N_10090,N_10048);
nand U10273 (N_10273,N_10093,N_10063);
nor U10274 (N_10274,N_10195,N_10060);
xnor U10275 (N_10275,N_10152,N_10137);
nor U10276 (N_10276,N_10014,N_10084);
nand U10277 (N_10277,N_10151,N_10119);
xnor U10278 (N_10278,N_10159,N_10118);
xor U10279 (N_10279,N_10167,N_10031);
nand U10280 (N_10280,N_10080,N_10074);
xnor U10281 (N_10281,N_10106,N_10032);
nor U10282 (N_10282,N_10092,N_10079);
or U10283 (N_10283,N_10078,N_10136);
or U10284 (N_10284,N_10077,N_10183);
and U10285 (N_10285,N_10131,N_10139);
nand U10286 (N_10286,N_10054,N_10138);
nand U10287 (N_10287,N_10174,N_10059);
xnor U10288 (N_10288,N_10045,N_10039);
or U10289 (N_10289,N_10175,N_10123);
xnor U10290 (N_10290,N_10025,N_10158);
or U10291 (N_10291,N_10125,N_10015);
and U10292 (N_10292,N_10150,N_10143);
and U10293 (N_10293,N_10081,N_10010);
or U10294 (N_10294,N_10171,N_10156);
nor U10295 (N_10295,N_10196,N_10058);
xnor U10296 (N_10296,N_10187,N_10177);
nor U10297 (N_10297,N_10043,N_10033);
and U10298 (N_10298,N_10116,N_10030);
xnor U10299 (N_10299,N_10193,N_10121);
or U10300 (N_10300,N_10139,N_10120);
and U10301 (N_10301,N_10065,N_10063);
or U10302 (N_10302,N_10176,N_10150);
nand U10303 (N_10303,N_10156,N_10021);
nor U10304 (N_10304,N_10083,N_10065);
nor U10305 (N_10305,N_10009,N_10190);
xnor U10306 (N_10306,N_10178,N_10158);
xnor U10307 (N_10307,N_10082,N_10137);
nand U10308 (N_10308,N_10184,N_10079);
or U10309 (N_10309,N_10023,N_10198);
xor U10310 (N_10310,N_10156,N_10143);
and U10311 (N_10311,N_10055,N_10142);
xnor U10312 (N_10312,N_10195,N_10067);
nand U10313 (N_10313,N_10125,N_10159);
xnor U10314 (N_10314,N_10098,N_10140);
nor U10315 (N_10315,N_10058,N_10091);
nor U10316 (N_10316,N_10049,N_10129);
xor U10317 (N_10317,N_10139,N_10146);
nand U10318 (N_10318,N_10109,N_10129);
or U10319 (N_10319,N_10151,N_10199);
xnor U10320 (N_10320,N_10161,N_10130);
and U10321 (N_10321,N_10134,N_10117);
nor U10322 (N_10322,N_10106,N_10150);
or U10323 (N_10323,N_10055,N_10038);
nand U10324 (N_10324,N_10154,N_10131);
nor U10325 (N_10325,N_10020,N_10060);
nor U10326 (N_10326,N_10008,N_10130);
xnor U10327 (N_10327,N_10025,N_10055);
or U10328 (N_10328,N_10141,N_10081);
and U10329 (N_10329,N_10162,N_10105);
nand U10330 (N_10330,N_10029,N_10065);
xor U10331 (N_10331,N_10022,N_10009);
nor U10332 (N_10332,N_10066,N_10022);
or U10333 (N_10333,N_10095,N_10143);
or U10334 (N_10334,N_10147,N_10176);
nor U10335 (N_10335,N_10191,N_10189);
xnor U10336 (N_10336,N_10148,N_10194);
and U10337 (N_10337,N_10101,N_10154);
nor U10338 (N_10338,N_10156,N_10141);
nor U10339 (N_10339,N_10144,N_10176);
nor U10340 (N_10340,N_10008,N_10090);
and U10341 (N_10341,N_10050,N_10142);
or U10342 (N_10342,N_10154,N_10199);
nor U10343 (N_10343,N_10061,N_10002);
or U10344 (N_10344,N_10100,N_10054);
nand U10345 (N_10345,N_10144,N_10024);
and U10346 (N_10346,N_10090,N_10026);
or U10347 (N_10347,N_10139,N_10115);
nor U10348 (N_10348,N_10193,N_10156);
nor U10349 (N_10349,N_10150,N_10188);
nand U10350 (N_10350,N_10171,N_10012);
or U10351 (N_10351,N_10006,N_10070);
and U10352 (N_10352,N_10117,N_10047);
and U10353 (N_10353,N_10182,N_10086);
or U10354 (N_10354,N_10172,N_10177);
nand U10355 (N_10355,N_10031,N_10075);
nor U10356 (N_10356,N_10071,N_10006);
nand U10357 (N_10357,N_10024,N_10036);
nor U10358 (N_10358,N_10090,N_10020);
xnor U10359 (N_10359,N_10025,N_10195);
and U10360 (N_10360,N_10087,N_10153);
xnor U10361 (N_10361,N_10037,N_10029);
or U10362 (N_10362,N_10011,N_10091);
or U10363 (N_10363,N_10140,N_10176);
and U10364 (N_10364,N_10061,N_10137);
or U10365 (N_10365,N_10168,N_10187);
nor U10366 (N_10366,N_10059,N_10191);
nand U10367 (N_10367,N_10198,N_10180);
xnor U10368 (N_10368,N_10177,N_10179);
xor U10369 (N_10369,N_10100,N_10197);
and U10370 (N_10370,N_10040,N_10119);
or U10371 (N_10371,N_10076,N_10066);
and U10372 (N_10372,N_10159,N_10187);
or U10373 (N_10373,N_10099,N_10087);
nor U10374 (N_10374,N_10168,N_10147);
or U10375 (N_10375,N_10010,N_10018);
nand U10376 (N_10376,N_10102,N_10041);
nor U10377 (N_10377,N_10001,N_10174);
xor U10378 (N_10378,N_10086,N_10166);
xnor U10379 (N_10379,N_10079,N_10112);
nand U10380 (N_10380,N_10085,N_10055);
and U10381 (N_10381,N_10082,N_10038);
or U10382 (N_10382,N_10068,N_10114);
nor U10383 (N_10383,N_10156,N_10187);
or U10384 (N_10384,N_10113,N_10083);
xnor U10385 (N_10385,N_10043,N_10002);
nand U10386 (N_10386,N_10118,N_10027);
nor U10387 (N_10387,N_10115,N_10129);
nand U10388 (N_10388,N_10138,N_10090);
nand U10389 (N_10389,N_10073,N_10053);
or U10390 (N_10390,N_10085,N_10028);
xnor U10391 (N_10391,N_10072,N_10138);
and U10392 (N_10392,N_10101,N_10084);
and U10393 (N_10393,N_10197,N_10080);
or U10394 (N_10394,N_10001,N_10114);
nor U10395 (N_10395,N_10100,N_10084);
and U10396 (N_10396,N_10183,N_10173);
nor U10397 (N_10397,N_10198,N_10181);
nand U10398 (N_10398,N_10112,N_10118);
or U10399 (N_10399,N_10127,N_10136);
nand U10400 (N_10400,N_10361,N_10310);
nand U10401 (N_10401,N_10386,N_10237);
nor U10402 (N_10402,N_10352,N_10294);
and U10403 (N_10403,N_10394,N_10288);
or U10404 (N_10404,N_10322,N_10220);
nor U10405 (N_10405,N_10324,N_10295);
or U10406 (N_10406,N_10258,N_10279);
or U10407 (N_10407,N_10216,N_10362);
nand U10408 (N_10408,N_10387,N_10293);
xor U10409 (N_10409,N_10321,N_10340);
nand U10410 (N_10410,N_10378,N_10360);
xor U10411 (N_10411,N_10350,N_10359);
xor U10412 (N_10412,N_10357,N_10229);
nand U10413 (N_10413,N_10219,N_10239);
nor U10414 (N_10414,N_10243,N_10327);
nor U10415 (N_10415,N_10210,N_10349);
or U10416 (N_10416,N_10286,N_10365);
nand U10417 (N_10417,N_10308,N_10265);
and U10418 (N_10418,N_10371,N_10254);
xnor U10419 (N_10419,N_10341,N_10381);
nor U10420 (N_10420,N_10261,N_10235);
nor U10421 (N_10421,N_10301,N_10224);
or U10422 (N_10422,N_10347,N_10372);
nand U10423 (N_10423,N_10226,N_10328);
and U10424 (N_10424,N_10373,N_10281);
xor U10425 (N_10425,N_10251,N_10259);
or U10426 (N_10426,N_10344,N_10364);
or U10427 (N_10427,N_10398,N_10233);
nand U10428 (N_10428,N_10214,N_10306);
xor U10429 (N_10429,N_10366,N_10255);
nand U10430 (N_10430,N_10207,N_10345);
and U10431 (N_10431,N_10354,N_10309);
nor U10432 (N_10432,N_10331,N_10267);
or U10433 (N_10433,N_10223,N_10213);
nor U10434 (N_10434,N_10316,N_10273);
nand U10435 (N_10435,N_10377,N_10333);
xor U10436 (N_10436,N_10289,N_10257);
nand U10437 (N_10437,N_10329,N_10247);
xor U10438 (N_10438,N_10291,N_10218);
nor U10439 (N_10439,N_10205,N_10278);
and U10440 (N_10440,N_10319,N_10264);
xnor U10441 (N_10441,N_10379,N_10248);
nor U10442 (N_10442,N_10249,N_10225);
or U10443 (N_10443,N_10270,N_10245);
nor U10444 (N_10444,N_10363,N_10388);
nand U10445 (N_10445,N_10274,N_10397);
or U10446 (N_10446,N_10358,N_10266);
or U10447 (N_10447,N_10238,N_10228);
xor U10448 (N_10448,N_10221,N_10368);
and U10449 (N_10449,N_10339,N_10314);
nor U10450 (N_10450,N_10334,N_10298);
and U10451 (N_10451,N_10302,N_10353);
and U10452 (N_10452,N_10337,N_10382);
xnor U10453 (N_10453,N_10280,N_10338);
and U10454 (N_10454,N_10299,N_10241);
xnor U10455 (N_10455,N_10209,N_10282);
and U10456 (N_10456,N_10263,N_10304);
xor U10457 (N_10457,N_10385,N_10287);
and U10458 (N_10458,N_10305,N_10203);
nor U10459 (N_10459,N_10312,N_10351);
or U10460 (N_10460,N_10384,N_10318);
nor U10461 (N_10461,N_10330,N_10202);
xor U10462 (N_10462,N_10200,N_10391);
or U10463 (N_10463,N_10284,N_10244);
nand U10464 (N_10464,N_10242,N_10315);
nand U10465 (N_10465,N_10380,N_10271);
nand U10466 (N_10466,N_10201,N_10283);
or U10467 (N_10467,N_10311,N_10300);
or U10468 (N_10468,N_10393,N_10375);
or U10469 (N_10469,N_10246,N_10206);
or U10470 (N_10470,N_10260,N_10275);
xor U10471 (N_10471,N_10313,N_10332);
and U10472 (N_10472,N_10323,N_10383);
xor U10473 (N_10473,N_10290,N_10204);
nor U10474 (N_10474,N_10296,N_10253);
or U10475 (N_10475,N_10272,N_10231);
nor U10476 (N_10476,N_10303,N_10399);
or U10477 (N_10477,N_10369,N_10232);
nor U10478 (N_10478,N_10292,N_10262);
and U10479 (N_10479,N_10252,N_10269);
and U10480 (N_10480,N_10256,N_10367);
nor U10481 (N_10481,N_10395,N_10374);
or U10482 (N_10482,N_10240,N_10277);
xnor U10483 (N_10483,N_10285,N_10227);
nand U10484 (N_10484,N_10396,N_10335);
nor U10485 (N_10485,N_10234,N_10307);
nor U10486 (N_10486,N_10336,N_10376);
and U10487 (N_10487,N_10208,N_10236);
or U10488 (N_10488,N_10268,N_10217);
and U10489 (N_10489,N_10276,N_10348);
or U10490 (N_10490,N_10389,N_10317);
nand U10491 (N_10491,N_10370,N_10356);
or U10492 (N_10492,N_10326,N_10325);
nand U10493 (N_10493,N_10215,N_10250);
or U10494 (N_10494,N_10320,N_10390);
nand U10495 (N_10495,N_10392,N_10230);
nor U10496 (N_10496,N_10222,N_10211);
or U10497 (N_10497,N_10343,N_10342);
and U10498 (N_10498,N_10355,N_10346);
and U10499 (N_10499,N_10297,N_10212);
nand U10500 (N_10500,N_10286,N_10363);
nand U10501 (N_10501,N_10270,N_10308);
or U10502 (N_10502,N_10395,N_10259);
or U10503 (N_10503,N_10346,N_10273);
or U10504 (N_10504,N_10329,N_10345);
nor U10505 (N_10505,N_10385,N_10331);
and U10506 (N_10506,N_10394,N_10363);
xor U10507 (N_10507,N_10213,N_10328);
nor U10508 (N_10508,N_10396,N_10219);
or U10509 (N_10509,N_10223,N_10383);
nor U10510 (N_10510,N_10367,N_10363);
nor U10511 (N_10511,N_10333,N_10382);
and U10512 (N_10512,N_10399,N_10280);
nor U10513 (N_10513,N_10302,N_10206);
or U10514 (N_10514,N_10247,N_10377);
and U10515 (N_10515,N_10339,N_10297);
nor U10516 (N_10516,N_10391,N_10274);
nor U10517 (N_10517,N_10258,N_10368);
nand U10518 (N_10518,N_10313,N_10212);
and U10519 (N_10519,N_10300,N_10259);
xor U10520 (N_10520,N_10229,N_10288);
nand U10521 (N_10521,N_10204,N_10286);
nand U10522 (N_10522,N_10387,N_10322);
or U10523 (N_10523,N_10240,N_10296);
nand U10524 (N_10524,N_10351,N_10237);
or U10525 (N_10525,N_10287,N_10363);
nor U10526 (N_10526,N_10305,N_10368);
xor U10527 (N_10527,N_10304,N_10323);
and U10528 (N_10528,N_10278,N_10247);
xor U10529 (N_10529,N_10385,N_10333);
or U10530 (N_10530,N_10275,N_10279);
nand U10531 (N_10531,N_10306,N_10266);
nand U10532 (N_10532,N_10272,N_10310);
and U10533 (N_10533,N_10206,N_10320);
nand U10534 (N_10534,N_10264,N_10204);
or U10535 (N_10535,N_10395,N_10203);
nand U10536 (N_10536,N_10321,N_10302);
or U10537 (N_10537,N_10278,N_10396);
nand U10538 (N_10538,N_10294,N_10345);
and U10539 (N_10539,N_10397,N_10349);
nor U10540 (N_10540,N_10304,N_10367);
xnor U10541 (N_10541,N_10360,N_10257);
xor U10542 (N_10542,N_10247,N_10238);
and U10543 (N_10543,N_10311,N_10315);
nand U10544 (N_10544,N_10398,N_10283);
or U10545 (N_10545,N_10310,N_10398);
or U10546 (N_10546,N_10359,N_10314);
and U10547 (N_10547,N_10225,N_10348);
or U10548 (N_10548,N_10231,N_10299);
nand U10549 (N_10549,N_10220,N_10218);
xnor U10550 (N_10550,N_10292,N_10354);
and U10551 (N_10551,N_10248,N_10314);
or U10552 (N_10552,N_10300,N_10268);
xor U10553 (N_10553,N_10220,N_10260);
nand U10554 (N_10554,N_10372,N_10326);
or U10555 (N_10555,N_10367,N_10396);
and U10556 (N_10556,N_10298,N_10280);
and U10557 (N_10557,N_10352,N_10379);
nand U10558 (N_10558,N_10230,N_10389);
xnor U10559 (N_10559,N_10233,N_10397);
or U10560 (N_10560,N_10235,N_10300);
nor U10561 (N_10561,N_10283,N_10232);
nor U10562 (N_10562,N_10258,N_10242);
and U10563 (N_10563,N_10336,N_10214);
nand U10564 (N_10564,N_10384,N_10387);
or U10565 (N_10565,N_10223,N_10271);
and U10566 (N_10566,N_10299,N_10283);
or U10567 (N_10567,N_10266,N_10350);
xnor U10568 (N_10568,N_10371,N_10352);
nor U10569 (N_10569,N_10297,N_10285);
nor U10570 (N_10570,N_10347,N_10202);
or U10571 (N_10571,N_10241,N_10353);
nor U10572 (N_10572,N_10306,N_10396);
nand U10573 (N_10573,N_10218,N_10381);
xnor U10574 (N_10574,N_10395,N_10218);
or U10575 (N_10575,N_10262,N_10291);
xnor U10576 (N_10576,N_10340,N_10374);
xor U10577 (N_10577,N_10334,N_10297);
and U10578 (N_10578,N_10340,N_10203);
nor U10579 (N_10579,N_10277,N_10365);
nor U10580 (N_10580,N_10354,N_10320);
or U10581 (N_10581,N_10344,N_10228);
xnor U10582 (N_10582,N_10284,N_10382);
and U10583 (N_10583,N_10254,N_10206);
or U10584 (N_10584,N_10265,N_10304);
nor U10585 (N_10585,N_10396,N_10263);
nand U10586 (N_10586,N_10276,N_10210);
xor U10587 (N_10587,N_10200,N_10360);
nor U10588 (N_10588,N_10257,N_10214);
and U10589 (N_10589,N_10280,N_10271);
xor U10590 (N_10590,N_10203,N_10233);
xnor U10591 (N_10591,N_10344,N_10318);
or U10592 (N_10592,N_10235,N_10395);
xnor U10593 (N_10593,N_10214,N_10363);
nor U10594 (N_10594,N_10350,N_10267);
nor U10595 (N_10595,N_10208,N_10316);
nor U10596 (N_10596,N_10306,N_10391);
or U10597 (N_10597,N_10293,N_10365);
nor U10598 (N_10598,N_10295,N_10397);
or U10599 (N_10599,N_10313,N_10375);
and U10600 (N_10600,N_10598,N_10515);
or U10601 (N_10601,N_10562,N_10535);
or U10602 (N_10602,N_10537,N_10549);
or U10603 (N_10603,N_10577,N_10468);
nand U10604 (N_10604,N_10529,N_10405);
or U10605 (N_10605,N_10566,N_10472);
or U10606 (N_10606,N_10439,N_10493);
nor U10607 (N_10607,N_10499,N_10442);
xnor U10608 (N_10608,N_10553,N_10411);
nor U10609 (N_10609,N_10555,N_10464);
xnor U10610 (N_10610,N_10526,N_10436);
nor U10611 (N_10611,N_10423,N_10528);
xnor U10612 (N_10612,N_10561,N_10434);
nor U10613 (N_10613,N_10587,N_10443);
xnor U10614 (N_10614,N_10534,N_10597);
or U10615 (N_10615,N_10498,N_10510);
xnor U10616 (N_10616,N_10487,N_10572);
or U10617 (N_10617,N_10560,N_10418);
or U10618 (N_10618,N_10410,N_10412);
or U10619 (N_10619,N_10455,N_10491);
xnor U10620 (N_10620,N_10582,N_10429);
or U10621 (N_10621,N_10589,N_10478);
nor U10622 (N_10622,N_10511,N_10565);
and U10623 (N_10623,N_10540,N_10452);
or U10624 (N_10624,N_10596,N_10538);
and U10625 (N_10625,N_10557,N_10466);
or U10626 (N_10626,N_10520,N_10407);
xnor U10627 (N_10627,N_10408,N_10471);
or U10628 (N_10628,N_10521,N_10579);
nand U10629 (N_10629,N_10469,N_10531);
nand U10630 (N_10630,N_10420,N_10430);
nor U10631 (N_10631,N_10554,N_10522);
nor U10632 (N_10632,N_10482,N_10433);
nand U10633 (N_10633,N_10451,N_10504);
or U10634 (N_10634,N_10525,N_10492);
xnor U10635 (N_10635,N_10427,N_10447);
nor U10636 (N_10636,N_10403,N_10437);
xnor U10637 (N_10637,N_10497,N_10507);
nor U10638 (N_10638,N_10574,N_10517);
xnor U10639 (N_10639,N_10402,N_10424);
or U10640 (N_10640,N_10494,N_10404);
and U10641 (N_10641,N_10519,N_10580);
nor U10642 (N_10642,N_10475,N_10435);
and U10643 (N_10643,N_10514,N_10432);
nand U10644 (N_10644,N_10480,N_10542);
xor U10645 (N_10645,N_10417,N_10476);
nor U10646 (N_10646,N_10415,N_10573);
xor U10647 (N_10647,N_10413,N_10474);
xor U10648 (N_10648,N_10594,N_10569);
nand U10649 (N_10649,N_10546,N_10462);
nand U10650 (N_10650,N_10595,N_10467);
and U10651 (N_10651,N_10438,N_10496);
or U10652 (N_10652,N_10501,N_10545);
nor U10653 (N_10653,N_10465,N_10416);
nor U10654 (N_10654,N_10448,N_10426);
and U10655 (N_10655,N_10453,N_10500);
or U10656 (N_10656,N_10479,N_10571);
nor U10657 (N_10657,N_10401,N_10536);
nor U10658 (N_10658,N_10486,N_10461);
or U10659 (N_10659,N_10590,N_10446);
nor U10660 (N_10660,N_10456,N_10543);
nand U10661 (N_10661,N_10422,N_10541);
nor U10662 (N_10662,N_10524,N_10576);
nor U10663 (N_10663,N_10495,N_10518);
nand U10664 (N_10664,N_10552,N_10444);
nand U10665 (N_10665,N_10513,N_10400);
or U10666 (N_10666,N_10583,N_10502);
xor U10667 (N_10667,N_10489,N_10506);
nand U10668 (N_10668,N_10463,N_10516);
nand U10669 (N_10669,N_10550,N_10445);
nand U10670 (N_10670,N_10585,N_10473);
nand U10671 (N_10671,N_10421,N_10488);
nor U10672 (N_10672,N_10530,N_10586);
nor U10673 (N_10673,N_10548,N_10477);
nand U10674 (N_10674,N_10485,N_10547);
and U10675 (N_10675,N_10539,N_10581);
nand U10676 (N_10676,N_10578,N_10470);
or U10677 (N_10677,N_10544,N_10460);
xnor U10678 (N_10678,N_10431,N_10509);
nand U10679 (N_10679,N_10556,N_10533);
or U10680 (N_10680,N_10563,N_10551);
and U10681 (N_10681,N_10567,N_10512);
xnor U10682 (N_10682,N_10503,N_10406);
nor U10683 (N_10683,N_10559,N_10414);
nor U10684 (N_10684,N_10505,N_10532);
or U10685 (N_10685,N_10592,N_10481);
xor U10686 (N_10686,N_10458,N_10575);
xor U10687 (N_10687,N_10457,N_10440);
nand U10688 (N_10688,N_10419,N_10570);
nor U10689 (N_10689,N_10484,N_10459);
xor U10690 (N_10690,N_10564,N_10527);
or U10691 (N_10691,N_10449,N_10584);
and U10692 (N_10692,N_10409,N_10454);
nand U10693 (N_10693,N_10490,N_10568);
or U10694 (N_10694,N_10593,N_10591);
xor U10695 (N_10695,N_10558,N_10588);
xnor U10696 (N_10696,N_10441,N_10425);
xor U10697 (N_10697,N_10523,N_10599);
and U10698 (N_10698,N_10508,N_10483);
nand U10699 (N_10699,N_10450,N_10428);
nor U10700 (N_10700,N_10463,N_10553);
and U10701 (N_10701,N_10591,N_10584);
and U10702 (N_10702,N_10541,N_10417);
and U10703 (N_10703,N_10571,N_10411);
nor U10704 (N_10704,N_10531,N_10477);
nor U10705 (N_10705,N_10514,N_10412);
and U10706 (N_10706,N_10512,N_10414);
or U10707 (N_10707,N_10598,N_10569);
nor U10708 (N_10708,N_10504,N_10577);
nor U10709 (N_10709,N_10484,N_10482);
nor U10710 (N_10710,N_10402,N_10516);
nor U10711 (N_10711,N_10448,N_10512);
nand U10712 (N_10712,N_10528,N_10421);
nand U10713 (N_10713,N_10527,N_10419);
nand U10714 (N_10714,N_10546,N_10449);
xor U10715 (N_10715,N_10481,N_10563);
nand U10716 (N_10716,N_10554,N_10581);
and U10717 (N_10717,N_10567,N_10464);
xor U10718 (N_10718,N_10468,N_10571);
nor U10719 (N_10719,N_10435,N_10426);
nor U10720 (N_10720,N_10429,N_10507);
and U10721 (N_10721,N_10408,N_10531);
or U10722 (N_10722,N_10430,N_10491);
nor U10723 (N_10723,N_10527,N_10423);
nor U10724 (N_10724,N_10543,N_10556);
nor U10725 (N_10725,N_10559,N_10495);
nand U10726 (N_10726,N_10407,N_10540);
xor U10727 (N_10727,N_10458,N_10561);
and U10728 (N_10728,N_10510,N_10464);
and U10729 (N_10729,N_10588,N_10519);
or U10730 (N_10730,N_10597,N_10549);
xor U10731 (N_10731,N_10497,N_10436);
or U10732 (N_10732,N_10491,N_10452);
nor U10733 (N_10733,N_10470,N_10544);
nor U10734 (N_10734,N_10416,N_10453);
nand U10735 (N_10735,N_10450,N_10429);
or U10736 (N_10736,N_10557,N_10571);
or U10737 (N_10737,N_10595,N_10464);
nor U10738 (N_10738,N_10426,N_10408);
nor U10739 (N_10739,N_10528,N_10592);
xnor U10740 (N_10740,N_10586,N_10432);
nor U10741 (N_10741,N_10529,N_10472);
and U10742 (N_10742,N_10429,N_10508);
xnor U10743 (N_10743,N_10404,N_10547);
and U10744 (N_10744,N_10499,N_10430);
nand U10745 (N_10745,N_10419,N_10568);
xor U10746 (N_10746,N_10429,N_10546);
nor U10747 (N_10747,N_10521,N_10581);
or U10748 (N_10748,N_10569,N_10505);
xor U10749 (N_10749,N_10519,N_10592);
or U10750 (N_10750,N_10408,N_10487);
nand U10751 (N_10751,N_10424,N_10455);
nor U10752 (N_10752,N_10596,N_10453);
xor U10753 (N_10753,N_10576,N_10570);
nor U10754 (N_10754,N_10430,N_10538);
and U10755 (N_10755,N_10487,N_10452);
xnor U10756 (N_10756,N_10414,N_10567);
or U10757 (N_10757,N_10554,N_10402);
nand U10758 (N_10758,N_10514,N_10556);
xnor U10759 (N_10759,N_10571,N_10524);
and U10760 (N_10760,N_10446,N_10533);
and U10761 (N_10761,N_10526,N_10570);
and U10762 (N_10762,N_10537,N_10467);
xor U10763 (N_10763,N_10569,N_10519);
or U10764 (N_10764,N_10466,N_10524);
nand U10765 (N_10765,N_10569,N_10424);
or U10766 (N_10766,N_10443,N_10548);
and U10767 (N_10767,N_10511,N_10522);
and U10768 (N_10768,N_10438,N_10551);
nand U10769 (N_10769,N_10571,N_10419);
and U10770 (N_10770,N_10572,N_10537);
or U10771 (N_10771,N_10479,N_10416);
xor U10772 (N_10772,N_10532,N_10523);
and U10773 (N_10773,N_10460,N_10458);
nor U10774 (N_10774,N_10563,N_10501);
nor U10775 (N_10775,N_10484,N_10587);
xor U10776 (N_10776,N_10586,N_10412);
and U10777 (N_10777,N_10503,N_10498);
nand U10778 (N_10778,N_10492,N_10575);
nor U10779 (N_10779,N_10430,N_10400);
nand U10780 (N_10780,N_10410,N_10584);
or U10781 (N_10781,N_10468,N_10496);
nor U10782 (N_10782,N_10520,N_10549);
xor U10783 (N_10783,N_10404,N_10426);
or U10784 (N_10784,N_10540,N_10591);
or U10785 (N_10785,N_10448,N_10465);
xor U10786 (N_10786,N_10580,N_10565);
xor U10787 (N_10787,N_10457,N_10403);
nand U10788 (N_10788,N_10581,N_10550);
and U10789 (N_10789,N_10492,N_10463);
nor U10790 (N_10790,N_10420,N_10549);
nor U10791 (N_10791,N_10489,N_10578);
or U10792 (N_10792,N_10492,N_10475);
and U10793 (N_10793,N_10539,N_10474);
and U10794 (N_10794,N_10483,N_10529);
nand U10795 (N_10795,N_10483,N_10543);
xnor U10796 (N_10796,N_10595,N_10455);
nand U10797 (N_10797,N_10493,N_10521);
nand U10798 (N_10798,N_10502,N_10478);
nand U10799 (N_10799,N_10580,N_10518);
nor U10800 (N_10800,N_10757,N_10739);
and U10801 (N_10801,N_10732,N_10616);
nor U10802 (N_10802,N_10665,N_10726);
or U10803 (N_10803,N_10646,N_10678);
nand U10804 (N_10804,N_10743,N_10668);
xor U10805 (N_10805,N_10642,N_10720);
or U10806 (N_10806,N_10606,N_10695);
nand U10807 (N_10807,N_10681,N_10765);
nor U10808 (N_10808,N_10618,N_10756);
xor U10809 (N_10809,N_10706,N_10745);
or U10810 (N_10810,N_10785,N_10603);
nand U10811 (N_10811,N_10685,N_10684);
xnor U10812 (N_10812,N_10741,N_10762);
nor U10813 (N_10813,N_10631,N_10654);
nand U10814 (N_10814,N_10620,N_10693);
xor U10815 (N_10815,N_10766,N_10664);
xor U10816 (N_10816,N_10612,N_10683);
nand U10817 (N_10817,N_10669,N_10780);
or U10818 (N_10818,N_10690,N_10666);
nor U10819 (N_10819,N_10600,N_10749);
nor U10820 (N_10820,N_10622,N_10751);
or U10821 (N_10821,N_10728,N_10737);
and U10822 (N_10822,N_10723,N_10602);
or U10823 (N_10823,N_10691,N_10713);
and U10824 (N_10824,N_10768,N_10790);
or U10825 (N_10825,N_10680,N_10722);
nand U10826 (N_10826,N_10619,N_10778);
or U10827 (N_10827,N_10747,N_10625);
or U10828 (N_10828,N_10609,N_10736);
or U10829 (N_10829,N_10613,N_10704);
xor U10830 (N_10830,N_10676,N_10639);
nor U10831 (N_10831,N_10742,N_10659);
or U10832 (N_10832,N_10675,N_10627);
nor U10833 (N_10833,N_10637,N_10754);
or U10834 (N_10834,N_10774,N_10764);
and U10835 (N_10835,N_10645,N_10710);
or U10836 (N_10836,N_10759,N_10791);
and U10837 (N_10837,N_10661,N_10730);
xnor U10838 (N_10838,N_10688,N_10655);
and U10839 (N_10839,N_10636,N_10779);
nand U10840 (N_10840,N_10799,N_10750);
and U10841 (N_10841,N_10748,N_10647);
or U10842 (N_10842,N_10628,N_10601);
or U10843 (N_10843,N_10672,N_10717);
xor U10844 (N_10844,N_10662,N_10776);
nor U10845 (N_10845,N_10740,N_10698);
nand U10846 (N_10846,N_10692,N_10657);
nand U10847 (N_10847,N_10670,N_10648);
xor U10848 (N_10848,N_10798,N_10604);
nand U10849 (N_10849,N_10772,N_10796);
or U10850 (N_10850,N_10608,N_10658);
or U10851 (N_10851,N_10701,N_10738);
and U10852 (N_10852,N_10682,N_10663);
nand U10853 (N_10853,N_10630,N_10746);
and U10854 (N_10854,N_10615,N_10786);
nor U10855 (N_10855,N_10715,N_10707);
or U10856 (N_10856,N_10641,N_10699);
xnor U10857 (N_10857,N_10649,N_10679);
or U10858 (N_10858,N_10703,N_10623);
nor U10859 (N_10859,N_10660,N_10714);
nand U10860 (N_10860,N_10752,N_10731);
nor U10861 (N_10861,N_10626,N_10610);
and U10862 (N_10862,N_10694,N_10783);
and U10863 (N_10863,N_10753,N_10797);
nor U10864 (N_10864,N_10696,N_10716);
or U10865 (N_10865,N_10640,N_10793);
or U10866 (N_10866,N_10725,N_10629);
nand U10867 (N_10867,N_10697,N_10673);
nand U10868 (N_10868,N_10607,N_10773);
nor U10869 (N_10869,N_10729,N_10687);
nand U10870 (N_10870,N_10769,N_10718);
and U10871 (N_10871,N_10605,N_10788);
nor U10872 (N_10872,N_10677,N_10643);
xnor U10873 (N_10873,N_10653,N_10724);
and U10874 (N_10874,N_10650,N_10667);
xor U10875 (N_10875,N_10775,N_10686);
xor U10876 (N_10876,N_10635,N_10763);
xnor U10877 (N_10877,N_10689,N_10709);
xor U10878 (N_10878,N_10767,N_10712);
nand U10879 (N_10879,N_10795,N_10789);
xnor U10880 (N_10880,N_10621,N_10634);
nor U10881 (N_10881,N_10651,N_10652);
xor U10882 (N_10882,N_10719,N_10782);
nor U10883 (N_10883,N_10656,N_10787);
and U10884 (N_10884,N_10708,N_10632);
or U10885 (N_10885,N_10735,N_10784);
nand U10886 (N_10886,N_10700,N_10761);
nand U10887 (N_10887,N_10771,N_10760);
or U10888 (N_10888,N_10721,N_10611);
and U10889 (N_10889,N_10770,N_10671);
nand U10890 (N_10890,N_10734,N_10633);
nor U10891 (N_10891,N_10792,N_10711);
and U10892 (N_10892,N_10727,N_10733);
xnor U10893 (N_10893,N_10624,N_10777);
nand U10894 (N_10894,N_10644,N_10617);
nor U10895 (N_10895,N_10674,N_10744);
nor U10896 (N_10896,N_10758,N_10638);
xnor U10897 (N_10897,N_10781,N_10794);
and U10898 (N_10898,N_10614,N_10755);
and U10899 (N_10899,N_10705,N_10702);
nor U10900 (N_10900,N_10680,N_10688);
nor U10901 (N_10901,N_10772,N_10769);
xor U10902 (N_10902,N_10785,N_10611);
or U10903 (N_10903,N_10690,N_10732);
nor U10904 (N_10904,N_10752,N_10730);
or U10905 (N_10905,N_10745,N_10651);
nor U10906 (N_10906,N_10639,N_10741);
xor U10907 (N_10907,N_10632,N_10787);
xor U10908 (N_10908,N_10784,N_10764);
nand U10909 (N_10909,N_10756,N_10743);
xnor U10910 (N_10910,N_10703,N_10796);
xnor U10911 (N_10911,N_10731,N_10737);
nand U10912 (N_10912,N_10702,N_10731);
and U10913 (N_10913,N_10696,N_10746);
or U10914 (N_10914,N_10769,N_10764);
and U10915 (N_10915,N_10757,N_10751);
and U10916 (N_10916,N_10605,N_10631);
xnor U10917 (N_10917,N_10688,N_10604);
nor U10918 (N_10918,N_10637,N_10733);
or U10919 (N_10919,N_10762,N_10682);
nand U10920 (N_10920,N_10716,N_10631);
nor U10921 (N_10921,N_10726,N_10630);
nand U10922 (N_10922,N_10663,N_10619);
and U10923 (N_10923,N_10793,N_10746);
or U10924 (N_10924,N_10682,N_10673);
or U10925 (N_10925,N_10642,N_10628);
or U10926 (N_10926,N_10635,N_10771);
nor U10927 (N_10927,N_10687,N_10733);
xnor U10928 (N_10928,N_10720,N_10615);
nand U10929 (N_10929,N_10797,N_10751);
or U10930 (N_10930,N_10686,N_10670);
nor U10931 (N_10931,N_10628,N_10734);
and U10932 (N_10932,N_10649,N_10683);
xor U10933 (N_10933,N_10697,N_10656);
nor U10934 (N_10934,N_10602,N_10690);
nor U10935 (N_10935,N_10709,N_10742);
xor U10936 (N_10936,N_10652,N_10771);
and U10937 (N_10937,N_10794,N_10696);
nand U10938 (N_10938,N_10708,N_10691);
nor U10939 (N_10939,N_10745,N_10730);
and U10940 (N_10940,N_10601,N_10660);
and U10941 (N_10941,N_10646,N_10724);
nor U10942 (N_10942,N_10640,N_10604);
nand U10943 (N_10943,N_10754,N_10686);
or U10944 (N_10944,N_10678,N_10606);
and U10945 (N_10945,N_10755,N_10746);
and U10946 (N_10946,N_10610,N_10748);
or U10947 (N_10947,N_10613,N_10701);
or U10948 (N_10948,N_10749,N_10636);
nor U10949 (N_10949,N_10788,N_10675);
nand U10950 (N_10950,N_10613,N_10609);
or U10951 (N_10951,N_10678,N_10751);
xnor U10952 (N_10952,N_10728,N_10673);
nor U10953 (N_10953,N_10789,N_10687);
xor U10954 (N_10954,N_10695,N_10742);
xnor U10955 (N_10955,N_10650,N_10744);
nand U10956 (N_10956,N_10784,N_10640);
xor U10957 (N_10957,N_10617,N_10646);
nor U10958 (N_10958,N_10733,N_10718);
nor U10959 (N_10959,N_10785,N_10604);
nor U10960 (N_10960,N_10606,N_10616);
xor U10961 (N_10961,N_10700,N_10698);
xnor U10962 (N_10962,N_10697,N_10643);
and U10963 (N_10963,N_10787,N_10765);
and U10964 (N_10964,N_10753,N_10674);
nand U10965 (N_10965,N_10770,N_10745);
and U10966 (N_10966,N_10763,N_10735);
nor U10967 (N_10967,N_10761,N_10628);
nand U10968 (N_10968,N_10600,N_10608);
or U10969 (N_10969,N_10625,N_10665);
or U10970 (N_10970,N_10639,N_10699);
xor U10971 (N_10971,N_10768,N_10731);
xnor U10972 (N_10972,N_10785,N_10751);
xor U10973 (N_10973,N_10740,N_10627);
nand U10974 (N_10974,N_10753,N_10683);
nor U10975 (N_10975,N_10725,N_10789);
or U10976 (N_10976,N_10602,N_10670);
nor U10977 (N_10977,N_10753,N_10611);
or U10978 (N_10978,N_10631,N_10673);
xnor U10979 (N_10979,N_10642,N_10657);
and U10980 (N_10980,N_10797,N_10720);
or U10981 (N_10981,N_10694,N_10620);
xnor U10982 (N_10982,N_10619,N_10719);
nor U10983 (N_10983,N_10650,N_10713);
and U10984 (N_10984,N_10677,N_10788);
nor U10985 (N_10985,N_10788,N_10648);
and U10986 (N_10986,N_10661,N_10731);
and U10987 (N_10987,N_10704,N_10627);
xnor U10988 (N_10988,N_10725,N_10780);
or U10989 (N_10989,N_10740,N_10695);
or U10990 (N_10990,N_10603,N_10761);
or U10991 (N_10991,N_10677,N_10701);
nor U10992 (N_10992,N_10701,N_10639);
or U10993 (N_10993,N_10648,N_10715);
nand U10994 (N_10994,N_10622,N_10750);
or U10995 (N_10995,N_10789,N_10649);
nand U10996 (N_10996,N_10678,N_10652);
and U10997 (N_10997,N_10650,N_10742);
xnor U10998 (N_10998,N_10738,N_10613);
and U10999 (N_10999,N_10671,N_10714);
or U11000 (N_11000,N_10847,N_10848);
or U11001 (N_11001,N_10886,N_10835);
or U11002 (N_11002,N_10809,N_10918);
and U11003 (N_11003,N_10859,N_10868);
and U11004 (N_11004,N_10992,N_10873);
xnor U11005 (N_11005,N_10861,N_10857);
and U11006 (N_11006,N_10910,N_10947);
xor U11007 (N_11007,N_10860,N_10998);
and U11008 (N_11008,N_10999,N_10872);
xor U11009 (N_11009,N_10936,N_10834);
nand U11010 (N_11010,N_10993,N_10916);
and U11011 (N_11011,N_10802,N_10813);
or U11012 (N_11012,N_10931,N_10980);
xor U11013 (N_11013,N_10829,N_10850);
nand U11014 (N_11014,N_10865,N_10969);
or U11015 (N_11015,N_10823,N_10811);
nor U11016 (N_11016,N_10909,N_10880);
xnor U11017 (N_11017,N_10946,N_10950);
and U11018 (N_11018,N_10952,N_10884);
xnor U11019 (N_11019,N_10849,N_10994);
and U11020 (N_11020,N_10995,N_10845);
nand U11021 (N_11021,N_10854,N_10954);
or U11022 (N_11022,N_10907,N_10912);
nand U11023 (N_11023,N_10897,N_10940);
nand U11024 (N_11024,N_10807,N_10958);
and U11025 (N_11025,N_10824,N_10917);
or U11026 (N_11026,N_10810,N_10836);
nand U11027 (N_11027,N_10948,N_10890);
and U11028 (N_11028,N_10988,N_10830);
nor U11029 (N_11029,N_10817,N_10800);
and U11030 (N_11030,N_10899,N_10882);
xnor U11031 (N_11031,N_10806,N_10875);
nand U11032 (N_11032,N_10844,N_10920);
and U11033 (N_11033,N_10826,N_10957);
and U11034 (N_11034,N_10972,N_10922);
nand U11035 (N_11035,N_10989,N_10891);
or U11036 (N_11036,N_10963,N_10951);
nand U11037 (N_11037,N_10863,N_10964);
nor U11038 (N_11038,N_10961,N_10892);
xnor U11039 (N_11039,N_10828,N_10820);
xor U11040 (N_11040,N_10911,N_10938);
xor U11041 (N_11041,N_10943,N_10979);
or U11042 (N_11042,N_10804,N_10887);
and U11043 (N_11043,N_10852,N_10978);
and U11044 (N_11044,N_10855,N_10827);
nand U11045 (N_11045,N_10864,N_10839);
xor U11046 (N_11046,N_10831,N_10926);
and U11047 (N_11047,N_10895,N_10900);
or U11048 (N_11048,N_10984,N_10846);
nor U11049 (N_11049,N_10919,N_10945);
xnor U11050 (N_11050,N_10906,N_10930);
nand U11051 (N_11051,N_10959,N_10986);
xnor U11052 (N_11052,N_10808,N_10935);
nor U11053 (N_11053,N_10915,N_10966);
and U11054 (N_11054,N_10821,N_10944);
xnor U11055 (N_11055,N_10866,N_10914);
nor U11056 (N_11056,N_10801,N_10965);
or U11057 (N_11057,N_10840,N_10949);
and U11058 (N_11058,N_10924,N_10903);
xnor U11059 (N_11059,N_10913,N_10990);
nor U11060 (N_11060,N_10894,N_10888);
nor U11061 (N_11061,N_10832,N_10838);
or U11062 (N_11062,N_10968,N_10904);
or U11063 (N_11063,N_10960,N_10869);
nand U11064 (N_11064,N_10837,N_10973);
and U11065 (N_11065,N_10982,N_10893);
or U11066 (N_11066,N_10889,N_10997);
and U11067 (N_11067,N_10833,N_10942);
nor U11068 (N_11068,N_10929,N_10883);
nand U11069 (N_11069,N_10853,N_10812);
xor U11070 (N_11070,N_10939,N_10941);
or U11071 (N_11071,N_10885,N_10843);
and U11072 (N_11072,N_10953,N_10818);
and U11073 (N_11073,N_10921,N_10923);
or U11074 (N_11074,N_10876,N_10819);
nand U11075 (N_11075,N_10967,N_10970);
or U11076 (N_11076,N_10987,N_10825);
nor U11077 (N_11077,N_10908,N_10955);
or U11078 (N_11078,N_10983,N_10996);
nor U11079 (N_11079,N_10932,N_10977);
nand U11080 (N_11080,N_10878,N_10871);
nor U11081 (N_11081,N_10803,N_10816);
xnor U11082 (N_11082,N_10877,N_10856);
nand U11083 (N_11083,N_10974,N_10862);
xnor U11084 (N_11084,N_10822,N_10896);
nand U11085 (N_11085,N_10934,N_10933);
xor U11086 (N_11086,N_10962,N_10805);
nand U11087 (N_11087,N_10981,N_10901);
or U11088 (N_11088,N_10902,N_10975);
nor U11089 (N_11089,N_10905,N_10925);
xnor U11090 (N_11090,N_10985,N_10991);
and U11091 (N_11091,N_10956,N_10842);
or U11092 (N_11092,N_10976,N_10879);
and U11093 (N_11093,N_10928,N_10927);
xor U11094 (N_11094,N_10881,N_10814);
or U11095 (N_11095,N_10971,N_10898);
xnor U11096 (N_11096,N_10874,N_10937);
or U11097 (N_11097,N_10841,N_10851);
or U11098 (N_11098,N_10867,N_10858);
nand U11099 (N_11099,N_10815,N_10870);
or U11100 (N_11100,N_10831,N_10907);
nand U11101 (N_11101,N_10839,N_10927);
xor U11102 (N_11102,N_10808,N_10877);
xor U11103 (N_11103,N_10818,N_10805);
nand U11104 (N_11104,N_10807,N_10881);
xnor U11105 (N_11105,N_10911,N_10988);
or U11106 (N_11106,N_10853,N_10911);
xnor U11107 (N_11107,N_10879,N_10979);
or U11108 (N_11108,N_10957,N_10851);
nor U11109 (N_11109,N_10871,N_10910);
and U11110 (N_11110,N_10878,N_10993);
nand U11111 (N_11111,N_10839,N_10866);
or U11112 (N_11112,N_10829,N_10801);
and U11113 (N_11113,N_10941,N_10857);
xor U11114 (N_11114,N_10975,N_10910);
or U11115 (N_11115,N_10894,N_10825);
xor U11116 (N_11116,N_10815,N_10993);
and U11117 (N_11117,N_10872,N_10907);
nand U11118 (N_11118,N_10910,N_10821);
nand U11119 (N_11119,N_10962,N_10985);
or U11120 (N_11120,N_10894,N_10927);
nor U11121 (N_11121,N_10900,N_10842);
or U11122 (N_11122,N_10917,N_10934);
xnor U11123 (N_11123,N_10975,N_10988);
and U11124 (N_11124,N_10902,N_10994);
and U11125 (N_11125,N_10862,N_10900);
nor U11126 (N_11126,N_10973,N_10926);
or U11127 (N_11127,N_10834,N_10973);
or U11128 (N_11128,N_10877,N_10969);
and U11129 (N_11129,N_10957,N_10968);
nand U11130 (N_11130,N_10962,N_10954);
or U11131 (N_11131,N_10818,N_10971);
xor U11132 (N_11132,N_10969,N_10947);
and U11133 (N_11133,N_10884,N_10906);
and U11134 (N_11134,N_10857,N_10836);
or U11135 (N_11135,N_10876,N_10965);
nor U11136 (N_11136,N_10961,N_10918);
xor U11137 (N_11137,N_10818,N_10895);
and U11138 (N_11138,N_10851,N_10816);
and U11139 (N_11139,N_10878,N_10891);
and U11140 (N_11140,N_10914,N_10833);
xnor U11141 (N_11141,N_10904,N_10851);
nand U11142 (N_11142,N_10858,N_10961);
xor U11143 (N_11143,N_10960,N_10957);
xor U11144 (N_11144,N_10863,N_10933);
nand U11145 (N_11145,N_10885,N_10810);
nand U11146 (N_11146,N_10837,N_10956);
or U11147 (N_11147,N_10858,N_10933);
nor U11148 (N_11148,N_10885,N_10837);
xor U11149 (N_11149,N_10832,N_10826);
or U11150 (N_11150,N_10936,N_10945);
nor U11151 (N_11151,N_10826,N_10827);
nor U11152 (N_11152,N_10933,N_10809);
and U11153 (N_11153,N_10999,N_10887);
nor U11154 (N_11154,N_10865,N_10872);
and U11155 (N_11155,N_10829,N_10817);
and U11156 (N_11156,N_10944,N_10969);
nand U11157 (N_11157,N_10872,N_10822);
or U11158 (N_11158,N_10862,N_10865);
nor U11159 (N_11159,N_10801,N_10824);
or U11160 (N_11160,N_10830,N_10962);
nand U11161 (N_11161,N_10955,N_10873);
or U11162 (N_11162,N_10879,N_10857);
nand U11163 (N_11163,N_10841,N_10861);
and U11164 (N_11164,N_10884,N_10822);
xor U11165 (N_11165,N_10856,N_10804);
nand U11166 (N_11166,N_10970,N_10840);
or U11167 (N_11167,N_10875,N_10952);
and U11168 (N_11168,N_10981,N_10875);
or U11169 (N_11169,N_10939,N_10874);
xor U11170 (N_11170,N_10821,N_10984);
or U11171 (N_11171,N_10895,N_10846);
nor U11172 (N_11172,N_10953,N_10817);
nor U11173 (N_11173,N_10992,N_10865);
and U11174 (N_11174,N_10872,N_10838);
and U11175 (N_11175,N_10899,N_10800);
xor U11176 (N_11176,N_10920,N_10867);
xnor U11177 (N_11177,N_10939,N_10825);
nand U11178 (N_11178,N_10928,N_10806);
xor U11179 (N_11179,N_10803,N_10926);
and U11180 (N_11180,N_10839,N_10826);
xor U11181 (N_11181,N_10890,N_10931);
and U11182 (N_11182,N_10983,N_10969);
nor U11183 (N_11183,N_10890,N_10927);
or U11184 (N_11184,N_10976,N_10890);
nor U11185 (N_11185,N_10844,N_10950);
xor U11186 (N_11186,N_10835,N_10978);
xor U11187 (N_11187,N_10834,N_10839);
and U11188 (N_11188,N_10923,N_10823);
nor U11189 (N_11189,N_10897,N_10974);
and U11190 (N_11190,N_10856,N_10955);
nor U11191 (N_11191,N_10839,N_10972);
and U11192 (N_11192,N_10953,N_10861);
or U11193 (N_11193,N_10991,N_10992);
and U11194 (N_11194,N_10936,N_10967);
or U11195 (N_11195,N_10815,N_10878);
and U11196 (N_11196,N_10999,N_10938);
nand U11197 (N_11197,N_10989,N_10831);
and U11198 (N_11198,N_10889,N_10941);
or U11199 (N_11199,N_10922,N_10841);
nand U11200 (N_11200,N_11065,N_11145);
nand U11201 (N_11201,N_11054,N_11039);
xnor U11202 (N_11202,N_11155,N_11128);
and U11203 (N_11203,N_11001,N_11186);
nand U11204 (N_11204,N_11104,N_11025);
nand U11205 (N_11205,N_11179,N_11116);
xnor U11206 (N_11206,N_11092,N_11082);
or U11207 (N_11207,N_11070,N_11156);
xnor U11208 (N_11208,N_11122,N_11166);
or U11209 (N_11209,N_11002,N_11044);
nand U11210 (N_11210,N_11120,N_11137);
nor U11211 (N_11211,N_11091,N_11098);
xor U11212 (N_11212,N_11124,N_11151);
nand U11213 (N_11213,N_11060,N_11078);
and U11214 (N_11214,N_11071,N_11014);
xor U11215 (N_11215,N_11132,N_11084);
and U11216 (N_11216,N_11051,N_11168);
or U11217 (N_11217,N_11093,N_11004);
nor U11218 (N_11218,N_11135,N_11141);
nor U11219 (N_11219,N_11022,N_11152);
nor U11220 (N_11220,N_11016,N_11094);
nand U11221 (N_11221,N_11008,N_11089);
xnor U11222 (N_11222,N_11198,N_11000);
xor U11223 (N_11223,N_11061,N_11036);
xor U11224 (N_11224,N_11123,N_11131);
nand U11225 (N_11225,N_11020,N_11046);
xor U11226 (N_11226,N_11146,N_11011);
xnor U11227 (N_11227,N_11043,N_11075);
or U11228 (N_11228,N_11118,N_11047);
xor U11229 (N_11229,N_11096,N_11176);
and U11230 (N_11230,N_11073,N_11191);
or U11231 (N_11231,N_11095,N_11041);
xor U11232 (N_11232,N_11068,N_11045);
and U11233 (N_11233,N_11019,N_11052);
nor U11234 (N_11234,N_11110,N_11090);
nor U11235 (N_11235,N_11017,N_11050);
or U11236 (N_11236,N_11064,N_11030);
xor U11237 (N_11237,N_11149,N_11144);
xor U11238 (N_11238,N_11088,N_11150);
nand U11239 (N_11239,N_11180,N_11081);
xor U11240 (N_11240,N_11021,N_11034);
xnor U11241 (N_11241,N_11188,N_11049);
nor U11242 (N_11242,N_11080,N_11109);
and U11243 (N_11243,N_11053,N_11174);
or U11244 (N_11244,N_11038,N_11035);
or U11245 (N_11245,N_11161,N_11063);
nand U11246 (N_11246,N_11074,N_11157);
nand U11247 (N_11247,N_11140,N_11076);
nand U11248 (N_11248,N_11024,N_11115);
and U11249 (N_11249,N_11029,N_11077);
nor U11250 (N_11250,N_11005,N_11111);
nor U11251 (N_11251,N_11102,N_11165);
or U11252 (N_11252,N_11187,N_11085);
and U11253 (N_11253,N_11028,N_11100);
or U11254 (N_11254,N_11164,N_11015);
and U11255 (N_11255,N_11169,N_11127);
nor U11256 (N_11256,N_11117,N_11108);
nand U11257 (N_11257,N_11101,N_11148);
and U11258 (N_11258,N_11172,N_11113);
and U11259 (N_11259,N_11107,N_11125);
xnor U11260 (N_11260,N_11066,N_11031);
and U11261 (N_11261,N_11196,N_11190);
xor U11262 (N_11262,N_11097,N_11010);
nand U11263 (N_11263,N_11106,N_11193);
nand U11264 (N_11264,N_11033,N_11087);
nor U11265 (N_11265,N_11099,N_11136);
or U11266 (N_11266,N_11121,N_11163);
nand U11267 (N_11267,N_11027,N_11194);
xnor U11268 (N_11268,N_11129,N_11167);
xor U11269 (N_11269,N_11197,N_11042);
xor U11270 (N_11270,N_11086,N_11184);
nor U11271 (N_11271,N_11160,N_11055);
and U11272 (N_11272,N_11143,N_11079);
xor U11273 (N_11273,N_11026,N_11009);
nand U11274 (N_11274,N_11181,N_11040);
or U11275 (N_11275,N_11185,N_11175);
or U11276 (N_11276,N_11006,N_11199);
and U11277 (N_11277,N_11139,N_11147);
nand U11278 (N_11278,N_11057,N_11032);
and U11279 (N_11279,N_11067,N_11062);
xnor U11280 (N_11280,N_11134,N_11153);
nand U11281 (N_11281,N_11182,N_11112);
and U11282 (N_11282,N_11171,N_11119);
or U11283 (N_11283,N_11058,N_11007);
nand U11284 (N_11284,N_11023,N_11012);
xnor U11285 (N_11285,N_11083,N_11142);
or U11286 (N_11286,N_11003,N_11130);
nand U11287 (N_11287,N_11114,N_11013);
nand U11288 (N_11288,N_11059,N_11105);
nand U11289 (N_11289,N_11126,N_11189);
or U11290 (N_11290,N_11103,N_11133);
nor U11291 (N_11291,N_11192,N_11154);
xor U11292 (N_11292,N_11173,N_11195);
and U11293 (N_11293,N_11037,N_11158);
nand U11294 (N_11294,N_11056,N_11069);
nor U11295 (N_11295,N_11177,N_11162);
nand U11296 (N_11296,N_11178,N_11018);
nand U11297 (N_11297,N_11072,N_11170);
nand U11298 (N_11298,N_11183,N_11138);
xor U11299 (N_11299,N_11159,N_11048);
xnor U11300 (N_11300,N_11166,N_11025);
or U11301 (N_11301,N_11038,N_11150);
nand U11302 (N_11302,N_11082,N_11136);
and U11303 (N_11303,N_11153,N_11183);
xor U11304 (N_11304,N_11122,N_11033);
xor U11305 (N_11305,N_11006,N_11170);
xor U11306 (N_11306,N_11096,N_11123);
xnor U11307 (N_11307,N_11094,N_11088);
or U11308 (N_11308,N_11159,N_11023);
and U11309 (N_11309,N_11148,N_11199);
nand U11310 (N_11310,N_11011,N_11170);
nand U11311 (N_11311,N_11068,N_11100);
xnor U11312 (N_11312,N_11137,N_11192);
or U11313 (N_11313,N_11122,N_11109);
xnor U11314 (N_11314,N_11125,N_11070);
nand U11315 (N_11315,N_11015,N_11081);
nand U11316 (N_11316,N_11117,N_11086);
nor U11317 (N_11317,N_11058,N_11181);
nor U11318 (N_11318,N_11091,N_11137);
and U11319 (N_11319,N_11178,N_11120);
nand U11320 (N_11320,N_11115,N_11113);
nor U11321 (N_11321,N_11177,N_11016);
or U11322 (N_11322,N_11182,N_11197);
nand U11323 (N_11323,N_11071,N_11074);
nor U11324 (N_11324,N_11044,N_11189);
or U11325 (N_11325,N_11183,N_11165);
nand U11326 (N_11326,N_11022,N_11050);
xnor U11327 (N_11327,N_11098,N_11147);
xnor U11328 (N_11328,N_11027,N_11112);
xor U11329 (N_11329,N_11085,N_11074);
nor U11330 (N_11330,N_11021,N_11032);
and U11331 (N_11331,N_11098,N_11188);
and U11332 (N_11332,N_11158,N_11083);
nor U11333 (N_11333,N_11053,N_11022);
xnor U11334 (N_11334,N_11051,N_11108);
nor U11335 (N_11335,N_11125,N_11010);
xnor U11336 (N_11336,N_11103,N_11145);
or U11337 (N_11337,N_11076,N_11037);
or U11338 (N_11338,N_11035,N_11171);
or U11339 (N_11339,N_11092,N_11107);
nor U11340 (N_11340,N_11094,N_11145);
nand U11341 (N_11341,N_11016,N_11100);
nor U11342 (N_11342,N_11128,N_11031);
nand U11343 (N_11343,N_11013,N_11186);
or U11344 (N_11344,N_11127,N_11096);
nor U11345 (N_11345,N_11145,N_11154);
nor U11346 (N_11346,N_11024,N_11013);
nor U11347 (N_11347,N_11162,N_11155);
and U11348 (N_11348,N_11155,N_11096);
xor U11349 (N_11349,N_11109,N_11160);
xnor U11350 (N_11350,N_11170,N_11091);
nand U11351 (N_11351,N_11076,N_11039);
or U11352 (N_11352,N_11188,N_11169);
xor U11353 (N_11353,N_11021,N_11091);
and U11354 (N_11354,N_11112,N_11143);
xnor U11355 (N_11355,N_11032,N_11161);
and U11356 (N_11356,N_11052,N_11036);
nor U11357 (N_11357,N_11059,N_11165);
and U11358 (N_11358,N_11029,N_11110);
nand U11359 (N_11359,N_11180,N_11094);
xnor U11360 (N_11360,N_11031,N_11077);
xor U11361 (N_11361,N_11131,N_11073);
xor U11362 (N_11362,N_11065,N_11176);
or U11363 (N_11363,N_11028,N_11083);
and U11364 (N_11364,N_11056,N_11151);
nor U11365 (N_11365,N_11112,N_11066);
and U11366 (N_11366,N_11022,N_11074);
or U11367 (N_11367,N_11171,N_11010);
nand U11368 (N_11368,N_11088,N_11139);
nand U11369 (N_11369,N_11185,N_11067);
nand U11370 (N_11370,N_11005,N_11138);
xnor U11371 (N_11371,N_11118,N_11155);
nand U11372 (N_11372,N_11078,N_11067);
and U11373 (N_11373,N_11012,N_11118);
xnor U11374 (N_11374,N_11189,N_11187);
xor U11375 (N_11375,N_11141,N_11116);
xor U11376 (N_11376,N_11164,N_11078);
and U11377 (N_11377,N_11151,N_11139);
nor U11378 (N_11378,N_11141,N_11054);
nor U11379 (N_11379,N_11011,N_11061);
nand U11380 (N_11380,N_11066,N_11178);
nor U11381 (N_11381,N_11084,N_11062);
nor U11382 (N_11382,N_11190,N_11099);
and U11383 (N_11383,N_11169,N_11082);
nand U11384 (N_11384,N_11132,N_11003);
nor U11385 (N_11385,N_11183,N_11159);
nor U11386 (N_11386,N_11026,N_11178);
nand U11387 (N_11387,N_11024,N_11193);
or U11388 (N_11388,N_11084,N_11102);
nor U11389 (N_11389,N_11027,N_11069);
or U11390 (N_11390,N_11132,N_11021);
and U11391 (N_11391,N_11056,N_11063);
or U11392 (N_11392,N_11127,N_11107);
nand U11393 (N_11393,N_11136,N_11024);
nor U11394 (N_11394,N_11084,N_11044);
nor U11395 (N_11395,N_11051,N_11172);
and U11396 (N_11396,N_11026,N_11008);
or U11397 (N_11397,N_11175,N_11154);
or U11398 (N_11398,N_11091,N_11120);
xor U11399 (N_11399,N_11015,N_11098);
or U11400 (N_11400,N_11235,N_11222);
and U11401 (N_11401,N_11319,N_11278);
nor U11402 (N_11402,N_11224,N_11265);
nand U11403 (N_11403,N_11399,N_11277);
or U11404 (N_11404,N_11321,N_11322);
and U11405 (N_11405,N_11326,N_11226);
nand U11406 (N_11406,N_11266,N_11395);
and U11407 (N_11407,N_11203,N_11288);
xnor U11408 (N_11408,N_11295,N_11343);
and U11409 (N_11409,N_11306,N_11355);
and U11410 (N_11410,N_11251,N_11318);
or U11411 (N_11411,N_11280,N_11334);
xor U11412 (N_11412,N_11371,N_11365);
xor U11413 (N_11413,N_11219,N_11383);
and U11414 (N_11414,N_11254,N_11381);
or U11415 (N_11415,N_11230,N_11216);
and U11416 (N_11416,N_11303,N_11373);
or U11417 (N_11417,N_11301,N_11210);
or U11418 (N_11418,N_11233,N_11349);
nor U11419 (N_11419,N_11332,N_11357);
xnor U11420 (N_11420,N_11236,N_11243);
nand U11421 (N_11421,N_11356,N_11275);
or U11422 (N_11422,N_11341,N_11229);
and U11423 (N_11423,N_11300,N_11329);
xor U11424 (N_11424,N_11220,N_11264);
or U11425 (N_11425,N_11297,N_11271);
or U11426 (N_11426,N_11209,N_11268);
nor U11427 (N_11427,N_11377,N_11286);
nand U11428 (N_11428,N_11363,N_11388);
or U11429 (N_11429,N_11270,N_11259);
or U11430 (N_11430,N_11240,N_11281);
and U11431 (N_11431,N_11354,N_11232);
xor U11432 (N_11432,N_11390,N_11276);
or U11433 (N_11433,N_11228,N_11338);
or U11434 (N_11434,N_11227,N_11316);
and U11435 (N_11435,N_11342,N_11244);
and U11436 (N_11436,N_11293,N_11258);
or U11437 (N_11437,N_11290,N_11215);
xor U11438 (N_11438,N_11375,N_11246);
nand U11439 (N_11439,N_11282,N_11291);
nand U11440 (N_11440,N_11211,N_11292);
xnor U11441 (N_11441,N_11328,N_11369);
xnor U11442 (N_11442,N_11320,N_11335);
nor U11443 (N_11443,N_11362,N_11393);
nor U11444 (N_11444,N_11304,N_11392);
or U11445 (N_11445,N_11336,N_11340);
nor U11446 (N_11446,N_11376,N_11380);
or U11447 (N_11447,N_11249,N_11333);
xor U11448 (N_11448,N_11253,N_11361);
and U11449 (N_11449,N_11331,N_11315);
and U11450 (N_11450,N_11261,N_11242);
nand U11451 (N_11451,N_11346,N_11269);
nor U11452 (N_11452,N_11372,N_11260);
and U11453 (N_11453,N_11311,N_11370);
xor U11454 (N_11454,N_11379,N_11359);
xor U11455 (N_11455,N_11206,N_11223);
xnor U11456 (N_11456,N_11284,N_11348);
xnor U11457 (N_11457,N_11294,N_11386);
nand U11458 (N_11458,N_11207,N_11391);
xnor U11459 (N_11459,N_11201,N_11307);
nor U11460 (N_11460,N_11360,N_11325);
and U11461 (N_11461,N_11274,N_11323);
xor U11462 (N_11462,N_11263,N_11313);
nand U11463 (N_11463,N_11256,N_11353);
or U11464 (N_11464,N_11351,N_11324);
nand U11465 (N_11465,N_11345,N_11279);
and U11466 (N_11466,N_11344,N_11218);
xnor U11467 (N_11467,N_11250,N_11289);
nand U11468 (N_11468,N_11204,N_11382);
nand U11469 (N_11469,N_11337,N_11396);
and U11470 (N_11470,N_11225,N_11310);
xor U11471 (N_11471,N_11364,N_11330);
and U11472 (N_11472,N_11299,N_11394);
nand U11473 (N_11473,N_11398,N_11366);
nor U11474 (N_11474,N_11314,N_11385);
nand U11475 (N_11475,N_11285,N_11298);
nand U11476 (N_11476,N_11309,N_11257);
xnor U11477 (N_11477,N_11214,N_11212);
nand U11478 (N_11478,N_11208,N_11241);
or U11479 (N_11479,N_11272,N_11384);
or U11480 (N_11480,N_11327,N_11347);
nor U11481 (N_11481,N_11374,N_11273);
or U11482 (N_11482,N_11202,N_11287);
nand U11483 (N_11483,N_11317,N_11387);
nand U11484 (N_11484,N_11248,N_11283);
nor U11485 (N_11485,N_11238,N_11247);
and U11486 (N_11486,N_11255,N_11308);
xnor U11487 (N_11487,N_11267,N_11231);
xnor U11488 (N_11488,N_11217,N_11221);
nor U11489 (N_11489,N_11312,N_11262);
and U11490 (N_11490,N_11389,N_11358);
and U11491 (N_11491,N_11296,N_11367);
and U11492 (N_11492,N_11237,N_11368);
xnor U11493 (N_11493,N_11302,N_11397);
and U11494 (N_11494,N_11200,N_11378);
and U11495 (N_11495,N_11305,N_11252);
nand U11496 (N_11496,N_11239,N_11245);
nand U11497 (N_11497,N_11213,N_11339);
nand U11498 (N_11498,N_11205,N_11234);
and U11499 (N_11499,N_11352,N_11350);
or U11500 (N_11500,N_11202,N_11378);
nor U11501 (N_11501,N_11302,N_11329);
and U11502 (N_11502,N_11391,N_11242);
nor U11503 (N_11503,N_11369,N_11363);
and U11504 (N_11504,N_11219,N_11366);
or U11505 (N_11505,N_11290,N_11216);
nand U11506 (N_11506,N_11313,N_11354);
and U11507 (N_11507,N_11244,N_11236);
nor U11508 (N_11508,N_11334,N_11239);
nor U11509 (N_11509,N_11255,N_11299);
nor U11510 (N_11510,N_11202,N_11364);
nand U11511 (N_11511,N_11284,N_11393);
or U11512 (N_11512,N_11277,N_11243);
xor U11513 (N_11513,N_11205,N_11302);
and U11514 (N_11514,N_11350,N_11367);
and U11515 (N_11515,N_11378,N_11335);
xnor U11516 (N_11516,N_11250,N_11333);
or U11517 (N_11517,N_11265,N_11319);
or U11518 (N_11518,N_11379,N_11317);
nor U11519 (N_11519,N_11302,N_11218);
and U11520 (N_11520,N_11315,N_11300);
or U11521 (N_11521,N_11228,N_11330);
nor U11522 (N_11522,N_11380,N_11304);
or U11523 (N_11523,N_11274,N_11310);
xnor U11524 (N_11524,N_11325,N_11311);
nand U11525 (N_11525,N_11258,N_11220);
nor U11526 (N_11526,N_11361,N_11227);
nand U11527 (N_11527,N_11201,N_11351);
and U11528 (N_11528,N_11363,N_11361);
nand U11529 (N_11529,N_11294,N_11221);
and U11530 (N_11530,N_11351,N_11290);
xor U11531 (N_11531,N_11281,N_11354);
nor U11532 (N_11532,N_11311,N_11379);
and U11533 (N_11533,N_11336,N_11341);
nor U11534 (N_11534,N_11342,N_11209);
and U11535 (N_11535,N_11341,N_11347);
xor U11536 (N_11536,N_11282,N_11373);
and U11537 (N_11537,N_11260,N_11364);
nand U11538 (N_11538,N_11274,N_11209);
and U11539 (N_11539,N_11371,N_11323);
or U11540 (N_11540,N_11303,N_11306);
xnor U11541 (N_11541,N_11313,N_11256);
xor U11542 (N_11542,N_11295,N_11262);
nor U11543 (N_11543,N_11398,N_11389);
xor U11544 (N_11544,N_11379,N_11336);
or U11545 (N_11545,N_11271,N_11334);
and U11546 (N_11546,N_11297,N_11313);
and U11547 (N_11547,N_11321,N_11338);
and U11548 (N_11548,N_11309,N_11294);
or U11549 (N_11549,N_11267,N_11248);
nor U11550 (N_11550,N_11303,N_11285);
xor U11551 (N_11551,N_11238,N_11278);
or U11552 (N_11552,N_11334,N_11266);
and U11553 (N_11553,N_11294,N_11232);
nor U11554 (N_11554,N_11301,N_11309);
nor U11555 (N_11555,N_11232,N_11269);
and U11556 (N_11556,N_11238,N_11383);
and U11557 (N_11557,N_11356,N_11253);
nand U11558 (N_11558,N_11322,N_11225);
xor U11559 (N_11559,N_11284,N_11232);
nand U11560 (N_11560,N_11351,N_11241);
nor U11561 (N_11561,N_11262,N_11290);
or U11562 (N_11562,N_11353,N_11324);
or U11563 (N_11563,N_11350,N_11210);
nand U11564 (N_11564,N_11384,N_11287);
nand U11565 (N_11565,N_11215,N_11390);
nor U11566 (N_11566,N_11299,N_11359);
nor U11567 (N_11567,N_11361,N_11378);
nand U11568 (N_11568,N_11328,N_11390);
and U11569 (N_11569,N_11323,N_11346);
nor U11570 (N_11570,N_11309,N_11339);
and U11571 (N_11571,N_11392,N_11292);
nand U11572 (N_11572,N_11220,N_11295);
and U11573 (N_11573,N_11322,N_11323);
nand U11574 (N_11574,N_11282,N_11398);
or U11575 (N_11575,N_11321,N_11373);
nor U11576 (N_11576,N_11316,N_11290);
nor U11577 (N_11577,N_11275,N_11389);
and U11578 (N_11578,N_11384,N_11387);
and U11579 (N_11579,N_11266,N_11275);
and U11580 (N_11580,N_11253,N_11337);
or U11581 (N_11581,N_11365,N_11349);
or U11582 (N_11582,N_11394,N_11303);
xnor U11583 (N_11583,N_11326,N_11282);
nor U11584 (N_11584,N_11384,N_11363);
and U11585 (N_11585,N_11319,N_11246);
xnor U11586 (N_11586,N_11373,N_11257);
xnor U11587 (N_11587,N_11311,N_11237);
xnor U11588 (N_11588,N_11217,N_11345);
or U11589 (N_11589,N_11292,N_11299);
xor U11590 (N_11590,N_11285,N_11205);
nand U11591 (N_11591,N_11359,N_11384);
nor U11592 (N_11592,N_11366,N_11302);
xor U11593 (N_11593,N_11358,N_11329);
nand U11594 (N_11594,N_11290,N_11375);
or U11595 (N_11595,N_11372,N_11337);
or U11596 (N_11596,N_11283,N_11384);
nor U11597 (N_11597,N_11271,N_11266);
or U11598 (N_11598,N_11307,N_11203);
nand U11599 (N_11599,N_11348,N_11343);
and U11600 (N_11600,N_11528,N_11516);
nor U11601 (N_11601,N_11475,N_11535);
or U11602 (N_11602,N_11546,N_11442);
nor U11603 (N_11603,N_11463,N_11555);
nand U11604 (N_11604,N_11542,N_11428);
and U11605 (N_11605,N_11552,N_11510);
nand U11606 (N_11606,N_11511,N_11400);
and U11607 (N_11607,N_11583,N_11533);
or U11608 (N_11608,N_11570,N_11518);
and U11609 (N_11609,N_11407,N_11461);
and U11610 (N_11610,N_11573,N_11596);
or U11611 (N_11611,N_11543,N_11544);
or U11612 (N_11612,N_11598,N_11450);
and U11613 (N_11613,N_11416,N_11556);
and U11614 (N_11614,N_11430,N_11575);
xnor U11615 (N_11615,N_11531,N_11420);
or U11616 (N_11616,N_11480,N_11433);
nand U11617 (N_11617,N_11589,N_11427);
nand U11618 (N_11618,N_11536,N_11486);
nand U11619 (N_11619,N_11523,N_11561);
or U11620 (N_11620,N_11484,N_11576);
xor U11621 (N_11621,N_11425,N_11452);
or U11622 (N_11622,N_11497,N_11448);
xnor U11623 (N_11623,N_11483,N_11567);
and U11624 (N_11624,N_11401,N_11588);
xnor U11625 (N_11625,N_11548,N_11421);
xnor U11626 (N_11626,N_11443,N_11537);
xor U11627 (N_11627,N_11566,N_11584);
nor U11628 (N_11628,N_11557,N_11469);
and U11629 (N_11629,N_11572,N_11585);
and U11630 (N_11630,N_11571,N_11597);
and U11631 (N_11631,N_11514,N_11446);
or U11632 (N_11632,N_11564,N_11599);
or U11633 (N_11633,N_11495,N_11466);
xnor U11634 (N_11634,N_11504,N_11411);
and U11635 (N_11635,N_11481,N_11476);
and U11636 (N_11636,N_11454,N_11581);
nand U11637 (N_11637,N_11436,N_11478);
nand U11638 (N_11638,N_11591,N_11474);
xnor U11639 (N_11639,N_11530,N_11580);
xor U11640 (N_11640,N_11489,N_11538);
and U11641 (N_11641,N_11574,N_11526);
and U11642 (N_11642,N_11457,N_11592);
and U11643 (N_11643,N_11499,N_11565);
nor U11644 (N_11644,N_11540,N_11455);
or U11645 (N_11645,N_11435,N_11473);
nand U11646 (N_11646,N_11440,N_11513);
and U11647 (N_11647,N_11507,N_11406);
or U11648 (N_11648,N_11451,N_11568);
or U11649 (N_11649,N_11403,N_11445);
xor U11650 (N_11650,N_11415,N_11417);
xnor U11651 (N_11651,N_11409,N_11419);
and U11652 (N_11652,N_11460,N_11553);
or U11653 (N_11653,N_11485,N_11500);
xnor U11654 (N_11654,N_11468,N_11470);
xor U11655 (N_11655,N_11432,N_11402);
nor U11656 (N_11656,N_11498,N_11458);
or U11657 (N_11657,N_11520,N_11578);
and U11658 (N_11658,N_11527,N_11467);
xor U11659 (N_11659,N_11459,N_11479);
and U11660 (N_11660,N_11444,N_11426);
nor U11661 (N_11661,N_11560,N_11477);
or U11662 (N_11662,N_11595,N_11593);
nor U11663 (N_11663,N_11472,N_11438);
and U11664 (N_11664,N_11577,N_11441);
nand U11665 (N_11665,N_11503,N_11453);
nor U11666 (N_11666,N_11594,N_11496);
xnor U11667 (N_11667,N_11545,N_11437);
nor U11668 (N_11668,N_11563,N_11586);
nor U11669 (N_11669,N_11482,N_11554);
or U11670 (N_11670,N_11541,N_11558);
nor U11671 (N_11671,N_11521,N_11547);
or U11672 (N_11672,N_11534,N_11429);
xor U11673 (N_11673,N_11493,N_11413);
nand U11674 (N_11674,N_11490,N_11405);
nand U11675 (N_11675,N_11431,N_11449);
nor U11676 (N_11676,N_11410,N_11508);
nor U11677 (N_11677,N_11549,N_11587);
xor U11678 (N_11678,N_11569,N_11434);
xnor U11679 (N_11679,N_11506,N_11494);
nor U11680 (N_11680,N_11447,N_11439);
nor U11681 (N_11681,N_11502,N_11464);
and U11682 (N_11682,N_11487,N_11582);
or U11683 (N_11683,N_11517,N_11471);
and U11684 (N_11684,N_11414,N_11462);
nor U11685 (N_11685,N_11524,N_11515);
xor U11686 (N_11686,N_11424,N_11491);
or U11687 (N_11687,N_11488,N_11529);
nand U11688 (N_11688,N_11519,N_11539);
nor U11689 (N_11689,N_11422,N_11512);
or U11690 (N_11690,N_11525,N_11559);
nand U11691 (N_11691,N_11551,N_11492);
and U11692 (N_11692,N_11418,N_11562);
and U11693 (N_11693,N_11501,N_11412);
xor U11694 (N_11694,N_11465,N_11456);
nor U11695 (N_11695,N_11509,N_11404);
or U11696 (N_11696,N_11579,N_11408);
nor U11697 (N_11697,N_11522,N_11423);
and U11698 (N_11698,N_11550,N_11532);
or U11699 (N_11699,N_11590,N_11505);
or U11700 (N_11700,N_11597,N_11456);
and U11701 (N_11701,N_11504,N_11588);
nand U11702 (N_11702,N_11578,N_11432);
nor U11703 (N_11703,N_11506,N_11400);
nor U11704 (N_11704,N_11403,N_11560);
nand U11705 (N_11705,N_11518,N_11596);
and U11706 (N_11706,N_11538,N_11453);
nand U11707 (N_11707,N_11547,N_11546);
nor U11708 (N_11708,N_11470,N_11517);
and U11709 (N_11709,N_11539,N_11403);
or U11710 (N_11710,N_11565,N_11531);
and U11711 (N_11711,N_11476,N_11509);
nor U11712 (N_11712,N_11450,N_11566);
nand U11713 (N_11713,N_11554,N_11541);
nand U11714 (N_11714,N_11483,N_11412);
xor U11715 (N_11715,N_11427,N_11516);
and U11716 (N_11716,N_11598,N_11472);
nand U11717 (N_11717,N_11454,N_11592);
and U11718 (N_11718,N_11407,N_11459);
nor U11719 (N_11719,N_11523,N_11462);
nor U11720 (N_11720,N_11458,N_11433);
and U11721 (N_11721,N_11596,N_11475);
or U11722 (N_11722,N_11582,N_11551);
nand U11723 (N_11723,N_11557,N_11527);
and U11724 (N_11724,N_11577,N_11522);
xnor U11725 (N_11725,N_11403,N_11497);
or U11726 (N_11726,N_11565,N_11550);
nand U11727 (N_11727,N_11518,N_11401);
and U11728 (N_11728,N_11462,N_11566);
nand U11729 (N_11729,N_11550,N_11507);
nor U11730 (N_11730,N_11453,N_11553);
or U11731 (N_11731,N_11495,N_11519);
and U11732 (N_11732,N_11506,N_11406);
xnor U11733 (N_11733,N_11486,N_11570);
xnor U11734 (N_11734,N_11478,N_11416);
or U11735 (N_11735,N_11422,N_11519);
nor U11736 (N_11736,N_11599,N_11440);
nand U11737 (N_11737,N_11594,N_11466);
nor U11738 (N_11738,N_11540,N_11508);
or U11739 (N_11739,N_11418,N_11570);
xnor U11740 (N_11740,N_11547,N_11425);
nand U11741 (N_11741,N_11559,N_11429);
nor U11742 (N_11742,N_11532,N_11541);
xor U11743 (N_11743,N_11499,N_11574);
or U11744 (N_11744,N_11568,N_11402);
or U11745 (N_11745,N_11598,N_11484);
and U11746 (N_11746,N_11593,N_11470);
nor U11747 (N_11747,N_11520,N_11498);
xnor U11748 (N_11748,N_11548,N_11539);
nor U11749 (N_11749,N_11549,N_11523);
nand U11750 (N_11750,N_11585,N_11426);
nor U11751 (N_11751,N_11461,N_11599);
nor U11752 (N_11752,N_11442,N_11586);
xnor U11753 (N_11753,N_11439,N_11540);
nor U11754 (N_11754,N_11436,N_11594);
nor U11755 (N_11755,N_11556,N_11578);
nor U11756 (N_11756,N_11418,N_11559);
nor U11757 (N_11757,N_11545,N_11415);
and U11758 (N_11758,N_11493,N_11506);
or U11759 (N_11759,N_11533,N_11446);
or U11760 (N_11760,N_11590,N_11462);
nand U11761 (N_11761,N_11452,N_11400);
xnor U11762 (N_11762,N_11494,N_11482);
and U11763 (N_11763,N_11450,N_11571);
xor U11764 (N_11764,N_11486,N_11454);
nand U11765 (N_11765,N_11505,N_11516);
nor U11766 (N_11766,N_11441,N_11480);
or U11767 (N_11767,N_11427,N_11559);
nand U11768 (N_11768,N_11477,N_11541);
and U11769 (N_11769,N_11475,N_11407);
nor U11770 (N_11770,N_11462,N_11451);
nand U11771 (N_11771,N_11456,N_11429);
or U11772 (N_11772,N_11450,N_11410);
and U11773 (N_11773,N_11459,N_11571);
nor U11774 (N_11774,N_11428,N_11498);
or U11775 (N_11775,N_11414,N_11486);
and U11776 (N_11776,N_11567,N_11533);
or U11777 (N_11777,N_11486,N_11494);
or U11778 (N_11778,N_11430,N_11509);
nand U11779 (N_11779,N_11556,N_11437);
nand U11780 (N_11780,N_11420,N_11479);
xor U11781 (N_11781,N_11494,N_11444);
nand U11782 (N_11782,N_11442,N_11509);
or U11783 (N_11783,N_11554,N_11461);
nand U11784 (N_11784,N_11449,N_11470);
and U11785 (N_11785,N_11475,N_11542);
nand U11786 (N_11786,N_11502,N_11536);
or U11787 (N_11787,N_11435,N_11405);
xor U11788 (N_11788,N_11518,N_11504);
and U11789 (N_11789,N_11531,N_11549);
and U11790 (N_11790,N_11567,N_11528);
nand U11791 (N_11791,N_11420,N_11424);
or U11792 (N_11792,N_11424,N_11459);
and U11793 (N_11793,N_11479,N_11515);
or U11794 (N_11794,N_11450,N_11550);
xor U11795 (N_11795,N_11407,N_11560);
nand U11796 (N_11796,N_11558,N_11507);
nand U11797 (N_11797,N_11423,N_11404);
nand U11798 (N_11798,N_11424,N_11521);
nor U11799 (N_11799,N_11499,N_11463);
xnor U11800 (N_11800,N_11770,N_11627);
or U11801 (N_11801,N_11720,N_11676);
xnor U11802 (N_11802,N_11683,N_11781);
xor U11803 (N_11803,N_11643,N_11701);
or U11804 (N_11804,N_11644,N_11746);
and U11805 (N_11805,N_11664,N_11687);
xor U11806 (N_11806,N_11740,N_11759);
xor U11807 (N_11807,N_11709,N_11622);
and U11808 (N_11808,N_11642,N_11693);
or U11809 (N_11809,N_11652,N_11714);
xor U11810 (N_11810,N_11617,N_11610);
xnor U11811 (N_11811,N_11771,N_11667);
or U11812 (N_11812,N_11707,N_11658);
nor U11813 (N_11813,N_11719,N_11711);
nand U11814 (N_11814,N_11739,N_11689);
nand U11815 (N_11815,N_11608,N_11692);
nand U11816 (N_11816,N_11737,N_11708);
nand U11817 (N_11817,N_11797,N_11705);
and U11818 (N_11818,N_11626,N_11679);
and U11819 (N_11819,N_11731,N_11744);
nand U11820 (N_11820,N_11767,N_11680);
and U11821 (N_11821,N_11764,N_11620);
and U11822 (N_11822,N_11779,N_11735);
xnor U11823 (N_11823,N_11757,N_11784);
and U11824 (N_11824,N_11745,N_11718);
and U11825 (N_11825,N_11752,N_11654);
nand U11826 (N_11826,N_11732,N_11639);
nand U11827 (N_11827,N_11619,N_11602);
xnor U11828 (N_11828,N_11756,N_11690);
nor U11829 (N_11829,N_11695,N_11754);
nand U11830 (N_11830,N_11741,N_11647);
nor U11831 (N_11831,N_11710,N_11793);
and U11832 (N_11832,N_11743,N_11789);
and U11833 (N_11833,N_11721,N_11673);
nor U11834 (N_11834,N_11645,N_11715);
xor U11835 (N_11835,N_11678,N_11691);
nor U11836 (N_11836,N_11661,N_11636);
nand U11837 (N_11837,N_11650,N_11734);
nand U11838 (N_11838,N_11663,N_11786);
xnor U11839 (N_11839,N_11641,N_11723);
or U11840 (N_11840,N_11606,N_11787);
nand U11841 (N_11841,N_11688,N_11760);
nand U11842 (N_11842,N_11726,N_11616);
nor U11843 (N_11843,N_11698,N_11765);
and U11844 (N_11844,N_11640,N_11660);
and U11845 (N_11845,N_11646,N_11727);
and U11846 (N_11846,N_11794,N_11772);
nor U11847 (N_11847,N_11677,N_11668);
xor U11848 (N_11848,N_11730,N_11628);
nand U11849 (N_11849,N_11736,N_11738);
nor U11850 (N_11850,N_11638,N_11603);
or U11851 (N_11851,N_11774,N_11799);
xor U11852 (N_11852,N_11637,N_11775);
and U11853 (N_11853,N_11750,N_11607);
nand U11854 (N_11854,N_11632,N_11666);
and U11855 (N_11855,N_11621,N_11684);
nor U11856 (N_11856,N_11623,N_11699);
nor U11857 (N_11857,N_11653,N_11725);
or U11858 (N_11858,N_11704,N_11783);
xor U11859 (N_11859,N_11696,N_11747);
or U11860 (N_11860,N_11763,N_11674);
nand U11861 (N_11861,N_11702,N_11791);
and U11862 (N_11862,N_11751,N_11713);
nor U11863 (N_11863,N_11758,N_11614);
xor U11864 (N_11864,N_11601,N_11604);
or U11865 (N_11865,N_11722,N_11755);
and U11866 (N_11866,N_11612,N_11716);
nand U11867 (N_11867,N_11670,N_11675);
nor U11868 (N_11868,N_11649,N_11686);
and U11869 (N_11869,N_11749,N_11648);
xnor U11870 (N_11870,N_11706,N_11600);
xor U11871 (N_11871,N_11631,N_11656);
nand U11872 (N_11872,N_11618,N_11768);
and U11873 (N_11873,N_11798,N_11729);
nor U11874 (N_11874,N_11717,N_11703);
nand U11875 (N_11875,N_11672,N_11624);
and U11876 (N_11876,N_11778,N_11777);
xor U11877 (N_11877,N_11682,N_11662);
xor U11878 (N_11878,N_11655,N_11659);
xnor U11879 (N_11879,N_11712,N_11796);
nor U11880 (N_11880,N_11613,N_11761);
nor U11881 (N_11881,N_11685,N_11742);
or U11882 (N_11882,N_11733,N_11776);
or U11883 (N_11883,N_11728,N_11753);
xor U11884 (N_11884,N_11615,N_11762);
nand U11885 (N_11885,N_11605,N_11780);
nor U11886 (N_11886,N_11773,N_11657);
nand U11887 (N_11887,N_11700,N_11724);
and U11888 (N_11888,N_11671,N_11782);
nor U11889 (N_11889,N_11665,N_11629);
and U11890 (N_11890,N_11635,N_11609);
nor U11891 (N_11891,N_11748,N_11694);
and U11892 (N_11892,N_11785,N_11630);
nor U11893 (N_11893,N_11633,N_11769);
nor U11894 (N_11894,N_11795,N_11697);
nand U11895 (N_11895,N_11625,N_11634);
and U11896 (N_11896,N_11766,N_11790);
and U11897 (N_11897,N_11792,N_11669);
and U11898 (N_11898,N_11651,N_11681);
nand U11899 (N_11899,N_11788,N_11611);
or U11900 (N_11900,N_11724,N_11740);
and U11901 (N_11901,N_11765,N_11773);
nor U11902 (N_11902,N_11657,N_11699);
nand U11903 (N_11903,N_11634,N_11769);
or U11904 (N_11904,N_11614,N_11757);
nor U11905 (N_11905,N_11699,N_11616);
nor U11906 (N_11906,N_11739,N_11791);
nor U11907 (N_11907,N_11764,N_11748);
or U11908 (N_11908,N_11696,N_11619);
nand U11909 (N_11909,N_11655,N_11603);
nor U11910 (N_11910,N_11668,N_11777);
nor U11911 (N_11911,N_11603,N_11663);
nor U11912 (N_11912,N_11602,N_11772);
nor U11913 (N_11913,N_11653,N_11694);
nand U11914 (N_11914,N_11687,N_11633);
nand U11915 (N_11915,N_11741,N_11775);
or U11916 (N_11916,N_11773,N_11723);
and U11917 (N_11917,N_11645,N_11630);
nor U11918 (N_11918,N_11769,N_11798);
nor U11919 (N_11919,N_11619,N_11644);
or U11920 (N_11920,N_11760,N_11752);
or U11921 (N_11921,N_11754,N_11770);
or U11922 (N_11922,N_11739,N_11610);
and U11923 (N_11923,N_11782,N_11770);
nor U11924 (N_11924,N_11654,N_11765);
and U11925 (N_11925,N_11707,N_11769);
and U11926 (N_11926,N_11661,N_11787);
and U11927 (N_11927,N_11796,N_11606);
and U11928 (N_11928,N_11798,N_11735);
and U11929 (N_11929,N_11614,N_11743);
xor U11930 (N_11930,N_11671,N_11664);
nor U11931 (N_11931,N_11667,N_11637);
or U11932 (N_11932,N_11653,N_11671);
or U11933 (N_11933,N_11706,N_11707);
nand U11934 (N_11934,N_11688,N_11719);
nand U11935 (N_11935,N_11796,N_11797);
or U11936 (N_11936,N_11743,N_11663);
xnor U11937 (N_11937,N_11673,N_11649);
xor U11938 (N_11938,N_11657,N_11658);
and U11939 (N_11939,N_11682,N_11781);
xor U11940 (N_11940,N_11728,N_11682);
and U11941 (N_11941,N_11697,N_11676);
xnor U11942 (N_11942,N_11781,N_11654);
and U11943 (N_11943,N_11672,N_11710);
nand U11944 (N_11944,N_11749,N_11782);
nand U11945 (N_11945,N_11738,N_11778);
and U11946 (N_11946,N_11708,N_11634);
and U11947 (N_11947,N_11778,N_11769);
nor U11948 (N_11948,N_11621,N_11795);
nor U11949 (N_11949,N_11754,N_11783);
nand U11950 (N_11950,N_11615,N_11634);
and U11951 (N_11951,N_11611,N_11669);
nor U11952 (N_11952,N_11682,N_11738);
nand U11953 (N_11953,N_11784,N_11701);
or U11954 (N_11954,N_11659,N_11646);
nor U11955 (N_11955,N_11652,N_11621);
nand U11956 (N_11956,N_11750,N_11777);
and U11957 (N_11957,N_11775,N_11679);
nand U11958 (N_11958,N_11648,N_11720);
nand U11959 (N_11959,N_11773,N_11754);
and U11960 (N_11960,N_11762,N_11629);
nand U11961 (N_11961,N_11718,N_11730);
nand U11962 (N_11962,N_11757,N_11723);
or U11963 (N_11963,N_11750,N_11763);
xor U11964 (N_11964,N_11643,N_11736);
nand U11965 (N_11965,N_11710,N_11703);
nand U11966 (N_11966,N_11722,N_11764);
xor U11967 (N_11967,N_11618,N_11774);
and U11968 (N_11968,N_11654,N_11690);
or U11969 (N_11969,N_11657,N_11647);
xnor U11970 (N_11970,N_11706,N_11724);
and U11971 (N_11971,N_11737,N_11694);
or U11972 (N_11972,N_11605,N_11607);
and U11973 (N_11973,N_11790,N_11777);
xnor U11974 (N_11974,N_11733,N_11735);
nor U11975 (N_11975,N_11661,N_11670);
and U11976 (N_11976,N_11607,N_11718);
and U11977 (N_11977,N_11723,N_11737);
xor U11978 (N_11978,N_11689,N_11652);
nor U11979 (N_11979,N_11772,N_11606);
and U11980 (N_11980,N_11694,N_11660);
and U11981 (N_11981,N_11634,N_11603);
xnor U11982 (N_11982,N_11772,N_11678);
nand U11983 (N_11983,N_11659,N_11662);
nand U11984 (N_11984,N_11781,N_11634);
and U11985 (N_11985,N_11784,N_11712);
and U11986 (N_11986,N_11628,N_11715);
nor U11987 (N_11987,N_11771,N_11706);
xor U11988 (N_11988,N_11686,N_11713);
nor U11989 (N_11989,N_11603,N_11770);
nand U11990 (N_11990,N_11712,N_11738);
or U11991 (N_11991,N_11731,N_11689);
or U11992 (N_11992,N_11774,N_11680);
nor U11993 (N_11993,N_11718,N_11754);
and U11994 (N_11994,N_11660,N_11726);
and U11995 (N_11995,N_11721,N_11777);
xnor U11996 (N_11996,N_11778,N_11675);
xor U11997 (N_11997,N_11654,N_11615);
or U11998 (N_11998,N_11663,N_11604);
nor U11999 (N_11999,N_11638,N_11724);
xor U12000 (N_12000,N_11882,N_11870);
nor U12001 (N_12001,N_11972,N_11811);
and U12002 (N_12002,N_11874,N_11981);
xor U12003 (N_12003,N_11852,N_11839);
or U12004 (N_12004,N_11909,N_11939);
nand U12005 (N_12005,N_11830,N_11840);
nor U12006 (N_12006,N_11866,N_11897);
xnor U12007 (N_12007,N_11846,N_11932);
or U12008 (N_12008,N_11979,N_11957);
xnor U12009 (N_12009,N_11994,N_11851);
and U12010 (N_12010,N_11956,N_11809);
or U12011 (N_12011,N_11969,N_11944);
xnor U12012 (N_12012,N_11964,N_11893);
and U12013 (N_12013,N_11857,N_11919);
nand U12014 (N_12014,N_11875,N_11843);
xor U12015 (N_12015,N_11829,N_11982);
nor U12016 (N_12016,N_11966,N_11959);
xor U12017 (N_12017,N_11947,N_11825);
nor U12018 (N_12018,N_11847,N_11824);
or U12019 (N_12019,N_11978,N_11810);
nand U12020 (N_12020,N_11987,N_11918);
and U12021 (N_12021,N_11908,N_11968);
nor U12022 (N_12022,N_11802,N_11855);
nand U12023 (N_12023,N_11949,N_11807);
nand U12024 (N_12024,N_11928,N_11996);
and U12025 (N_12025,N_11877,N_11826);
nor U12026 (N_12026,N_11817,N_11806);
or U12027 (N_12027,N_11936,N_11833);
or U12028 (N_12028,N_11962,N_11838);
nand U12029 (N_12029,N_11813,N_11886);
and U12030 (N_12030,N_11803,N_11940);
and U12031 (N_12031,N_11894,N_11812);
xor U12032 (N_12032,N_11864,N_11960);
nor U12033 (N_12033,N_11902,N_11845);
or U12034 (N_12034,N_11848,N_11863);
and U12035 (N_12035,N_11973,N_11819);
nand U12036 (N_12036,N_11827,N_11943);
and U12037 (N_12037,N_11834,N_11977);
or U12038 (N_12038,N_11991,N_11913);
nand U12039 (N_12039,N_11879,N_11873);
nor U12040 (N_12040,N_11999,N_11917);
and U12041 (N_12041,N_11853,N_11974);
nand U12042 (N_12042,N_11976,N_11841);
xnor U12043 (N_12043,N_11872,N_11849);
nor U12044 (N_12044,N_11912,N_11905);
or U12045 (N_12045,N_11896,N_11860);
nor U12046 (N_12046,N_11998,N_11980);
or U12047 (N_12047,N_11821,N_11859);
xnor U12048 (N_12048,N_11921,N_11814);
nand U12049 (N_12049,N_11970,N_11800);
nand U12050 (N_12050,N_11881,N_11923);
nand U12051 (N_12051,N_11891,N_11836);
or U12052 (N_12052,N_11942,N_11946);
or U12053 (N_12053,N_11967,N_11871);
nand U12054 (N_12054,N_11804,N_11892);
or U12055 (N_12055,N_11945,N_11832);
or U12056 (N_12056,N_11883,N_11861);
xnor U12057 (N_12057,N_11869,N_11941);
nor U12058 (N_12058,N_11805,N_11822);
or U12059 (N_12059,N_11951,N_11900);
xnor U12060 (N_12060,N_11895,N_11914);
and U12061 (N_12061,N_11925,N_11990);
or U12062 (N_12062,N_11961,N_11911);
and U12063 (N_12063,N_11837,N_11818);
nand U12064 (N_12064,N_11801,N_11898);
nand U12065 (N_12065,N_11868,N_11971);
nor U12066 (N_12066,N_11828,N_11955);
and U12067 (N_12067,N_11835,N_11816);
or U12068 (N_12068,N_11885,N_11988);
nand U12069 (N_12069,N_11878,N_11820);
nand U12070 (N_12070,N_11986,N_11953);
nor U12071 (N_12071,N_11850,N_11856);
xor U12072 (N_12072,N_11862,N_11889);
xor U12073 (N_12073,N_11933,N_11992);
nor U12074 (N_12074,N_11906,N_11931);
or U12075 (N_12075,N_11984,N_11950);
and U12076 (N_12076,N_11926,N_11983);
or U12077 (N_12077,N_11920,N_11948);
and U12078 (N_12078,N_11915,N_11995);
nor U12079 (N_12079,N_11930,N_11901);
nor U12080 (N_12080,N_11985,N_11899);
nor U12081 (N_12081,N_11937,N_11842);
nor U12082 (N_12082,N_11934,N_11993);
nor U12083 (N_12083,N_11904,N_11867);
nand U12084 (N_12084,N_11887,N_11929);
xnor U12085 (N_12085,N_11922,N_11815);
and U12086 (N_12086,N_11858,N_11958);
nor U12087 (N_12087,N_11924,N_11997);
xnor U12088 (N_12088,N_11954,N_11938);
and U12089 (N_12089,N_11989,N_11927);
or U12090 (N_12090,N_11880,N_11884);
xor U12091 (N_12091,N_11876,N_11903);
and U12092 (N_12092,N_11910,N_11865);
or U12093 (N_12093,N_11952,N_11888);
nor U12094 (N_12094,N_11963,N_11935);
and U12095 (N_12095,N_11808,N_11890);
xor U12096 (N_12096,N_11965,N_11823);
and U12097 (N_12097,N_11854,N_11975);
nor U12098 (N_12098,N_11907,N_11916);
and U12099 (N_12099,N_11831,N_11844);
or U12100 (N_12100,N_11872,N_11889);
xor U12101 (N_12101,N_11951,N_11835);
xnor U12102 (N_12102,N_11804,N_11829);
nand U12103 (N_12103,N_11995,N_11830);
xor U12104 (N_12104,N_11891,N_11911);
and U12105 (N_12105,N_11915,N_11994);
or U12106 (N_12106,N_11863,N_11908);
and U12107 (N_12107,N_11902,N_11890);
nand U12108 (N_12108,N_11991,N_11892);
nor U12109 (N_12109,N_11948,N_11941);
nor U12110 (N_12110,N_11865,N_11832);
and U12111 (N_12111,N_11911,N_11852);
nand U12112 (N_12112,N_11949,N_11904);
or U12113 (N_12113,N_11933,N_11962);
nor U12114 (N_12114,N_11947,N_11927);
xor U12115 (N_12115,N_11880,N_11914);
xor U12116 (N_12116,N_11849,N_11918);
or U12117 (N_12117,N_11948,N_11968);
and U12118 (N_12118,N_11808,N_11969);
or U12119 (N_12119,N_11869,N_11969);
nand U12120 (N_12120,N_11910,N_11862);
xor U12121 (N_12121,N_11960,N_11977);
nor U12122 (N_12122,N_11824,N_11905);
and U12123 (N_12123,N_11908,N_11956);
nand U12124 (N_12124,N_11818,N_11893);
nor U12125 (N_12125,N_11852,N_11851);
and U12126 (N_12126,N_11803,N_11992);
nor U12127 (N_12127,N_11995,N_11911);
nor U12128 (N_12128,N_11922,N_11824);
xor U12129 (N_12129,N_11814,N_11922);
and U12130 (N_12130,N_11823,N_11977);
nand U12131 (N_12131,N_11961,N_11904);
and U12132 (N_12132,N_11880,N_11970);
or U12133 (N_12133,N_11999,N_11913);
or U12134 (N_12134,N_11865,N_11984);
xor U12135 (N_12135,N_11870,N_11836);
nor U12136 (N_12136,N_11992,N_11804);
nand U12137 (N_12137,N_11981,N_11830);
xor U12138 (N_12138,N_11830,N_11860);
nand U12139 (N_12139,N_11895,N_11913);
nand U12140 (N_12140,N_11959,N_11961);
nand U12141 (N_12141,N_11913,N_11938);
or U12142 (N_12142,N_11969,N_11907);
nor U12143 (N_12143,N_11947,N_11938);
xnor U12144 (N_12144,N_11908,N_11880);
and U12145 (N_12145,N_11986,N_11895);
nand U12146 (N_12146,N_11814,N_11956);
nor U12147 (N_12147,N_11923,N_11987);
nor U12148 (N_12148,N_11938,N_11830);
nand U12149 (N_12149,N_11913,N_11879);
or U12150 (N_12150,N_11971,N_11836);
nor U12151 (N_12151,N_11819,N_11879);
and U12152 (N_12152,N_11814,N_11942);
and U12153 (N_12153,N_11835,N_11945);
or U12154 (N_12154,N_11808,N_11907);
nand U12155 (N_12155,N_11890,N_11887);
or U12156 (N_12156,N_11892,N_11924);
nand U12157 (N_12157,N_11933,N_11939);
xor U12158 (N_12158,N_11942,N_11850);
nand U12159 (N_12159,N_11949,N_11939);
xor U12160 (N_12160,N_11957,N_11838);
nand U12161 (N_12161,N_11845,N_11953);
nor U12162 (N_12162,N_11886,N_11956);
nand U12163 (N_12163,N_11819,N_11803);
nor U12164 (N_12164,N_11855,N_11962);
or U12165 (N_12165,N_11875,N_11959);
nand U12166 (N_12166,N_11808,N_11926);
xor U12167 (N_12167,N_11890,N_11850);
or U12168 (N_12168,N_11824,N_11814);
or U12169 (N_12169,N_11893,N_11993);
nand U12170 (N_12170,N_11992,N_11844);
nand U12171 (N_12171,N_11953,N_11891);
nand U12172 (N_12172,N_11934,N_11992);
nand U12173 (N_12173,N_11974,N_11870);
or U12174 (N_12174,N_11924,N_11869);
or U12175 (N_12175,N_11876,N_11803);
xor U12176 (N_12176,N_11950,N_11914);
xor U12177 (N_12177,N_11911,N_11834);
xnor U12178 (N_12178,N_11975,N_11871);
or U12179 (N_12179,N_11927,N_11952);
xnor U12180 (N_12180,N_11819,N_11831);
nand U12181 (N_12181,N_11921,N_11916);
or U12182 (N_12182,N_11987,N_11824);
xnor U12183 (N_12183,N_11937,N_11873);
xnor U12184 (N_12184,N_11897,N_11873);
nor U12185 (N_12185,N_11940,N_11959);
or U12186 (N_12186,N_11889,N_11833);
and U12187 (N_12187,N_11880,N_11992);
nor U12188 (N_12188,N_11919,N_11972);
and U12189 (N_12189,N_11853,N_11926);
nor U12190 (N_12190,N_11838,N_11826);
or U12191 (N_12191,N_11957,N_11988);
nand U12192 (N_12192,N_11942,N_11955);
and U12193 (N_12193,N_11858,N_11982);
and U12194 (N_12194,N_11953,N_11824);
xnor U12195 (N_12195,N_11958,N_11971);
nand U12196 (N_12196,N_11857,N_11986);
nand U12197 (N_12197,N_11925,N_11946);
nand U12198 (N_12198,N_11829,N_11929);
nand U12199 (N_12199,N_11910,N_11844);
and U12200 (N_12200,N_12011,N_12197);
xnor U12201 (N_12201,N_12038,N_12067);
nor U12202 (N_12202,N_12078,N_12185);
xnor U12203 (N_12203,N_12192,N_12088);
nand U12204 (N_12204,N_12033,N_12083);
or U12205 (N_12205,N_12095,N_12027);
and U12206 (N_12206,N_12111,N_12056);
or U12207 (N_12207,N_12004,N_12184);
or U12208 (N_12208,N_12124,N_12041);
or U12209 (N_12209,N_12163,N_12016);
nor U12210 (N_12210,N_12122,N_12049);
xnor U12211 (N_12211,N_12058,N_12189);
nor U12212 (N_12212,N_12107,N_12164);
nor U12213 (N_12213,N_12132,N_12128);
xnor U12214 (N_12214,N_12142,N_12134);
and U12215 (N_12215,N_12026,N_12168);
or U12216 (N_12216,N_12172,N_12195);
xor U12217 (N_12217,N_12141,N_12113);
or U12218 (N_12218,N_12025,N_12008);
nand U12219 (N_12219,N_12007,N_12069);
or U12220 (N_12220,N_12152,N_12100);
nand U12221 (N_12221,N_12166,N_12047);
or U12222 (N_12222,N_12042,N_12193);
nand U12223 (N_12223,N_12061,N_12138);
or U12224 (N_12224,N_12074,N_12179);
or U12225 (N_12225,N_12029,N_12148);
xnor U12226 (N_12226,N_12040,N_12043);
nand U12227 (N_12227,N_12009,N_12190);
nor U12228 (N_12228,N_12050,N_12120);
nand U12229 (N_12229,N_12096,N_12054);
or U12230 (N_12230,N_12196,N_12114);
nand U12231 (N_12231,N_12112,N_12020);
xnor U12232 (N_12232,N_12115,N_12015);
and U12233 (N_12233,N_12139,N_12045);
nor U12234 (N_12234,N_12109,N_12019);
or U12235 (N_12235,N_12167,N_12079);
and U12236 (N_12236,N_12121,N_12082);
xnor U12237 (N_12237,N_12046,N_12071);
nand U12238 (N_12238,N_12104,N_12003);
xor U12239 (N_12239,N_12017,N_12191);
xnor U12240 (N_12240,N_12145,N_12123);
and U12241 (N_12241,N_12080,N_12144);
or U12242 (N_12242,N_12024,N_12186);
nor U12243 (N_12243,N_12102,N_12028);
and U12244 (N_12244,N_12014,N_12076);
and U12245 (N_12245,N_12089,N_12064);
and U12246 (N_12246,N_12063,N_12156);
and U12247 (N_12247,N_12002,N_12133);
nor U12248 (N_12248,N_12087,N_12012);
and U12249 (N_12249,N_12086,N_12177);
xnor U12250 (N_12250,N_12098,N_12155);
nor U12251 (N_12251,N_12188,N_12117);
and U12252 (N_12252,N_12062,N_12022);
or U12253 (N_12253,N_12093,N_12146);
xor U12254 (N_12254,N_12131,N_12034);
and U12255 (N_12255,N_12199,N_12037);
or U12256 (N_12256,N_12053,N_12182);
nand U12257 (N_12257,N_12090,N_12073);
nor U12258 (N_12258,N_12052,N_12092);
nand U12259 (N_12259,N_12165,N_12000);
nand U12260 (N_12260,N_12118,N_12103);
nor U12261 (N_12261,N_12175,N_12187);
nand U12262 (N_12262,N_12181,N_12178);
xnor U12263 (N_12263,N_12159,N_12072);
nor U12264 (N_12264,N_12055,N_12105);
nor U12265 (N_12265,N_12057,N_12085);
xor U12266 (N_12266,N_12035,N_12161);
nor U12267 (N_12267,N_12154,N_12001);
nand U12268 (N_12268,N_12048,N_12180);
nor U12269 (N_12269,N_12110,N_12130);
xor U12270 (N_12270,N_12070,N_12030);
or U12271 (N_12271,N_12068,N_12006);
xnor U12272 (N_12272,N_12174,N_12171);
nand U12273 (N_12273,N_12127,N_12066);
nor U12274 (N_12274,N_12116,N_12099);
and U12275 (N_12275,N_12143,N_12084);
nand U12276 (N_12276,N_12091,N_12198);
or U12277 (N_12277,N_12169,N_12135);
or U12278 (N_12278,N_12039,N_12108);
or U12279 (N_12279,N_12097,N_12136);
and U12280 (N_12280,N_12137,N_12129);
nand U12281 (N_12281,N_12051,N_12183);
xor U12282 (N_12282,N_12150,N_12101);
and U12283 (N_12283,N_12125,N_12036);
nor U12284 (N_12284,N_12065,N_12158);
nand U12285 (N_12285,N_12031,N_12106);
or U12286 (N_12286,N_12021,N_12149);
nor U12287 (N_12287,N_12094,N_12160);
nand U12288 (N_12288,N_12010,N_12075);
and U12289 (N_12289,N_12157,N_12153);
and U12290 (N_12290,N_12151,N_12140);
and U12291 (N_12291,N_12176,N_12194);
and U12292 (N_12292,N_12173,N_12162);
nand U12293 (N_12293,N_12077,N_12044);
or U12294 (N_12294,N_12147,N_12032);
xnor U12295 (N_12295,N_12060,N_12170);
nor U12296 (N_12296,N_12119,N_12081);
or U12297 (N_12297,N_12013,N_12059);
xnor U12298 (N_12298,N_12126,N_12005);
and U12299 (N_12299,N_12018,N_12023);
nand U12300 (N_12300,N_12023,N_12070);
nand U12301 (N_12301,N_12168,N_12102);
nand U12302 (N_12302,N_12033,N_12104);
nand U12303 (N_12303,N_12070,N_12176);
xor U12304 (N_12304,N_12065,N_12057);
nand U12305 (N_12305,N_12186,N_12153);
and U12306 (N_12306,N_12174,N_12195);
xnor U12307 (N_12307,N_12098,N_12118);
xnor U12308 (N_12308,N_12154,N_12028);
xnor U12309 (N_12309,N_12072,N_12107);
xor U12310 (N_12310,N_12190,N_12079);
and U12311 (N_12311,N_12022,N_12046);
and U12312 (N_12312,N_12058,N_12164);
or U12313 (N_12313,N_12082,N_12164);
and U12314 (N_12314,N_12109,N_12171);
nand U12315 (N_12315,N_12133,N_12081);
or U12316 (N_12316,N_12073,N_12109);
nand U12317 (N_12317,N_12044,N_12184);
and U12318 (N_12318,N_12183,N_12149);
nand U12319 (N_12319,N_12024,N_12125);
nand U12320 (N_12320,N_12033,N_12064);
nand U12321 (N_12321,N_12032,N_12130);
xor U12322 (N_12322,N_12145,N_12090);
xor U12323 (N_12323,N_12154,N_12073);
nor U12324 (N_12324,N_12125,N_12105);
or U12325 (N_12325,N_12113,N_12075);
nand U12326 (N_12326,N_12124,N_12167);
nand U12327 (N_12327,N_12106,N_12100);
xor U12328 (N_12328,N_12073,N_12020);
and U12329 (N_12329,N_12078,N_12108);
and U12330 (N_12330,N_12059,N_12041);
nand U12331 (N_12331,N_12070,N_12147);
xnor U12332 (N_12332,N_12128,N_12199);
or U12333 (N_12333,N_12137,N_12088);
or U12334 (N_12334,N_12003,N_12183);
xnor U12335 (N_12335,N_12141,N_12142);
nand U12336 (N_12336,N_12193,N_12108);
and U12337 (N_12337,N_12103,N_12094);
or U12338 (N_12338,N_12003,N_12016);
nor U12339 (N_12339,N_12035,N_12197);
or U12340 (N_12340,N_12128,N_12021);
and U12341 (N_12341,N_12168,N_12195);
or U12342 (N_12342,N_12037,N_12097);
nand U12343 (N_12343,N_12149,N_12165);
and U12344 (N_12344,N_12199,N_12027);
and U12345 (N_12345,N_12103,N_12097);
nor U12346 (N_12346,N_12049,N_12157);
xor U12347 (N_12347,N_12009,N_12047);
or U12348 (N_12348,N_12148,N_12072);
and U12349 (N_12349,N_12013,N_12140);
and U12350 (N_12350,N_12180,N_12147);
nand U12351 (N_12351,N_12110,N_12013);
and U12352 (N_12352,N_12168,N_12097);
or U12353 (N_12353,N_12186,N_12127);
or U12354 (N_12354,N_12064,N_12184);
nand U12355 (N_12355,N_12054,N_12030);
xor U12356 (N_12356,N_12060,N_12022);
nor U12357 (N_12357,N_12049,N_12146);
or U12358 (N_12358,N_12124,N_12088);
nor U12359 (N_12359,N_12196,N_12079);
and U12360 (N_12360,N_12000,N_12008);
or U12361 (N_12361,N_12075,N_12085);
xnor U12362 (N_12362,N_12186,N_12137);
xnor U12363 (N_12363,N_12019,N_12032);
xor U12364 (N_12364,N_12133,N_12050);
and U12365 (N_12365,N_12098,N_12179);
nor U12366 (N_12366,N_12028,N_12031);
nor U12367 (N_12367,N_12159,N_12145);
nand U12368 (N_12368,N_12010,N_12171);
and U12369 (N_12369,N_12031,N_12183);
nor U12370 (N_12370,N_12181,N_12005);
and U12371 (N_12371,N_12065,N_12191);
nor U12372 (N_12372,N_12069,N_12053);
xnor U12373 (N_12373,N_12037,N_12047);
nand U12374 (N_12374,N_12021,N_12108);
nand U12375 (N_12375,N_12048,N_12172);
xor U12376 (N_12376,N_12152,N_12000);
and U12377 (N_12377,N_12024,N_12068);
nor U12378 (N_12378,N_12023,N_12099);
nor U12379 (N_12379,N_12047,N_12181);
or U12380 (N_12380,N_12167,N_12160);
or U12381 (N_12381,N_12106,N_12167);
and U12382 (N_12382,N_12124,N_12101);
or U12383 (N_12383,N_12085,N_12158);
xnor U12384 (N_12384,N_12064,N_12139);
and U12385 (N_12385,N_12053,N_12036);
or U12386 (N_12386,N_12162,N_12091);
nor U12387 (N_12387,N_12041,N_12092);
or U12388 (N_12388,N_12003,N_12195);
or U12389 (N_12389,N_12177,N_12172);
xnor U12390 (N_12390,N_12100,N_12109);
nor U12391 (N_12391,N_12109,N_12000);
xnor U12392 (N_12392,N_12116,N_12035);
nor U12393 (N_12393,N_12023,N_12054);
or U12394 (N_12394,N_12007,N_12142);
nand U12395 (N_12395,N_12172,N_12128);
or U12396 (N_12396,N_12065,N_12000);
or U12397 (N_12397,N_12146,N_12055);
xor U12398 (N_12398,N_12194,N_12192);
nor U12399 (N_12399,N_12094,N_12176);
nand U12400 (N_12400,N_12257,N_12327);
or U12401 (N_12401,N_12256,N_12361);
and U12402 (N_12402,N_12241,N_12334);
or U12403 (N_12403,N_12397,N_12291);
or U12404 (N_12404,N_12212,N_12399);
xnor U12405 (N_12405,N_12236,N_12274);
or U12406 (N_12406,N_12218,N_12366);
xor U12407 (N_12407,N_12379,N_12322);
and U12408 (N_12408,N_12223,N_12333);
xor U12409 (N_12409,N_12297,N_12266);
and U12410 (N_12410,N_12205,N_12395);
and U12411 (N_12411,N_12341,N_12259);
xnor U12412 (N_12412,N_12295,N_12306);
xor U12413 (N_12413,N_12261,N_12237);
nand U12414 (N_12414,N_12359,N_12284);
nand U12415 (N_12415,N_12302,N_12340);
or U12416 (N_12416,N_12367,N_12248);
xor U12417 (N_12417,N_12381,N_12390);
nand U12418 (N_12418,N_12326,N_12225);
and U12419 (N_12419,N_12254,N_12283);
nand U12420 (N_12420,N_12324,N_12290);
and U12421 (N_12421,N_12272,N_12364);
xnor U12422 (N_12422,N_12385,N_12353);
xnor U12423 (N_12423,N_12360,N_12298);
or U12424 (N_12424,N_12378,N_12255);
nand U12425 (N_12425,N_12380,N_12240);
or U12426 (N_12426,N_12300,N_12200);
or U12427 (N_12427,N_12271,N_12214);
or U12428 (N_12428,N_12228,N_12277);
xnor U12429 (N_12429,N_12211,N_12202);
nand U12430 (N_12430,N_12346,N_12219);
nand U12431 (N_12431,N_12321,N_12229);
xnor U12432 (N_12432,N_12313,N_12258);
nand U12433 (N_12433,N_12316,N_12392);
and U12434 (N_12434,N_12250,N_12233);
or U12435 (N_12435,N_12285,N_12263);
xor U12436 (N_12436,N_12294,N_12239);
or U12437 (N_12437,N_12351,N_12207);
nand U12438 (N_12438,N_12282,N_12309);
nor U12439 (N_12439,N_12269,N_12244);
nor U12440 (N_12440,N_12349,N_12374);
nor U12441 (N_12441,N_12227,N_12221);
xnor U12442 (N_12442,N_12220,N_12330);
nand U12443 (N_12443,N_12368,N_12301);
or U12444 (N_12444,N_12362,N_12230);
nand U12445 (N_12445,N_12387,N_12216);
xnor U12446 (N_12446,N_12339,N_12396);
xor U12447 (N_12447,N_12231,N_12311);
and U12448 (N_12448,N_12264,N_12356);
and U12449 (N_12449,N_12312,N_12235);
or U12450 (N_12450,N_12296,N_12344);
nand U12451 (N_12451,N_12304,N_12391);
and U12452 (N_12452,N_12210,N_12206);
nor U12453 (N_12453,N_12224,N_12208);
nand U12454 (N_12454,N_12347,N_12292);
xnor U12455 (N_12455,N_12232,N_12310);
nor U12456 (N_12456,N_12281,N_12343);
nand U12457 (N_12457,N_12345,N_12315);
xnor U12458 (N_12458,N_12245,N_12319);
nor U12459 (N_12459,N_12222,N_12242);
and U12460 (N_12460,N_12372,N_12377);
or U12461 (N_12461,N_12398,N_12260);
nand U12462 (N_12462,N_12249,N_12273);
nand U12463 (N_12463,N_12358,N_12363);
and U12464 (N_12464,N_12252,N_12215);
nand U12465 (N_12465,N_12371,N_12338);
xnor U12466 (N_12466,N_12203,N_12288);
and U12467 (N_12467,N_12251,N_12267);
and U12468 (N_12468,N_12342,N_12328);
or U12469 (N_12469,N_12299,N_12376);
or U12470 (N_12470,N_12307,N_12365);
or U12471 (N_12471,N_12355,N_12384);
and U12472 (N_12472,N_12280,N_12201);
or U12473 (N_12473,N_12348,N_12383);
xor U12474 (N_12474,N_12352,N_12308);
nor U12475 (N_12475,N_12388,N_12331);
or U12476 (N_12476,N_12279,N_12293);
and U12477 (N_12477,N_12350,N_12253);
nand U12478 (N_12478,N_12394,N_12289);
nor U12479 (N_12479,N_12234,N_12204);
and U12480 (N_12480,N_12317,N_12209);
nand U12481 (N_12481,N_12323,N_12275);
nor U12482 (N_12482,N_12329,N_12354);
and U12483 (N_12483,N_12238,N_12213);
nand U12484 (N_12484,N_12393,N_12336);
and U12485 (N_12485,N_12373,N_12270);
or U12486 (N_12486,N_12369,N_12303);
and U12487 (N_12487,N_12386,N_12335);
xor U12488 (N_12488,N_12382,N_12286);
nand U12489 (N_12489,N_12337,N_12268);
xor U12490 (N_12490,N_12357,N_12217);
and U12491 (N_12491,N_12325,N_12389);
nand U12492 (N_12492,N_12226,N_12332);
or U12493 (N_12493,N_12243,N_12320);
nand U12494 (N_12494,N_12318,N_12278);
and U12495 (N_12495,N_12247,N_12276);
nor U12496 (N_12496,N_12287,N_12314);
or U12497 (N_12497,N_12262,N_12265);
or U12498 (N_12498,N_12246,N_12305);
or U12499 (N_12499,N_12375,N_12370);
nand U12500 (N_12500,N_12303,N_12306);
nor U12501 (N_12501,N_12272,N_12258);
nand U12502 (N_12502,N_12262,N_12303);
nand U12503 (N_12503,N_12302,N_12285);
xor U12504 (N_12504,N_12329,N_12219);
and U12505 (N_12505,N_12264,N_12312);
nor U12506 (N_12506,N_12211,N_12330);
or U12507 (N_12507,N_12206,N_12397);
nor U12508 (N_12508,N_12322,N_12303);
nor U12509 (N_12509,N_12257,N_12344);
nor U12510 (N_12510,N_12380,N_12302);
nor U12511 (N_12511,N_12220,N_12265);
and U12512 (N_12512,N_12258,N_12276);
nor U12513 (N_12513,N_12241,N_12336);
or U12514 (N_12514,N_12318,N_12367);
nand U12515 (N_12515,N_12363,N_12380);
or U12516 (N_12516,N_12339,N_12309);
or U12517 (N_12517,N_12396,N_12299);
xor U12518 (N_12518,N_12229,N_12339);
nand U12519 (N_12519,N_12268,N_12343);
or U12520 (N_12520,N_12229,N_12385);
and U12521 (N_12521,N_12315,N_12281);
or U12522 (N_12522,N_12241,N_12259);
or U12523 (N_12523,N_12261,N_12297);
nand U12524 (N_12524,N_12361,N_12232);
or U12525 (N_12525,N_12299,N_12342);
or U12526 (N_12526,N_12325,N_12217);
nand U12527 (N_12527,N_12212,N_12247);
xor U12528 (N_12528,N_12285,N_12222);
xnor U12529 (N_12529,N_12246,N_12285);
nand U12530 (N_12530,N_12377,N_12243);
xor U12531 (N_12531,N_12226,N_12364);
xor U12532 (N_12532,N_12212,N_12286);
nor U12533 (N_12533,N_12247,N_12354);
or U12534 (N_12534,N_12391,N_12292);
xor U12535 (N_12535,N_12364,N_12247);
or U12536 (N_12536,N_12297,N_12288);
nand U12537 (N_12537,N_12328,N_12216);
nor U12538 (N_12538,N_12396,N_12366);
nor U12539 (N_12539,N_12302,N_12252);
xor U12540 (N_12540,N_12248,N_12259);
nand U12541 (N_12541,N_12268,N_12316);
and U12542 (N_12542,N_12392,N_12246);
xnor U12543 (N_12543,N_12250,N_12205);
nand U12544 (N_12544,N_12304,N_12255);
nand U12545 (N_12545,N_12345,N_12304);
nand U12546 (N_12546,N_12210,N_12266);
nor U12547 (N_12547,N_12231,N_12387);
xnor U12548 (N_12548,N_12323,N_12341);
and U12549 (N_12549,N_12373,N_12252);
nor U12550 (N_12550,N_12225,N_12366);
and U12551 (N_12551,N_12223,N_12315);
and U12552 (N_12552,N_12294,N_12275);
or U12553 (N_12553,N_12352,N_12236);
and U12554 (N_12554,N_12245,N_12239);
xnor U12555 (N_12555,N_12236,N_12373);
nand U12556 (N_12556,N_12365,N_12227);
and U12557 (N_12557,N_12356,N_12376);
nor U12558 (N_12558,N_12370,N_12309);
xnor U12559 (N_12559,N_12227,N_12206);
nor U12560 (N_12560,N_12251,N_12278);
xnor U12561 (N_12561,N_12272,N_12357);
and U12562 (N_12562,N_12390,N_12219);
nand U12563 (N_12563,N_12220,N_12389);
nor U12564 (N_12564,N_12394,N_12357);
and U12565 (N_12565,N_12260,N_12351);
xor U12566 (N_12566,N_12281,N_12231);
and U12567 (N_12567,N_12229,N_12388);
xnor U12568 (N_12568,N_12219,N_12393);
nor U12569 (N_12569,N_12383,N_12339);
nor U12570 (N_12570,N_12241,N_12305);
nand U12571 (N_12571,N_12256,N_12212);
or U12572 (N_12572,N_12357,N_12265);
and U12573 (N_12573,N_12282,N_12211);
nand U12574 (N_12574,N_12230,N_12295);
and U12575 (N_12575,N_12396,N_12282);
xor U12576 (N_12576,N_12384,N_12374);
nand U12577 (N_12577,N_12276,N_12342);
nand U12578 (N_12578,N_12354,N_12288);
and U12579 (N_12579,N_12341,N_12290);
and U12580 (N_12580,N_12219,N_12387);
nand U12581 (N_12581,N_12377,N_12230);
or U12582 (N_12582,N_12317,N_12281);
xnor U12583 (N_12583,N_12369,N_12266);
nand U12584 (N_12584,N_12384,N_12243);
or U12585 (N_12585,N_12398,N_12287);
nand U12586 (N_12586,N_12277,N_12345);
or U12587 (N_12587,N_12288,N_12338);
xnor U12588 (N_12588,N_12397,N_12332);
nand U12589 (N_12589,N_12372,N_12285);
nand U12590 (N_12590,N_12209,N_12278);
or U12591 (N_12591,N_12361,N_12289);
nor U12592 (N_12592,N_12399,N_12228);
xnor U12593 (N_12593,N_12255,N_12375);
nand U12594 (N_12594,N_12278,N_12236);
nor U12595 (N_12595,N_12301,N_12282);
xor U12596 (N_12596,N_12331,N_12316);
nor U12597 (N_12597,N_12230,N_12348);
nand U12598 (N_12598,N_12338,N_12277);
nor U12599 (N_12599,N_12361,N_12307);
or U12600 (N_12600,N_12522,N_12526);
and U12601 (N_12601,N_12439,N_12514);
xor U12602 (N_12602,N_12469,N_12585);
and U12603 (N_12603,N_12550,N_12472);
and U12604 (N_12604,N_12404,N_12494);
nor U12605 (N_12605,N_12425,N_12403);
and U12606 (N_12606,N_12542,N_12571);
and U12607 (N_12607,N_12449,N_12597);
xnor U12608 (N_12608,N_12578,N_12445);
nor U12609 (N_12609,N_12570,N_12553);
and U12610 (N_12610,N_12525,N_12595);
or U12611 (N_12611,N_12464,N_12560);
nand U12612 (N_12612,N_12531,N_12503);
and U12613 (N_12613,N_12457,N_12406);
nor U12614 (N_12614,N_12428,N_12567);
nand U12615 (N_12615,N_12545,N_12465);
and U12616 (N_12616,N_12440,N_12476);
xor U12617 (N_12617,N_12437,N_12539);
or U12618 (N_12618,N_12442,N_12549);
nand U12619 (N_12619,N_12450,N_12474);
and U12620 (N_12620,N_12552,N_12482);
or U12621 (N_12621,N_12584,N_12468);
nand U12622 (N_12622,N_12540,N_12462);
xor U12623 (N_12623,N_12455,N_12438);
nand U12624 (N_12624,N_12454,N_12496);
nand U12625 (N_12625,N_12470,N_12458);
xor U12626 (N_12626,N_12575,N_12599);
and U12627 (N_12627,N_12573,N_12556);
nor U12628 (N_12628,N_12590,N_12528);
xor U12629 (N_12629,N_12583,N_12518);
nand U12630 (N_12630,N_12489,N_12490);
or U12631 (N_12631,N_12419,N_12441);
xnor U12632 (N_12632,N_12409,N_12416);
nor U12633 (N_12633,N_12460,N_12484);
or U12634 (N_12634,N_12497,N_12402);
nor U12635 (N_12635,N_12593,N_12405);
and U12636 (N_12636,N_12420,N_12579);
and U12637 (N_12637,N_12511,N_12480);
nor U12638 (N_12638,N_12475,N_12557);
nand U12639 (N_12639,N_12565,N_12461);
and U12640 (N_12640,N_12431,N_12411);
nand U12641 (N_12641,N_12407,N_12400);
nor U12642 (N_12642,N_12519,N_12541);
or U12643 (N_12643,N_12499,N_12537);
and U12644 (N_12644,N_12598,N_12546);
nor U12645 (N_12645,N_12401,N_12478);
nand U12646 (N_12646,N_12543,N_12418);
and U12647 (N_12647,N_12434,N_12424);
or U12648 (N_12648,N_12417,N_12517);
nor U12649 (N_12649,N_12534,N_12566);
nor U12650 (N_12650,N_12422,N_12547);
or U12651 (N_12651,N_12483,N_12562);
nand U12652 (N_12652,N_12436,N_12500);
nor U12653 (N_12653,N_12529,N_12558);
nand U12654 (N_12654,N_12477,N_12555);
xor U12655 (N_12655,N_12524,N_12533);
or U12656 (N_12656,N_12479,N_12423);
and U12657 (N_12657,N_12433,N_12448);
or U12658 (N_12658,N_12574,N_12451);
nand U12659 (N_12659,N_12492,N_12426);
xor U12660 (N_12660,N_12513,N_12530);
nand U12661 (N_12661,N_12444,N_12527);
nand U12662 (N_12662,N_12435,N_12591);
or U12663 (N_12663,N_12410,N_12587);
nand U12664 (N_12664,N_12443,N_12592);
or U12665 (N_12665,N_12413,N_12430);
nand U12666 (N_12666,N_12551,N_12487);
and U12667 (N_12667,N_12576,N_12559);
nand U12668 (N_12668,N_12456,N_12532);
nor U12669 (N_12669,N_12544,N_12427);
and U12670 (N_12670,N_12509,N_12488);
and U12671 (N_12671,N_12596,N_12538);
nor U12672 (N_12672,N_12467,N_12481);
xnor U12673 (N_12673,N_12485,N_12408);
and U12674 (N_12674,N_12498,N_12508);
nand U12675 (N_12675,N_12414,N_12563);
nand U12676 (N_12676,N_12502,N_12569);
nor U12677 (N_12677,N_12432,N_12491);
nor U12678 (N_12678,N_12521,N_12493);
xnor U12679 (N_12679,N_12447,N_12586);
nor U12680 (N_12680,N_12505,N_12495);
and U12681 (N_12681,N_12507,N_12473);
nand U12682 (N_12682,N_12486,N_12421);
or U12683 (N_12683,N_12580,N_12582);
and U12684 (N_12684,N_12535,N_12412);
and U12685 (N_12685,N_12561,N_12548);
xor U12686 (N_12686,N_12504,N_12523);
nor U12687 (N_12687,N_12568,N_12471);
or U12688 (N_12688,N_12510,N_12572);
and U12689 (N_12689,N_12501,N_12459);
nand U12690 (N_12690,N_12564,N_12515);
xor U12691 (N_12691,N_12520,N_12429);
nor U12692 (N_12692,N_12588,N_12577);
nand U12693 (N_12693,N_12516,N_12554);
and U12694 (N_12694,N_12466,N_12512);
xor U12695 (N_12695,N_12589,N_12446);
nand U12696 (N_12696,N_12453,N_12594);
xnor U12697 (N_12697,N_12506,N_12581);
and U12698 (N_12698,N_12452,N_12415);
or U12699 (N_12699,N_12536,N_12463);
nor U12700 (N_12700,N_12575,N_12523);
xor U12701 (N_12701,N_12559,N_12563);
or U12702 (N_12702,N_12411,N_12570);
or U12703 (N_12703,N_12500,N_12458);
or U12704 (N_12704,N_12525,N_12428);
and U12705 (N_12705,N_12592,N_12571);
xnor U12706 (N_12706,N_12576,N_12418);
nand U12707 (N_12707,N_12468,N_12522);
xnor U12708 (N_12708,N_12589,N_12534);
nor U12709 (N_12709,N_12470,N_12444);
nand U12710 (N_12710,N_12542,N_12512);
nor U12711 (N_12711,N_12556,N_12525);
and U12712 (N_12712,N_12419,N_12557);
nand U12713 (N_12713,N_12594,N_12481);
and U12714 (N_12714,N_12492,N_12449);
xor U12715 (N_12715,N_12524,N_12573);
xor U12716 (N_12716,N_12536,N_12531);
nor U12717 (N_12717,N_12452,N_12409);
or U12718 (N_12718,N_12573,N_12551);
xnor U12719 (N_12719,N_12459,N_12452);
or U12720 (N_12720,N_12571,N_12565);
nand U12721 (N_12721,N_12596,N_12485);
and U12722 (N_12722,N_12551,N_12490);
xnor U12723 (N_12723,N_12528,N_12521);
nand U12724 (N_12724,N_12509,N_12570);
nand U12725 (N_12725,N_12460,N_12438);
and U12726 (N_12726,N_12414,N_12495);
xnor U12727 (N_12727,N_12511,N_12459);
nand U12728 (N_12728,N_12486,N_12573);
or U12729 (N_12729,N_12552,N_12574);
nand U12730 (N_12730,N_12555,N_12487);
nand U12731 (N_12731,N_12469,N_12546);
xor U12732 (N_12732,N_12538,N_12477);
xor U12733 (N_12733,N_12578,N_12541);
nor U12734 (N_12734,N_12486,N_12504);
and U12735 (N_12735,N_12559,N_12450);
nor U12736 (N_12736,N_12476,N_12493);
nor U12737 (N_12737,N_12426,N_12480);
nand U12738 (N_12738,N_12404,N_12457);
xnor U12739 (N_12739,N_12506,N_12563);
and U12740 (N_12740,N_12401,N_12530);
or U12741 (N_12741,N_12484,N_12571);
and U12742 (N_12742,N_12470,N_12585);
nor U12743 (N_12743,N_12458,N_12541);
nor U12744 (N_12744,N_12414,N_12465);
and U12745 (N_12745,N_12582,N_12512);
nor U12746 (N_12746,N_12545,N_12564);
xnor U12747 (N_12747,N_12485,N_12528);
and U12748 (N_12748,N_12409,N_12446);
nor U12749 (N_12749,N_12445,N_12455);
nor U12750 (N_12750,N_12520,N_12413);
xor U12751 (N_12751,N_12422,N_12577);
and U12752 (N_12752,N_12481,N_12528);
and U12753 (N_12753,N_12487,N_12581);
xnor U12754 (N_12754,N_12492,N_12584);
nor U12755 (N_12755,N_12565,N_12543);
nand U12756 (N_12756,N_12479,N_12450);
nand U12757 (N_12757,N_12483,N_12574);
and U12758 (N_12758,N_12515,N_12415);
and U12759 (N_12759,N_12519,N_12587);
or U12760 (N_12760,N_12443,N_12571);
nor U12761 (N_12761,N_12533,N_12450);
nor U12762 (N_12762,N_12555,N_12585);
and U12763 (N_12763,N_12484,N_12450);
and U12764 (N_12764,N_12507,N_12407);
xnor U12765 (N_12765,N_12406,N_12456);
xor U12766 (N_12766,N_12552,N_12414);
or U12767 (N_12767,N_12530,N_12501);
and U12768 (N_12768,N_12436,N_12526);
and U12769 (N_12769,N_12437,N_12554);
nand U12770 (N_12770,N_12549,N_12586);
or U12771 (N_12771,N_12585,N_12400);
xnor U12772 (N_12772,N_12520,N_12457);
nand U12773 (N_12773,N_12405,N_12528);
nand U12774 (N_12774,N_12471,N_12545);
or U12775 (N_12775,N_12545,N_12587);
and U12776 (N_12776,N_12534,N_12538);
xor U12777 (N_12777,N_12519,N_12573);
nand U12778 (N_12778,N_12491,N_12589);
nand U12779 (N_12779,N_12443,N_12595);
or U12780 (N_12780,N_12426,N_12589);
nor U12781 (N_12781,N_12505,N_12405);
nor U12782 (N_12782,N_12475,N_12547);
xor U12783 (N_12783,N_12455,N_12415);
nand U12784 (N_12784,N_12509,N_12514);
and U12785 (N_12785,N_12519,N_12513);
nor U12786 (N_12786,N_12432,N_12497);
xor U12787 (N_12787,N_12488,N_12588);
nand U12788 (N_12788,N_12482,N_12547);
or U12789 (N_12789,N_12588,N_12512);
nand U12790 (N_12790,N_12534,N_12593);
or U12791 (N_12791,N_12404,N_12441);
nand U12792 (N_12792,N_12587,N_12472);
xnor U12793 (N_12793,N_12491,N_12553);
nor U12794 (N_12794,N_12490,N_12574);
xnor U12795 (N_12795,N_12443,N_12542);
nand U12796 (N_12796,N_12556,N_12427);
nand U12797 (N_12797,N_12469,N_12402);
or U12798 (N_12798,N_12508,N_12589);
nand U12799 (N_12799,N_12598,N_12457);
nor U12800 (N_12800,N_12797,N_12671);
or U12801 (N_12801,N_12756,N_12728);
or U12802 (N_12802,N_12672,N_12690);
or U12803 (N_12803,N_12784,N_12652);
xnor U12804 (N_12804,N_12712,N_12739);
nor U12805 (N_12805,N_12637,N_12703);
xor U12806 (N_12806,N_12664,N_12693);
xor U12807 (N_12807,N_12679,N_12767);
and U12808 (N_12808,N_12638,N_12613);
nor U12809 (N_12809,N_12749,N_12697);
and U12810 (N_12810,N_12620,N_12622);
and U12811 (N_12811,N_12796,N_12798);
nand U12812 (N_12812,N_12619,N_12650);
nor U12813 (N_12813,N_12724,N_12727);
or U12814 (N_12814,N_12665,N_12774);
nor U12815 (N_12815,N_12631,N_12759);
or U12816 (N_12816,N_12709,N_12778);
or U12817 (N_12817,N_12736,N_12621);
nor U12818 (N_12818,N_12625,N_12741);
xor U12819 (N_12819,N_12773,N_12655);
and U12820 (N_12820,N_12639,N_12794);
and U12821 (N_12821,N_12681,N_12731);
nand U12822 (N_12822,N_12707,N_12722);
nor U12823 (N_12823,N_12701,N_12632);
or U12824 (N_12824,N_12602,N_12691);
nand U12825 (N_12825,N_12624,N_12603);
nand U12826 (N_12826,N_12667,N_12725);
xor U12827 (N_12827,N_12623,N_12721);
or U12828 (N_12828,N_12716,N_12641);
nor U12829 (N_12829,N_12744,N_12666);
or U12830 (N_12830,N_12788,N_12777);
or U12831 (N_12831,N_12713,N_12730);
nor U12832 (N_12832,N_12685,N_12766);
xnor U12833 (N_12833,N_12752,N_12740);
or U12834 (N_12834,N_12670,N_12699);
xor U12835 (N_12835,N_12644,N_12710);
nand U12836 (N_12836,N_12769,N_12763);
nand U12837 (N_12837,N_12694,N_12618);
nand U12838 (N_12838,N_12706,N_12792);
and U12839 (N_12839,N_12682,N_12735);
and U12840 (N_12840,N_12771,N_12649);
xor U12841 (N_12841,N_12745,N_12686);
xor U12842 (N_12842,N_12711,N_12714);
nor U12843 (N_12843,N_12733,N_12635);
and U12844 (N_12844,N_12680,N_12669);
xor U12845 (N_12845,N_12646,N_12791);
nor U12846 (N_12846,N_12726,N_12761);
nand U12847 (N_12847,N_12729,N_12606);
nor U12848 (N_12848,N_12781,N_12643);
nand U12849 (N_12849,N_12692,N_12628);
or U12850 (N_12850,N_12734,N_12787);
xor U12851 (N_12851,N_12698,N_12687);
nor U12852 (N_12852,N_12660,N_12684);
nand U12853 (N_12853,N_12786,N_12668);
or U12854 (N_12854,N_12732,N_12799);
nand U12855 (N_12855,N_12717,N_12695);
nor U12856 (N_12856,N_12674,N_12783);
nand U12857 (N_12857,N_12755,N_12765);
and U12858 (N_12858,N_12762,N_12617);
and U12859 (N_12859,N_12636,N_12757);
or U12860 (N_12860,N_12675,N_12758);
nor U12861 (N_12861,N_12612,N_12723);
or U12862 (N_12862,N_12683,N_12779);
nor U12863 (N_12863,N_12688,N_12656);
xor U12864 (N_12864,N_12626,N_12746);
or U12865 (N_12865,N_12600,N_12751);
nand U12866 (N_12866,N_12604,N_12795);
and U12867 (N_12867,N_12648,N_12676);
and U12868 (N_12868,N_12614,N_12719);
xor U12869 (N_12869,N_12673,N_12768);
nand U12870 (N_12870,N_12651,N_12702);
and U12871 (N_12871,N_12760,N_12677);
or U12872 (N_12872,N_12708,N_12607);
nand U12873 (N_12873,N_12782,N_12640);
or U12874 (N_12874,N_12654,N_12659);
nand U12875 (N_12875,N_12663,N_12657);
and U12876 (N_12876,N_12775,N_12601);
or U12877 (N_12877,N_12634,N_12610);
nor U12878 (N_12878,N_12718,N_12700);
xor U12879 (N_12879,N_12658,N_12653);
nor U12880 (N_12880,N_12790,N_12645);
nor U12881 (N_12881,N_12630,N_12753);
nor U12882 (N_12882,N_12793,N_12780);
and U12883 (N_12883,N_12704,N_12747);
nor U12884 (N_12884,N_12720,N_12705);
nand U12885 (N_12885,N_12642,N_12789);
or U12886 (N_12886,N_12785,N_12748);
or U12887 (N_12887,N_12715,N_12609);
and U12888 (N_12888,N_12678,N_12743);
nand U12889 (N_12889,N_12661,N_12611);
nand U12890 (N_12890,N_12764,N_12750);
and U12891 (N_12891,N_12633,N_12742);
xnor U12892 (N_12892,N_12615,N_12737);
and U12893 (N_12893,N_12605,N_12696);
and U12894 (N_12894,N_12689,N_12770);
nor U12895 (N_12895,N_12662,N_12738);
xor U12896 (N_12896,N_12616,N_12627);
and U12897 (N_12897,N_12647,N_12776);
or U12898 (N_12898,N_12754,N_12629);
nand U12899 (N_12899,N_12608,N_12772);
xnor U12900 (N_12900,N_12738,N_12614);
nand U12901 (N_12901,N_12739,N_12765);
or U12902 (N_12902,N_12672,N_12657);
nor U12903 (N_12903,N_12700,N_12644);
and U12904 (N_12904,N_12672,N_12742);
or U12905 (N_12905,N_12772,N_12763);
nand U12906 (N_12906,N_12734,N_12728);
xor U12907 (N_12907,N_12725,N_12646);
nor U12908 (N_12908,N_12754,N_12672);
and U12909 (N_12909,N_12761,N_12791);
nor U12910 (N_12910,N_12697,N_12747);
nand U12911 (N_12911,N_12724,N_12609);
xnor U12912 (N_12912,N_12729,N_12620);
nand U12913 (N_12913,N_12779,N_12687);
or U12914 (N_12914,N_12622,N_12778);
or U12915 (N_12915,N_12650,N_12610);
xnor U12916 (N_12916,N_12667,N_12705);
and U12917 (N_12917,N_12769,N_12768);
nor U12918 (N_12918,N_12797,N_12647);
nand U12919 (N_12919,N_12675,N_12729);
and U12920 (N_12920,N_12693,N_12685);
nor U12921 (N_12921,N_12607,N_12694);
nand U12922 (N_12922,N_12707,N_12692);
xnor U12923 (N_12923,N_12624,N_12711);
or U12924 (N_12924,N_12797,N_12684);
or U12925 (N_12925,N_12718,N_12706);
nand U12926 (N_12926,N_12645,N_12757);
or U12927 (N_12927,N_12688,N_12785);
or U12928 (N_12928,N_12625,N_12798);
and U12929 (N_12929,N_12727,N_12636);
nand U12930 (N_12930,N_12776,N_12764);
nand U12931 (N_12931,N_12669,N_12652);
nor U12932 (N_12932,N_12678,N_12717);
nor U12933 (N_12933,N_12687,N_12669);
nand U12934 (N_12934,N_12665,N_12734);
xnor U12935 (N_12935,N_12665,N_12775);
nor U12936 (N_12936,N_12761,N_12723);
and U12937 (N_12937,N_12644,N_12656);
nor U12938 (N_12938,N_12742,N_12756);
and U12939 (N_12939,N_12676,N_12634);
or U12940 (N_12940,N_12719,N_12788);
xor U12941 (N_12941,N_12616,N_12746);
xnor U12942 (N_12942,N_12668,N_12694);
or U12943 (N_12943,N_12690,N_12630);
nand U12944 (N_12944,N_12703,N_12636);
nor U12945 (N_12945,N_12780,N_12763);
and U12946 (N_12946,N_12600,N_12755);
nor U12947 (N_12947,N_12657,N_12762);
nor U12948 (N_12948,N_12604,N_12620);
nor U12949 (N_12949,N_12715,N_12686);
xnor U12950 (N_12950,N_12706,N_12677);
and U12951 (N_12951,N_12604,N_12713);
nand U12952 (N_12952,N_12636,N_12685);
xnor U12953 (N_12953,N_12789,N_12634);
nand U12954 (N_12954,N_12771,N_12691);
and U12955 (N_12955,N_12704,N_12678);
nor U12956 (N_12956,N_12638,N_12696);
nand U12957 (N_12957,N_12728,N_12656);
nor U12958 (N_12958,N_12783,N_12612);
or U12959 (N_12959,N_12783,N_12620);
and U12960 (N_12960,N_12634,N_12667);
nand U12961 (N_12961,N_12770,N_12668);
xor U12962 (N_12962,N_12726,N_12719);
or U12963 (N_12963,N_12683,N_12634);
or U12964 (N_12964,N_12638,N_12792);
or U12965 (N_12965,N_12694,N_12772);
nor U12966 (N_12966,N_12605,N_12660);
nor U12967 (N_12967,N_12709,N_12686);
and U12968 (N_12968,N_12757,N_12763);
nor U12969 (N_12969,N_12667,N_12716);
xor U12970 (N_12970,N_12683,N_12717);
and U12971 (N_12971,N_12605,N_12724);
xnor U12972 (N_12972,N_12787,N_12621);
nor U12973 (N_12973,N_12673,N_12778);
nor U12974 (N_12974,N_12747,N_12723);
nor U12975 (N_12975,N_12762,N_12636);
or U12976 (N_12976,N_12666,N_12794);
xnor U12977 (N_12977,N_12646,N_12733);
or U12978 (N_12978,N_12643,N_12655);
or U12979 (N_12979,N_12687,N_12694);
and U12980 (N_12980,N_12675,N_12639);
xnor U12981 (N_12981,N_12614,N_12720);
or U12982 (N_12982,N_12635,N_12729);
nor U12983 (N_12983,N_12637,N_12611);
xnor U12984 (N_12984,N_12703,N_12640);
nor U12985 (N_12985,N_12657,N_12765);
nand U12986 (N_12986,N_12672,N_12628);
xor U12987 (N_12987,N_12633,N_12786);
xnor U12988 (N_12988,N_12689,N_12752);
nor U12989 (N_12989,N_12794,N_12768);
and U12990 (N_12990,N_12672,N_12769);
nor U12991 (N_12991,N_12693,N_12765);
nor U12992 (N_12992,N_12678,N_12752);
nor U12993 (N_12993,N_12730,N_12779);
or U12994 (N_12994,N_12768,N_12647);
or U12995 (N_12995,N_12730,N_12665);
nand U12996 (N_12996,N_12639,N_12765);
nor U12997 (N_12997,N_12638,N_12733);
or U12998 (N_12998,N_12662,N_12718);
and U12999 (N_12999,N_12687,N_12630);
or U13000 (N_13000,N_12894,N_12982);
xnor U13001 (N_13001,N_12803,N_12801);
xnor U13002 (N_13002,N_12822,N_12950);
nor U13003 (N_13003,N_12948,N_12964);
nor U13004 (N_13004,N_12813,N_12910);
and U13005 (N_13005,N_12892,N_12960);
or U13006 (N_13006,N_12904,N_12805);
and U13007 (N_13007,N_12937,N_12821);
nor U13008 (N_13008,N_12958,N_12853);
or U13009 (N_13009,N_12846,N_12997);
or U13010 (N_13010,N_12935,N_12852);
xor U13011 (N_13011,N_12945,N_12902);
and U13012 (N_13012,N_12978,N_12876);
nor U13013 (N_13013,N_12838,N_12856);
nand U13014 (N_13014,N_12925,N_12919);
and U13015 (N_13015,N_12927,N_12848);
nor U13016 (N_13016,N_12827,N_12824);
and U13017 (N_13017,N_12946,N_12979);
and U13018 (N_13018,N_12977,N_12845);
and U13019 (N_13019,N_12847,N_12855);
or U13020 (N_13020,N_12888,N_12939);
nor U13021 (N_13021,N_12943,N_12980);
nand U13022 (N_13022,N_12859,N_12951);
or U13023 (N_13023,N_12870,N_12899);
and U13024 (N_13024,N_12913,N_12895);
nor U13025 (N_13025,N_12998,N_12915);
nor U13026 (N_13026,N_12933,N_12885);
or U13027 (N_13027,N_12952,N_12893);
or U13028 (N_13028,N_12889,N_12802);
nand U13029 (N_13029,N_12944,N_12834);
or U13030 (N_13030,N_12861,N_12879);
nand U13031 (N_13031,N_12955,N_12994);
nand U13032 (N_13032,N_12832,N_12934);
xor U13033 (N_13033,N_12873,N_12975);
and U13034 (N_13034,N_12909,N_12971);
nor U13035 (N_13035,N_12901,N_12996);
xnor U13036 (N_13036,N_12966,N_12981);
nor U13037 (N_13037,N_12911,N_12804);
nor U13038 (N_13038,N_12867,N_12860);
nor U13039 (N_13039,N_12941,N_12961);
and U13040 (N_13040,N_12983,N_12825);
xor U13041 (N_13041,N_12840,N_12988);
nand U13042 (N_13042,N_12865,N_12884);
xor U13043 (N_13043,N_12849,N_12854);
nand U13044 (N_13044,N_12828,N_12863);
or U13045 (N_13045,N_12842,N_12914);
xor U13046 (N_13046,N_12918,N_12932);
xnor U13047 (N_13047,N_12800,N_12875);
xor U13048 (N_13048,N_12999,N_12831);
nor U13049 (N_13049,N_12833,N_12886);
or U13050 (N_13050,N_12819,N_12923);
or U13051 (N_13051,N_12816,N_12940);
or U13052 (N_13052,N_12986,N_12924);
and U13053 (N_13053,N_12807,N_12829);
xnor U13054 (N_13054,N_12817,N_12968);
nor U13055 (N_13055,N_12903,N_12905);
nand U13056 (N_13056,N_12898,N_12992);
xor U13057 (N_13057,N_12844,N_12922);
or U13058 (N_13058,N_12841,N_12972);
xor U13059 (N_13059,N_12928,N_12862);
nand U13060 (N_13060,N_12814,N_12976);
nand U13061 (N_13061,N_12957,N_12987);
and U13062 (N_13062,N_12880,N_12823);
xor U13063 (N_13063,N_12811,N_12947);
and U13064 (N_13064,N_12920,N_12912);
or U13065 (N_13065,N_12869,N_12967);
nand U13066 (N_13066,N_12820,N_12916);
and U13067 (N_13067,N_12985,N_12890);
xnor U13068 (N_13068,N_12974,N_12926);
nor U13069 (N_13069,N_12929,N_12871);
or U13070 (N_13070,N_12942,N_12995);
xnor U13071 (N_13071,N_12868,N_12872);
and U13072 (N_13072,N_12962,N_12897);
nor U13073 (N_13073,N_12857,N_12883);
nor U13074 (N_13074,N_12993,N_12949);
or U13075 (N_13075,N_12837,N_12954);
nor U13076 (N_13076,N_12850,N_12806);
xnor U13077 (N_13077,N_12815,N_12808);
nand U13078 (N_13078,N_12956,N_12931);
or U13079 (N_13079,N_12917,N_12830);
nor U13080 (N_13080,N_12836,N_12930);
nor U13081 (N_13081,N_12877,N_12858);
xnor U13082 (N_13082,N_12906,N_12843);
or U13083 (N_13083,N_12908,N_12864);
or U13084 (N_13084,N_12810,N_12826);
nor U13085 (N_13085,N_12907,N_12835);
xor U13086 (N_13086,N_12990,N_12984);
xor U13087 (N_13087,N_12812,N_12851);
or U13088 (N_13088,N_12882,N_12809);
and U13089 (N_13089,N_12839,N_12973);
xnor U13090 (N_13090,N_12938,N_12921);
nor U13091 (N_13091,N_12959,N_12953);
nand U13092 (N_13092,N_12818,N_12896);
nor U13093 (N_13093,N_12989,N_12881);
nor U13094 (N_13094,N_12936,N_12887);
nand U13095 (N_13095,N_12965,N_12878);
xnor U13096 (N_13096,N_12991,N_12969);
xor U13097 (N_13097,N_12866,N_12970);
nand U13098 (N_13098,N_12900,N_12963);
xnor U13099 (N_13099,N_12874,N_12891);
nand U13100 (N_13100,N_12960,N_12831);
or U13101 (N_13101,N_12929,N_12811);
or U13102 (N_13102,N_12996,N_12983);
and U13103 (N_13103,N_12839,N_12937);
and U13104 (N_13104,N_12891,N_12855);
nor U13105 (N_13105,N_12952,N_12845);
nor U13106 (N_13106,N_12893,N_12823);
or U13107 (N_13107,N_12931,N_12964);
and U13108 (N_13108,N_12916,N_12804);
nor U13109 (N_13109,N_12883,N_12833);
nand U13110 (N_13110,N_12949,N_12810);
or U13111 (N_13111,N_12876,N_12861);
xor U13112 (N_13112,N_12820,N_12910);
or U13113 (N_13113,N_12832,N_12940);
nand U13114 (N_13114,N_12899,N_12847);
or U13115 (N_13115,N_12929,N_12907);
nor U13116 (N_13116,N_12888,N_12933);
nor U13117 (N_13117,N_12973,N_12900);
xor U13118 (N_13118,N_12909,N_12880);
nor U13119 (N_13119,N_12908,N_12800);
nor U13120 (N_13120,N_12950,N_12995);
xnor U13121 (N_13121,N_12950,N_12845);
or U13122 (N_13122,N_12928,N_12904);
or U13123 (N_13123,N_12834,N_12919);
nor U13124 (N_13124,N_12930,N_12858);
nor U13125 (N_13125,N_12969,N_12934);
xnor U13126 (N_13126,N_12912,N_12950);
and U13127 (N_13127,N_12942,N_12867);
nand U13128 (N_13128,N_12872,N_12810);
nor U13129 (N_13129,N_12903,N_12938);
nand U13130 (N_13130,N_12982,N_12979);
nor U13131 (N_13131,N_12966,N_12931);
or U13132 (N_13132,N_12919,N_12886);
nand U13133 (N_13133,N_12831,N_12990);
and U13134 (N_13134,N_12862,N_12955);
nor U13135 (N_13135,N_12992,N_12956);
xor U13136 (N_13136,N_12973,N_12895);
or U13137 (N_13137,N_12964,N_12803);
or U13138 (N_13138,N_12801,N_12965);
and U13139 (N_13139,N_12872,N_12916);
xnor U13140 (N_13140,N_12940,N_12977);
nor U13141 (N_13141,N_12977,N_12922);
nand U13142 (N_13142,N_12923,N_12825);
and U13143 (N_13143,N_12953,N_12966);
nand U13144 (N_13144,N_12911,N_12809);
xnor U13145 (N_13145,N_12878,N_12827);
and U13146 (N_13146,N_12855,N_12811);
and U13147 (N_13147,N_12865,N_12943);
nor U13148 (N_13148,N_12938,N_12927);
and U13149 (N_13149,N_12839,N_12929);
nor U13150 (N_13150,N_12982,N_12876);
nor U13151 (N_13151,N_12832,N_12978);
nand U13152 (N_13152,N_12871,N_12890);
nand U13153 (N_13153,N_12860,N_12829);
xor U13154 (N_13154,N_12855,N_12974);
or U13155 (N_13155,N_12822,N_12807);
or U13156 (N_13156,N_12888,N_12928);
or U13157 (N_13157,N_12853,N_12823);
and U13158 (N_13158,N_12918,N_12850);
nand U13159 (N_13159,N_12880,N_12920);
xnor U13160 (N_13160,N_12878,N_12818);
and U13161 (N_13161,N_12917,N_12969);
or U13162 (N_13162,N_12998,N_12913);
nand U13163 (N_13163,N_12842,N_12926);
nor U13164 (N_13164,N_12972,N_12838);
nand U13165 (N_13165,N_12899,N_12868);
nand U13166 (N_13166,N_12818,N_12938);
or U13167 (N_13167,N_12801,N_12852);
or U13168 (N_13168,N_12966,N_12821);
and U13169 (N_13169,N_12953,N_12981);
and U13170 (N_13170,N_12972,N_12960);
nor U13171 (N_13171,N_12998,N_12941);
nand U13172 (N_13172,N_12924,N_12851);
nor U13173 (N_13173,N_12862,N_12847);
or U13174 (N_13174,N_12980,N_12834);
or U13175 (N_13175,N_12932,N_12887);
nor U13176 (N_13176,N_12964,N_12801);
or U13177 (N_13177,N_12936,N_12822);
nor U13178 (N_13178,N_12939,N_12897);
nand U13179 (N_13179,N_12962,N_12917);
nor U13180 (N_13180,N_12924,N_12869);
xnor U13181 (N_13181,N_12930,N_12886);
nand U13182 (N_13182,N_12816,N_12815);
and U13183 (N_13183,N_12918,N_12921);
nand U13184 (N_13184,N_12928,N_12909);
xor U13185 (N_13185,N_12909,N_12913);
nor U13186 (N_13186,N_12856,N_12809);
nor U13187 (N_13187,N_12877,N_12801);
nand U13188 (N_13188,N_12908,N_12977);
nor U13189 (N_13189,N_12861,N_12830);
or U13190 (N_13190,N_12822,N_12946);
and U13191 (N_13191,N_12811,N_12943);
xor U13192 (N_13192,N_12973,N_12981);
nand U13193 (N_13193,N_12905,N_12811);
nor U13194 (N_13194,N_12927,N_12954);
nor U13195 (N_13195,N_12989,N_12944);
nand U13196 (N_13196,N_12848,N_12804);
and U13197 (N_13197,N_12868,N_12871);
and U13198 (N_13198,N_12933,N_12956);
and U13199 (N_13199,N_12940,N_12903);
or U13200 (N_13200,N_13091,N_13186);
nand U13201 (N_13201,N_13157,N_13095);
nand U13202 (N_13202,N_13083,N_13183);
nand U13203 (N_13203,N_13193,N_13060);
nor U13204 (N_13204,N_13122,N_13144);
nor U13205 (N_13205,N_13132,N_13125);
nor U13206 (N_13206,N_13079,N_13156);
xnor U13207 (N_13207,N_13053,N_13021);
or U13208 (N_13208,N_13191,N_13048);
xor U13209 (N_13209,N_13008,N_13100);
xnor U13210 (N_13210,N_13196,N_13116);
and U13211 (N_13211,N_13107,N_13113);
and U13212 (N_13212,N_13050,N_13019);
nor U13213 (N_13213,N_13141,N_13198);
nor U13214 (N_13214,N_13173,N_13080);
nand U13215 (N_13215,N_13180,N_13064);
or U13216 (N_13216,N_13162,N_13020);
and U13217 (N_13217,N_13015,N_13031);
or U13218 (N_13218,N_13160,N_13046);
and U13219 (N_13219,N_13087,N_13004);
or U13220 (N_13220,N_13149,N_13138);
xnor U13221 (N_13221,N_13176,N_13197);
nor U13222 (N_13222,N_13104,N_13045);
and U13223 (N_13223,N_13047,N_13136);
and U13224 (N_13224,N_13121,N_13185);
nor U13225 (N_13225,N_13102,N_13188);
and U13226 (N_13226,N_13145,N_13076);
xor U13227 (N_13227,N_13163,N_13052);
xnor U13228 (N_13228,N_13135,N_13119);
and U13229 (N_13229,N_13118,N_13130);
and U13230 (N_13230,N_13093,N_13187);
and U13231 (N_13231,N_13195,N_13101);
and U13232 (N_13232,N_13131,N_13098);
and U13233 (N_13233,N_13063,N_13075);
or U13234 (N_13234,N_13124,N_13061);
or U13235 (N_13235,N_13159,N_13105);
nor U13236 (N_13236,N_13000,N_13133);
nor U13237 (N_13237,N_13024,N_13073);
nor U13238 (N_13238,N_13151,N_13117);
and U13239 (N_13239,N_13114,N_13088);
xnor U13240 (N_13240,N_13171,N_13011);
or U13241 (N_13241,N_13152,N_13090);
nor U13242 (N_13242,N_13174,N_13178);
or U13243 (N_13243,N_13194,N_13085);
xnor U13244 (N_13244,N_13054,N_13150);
nor U13245 (N_13245,N_13097,N_13143);
and U13246 (N_13246,N_13014,N_13140);
or U13247 (N_13247,N_13057,N_13018);
xnor U13248 (N_13248,N_13148,N_13153);
nor U13249 (N_13249,N_13072,N_13103);
nor U13250 (N_13250,N_13169,N_13016);
and U13251 (N_13251,N_13033,N_13165);
nand U13252 (N_13252,N_13170,N_13168);
or U13253 (N_13253,N_13042,N_13077);
nor U13254 (N_13254,N_13071,N_13161);
or U13255 (N_13255,N_13115,N_13081);
xnor U13256 (N_13256,N_13084,N_13059);
xnor U13257 (N_13257,N_13025,N_13036);
nand U13258 (N_13258,N_13089,N_13123);
nor U13259 (N_13259,N_13109,N_13041);
xor U13260 (N_13260,N_13039,N_13037);
and U13261 (N_13261,N_13128,N_13012);
or U13262 (N_13262,N_13044,N_13108);
or U13263 (N_13263,N_13074,N_13003);
and U13264 (N_13264,N_13070,N_13184);
or U13265 (N_13265,N_13001,N_13129);
or U13266 (N_13266,N_13106,N_13055);
nor U13267 (N_13267,N_13086,N_13142);
or U13268 (N_13268,N_13049,N_13032);
nand U13269 (N_13269,N_13043,N_13137);
and U13270 (N_13270,N_13026,N_13094);
or U13271 (N_13271,N_13154,N_13111);
nand U13272 (N_13272,N_13038,N_13002);
nand U13273 (N_13273,N_13164,N_13120);
xor U13274 (N_13274,N_13190,N_13167);
xor U13275 (N_13275,N_13181,N_13127);
or U13276 (N_13276,N_13022,N_13189);
and U13277 (N_13277,N_13166,N_13030);
or U13278 (N_13278,N_13062,N_13010);
or U13279 (N_13279,N_13027,N_13110);
xor U13280 (N_13280,N_13177,N_13067);
nand U13281 (N_13281,N_13017,N_13023);
xnor U13282 (N_13282,N_13139,N_13146);
nor U13283 (N_13283,N_13013,N_13028);
xor U13284 (N_13284,N_13034,N_13179);
nand U13285 (N_13285,N_13112,N_13182);
nor U13286 (N_13286,N_13192,N_13006);
or U13287 (N_13287,N_13155,N_13126);
or U13288 (N_13288,N_13051,N_13040);
and U13289 (N_13289,N_13099,N_13029);
nand U13290 (N_13290,N_13058,N_13158);
nand U13291 (N_13291,N_13092,N_13007);
and U13292 (N_13292,N_13172,N_13147);
nor U13293 (N_13293,N_13096,N_13078);
nand U13294 (N_13294,N_13069,N_13056);
xnor U13295 (N_13295,N_13068,N_13035);
or U13296 (N_13296,N_13082,N_13066);
or U13297 (N_13297,N_13005,N_13009);
and U13298 (N_13298,N_13065,N_13175);
nor U13299 (N_13299,N_13199,N_13134);
nand U13300 (N_13300,N_13160,N_13117);
nand U13301 (N_13301,N_13071,N_13119);
nand U13302 (N_13302,N_13148,N_13055);
nor U13303 (N_13303,N_13012,N_13162);
or U13304 (N_13304,N_13070,N_13134);
nand U13305 (N_13305,N_13196,N_13041);
or U13306 (N_13306,N_13045,N_13082);
xnor U13307 (N_13307,N_13096,N_13066);
nand U13308 (N_13308,N_13080,N_13112);
nor U13309 (N_13309,N_13095,N_13050);
xnor U13310 (N_13310,N_13107,N_13196);
and U13311 (N_13311,N_13076,N_13058);
xnor U13312 (N_13312,N_13029,N_13149);
nand U13313 (N_13313,N_13144,N_13012);
nand U13314 (N_13314,N_13026,N_13057);
or U13315 (N_13315,N_13083,N_13191);
nand U13316 (N_13316,N_13162,N_13079);
xor U13317 (N_13317,N_13191,N_13168);
xor U13318 (N_13318,N_13055,N_13145);
or U13319 (N_13319,N_13188,N_13066);
nand U13320 (N_13320,N_13158,N_13149);
or U13321 (N_13321,N_13125,N_13011);
nor U13322 (N_13322,N_13057,N_13150);
nand U13323 (N_13323,N_13071,N_13015);
and U13324 (N_13324,N_13008,N_13021);
xor U13325 (N_13325,N_13123,N_13137);
nor U13326 (N_13326,N_13196,N_13018);
nand U13327 (N_13327,N_13152,N_13059);
or U13328 (N_13328,N_13114,N_13106);
and U13329 (N_13329,N_13191,N_13108);
or U13330 (N_13330,N_13031,N_13052);
nor U13331 (N_13331,N_13022,N_13169);
or U13332 (N_13332,N_13081,N_13107);
and U13333 (N_13333,N_13127,N_13014);
or U13334 (N_13334,N_13164,N_13076);
or U13335 (N_13335,N_13091,N_13057);
nand U13336 (N_13336,N_13054,N_13124);
nor U13337 (N_13337,N_13031,N_13077);
or U13338 (N_13338,N_13114,N_13115);
or U13339 (N_13339,N_13130,N_13160);
and U13340 (N_13340,N_13043,N_13172);
xor U13341 (N_13341,N_13066,N_13123);
xor U13342 (N_13342,N_13022,N_13094);
and U13343 (N_13343,N_13157,N_13108);
and U13344 (N_13344,N_13070,N_13162);
nor U13345 (N_13345,N_13050,N_13014);
nor U13346 (N_13346,N_13012,N_13014);
xor U13347 (N_13347,N_13068,N_13180);
xor U13348 (N_13348,N_13117,N_13125);
nand U13349 (N_13349,N_13008,N_13048);
nor U13350 (N_13350,N_13192,N_13187);
xor U13351 (N_13351,N_13128,N_13076);
or U13352 (N_13352,N_13154,N_13007);
nand U13353 (N_13353,N_13112,N_13097);
xnor U13354 (N_13354,N_13159,N_13187);
and U13355 (N_13355,N_13145,N_13141);
xor U13356 (N_13356,N_13084,N_13191);
xnor U13357 (N_13357,N_13118,N_13147);
or U13358 (N_13358,N_13190,N_13112);
and U13359 (N_13359,N_13151,N_13108);
and U13360 (N_13360,N_13168,N_13043);
nor U13361 (N_13361,N_13005,N_13169);
xor U13362 (N_13362,N_13043,N_13045);
nor U13363 (N_13363,N_13119,N_13022);
xnor U13364 (N_13364,N_13114,N_13016);
xnor U13365 (N_13365,N_13018,N_13002);
nand U13366 (N_13366,N_13050,N_13098);
xnor U13367 (N_13367,N_13143,N_13137);
or U13368 (N_13368,N_13141,N_13082);
and U13369 (N_13369,N_13070,N_13119);
or U13370 (N_13370,N_13151,N_13165);
nand U13371 (N_13371,N_13182,N_13088);
or U13372 (N_13372,N_13046,N_13087);
and U13373 (N_13373,N_13154,N_13023);
nand U13374 (N_13374,N_13184,N_13198);
nor U13375 (N_13375,N_13183,N_13196);
nor U13376 (N_13376,N_13028,N_13139);
and U13377 (N_13377,N_13178,N_13055);
or U13378 (N_13378,N_13092,N_13090);
nand U13379 (N_13379,N_13048,N_13095);
xnor U13380 (N_13380,N_13039,N_13129);
or U13381 (N_13381,N_13186,N_13039);
xor U13382 (N_13382,N_13041,N_13038);
nand U13383 (N_13383,N_13178,N_13188);
or U13384 (N_13384,N_13080,N_13036);
xnor U13385 (N_13385,N_13001,N_13006);
nor U13386 (N_13386,N_13027,N_13130);
and U13387 (N_13387,N_13154,N_13161);
nand U13388 (N_13388,N_13175,N_13114);
and U13389 (N_13389,N_13163,N_13150);
or U13390 (N_13390,N_13021,N_13182);
or U13391 (N_13391,N_13125,N_13097);
or U13392 (N_13392,N_13066,N_13049);
nor U13393 (N_13393,N_13184,N_13024);
xor U13394 (N_13394,N_13156,N_13078);
and U13395 (N_13395,N_13075,N_13181);
nand U13396 (N_13396,N_13080,N_13073);
xor U13397 (N_13397,N_13059,N_13090);
and U13398 (N_13398,N_13146,N_13182);
and U13399 (N_13399,N_13072,N_13198);
nor U13400 (N_13400,N_13252,N_13271);
nand U13401 (N_13401,N_13264,N_13256);
nand U13402 (N_13402,N_13398,N_13274);
and U13403 (N_13403,N_13288,N_13211);
and U13404 (N_13404,N_13204,N_13386);
nand U13405 (N_13405,N_13214,N_13320);
or U13406 (N_13406,N_13323,N_13381);
nand U13407 (N_13407,N_13321,N_13331);
nor U13408 (N_13408,N_13282,N_13290);
nand U13409 (N_13409,N_13266,N_13203);
xor U13410 (N_13410,N_13350,N_13361);
or U13411 (N_13411,N_13393,N_13324);
nand U13412 (N_13412,N_13226,N_13305);
and U13413 (N_13413,N_13212,N_13333);
or U13414 (N_13414,N_13246,N_13276);
xnor U13415 (N_13415,N_13216,N_13249);
xnor U13416 (N_13416,N_13313,N_13255);
or U13417 (N_13417,N_13294,N_13311);
xor U13418 (N_13418,N_13353,N_13210);
nor U13419 (N_13419,N_13248,N_13316);
and U13420 (N_13420,N_13222,N_13259);
or U13421 (N_13421,N_13209,N_13231);
or U13422 (N_13422,N_13382,N_13301);
or U13423 (N_13423,N_13205,N_13357);
or U13424 (N_13424,N_13317,N_13201);
xor U13425 (N_13425,N_13367,N_13227);
nor U13426 (N_13426,N_13267,N_13335);
xnor U13427 (N_13427,N_13303,N_13218);
nor U13428 (N_13428,N_13258,N_13396);
or U13429 (N_13429,N_13340,N_13334);
nor U13430 (N_13430,N_13383,N_13235);
nor U13431 (N_13431,N_13338,N_13379);
and U13432 (N_13432,N_13354,N_13336);
nand U13433 (N_13433,N_13215,N_13344);
or U13434 (N_13434,N_13360,N_13224);
xnor U13435 (N_13435,N_13208,N_13318);
or U13436 (N_13436,N_13332,N_13314);
or U13437 (N_13437,N_13388,N_13343);
or U13438 (N_13438,N_13241,N_13238);
xor U13439 (N_13439,N_13217,N_13346);
nand U13440 (N_13440,N_13319,N_13348);
nor U13441 (N_13441,N_13355,N_13300);
or U13442 (N_13442,N_13397,N_13244);
nor U13443 (N_13443,N_13251,N_13395);
or U13444 (N_13444,N_13368,N_13376);
nor U13445 (N_13445,N_13234,N_13351);
xor U13446 (N_13446,N_13265,N_13296);
nand U13447 (N_13447,N_13391,N_13375);
or U13448 (N_13448,N_13371,N_13229);
xor U13449 (N_13449,N_13247,N_13253);
or U13450 (N_13450,N_13387,N_13281);
nand U13451 (N_13451,N_13330,N_13306);
or U13452 (N_13452,N_13292,N_13365);
nand U13453 (N_13453,N_13279,N_13399);
or U13454 (N_13454,N_13342,N_13349);
xor U13455 (N_13455,N_13322,N_13219);
nor U13456 (N_13456,N_13325,N_13299);
and U13457 (N_13457,N_13202,N_13270);
nand U13458 (N_13458,N_13287,N_13254);
nor U13459 (N_13459,N_13372,N_13260);
xnor U13460 (N_13460,N_13286,N_13230);
nand U13461 (N_13461,N_13232,N_13263);
nand U13462 (N_13462,N_13378,N_13328);
nor U13463 (N_13463,N_13312,N_13297);
nor U13464 (N_13464,N_13239,N_13278);
xor U13465 (N_13465,N_13285,N_13289);
nor U13466 (N_13466,N_13250,N_13302);
nand U13467 (N_13467,N_13374,N_13394);
and U13468 (N_13468,N_13240,N_13310);
nand U13469 (N_13469,N_13277,N_13373);
nor U13470 (N_13470,N_13339,N_13315);
nor U13471 (N_13471,N_13298,N_13200);
and U13472 (N_13472,N_13280,N_13384);
nor U13473 (N_13473,N_13326,N_13304);
nor U13474 (N_13474,N_13207,N_13206);
nor U13475 (N_13475,N_13236,N_13257);
and U13476 (N_13476,N_13284,N_13362);
nand U13477 (N_13477,N_13295,N_13228);
nor U13478 (N_13478,N_13269,N_13345);
nand U13479 (N_13479,N_13329,N_13363);
nand U13480 (N_13480,N_13262,N_13242);
nand U13481 (N_13481,N_13392,N_13307);
or U13482 (N_13482,N_13272,N_13341);
xor U13483 (N_13483,N_13309,N_13275);
nor U13484 (N_13484,N_13389,N_13245);
and U13485 (N_13485,N_13233,N_13359);
nand U13486 (N_13486,N_13370,N_13327);
xnor U13487 (N_13487,N_13213,N_13366);
or U13488 (N_13488,N_13283,N_13377);
nand U13489 (N_13489,N_13358,N_13237);
nor U13490 (N_13490,N_13390,N_13347);
nand U13491 (N_13491,N_13308,N_13221);
xnor U13492 (N_13492,N_13364,N_13293);
or U13493 (N_13493,N_13337,N_13356);
nand U13494 (N_13494,N_13380,N_13220);
nor U13495 (N_13495,N_13268,N_13369);
or U13496 (N_13496,N_13273,N_13291);
and U13497 (N_13497,N_13352,N_13261);
nand U13498 (N_13498,N_13385,N_13223);
nand U13499 (N_13499,N_13225,N_13243);
or U13500 (N_13500,N_13324,N_13287);
nand U13501 (N_13501,N_13251,N_13220);
and U13502 (N_13502,N_13363,N_13322);
xnor U13503 (N_13503,N_13250,N_13322);
and U13504 (N_13504,N_13258,N_13385);
nand U13505 (N_13505,N_13360,N_13375);
xor U13506 (N_13506,N_13244,N_13325);
or U13507 (N_13507,N_13326,N_13267);
or U13508 (N_13508,N_13354,N_13238);
and U13509 (N_13509,N_13301,N_13341);
nor U13510 (N_13510,N_13279,N_13390);
and U13511 (N_13511,N_13293,N_13234);
nand U13512 (N_13512,N_13395,N_13222);
nor U13513 (N_13513,N_13350,N_13253);
or U13514 (N_13514,N_13365,N_13287);
or U13515 (N_13515,N_13267,N_13213);
and U13516 (N_13516,N_13226,N_13293);
and U13517 (N_13517,N_13233,N_13342);
and U13518 (N_13518,N_13398,N_13312);
nand U13519 (N_13519,N_13334,N_13344);
or U13520 (N_13520,N_13353,N_13301);
or U13521 (N_13521,N_13348,N_13246);
nor U13522 (N_13522,N_13380,N_13322);
or U13523 (N_13523,N_13266,N_13263);
and U13524 (N_13524,N_13366,N_13352);
nor U13525 (N_13525,N_13372,N_13382);
nand U13526 (N_13526,N_13296,N_13350);
nor U13527 (N_13527,N_13283,N_13263);
or U13528 (N_13528,N_13310,N_13275);
or U13529 (N_13529,N_13379,N_13216);
nand U13530 (N_13530,N_13228,N_13208);
or U13531 (N_13531,N_13253,N_13208);
nor U13532 (N_13532,N_13392,N_13399);
or U13533 (N_13533,N_13335,N_13226);
and U13534 (N_13534,N_13306,N_13254);
or U13535 (N_13535,N_13343,N_13328);
nor U13536 (N_13536,N_13346,N_13332);
nor U13537 (N_13537,N_13248,N_13341);
and U13538 (N_13538,N_13269,N_13373);
nor U13539 (N_13539,N_13200,N_13221);
xnor U13540 (N_13540,N_13385,N_13264);
or U13541 (N_13541,N_13242,N_13337);
and U13542 (N_13542,N_13288,N_13349);
nand U13543 (N_13543,N_13336,N_13380);
xnor U13544 (N_13544,N_13200,N_13327);
or U13545 (N_13545,N_13276,N_13312);
xnor U13546 (N_13546,N_13239,N_13332);
nor U13547 (N_13547,N_13324,N_13339);
or U13548 (N_13548,N_13318,N_13231);
and U13549 (N_13549,N_13311,N_13319);
nor U13550 (N_13550,N_13369,N_13368);
xor U13551 (N_13551,N_13340,N_13228);
xnor U13552 (N_13552,N_13259,N_13305);
nand U13553 (N_13553,N_13279,N_13387);
nor U13554 (N_13554,N_13380,N_13364);
or U13555 (N_13555,N_13287,N_13232);
nor U13556 (N_13556,N_13386,N_13244);
and U13557 (N_13557,N_13271,N_13231);
nand U13558 (N_13558,N_13325,N_13395);
xnor U13559 (N_13559,N_13215,N_13342);
and U13560 (N_13560,N_13256,N_13268);
nor U13561 (N_13561,N_13383,N_13380);
xor U13562 (N_13562,N_13372,N_13237);
and U13563 (N_13563,N_13298,N_13286);
nor U13564 (N_13564,N_13359,N_13222);
nor U13565 (N_13565,N_13348,N_13210);
or U13566 (N_13566,N_13334,N_13353);
nand U13567 (N_13567,N_13349,N_13274);
nor U13568 (N_13568,N_13286,N_13290);
xor U13569 (N_13569,N_13275,N_13339);
nand U13570 (N_13570,N_13215,N_13202);
or U13571 (N_13571,N_13269,N_13238);
nor U13572 (N_13572,N_13268,N_13355);
or U13573 (N_13573,N_13265,N_13351);
xnor U13574 (N_13574,N_13344,N_13200);
xor U13575 (N_13575,N_13255,N_13361);
and U13576 (N_13576,N_13376,N_13275);
nor U13577 (N_13577,N_13392,N_13225);
and U13578 (N_13578,N_13268,N_13376);
xnor U13579 (N_13579,N_13241,N_13382);
nand U13580 (N_13580,N_13224,N_13383);
nor U13581 (N_13581,N_13202,N_13325);
and U13582 (N_13582,N_13277,N_13396);
or U13583 (N_13583,N_13331,N_13271);
and U13584 (N_13584,N_13214,N_13270);
nor U13585 (N_13585,N_13315,N_13230);
and U13586 (N_13586,N_13211,N_13287);
and U13587 (N_13587,N_13392,N_13250);
xnor U13588 (N_13588,N_13361,N_13231);
nor U13589 (N_13589,N_13256,N_13273);
nor U13590 (N_13590,N_13376,N_13311);
nand U13591 (N_13591,N_13241,N_13251);
nor U13592 (N_13592,N_13395,N_13217);
nand U13593 (N_13593,N_13330,N_13212);
and U13594 (N_13594,N_13214,N_13329);
nand U13595 (N_13595,N_13202,N_13344);
and U13596 (N_13596,N_13379,N_13214);
xnor U13597 (N_13597,N_13299,N_13309);
and U13598 (N_13598,N_13332,N_13357);
xnor U13599 (N_13599,N_13275,N_13250);
and U13600 (N_13600,N_13515,N_13401);
nand U13601 (N_13601,N_13479,N_13454);
nand U13602 (N_13602,N_13480,N_13497);
and U13603 (N_13603,N_13566,N_13491);
nor U13604 (N_13604,N_13455,N_13518);
and U13605 (N_13605,N_13409,N_13481);
and U13606 (N_13606,N_13453,N_13505);
and U13607 (N_13607,N_13551,N_13537);
xnor U13608 (N_13608,N_13456,N_13584);
or U13609 (N_13609,N_13511,N_13528);
and U13610 (N_13610,N_13522,N_13460);
or U13611 (N_13611,N_13513,N_13527);
xor U13612 (N_13612,N_13525,N_13533);
xor U13613 (N_13613,N_13432,N_13568);
xnor U13614 (N_13614,N_13427,N_13572);
xor U13615 (N_13615,N_13571,N_13562);
or U13616 (N_13616,N_13557,N_13435);
nor U13617 (N_13617,N_13547,N_13578);
or U13618 (N_13618,N_13514,N_13421);
and U13619 (N_13619,N_13520,N_13532);
xnor U13620 (N_13620,N_13463,N_13471);
xnor U13621 (N_13621,N_13484,N_13508);
nand U13622 (N_13622,N_13443,N_13485);
nor U13623 (N_13623,N_13567,N_13549);
xnor U13624 (N_13624,N_13576,N_13498);
and U13625 (N_13625,N_13403,N_13465);
and U13626 (N_13626,N_13581,N_13441);
xnor U13627 (N_13627,N_13558,N_13534);
or U13628 (N_13628,N_13439,N_13506);
or U13629 (N_13629,N_13544,N_13406);
xnor U13630 (N_13630,N_13478,N_13473);
nor U13631 (N_13631,N_13433,N_13430);
xnor U13632 (N_13632,N_13467,N_13517);
nor U13633 (N_13633,N_13510,N_13414);
or U13634 (N_13634,N_13538,N_13555);
and U13635 (N_13635,N_13540,N_13516);
and U13636 (N_13636,N_13535,N_13599);
or U13637 (N_13637,N_13488,N_13446);
or U13638 (N_13638,N_13472,N_13561);
xor U13639 (N_13639,N_13489,N_13579);
xnor U13640 (N_13640,N_13586,N_13596);
nor U13641 (N_13641,N_13410,N_13422);
and U13642 (N_13642,N_13593,N_13449);
or U13643 (N_13643,N_13529,N_13470);
nor U13644 (N_13644,N_13512,N_13588);
nand U13645 (N_13645,N_13548,N_13483);
or U13646 (N_13646,N_13451,N_13424);
xor U13647 (N_13647,N_13541,N_13493);
nor U13648 (N_13648,N_13477,N_13425);
nor U13649 (N_13649,N_13530,N_13542);
nor U13650 (N_13650,N_13552,N_13560);
nand U13651 (N_13651,N_13595,N_13413);
or U13652 (N_13652,N_13444,N_13504);
xnor U13653 (N_13653,N_13445,N_13415);
or U13654 (N_13654,N_13400,N_13486);
xnor U13655 (N_13655,N_13447,N_13519);
xor U13656 (N_13656,N_13448,N_13587);
nor U13657 (N_13657,N_13407,N_13582);
xnor U13658 (N_13658,N_13553,N_13416);
nand U13659 (N_13659,N_13428,N_13458);
and U13660 (N_13660,N_13402,N_13482);
nor U13661 (N_13661,N_13487,N_13501);
and U13662 (N_13662,N_13412,N_13464);
or U13663 (N_13663,N_13452,N_13591);
xnor U13664 (N_13664,N_13426,N_13592);
or U13665 (N_13665,N_13550,N_13437);
or U13666 (N_13666,N_13503,N_13569);
and U13667 (N_13667,N_13434,N_13502);
nor U13668 (N_13668,N_13418,N_13583);
xor U13669 (N_13669,N_13580,N_13442);
xnor U13670 (N_13670,N_13438,N_13475);
xor U13671 (N_13671,N_13573,N_13594);
xor U13672 (N_13672,N_13590,N_13523);
or U13673 (N_13673,N_13597,N_13490);
and U13674 (N_13674,N_13417,N_13509);
and U13675 (N_13675,N_13536,N_13461);
and U13676 (N_13676,N_13570,N_13495);
nor U13677 (N_13677,N_13546,N_13543);
xnor U13678 (N_13678,N_13429,N_13462);
nor U13679 (N_13679,N_13404,N_13440);
xor U13680 (N_13680,N_13565,N_13419);
nor U13681 (N_13681,N_13524,N_13554);
nand U13682 (N_13682,N_13598,N_13526);
nor U13683 (N_13683,N_13431,N_13457);
and U13684 (N_13684,N_13423,N_13411);
nand U13685 (N_13685,N_13531,N_13408);
or U13686 (N_13686,N_13521,N_13585);
nor U13687 (N_13687,N_13496,N_13436);
and U13688 (N_13688,N_13492,N_13577);
xor U13689 (N_13689,N_13499,N_13507);
and U13690 (N_13690,N_13476,N_13420);
nand U13691 (N_13691,N_13589,N_13494);
or U13692 (N_13692,N_13564,N_13539);
nor U13693 (N_13693,N_13545,N_13500);
nor U13694 (N_13694,N_13556,N_13575);
or U13695 (N_13695,N_13466,N_13563);
and U13696 (N_13696,N_13468,N_13474);
nand U13697 (N_13697,N_13405,N_13574);
nand U13698 (N_13698,N_13559,N_13469);
nand U13699 (N_13699,N_13459,N_13450);
xnor U13700 (N_13700,N_13544,N_13473);
nor U13701 (N_13701,N_13439,N_13435);
or U13702 (N_13702,N_13418,N_13555);
nor U13703 (N_13703,N_13483,N_13577);
xor U13704 (N_13704,N_13592,N_13526);
xor U13705 (N_13705,N_13432,N_13526);
nand U13706 (N_13706,N_13570,N_13405);
nand U13707 (N_13707,N_13499,N_13529);
xor U13708 (N_13708,N_13450,N_13435);
and U13709 (N_13709,N_13400,N_13489);
and U13710 (N_13710,N_13494,N_13582);
or U13711 (N_13711,N_13553,N_13438);
or U13712 (N_13712,N_13434,N_13585);
or U13713 (N_13713,N_13512,N_13545);
and U13714 (N_13714,N_13400,N_13444);
xnor U13715 (N_13715,N_13426,N_13548);
xnor U13716 (N_13716,N_13551,N_13567);
or U13717 (N_13717,N_13437,N_13459);
nand U13718 (N_13718,N_13511,N_13584);
nor U13719 (N_13719,N_13487,N_13563);
nor U13720 (N_13720,N_13515,N_13594);
or U13721 (N_13721,N_13443,N_13467);
nand U13722 (N_13722,N_13474,N_13435);
xnor U13723 (N_13723,N_13543,N_13560);
or U13724 (N_13724,N_13594,N_13536);
xor U13725 (N_13725,N_13596,N_13573);
or U13726 (N_13726,N_13440,N_13500);
nor U13727 (N_13727,N_13445,N_13407);
nor U13728 (N_13728,N_13431,N_13470);
nand U13729 (N_13729,N_13553,N_13429);
and U13730 (N_13730,N_13484,N_13530);
nor U13731 (N_13731,N_13479,N_13573);
nor U13732 (N_13732,N_13406,N_13476);
and U13733 (N_13733,N_13559,N_13561);
nor U13734 (N_13734,N_13555,N_13565);
nor U13735 (N_13735,N_13409,N_13414);
nand U13736 (N_13736,N_13552,N_13522);
and U13737 (N_13737,N_13561,N_13450);
and U13738 (N_13738,N_13406,N_13437);
and U13739 (N_13739,N_13530,N_13407);
or U13740 (N_13740,N_13467,N_13515);
nand U13741 (N_13741,N_13495,N_13474);
xnor U13742 (N_13742,N_13583,N_13580);
or U13743 (N_13743,N_13547,N_13422);
nor U13744 (N_13744,N_13547,N_13579);
or U13745 (N_13745,N_13496,N_13548);
xor U13746 (N_13746,N_13442,N_13520);
and U13747 (N_13747,N_13460,N_13484);
nor U13748 (N_13748,N_13440,N_13461);
or U13749 (N_13749,N_13472,N_13581);
nor U13750 (N_13750,N_13573,N_13562);
and U13751 (N_13751,N_13561,N_13466);
nand U13752 (N_13752,N_13483,N_13587);
xnor U13753 (N_13753,N_13595,N_13460);
nor U13754 (N_13754,N_13489,N_13503);
nand U13755 (N_13755,N_13433,N_13454);
and U13756 (N_13756,N_13404,N_13413);
and U13757 (N_13757,N_13566,N_13542);
nor U13758 (N_13758,N_13420,N_13544);
and U13759 (N_13759,N_13413,N_13420);
xnor U13760 (N_13760,N_13415,N_13416);
and U13761 (N_13761,N_13578,N_13497);
xor U13762 (N_13762,N_13529,N_13537);
and U13763 (N_13763,N_13517,N_13498);
xor U13764 (N_13764,N_13571,N_13558);
xor U13765 (N_13765,N_13436,N_13522);
or U13766 (N_13766,N_13431,N_13454);
xnor U13767 (N_13767,N_13561,N_13497);
nand U13768 (N_13768,N_13592,N_13498);
and U13769 (N_13769,N_13449,N_13586);
xnor U13770 (N_13770,N_13468,N_13576);
nand U13771 (N_13771,N_13598,N_13430);
and U13772 (N_13772,N_13452,N_13411);
and U13773 (N_13773,N_13486,N_13401);
nand U13774 (N_13774,N_13597,N_13553);
nand U13775 (N_13775,N_13488,N_13479);
nor U13776 (N_13776,N_13460,N_13438);
xnor U13777 (N_13777,N_13502,N_13593);
xor U13778 (N_13778,N_13582,N_13544);
or U13779 (N_13779,N_13413,N_13498);
and U13780 (N_13780,N_13428,N_13475);
nand U13781 (N_13781,N_13424,N_13520);
or U13782 (N_13782,N_13587,N_13542);
nand U13783 (N_13783,N_13412,N_13450);
nor U13784 (N_13784,N_13498,N_13560);
and U13785 (N_13785,N_13505,N_13439);
nor U13786 (N_13786,N_13532,N_13450);
xnor U13787 (N_13787,N_13407,N_13490);
and U13788 (N_13788,N_13427,N_13542);
and U13789 (N_13789,N_13433,N_13510);
and U13790 (N_13790,N_13482,N_13565);
and U13791 (N_13791,N_13476,N_13512);
xor U13792 (N_13792,N_13574,N_13593);
and U13793 (N_13793,N_13574,N_13524);
or U13794 (N_13794,N_13542,N_13575);
nor U13795 (N_13795,N_13481,N_13523);
nor U13796 (N_13796,N_13439,N_13495);
nor U13797 (N_13797,N_13534,N_13502);
and U13798 (N_13798,N_13427,N_13433);
nor U13799 (N_13799,N_13574,N_13523);
nor U13800 (N_13800,N_13650,N_13668);
nor U13801 (N_13801,N_13645,N_13623);
nor U13802 (N_13802,N_13766,N_13773);
nor U13803 (N_13803,N_13666,N_13601);
or U13804 (N_13804,N_13711,N_13686);
nand U13805 (N_13805,N_13755,N_13626);
xnor U13806 (N_13806,N_13702,N_13691);
nand U13807 (N_13807,N_13646,N_13606);
nor U13808 (N_13808,N_13659,N_13731);
and U13809 (N_13809,N_13671,N_13776);
and U13810 (N_13810,N_13738,N_13724);
or U13811 (N_13811,N_13628,N_13750);
nor U13812 (N_13812,N_13609,N_13797);
or U13813 (N_13813,N_13665,N_13794);
nand U13814 (N_13814,N_13734,N_13789);
and U13815 (N_13815,N_13743,N_13658);
nor U13816 (N_13816,N_13703,N_13604);
or U13817 (N_13817,N_13726,N_13721);
or U13818 (N_13818,N_13661,N_13669);
or U13819 (N_13819,N_13792,N_13675);
and U13820 (N_13820,N_13602,N_13636);
or U13821 (N_13821,N_13633,N_13660);
and U13822 (N_13822,N_13782,N_13634);
xor U13823 (N_13823,N_13651,N_13764);
or U13824 (N_13824,N_13710,N_13662);
nor U13825 (N_13825,N_13713,N_13676);
nand U13826 (N_13826,N_13617,N_13629);
and U13827 (N_13827,N_13619,N_13765);
xnor U13828 (N_13828,N_13657,N_13689);
or U13829 (N_13829,N_13796,N_13677);
or U13830 (N_13830,N_13655,N_13674);
xnor U13831 (N_13831,N_13732,N_13608);
xor U13832 (N_13832,N_13644,N_13788);
nand U13833 (N_13833,N_13787,N_13762);
xor U13834 (N_13834,N_13699,N_13682);
and U13835 (N_13835,N_13716,N_13652);
nand U13836 (N_13836,N_13620,N_13610);
xnor U13837 (N_13837,N_13740,N_13630);
nor U13838 (N_13838,N_13714,N_13704);
and U13839 (N_13839,N_13763,N_13717);
and U13840 (N_13840,N_13775,N_13778);
or U13841 (N_13841,N_13678,N_13654);
and U13842 (N_13842,N_13745,N_13707);
xor U13843 (N_13843,N_13771,N_13767);
nand U13844 (N_13844,N_13719,N_13748);
nor U13845 (N_13845,N_13725,N_13799);
and U13846 (N_13846,N_13653,N_13643);
or U13847 (N_13847,N_13772,N_13697);
nand U13848 (N_13848,N_13600,N_13624);
nand U13849 (N_13849,N_13733,N_13736);
or U13850 (N_13850,N_13690,N_13605);
nand U13851 (N_13851,N_13780,N_13648);
nand U13852 (N_13852,N_13785,N_13688);
nor U13853 (N_13853,N_13779,N_13708);
and U13854 (N_13854,N_13685,N_13722);
xnor U13855 (N_13855,N_13712,N_13614);
nor U13856 (N_13856,N_13622,N_13761);
and U13857 (N_13857,N_13692,N_13752);
nor U13858 (N_13858,N_13656,N_13786);
and U13859 (N_13859,N_13611,N_13730);
and U13860 (N_13860,N_13663,N_13696);
and U13861 (N_13861,N_13744,N_13798);
xnor U13862 (N_13862,N_13640,N_13681);
xnor U13863 (N_13863,N_13760,N_13757);
and U13864 (N_13864,N_13747,N_13753);
xnor U13865 (N_13865,N_13695,N_13741);
nand U13866 (N_13866,N_13729,N_13720);
nand U13867 (N_13867,N_13672,N_13687);
or U13868 (N_13868,N_13774,N_13737);
xor U13869 (N_13869,N_13700,N_13615);
nand U13870 (N_13870,N_13621,N_13612);
nand U13871 (N_13871,N_13647,N_13607);
or U13872 (N_13872,N_13735,N_13758);
xnor U13873 (N_13873,N_13670,N_13613);
xor U13874 (N_13874,N_13723,N_13698);
nor U13875 (N_13875,N_13632,N_13641);
or U13876 (N_13876,N_13784,N_13751);
nand U13877 (N_13877,N_13705,N_13684);
nor U13878 (N_13878,N_13639,N_13783);
or U13879 (N_13879,N_13664,N_13742);
and U13880 (N_13880,N_13603,N_13625);
nand U13881 (N_13881,N_13739,N_13769);
and U13882 (N_13882,N_13683,N_13749);
or U13883 (N_13883,N_13627,N_13791);
xor U13884 (N_13884,N_13693,N_13795);
xnor U13885 (N_13885,N_13635,N_13694);
nor U13886 (N_13886,N_13718,N_13709);
nor U13887 (N_13887,N_13679,N_13777);
nand U13888 (N_13888,N_13616,N_13618);
and U13889 (N_13889,N_13759,N_13673);
nand U13890 (N_13890,N_13680,N_13706);
and U13891 (N_13891,N_13727,N_13746);
xnor U13892 (N_13892,N_13770,N_13728);
xor U13893 (N_13893,N_13715,N_13790);
xor U13894 (N_13894,N_13754,N_13756);
nand U13895 (N_13895,N_13781,N_13649);
nor U13896 (N_13896,N_13631,N_13642);
or U13897 (N_13897,N_13637,N_13701);
and U13898 (N_13898,N_13667,N_13768);
xor U13899 (N_13899,N_13793,N_13638);
xnor U13900 (N_13900,N_13769,N_13666);
xor U13901 (N_13901,N_13763,N_13704);
nor U13902 (N_13902,N_13771,N_13752);
nor U13903 (N_13903,N_13775,N_13725);
and U13904 (N_13904,N_13781,N_13767);
xnor U13905 (N_13905,N_13785,N_13606);
xor U13906 (N_13906,N_13796,N_13643);
and U13907 (N_13907,N_13686,N_13658);
nor U13908 (N_13908,N_13694,N_13650);
nand U13909 (N_13909,N_13693,N_13666);
xnor U13910 (N_13910,N_13739,N_13678);
or U13911 (N_13911,N_13628,N_13767);
xor U13912 (N_13912,N_13756,N_13603);
nor U13913 (N_13913,N_13647,N_13612);
nor U13914 (N_13914,N_13729,N_13670);
and U13915 (N_13915,N_13697,N_13668);
nor U13916 (N_13916,N_13792,N_13704);
or U13917 (N_13917,N_13663,N_13646);
xnor U13918 (N_13918,N_13649,N_13627);
nand U13919 (N_13919,N_13791,N_13790);
xor U13920 (N_13920,N_13730,N_13700);
and U13921 (N_13921,N_13629,N_13679);
and U13922 (N_13922,N_13615,N_13607);
or U13923 (N_13923,N_13694,N_13662);
xnor U13924 (N_13924,N_13703,N_13764);
nor U13925 (N_13925,N_13746,N_13629);
and U13926 (N_13926,N_13774,N_13760);
or U13927 (N_13927,N_13703,N_13728);
and U13928 (N_13928,N_13682,N_13723);
nor U13929 (N_13929,N_13703,N_13727);
nand U13930 (N_13930,N_13795,N_13671);
xor U13931 (N_13931,N_13749,N_13680);
and U13932 (N_13932,N_13698,N_13681);
or U13933 (N_13933,N_13713,N_13718);
or U13934 (N_13934,N_13655,N_13603);
nor U13935 (N_13935,N_13657,N_13619);
or U13936 (N_13936,N_13604,N_13792);
xor U13937 (N_13937,N_13762,N_13602);
and U13938 (N_13938,N_13740,N_13752);
or U13939 (N_13939,N_13658,N_13703);
or U13940 (N_13940,N_13776,N_13758);
nand U13941 (N_13941,N_13712,N_13669);
xnor U13942 (N_13942,N_13604,N_13736);
or U13943 (N_13943,N_13724,N_13797);
or U13944 (N_13944,N_13750,N_13728);
nor U13945 (N_13945,N_13643,N_13628);
nor U13946 (N_13946,N_13727,N_13797);
or U13947 (N_13947,N_13694,N_13616);
nand U13948 (N_13948,N_13687,N_13767);
nor U13949 (N_13949,N_13760,N_13721);
nand U13950 (N_13950,N_13605,N_13627);
or U13951 (N_13951,N_13700,N_13670);
nand U13952 (N_13952,N_13740,N_13688);
or U13953 (N_13953,N_13713,N_13709);
and U13954 (N_13954,N_13786,N_13664);
nand U13955 (N_13955,N_13769,N_13681);
xor U13956 (N_13956,N_13796,N_13625);
xnor U13957 (N_13957,N_13619,N_13781);
xnor U13958 (N_13958,N_13617,N_13665);
or U13959 (N_13959,N_13610,N_13677);
nand U13960 (N_13960,N_13725,N_13682);
or U13961 (N_13961,N_13693,N_13732);
xor U13962 (N_13962,N_13705,N_13619);
and U13963 (N_13963,N_13649,N_13753);
and U13964 (N_13964,N_13770,N_13645);
nand U13965 (N_13965,N_13614,N_13691);
or U13966 (N_13966,N_13757,N_13741);
xor U13967 (N_13967,N_13747,N_13751);
xnor U13968 (N_13968,N_13657,N_13624);
xor U13969 (N_13969,N_13712,N_13774);
or U13970 (N_13970,N_13696,N_13684);
nor U13971 (N_13971,N_13726,N_13716);
or U13972 (N_13972,N_13613,N_13783);
and U13973 (N_13973,N_13692,N_13714);
and U13974 (N_13974,N_13747,N_13607);
and U13975 (N_13975,N_13640,N_13785);
or U13976 (N_13976,N_13640,N_13613);
xor U13977 (N_13977,N_13622,N_13763);
xor U13978 (N_13978,N_13654,N_13615);
nor U13979 (N_13979,N_13691,N_13615);
and U13980 (N_13980,N_13717,N_13675);
xnor U13981 (N_13981,N_13761,N_13703);
or U13982 (N_13982,N_13699,N_13675);
xnor U13983 (N_13983,N_13704,N_13718);
and U13984 (N_13984,N_13663,N_13796);
nand U13985 (N_13985,N_13620,N_13710);
xnor U13986 (N_13986,N_13657,N_13781);
nor U13987 (N_13987,N_13758,N_13730);
nand U13988 (N_13988,N_13725,N_13771);
nor U13989 (N_13989,N_13633,N_13738);
and U13990 (N_13990,N_13765,N_13741);
xnor U13991 (N_13991,N_13724,N_13621);
nand U13992 (N_13992,N_13775,N_13681);
or U13993 (N_13993,N_13642,N_13641);
xor U13994 (N_13994,N_13768,N_13642);
xnor U13995 (N_13995,N_13637,N_13774);
xnor U13996 (N_13996,N_13639,N_13715);
nor U13997 (N_13997,N_13653,N_13696);
and U13998 (N_13998,N_13723,N_13794);
and U13999 (N_13999,N_13728,N_13674);
nor U14000 (N_14000,N_13913,N_13817);
xor U14001 (N_14001,N_13984,N_13871);
and U14002 (N_14002,N_13907,N_13923);
xnor U14003 (N_14003,N_13902,N_13873);
nand U14004 (N_14004,N_13945,N_13967);
and U14005 (N_14005,N_13827,N_13999);
xor U14006 (N_14006,N_13953,N_13982);
or U14007 (N_14007,N_13892,N_13808);
xor U14008 (N_14008,N_13847,N_13861);
and U14009 (N_14009,N_13851,N_13849);
nand U14010 (N_14010,N_13813,N_13832);
and U14011 (N_14011,N_13826,N_13864);
and U14012 (N_14012,N_13835,N_13891);
nand U14013 (N_14013,N_13990,N_13841);
or U14014 (N_14014,N_13828,N_13981);
or U14015 (N_14015,N_13931,N_13908);
and U14016 (N_14016,N_13854,N_13863);
nand U14017 (N_14017,N_13932,N_13840);
or U14018 (N_14018,N_13852,N_13978);
or U14019 (N_14019,N_13927,N_13882);
and U14020 (N_14020,N_13941,N_13836);
or U14021 (N_14021,N_13874,N_13973);
xnor U14022 (N_14022,N_13918,N_13829);
and U14023 (N_14023,N_13938,N_13821);
or U14024 (N_14024,N_13991,N_13994);
nor U14025 (N_14025,N_13988,N_13911);
nand U14026 (N_14026,N_13860,N_13846);
xnor U14027 (N_14027,N_13905,N_13856);
or U14028 (N_14028,N_13920,N_13879);
xnor U14029 (N_14029,N_13859,N_13816);
and U14030 (N_14030,N_13928,N_13857);
and U14031 (N_14031,N_13899,N_13965);
or U14032 (N_14032,N_13893,N_13807);
nand U14033 (N_14033,N_13818,N_13983);
xor U14034 (N_14034,N_13955,N_13974);
and U14035 (N_14035,N_13940,N_13889);
or U14036 (N_14036,N_13888,N_13848);
and U14037 (N_14037,N_13900,N_13800);
or U14038 (N_14038,N_13964,N_13934);
or U14039 (N_14039,N_13937,N_13987);
nand U14040 (N_14040,N_13867,N_13868);
xor U14041 (N_14041,N_13972,N_13959);
nand U14042 (N_14042,N_13881,N_13930);
nand U14043 (N_14043,N_13947,N_13812);
xor U14044 (N_14044,N_13805,N_13939);
nor U14045 (N_14045,N_13989,N_13912);
nor U14046 (N_14046,N_13949,N_13825);
and U14047 (N_14047,N_13810,N_13995);
nand U14048 (N_14048,N_13942,N_13880);
nand U14049 (N_14049,N_13980,N_13976);
and U14050 (N_14050,N_13890,N_13914);
xor U14051 (N_14051,N_13929,N_13975);
or U14052 (N_14052,N_13977,N_13858);
and U14053 (N_14053,N_13935,N_13996);
and U14054 (N_14054,N_13870,N_13933);
and U14055 (N_14055,N_13993,N_13946);
nor U14056 (N_14056,N_13904,N_13971);
nand U14057 (N_14057,N_13887,N_13869);
and U14058 (N_14058,N_13903,N_13901);
nor U14059 (N_14059,N_13906,N_13992);
nor U14060 (N_14060,N_13804,N_13822);
or U14061 (N_14061,N_13963,N_13998);
or U14062 (N_14062,N_13958,N_13968);
xnor U14063 (N_14063,N_13824,N_13960);
and U14064 (N_14064,N_13910,N_13943);
or U14065 (N_14065,N_13834,N_13866);
nand U14066 (N_14066,N_13970,N_13952);
or U14067 (N_14067,N_13894,N_13957);
and U14068 (N_14068,N_13811,N_13806);
or U14069 (N_14069,N_13844,N_13819);
nand U14070 (N_14070,N_13830,N_13802);
nor U14071 (N_14071,N_13985,N_13919);
xor U14072 (N_14072,N_13916,N_13917);
xor U14073 (N_14073,N_13962,N_13839);
nor U14074 (N_14074,N_13925,N_13886);
nor U14075 (N_14075,N_13809,N_13850);
nor U14076 (N_14076,N_13948,N_13951);
xnor U14077 (N_14077,N_13961,N_13921);
or U14078 (N_14078,N_13954,N_13837);
and U14079 (N_14079,N_13986,N_13997);
or U14080 (N_14080,N_13926,N_13862);
xor U14081 (N_14081,N_13936,N_13803);
and U14082 (N_14082,N_13895,N_13853);
or U14083 (N_14083,N_13842,N_13944);
nor U14084 (N_14084,N_13898,N_13896);
nand U14085 (N_14085,N_13909,N_13875);
and U14086 (N_14086,N_13872,N_13883);
xor U14087 (N_14087,N_13884,N_13979);
and U14088 (N_14088,N_13950,N_13814);
and U14089 (N_14089,N_13838,N_13885);
nor U14090 (N_14090,N_13956,N_13876);
or U14091 (N_14091,N_13915,N_13922);
nand U14092 (N_14092,N_13833,N_13823);
and U14093 (N_14093,N_13966,N_13843);
xnor U14094 (N_14094,N_13897,N_13865);
or U14095 (N_14095,N_13969,N_13815);
xor U14096 (N_14096,N_13855,N_13801);
nand U14097 (N_14097,N_13845,N_13820);
nor U14098 (N_14098,N_13877,N_13831);
and U14099 (N_14099,N_13878,N_13924);
nor U14100 (N_14100,N_13938,N_13961);
nor U14101 (N_14101,N_13819,N_13866);
xor U14102 (N_14102,N_13851,N_13913);
or U14103 (N_14103,N_13803,N_13924);
xor U14104 (N_14104,N_13966,N_13857);
and U14105 (N_14105,N_13889,N_13964);
or U14106 (N_14106,N_13880,N_13879);
xor U14107 (N_14107,N_13986,N_13978);
nor U14108 (N_14108,N_13964,N_13838);
xor U14109 (N_14109,N_13998,N_13909);
nand U14110 (N_14110,N_13977,N_13993);
nor U14111 (N_14111,N_13887,N_13888);
or U14112 (N_14112,N_13896,N_13804);
nand U14113 (N_14113,N_13824,N_13971);
nor U14114 (N_14114,N_13991,N_13952);
and U14115 (N_14115,N_13919,N_13934);
nand U14116 (N_14116,N_13820,N_13899);
nor U14117 (N_14117,N_13936,N_13859);
or U14118 (N_14118,N_13950,N_13819);
nand U14119 (N_14119,N_13947,N_13823);
xnor U14120 (N_14120,N_13857,N_13816);
xor U14121 (N_14121,N_13840,N_13942);
nor U14122 (N_14122,N_13923,N_13857);
xor U14123 (N_14123,N_13895,N_13867);
nor U14124 (N_14124,N_13826,N_13984);
or U14125 (N_14125,N_13986,N_13944);
or U14126 (N_14126,N_13907,N_13838);
and U14127 (N_14127,N_13893,N_13936);
and U14128 (N_14128,N_13893,N_13968);
nand U14129 (N_14129,N_13906,N_13923);
xor U14130 (N_14130,N_13882,N_13960);
nand U14131 (N_14131,N_13931,N_13956);
or U14132 (N_14132,N_13915,N_13979);
and U14133 (N_14133,N_13927,N_13888);
nand U14134 (N_14134,N_13803,N_13986);
nand U14135 (N_14135,N_13894,N_13886);
or U14136 (N_14136,N_13912,N_13973);
nand U14137 (N_14137,N_13850,N_13919);
xor U14138 (N_14138,N_13975,N_13985);
nor U14139 (N_14139,N_13959,N_13828);
xor U14140 (N_14140,N_13935,N_13930);
and U14141 (N_14141,N_13993,N_13894);
or U14142 (N_14142,N_13883,N_13970);
or U14143 (N_14143,N_13819,N_13807);
and U14144 (N_14144,N_13936,N_13999);
and U14145 (N_14145,N_13873,N_13874);
and U14146 (N_14146,N_13820,N_13828);
xnor U14147 (N_14147,N_13846,N_13849);
xor U14148 (N_14148,N_13921,N_13861);
and U14149 (N_14149,N_13906,N_13945);
or U14150 (N_14150,N_13927,N_13853);
or U14151 (N_14151,N_13874,N_13985);
nand U14152 (N_14152,N_13840,N_13834);
and U14153 (N_14153,N_13883,N_13846);
xnor U14154 (N_14154,N_13975,N_13839);
or U14155 (N_14155,N_13899,N_13825);
and U14156 (N_14156,N_13837,N_13899);
xnor U14157 (N_14157,N_13974,N_13930);
or U14158 (N_14158,N_13814,N_13942);
nand U14159 (N_14159,N_13885,N_13925);
and U14160 (N_14160,N_13955,N_13801);
nand U14161 (N_14161,N_13997,N_13894);
or U14162 (N_14162,N_13821,N_13955);
xnor U14163 (N_14163,N_13854,N_13835);
or U14164 (N_14164,N_13821,N_13867);
or U14165 (N_14165,N_13803,N_13932);
nor U14166 (N_14166,N_13957,N_13949);
nand U14167 (N_14167,N_13831,N_13881);
or U14168 (N_14168,N_13966,N_13937);
xnor U14169 (N_14169,N_13839,N_13945);
nor U14170 (N_14170,N_13922,N_13926);
nand U14171 (N_14171,N_13852,N_13953);
xor U14172 (N_14172,N_13930,N_13808);
nor U14173 (N_14173,N_13961,N_13826);
xnor U14174 (N_14174,N_13953,N_13969);
nand U14175 (N_14175,N_13866,N_13871);
nand U14176 (N_14176,N_13805,N_13859);
nand U14177 (N_14177,N_13864,N_13991);
or U14178 (N_14178,N_13810,N_13910);
nor U14179 (N_14179,N_13947,N_13874);
xnor U14180 (N_14180,N_13994,N_13911);
nor U14181 (N_14181,N_13944,N_13975);
xnor U14182 (N_14182,N_13933,N_13972);
and U14183 (N_14183,N_13850,N_13989);
xor U14184 (N_14184,N_13855,N_13872);
nor U14185 (N_14185,N_13901,N_13840);
or U14186 (N_14186,N_13971,N_13885);
nand U14187 (N_14187,N_13873,N_13904);
nand U14188 (N_14188,N_13990,N_13823);
nand U14189 (N_14189,N_13964,N_13946);
nand U14190 (N_14190,N_13967,N_13901);
and U14191 (N_14191,N_13800,N_13805);
nor U14192 (N_14192,N_13970,N_13995);
xnor U14193 (N_14193,N_13887,N_13913);
and U14194 (N_14194,N_13977,N_13841);
and U14195 (N_14195,N_13859,N_13826);
nand U14196 (N_14196,N_13972,N_13846);
and U14197 (N_14197,N_13850,N_13808);
nor U14198 (N_14198,N_13940,N_13858);
nor U14199 (N_14199,N_13835,N_13888);
nand U14200 (N_14200,N_14150,N_14172);
and U14201 (N_14201,N_14021,N_14173);
and U14202 (N_14202,N_14052,N_14031);
xor U14203 (N_14203,N_14198,N_14004);
and U14204 (N_14204,N_14121,N_14103);
nand U14205 (N_14205,N_14066,N_14123);
xnor U14206 (N_14206,N_14026,N_14197);
nand U14207 (N_14207,N_14023,N_14055);
nor U14208 (N_14208,N_14098,N_14072);
and U14209 (N_14209,N_14027,N_14117);
xnor U14210 (N_14210,N_14094,N_14158);
and U14211 (N_14211,N_14115,N_14048);
nor U14212 (N_14212,N_14194,N_14057);
and U14213 (N_14213,N_14028,N_14032);
xnor U14214 (N_14214,N_14065,N_14030);
xnor U14215 (N_14215,N_14081,N_14082);
or U14216 (N_14216,N_14180,N_14167);
nand U14217 (N_14217,N_14073,N_14196);
or U14218 (N_14218,N_14176,N_14064);
xnor U14219 (N_14219,N_14067,N_14079);
xor U14220 (N_14220,N_14168,N_14029);
nand U14221 (N_14221,N_14033,N_14184);
xnor U14222 (N_14222,N_14142,N_14046);
nor U14223 (N_14223,N_14159,N_14022);
or U14224 (N_14224,N_14164,N_14089);
or U14225 (N_14225,N_14140,N_14091);
nor U14226 (N_14226,N_14149,N_14147);
xnor U14227 (N_14227,N_14136,N_14071);
and U14228 (N_14228,N_14043,N_14088);
xnor U14229 (N_14229,N_14144,N_14154);
and U14230 (N_14230,N_14097,N_14036);
nor U14231 (N_14231,N_14077,N_14095);
nor U14232 (N_14232,N_14010,N_14008);
xnor U14233 (N_14233,N_14069,N_14178);
nand U14234 (N_14234,N_14122,N_14135);
or U14235 (N_14235,N_14174,N_14001);
xor U14236 (N_14236,N_14085,N_14177);
and U14237 (N_14237,N_14024,N_14090);
nand U14238 (N_14238,N_14179,N_14160);
or U14239 (N_14239,N_14119,N_14131);
nor U14240 (N_14240,N_14084,N_14041);
nand U14241 (N_14241,N_14059,N_14009);
nand U14242 (N_14242,N_14053,N_14146);
nand U14243 (N_14243,N_14124,N_14037);
xnor U14244 (N_14244,N_14165,N_14025);
or U14245 (N_14245,N_14145,N_14003);
nand U14246 (N_14246,N_14039,N_14019);
or U14247 (N_14247,N_14070,N_14139);
xor U14248 (N_14248,N_14101,N_14083);
xnor U14249 (N_14249,N_14080,N_14186);
or U14250 (N_14250,N_14171,N_14148);
xnor U14251 (N_14251,N_14061,N_14130);
nor U14252 (N_14252,N_14011,N_14014);
nor U14253 (N_14253,N_14141,N_14060);
nor U14254 (N_14254,N_14106,N_14045);
nor U14255 (N_14255,N_14116,N_14040);
nor U14256 (N_14256,N_14181,N_14182);
nor U14257 (N_14257,N_14092,N_14086);
xor U14258 (N_14258,N_14005,N_14020);
nor U14259 (N_14259,N_14120,N_14000);
nand U14260 (N_14260,N_14151,N_14128);
and U14261 (N_14261,N_14109,N_14187);
xnor U14262 (N_14262,N_14015,N_14051);
nor U14263 (N_14263,N_14017,N_14016);
and U14264 (N_14264,N_14102,N_14034);
and U14265 (N_14265,N_14166,N_14087);
nand U14266 (N_14266,N_14035,N_14188);
or U14267 (N_14267,N_14058,N_14138);
and U14268 (N_14268,N_14107,N_14129);
nor U14269 (N_14269,N_14192,N_14161);
nor U14270 (N_14270,N_14133,N_14099);
nand U14271 (N_14271,N_14006,N_14199);
or U14272 (N_14272,N_14185,N_14125);
nand U14273 (N_14273,N_14042,N_14012);
and U14274 (N_14274,N_14074,N_14126);
nand U14275 (N_14275,N_14062,N_14104);
and U14276 (N_14276,N_14183,N_14093);
xor U14277 (N_14277,N_14163,N_14038);
nor U14278 (N_14278,N_14195,N_14156);
nor U14279 (N_14279,N_14162,N_14114);
or U14280 (N_14280,N_14152,N_14134);
xor U14281 (N_14281,N_14100,N_14170);
and U14282 (N_14282,N_14013,N_14175);
or U14283 (N_14283,N_14096,N_14137);
or U14284 (N_14284,N_14047,N_14108);
and U14285 (N_14285,N_14078,N_14127);
or U14286 (N_14286,N_14018,N_14002);
or U14287 (N_14287,N_14049,N_14110);
or U14288 (N_14288,N_14189,N_14056);
xor U14289 (N_14289,N_14155,N_14157);
nand U14290 (N_14290,N_14193,N_14113);
and U14291 (N_14291,N_14044,N_14132);
and U14292 (N_14292,N_14063,N_14105);
nand U14293 (N_14293,N_14118,N_14007);
or U14294 (N_14294,N_14111,N_14169);
nand U14295 (N_14295,N_14153,N_14112);
nor U14296 (N_14296,N_14050,N_14075);
nand U14297 (N_14297,N_14076,N_14191);
and U14298 (N_14298,N_14143,N_14190);
and U14299 (N_14299,N_14068,N_14054);
and U14300 (N_14300,N_14195,N_14015);
nor U14301 (N_14301,N_14188,N_14181);
nand U14302 (N_14302,N_14167,N_14179);
and U14303 (N_14303,N_14153,N_14141);
nor U14304 (N_14304,N_14124,N_14148);
nor U14305 (N_14305,N_14149,N_14044);
xor U14306 (N_14306,N_14193,N_14180);
nand U14307 (N_14307,N_14199,N_14073);
nand U14308 (N_14308,N_14177,N_14086);
and U14309 (N_14309,N_14156,N_14186);
nor U14310 (N_14310,N_14001,N_14152);
or U14311 (N_14311,N_14079,N_14061);
nor U14312 (N_14312,N_14033,N_14147);
and U14313 (N_14313,N_14065,N_14007);
nor U14314 (N_14314,N_14191,N_14090);
nor U14315 (N_14315,N_14075,N_14064);
or U14316 (N_14316,N_14012,N_14057);
nand U14317 (N_14317,N_14126,N_14195);
or U14318 (N_14318,N_14137,N_14121);
xnor U14319 (N_14319,N_14049,N_14094);
xor U14320 (N_14320,N_14011,N_14123);
nor U14321 (N_14321,N_14130,N_14192);
xor U14322 (N_14322,N_14051,N_14172);
nand U14323 (N_14323,N_14199,N_14140);
xnor U14324 (N_14324,N_14124,N_14186);
nor U14325 (N_14325,N_14029,N_14001);
nor U14326 (N_14326,N_14139,N_14073);
or U14327 (N_14327,N_14074,N_14151);
or U14328 (N_14328,N_14026,N_14134);
xor U14329 (N_14329,N_14134,N_14105);
or U14330 (N_14330,N_14172,N_14180);
xor U14331 (N_14331,N_14075,N_14157);
and U14332 (N_14332,N_14174,N_14083);
nor U14333 (N_14333,N_14086,N_14004);
or U14334 (N_14334,N_14030,N_14057);
nor U14335 (N_14335,N_14023,N_14173);
nor U14336 (N_14336,N_14177,N_14111);
or U14337 (N_14337,N_14152,N_14160);
nor U14338 (N_14338,N_14169,N_14171);
and U14339 (N_14339,N_14120,N_14046);
or U14340 (N_14340,N_14068,N_14154);
nor U14341 (N_14341,N_14038,N_14087);
nand U14342 (N_14342,N_14079,N_14131);
nor U14343 (N_14343,N_14114,N_14086);
nor U14344 (N_14344,N_14180,N_14042);
nand U14345 (N_14345,N_14191,N_14117);
nand U14346 (N_14346,N_14089,N_14132);
and U14347 (N_14347,N_14066,N_14031);
xnor U14348 (N_14348,N_14057,N_14032);
xor U14349 (N_14349,N_14004,N_14104);
nor U14350 (N_14350,N_14139,N_14161);
or U14351 (N_14351,N_14131,N_14072);
nand U14352 (N_14352,N_14015,N_14068);
or U14353 (N_14353,N_14141,N_14070);
nor U14354 (N_14354,N_14157,N_14103);
nand U14355 (N_14355,N_14114,N_14011);
nand U14356 (N_14356,N_14198,N_14009);
nand U14357 (N_14357,N_14141,N_14175);
or U14358 (N_14358,N_14171,N_14001);
xor U14359 (N_14359,N_14064,N_14098);
xor U14360 (N_14360,N_14103,N_14182);
and U14361 (N_14361,N_14172,N_14029);
nor U14362 (N_14362,N_14027,N_14191);
nor U14363 (N_14363,N_14136,N_14075);
and U14364 (N_14364,N_14127,N_14085);
and U14365 (N_14365,N_14070,N_14058);
nor U14366 (N_14366,N_14127,N_14064);
xor U14367 (N_14367,N_14006,N_14102);
xor U14368 (N_14368,N_14030,N_14132);
or U14369 (N_14369,N_14071,N_14177);
xnor U14370 (N_14370,N_14168,N_14138);
and U14371 (N_14371,N_14129,N_14007);
or U14372 (N_14372,N_14012,N_14144);
or U14373 (N_14373,N_14093,N_14066);
or U14374 (N_14374,N_14182,N_14195);
nor U14375 (N_14375,N_14068,N_14170);
xnor U14376 (N_14376,N_14131,N_14138);
xor U14377 (N_14377,N_14116,N_14085);
nand U14378 (N_14378,N_14180,N_14083);
or U14379 (N_14379,N_14085,N_14081);
nor U14380 (N_14380,N_14092,N_14051);
or U14381 (N_14381,N_14173,N_14124);
nand U14382 (N_14382,N_14005,N_14147);
or U14383 (N_14383,N_14097,N_14043);
or U14384 (N_14384,N_14116,N_14109);
xnor U14385 (N_14385,N_14189,N_14146);
or U14386 (N_14386,N_14108,N_14168);
xor U14387 (N_14387,N_14060,N_14070);
and U14388 (N_14388,N_14009,N_14095);
xor U14389 (N_14389,N_14105,N_14182);
xor U14390 (N_14390,N_14176,N_14130);
and U14391 (N_14391,N_14055,N_14015);
or U14392 (N_14392,N_14042,N_14119);
nor U14393 (N_14393,N_14047,N_14041);
nand U14394 (N_14394,N_14082,N_14179);
xor U14395 (N_14395,N_14140,N_14081);
nor U14396 (N_14396,N_14029,N_14123);
nor U14397 (N_14397,N_14185,N_14076);
nand U14398 (N_14398,N_14107,N_14093);
or U14399 (N_14399,N_14070,N_14022);
and U14400 (N_14400,N_14227,N_14241);
nand U14401 (N_14401,N_14296,N_14283);
nand U14402 (N_14402,N_14365,N_14262);
xnor U14403 (N_14403,N_14389,N_14315);
or U14404 (N_14404,N_14239,N_14325);
nand U14405 (N_14405,N_14361,N_14251);
or U14406 (N_14406,N_14379,N_14364);
or U14407 (N_14407,N_14248,N_14203);
and U14408 (N_14408,N_14351,N_14373);
nor U14409 (N_14409,N_14388,N_14369);
nand U14410 (N_14410,N_14356,N_14321);
and U14411 (N_14411,N_14281,N_14391);
and U14412 (N_14412,N_14270,N_14371);
xnor U14413 (N_14413,N_14316,N_14244);
nand U14414 (N_14414,N_14257,N_14243);
nor U14415 (N_14415,N_14255,N_14218);
and U14416 (N_14416,N_14215,N_14287);
xor U14417 (N_14417,N_14383,N_14336);
xor U14418 (N_14418,N_14392,N_14233);
nand U14419 (N_14419,N_14342,N_14224);
nor U14420 (N_14420,N_14355,N_14363);
and U14421 (N_14421,N_14252,N_14390);
and U14422 (N_14422,N_14204,N_14393);
nand U14423 (N_14423,N_14396,N_14220);
xnor U14424 (N_14424,N_14367,N_14305);
or U14425 (N_14425,N_14311,N_14293);
or U14426 (N_14426,N_14250,N_14275);
or U14427 (N_14427,N_14308,N_14231);
or U14428 (N_14428,N_14228,N_14352);
and U14429 (N_14429,N_14346,N_14205);
or U14430 (N_14430,N_14286,N_14278);
nor U14431 (N_14431,N_14242,N_14207);
or U14432 (N_14432,N_14282,N_14302);
xnor U14433 (N_14433,N_14214,N_14211);
and U14434 (N_14434,N_14345,N_14304);
xor U14435 (N_14435,N_14277,N_14290);
or U14436 (N_14436,N_14382,N_14294);
nor U14437 (N_14437,N_14347,N_14324);
nand U14438 (N_14438,N_14366,N_14377);
nand U14439 (N_14439,N_14263,N_14333);
xnor U14440 (N_14440,N_14354,N_14387);
and U14441 (N_14441,N_14232,N_14238);
and U14442 (N_14442,N_14398,N_14253);
nor U14443 (N_14443,N_14339,N_14299);
nor U14444 (N_14444,N_14301,N_14279);
or U14445 (N_14445,N_14213,N_14353);
nor U14446 (N_14446,N_14284,N_14269);
nor U14447 (N_14447,N_14378,N_14318);
or U14448 (N_14448,N_14313,N_14246);
or U14449 (N_14449,N_14298,N_14223);
xor U14450 (N_14450,N_14384,N_14376);
xor U14451 (N_14451,N_14261,N_14394);
and U14452 (N_14452,N_14285,N_14289);
nor U14453 (N_14453,N_14327,N_14349);
nor U14454 (N_14454,N_14288,N_14350);
and U14455 (N_14455,N_14303,N_14222);
nand U14456 (N_14456,N_14397,N_14306);
xnor U14457 (N_14457,N_14271,N_14337);
and U14458 (N_14458,N_14341,N_14276);
nand U14459 (N_14459,N_14343,N_14309);
xor U14460 (N_14460,N_14260,N_14338);
nor U14461 (N_14461,N_14219,N_14280);
nand U14462 (N_14462,N_14344,N_14358);
or U14463 (N_14463,N_14374,N_14320);
nand U14464 (N_14464,N_14359,N_14297);
or U14465 (N_14465,N_14335,N_14259);
or U14466 (N_14466,N_14330,N_14216);
nand U14467 (N_14467,N_14399,N_14340);
xor U14468 (N_14468,N_14368,N_14334);
and U14469 (N_14469,N_14200,N_14221);
xnor U14470 (N_14470,N_14319,N_14362);
nor U14471 (N_14471,N_14236,N_14249);
nor U14472 (N_14472,N_14385,N_14209);
nand U14473 (N_14473,N_14395,N_14292);
xnor U14474 (N_14474,N_14332,N_14386);
or U14475 (N_14475,N_14234,N_14317);
nand U14476 (N_14476,N_14230,N_14264);
nor U14477 (N_14477,N_14273,N_14326);
xor U14478 (N_14478,N_14217,N_14323);
nand U14479 (N_14479,N_14307,N_14375);
and U14480 (N_14480,N_14210,N_14266);
xor U14481 (N_14481,N_14322,N_14295);
and U14482 (N_14482,N_14331,N_14380);
nor U14483 (N_14483,N_14372,N_14256);
nand U14484 (N_14484,N_14247,N_14237);
nor U14485 (N_14485,N_14267,N_14226);
nand U14486 (N_14486,N_14312,N_14348);
nand U14487 (N_14487,N_14208,N_14300);
xnor U14488 (N_14488,N_14225,N_14254);
or U14489 (N_14489,N_14314,N_14360);
nand U14490 (N_14490,N_14229,N_14370);
or U14491 (N_14491,N_14202,N_14268);
xnor U14492 (N_14492,N_14265,N_14381);
and U14493 (N_14493,N_14310,N_14328);
or U14494 (N_14494,N_14240,N_14258);
xnor U14495 (N_14495,N_14357,N_14272);
and U14496 (N_14496,N_14245,N_14212);
nand U14497 (N_14497,N_14291,N_14201);
and U14498 (N_14498,N_14206,N_14235);
nand U14499 (N_14499,N_14274,N_14329);
nand U14500 (N_14500,N_14343,N_14374);
nor U14501 (N_14501,N_14357,N_14278);
or U14502 (N_14502,N_14323,N_14368);
nor U14503 (N_14503,N_14314,N_14364);
and U14504 (N_14504,N_14216,N_14241);
or U14505 (N_14505,N_14374,N_14206);
or U14506 (N_14506,N_14357,N_14378);
xor U14507 (N_14507,N_14325,N_14393);
xor U14508 (N_14508,N_14369,N_14337);
nand U14509 (N_14509,N_14359,N_14222);
and U14510 (N_14510,N_14234,N_14387);
and U14511 (N_14511,N_14338,N_14214);
nor U14512 (N_14512,N_14288,N_14212);
or U14513 (N_14513,N_14256,N_14351);
nor U14514 (N_14514,N_14389,N_14279);
nor U14515 (N_14515,N_14336,N_14311);
xor U14516 (N_14516,N_14243,N_14240);
xnor U14517 (N_14517,N_14233,N_14283);
nand U14518 (N_14518,N_14305,N_14210);
and U14519 (N_14519,N_14342,N_14301);
or U14520 (N_14520,N_14260,N_14289);
and U14521 (N_14521,N_14395,N_14369);
nand U14522 (N_14522,N_14261,N_14284);
nand U14523 (N_14523,N_14317,N_14385);
and U14524 (N_14524,N_14229,N_14319);
nor U14525 (N_14525,N_14388,N_14303);
or U14526 (N_14526,N_14365,N_14372);
nor U14527 (N_14527,N_14392,N_14361);
nor U14528 (N_14528,N_14228,N_14296);
xnor U14529 (N_14529,N_14301,N_14254);
xor U14530 (N_14530,N_14265,N_14333);
and U14531 (N_14531,N_14357,N_14370);
or U14532 (N_14532,N_14214,N_14285);
xnor U14533 (N_14533,N_14206,N_14347);
and U14534 (N_14534,N_14293,N_14295);
nor U14535 (N_14535,N_14398,N_14291);
and U14536 (N_14536,N_14298,N_14301);
or U14537 (N_14537,N_14298,N_14363);
or U14538 (N_14538,N_14341,N_14295);
or U14539 (N_14539,N_14387,N_14389);
nand U14540 (N_14540,N_14332,N_14288);
xor U14541 (N_14541,N_14261,N_14320);
nand U14542 (N_14542,N_14203,N_14326);
nor U14543 (N_14543,N_14314,N_14313);
nand U14544 (N_14544,N_14231,N_14230);
nand U14545 (N_14545,N_14399,N_14295);
xor U14546 (N_14546,N_14248,N_14366);
xor U14547 (N_14547,N_14235,N_14333);
nor U14548 (N_14548,N_14378,N_14297);
or U14549 (N_14549,N_14252,N_14217);
xnor U14550 (N_14550,N_14340,N_14221);
nand U14551 (N_14551,N_14285,N_14251);
or U14552 (N_14552,N_14271,N_14256);
xnor U14553 (N_14553,N_14222,N_14336);
nor U14554 (N_14554,N_14389,N_14211);
and U14555 (N_14555,N_14291,N_14290);
xor U14556 (N_14556,N_14261,N_14209);
nand U14557 (N_14557,N_14213,N_14351);
or U14558 (N_14558,N_14386,N_14374);
xnor U14559 (N_14559,N_14211,N_14371);
xnor U14560 (N_14560,N_14280,N_14334);
or U14561 (N_14561,N_14234,N_14289);
and U14562 (N_14562,N_14209,N_14357);
nor U14563 (N_14563,N_14366,N_14294);
nor U14564 (N_14564,N_14301,N_14350);
nand U14565 (N_14565,N_14212,N_14349);
nand U14566 (N_14566,N_14220,N_14371);
xor U14567 (N_14567,N_14399,N_14240);
or U14568 (N_14568,N_14249,N_14347);
and U14569 (N_14569,N_14210,N_14203);
or U14570 (N_14570,N_14282,N_14363);
nor U14571 (N_14571,N_14394,N_14295);
nor U14572 (N_14572,N_14337,N_14267);
nor U14573 (N_14573,N_14286,N_14375);
nand U14574 (N_14574,N_14284,N_14250);
or U14575 (N_14575,N_14262,N_14273);
and U14576 (N_14576,N_14237,N_14228);
nand U14577 (N_14577,N_14290,N_14246);
and U14578 (N_14578,N_14308,N_14274);
nand U14579 (N_14579,N_14350,N_14342);
and U14580 (N_14580,N_14351,N_14301);
nor U14581 (N_14581,N_14213,N_14239);
and U14582 (N_14582,N_14224,N_14372);
nor U14583 (N_14583,N_14295,N_14208);
nand U14584 (N_14584,N_14349,N_14369);
and U14585 (N_14585,N_14372,N_14344);
nand U14586 (N_14586,N_14208,N_14354);
nand U14587 (N_14587,N_14385,N_14213);
nand U14588 (N_14588,N_14223,N_14249);
nand U14589 (N_14589,N_14219,N_14390);
or U14590 (N_14590,N_14214,N_14363);
nor U14591 (N_14591,N_14252,N_14315);
xnor U14592 (N_14592,N_14263,N_14378);
nor U14593 (N_14593,N_14334,N_14307);
nand U14594 (N_14594,N_14305,N_14358);
nor U14595 (N_14595,N_14318,N_14213);
and U14596 (N_14596,N_14369,N_14309);
nand U14597 (N_14597,N_14210,N_14375);
xnor U14598 (N_14598,N_14249,N_14378);
or U14599 (N_14599,N_14337,N_14316);
and U14600 (N_14600,N_14437,N_14587);
and U14601 (N_14601,N_14554,N_14475);
xor U14602 (N_14602,N_14426,N_14532);
xnor U14603 (N_14603,N_14581,N_14534);
or U14604 (N_14604,N_14521,N_14570);
nor U14605 (N_14605,N_14588,N_14543);
nor U14606 (N_14606,N_14580,N_14419);
and U14607 (N_14607,N_14582,N_14486);
nand U14608 (N_14608,N_14523,N_14423);
xnor U14609 (N_14609,N_14432,N_14509);
and U14610 (N_14610,N_14415,N_14411);
xnor U14611 (N_14611,N_14453,N_14577);
xor U14612 (N_14612,N_14428,N_14400);
xor U14613 (N_14613,N_14545,N_14476);
and U14614 (N_14614,N_14540,N_14406);
and U14615 (N_14615,N_14416,N_14535);
or U14616 (N_14616,N_14434,N_14562);
or U14617 (N_14617,N_14538,N_14592);
nand U14618 (N_14618,N_14493,N_14414);
xnor U14619 (N_14619,N_14441,N_14550);
and U14620 (N_14620,N_14433,N_14444);
xnor U14621 (N_14621,N_14422,N_14408);
nor U14622 (N_14622,N_14561,N_14527);
nor U14623 (N_14623,N_14492,N_14495);
xor U14624 (N_14624,N_14496,N_14478);
nor U14625 (N_14625,N_14536,N_14481);
nand U14626 (N_14626,N_14553,N_14514);
nand U14627 (N_14627,N_14460,N_14508);
xor U14628 (N_14628,N_14515,N_14407);
and U14629 (N_14629,N_14436,N_14420);
nand U14630 (N_14630,N_14404,N_14524);
and U14631 (N_14631,N_14499,N_14502);
or U14632 (N_14632,N_14425,N_14480);
xnor U14633 (N_14633,N_14410,N_14551);
nand U14634 (N_14634,N_14468,N_14572);
or U14635 (N_14635,N_14442,N_14576);
or U14636 (N_14636,N_14517,N_14528);
or U14637 (N_14637,N_14405,N_14511);
nand U14638 (N_14638,N_14457,N_14547);
and U14639 (N_14639,N_14539,N_14563);
or U14640 (N_14640,N_14461,N_14503);
or U14641 (N_14641,N_14459,N_14465);
and U14642 (N_14642,N_14599,N_14526);
or U14643 (N_14643,N_14421,N_14424);
xor U14644 (N_14644,N_14567,N_14485);
nor U14645 (N_14645,N_14586,N_14418);
xnor U14646 (N_14646,N_14578,N_14491);
nor U14647 (N_14647,N_14546,N_14525);
nand U14648 (N_14648,N_14564,N_14552);
xnor U14649 (N_14649,N_14470,N_14593);
or U14650 (N_14650,N_14565,N_14591);
nor U14651 (N_14651,N_14589,N_14575);
or U14652 (N_14652,N_14439,N_14448);
nor U14653 (N_14653,N_14450,N_14574);
and U14654 (N_14654,N_14462,N_14573);
or U14655 (N_14655,N_14440,N_14529);
or U14656 (N_14656,N_14500,N_14598);
and U14657 (N_14657,N_14438,N_14568);
and U14658 (N_14658,N_14544,N_14473);
nor U14659 (N_14659,N_14445,N_14472);
xor U14660 (N_14660,N_14412,N_14447);
and U14661 (N_14661,N_14519,N_14594);
nand U14662 (N_14662,N_14571,N_14510);
xor U14663 (N_14663,N_14464,N_14559);
and U14664 (N_14664,N_14474,N_14531);
nor U14665 (N_14665,N_14401,N_14555);
nor U14666 (N_14666,N_14417,N_14467);
and U14667 (N_14667,N_14548,N_14530);
nor U14668 (N_14668,N_14490,N_14482);
and U14669 (N_14669,N_14449,N_14579);
nand U14670 (N_14670,N_14452,N_14516);
xnor U14671 (N_14671,N_14557,N_14466);
nor U14672 (N_14672,N_14505,N_14584);
and U14673 (N_14673,N_14446,N_14487);
xor U14674 (N_14674,N_14596,N_14597);
xnor U14675 (N_14675,N_14463,N_14512);
and U14676 (N_14676,N_14471,N_14455);
and U14677 (N_14677,N_14513,N_14409);
and U14678 (N_14678,N_14483,N_14520);
nor U14679 (N_14679,N_14590,N_14541);
or U14680 (N_14680,N_14518,N_14507);
nand U14681 (N_14681,N_14498,N_14506);
nand U14682 (N_14682,N_14542,N_14585);
and U14683 (N_14683,N_14458,N_14556);
nor U14684 (N_14684,N_14413,N_14583);
xor U14685 (N_14685,N_14469,N_14427);
or U14686 (N_14686,N_14477,N_14560);
and U14687 (N_14687,N_14488,N_14569);
and U14688 (N_14688,N_14435,N_14558);
xor U14689 (N_14689,N_14402,N_14537);
xnor U14690 (N_14690,N_14403,N_14454);
or U14691 (N_14691,N_14456,N_14430);
or U14692 (N_14692,N_14522,N_14566);
and U14693 (N_14693,N_14494,N_14549);
or U14694 (N_14694,N_14504,N_14429);
and U14695 (N_14695,N_14431,N_14484);
nand U14696 (N_14696,N_14501,N_14479);
or U14697 (N_14697,N_14497,N_14533);
xnor U14698 (N_14698,N_14443,N_14489);
nor U14699 (N_14699,N_14595,N_14451);
nand U14700 (N_14700,N_14518,N_14550);
xnor U14701 (N_14701,N_14416,N_14565);
nor U14702 (N_14702,N_14507,N_14578);
xor U14703 (N_14703,N_14491,N_14538);
nand U14704 (N_14704,N_14567,N_14424);
xor U14705 (N_14705,N_14494,N_14554);
nand U14706 (N_14706,N_14565,N_14491);
nand U14707 (N_14707,N_14594,N_14580);
nor U14708 (N_14708,N_14583,N_14450);
nand U14709 (N_14709,N_14570,N_14497);
xnor U14710 (N_14710,N_14547,N_14430);
nand U14711 (N_14711,N_14436,N_14501);
or U14712 (N_14712,N_14520,N_14471);
or U14713 (N_14713,N_14479,N_14453);
nor U14714 (N_14714,N_14515,N_14546);
nand U14715 (N_14715,N_14534,N_14477);
nor U14716 (N_14716,N_14453,N_14473);
nor U14717 (N_14717,N_14562,N_14554);
nand U14718 (N_14718,N_14437,N_14453);
nand U14719 (N_14719,N_14571,N_14578);
or U14720 (N_14720,N_14504,N_14446);
nand U14721 (N_14721,N_14444,N_14406);
and U14722 (N_14722,N_14567,N_14558);
or U14723 (N_14723,N_14484,N_14543);
nand U14724 (N_14724,N_14527,N_14574);
and U14725 (N_14725,N_14425,N_14409);
nand U14726 (N_14726,N_14534,N_14564);
xnor U14727 (N_14727,N_14545,N_14500);
and U14728 (N_14728,N_14429,N_14579);
xor U14729 (N_14729,N_14420,N_14587);
and U14730 (N_14730,N_14515,N_14539);
nand U14731 (N_14731,N_14551,N_14498);
and U14732 (N_14732,N_14562,N_14525);
or U14733 (N_14733,N_14545,N_14410);
nand U14734 (N_14734,N_14525,N_14566);
or U14735 (N_14735,N_14483,N_14514);
nor U14736 (N_14736,N_14468,N_14423);
or U14737 (N_14737,N_14486,N_14554);
nor U14738 (N_14738,N_14496,N_14499);
nand U14739 (N_14739,N_14431,N_14443);
xor U14740 (N_14740,N_14447,N_14406);
and U14741 (N_14741,N_14597,N_14559);
or U14742 (N_14742,N_14572,N_14452);
nand U14743 (N_14743,N_14495,N_14528);
nand U14744 (N_14744,N_14527,N_14490);
nand U14745 (N_14745,N_14494,N_14568);
nor U14746 (N_14746,N_14596,N_14481);
xor U14747 (N_14747,N_14456,N_14475);
and U14748 (N_14748,N_14586,N_14411);
xor U14749 (N_14749,N_14433,N_14577);
and U14750 (N_14750,N_14562,N_14530);
nand U14751 (N_14751,N_14468,N_14460);
nand U14752 (N_14752,N_14544,N_14459);
nand U14753 (N_14753,N_14482,N_14477);
or U14754 (N_14754,N_14542,N_14574);
and U14755 (N_14755,N_14470,N_14506);
and U14756 (N_14756,N_14528,N_14401);
nand U14757 (N_14757,N_14523,N_14434);
or U14758 (N_14758,N_14424,N_14405);
and U14759 (N_14759,N_14415,N_14461);
nand U14760 (N_14760,N_14536,N_14438);
or U14761 (N_14761,N_14522,N_14430);
nand U14762 (N_14762,N_14404,N_14578);
nor U14763 (N_14763,N_14567,N_14578);
or U14764 (N_14764,N_14537,N_14587);
xnor U14765 (N_14765,N_14404,N_14483);
or U14766 (N_14766,N_14407,N_14429);
or U14767 (N_14767,N_14487,N_14482);
or U14768 (N_14768,N_14471,N_14580);
nor U14769 (N_14769,N_14425,N_14448);
nand U14770 (N_14770,N_14474,N_14553);
or U14771 (N_14771,N_14498,N_14477);
and U14772 (N_14772,N_14487,N_14413);
nor U14773 (N_14773,N_14482,N_14522);
or U14774 (N_14774,N_14537,N_14522);
xor U14775 (N_14775,N_14433,N_14569);
nor U14776 (N_14776,N_14582,N_14415);
nor U14777 (N_14777,N_14563,N_14553);
xnor U14778 (N_14778,N_14410,N_14487);
or U14779 (N_14779,N_14543,N_14564);
or U14780 (N_14780,N_14540,N_14598);
and U14781 (N_14781,N_14443,N_14579);
and U14782 (N_14782,N_14520,N_14536);
or U14783 (N_14783,N_14423,N_14515);
nand U14784 (N_14784,N_14457,N_14599);
and U14785 (N_14785,N_14584,N_14509);
nand U14786 (N_14786,N_14426,N_14460);
and U14787 (N_14787,N_14542,N_14524);
nand U14788 (N_14788,N_14467,N_14492);
and U14789 (N_14789,N_14570,N_14454);
xor U14790 (N_14790,N_14551,N_14495);
or U14791 (N_14791,N_14541,N_14598);
and U14792 (N_14792,N_14506,N_14523);
or U14793 (N_14793,N_14551,N_14413);
nand U14794 (N_14794,N_14418,N_14550);
nor U14795 (N_14795,N_14416,N_14476);
nor U14796 (N_14796,N_14581,N_14583);
or U14797 (N_14797,N_14495,N_14549);
or U14798 (N_14798,N_14463,N_14423);
nor U14799 (N_14799,N_14422,N_14434);
nor U14800 (N_14800,N_14753,N_14781);
and U14801 (N_14801,N_14794,N_14770);
and U14802 (N_14802,N_14752,N_14746);
or U14803 (N_14803,N_14774,N_14749);
xnor U14804 (N_14804,N_14674,N_14762);
and U14805 (N_14805,N_14754,N_14757);
or U14806 (N_14806,N_14679,N_14663);
nand U14807 (N_14807,N_14645,N_14722);
nor U14808 (N_14808,N_14783,N_14650);
or U14809 (N_14809,N_14710,N_14793);
nand U14810 (N_14810,N_14639,N_14615);
nand U14811 (N_14811,N_14718,N_14621);
or U14812 (N_14812,N_14622,N_14692);
xor U14813 (N_14813,N_14619,N_14716);
xnor U14814 (N_14814,N_14741,N_14703);
or U14815 (N_14815,N_14792,N_14728);
nand U14816 (N_14816,N_14667,N_14785);
xor U14817 (N_14817,N_14705,N_14763);
xor U14818 (N_14818,N_14613,N_14605);
nand U14819 (N_14819,N_14623,N_14702);
or U14820 (N_14820,N_14744,N_14648);
nor U14821 (N_14821,N_14651,N_14712);
nor U14822 (N_14822,N_14726,N_14777);
nor U14823 (N_14823,N_14796,N_14609);
xnor U14824 (N_14824,N_14683,N_14698);
nor U14825 (N_14825,N_14771,N_14638);
nand U14826 (N_14826,N_14682,N_14656);
and U14827 (N_14827,N_14799,N_14734);
and U14828 (N_14828,N_14617,N_14695);
nand U14829 (N_14829,N_14798,N_14606);
nand U14830 (N_14830,N_14769,N_14602);
nor U14831 (N_14831,N_14611,N_14701);
or U14832 (N_14832,N_14659,N_14642);
xor U14833 (N_14833,N_14664,N_14691);
and U14834 (N_14834,N_14790,N_14677);
nand U14835 (N_14835,N_14748,N_14687);
or U14836 (N_14836,N_14612,N_14704);
and U14837 (N_14837,N_14660,N_14626);
and U14838 (N_14838,N_14779,N_14789);
nand U14839 (N_14839,N_14782,N_14665);
xor U14840 (N_14840,N_14707,N_14747);
xnor U14841 (N_14841,N_14733,N_14641);
xor U14842 (N_14842,N_14644,N_14717);
xor U14843 (N_14843,N_14773,N_14647);
or U14844 (N_14844,N_14666,N_14624);
or U14845 (N_14845,N_14678,N_14689);
nand U14846 (N_14846,N_14618,N_14725);
nor U14847 (N_14847,N_14672,N_14696);
or U14848 (N_14848,N_14751,N_14766);
or U14849 (N_14849,N_14632,N_14688);
nor U14850 (N_14850,N_14727,N_14699);
nand U14851 (N_14851,N_14742,N_14649);
xnor U14852 (N_14852,N_14608,N_14738);
nand U14853 (N_14853,N_14604,N_14690);
or U14854 (N_14854,N_14640,N_14765);
nor U14855 (N_14855,N_14700,N_14634);
nor U14856 (N_14856,N_14711,N_14631);
or U14857 (N_14857,N_14643,N_14750);
nor U14858 (N_14858,N_14708,N_14732);
or U14859 (N_14859,N_14715,N_14670);
nand U14860 (N_14860,N_14720,N_14668);
nand U14861 (N_14861,N_14614,N_14795);
xor U14862 (N_14862,N_14637,N_14697);
and U14863 (N_14863,N_14719,N_14714);
nand U14864 (N_14864,N_14654,N_14646);
nand U14865 (N_14865,N_14778,N_14709);
and U14866 (N_14866,N_14764,N_14610);
nor U14867 (N_14867,N_14657,N_14603);
xnor U14868 (N_14868,N_14693,N_14772);
nor U14869 (N_14869,N_14731,N_14635);
nor U14870 (N_14870,N_14784,N_14780);
nand U14871 (N_14871,N_14745,N_14758);
and U14872 (N_14872,N_14787,N_14655);
and U14873 (N_14873,N_14601,N_14627);
nor U14874 (N_14874,N_14776,N_14661);
xnor U14875 (N_14875,N_14723,N_14729);
nand U14876 (N_14876,N_14761,N_14652);
nor U14877 (N_14877,N_14686,N_14673);
xor U14878 (N_14878,N_14600,N_14658);
nand U14879 (N_14879,N_14788,N_14736);
and U14880 (N_14880,N_14797,N_14767);
xnor U14881 (N_14881,N_14636,N_14760);
or U14882 (N_14882,N_14629,N_14724);
xor U14883 (N_14883,N_14713,N_14740);
or U14884 (N_14884,N_14633,N_14625);
nor U14885 (N_14885,N_14786,N_14680);
xnor U14886 (N_14886,N_14721,N_14620);
nand U14887 (N_14887,N_14653,N_14755);
nor U14888 (N_14888,N_14768,N_14775);
and U14889 (N_14889,N_14676,N_14681);
and U14890 (N_14890,N_14669,N_14739);
nand U14891 (N_14891,N_14684,N_14671);
and U14892 (N_14892,N_14756,N_14759);
nand U14893 (N_14893,N_14616,N_14630);
and U14894 (N_14894,N_14730,N_14694);
and U14895 (N_14895,N_14685,N_14628);
and U14896 (N_14896,N_14791,N_14737);
nor U14897 (N_14897,N_14675,N_14706);
nand U14898 (N_14898,N_14743,N_14662);
or U14899 (N_14899,N_14607,N_14735);
nand U14900 (N_14900,N_14776,N_14735);
nor U14901 (N_14901,N_14675,N_14682);
xnor U14902 (N_14902,N_14609,N_14647);
or U14903 (N_14903,N_14718,N_14701);
and U14904 (N_14904,N_14741,N_14624);
or U14905 (N_14905,N_14640,N_14775);
and U14906 (N_14906,N_14749,N_14602);
nand U14907 (N_14907,N_14763,N_14725);
and U14908 (N_14908,N_14660,N_14652);
or U14909 (N_14909,N_14746,N_14631);
and U14910 (N_14910,N_14656,N_14732);
and U14911 (N_14911,N_14708,N_14743);
or U14912 (N_14912,N_14713,N_14622);
and U14913 (N_14913,N_14689,N_14621);
and U14914 (N_14914,N_14784,N_14695);
or U14915 (N_14915,N_14706,N_14722);
and U14916 (N_14916,N_14780,N_14703);
xor U14917 (N_14917,N_14650,N_14635);
xnor U14918 (N_14918,N_14774,N_14721);
nand U14919 (N_14919,N_14740,N_14782);
and U14920 (N_14920,N_14756,N_14700);
or U14921 (N_14921,N_14690,N_14796);
nand U14922 (N_14922,N_14725,N_14721);
xor U14923 (N_14923,N_14602,N_14617);
nand U14924 (N_14924,N_14729,N_14722);
and U14925 (N_14925,N_14779,N_14702);
and U14926 (N_14926,N_14727,N_14631);
nor U14927 (N_14927,N_14700,N_14751);
and U14928 (N_14928,N_14687,N_14693);
or U14929 (N_14929,N_14630,N_14707);
nand U14930 (N_14930,N_14601,N_14634);
and U14931 (N_14931,N_14605,N_14614);
and U14932 (N_14932,N_14625,N_14711);
nand U14933 (N_14933,N_14608,N_14757);
and U14934 (N_14934,N_14789,N_14743);
and U14935 (N_14935,N_14780,N_14734);
nor U14936 (N_14936,N_14761,N_14735);
nor U14937 (N_14937,N_14678,N_14639);
or U14938 (N_14938,N_14744,N_14637);
or U14939 (N_14939,N_14683,N_14602);
xor U14940 (N_14940,N_14798,N_14719);
xnor U14941 (N_14941,N_14668,N_14683);
nand U14942 (N_14942,N_14776,N_14789);
xor U14943 (N_14943,N_14649,N_14662);
nand U14944 (N_14944,N_14760,N_14620);
nor U14945 (N_14945,N_14719,N_14679);
or U14946 (N_14946,N_14724,N_14704);
or U14947 (N_14947,N_14781,N_14707);
nand U14948 (N_14948,N_14738,N_14619);
or U14949 (N_14949,N_14662,N_14723);
nand U14950 (N_14950,N_14649,N_14799);
xnor U14951 (N_14951,N_14715,N_14735);
and U14952 (N_14952,N_14669,N_14749);
nor U14953 (N_14953,N_14708,N_14625);
nor U14954 (N_14954,N_14649,N_14704);
or U14955 (N_14955,N_14774,N_14604);
and U14956 (N_14956,N_14760,N_14629);
and U14957 (N_14957,N_14704,N_14668);
and U14958 (N_14958,N_14779,N_14670);
xnor U14959 (N_14959,N_14689,N_14737);
and U14960 (N_14960,N_14714,N_14669);
nand U14961 (N_14961,N_14621,N_14735);
or U14962 (N_14962,N_14723,N_14665);
or U14963 (N_14963,N_14715,N_14658);
nor U14964 (N_14964,N_14693,N_14699);
or U14965 (N_14965,N_14715,N_14661);
xor U14966 (N_14966,N_14645,N_14799);
xor U14967 (N_14967,N_14608,N_14635);
nor U14968 (N_14968,N_14720,N_14698);
and U14969 (N_14969,N_14734,N_14745);
or U14970 (N_14970,N_14712,N_14601);
nand U14971 (N_14971,N_14645,N_14652);
nand U14972 (N_14972,N_14620,N_14785);
nand U14973 (N_14973,N_14677,N_14650);
xor U14974 (N_14974,N_14625,N_14691);
xor U14975 (N_14975,N_14642,N_14611);
nand U14976 (N_14976,N_14753,N_14664);
xor U14977 (N_14977,N_14614,N_14733);
and U14978 (N_14978,N_14713,N_14775);
nand U14979 (N_14979,N_14788,N_14775);
nand U14980 (N_14980,N_14639,N_14773);
xor U14981 (N_14981,N_14603,N_14733);
and U14982 (N_14982,N_14619,N_14721);
nor U14983 (N_14983,N_14797,N_14684);
nand U14984 (N_14984,N_14604,N_14664);
xnor U14985 (N_14985,N_14738,N_14740);
or U14986 (N_14986,N_14756,N_14670);
xnor U14987 (N_14987,N_14728,N_14775);
xnor U14988 (N_14988,N_14600,N_14761);
or U14989 (N_14989,N_14690,N_14793);
and U14990 (N_14990,N_14781,N_14603);
or U14991 (N_14991,N_14795,N_14618);
nor U14992 (N_14992,N_14682,N_14648);
and U14993 (N_14993,N_14670,N_14644);
nor U14994 (N_14994,N_14679,N_14786);
and U14995 (N_14995,N_14618,N_14781);
nand U14996 (N_14996,N_14781,N_14683);
nor U14997 (N_14997,N_14614,N_14630);
or U14998 (N_14998,N_14671,N_14796);
xnor U14999 (N_14999,N_14649,N_14708);
and U15000 (N_15000,N_14883,N_14902);
or U15001 (N_15001,N_14826,N_14928);
or U15002 (N_15002,N_14980,N_14965);
nor U15003 (N_15003,N_14945,N_14802);
nor U15004 (N_15004,N_14946,N_14953);
and U15005 (N_15005,N_14803,N_14874);
and U15006 (N_15006,N_14801,N_14866);
xnor U15007 (N_15007,N_14824,N_14934);
or U15008 (N_15008,N_14811,N_14950);
nand U15009 (N_15009,N_14877,N_14895);
and U15010 (N_15010,N_14920,N_14988);
nand U15011 (N_15011,N_14851,N_14871);
or U15012 (N_15012,N_14807,N_14964);
nor U15013 (N_15013,N_14848,N_14994);
and U15014 (N_15014,N_14918,N_14832);
nor U15015 (N_15015,N_14907,N_14911);
or U15016 (N_15016,N_14843,N_14898);
and U15017 (N_15017,N_14910,N_14815);
xnor U15018 (N_15018,N_14862,N_14927);
nor U15019 (N_15019,N_14809,N_14859);
nand U15020 (N_15020,N_14818,N_14998);
or U15021 (N_15021,N_14925,N_14954);
nor U15022 (N_15022,N_14916,N_14814);
nand U15023 (N_15023,N_14905,N_14880);
nand U15024 (N_15024,N_14960,N_14942);
or U15025 (N_15025,N_14894,N_14888);
xnor U15026 (N_15026,N_14836,N_14924);
xnor U15027 (N_15027,N_14979,N_14992);
nor U15028 (N_15028,N_14921,N_14854);
or U15029 (N_15029,N_14975,N_14829);
xnor U15030 (N_15030,N_14861,N_14878);
or U15031 (N_15031,N_14914,N_14891);
or U15032 (N_15032,N_14837,N_14890);
nand U15033 (N_15033,N_14856,N_14984);
nor U15034 (N_15034,N_14983,N_14899);
and U15035 (N_15035,N_14923,N_14959);
xnor U15036 (N_15036,N_14839,N_14903);
nand U15037 (N_15037,N_14996,N_14932);
or U15038 (N_15038,N_14834,N_14830);
xnor U15039 (N_15039,N_14936,N_14944);
xnor U15040 (N_15040,N_14972,N_14967);
or U15041 (N_15041,N_14971,N_14976);
or U15042 (N_15042,N_14985,N_14886);
nand U15043 (N_15043,N_14987,N_14991);
and U15044 (N_15044,N_14828,N_14947);
nand U15045 (N_15045,N_14840,N_14943);
nor U15046 (N_15046,N_14864,N_14901);
or U15047 (N_15047,N_14847,N_14995);
nand U15048 (N_15048,N_14827,N_14937);
xor U15049 (N_15049,N_14845,N_14821);
nand U15050 (N_15050,N_14889,N_14812);
and U15051 (N_15051,N_14917,N_14966);
nand U15052 (N_15052,N_14969,N_14858);
and U15053 (N_15053,N_14893,N_14838);
xor U15054 (N_15054,N_14974,N_14900);
nor U15055 (N_15055,N_14875,N_14800);
xor U15056 (N_15056,N_14879,N_14813);
nor U15057 (N_15057,N_14844,N_14850);
or U15058 (N_15058,N_14926,N_14908);
nand U15059 (N_15059,N_14948,N_14993);
nor U15060 (N_15060,N_14863,N_14939);
and U15061 (N_15061,N_14931,N_14940);
and U15062 (N_15062,N_14961,N_14892);
and U15063 (N_15063,N_14842,N_14951);
xor U15064 (N_15064,N_14804,N_14805);
or U15065 (N_15065,N_14955,N_14922);
or U15066 (N_15066,N_14904,N_14956);
or U15067 (N_15067,N_14876,N_14881);
or U15068 (N_15068,N_14855,N_14816);
nor U15069 (N_15069,N_14887,N_14825);
xor U15070 (N_15070,N_14873,N_14935);
or U15071 (N_15071,N_14870,N_14957);
and U15072 (N_15072,N_14817,N_14912);
xor U15073 (N_15073,N_14868,N_14819);
xnor U15074 (N_15074,N_14915,N_14882);
or U15075 (N_15075,N_14938,N_14973);
nor U15076 (N_15076,N_14857,N_14913);
and U15077 (N_15077,N_14929,N_14919);
or U15078 (N_15078,N_14835,N_14982);
xnor U15079 (N_15079,N_14906,N_14869);
or U15080 (N_15080,N_14990,N_14823);
xnor U15081 (N_15081,N_14806,N_14909);
nor U15082 (N_15082,N_14930,N_14999);
or U15083 (N_15083,N_14860,N_14841);
nand U15084 (N_15084,N_14970,N_14884);
xnor U15085 (N_15085,N_14933,N_14867);
and U15086 (N_15086,N_14872,N_14896);
nand U15087 (N_15087,N_14852,N_14958);
or U15088 (N_15088,N_14962,N_14977);
nand U15089 (N_15089,N_14989,N_14808);
xor U15090 (N_15090,N_14831,N_14846);
xnor U15091 (N_15091,N_14952,N_14833);
and U15092 (N_15092,N_14849,N_14810);
and U15093 (N_15093,N_14978,N_14968);
nand U15094 (N_15094,N_14963,N_14820);
or U15095 (N_15095,N_14885,N_14949);
nand U15096 (N_15096,N_14853,N_14897);
xor U15097 (N_15097,N_14997,N_14986);
and U15098 (N_15098,N_14865,N_14981);
nand U15099 (N_15099,N_14941,N_14822);
xnor U15100 (N_15100,N_14959,N_14999);
nand U15101 (N_15101,N_14864,N_14944);
nand U15102 (N_15102,N_14876,N_14828);
or U15103 (N_15103,N_14825,N_14897);
nor U15104 (N_15104,N_14930,N_14918);
and U15105 (N_15105,N_14873,N_14924);
or U15106 (N_15106,N_14994,N_14810);
nor U15107 (N_15107,N_14827,N_14814);
and U15108 (N_15108,N_14843,N_14858);
or U15109 (N_15109,N_14805,N_14985);
nand U15110 (N_15110,N_14914,N_14952);
nand U15111 (N_15111,N_14898,N_14899);
xor U15112 (N_15112,N_14992,N_14922);
nor U15113 (N_15113,N_14971,N_14984);
nand U15114 (N_15114,N_14941,N_14902);
xor U15115 (N_15115,N_14868,N_14844);
nand U15116 (N_15116,N_14943,N_14991);
nor U15117 (N_15117,N_14948,N_14938);
or U15118 (N_15118,N_14982,N_14996);
or U15119 (N_15119,N_14905,N_14861);
nand U15120 (N_15120,N_14902,N_14958);
and U15121 (N_15121,N_14924,N_14808);
nand U15122 (N_15122,N_14949,N_14950);
or U15123 (N_15123,N_14931,N_14800);
nor U15124 (N_15124,N_14951,N_14993);
xnor U15125 (N_15125,N_14909,N_14977);
nand U15126 (N_15126,N_14865,N_14856);
and U15127 (N_15127,N_14857,N_14952);
nand U15128 (N_15128,N_14960,N_14878);
nand U15129 (N_15129,N_14846,N_14856);
nand U15130 (N_15130,N_14917,N_14826);
nand U15131 (N_15131,N_14860,N_14970);
nor U15132 (N_15132,N_14904,N_14841);
or U15133 (N_15133,N_14832,N_14970);
or U15134 (N_15134,N_14858,N_14942);
and U15135 (N_15135,N_14921,N_14922);
xor U15136 (N_15136,N_14887,N_14802);
xor U15137 (N_15137,N_14933,N_14916);
and U15138 (N_15138,N_14801,N_14823);
nand U15139 (N_15139,N_14907,N_14924);
nor U15140 (N_15140,N_14866,N_14869);
or U15141 (N_15141,N_14890,N_14917);
or U15142 (N_15142,N_14803,N_14976);
xor U15143 (N_15143,N_14800,N_14881);
or U15144 (N_15144,N_14905,N_14879);
nand U15145 (N_15145,N_14877,N_14846);
and U15146 (N_15146,N_14893,N_14888);
and U15147 (N_15147,N_14891,N_14928);
nor U15148 (N_15148,N_14925,N_14854);
nor U15149 (N_15149,N_14836,N_14943);
or U15150 (N_15150,N_14825,N_14927);
or U15151 (N_15151,N_14892,N_14988);
and U15152 (N_15152,N_14943,N_14918);
nand U15153 (N_15153,N_14889,N_14839);
nand U15154 (N_15154,N_14917,N_14984);
nor U15155 (N_15155,N_14992,N_14938);
nor U15156 (N_15156,N_14804,N_14980);
and U15157 (N_15157,N_14854,N_14800);
and U15158 (N_15158,N_14885,N_14876);
nor U15159 (N_15159,N_14985,N_14978);
xnor U15160 (N_15160,N_14804,N_14914);
xnor U15161 (N_15161,N_14901,N_14839);
and U15162 (N_15162,N_14824,N_14984);
xnor U15163 (N_15163,N_14993,N_14942);
or U15164 (N_15164,N_14924,N_14816);
nor U15165 (N_15165,N_14995,N_14857);
or U15166 (N_15166,N_14955,N_14850);
nand U15167 (N_15167,N_14850,N_14801);
nand U15168 (N_15168,N_14811,N_14832);
and U15169 (N_15169,N_14965,N_14916);
nor U15170 (N_15170,N_14969,N_14973);
nand U15171 (N_15171,N_14823,N_14854);
and U15172 (N_15172,N_14812,N_14882);
xnor U15173 (N_15173,N_14925,N_14841);
nand U15174 (N_15174,N_14875,N_14955);
xor U15175 (N_15175,N_14905,N_14906);
nand U15176 (N_15176,N_14808,N_14882);
nor U15177 (N_15177,N_14811,N_14922);
or U15178 (N_15178,N_14836,N_14977);
nand U15179 (N_15179,N_14882,N_14896);
nand U15180 (N_15180,N_14935,N_14849);
xnor U15181 (N_15181,N_14840,N_14836);
and U15182 (N_15182,N_14827,N_14933);
and U15183 (N_15183,N_14905,N_14941);
or U15184 (N_15184,N_14953,N_14918);
xor U15185 (N_15185,N_14842,N_14929);
and U15186 (N_15186,N_14821,N_14863);
nor U15187 (N_15187,N_14878,N_14915);
and U15188 (N_15188,N_14864,N_14890);
and U15189 (N_15189,N_14861,N_14851);
and U15190 (N_15190,N_14955,N_14874);
and U15191 (N_15191,N_14970,N_14986);
or U15192 (N_15192,N_14885,N_14816);
nor U15193 (N_15193,N_14914,N_14960);
and U15194 (N_15194,N_14968,N_14832);
and U15195 (N_15195,N_14840,N_14928);
nor U15196 (N_15196,N_14940,N_14812);
and U15197 (N_15197,N_14885,N_14833);
and U15198 (N_15198,N_14941,N_14832);
nor U15199 (N_15199,N_14871,N_14870);
nor U15200 (N_15200,N_15047,N_15062);
xnor U15201 (N_15201,N_15100,N_15141);
or U15202 (N_15202,N_15139,N_15165);
or U15203 (N_15203,N_15096,N_15038);
and U15204 (N_15204,N_15164,N_15036);
xor U15205 (N_15205,N_15028,N_15056);
and U15206 (N_15206,N_15173,N_15019);
nand U15207 (N_15207,N_15185,N_15060);
or U15208 (N_15208,N_15107,N_15127);
or U15209 (N_15209,N_15192,N_15188);
or U15210 (N_15210,N_15074,N_15154);
and U15211 (N_15211,N_15018,N_15061);
and U15212 (N_15212,N_15095,N_15104);
nand U15213 (N_15213,N_15042,N_15063);
and U15214 (N_15214,N_15172,N_15119);
nor U15215 (N_15215,N_15026,N_15130);
or U15216 (N_15216,N_15001,N_15147);
xor U15217 (N_15217,N_15076,N_15011);
nand U15218 (N_15218,N_15135,N_15123);
xnor U15219 (N_15219,N_15110,N_15020);
and U15220 (N_15220,N_15083,N_15044);
nand U15221 (N_15221,N_15108,N_15166);
xnor U15222 (N_15222,N_15057,N_15087);
nor U15223 (N_15223,N_15089,N_15189);
xor U15224 (N_15224,N_15071,N_15037);
nand U15225 (N_15225,N_15004,N_15190);
nor U15226 (N_15226,N_15053,N_15181);
nand U15227 (N_15227,N_15050,N_15149);
xor U15228 (N_15228,N_15081,N_15099);
or U15229 (N_15229,N_15178,N_15159);
or U15230 (N_15230,N_15010,N_15041);
nor U15231 (N_15231,N_15093,N_15128);
nand U15232 (N_15232,N_15151,N_15084);
xor U15233 (N_15233,N_15196,N_15117);
xnor U15234 (N_15234,N_15034,N_15145);
xor U15235 (N_15235,N_15163,N_15046);
nor U15236 (N_15236,N_15143,N_15186);
or U15237 (N_15237,N_15058,N_15000);
or U15238 (N_15238,N_15126,N_15155);
and U15239 (N_15239,N_15065,N_15003);
and U15240 (N_15240,N_15184,N_15152);
xor U15241 (N_15241,N_15106,N_15140);
or U15242 (N_15242,N_15175,N_15109);
nor U15243 (N_15243,N_15022,N_15015);
nand U15244 (N_15244,N_15124,N_15176);
and U15245 (N_15245,N_15170,N_15021);
and U15246 (N_15246,N_15002,N_15198);
xor U15247 (N_15247,N_15054,N_15171);
nand U15248 (N_15248,N_15146,N_15191);
and U15249 (N_15249,N_15136,N_15059);
or U15250 (N_15250,N_15160,N_15067);
xnor U15251 (N_15251,N_15051,N_15162);
or U15252 (N_15252,N_15137,N_15072);
nand U15253 (N_15253,N_15009,N_15193);
or U15254 (N_15254,N_15086,N_15088);
nor U15255 (N_15255,N_15014,N_15097);
nand U15256 (N_15256,N_15027,N_15156);
nand U15257 (N_15257,N_15066,N_15069);
and U15258 (N_15258,N_15134,N_15174);
nor U15259 (N_15259,N_15079,N_15129);
nor U15260 (N_15260,N_15132,N_15007);
nand U15261 (N_15261,N_15029,N_15094);
nand U15262 (N_15262,N_15052,N_15024);
xor U15263 (N_15263,N_15103,N_15118);
and U15264 (N_15264,N_15187,N_15180);
xor U15265 (N_15265,N_15114,N_15092);
xnor U15266 (N_15266,N_15030,N_15197);
nor U15267 (N_15267,N_15025,N_15144);
and U15268 (N_15268,N_15199,N_15070);
xor U15269 (N_15269,N_15138,N_15040);
or U15270 (N_15270,N_15016,N_15091);
and U15271 (N_15271,N_15085,N_15150);
nand U15272 (N_15272,N_15194,N_15121);
nand U15273 (N_15273,N_15033,N_15195);
nor U15274 (N_15274,N_15064,N_15090);
and U15275 (N_15275,N_15161,N_15115);
and U15276 (N_15276,N_15158,N_15133);
and U15277 (N_15277,N_15023,N_15031);
xor U15278 (N_15278,N_15167,N_15111);
nand U15279 (N_15279,N_15157,N_15125);
xnor U15280 (N_15280,N_15168,N_15179);
xnor U15281 (N_15281,N_15142,N_15169);
xnor U15282 (N_15282,N_15102,N_15073);
or U15283 (N_15283,N_15005,N_15078);
nand U15284 (N_15284,N_15077,N_15008);
or U15285 (N_15285,N_15039,N_15105);
nor U15286 (N_15286,N_15153,N_15045);
nand U15287 (N_15287,N_15049,N_15182);
or U15288 (N_15288,N_15112,N_15101);
xnor U15289 (N_15289,N_15035,N_15032);
xnor U15290 (N_15290,N_15017,N_15148);
xnor U15291 (N_15291,N_15131,N_15116);
xor U15292 (N_15292,N_15006,N_15122);
or U15293 (N_15293,N_15080,N_15082);
and U15294 (N_15294,N_15012,N_15048);
and U15295 (N_15295,N_15120,N_15183);
nand U15296 (N_15296,N_15075,N_15098);
xnor U15297 (N_15297,N_15013,N_15177);
nor U15298 (N_15298,N_15055,N_15043);
or U15299 (N_15299,N_15068,N_15113);
and U15300 (N_15300,N_15000,N_15134);
nor U15301 (N_15301,N_15142,N_15097);
nor U15302 (N_15302,N_15171,N_15002);
or U15303 (N_15303,N_15100,N_15150);
nand U15304 (N_15304,N_15080,N_15128);
and U15305 (N_15305,N_15102,N_15041);
xor U15306 (N_15306,N_15045,N_15055);
and U15307 (N_15307,N_15023,N_15130);
nor U15308 (N_15308,N_15089,N_15011);
or U15309 (N_15309,N_15072,N_15186);
nor U15310 (N_15310,N_15120,N_15131);
xor U15311 (N_15311,N_15097,N_15046);
or U15312 (N_15312,N_15163,N_15079);
and U15313 (N_15313,N_15193,N_15134);
or U15314 (N_15314,N_15006,N_15042);
nand U15315 (N_15315,N_15010,N_15081);
and U15316 (N_15316,N_15163,N_15027);
xor U15317 (N_15317,N_15093,N_15050);
or U15318 (N_15318,N_15113,N_15146);
or U15319 (N_15319,N_15101,N_15159);
or U15320 (N_15320,N_15130,N_15022);
xor U15321 (N_15321,N_15090,N_15093);
xor U15322 (N_15322,N_15105,N_15044);
or U15323 (N_15323,N_15122,N_15024);
nor U15324 (N_15324,N_15070,N_15041);
nand U15325 (N_15325,N_15019,N_15008);
and U15326 (N_15326,N_15092,N_15165);
xor U15327 (N_15327,N_15161,N_15186);
nor U15328 (N_15328,N_15037,N_15148);
nor U15329 (N_15329,N_15079,N_15111);
xor U15330 (N_15330,N_15047,N_15183);
nand U15331 (N_15331,N_15004,N_15142);
nand U15332 (N_15332,N_15135,N_15097);
nand U15333 (N_15333,N_15161,N_15039);
and U15334 (N_15334,N_15162,N_15025);
or U15335 (N_15335,N_15015,N_15068);
nor U15336 (N_15336,N_15045,N_15137);
or U15337 (N_15337,N_15069,N_15195);
nor U15338 (N_15338,N_15143,N_15013);
or U15339 (N_15339,N_15142,N_15181);
nor U15340 (N_15340,N_15128,N_15133);
xnor U15341 (N_15341,N_15046,N_15146);
xor U15342 (N_15342,N_15072,N_15177);
or U15343 (N_15343,N_15176,N_15095);
xnor U15344 (N_15344,N_15189,N_15099);
nor U15345 (N_15345,N_15072,N_15123);
or U15346 (N_15346,N_15016,N_15136);
and U15347 (N_15347,N_15089,N_15017);
nor U15348 (N_15348,N_15111,N_15164);
xnor U15349 (N_15349,N_15155,N_15121);
nand U15350 (N_15350,N_15194,N_15005);
xnor U15351 (N_15351,N_15161,N_15130);
xnor U15352 (N_15352,N_15107,N_15117);
or U15353 (N_15353,N_15166,N_15160);
and U15354 (N_15354,N_15002,N_15084);
and U15355 (N_15355,N_15140,N_15008);
and U15356 (N_15356,N_15095,N_15034);
or U15357 (N_15357,N_15104,N_15024);
nor U15358 (N_15358,N_15057,N_15124);
or U15359 (N_15359,N_15047,N_15142);
nand U15360 (N_15360,N_15106,N_15156);
nand U15361 (N_15361,N_15129,N_15057);
xor U15362 (N_15362,N_15025,N_15111);
or U15363 (N_15363,N_15159,N_15036);
or U15364 (N_15364,N_15151,N_15194);
xor U15365 (N_15365,N_15042,N_15070);
nor U15366 (N_15366,N_15037,N_15109);
xor U15367 (N_15367,N_15198,N_15062);
and U15368 (N_15368,N_15000,N_15051);
or U15369 (N_15369,N_15066,N_15170);
nand U15370 (N_15370,N_15145,N_15008);
nor U15371 (N_15371,N_15019,N_15108);
nand U15372 (N_15372,N_15090,N_15177);
or U15373 (N_15373,N_15066,N_15161);
nand U15374 (N_15374,N_15016,N_15119);
nand U15375 (N_15375,N_15166,N_15149);
and U15376 (N_15376,N_15100,N_15079);
xor U15377 (N_15377,N_15151,N_15175);
or U15378 (N_15378,N_15177,N_15125);
or U15379 (N_15379,N_15074,N_15145);
or U15380 (N_15380,N_15185,N_15141);
or U15381 (N_15381,N_15047,N_15021);
or U15382 (N_15382,N_15175,N_15147);
or U15383 (N_15383,N_15190,N_15199);
xnor U15384 (N_15384,N_15130,N_15025);
nor U15385 (N_15385,N_15081,N_15014);
and U15386 (N_15386,N_15038,N_15125);
nor U15387 (N_15387,N_15082,N_15041);
and U15388 (N_15388,N_15088,N_15175);
nor U15389 (N_15389,N_15128,N_15075);
or U15390 (N_15390,N_15061,N_15164);
xor U15391 (N_15391,N_15069,N_15196);
nor U15392 (N_15392,N_15166,N_15196);
and U15393 (N_15393,N_15100,N_15174);
xnor U15394 (N_15394,N_15021,N_15056);
nand U15395 (N_15395,N_15005,N_15022);
nand U15396 (N_15396,N_15035,N_15004);
and U15397 (N_15397,N_15172,N_15110);
xnor U15398 (N_15398,N_15161,N_15157);
or U15399 (N_15399,N_15191,N_15120);
xor U15400 (N_15400,N_15369,N_15372);
xor U15401 (N_15401,N_15321,N_15301);
and U15402 (N_15402,N_15213,N_15240);
or U15403 (N_15403,N_15352,N_15297);
xnor U15404 (N_15404,N_15245,N_15223);
or U15405 (N_15405,N_15329,N_15258);
xor U15406 (N_15406,N_15296,N_15309);
nor U15407 (N_15407,N_15212,N_15356);
nor U15408 (N_15408,N_15232,N_15376);
nor U15409 (N_15409,N_15339,N_15330);
nand U15410 (N_15410,N_15322,N_15397);
nor U15411 (N_15411,N_15226,N_15365);
nor U15412 (N_15412,N_15327,N_15255);
or U15413 (N_15413,N_15277,N_15314);
nor U15414 (N_15414,N_15293,N_15295);
nor U15415 (N_15415,N_15391,N_15249);
xor U15416 (N_15416,N_15209,N_15334);
or U15417 (N_15417,N_15253,N_15379);
nor U15418 (N_15418,N_15236,N_15267);
nor U15419 (N_15419,N_15351,N_15264);
xnor U15420 (N_15420,N_15370,N_15384);
and U15421 (N_15421,N_15299,N_15202);
and U15422 (N_15422,N_15211,N_15333);
or U15423 (N_15423,N_15221,N_15392);
and U15424 (N_15424,N_15325,N_15323);
or U15425 (N_15425,N_15399,N_15373);
or U15426 (N_15426,N_15252,N_15305);
nand U15427 (N_15427,N_15225,N_15335);
xnor U15428 (N_15428,N_15341,N_15260);
nand U15429 (N_15429,N_15316,N_15265);
or U15430 (N_15430,N_15272,N_15389);
nor U15431 (N_15431,N_15347,N_15227);
nor U15432 (N_15432,N_15308,N_15300);
nor U15433 (N_15433,N_15210,N_15248);
xor U15434 (N_15434,N_15378,N_15233);
xor U15435 (N_15435,N_15381,N_15320);
or U15436 (N_15436,N_15224,N_15288);
nor U15437 (N_15437,N_15286,N_15336);
and U15438 (N_15438,N_15219,N_15387);
xor U15439 (N_15439,N_15241,N_15244);
and U15440 (N_15440,N_15268,N_15310);
nor U15441 (N_15441,N_15386,N_15349);
and U15442 (N_15442,N_15313,N_15396);
nor U15443 (N_15443,N_15340,N_15229);
nand U15444 (N_15444,N_15385,N_15200);
nor U15445 (N_15445,N_15216,N_15243);
and U15446 (N_15446,N_15254,N_15266);
or U15447 (N_15447,N_15292,N_15263);
nand U15448 (N_15448,N_15382,N_15283);
or U15449 (N_15449,N_15375,N_15319);
and U15450 (N_15450,N_15353,N_15261);
nand U15451 (N_15451,N_15218,N_15357);
xor U15452 (N_15452,N_15355,N_15311);
nor U15453 (N_15453,N_15332,N_15383);
nand U15454 (N_15454,N_15360,N_15328);
xnor U15455 (N_15455,N_15291,N_15280);
and U15456 (N_15456,N_15228,N_15324);
and U15457 (N_15457,N_15303,N_15207);
xor U15458 (N_15458,N_15269,N_15388);
or U15459 (N_15459,N_15251,N_15214);
and U15460 (N_15460,N_15281,N_15206);
and U15461 (N_15461,N_15354,N_15398);
and U15462 (N_15462,N_15304,N_15274);
or U15463 (N_15463,N_15393,N_15395);
xnor U15464 (N_15464,N_15284,N_15390);
and U15465 (N_15465,N_15362,N_15394);
xor U15466 (N_15466,N_15279,N_15235);
and U15467 (N_15467,N_15306,N_15239);
or U15468 (N_15468,N_15256,N_15363);
and U15469 (N_15469,N_15312,N_15282);
and U15470 (N_15470,N_15290,N_15262);
nor U15471 (N_15471,N_15337,N_15271);
and U15472 (N_15472,N_15342,N_15231);
nor U15473 (N_15473,N_15204,N_15222);
nand U15474 (N_15474,N_15298,N_15230);
and U15475 (N_15475,N_15366,N_15270);
or U15476 (N_15476,N_15276,N_15318);
and U15477 (N_15477,N_15343,N_15237);
nor U15478 (N_15478,N_15201,N_15361);
nand U15479 (N_15479,N_15257,N_15377);
or U15480 (N_15480,N_15326,N_15246);
and U15481 (N_15481,N_15203,N_15250);
nand U15482 (N_15482,N_15315,N_15220);
nand U15483 (N_15483,N_15208,N_15215);
and U15484 (N_15484,N_15238,N_15338);
and U15485 (N_15485,N_15217,N_15350);
nor U15486 (N_15486,N_15302,N_15359);
and U15487 (N_15487,N_15287,N_15234);
nand U15488 (N_15488,N_15380,N_15364);
nand U15489 (N_15489,N_15294,N_15273);
nand U15490 (N_15490,N_15307,N_15278);
nor U15491 (N_15491,N_15317,N_15285);
nor U15492 (N_15492,N_15345,N_15346);
xnor U15493 (N_15493,N_15331,N_15374);
or U15494 (N_15494,N_15289,N_15371);
or U15495 (N_15495,N_15368,N_15242);
and U15496 (N_15496,N_15275,N_15205);
nand U15497 (N_15497,N_15348,N_15344);
nor U15498 (N_15498,N_15358,N_15259);
nand U15499 (N_15499,N_15247,N_15367);
or U15500 (N_15500,N_15395,N_15251);
xor U15501 (N_15501,N_15243,N_15296);
nand U15502 (N_15502,N_15264,N_15253);
or U15503 (N_15503,N_15397,N_15339);
and U15504 (N_15504,N_15336,N_15387);
xor U15505 (N_15505,N_15384,N_15302);
nand U15506 (N_15506,N_15264,N_15349);
xnor U15507 (N_15507,N_15371,N_15380);
and U15508 (N_15508,N_15330,N_15201);
nand U15509 (N_15509,N_15235,N_15394);
or U15510 (N_15510,N_15381,N_15207);
or U15511 (N_15511,N_15381,N_15353);
xor U15512 (N_15512,N_15347,N_15348);
nor U15513 (N_15513,N_15216,N_15380);
nand U15514 (N_15514,N_15381,N_15214);
nor U15515 (N_15515,N_15253,N_15227);
or U15516 (N_15516,N_15205,N_15242);
nor U15517 (N_15517,N_15305,N_15271);
nor U15518 (N_15518,N_15217,N_15346);
and U15519 (N_15519,N_15318,N_15320);
nor U15520 (N_15520,N_15274,N_15251);
xnor U15521 (N_15521,N_15220,N_15336);
xor U15522 (N_15522,N_15296,N_15236);
xor U15523 (N_15523,N_15299,N_15258);
and U15524 (N_15524,N_15305,N_15361);
nand U15525 (N_15525,N_15346,N_15321);
xnor U15526 (N_15526,N_15213,N_15351);
or U15527 (N_15527,N_15208,N_15338);
and U15528 (N_15528,N_15353,N_15252);
and U15529 (N_15529,N_15202,N_15364);
and U15530 (N_15530,N_15333,N_15232);
nand U15531 (N_15531,N_15359,N_15333);
xnor U15532 (N_15532,N_15279,N_15302);
nor U15533 (N_15533,N_15345,N_15235);
and U15534 (N_15534,N_15391,N_15357);
or U15535 (N_15535,N_15303,N_15241);
xnor U15536 (N_15536,N_15353,N_15331);
and U15537 (N_15537,N_15378,N_15225);
xor U15538 (N_15538,N_15320,N_15292);
nor U15539 (N_15539,N_15261,N_15340);
nand U15540 (N_15540,N_15390,N_15251);
nand U15541 (N_15541,N_15295,N_15254);
or U15542 (N_15542,N_15326,N_15324);
xor U15543 (N_15543,N_15274,N_15242);
nor U15544 (N_15544,N_15332,N_15273);
nand U15545 (N_15545,N_15312,N_15386);
or U15546 (N_15546,N_15222,N_15339);
xor U15547 (N_15547,N_15384,N_15304);
xor U15548 (N_15548,N_15349,N_15368);
nor U15549 (N_15549,N_15224,N_15366);
nand U15550 (N_15550,N_15310,N_15315);
and U15551 (N_15551,N_15227,N_15274);
nand U15552 (N_15552,N_15264,N_15266);
nand U15553 (N_15553,N_15272,N_15240);
nand U15554 (N_15554,N_15205,N_15326);
and U15555 (N_15555,N_15280,N_15296);
and U15556 (N_15556,N_15245,N_15371);
xor U15557 (N_15557,N_15363,N_15340);
and U15558 (N_15558,N_15347,N_15321);
and U15559 (N_15559,N_15321,N_15341);
and U15560 (N_15560,N_15250,N_15298);
nand U15561 (N_15561,N_15385,N_15220);
xnor U15562 (N_15562,N_15236,N_15358);
and U15563 (N_15563,N_15211,N_15234);
or U15564 (N_15564,N_15291,N_15211);
nor U15565 (N_15565,N_15264,N_15353);
nor U15566 (N_15566,N_15221,N_15314);
or U15567 (N_15567,N_15353,N_15277);
nor U15568 (N_15568,N_15261,N_15222);
nand U15569 (N_15569,N_15310,N_15316);
and U15570 (N_15570,N_15262,N_15343);
nand U15571 (N_15571,N_15314,N_15363);
xor U15572 (N_15572,N_15353,N_15260);
or U15573 (N_15573,N_15262,N_15353);
xnor U15574 (N_15574,N_15241,N_15320);
xor U15575 (N_15575,N_15288,N_15343);
xor U15576 (N_15576,N_15213,N_15383);
or U15577 (N_15577,N_15331,N_15310);
and U15578 (N_15578,N_15358,N_15253);
or U15579 (N_15579,N_15392,N_15368);
and U15580 (N_15580,N_15214,N_15240);
or U15581 (N_15581,N_15358,N_15381);
and U15582 (N_15582,N_15389,N_15321);
or U15583 (N_15583,N_15332,N_15364);
or U15584 (N_15584,N_15281,N_15299);
and U15585 (N_15585,N_15369,N_15264);
or U15586 (N_15586,N_15346,N_15328);
and U15587 (N_15587,N_15276,N_15358);
nand U15588 (N_15588,N_15340,N_15323);
nand U15589 (N_15589,N_15282,N_15343);
nand U15590 (N_15590,N_15289,N_15252);
and U15591 (N_15591,N_15242,N_15295);
or U15592 (N_15592,N_15342,N_15328);
xor U15593 (N_15593,N_15338,N_15282);
xor U15594 (N_15594,N_15267,N_15351);
and U15595 (N_15595,N_15293,N_15205);
and U15596 (N_15596,N_15279,N_15310);
and U15597 (N_15597,N_15304,N_15393);
nand U15598 (N_15598,N_15301,N_15222);
xnor U15599 (N_15599,N_15291,N_15250);
nor U15600 (N_15600,N_15515,N_15548);
xor U15601 (N_15601,N_15406,N_15468);
or U15602 (N_15602,N_15440,N_15504);
nor U15603 (N_15603,N_15453,N_15461);
or U15604 (N_15604,N_15452,N_15567);
nand U15605 (N_15605,N_15525,N_15427);
or U15606 (N_15606,N_15500,N_15550);
nor U15607 (N_15607,N_15517,N_15539);
or U15608 (N_15608,N_15422,N_15435);
or U15609 (N_15609,N_15491,N_15527);
xor U15610 (N_15610,N_15535,N_15488);
nor U15611 (N_15611,N_15547,N_15594);
and U15612 (N_15612,N_15465,N_15580);
and U15613 (N_15613,N_15596,N_15450);
nor U15614 (N_15614,N_15416,N_15560);
and U15615 (N_15615,N_15519,N_15474);
and U15616 (N_15616,N_15446,N_15480);
and U15617 (N_15617,N_15593,N_15469);
nor U15618 (N_15618,N_15569,N_15551);
xnor U15619 (N_15619,N_15419,N_15423);
nor U15620 (N_15620,N_15499,N_15520);
or U15621 (N_15621,N_15415,N_15505);
xnor U15622 (N_15622,N_15591,N_15512);
or U15623 (N_15623,N_15451,N_15431);
nand U15624 (N_15624,N_15534,N_15510);
or U15625 (N_15625,N_15475,N_15570);
nor U15626 (N_15626,N_15555,N_15574);
nand U15627 (N_15627,N_15564,N_15442);
nand U15628 (N_15628,N_15434,N_15439);
and U15629 (N_15629,N_15577,N_15585);
and U15630 (N_15630,N_15409,N_15497);
nand U15631 (N_15631,N_15443,N_15565);
and U15632 (N_15632,N_15455,N_15546);
nor U15633 (N_15633,N_15587,N_15522);
xnor U15634 (N_15634,N_15552,N_15405);
nand U15635 (N_15635,N_15496,N_15595);
and U15636 (N_15636,N_15597,N_15572);
and U15637 (N_15637,N_15473,N_15432);
nor U15638 (N_15638,N_15449,N_15454);
nand U15639 (N_15639,N_15470,N_15411);
xor U15640 (N_15640,N_15575,N_15403);
nand U15641 (N_15641,N_15563,N_15457);
nand U15642 (N_15642,N_15589,N_15479);
xnor U15643 (N_15643,N_15420,N_15521);
and U15644 (N_15644,N_15489,N_15506);
and U15645 (N_15645,N_15476,N_15400);
and U15646 (N_15646,N_15471,N_15509);
nor U15647 (N_15647,N_15428,N_15583);
or U15648 (N_15648,N_15456,N_15484);
nor U15649 (N_15649,N_15542,N_15503);
nand U15650 (N_15650,N_15472,N_15573);
nor U15651 (N_15651,N_15516,N_15407);
nand U15652 (N_15652,N_15507,N_15414);
nand U15653 (N_15653,N_15561,N_15498);
xnor U15654 (N_15654,N_15424,N_15538);
xnor U15655 (N_15655,N_15557,N_15501);
nand U15656 (N_15656,N_15448,N_15586);
or U15657 (N_15657,N_15438,N_15523);
and U15658 (N_15658,N_15466,N_15578);
and U15659 (N_15659,N_15486,N_15447);
nand U15660 (N_15660,N_15531,N_15410);
nand U15661 (N_15661,N_15502,N_15459);
xor U15662 (N_15662,N_15462,N_15558);
nor U15663 (N_15663,N_15529,N_15599);
nor U15664 (N_15664,N_15544,N_15566);
or U15665 (N_15665,N_15463,N_15549);
and U15666 (N_15666,N_15437,N_15545);
nand U15667 (N_15667,N_15537,N_15518);
nand U15668 (N_15668,N_15576,N_15458);
nand U15669 (N_15669,N_15408,N_15444);
nand U15670 (N_15670,N_15426,N_15553);
xor U15671 (N_15671,N_15532,N_15483);
or U15672 (N_15672,N_15592,N_15579);
nand U15673 (N_15673,N_15464,N_15588);
xor U15674 (N_15674,N_15495,N_15477);
xnor U15675 (N_15675,N_15430,N_15485);
xnor U15676 (N_15676,N_15524,N_15540);
xnor U15677 (N_15677,N_15493,N_15559);
xor U15678 (N_15678,N_15413,N_15433);
or U15679 (N_15679,N_15460,N_15436);
nor U15680 (N_15680,N_15481,N_15429);
nand U15681 (N_15681,N_15417,N_15494);
nor U15682 (N_15682,N_15590,N_15402);
nor U15683 (N_15683,N_15582,N_15445);
nand U15684 (N_15684,N_15554,N_15543);
xor U15685 (N_15685,N_15571,N_15418);
or U15686 (N_15686,N_15404,N_15401);
nand U15687 (N_15687,N_15556,N_15528);
xor U15688 (N_15688,N_15530,N_15482);
xor U15689 (N_15689,N_15598,N_15412);
and U15690 (N_15690,N_15533,N_15513);
nand U15691 (N_15691,N_15584,N_15511);
and U15692 (N_15692,N_15425,N_15478);
or U15693 (N_15693,N_15568,N_15581);
xor U15694 (N_15694,N_15467,N_15487);
and U15695 (N_15695,N_15541,N_15441);
and U15696 (N_15696,N_15526,N_15490);
xnor U15697 (N_15697,N_15508,N_15492);
xnor U15698 (N_15698,N_15562,N_15421);
or U15699 (N_15699,N_15514,N_15536);
nor U15700 (N_15700,N_15527,N_15405);
xor U15701 (N_15701,N_15517,N_15593);
nand U15702 (N_15702,N_15557,N_15516);
nor U15703 (N_15703,N_15490,N_15586);
nand U15704 (N_15704,N_15402,N_15535);
xnor U15705 (N_15705,N_15418,N_15432);
nor U15706 (N_15706,N_15514,N_15435);
nor U15707 (N_15707,N_15552,N_15528);
or U15708 (N_15708,N_15448,N_15479);
nand U15709 (N_15709,N_15517,N_15556);
xnor U15710 (N_15710,N_15565,N_15584);
nand U15711 (N_15711,N_15547,N_15548);
nand U15712 (N_15712,N_15447,N_15572);
or U15713 (N_15713,N_15451,N_15475);
nand U15714 (N_15714,N_15469,N_15411);
nor U15715 (N_15715,N_15553,N_15531);
nor U15716 (N_15716,N_15453,N_15444);
and U15717 (N_15717,N_15524,N_15599);
and U15718 (N_15718,N_15405,N_15426);
nand U15719 (N_15719,N_15533,N_15570);
nand U15720 (N_15720,N_15402,N_15536);
nor U15721 (N_15721,N_15553,N_15561);
nor U15722 (N_15722,N_15414,N_15432);
or U15723 (N_15723,N_15521,N_15598);
nor U15724 (N_15724,N_15492,N_15593);
xnor U15725 (N_15725,N_15456,N_15414);
nand U15726 (N_15726,N_15509,N_15408);
nand U15727 (N_15727,N_15561,N_15487);
nor U15728 (N_15728,N_15450,N_15505);
xnor U15729 (N_15729,N_15473,N_15448);
and U15730 (N_15730,N_15535,N_15482);
nor U15731 (N_15731,N_15500,N_15456);
nor U15732 (N_15732,N_15545,N_15528);
or U15733 (N_15733,N_15411,N_15523);
nand U15734 (N_15734,N_15465,N_15515);
or U15735 (N_15735,N_15480,N_15421);
nand U15736 (N_15736,N_15560,N_15408);
nand U15737 (N_15737,N_15556,N_15571);
nand U15738 (N_15738,N_15550,N_15425);
nor U15739 (N_15739,N_15491,N_15457);
or U15740 (N_15740,N_15511,N_15596);
xor U15741 (N_15741,N_15500,N_15507);
or U15742 (N_15742,N_15579,N_15489);
or U15743 (N_15743,N_15521,N_15422);
or U15744 (N_15744,N_15568,N_15590);
nor U15745 (N_15745,N_15455,N_15562);
nand U15746 (N_15746,N_15568,N_15551);
or U15747 (N_15747,N_15507,N_15525);
xnor U15748 (N_15748,N_15493,N_15573);
nand U15749 (N_15749,N_15540,N_15419);
nor U15750 (N_15750,N_15560,N_15465);
or U15751 (N_15751,N_15503,N_15516);
or U15752 (N_15752,N_15503,N_15410);
xnor U15753 (N_15753,N_15404,N_15499);
nand U15754 (N_15754,N_15559,N_15553);
and U15755 (N_15755,N_15540,N_15577);
xor U15756 (N_15756,N_15432,N_15531);
and U15757 (N_15757,N_15538,N_15446);
nor U15758 (N_15758,N_15592,N_15553);
and U15759 (N_15759,N_15566,N_15477);
nor U15760 (N_15760,N_15422,N_15497);
or U15761 (N_15761,N_15579,N_15433);
nor U15762 (N_15762,N_15520,N_15495);
and U15763 (N_15763,N_15550,N_15431);
and U15764 (N_15764,N_15515,N_15574);
or U15765 (N_15765,N_15537,N_15502);
xor U15766 (N_15766,N_15565,N_15506);
xor U15767 (N_15767,N_15565,N_15454);
xnor U15768 (N_15768,N_15506,N_15406);
nor U15769 (N_15769,N_15549,N_15422);
nand U15770 (N_15770,N_15522,N_15589);
xnor U15771 (N_15771,N_15540,N_15475);
nand U15772 (N_15772,N_15436,N_15470);
or U15773 (N_15773,N_15514,N_15448);
xor U15774 (N_15774,N_15465,N_15556);
nand U15775 (N_15775,N_15446,N_15524);
xnor U15776 (N_15776,N_15548,N_15428);
nor U15777 (N_15777,N_15536,N_15471);
nor U15778 (N_15778,N_15465,N_15431);
xnor U15779 (N_15779,N_15499,N_15531);
nor U15780 (N_15780,N_15477,N_15409);
xnor U15781 (N_15781,N_15587,N_15569);
nor U15782 (N_15782,N_15532,N_15577);
xor U15783 (N_15783,N_15492,N_15554);
nand U15784 (N_15784,N_15589,N_15533);
xnor U15785 (N_15785,N_15551,N_15440);
nand U15786 (N_15786,N_15545,N_15483);
or U15787 (N_15787,N_15521,N_15573);
xnor U15788 (N_15788,N_15559,N_15573);
and U15789 (N_15789,N_15469,N_15518);
xor U15790 (N_15790,N_15592,N_15433);
and U15791 (N_15791,N_15494,N_15461);
nor U15792 (N_15792,N_15493,N_15472);
nand U15793 (N_15793,N_15519,N_15478);
nand U15794 (N_15794,N_15524,N_15405);
or U15795 (N_15795,N_15534,N_15486);
nor U15796 (N_15796,N_15494,N_15489);
and U15797 (N_15797,N_15547,N_15419);
xor U15798 (N_15798,N_15497,N_15402);
or U15799 (N_15799,N_15549,N_15521);
xnor U15800 (N_15800,N_15683,N_15646);
or U15801 (N_15801,N_15752,N_15745);
xnor U15802 (N_15802,N_15761,N_15739);
and U15803 (N_15803,N_15712,N_15648);
and U15804 (N_15804,N_15630,N_15792);
xnor U15805 (N_15805,N_15795,N_15654);
or U15806 (N_15806,N_15604,N_15643);
xnor U15807 (N_15807,N_15605,N_15673);
nor U15808 (N_15808,N_15627,N_15798);
nor U15809 (N_15809,N_15772,N_15771);
or U15810 (N_15810,N_15600,N_15621);
and U15811 (N_15811,N_15642,N_15791);
nand U15812 (N_15812,N_15733,N_15715);
xnor U15813 (N_15813,N_15665,N_15725);
xor U15814 (N_15814,N_15703,N_15625);
xor U15815 (N_15815,N_15607,N_15731);
or U15816 (N_15816,N_15777,N_15714);
nand U15817 (N_15817,N_15697,N_15672);
xor U15818 (N_15818,N_15664,N_15743);
nand U15819 (N_15819,N_15732,N_15649);
xor U15820 (N_15820,N_15754,N_15736);
nand U15821 (N_15821,N_15787,N_15685);
nand U15822 (N_15822,N_15602,N_15684);
nand U15823 (N_15823,N_15629,N_15723);
or U15824 (N_15824,N_15615,N_15652);
nor U15825 (N_15825,N_15738,N_15681);
or U15826 (N_15826,N_15679,N_15663);
xnor U15827 (N_15827,N_15770,N_15666);
xor U15828 (N_15828,N_15786,N_15693);
xor U15829 (N_15829,N_15616,N_15634);
nor U15830 (N_15830,N_15617,N_15780);
or U15831 (N_15831,N_15656,N_15775);
nor U15832 (N_15832,N_15718,N_15701);
or U15833 (N_15833,N_15620,N_15794);
nand U15834 (N_15834,N_15692,N_15610);
xnor U15835 (N_15835,N_15707,N_15719);
xor U15836 (N_15836,N_15769,N_15660);
nor U15837 (N_15837,N_15614,N_15698);
xor U15838 (N_15838,N_15713,N_15609);
nand U15839 (N_15839,N_15789,N_15678);
and U15840 (N_15840,N_15662,N_15767);
nand U15841 (N_15841,N_15696,N_15647);
nor U15842 (N_15842,N_15766,N_15682);
xor U15843 (N_15843,N_15776,N_15690);
or U15844 (N_15844,N_15758,N_15782);
nand U15845 (N_15845,N_15717,N_15751);
or U15846 (N_15846,N_15760,N_15637);
nand U15847 (N_15847,N_15608,N_15705);
nor U15848 (N_15848,N_15710,N_15757);
or U15849 (N_15849,N_15730,N_15675);
nand U15850 (N_15850,N_15603,N_15623);
nor U15851 (N_15851,N_15756,N_15774);
or U15852 (N_15852,N_15626,N_15727);
nand U15853 (N_15853,N_15635,N_15742);
xor U15854 (N_15854,N_15677,N_15721);
and U15855 (N_15855,N_15778,N_15686);
nand U15856 (N_15856,N_15773,N_15618);
xor U15857 (N_15857,N_15764,N_15781);
and U15858 (N_15858,N_15688,N_15657);
or U15859 (N_15859,N_15613,N_15601);
nor U15860 (N_15860,N_15729,N_15612);
xor U15861 (N_15861,N_15793,N_15711);
or U15862 (N_15862,N_15728,N_15628);
or U15863 (N_15863,N_15785,N_15645);
and U15864 (N_15864,N_15661,N_15633);
or U15865 (N_15865,N_15768,N_15651);
or U15866 (N_15866,N_15783,N_15748);
xor U15867 (N_15867,N_15640,N_15708);
or U15868 (N_15868,N_15765,N_15691);
nand U15869 (N_15869,N_15716,N_15650);
nor U15870 (N_15870,N_15779,N_15655);
or U15871 (N_15871,N_15644,N_15636);
nor U15872 (N_15872,N_15659,N_15671);
or U15873 (N_15873,N_15709,N_15741);
nand U15874 (N_15874,N_15668,N_15759);
or U15875 (N_15875,N_15670,N_15796);
nor U15876 (N_15876,N_15658,N_15747);
nand U15877 (N_15877,N_15797,N_15611);
xnor U15878 (N_15878,N_15750,N_15746);
nor U15879 (N_15879,N_15619,N_15734);
nand U15880 (N_15880,N_15622,N_15694);
and U15881 (N_15881,N_15689,N_15638);
and U15882 (N_15882,N_15744,N_15702);
and U15883 (N_15883,N_15749,N_15755);
and U15884 (N_15884,N_15722,N_15706);
and U15885 (N_15885,N_15680,N_15720);
or U15886 (N_15886,N_15790,N_15740);
and U15887 (N_15887,N_15737,N_15669);
nand U15888 (N_15888,N_15788,N_15726);
nand U15889 (N_15889,N_15641,N_15624);
or U15890 (N_15890,N_15687,N_15763);
and U15891 (N_15891,N_15632,N_15784);
xnor U15892 (N_15892,N_15695,N_15639);
nand U15893 (N_15893,N_15724,N_15699);
nor U15894 (N_15894,N_15753,N_15667);
nand U15895 (N_15895,N_15762,N_15676);
nand U15896 (N_15896,N_15704,N_15700);
xnor U15897 (N_15897,N_15653,N_15631);
xor U15898 (N_15898,N_15799,N_15674);
xnor U15899 (N_15899,N_15735,N_15606);
or U15900 (N_15900,N_15726,N_15763);
and U15901 (N_15901,N_15671,N_15643);
xnor U15902 (N_15902,N_15644,N_15623);
xor U15903 (N_15903,N_15702,N_15773);
and U15904 (N_15904,N_15738,N_15752);
and U15905 (N_15905,N_15751,N_15744);
or U15906 (N_15906,N_15719,N_15720);
and U15907 (N_15907,N_15690,N_15696);
or U15908 (N_15908,N_15763,N_15622);
xnor U15909 (N_15909,N_15682,N_15613);
xor U15910 (N_15910,N_15637,N_15627);
or U15911 (N_15911,N_15659,N_15636);
nor U15912 (N_15912,N_15661,N_15646);
and U15913 (N_15913,N_15737,N_15636);
xor U15914 (N_15914,N_15751,N_15608);
or U15915 (N_15915,N_15769,N_15775);
or U15916 (N_15916,N_15689,N_15656);
nor U15917 (N_15917,N_15760,N_15754);
nand U15918 (N_15918,N_15601,N_15605);
and U15919 (N_15919,N_15747,N_15772);
nand U15920 (N_15920,N_15635,N_15676);
and U15921 (N_15921,N_15648,N_15779);
or U15922 (N_15922,N_15612,N_15677);
and U15923 (N_15923,N_15694,N_15704);
nor U15924 (N_15924,N_15790,N_15650);
nand U15925 (N_15925,N_15709,N_15711);
nor U15926 (N_15926,N_15655,N_15689);
xnor U15927 (N_15927,N_15759,N_15654);
or U15928 (N_15928,N_15622,N_15601);
nand U15929 (N_15929,N_15600,N_15791);
nor U15930 (N_15930,N_15740,N_15779);
and U15931 (N_15931,N_15680,N_15736);
nand U15932 (N_15932,N_15656,N_15749);
and U15933 (N_15933,N_15605,N_15799);
nor U15934 (N_15934,N_15643,N_15758);
xnor U15935 (N_15935,N_15770,N_15748);
xor U15936 (N_15936,N_15659,N_15623);
xor U15937 (N_15937,N_15666,N_15775);
xnor U15938 (N_15938,N_15779,N_15716);
nand U15939 (N_15939,N_15601,N_15686);
nor U15940 (N_15940,N_15693,N_15689);
nor U15941 (N_15941,N_15687,N_15764);
nand U15942 (N_15942,N_15702,N_15627);
xor U15943 (N_15943,N_15653,N_15742);
and U15944 (N_15944,N_15770,N_15772);
nand U15945 (N_15945,N_15779,N_15726);
and U15946 (N_15946,N_15788,N_15642);
or U15947 (N_15947,N_15666,N_15655);
nand U15948 (N_15948,N_15658,N_15762);
or U15949 (N_15949,N_15658,N_15608);
or U15950 (N_15950,N_15717,N_15668);
nor U15951 (N_15951,N_15738,N_15723);
nand U15952 (N_15952,N_15771,N_15611);
nand U15953 (N_15953,N_15735,N_15618);
xnor U15954 (N_15954,N_15734,N_15637);
xnor U15955 (N_15955,N_15635,N_15625);
nor U15956 (N_15956,N_15603,N_15650);
xnor U15957 (N_15957,N_15783,N_15651);
nand U15958 (N_15958,N_15623,N_15756);
nand U15959 (N_15959,N_15746,N_15769);
nor U15960 (N_15960,N_15741,N_15653);
and U15961 (N_15961,N_15710,N_15612);
nand U15962 (N_15962,N_15611,N_15607);
nand U15963 (N_15963,N_15698,N_15669);
nor U15964 (N_15964,N_15696,N_15758);
and U15965 (N_15965,N_15784,N_15792);
xnor U15966 (N_15966,N_15670,N_15794);
nand U15967 (N_15967,N_15624,N_15623);
nor U15968 (N_15968,N_15703,N_15678);
xnor U15969 (N_15969,N_15606,N_15638);
nand U15970 (N_15970,N_15659,N_15645);
nand U15971 (N_15971,N_15798,N_15692);
xor U15972 (N_15972,N_15764,N_15645);
xnor U15973 (N_15973,N_15650,N_15737);
and U15974 (N_15974,N_15757,N_15727);
nand U15975 (N_15975,N_15706,N_15787);
or U15976 (N_15976,N_15646,N_15696);
or U15977 (N_15977,N_15748,N_15667);
nand U15978 (N_15978,N_15693,N_15730);
nor U15979 (N_15979,N_15660,N_15765);
xnor U15980 (N_15980,N_15788,N_15693);
and U15981 (N_15981,N_15615,N_15780);
xor U15982 (N_15982,N_15779,N_15766);
or U15983 (N_15983,N_15660,N_15608);
or U15984 (N_15984,N_15610,N_15770);
and U15985 (N_15985,N_15659,N_15667);
xor U15986 (N_15986,N_15735,N_15727);
nand U15987 (N_15987,N_15615,N_15698);
nand U15988 (N_15988,N_15740,N_15781);
xnor U15989 (N_15989,N_15779,N_15614);
xor U15990 (N_15990,N_15648,N_15705);
and U15991 (N_15991,N_15706,N_15684);
nor U15992 (N_15992,N_15631,N_15645);
or U15993 (N_15993,N_15727,N_15765);
nor U15994 (N_15994,N_15685,N_15719);
nor U15995 (N_15995,N_15767,N_15670);
xnor U15996 (N_15996,N_15675,N_15610);
or U15997 (N_15997,N_15714,N_15778);
or U15998 (N_15998,N_15795,N_15613);
or U15999 (N_15999,N_15649,N_15655);
nor U16000 (N_16000,N_15884,N_15960);
and U16001 (N_16001,N_15907,N_15868);
and U16002 (N_16002,N_15895,N_15961);
nand U16003 (N_16003,N_15919,N_15874);
nor U16004 (N_16004,N_15940,N_15914);
or U16005 (N_16005,N_15927,N_15891);
or U16006 (N_16006,N_15879,N_15885);
or U16007 (N_16007,N_15970,N_15854);
nand U16008 (N_16008,N_15807,N_15815);
nand U16009 (N_16009,N_15838,N_15865);
xor U16010 (N_16010,N_15930,N_15812);
nor U16011 (N_16011,N_15902,N_15996);
xor U16012 (N_16012,N_15915,N_15999);
nor U16013 (N_16013,N_15908,N_15934);
and U16014 (N_16014,N_15889,N_15988);
nand U16015 (N_16015,N_15836,N_15993);
xnor U16016 (N_16016,N_15949,N_15849);
xor U16017 (N_16017,N_15989,N_15911);
nor U16018 (N_16018,N_15892,N_15916);
and U16019 (N_16019,N_15931,N_15984);
nor U16020 (N_16020,N_15852,N_15969);
nor U16021 (N_16021,N_15851,N_15867);
or U16022 (N_16022,N_15894,N_15944);
xor U16023 (N_16023,N_15841,N_15901);
xnor U16024 (N_16024,N_15802,N_15906);
nand U16025 (N_16025,N_15821,N_15848);
nand U16026 (N_16026,N_15805,N_15942);
nand U16027 (N_16027,N_15832,N_15847);
xnor U16028 (N_16028,N_15987,N_15939);
xnor U16029 (N_16029,N_15972,N_15962);
nor U16030 (N_16030,N_15910,N_15973);
xor U16031 (N_16031,N_15816,N_15982);
nor U16032 (N_16032,N_15955,N_15880);
xnor U16033 (N_16033,N_15951,N_15866);
and U16034 (N_16034,N_15829,N_15935);
nor U16035 (N_16035,N_15921,N_15978);
xnor U16036 (N_16036,N_15819,N_15967);
or U16037 (N_16037,N_15971,N_15976);
and U16038 (N_16038,N_15823,N_15888);
xnor U16039 (N_16039,N_15997,N_15990);
nor U16040 (N_16040,N_15881,N_15833);
nor U16041 (N_16041,N_15947,N_15963);
and U16042 (N_16042,N_15995,N_15922);
or U16043 (N_16043,N_15898,N_15992);
or U16044 (N_16044,N_15820,N_15965);
xnor U16045 (N_16045,N_15900,N_15909);
nand U16046 (N_16046,N_15905,N_15862);
xnor U16047 (N_16047,N_15818,N_15856);
nand U16048 (N_16048,N_15861,N_15804);
nand U16049 (N_16049,N_15958,N_15946);
nand U16050 (N_16050,N_15873,N_15893);
nor U16051 (N_16051,N_15814,N_15913);
nor U16052 (N_16052,N_15860,N_15869);
or U16053 (N_16053,N_15839,N_15857);
or U16054 (N_16054,N_15903,N_15932);
and U16055 (N_16055,N_15923,N_15986);
nor U16056 (N_16056,N_15887,N_15878);
xor U16057 (N_16057,N_15801,N_15974);
or U16058 (N_16058,N_15863,N_15834);
nor U16059 (N_16059,N_15813,N_15803);
or U16060 (N_16060,N_15825,N_15844);
nor U16061 (N_16061,N_15808,N_15864);
nand U16062 (N_16062,N_15985,N_15850);
nor U16063 (N_16063,N_15966,N_15979);
or U16064 (N_16064,N_15870,N_15918);
and U16065 (N_16065,N_15830,N_15842);
or U16066 (N_16066,N_15883,N_15877);
xor U16067 (N_16067,N_15991,N_15924);
nor U16068 (N_16068,N_15875,N_15837);
and U16069 (N_16069,N_15933,N_15952);
and U16070 (N_16070,N_15840,N_15994);
or U16071 (N_16071,N_15920,N_15959);
and U16072 (N_16072,N_15811,N_15956);
nor U16073 (N_16073,N_15843,N_15938);
xnor U16074 (N_16074,N_15859,N_15846);
xnor U16075 (N_16075,N_15981,N_15928);
nand U16076 (N_16076,N_15822,N_15904);
nand U16077 (N_16077,N_15817,N_15827);
nand U16078 (N_16078,N_15897,N_15983);
nand U16079 (N_16079,N_15926,N_15809);
nand U16080 (N_16080,N_15925,N_15871);
and U16081 (N_16081,N_15890,N_15948);
and U16082 (N_16082,N_15917,N_15929);
or U16083 (N_16083,N_15824,N_15826);
or U16084 (N_16084,N_15977,N_15858);
nor U16085 (N_16085,N_15975,N_15937);
nand U16086 (N_16086,N_15828,N_15800);
or U16087 (N_16087,N_15950,N_15957);
or U16088 (N_16088,N_15941,N_15980);
nor U16089 (N_16089,N_15896,N_15943);
or U16090 (N_16090,N_15945,N_15845);
nand U16091 (N_16091,N_15806,N_15954);
xor U16092 (N_16092,N_15835,N_15998);
and U16093 (N_16093,N_15953,N_15882);
nor U16094 (N_16094,N_15810,N_15886);
and U16095 (N_16095,N_15853,N_15872);
xnor U16096 (N_16096,N_15876,N_15912);
nand U16097 (N_16097,N_15855,N_15831);
xnor U16098 (N_16098,N_15968,N_15899);
and U16099 (N_16099,N_15936,N_15964);
xor U16100 (N_16100,N_15998,N_15981);
xor U16101 (N_16101,N_15911,N_15817);
or U16102 (N_16102,N_15957,N_15866);
nor U16103 (N_16103,N_15923,N_15858);
nor U16104 (N_16104,N_15827,N_15959);
nand U16105 (N_16105,N_15971,N_15946);
and U16106 (N_16106,N_15877,N_15892);
xnor U16107 (N_16107,N_15978,N_15953);
and U16108 (N_16108,N_15879,N_15905);
and U16109 (N_16109,N_15924,N_15844);
nand U16110 (N_16110,N_15837,N_15914);
nand U16111 (N_16111,N_15983,N_15988);
nor U16112 (N_16112,N_15920,N_15843);
nor U16113 (N_16113,N_15803,N_15983);
or U16114 (N_16114,N_15920,N_15859);
nand U16115 (N_16115,N_15846,N_15994);
xor U16116 (N_16116,N_15944,N_15818);
or U16117 (N_16117,N_15861,N_15932);
and U16118 (N_16118,N_15871,N_15998);
xnor U16119 (N_16119,N_15834,N_15821);
nor U16120 (N_16120,N_15809,N_15919);
and U16121 (N_16121,N_15908,N_15807);
nand U16122 (N_16122,N_15953,N_15844);
or U16123 (N_16123,N_15874,N_15974);
xnor U16124 (N_16124,N_15885,N_15875);
nor U16125 (N_16125,N_15852,N_15828);
xor U16126 (N_16126,N_15958,N_15819);
nand U16127 (N_16127,N_15987,N_15875);
nor U16128 (N_16128,N_15915,N_15972);
nand U16129 (N_16129,N_15869,N_15837);
and U16130 (N_16130,N_15986,N_15914);
nor U16131 (N_16131,N_15882,N_15809);
and U16132 (N_16132,N_15943,N_15879);
nor U16133 (N_16133,N_15878,N_15879);
or U16134 (N_16134,N_15804,N_15867);
nor U16135 (N_16135,N_15915,N_15826);
or U16136 (N_16136,N_15839,N_15884);
and U16137 (N_16137,N_15852,N_15987);
xnor U16138 (N_16138,N_15940,N_15934);
or U16139 (N_16139,N_15806,N_15906);
and U16140 (N_16140,N_15811,N_15836);
or U16141 (N_16141,N_15860,N_15933);
or U16142 (N_16142,N_15886,N_15924);
or U16143 (N_16143,N_15910,N_15840);
nor U16144 (N_16144,N_15860,N_15991);
or U16145 (N_16145,N_15996,N_15812);
nand U16146 (N_16146,N_15918,N_15977);
and U16147 (N_16147,N_15821,N_15932);
nand U16148 (N_16148,N_15958,N_15913);
nand U16149 (N_16149,N_15807,N_15834);
or U16150 (N_16150,N_15979,N_15969);
and U16151 (N_16151,N_15910,N_15819);
nor U16152 (N_16152,N_15991,N_15925);
and U16153 (N_16153,N_15976,N_15887);
or U16154 (N_16154,N_15897,N_15849);
and U16155 (N_16155,N_15993,N_15992);
xor U16156 (N_16156,N_15957,N_15825);
xor U16157 (N_16157,N_15817,N_15978);
and U16158 (N_16158,N_15913,N_15851);
nand U16159 (N_16159,N_15821,N_15859);
or U16160 (N_16160,N_15916,N_15962);
or U16161 (N_16161,N_15805,N_15928);
nand U16162 (N_16162,N_15903,N_15823);
nand U16163 (N_16163,N_15956,N_15953);
nor U16164 (N_16164,N_15909,N_15853);
xor U16165 (N_16165,N_15968,N_15989);
and U16166 (N_16166,N_15980,N_15872);
or U16167 (N_16167,N_15987,N_15878);
nor U16168 (N_16168,N_15895,N_15904);
nor U16169 (N_16169,N_15851,N_15968);
xnor U16170 (N_16170,N_15967,N_15834);
or U16171 (N_16171,N_15841,N_15825);
or U16172 (N_16172,N_15938,N_15873);
nand U16173 (N_16173,N_15907,N_15875);
xor U16174 (N_16174,N_15929,N_15977);
and U16175 (N_16175,N_15911,N_15864);
xnor U16176 (N_16176,N_15801,N_15996);
xnor U16177 (N_16177,N_15812,N_15880);
xnor U16178 (N_16178,N_15856,N_15893);
nor U16179 (N_16179,N_15961,N_15931);
nor U16180 (N_16180,N_15973,N_15962);
nor U16181 (N_16181,N_15918,N_15999);
xnor U16182 (N_16182,N_15911,N_15918);
nand U16183 (N_16183,N_15874,N_15923);
xnor U16184 (N_16184,N_15817,N_15967);
and U16185 (N_16185,N_15801,N_15982);
nor U16186 (N_16186,N_15834,N_15861);
xor U16187 (N_16187,N_15995,N_15911);
nand U16188 (N_16188,N_15830,N_15857);
xnor U16189 (N_16189,N_15815,N_15927);
or U16190 (N_16190,N_15958,N_15820);
or U16191 (N_16191,N_15896,N_15912);
and U16192 (N_16192,N_15851,N_15919);
xor U16193 (N_16193,N_15858,N_15872);
and U16194 (N_16194,N_15909,N_15865);
xor U16195 (N_16195,N_15950,N_15850);
or U16196 (N_16196,N_15919,N_15993);
nor U16197 (N_16197,N_15902,N_15954);
nor U16198 (N_16198,N_15874,N_15854);
nand U16199 (N_16199,N_15925,N_15873);
xor U16200 (N_16200,N_16156,N_16157);
nor U16201 (N_16201,N_16183,N_16180);
nand U16202 (N_16202,N_16012,N_16016);
and U16203 (N_16203,N_16017,N_16165);
xor U16204 (N_16204,N_16075,N_16029);
nand U16205 (N_16205,N_16086,N_16138);
nand U16206 (N_16206,N_16044,N_16167);
nand U16207 (N_16207,N_16110,N_16142);
or U16208 (N_16208,N_16126,N_16105);
and U16209 (N_16209,N_16198,N_16137);
nor U16210 (N_16210,N_16127,N_16027);
nand U16211 (N_16211,N_16085,N_16149);
nand U16212 (N_16212,N_16010,N_16061);
and U16213 (N_16213,N_16195,N_16095);
xnor U16214 (N_16214,N_16119,N_16045);
nor U16215 (N_16215,N_16152,N_16070);
nor U16216 (N_16216,N_16186,N_16094);
and U16217 (N_16217,N_16108,N_16199);
and U16218 (N_16218,N_16125,N_16065);
or U16219 (N_16219,N_16058,N_16161);
nand U16220 (N_16220,N_16054,N_16043);
nand U16221 (N_16221,N_16109,N_16158);
xnor U16222 (N_16222,N_16041,N_16118);
nor U16223 (N_16223,N_16196,N_16068);
or U16224 (N_16224,N_16064,N_16123);
nand U16225 (N_16225,N_16194,N_16100);
xnor U16226 (N_16226,N_16114,N_16013);
or U16227 (N_16227,N_16188,N_16038);
nor U16228 (N_16228,N_16000,N_16185);
or U16229 (N_16229,N_16116,N_16021);
or U16230 (N_16230,N_16088,N_16117);
nand U16231 (N_16231,N_16024,N_16059);
nand U16232 (N_16232,N_16187,N_16122);
nand U16233 (N_16233,N_16023,N_16092);
or U16234 (N_16234,N_16164,N_16020);
nor U16235 (N_16235,N_16083,N_16028);
and U16236 (N_16236,N_16177,N_16015);
or U16237 (N_16237,N_16079,N_16022);
xor U16238 (N_16238,N_16145,N_16004);
xor U16239 (N_16239,N_16066,N_16076);
and U16240 (N_16240,N_16090,N_16036);
nand U16241 (N_16241,N_16169,N_16046);
or U16242 (N_16242,N_16166,N_16097);
and U16243 (N_16243,N_16101,N_16160);
or U16244 (N_16244,N_16153,N_16001);
and U16245 (N_16245,N_16143,N_16191);
and U16246 (N_16246,N_16121,N_16175);
and U16247 (N_16247,N_16031,N_16019);
nor U16248 (N_16248,N_16128,N_16071);
xor U16249 (N_16249,N_16089,N_16112);
nand U16250 (N_16250,N_16179,N_16174);
or U16251 (N_16251,N_16002,N_16129);
nor U16252 (N_16252,N_16163,N_16077);
nand U16253 (N_16253,N_16104,N_16181);
and U16254 (N_16254,N_16113,N_16078);
nor U16255 (N_16255,N_16155,N_16147);
or U16256 (N_16256,N_16193,N_16154);
or U16257 (N_16257,N_16053,N_16096);
nor U16258 (N_16258,N_16184,N_16074);
nor U16259 (N_16259,N_16069,N_16067);
and U16260 (N_16260,N_16190,N_16107);
xor U16261 (N_16261,N_16171,N_16146);
and U16262 (N_16262,N_16037,N_16047);
nor U16263 (N_16263,N_16150,N_16176);
nand U16264 (N_16264,N_16140,N_16049);
or U16265 (N_16265,N_16035,N_16081);
nand U16266 (N_16266,N_16093,N_16072);
or U16267 (N_16267,N_16111,N_16162);
nor U16268 (N_16268,N_16131,N_16073);
nor U16269 (N_16269,N_16011,N_16120);
or U16270 (N_16270,N_16141,N_16087);
nor U16271 (N_16271,N_16007,N_16026);
or U16272 (N_16272,N_16062,N_16008);
nand U16273 (N_16273,N_16042,N_16052);
nor U16274 (N_16274,N_16197,N_16148);
nor U16275 (N_16275,N_16056,N_16080);
nor U16276 (N_16276,N_16178,N_16084);
nor U16277 (N_16277,N_16103,N_16151);
and U16278 (N_16278,N_16034,N_16136);
nand U16279 (N_16279,N_16102,N_16014);
nor U16280 (N_16280,N_16005,N_16135);
nand U16281 (N_16281,N_16051,N_16057);
nor U16282 (N_16282,N_16050,N_16033);
nor U16283 (N_16283,N_16003,N_16099);
nor U16284 (N_16284,N_16130,N_16025);
and U16285 (N_16285,N_16055,N_16032);
xnor U16286 (N_16286,N_16132,N_16063);
nand U16287 (N_16287,N_16091,N_16168);
and U16288 (N_16288,N_16134,N_16139);
nor U16289 (N_16289,N_16006,N_16040);
or U16290 (N_16290,N_16039,N_16009);
nand U16291 (N_16291,N_16048,N_16133);
nor U16292 (N_16292,N_16170,N_16144);
and U16293 (N_16293,N_16060,N_16030);
nand U16294 (N_16294,N_16192,N_16124);
and U16295 (N_16295,N_16172,N_16115);
and U16296 (N_16296,N_16082,N_16018);
nor U16297 (N_16297,N_16159,N_16098);
and U16298 (N_16298,N_16106,N_16189);
nand U16299 (N_16299,N_16182,N_16173);
and U16300 (N_16300,N_16088,N_16150);
xor U16301 (N_16301,N_16111,N_16046);
nand U16302 (N_16302,N_16041,N_16119);
nor U16303 (N_16303,N_16107,N_16041);
and U16304 (N_16304,N_16148,N_16140);
nand U16305 (N_16305,N_16104,N_16171);
or U16306 (N_16306,N_16092,N_16122);
or U16307 (N_16307,N_16037,N_16126);
or U16308 (N_16308,N_16003,N_16076);
xnor U16309 (N_16309,N_16103,N_16002);
and U16310 (N_16310,N_16056,N_16104);
nand U16311 (N_16311,N_16110,N_16195);
or U16312 (N_16312,N_16086,N_16063);
and U16313 (N_16313,N_16106,N_16040);
xnor U16314 (N_16314,N_16057,N_16066);
xnor U16315 (N_16315,N_16166,N_16179);
xnor U16316 (N_16316,N_16114,N_16009);
or U16317 (N_16317,N_16195,N_16128);
xor U16318 (N_16318,N_16151,N_16121);
nand U16319 (N_16319,N_16013,N_16058);
or U16320 (N_16320,N_16164,N_16147);
or U16321 (N_16321,N_16045,N_16164);
nand U16322 (N_16322,N_16178,N_16161);
nor U16323 (N_16323,N_16095,N_16016);
xor U16324 (N_16324,N_16011,N_16129);
nor U16325 (N_16325,N_16114,N_16074);
or U16326 (N_16326,N_16097,N_16010);
or U16327 (N_16327,N_16020,N_16050);
and U16328 (N_16328,N_16009,N_16067);
nand U16329 (N_16329,N_16058,N_16059);
and U16330 (N_16330,N_16075,N_16199);
and U16331 (N_16331,N_16082,N_16076);
nor U16332 (N_16332,N_16108,N_16126);
nand U16333 (N_16333,N_16096,N_16124);
xnor U16334 (N_16334,N_16142,N_16067);
and U16335 (N_16335,N_16087,N_16075);
or U16336 (N_16336,N_16196,N_16059);
nor U16337 (N_16337,N_16067,N_16170);
or U16338 (N_16338,N_16167,N_16142);
or U16339 (N_16339,N_16179,N_16051);
or U16340 (N_16340,N_16077,N_16000);
and U16341 (N_16341,N_16175,N_16188);
nand U16342 (N_16342,N_16021,N_16041);
nand U16343 (N_16343,N_16105,N_16100);
nor U16344 (N_16344,N_16001,N_16197);
xor U16345 (N_16345,N_16002,N_16066);
nor U16346 (N_16346,N_16112,N_16077);
and U16347 (N_16347,N_16046,N_16135);
xor U16348 (N_16348,N_16145,N_16085);
and U16349 (N_16349,N_16040,N_16026);
nor U16350 (N_16350,N_16053,N_16009);
nor U16351 (N_16351,N_16078,N_16049);
and U16352 (N_16352,N_16192,N_16076);
nand U16353 (N_16353,N_16060,N_16154);
xnor U16354 (N_16354,N_16191,N_16007);
or U16355 (N_16355,N_16070,N_16095);
and U16356 (N_16356,N_16003,N_16187);
and U16357 (N_16357,N_16045,N_16189);
or U16358 (N_16358,N_16129,N_16198);
xor U16359 (N_16359,N_16061,N_16096);
nand U16360 (N_16360,N_16170,N_16106);
and U16361 (N_16361,N_16197,N_16150);
or U16362 (N_16362,N_16050,N_16026);
or U16363 (N_16363,N_16114,N_16085);
nand U16364 (N_16364,N_16041,N_16059);
nor U16365 (N_16365,N_16074,N_16164);
xnor U16366 (N_16366,N_16071,N_16143);
or U16367 (N_16367,N_16181,N_16080);
nand U16368 (N_16368,N_16038,N_16044);
and U16369 (N_16369,N_16112,N_16140);
and U16370 (N_16370,N_16036,N_16116);
and U16371 (N_16371,N_16142,N_16047);
nand U16372 (N_16372,N_16096,N_16071);
nand U16373 (N_16373,N_16169,N_16041);
and U16374 (N_16374,N_16053,N_16177);
or U16375 (N_16375,N_16025,N_16198);
nor U16376 (N_16376,N_16178,N_16127);
xnor U16377 (N_16377,N_16151,N_16140);
xor U16378 (N_16378,N_16060,N_16085);
or U16379 (N_16379,N_16169,N_16045);
or U16380 (N_16380,N_16125,N_16035);
nor U16381 (N_16381,N_16057,N_16129);
nor U16382 (N_16382,N_16024,N_16168);
nor U16383 (N_16383,N_16127,N_16089);
xnor U16384 (N_16384,N_16006,N_16071);
or U16385 (N_16385,N_16016,N_16003);
or U16386 (N_16386,N_16098,N_16168);
or U16387 (N_16387,N_16105,N_16079);
xnor U16388 (N_16388,N_16044,N_16026);
nor U16389 (N_16389,N_16013,N_16003);
nand U16390 (N_16390,N_16140,N_16163);
and U16391 (N_16391,N_16165,N_16195);
nor U16392 (N_16392,N_16139,N_16089);
xnor U16393 (N_16393,N_16176,N_16172);
or U16394 (N_16394,N_16137,N_16072);
or U16395 (N_16395,N_16082,N_16074);
nand U16396 (N_16396,N_16050,N_16101);
xor U16397 (N_16397,N_16176,N_16164);
xnor U16398 (N_16398,N_16059,N_16066);
or U16399 (N_16399,N_16012,N_16175);
and U16400 (N_16400,N_16237,N_16245);
nand U16401 (N_16401,N_16262,N_16282);
or U16402 (N_16402,N_16345,N_16387);
or U16403 (N_16403,N_16312,N_16353);
nand U16404 (N_16404,N_16214,N_16221);
or U16405 (N_16405,N_16362,N_16390);
nor U16406 (N_16406,N_16256,N_16205);
xor U16407 (N_16407,N_16244,N_16233);
nor U16408 (N_16408,N_16218,N_16377);
xnor U16409 (N_16409,N_16324,N_16286);
and U16410 (N_16410,N_16287,N_16276);
nor U16411 (N_16411,N_16326,N_16241);
and U16412 (N_16412,N_16348,N_16242);
and U16413 (N_16413,N_16372,N_16229);
nor U16414 (N_16414,N_16289,N_16341);
xnor U16415 (N_16415,N_16263,N_16391);
or U16416 (N_16416,N_16291,N_16250);
xnor U16417 (N_16417,N_16223,N_16269);
nor U16418 (N_16418,N_16302,N_16264);
nand U16419 (N_16419,N_16319,N_16292);
or U16420 (N_16420,N_16265,N_16358);
nand U16421 (N_16421,N_16212,N_16274);
xnor U16422 (N_16422,N_16398,N_16337);
nand U16423 (N_16423,N_16318,N_16379);
or U16424 (N_16424,N_16283,N_16365);
and U16425 (N_16425,N_16222,N_16267);
nor U16426 (N_16426,N_16230,N_16378);
or U16427 (N_16427,N_16369,N_16299);
nor U16428 (N_16428,N_16311,N_16327);
nor U16429 (N_16429,N_16331,N_16220);
nor U16430 (N_16430,N_16397,N_16272);
or U16431 (N_16431,N_16297,N_16309);
nor U16432 (N_16432,N_16330,N_16320);
or U16433 (N_16433,N_16239,N_16367);
or U16434 (N_16434,N_16322,N_16259);
or U16435 (N_16435,N_16342,N_16228);
nand U16436 (N_16436,N_16364,N_16316);
nor U16437 (N_16437,N_16258,N_16217);
nand U16438 (N_16438,N_16293,N_16207);
xnor U16439 (N_16439,N_16211,N_16254);
nor U16440 (N_16440,N_16248,N_16317);
or U16441 (N_16441,N_16224,N_16209);
nand U16442 (N_16442,N_16251,N_16306);
and U16443 (N_16443,N_16252,N_16357);
xnor U16444 (N_16444,N_16304,N_16352);
nand U16445 (N_16445,N_16366,N_16334);
nor U16446 (N_16446,N_16346,N_16376);
xnor U16447 (N_16447,N_16392,N_16200);
xor U16448 (N_16448,N_16396,N_16307);
nor U16449 (N_16449,N_16310,N_16355);
and U16450 (N_16450,N_16275,N_16384);
and U16451 (N_16451,N_16314,N_16278);
or U16452 (N_16452,N_16270,N_16359);
and U16453 (N_16453,N_16273,N_16255);
or U16454 (N_16454,N_16399,N_16271);
xor U16455 (N_16455,N_16285,N_16395);
xnor U16456 (N_16456,N_16380,N_16338);
nor U16457 (N_16457,N_16281,N_16288);
xor U16458 (N_16458,N_16333,N_16371);
or U16459 (N_16459,N_16204,N_16243);
or U16460 (N_16460,N_16235,N_16201);
nand U16461 (N_16461,N_16386,N_16370);
nand U16462 (N_16462,N_16329,N_16210);
nand U16463 (N_16463,N_16361,N_16298);
nor U16464 (N_16464,N_16360,N_16368);
nor U16465 (N_16465,N_16385,N_16350);
and U16466 (N_16466,N_16279,N_16234);
nand U16467 (N_16467,N_16226,N_16305);
nor U16468 (N_16468,N_16240,N_16354);
nor U16469 (N_16469,N_16344,N_16303);
or U16470 (N_16470,N_16315,N_16206);
nor U16471 (N_16471,N_16332,N_16257);
or U16472 (N_16472,N_16202,N_16284);
or U16473 (N_16473,N_16343,N_16280);
nand U16474 (N_16474,N_16295,N_16389);
and U16475 (N_16475,N_16231,N_16216);
nand U16476 (N_16476,N_16247,N_16260);
nor U16477 (N_16477,N_16266,N_16300);
xor U16478 (N_16478,N_16325,N_16394);
xor U16479 (N_16479,N_16383,N_16328);
and U16480 (N_16480,N_16294,N_16340);
or U16481 (N_16481,N_16208,N_16308);
nor U16482 (N_16482,N_16336,N_16374);
nor U16483 (N_16483,N_16236,N_16375);
nand U16484 (N_16484,N_16261,N_16382);
nor U16485 (N_16485,N_16335,N_16249);
nand U16486 (N_16486,N_16277,N_16232);
nor U16487 (N_16487,N_16356,N_16393);
nor U16488 (N_16488,N_16225,N_16349);
nor U16489 (N_16489,N_16363,N_16213);
xor U16490 (N_16490,N_16301,N_16351);
xnor U16491 (N_16491,N_16381,N_16203);
and U16492 (N_16492,N_16268,N_16253);
xnor U16493 (N_16493,N_16347,N_16246);
nor U16494 (N_16494,N_16373,N_16339);
nor U16495 (N_16495,N_16290,N_16323);
nand U16496 (N_16496,N_16238,N_16227);
nand U16497 (N_16497,N_16388,N_16219);
xnor U16498 (N_16498,N_16313,N_16296);
nor U16499 (N_16499,N_16215,N_16321);
xor U16500 (N_16500,N_16351,N_16288);
and U16501 (N_16501,N_16259,N_16300);
and U16502 (N_16502,N_16253,N_16323);
or U16503 (N_16503,N_16379,N_16220);
nor U16504 (N_16504,N_16245,N_16358);
nor U16505 (N_16505,N_16351,N_16218);
nor U16506 (N_16506,N_16305,N_16340);
or U16507 (N_16507,N_16258,N_16243);
and U16508 (N_16508,N_16353,N_16280);
xor U16509 (N_16509,N_16211,N_16273);
xnor U16510 (N_16510,N_16305,N_16235);
and U16511 (N_16511,N_16275,N_16262);
xnor U16512 (N_16512,N_16391,N_16213);
nor U16513 (N_16513,N_16209,N_16344);
xor U16514 (N_16514,N_16382,N_16317);
xnor U16515 (N_16515,N_16231,N_16380);
or U16516 (N_16516,N_16393,N_16276);
nor U16517 (N_16517,N_16349,N_16215);
nand U16518 (N_16518,N_16285,N_16242);
or U16519 (N_16519,N_16227,N_16342);
and U16520 (N_16520,N_16241,N_16267);
nor U16521 (N_16521,N_16304,N_16322);
nand U16522 (N_16522,N_16331,N_16356);
nor U16523 (N_16523,N_16289,N_16366);
nor U16524 (N_16524,N_16345,N_16272);
and U16525 (N_16525,N_16268,N_16355);
nand U16526 (N_16526,N_16384,N_16379);
or U16527 (N_16527,N_16334,N_16252);
or U16528 (N_16528,N_16378,N_16307);
xnor U16529 (N_16529,N_16375,N_16208);
and U16530 (N_16530,N_16343,N_16368);
and U16531 (N_16531,N_16261,N_16254);
or U16532 (N_16532,N_16353,N_16378);
nor U16533 (N_16533,N_16277,N_16354);
nor U16534 (N_16534,N_16330,N_16324);
nand U16535 (N_16535,N_16296,N_16248);
and U16536 (N_16536,N_16392,N_16338);
nand U16537 (N_16537,N_16268,N_16231);
nor U16538 (N_16538,N_16349,N_16291);
nor U16539 (N_16539,N_16278,N_16301);
nor U16540 (N_16540,N_16262,N_16352);
and U16541 (N_16541,N_16285,N_16303);
nor U16542 (N_16542,N_16248,N_16363);
or U16543 (N_16543,N_16332,N_16262);
nor U16544 (N_16544,N_16291,N_16277);
nor U16545 (N_16545,N_16229,N_16289);
nand U16546 (N_16546,N_16254,N_16339);
xor U16547 (N_16547,N_16264,N_16207);
and U16548 (N_16548,N_16361,N_16244);
and U16549 (N_16549,N_16399,N_16293);
nor U16550 (N_16550,N_16219,N_16320);
xnor U16551 (N_16551,N_16291,N_16320);
and U16552 (N_16552,N_16214,N_16257);
nor U16553 (N_16553,N_16219,N_16278);
nand U16554 (N_16554,N_16334,N_16335);
nor U16555 (N_16555,N_16266,N_16263);
nand U16556 (N_16556,N_16201,N_16387);
and U16557 (N_16557,N_16389,N_16369);
and U16558 (N_16558,N_16250,N_16218);
xor U16559 (N_16559,N_16320,N_16342);
xor U16560 (N_16560,N_16344,N_16256);
and U16561 (N_16561,N_16214,N_16392);
nand U16562 (N_16562,N_16332,N_16353);
and U16563 (N_16563,N_16224,N_16376);
nor U16564 (N_16564,N_16256,N_16329);
nor U16565 (N_16565,N_16234,N_16206);
nand U16566 (N_16566,N_16200,N_16228);
or U16567 (N_16567,N_16351,N_16350);
nand U16568 (N_16568,N_16397,N_16344);
or U16569 (N_16569,N_16265,N_16272);
and U16570 (N_16570,N_16214,N_16330);
and U16571 (N_16571,N_16212,N_16315);
nor U16572 (N_16572,N_16294,N_16296);
nor U16573 (N_16573,N_16293,N_16229);
nor U16574 (N_16574,N_16399,N_16250);
nand U16575 (N_16575,N_16237,N_16370);
or U16576 (N_16576,N_16221,N_16205);
xnor U16577 (N_16577,N_16264,N_16245);
and U16578 (N_16578,N_16201,N_16212);
nor U16579 (N_16579,N_16220,N_16319);
nor U16580 (N_16580,N_16372,N_16348);
and U16581 (N_16581,N_16312,N_16369);
nand U16582 (N_16582,N_16324,N_16270);
nand U16583 (N_16583,N_16284,N_16251);
nand U16584 (N_16584,N_16287,N_16374);
and U16585 (N_16585,N_16252,N_16364);
nor U16586 (N_16586,N_16312,N_16227);
xor U16587 (N_16587,N_16301,N_16371);
xor U16588 (N_16588,N_16274,N_16318);
nor U16589 (N_16589,N_16347,N_16369);
nor U16590 (N_16590,N_16215,N_16369);
and U16591 (N_16591,N_16202,N_16321);
nand U16592 (N_16592,N_16357,N_16296);
or U16593 (N_16593,N_16393,N_16299);
and U16594 (N_16594,N_16395,N_16312);
or U16595 (N_16595,N_16349,N_16255);
xnor U16596 (N_16596,N_16253,N_16274);
or U16597 (N_16597,N_16261,N_16307);
and U16598 (N_16598,N_16206,N_16368);
nor U16599 (N_16599,N_16239,N_16204);
nand U16600 (N_16600,N_16462,N_16546);
nand U16601 (N_16601,N_16418,N_16561);
or U16602 (N_16602,N_16467,N_16559);
xnor U16603 (N_16603,N_16479,N_16461);
nand U16604 (N_16604,N_16450,N_16523);
nor U16605 (N_16605,N_16595,N_16425);
nand U16606 (N_16606,N_16496,N_16516);
or U16607 (N_16607,N_16517,N_16430);
and U16608 (N_16608,N_16481,N_16515);
or U16609 (N_16609,N_16484,N_16447);
xor U16610 (N_16610,N_16514,N_16485);
nand U16611 (N_16611,N_16531,N_16534);
xor U16612 (N_16612,N_16544,N_16573);
nand U16613 (N_16613,N_16588,N_16564);
and U16614 (N_16614,N_16477,N_16550);
or U16615 (N_16615,N_16527,N_16429);
or U16616 (N_16616,N_16555,N_16518);
nand U16617 (N_16617,N_16420,N_16431);
nand U16618 (N_16618,N_16465,N_16422);
nand U16619 (N_16619,N_16437,N_16410);
xor U16620 (N_16620,N_16511,N_16582);
xor U16621 (N_16621,N_16557,N_16469);
nand U16622 (N_16622,N_16509,N_16590);
or U16623 (N_16623,N_16442,N_16565);
and U16624 (N_16624,N_16497,N_16405);
nand U16625 (N_16625,N_16597,N_16592);
nand U16626 (N_16626,N_16417,N_16413);
nand U16627 (N_16627,N_16476,N_16554);
and U16628 (N_16628,N_16505,N_16500);
and U16629 (N_16629,N_16568,N_16545);
xor U16630 (N_16630,N_16407,N_16507);
nand U16631 (N_16631,N_16444,N_16503);
xor U16632 (N_16632,N_16501,N_16401);
or U16633 (N_16633,N_16574,N_16508);
nand U16634 (N_16634,N_16400,N_16510);
and U16635 (N_16635,N_16540,N_16406);
nor U16636 (N_16636,N_16502,N_16435);
xor U16637 (N_16637,N_16530,N_16598);
xor U16638 (N_16638,N_16486,N_16542);
xnor U16639 (N_16639,N_16553,N_16424);
nor U16640 (N_16640,N_16535,N_16490);
xor U16641 (N_16641,N_16566,N_16423);
xnor U16642 (N_16642,N_16551,N_16416);
xnor U16643 (N_16643,N_16524,N_16512);
and U16644 (N_16644,N_16529,N_16414);
and U16645 (N_16645,N_16495,N_16441);
or U16646 (N_16646,N_16464,N_16532);
nand U16647 (N_16647,N_16458,N_16528);
nand U16648 (N_16648,N_16428,N_16533);
xor U16649 (N_16649,N_16549,N_16468);
nand U16650 (N_16650,N_16599,N_16591);
xor U16651 (N_16651,N_16419,N_16572);
xnor U16652 (N_16652,N_16536,N_16473);
xor U16653 (N_16653,N_16459,N_16579);
nor U16654 (N_16654,N_16570,N_16594);
and U16655 (N_16655,N_16434,N_16576);
nand U16656 (N_16656,N_16499,N_16491);
nor U16657 (N_16657,N_16415,N_16506);
or U16658 (N_16658,N_16454,N_16583);
nand U16659 (N_16659,N_16522,N_16548);
or U16660 (N_16660,N_16436,N_16433);
and U16661 (N_16661,N_16498,N_16593);
xor U16662 (N_16662,N_16408,N_16472);
nand U16663 (N_16663,N_16480,N_16525);
nand U16664 (N_16664,N_16562,N_16448);
nor U16665 (N_16665,N_16571,N_16541);
xor U16666 (N_16666,N_16521,N_16471);
or U16667 (N_16667,N_16446,N_16402);
xor U16668 (N_16668,N_16537,N_16409);
nor U16669 (N_16669,N_16478,N_16520);
nor U16670 (N_16670,N_16552,N_16403);
and U16671 (N_16671,N_16596,N_16513);
nor U16672 (N_16672,N_16463,N_16556);
nand U16673 (N_16673,N_16451,N_16455);
and U16674 (N_16674,N_16581,N_16470);
xor U16675 (N_16675,N_16567,N_16504);
nor U16676 (N_16676,N_16587,N_16466);
or U16677 (N_16677,N_16494,N_16483);
nor U16678 (N_16678,N_16580,N_16443);
nor U16679 (N_16679,N_16489,N_16586);
and U16680 (N_16680,N_16427,N_16577);
or U16681 (N_16681,N_16456,N_16543);
nand U16682 (N_16682,N_16460,N_16411);
xor U16683 (N_16683,N_16482,N_16457);
or U16684 (N_16684,N_16538,N_16493);
and U16685 (N_16685,N_16539,N_16563);
or U16686 (N_16686,N_16475,N_16492);
or U16687 (N_16687,N_16578,N_16452);
nand U16688 (N_16688,N_16589,N_16438);
or U16689 (N_16689,N_16404,N_16474);
nand U16690 (N_16690,N_16547,N_16432);
or U16691 (N_16691,N_16575,N_16453);
nand U16692 (N_16692,N_16584,N_16569);
and U16693 (N_16693,N_16445,N_16440);
nor U16694 (N_16694,N_16560,N_16488);
nand U16695 (N_16695,N_16439,N_16519);
nor U16696 (N_16696,N_16526,N_16421);
nor U16697 (N_16697,N_16585,N_16412);
nand U16698 (N_16698,N_16487,N_16426);
or U16699 (N_16699,N_16449,N_16558);
nor U16700 (N_16700,N_16528,N_16426);
xor U16701 (N_16701,N_16560,N_16520);
and U16702 (N_16702,N_16515,N_16576);
or U16703 (N_16703,N_16550,N_16447);
and U16704 (N_16704,N_16489,N_16594);
xor U16705 (N_16705,N_16461,N_16540);
or U16706 (N_16706,N_16557,N_16457);
xnor U16707 (N_16707,N_16408,N_16502);
nor U16708 (N_16708,N_16459,N_16499);
xor U16709 (N_16709,N_16407,N_16505);
xor U16710 (N_16710,N_16568,N_16498);
and U16711 (N_16711,N_16586,N_16487);
nand U16712 (N_16712,N_16527,N_16434);
xnor U16713 (N_16713,N_16507,N_16404);
and U16714 (N_16714,N_16511,N_16406);
or U16715 (N_16715,N_16487,N_16406);
nand U16716 (N_16716,N_16525,N_16487);
or U16717 (N_16717,N_16433,N_16553);
xnor U16718 (N_16718,N_16486,N_16426);
and U16719 (N_16719,N_16473,N_16525);
xnor U16720 (N_16720,N_16410,N_16552);
nand U16721 (N_16721,N_16548,N_16563);
or U16722 (N_16722,N_16432,N_16416);
and U16723 (N_16723,N_16409,N_16421);
and U16724 (N_16724,N_16469,N_16432);
xnor U16725 (N_16725,N_16436,N_16516);
nand U16726 (N_16726,N_16470,N_16556);
xnor U16727 (N_16727,N_16501,N_16531);
xor U16728 (N_16728,N_16552,N_16556);
and U16729 (N_16729,N_16537,N_16465);
or U16730 (N_16730,N_16528,N_16440);
nor U16731 (N_16731,N_16526,N_16515);
or U16732 (N_16732,N_16555,N_16524);
xor U16733 (N_16733,N_16424,N_16591);
xnor U16734 (N_16734,N_16422,N_16455);
nor U16735 (N_16735,N_16449,N_16539);
nor U16736 (N_16736,N_16407,N_16596);
and U16737 (N_16737,N_16411,N_16571);
nor U16738 (N_16738,N_16410,N_16576);
and U16739 (N_16739,N_16534,N_16581);
or U16740 (N_16740,N_16429,N_16451);
xnor U16741 (N_16741,N_16484,N_16541);
and U16742 (N_16742,N_16469,N_16521);
nor U16743 (N_16743,N_16595,N_16405);
nand U16744 (N_16744,N_16495,N_16593);
and U16745 (N_16745,N_16439,N_16437);
nand U16746 (N_16746,N_16495,N_16413);
xnor U16747 (N_16747,N_16512,N_16406);
xnor U16748 (N_16748,N_16527,N_16407);
and U16749 (N_16749,N_16421,N_16594);
nor U16750 (N_16750,N_16511,N_16469);
nor U16751 (N_16751,N_16548,N_16447);
or U16752 (N_16752,N_16528,N_16577);
nor U16753 (N_16753,N_16486,N_16513);
or U16754 (N_16754,N_16478,N_16482);
nor U16755 (N_16755,N_16554,N_16517);
or U16756 (N_16756,N_16562,N_16543);
and U16757 (N_16757,N_16520,N_16441);
xnor U16758 (N_16758,N_16444,N_16461);
and U16759 (N_16759,N_16508,N_16434);
or U16760 (N_16760,N_16487,N_16485);
or U16761 (N_16761,N_16589,N_16484);
xor U16762 (N_16762,N_16522,N_16508);
nor U16763 (N_16763,N_16510,N_16484);
and U16764 (N_16764,N_16516,N_16486);
nand U16765 (N_16765,N_16460,N_16504);
or U16766 (N_16766,N_16421,N_16454);
and U16767 (N_16767,N_16407,N_16498);
xor U16768 (N_16768,N_16582,N_16444);
or U16769 (N_16769,N_16492,N_16544);
xor U16770 (N_16770,N_16474,N_16440);
and U16771 (N_16771,N_16480,N_16446);
or U16772 (N_16772,N_16436,N_16486);
nor U16773 (N_16773,N_16490,N_16449);
nor U16774 (N_16774,N_16438,N_16454);
nor U16775 (N_16775,N_16552,N_16569);
or U16776 (N_16776,N_16587,N_16407);
nor U16777 (N_16777,N_16557,N_16416);
nand U16778 (N_16778,N_16563,N_16460);
or U16779 (N_16779,N_16454,N_16576);
nor U16780 (N_16780,N_16427,N_16500);
nor U16781 (N_16781,N_16577,N_16564);
nor U16782 (N_16782,N_16512,N_16405);
or U16783 (N_16783,N_16588,N_16496);
nor U16784 (N_16784,N_16496,N_16533);
or U16785 (N_16785,N_16442,N_16405);
and U16786 (N_16786,N_16478,N_16402);
and U16787 (N_16787,N_16439,N_16409);
xnor U16788 (N_16788,N_16461,N_16499);
and U16789 (N_16789,N_16418,N_16476);
or U16790 (N_16790,N_16461,N_16576);
xnor U16791 (N_16791,N_16492,N_16521);
and U16792 (N_16792,N_16589,N_16598);
nor U16793 (N_16793,N_16506,N_16553);
nor U16794 (N_16794,N_16596,N_16527);
xor U16795 (N_16795,N_16438,N_16415);
and U16796 (N_16796,N_16555,N_16469);
or U16797 (N_16797,N_16437,N_16470);
nor U16798 (N_16798,N_16507,N_16589);
xnor U16799 (N_16799,N_16543,N_16591);
or U16800 (N_16800,N_16793,N_16700);
or U16801 (N_16801,N_16710,N_16771);
nor U16802 (N_16802,N_16729,N_16759);
nand U16803 (N_16803,N_16630,N_16607);
nor U16804 (N_16804,N_16666,N_16746);
nand U16805 (N_16805,N_16715,N_16637);
nand U16806 (N_16806,N_16758,N_16732);
nor U16807 (N_16807,N_16652,N_16694);
nor U16808 (N_16808,N_16662,N_16720);
xnor U16809 (N_16809,N_16726,N_16724);
nor U16810 (N_16810,N_16717,N_16788);
nor U16811 (N_16811,N_16725,N_16684);
nor U16812 (N_16812,N_16625,N_16782);
or U16813 (N_16813,N_16740,N_16698);
and U16814 (N_16814,N_16754,N_16752);
nor U16815 (N_16815,N_16691,N_16617);
nor U16816 (N_16816,N_16604,N_16649);
xor U16817 (N_16817,N_16790,N_16753);
or U16818 (N_16818,N_16727,N_16688);
xor U16819 (N_16819,N_16663,N_16682);
and U16820 (N_16820,N_16749,N_16642);
or U16821 (N_16821,N_16766,N_16600);
and U16822 (N_16822,N_16747,N_16621);
nor U16823 (N_16823,N_16693,N_16728);
xnor U16824 (N_16824,N_16786,N_16692);
nor U16825 (N_16825,N_16647,N_16792);
nand U16826 (N_16826,N_16653,N_16639);
nor U16827 (N_16827,N_16708,N_16674);
xor U16828 (N_16828,N_16703,N_16613);
or U16829 (N_16829,N_16606,N_16660);
and U16830 (N_16830,N_16722,N_16744);
and U16831 (N_16831,N_16742,N_16709);
and U16832 (N_16832,N_16608,N_16787);
and U16833 (N_16833,N_16723,N_16629);
nor U16834 (N_16834,N_16781,N_16676);
or U16835 (N_16835,N_16737,N_16735);
xnor U16836 (N_16836,N_16797,N_16713);
nand U16837 (N_16837,N_16768,N_16774);
xor U16838 (N_16838,N_16603,N_16695);
xor U16839 (N_16839,N_16702,N_16770);
or U16840 (N_16840,N_16772,N_16773);
nor U16841 (N_16841,N_16670,N_16689);
nand U16842 (N_16842,N_16760,N_16669);
or U16843 (N_16843,N_16614,N_16736);
or U16844 (N_16844,N_16636,N_16632);
xor U16845 (N_16845,N_16767,N_16743);
xnor U16846 (N_16846,N_16657,N_16779);
nor U16847 (N_16847,N_16661,N_16650);
nor U16848 (N_16848,N_16761,N_16643);
and U16849 (N_16849,N_16762,N_16648);
or U16850 (N_16850,N_16704,N_16751);
nor U16851 (N_16851,N_16678,N_16690);
and U16852 (N_16852,N_16756,N_16795);
nand U16853 (N_16853,N_16699,N_16711);
nand U16854 (N_16854,N_16644,N_16796);
nor U16855 (N_16855,N_16671,N_16610);
and U16856 (N_16856,N_16664,N_16776);
and U16857 (N_16857,N_16683,N_16654);
nand U16858 (N_16858,N_16734,N_16721);
and U16859 (N_16859,N_16741,N_16780);
nor U16860 (N_16860,N_16665,N_16623);
nor U16861 (N_16861,N_16628,N_16641);
and U16862 (N_16862,N_16611,N_16656);
xnor U16863 (N_16863,N_16798,N_16731);
xor U16864 (N_16864,N_16616,N_16745);
or U16865 (N_16865,N_16687,N_16706);
nand U16866 (N_16866,N_16799,N_16764);
or U16867 (N_16867,N_16775,N_16696);
and U16868 (N_16868,N_16645,N_16626);
xnor U16869 (N_16869,N_16701,N_16739);
nor U16870 (N_16870,N_16633,N_16622);
xnor U16871 (N_16871,N_16697,N_16755);
and U16872 (N_16872,N_16769,N_16750);
nand U16873 (N_16873,N_16627,N_16624);
nor U16874 (N_16874,N_16791,N_16615);
nand U16875 (N_16875,N_16605,N_16667);
or U16876 (N_16876,N_16763,N_16778);
xnor U16877 (N_16877,N_16785,N_16686);
nand U16878 (N_16878,N_16672,N_16719);
xor U16879 (N_16879,N_16659,N_16634);
nand U16880 (N_16880,N_16609,N_16716);
or U16881 (N_16881,N_16618,N_16612);
and U16882 (N_16882,N_16651,N_16748);
xor U16883 (N_16883,N_16640,N_16794);
xor U16884 (N_16884,N_16602,N_16619);
and U16885 (N_16885,N_16707,N_16784);
or U16886 (N_16886,N_16730,N_16685);
or U16887 (N_16887,N_16733,N_16783);
nand U16888 (N_16888,N_16668,N_16675);
and U16889 (N_16889,N_16712,N_16646);
nand U16890 (N_16890,N_16631,N_16765);
xor U16891 (N_16891,N_16705,N_16718);
nor U16892 (N_16892,N_16635,N_16757);
xor U16893 (N_16893,N_16777,N_16655);
and U16894 (N_16894,N_16677,N_16601);
and U16895 (N_16895,N_16620,N_16680);
nand U16896 (N_16896,N_16658,N_16738);
nand U16897 (N_16897,N_16681,N_16789);
and U16898 (N_16898,N_16714,N_16638);
nand U16899 (N_16899,N_16673,N_16679);
nor U16900 (N_16900,N_16766,N_16763);
and U16901 (N_16901,N_16780,N_16609);
xnor U16902 (N_16902,N_16634,N_16755);
and U16903 (N_16903,N_16631,N_16762);
xnor U16904 (N_16904,N_16681,N_16716);
nand U16905 (N_16905,N_16655,N_16771);
or U16906 (N_16906,N_16616,N_16765);
xnor U16907 (N_16907,N_16642,N_16729);
xnor U16908 (N_16908,N_16679,N_16785);
nand U16909 (N_16909,N_16773,N_16784);
or U16910 (N_16910,N_16632,N_16625);
or U16911 (N_16911,N_16736,N_16735);
and U16912 (N_16912,N_16631,N_16714);
xor U16913 (N_16913,N_16609,N_16650);
or U16914 (N_16914,N_16742,N_16693);
xor U16915 (N_16915,N_16663,N_16734);
nor U16916 (N_16916,N_16642,N_16744);
nand U16917 (N_16917,N_16714,N_16741);
or U16918 (N_16918,N_16737,N_16622);
and U16919 (N_16919,N_16738,N_16736);
or U16920 (N_16920,N_16719,N_16652);
nor U16921 (N_16921,N_16621,N_16623);
nor U16922 (N_16922,N_16637,N_16719);
or U16923 (N_16923,N_16638,N_16742);
nand U16924 (N_16924,N_16717,N_16705);
xor U16925 (N_16925,N_16724,N_16727);
nor U16926 (N_16926,N_16618,N_16765);
nor U16927 (N_16927,N_16616,N_16720);
and U16928 (N_16928,N_16687,N_16703);
nor U16929 (N_16929,N_16745,N_16655);
and U16930 (N_16930,N_16711,N_16730);
or U16931 (N_16931,N_16652,N_16763);
and U16932 (N_16932,N_16743,N_16724);
nand U16933 (N_16933,N_16711,N_16759);
or U16934 (N_16934,N_16601,N_16684);
nor U16935 (N_16935,N_16763,N_16671);
and U16936 (N_16936,N_16684,N_16749);
or U16937 (N_16937,N_16698,N_16660);
xnor U16938 (N_16938,N_16676,N_16741);
nor U16939 (N_16939,N_16660,N_16609);
xnor U16940 (N_16940,N_16727,N_16678);
nor U16941 (N_16941,N_16744,N_16665);
or U16942 (N_16942,N_16762,N_16615);
nor U16943 (N_16943,N_16707,N_16757);
xor U16944 (N_16944,N_16651,N_16684);
nor U16945 (N_16945,N_16640,N_16737);
and U16946 (N_16946,N_16708,N_16645);
and U16947 (N_16947,N_16759,N_16667);
nand U16948 (N_16948,N_16759,N_16792);
xnor U16949 (N_16949,N_16756,N_16793);
and U16950 (N_16950,N_16679,N_16681);
xnor U16951 (N_16951,N_16623,N_16792);
nor U16952 (N_16952,N_16624,N_16720);
and U16953 (N_16953,N_16697,N_16728);
and U16954 (N_16954,N_16605,N_16655);
xnor U16955 (N_16955,N_16772,N_16629);
nor U16956 (N_16956,N_16708,N_16685);
nand U16957 (N_16957,N_16611,N_16653);
xor U16958 (N_16958,N_16786,N_16623);
and U16959 (N_16959,N_16744,N_16747);
nand U16960 (N_16960,N_16756,N_16623);
and U16961 (N_16961,N_16732,N_16679);
nor U16962 (N_16962,N_16670,N_16700);
xnor U16963 (N_16963,N_16765,N_16704);
and U16964 (N_16964,N_16761,N_16601);
nand U16965 (N_16965,N_16698,N_16721);
xor U16966 (N_16966,N_16796,N_16694);
and U16967 (N_16967,N_16748,N_16763);
xor U16968 (N_16968,N_16680,N_16667);
xnor U16969 (N_16969,N_16681,N_16702);
xor U16970 (N_16970,N_16753,N_16766);
nor U16971 (N_16971,N_16751,N_16681);
nand U16972 (N_16972,N_16607,N_16793);
and U16973 (N_16973,N_16636,N_16678);
nor U16974 (N_16974,N_16719,N_16737);
nand U16975 (N_16975,N_16797,N_16717);
xnor U16976 (N_16976,N_16665,N_16754);
nor U16977 (N_16977,N_16761,N_16674);
or U16978 (N_16978,N_16697,N_16739);
and U16979 (N_16979,N_16775,N_16663);
or U16980 (N_16980,N_16705,N_16747);
xor U16981 (N_16981,N_16789,N_16772);
nand U16982 (N_16982,N_16619,N_16610);
nor U16983 (N_16983,N_16606,N_16788);
or U16984 (N_16984,N_16669,N_16699);
nand U16985 (N_16985,N_16719,N_16629);
and U16986 (N_16986,N_16665,N_16658);
xnor U16987 (N_16987,N_16692,N_16679);
xnor U16988 (N_16988,N_16619,N_16727);
and U16989 (N_16989,N_16774,N_16738);
nand U16990 (N_16990,N_16765,N_16683);
nor U16991 (N_16991,N_16635,N_16756);
or U16992 (N_16992,N_16649,N_16786);
nor U16993 (N_16993,N_16752,N_16764);
nor U16994 (N_16994,N_16680,N_16767);
nand U16995 (N_16995,N_16785,N_16623);
or U16996 (N_16996,N_16767,N_16733);
nor U16997 (N_16997,N_16749,N_16622);
nor U16998 (N_16998,N_16723,N_16681);
nor U16999 (N_16999,N_16745,N_16719);
nor U17000 (N_17000,N_16876,N_16914);
xor U17001 (N_17001,N_16854,N_16827);
or U17002 (N_17002,N_16974,N_16831);
nand U17003 (N_17003,N_16921,N_16967);
and U17004 (N_17004,N_16990,N_16904);
nand U17005 (N_17005,N_16960,N_16905);
nor U17006 (N_17006,N_16947,N_16989);
or U17007 (N_17007,N_16871,N_16861);
nor U17008 (N_17008,N_16883,N_16924);
xnor U17009 (N_17009,N_16848,N_16822);
or U17010 (N_17010,N_16935,N_16913);
xor U17011 (N_17011,N_16872,N_16801);
and U17012 (N_17012,N_16925,N_16918);
nand U17013 (N_17013,N_16936,N_16865);
or U17014 (N_17014,N_16844,N_16922);
nand U17015 (N_17015,N_16968,N_16923);
and U17016 (N_17016,N_16893,N_16847);
or U17017 (N_17017,N_16881,N_16941);
and U17018 (N_17018,N_16972,N_16991);
nor U17019 (N_17019,N_16834,N_16851);
and U17020 (N_17020,N_16829,N_16812);
nand U17021 (N_17021,N_16869,N_16944);
nor U17022 (N_17022,N_16874,N_16815);
or U17023 (N_17023,N_16832,N_16840);
and U17024 (N_17024,N_16939,N_16973);
or U17025 (N_17025,N_16868,N_16819);
nand U17026 (N_17026,N_16825,N_16997);
nor U17027 (N_17027,N_16953,N_16928);
nand U17028 (N_17028,N_16965,N_16942);
nand U17029 (N_17029,N_16969,N_16954);
nand U17030 (N_17030,N_16889,N_16917);
xnor U17031 (N_17031,N_16836,N_16945);
nand U17032 (N_17032,N_16946,N_16977);
nor U17033 (N_17033,N_16826,N_16828);
and U17034 (N_17034,N_16891,N_16966);
nor U17035 (N_17035,N_16808,N_16982);
and U17036 (N_17036,N_16919,N_16994);
and U17037 (N_17037,N_16853,N_16882);
xnor U17038 (N_17038,N_16937,N_16906);
nand U17039 (N_17039,N_16897,N_16809);
and U17040 (N_17040,N_16863,N_16860);
nor U17041 (N_17041,N_16821,N_16800);
nor U17042 (N_17042,N_16956,N_16885);
nor U17043 (N_17043,N_16938,N_16858);
nand U17044 (N_17044,N_16817,N_16943);
or U17045 (N_17045,N_16988,N_16846);
and U17046 (N_17046,N_16807,N_16930);
xor U17047 (N_17047,N_16993,N_16830);
nand U17048 (N_17048,N_16892,N_16804);
or U17049 (N_17049,N_16979,N_16862);
or U17050 (N_17050,N_16903,N_16951);
nor U17051 (N_17051,N_16895,N_16835);
nand U17052 (N_17052,N_16856,N_16864);
xnor U17053 (N_17053,N_16996,N_16959);
nand U17054 (N_17054,N_16909,N_16983);
nor U17055 (N_17055,N_16987,N_16875);
nand U17056 (N_17056,N_16985,N_16998);
or U17057 (N_17057,N_16916,N_16837);
nor U17058 (N_17058,N_16887,N_16899);
nand U17059 (N_17059,N_16970,N_16870);
xor U17060 (N_17060,N_16908,N_16843);
or U17061 (N_17061,N_16984,N_16957);
xnor U17062 (N_17062,N_16890,N_16910);
xnor U17063 (N_17063,N_16912,N_16841);
nand U17064 (N_17064,N_16803,N_16879);
nor U17065 (N_17065,N_16961,N_16949);
nand U17066 (N_17066,N_16978,N_16878);
nor U17067 (N_17067,N_16896,N_16877);
and U17068 (N_17068,N_16839,N_16833);
nand U17069 (N_17069,N_16886,N_16915);
xnor U17070 (N_17070,N_16813,N_16981);
and U17071 (N_17071,N_16806,N_16898);
nand U17072 (N_17072,N_16995,N_16816);
xor U17073 (N_17073,N_16999,N_16880);
and U17074 (N_17074,N_16920,N_16986);
xnor U17075 (N_17075,N_16901,N_16838);
nor U17076 (N_17076,N_16902,N_16855);
xnor U17077 (N_17077,N_16824,N_16955);
nand U17078 (N_17078,N_16850,N_16964);
and U17079 (N_17079,N_16931,N_16911);
nand U17080 (N_17080,N_16810,N_16859);
nand U17081 (N_17081,N_16992,N_16805);
or U17082 (N_17082,N_16818,N_16948);
and U17083 (N_17083,N_16926,N_16971);
xnor U17084 (N_17084,N_16900,N_16823);
xor U17085 (N_17085,N_16811,N_16852);
nand U17086 (N_17086,N_16857,N_16933);
nor U17087 (N_17087,N_16958,N_16888);
or U17088 (N_17088,N_16963,N_16867);
xnor U17089 (N_17089,N_16976,N_16894);
or U17090 (N_17090,N_16845,N_16927);
nand U17091 (N_17091,N_16814,N_16952);
xor U17092 (N_17092,N_16802,N_16932);
xnor U17093 (N_17093,N_16934,N_16980);
xnor U17094 (N_17094,N_16950,N_16907);
or U17095 (N_17095,N_16849,N_16842);
nand U17096 (N_17096,N_16866,N_16884);
and U17097 (N_17097,N_16873,N_16929);
xor U17098 (N_17098,N_16940,N_16975);
nor U17099 (N_17099,N_16962,N_16820);
nand U17100 (N_17100,N_16951,N_16911);
and U17101 (N_17101,N_16966,N_16992);
or U17102 (N_17102,N_16815,N_16968);
nor U17103 (N_17103,N_16967,N_16809);
nor U17104 (N_17104,N_16894,N_16878);
and U17105 (N_17105,N_16835,N_16930);
or U17106 (N_17106,N_16949,N_16808);
and U17107 (N_17107,N_16977,N_16982);
nor U17108 (N_17108,N_16913,N_16993);
or U17109 (N_17109,N_16914,N_16942);
xor U17110 (N_17110,N_16957,N_16840);
nor U17111 (N_17111,N_16981,N_16841);
nor U17112 (N_17112,N_16814,N_16858);
nand U17113 (N_17113,N_16956,N_16935);
nand U17114 (N_17114,N_16986,N_16993);
or U17115 (N_17115,N_16929,N_16980);
nor U17116 (N_17116,N_16875,N_16899);
xnor U17117 (N_17117,N_16902,N_16926);
xor U17118 (N_17118,N_16937,N_16978);
nand U17119 (N_17119,N_16965,N_16976);
xnor U17120 (N_17120,N_16863,N_16837);
and U17121 (N_17121,N_16991,N_16854);
and U17122 (N_17122,N_16960,N_16891);
nor U17123 (N_17123,N_16896,N_16847);
nand U17124 (N_17124,N_16973,N_16854);
or U17125 (N_17125,N_16988,N_16882);
and U17126 (N_17126,N_16885,N_16837);
xor U17127 (N_17127,N_16860,N_16883);
xor U17128 (N_17128,N_16944,N_16871);
nand U17129 (N_17129,N_16820,N_16972);
xor U17130 (N_17130,N_16887,N_16897);
nand U17131 (N_17131,N_16807,N_16824);
xnor U17132 (N_17132,N_16952,N_16848);
xnor U17133 (N_17133,N_16803,N_16821);
nor U17134 (N_17134,N_16949,N_16896);
or U17135 (N_17135,N_16992,N_16923);
and U17136 (N_17136,N_16946,N_16905);
and U17137 (N_17137,N_16908,N_16871);
nand U17138 (N_17138,N_16811,N_16990);
nor U17139 (N_17139,N_16830,N_16920);
xor U17140 (N_17140,N_16938,N_16824);
xnor U17141 (N_17141,N_16887,N_16941);
and U17142 (N_17142,N_16965,N_16966);
or U17143 (N_17143,N_16815,N_16922);
and U17144 (N_17144,N_16868,N_16877);
and U17145 (N_17145,N_16947,N_16872);
xor U17146 (N_17146,N_16961,N_16881);
xor U17147 (N_17147,N_16843,N_16917);
nor U17148 (N_17148,N_16943,N_16883);
or U17149 (N_17149,N_16972,N_16807);
or U17150 (N_17150,N_16812,N_16965);
and U17151 (N_17151,N_16999,N_16822);
and U17152 (N_17152,N_16991,N_16893);
nor U17153 (N_17153,N_16955,N_16919);
and U17154 (N_17154,N_16954,N_16809);
and U17155 (N_17155,N_16876,N_16820);
nand U17156 (N_17156,N_16876,N_16879);
or U17157 (N_17157,N_16826,N_16978);
or U17158 (N_17158,N_16856,N_16903);
or U17159 (N_17159,N_16985,N_16905);
xor U17160 (N_17160,N_16960,N_16947);
xor U17161 (N_17161,N_16933,N_16929);
and U17162 (N_17162,N_16997,N_16969);
nand U17163 (N_17163,N_16817,N_16874);
nand U17164 (N_17164,N_16823,N_16878);
and U17165 (N_17165,N_16996,N_16932);
or U17166 (N_17166,N_16855,N_16830);
and U17167 (N_17167,N_16888,N_16850);
and U17168 (N_17168,N_16951,N_16912);
nor U17169 (N_17169,N_16926,N_16828);
nor U17170 (N_17170,N_16865,N_16883);
or U17171 (N_17171,N_16863,N_16881);
or U17172 (N_17172,N_16914,N_16964);
and U17173 (N_17173,N_16881,N_16970);
and U17174 (N_17174,N_16969,N_16917);
xor U17175 (N_17175,N_16893,N_16837);
or U17176 (N_17176,N_16840,N_16954);
or U17177 (N_17177,N_16970,N_16888);
xor U17178 (N_17178,N_16876,N_16970);
nor U17179 (N_17179,N_16848,N_16948);
or U17180 (N_17180,N_16893,N_16833);
and U17181 (N_17181,N_16881,N_16813);
xor U17182 (N_17182,N_16992,N_16990);
nand U17183 (N_17183,N_16809,N_16820);
nand U17184 (N_17184,N_16997,N_16881);
or U17185 (N_17185,N_16902,N_16991);
nor U17186 (N_17186,N_16829,N_16970);
or U17187 (N_17187,N_16980,N_16856);
or U17188 (N_17188,N_16960,N_16987);
nand U17189 (N_17189,N_16935,N_16933);
nor U17190 (N_17190,N_16899,N_16933);
or U17191 (N_17191,N_16874,N_16875);
nand U17192 (N_17192,N_16816,N_16877);
xor U17193 (N_17193,N_16921,N_16977);
nand U17194 (N_17194,N_16836,N_16888);
nand U17195 (N_17195,N_16987,N_16860);
nand U17196 (N_17196,N_16898,N_16935);
nor U17197 (N_17197,N_16931,N_16995);
xor U17198 (N_17198,N_16953,N_16806);
nand U17199 (N_17199,N_16889,N_16826);
or U17200 (N_17200,N_17005,N_17053);
nand U17201 (N_17201,N_17175,N_17024);
or U17202 (N_17202,N_17064,N_17004);
and U17203 (N_17203,N_17197,N_17145);
nor U17204 (N_17204,N_17109,N_17090);
xnor U17205 (N_17205,N_17104,N_17194);
nand U17206 (N_17206,N_17036,N_17164);
or U17207 (N_17207,N_17079,N_17050);
and U17208 (N_17208,N_17096,N_17022);
xnor U17209 (N_17209,N_17018,N_17103);
or U17210 (N_17210,N_17001,N_17159);
nor U17211 (N_17211,N_17180,N_17075);
nor U17212 (N_17212,N_17045,N_17150);
or U17213 (N_17213,N_17156,N_17152);
nand U17214 (N_17214,N_17111,N_17063);
or U17215 (N_17215,N_17049,N_17040);
nand U17216 (N_17216,N_17163,N_17089);
or U17217 (N_17217,N_17148,N_17085);
nor U17218 (N_17218,N_17121,N_17080);
xnor U17219 (N_17219,N_17171,N_17187);
nand U17220 (N_17220,N_17182,N_17110);
nor U17221 (N_17221,N_17174,N_17169);
nor U17222 (N_17222,N_17141,N_17155);
or U17223 (N_17223,N_17067,N_17165);
or U17224 (N_17224,N_17115,N_17077);
or U17225 (N_17225,N_17138,N_17170);
nor U17226 (N_17226,N_17195,N_17006);
or U17227 (N_17227,N_17123,N_17086);
or U17228 (N_17228,N_17037,N_17139);
or U17229 (N_17229,N_17062,N_17076);
nand U17230 (N_17230,N_17185,N_17114);
or U17231 (N_17231,N_17027,N_17088);
nand U17232 (N_17232,N_17012,N_17025);
or U17233 (N_17233,N_17199,N_17132);
nor U17234 (N_17234,N_17071,N_17052);
and U17235 (N_17235,N_17046,N_17124);
nor U17236 (N_17236,N_17003,N_17192);
and U17237 (N_17237,N_17065,N_17116);
or U17238 (N_17238,N_17140,N_17028);
nor U17239 (N_17239,N_17032,N_17078);
xnor U17240 (N_17240,N_17144,N_17134);
nor U17241 (N_17241,N_17157,N_17137);
nor U17242 (N_17242,N_17044,N_17007);
xnor U17243 (N_17243,N_17029,N_17017);
xor U17244 (N_17244,N_17033,N_17035);
xor U17245 (N_17245,N_17016,N_17122);
nand U17246 (N_17246,N_17011,N_17093);
nand U17247 (N_17247,N_17092,N_17095);
or U17248 (N_17248,N_17034,N_17055);
or U17249 (N_17249,N_17069,N_17191);
nand U17250 (N_17250,N_17048,N_17178);
nand U17251 (N_17251,N_17002,N_17162);
xnor U17252 (N_17252,N_17153,N_17060);
and U17253 (N_17253,N_17176,N_17146);
nand U17254 (N_17254,N_17151,N_17125);
nand U17255 (N_17255,N_17031,N_17010);
xor U17256 (N_17256,N_17008,N_17068);
or U17257 (N_17257,N_17105,N_17193);
nand U17258 (N_17258,N_17000,N_17158);
xor U17259 (N_17259,N_17147,N_17081);
or U17260 (N_17260,N_17177,N_17118);
nand U17261 (N_17261,N_17113,N_17117);
xnor U17262 (N_17262,N_17020,N_17043);
xor U17263 (N_17263,N_17098,N_17184);
or U17264 (N_17264,N_17106,N_17054);
xor U17265 (N_17265,N_17066,N_17051);
xor U17266 (N_17266,N_17021,N_17030);
xnor U17267 (N_17267,N_17131,N_17014);
xor U17268 (N_17268,N_17070,N_17019);
nand U17269 (N_17269,N_17057,N_17087);
nor U17270 (N_17270,N_17190,N_17179);
xor U17271 (N_17271,N_17058,N_17108);
xnor U17272 (N_17272,N_17059,N_17188);
nor U17273 (N_17273,N_17168,N_17133);
nand U17274 (N_17274,N_17130,N_17183);
and U17275 (N_17275,N_17099,N_17047);
nand U17276 (N_17276,N_17100,N_17026);
and U17277 (N_17277,N_17107,N_17112);
and U17278 (N_17278,N_17009,N_17102);
and U17279 (N_17279,N_17198,N_17042);
and U17280 (N_17280,N_17056,N_17142);
nor U17281 (N_17281,N_17120,N_17097);
and U17282 (N_17282,N_17082,N_17101);
or U17283 (N_17283,N_17166,N_17186);
nand U17284 (N_17284,N_17038,N_17084);
nor U17285 (N_17285,N_17160,N_17127);
and U17286 (N_17286,N_17074,N_17041);
and U17287 (N_17287,N_17083,N_17073);
nor U17288 (N_17288,N_17015,N_17167);
or U17289 (N_17289,N_17136,N_17172);
nor U17290 (N_17290,N_17061,N_17189);
or U17291 (N_17291,N_17143,N_17196);
or U17292 (N_17292,N_17135,N_17072);
nor U17293 (N_17293,N_17119,N_17173);
and U17294 (N_17294,N_17126,N_17129);
nor U17295 (N_17295,N_17154,N_17181);
nor U17296 (N_17296,N_17128,N_17161);
and U17297 (N_17297,N_17039,N_17013);
xnor U17298 (N_17298,N_17094,N_17149);
nand U17299 (N_17299,N_17091,N_17023);
or U17300 (N_17300,N_17194,N_17164);
and U17301 (N_17301,N_17039,N_17086);
or U17302 (N_17302,N_17126,N_17171);
nand U17303 (N_17303,N_17149,N_17167);
or U17304 (N_17304,N_17025,N_17142);
xor U17305 (N_17305,N_17091,N_17150);
nand U17306 (N_17306,N_17171,N_17014);
nor U17307 (N_17307,N_17077,N_17084);
nand U17308 (N_17308,N_17039,N_17176);
nand U17309 (N_17309,N_17081,N_17188);
nor U17310 (N_17310,N_17008,N_17140);
or U17311 (N_17311,N_17060,N_17054);
nand U17312 (N_17312,N_17199,N_17023);
or U17313 (N_17313,N_17178,N_17177);
or U17314 (N_17314,N_17030,N_17000);
xor U17315 (N_17315,N_17198,N_17033);
nor U17316 (N_17316,N_17083,N_17126);
nor U17317 (N_17317,N_17154,N_17015);
and U17318 (N_17318,N_17149,N_17119);
xnor U17319 (N_17319,N_17155,N_17086);
nor U17320 (N_17320,N_17013,N_17176);
or U17321 (N_17321,N_17059,N_17192);
nor U17322 (N_17322,N_17062,N_17150);
nor U17323 (N_17323,N_17102,N_17116);
xor U17324 (N_17324,N_17160,N_17055);
nand U17325 (N_17325,N_17005,N_17111);
xnor U17326 (N_17326,N_17134,N_17128);
nor U17327 (N_17327,N_17098,N_17171);
nor U17328 (N_17328,N_17084,N_17097);
or U17329 (N_17329,N_17028,N_17113);
xor U17330 (N_17330,N_17113,N_17002);
and U17331 (N_17331,N_17068,N_17035);
xor U17332 (N_17332,N_17084,N_17135);
and U17333 (N_17333,N_17042,N_17095);
and U17334 (N_17334,N_17084,N_17028);
xor U17335 (N_17335,N_17101,N_17139);
nand U17336 (N_17336,N_17139,N_17050);
xor U17337 (N_17337,N_17104,N_17010);
nor U17338 (N_17338,N_17019,N_17100);
and U17339 (N_17339,N_17158,N_17118);
and U17340 (N_17340,N_17120,N_17085);
or U17341 (N_17341,N_17055,N_17129);
nor U17342 (N_17342,N_17005,N_17083);
and U17343 (N_17343,N_17153,N_17072);
and U17344 (N_17344,N_17197,N_17083);
or U17345 (N_17345,N_17189,N_17185);
and U17346 (N_17346,N_17149,N_17024);
or U17347 (N_17347,N_17002,N_17034);
xor U17348 (N_17348,N_17007,N_17099);
nand U17349 (N_17349,N_17073,N_17031);
and U17350 (N_17350,N_17130,N_17173);
xnor U17351 (N_17351,N_17167,N_17196);
xnor U17352 (N_17352,N_17042,N_17069);
nor U17353 (N_17353,N_17127,N_17062);
xnor U17354 (N_17354,N_17018,N_17188);
nor U17355 (N_17355,N_17043,N_17105);
nor U17356 (N_17356,N_17185,N_17097);
nand U17357 (N_17357,N_17042,N_17178);
xor U17358 (N_17358,N_17089,N_17176);
nand U17359 (N_17359,N_17034,N_17162);
nand U17360 (N_17360,N_17066,N_17171);
or U17361 (N_17361,N_17066,N_17019);
nor U17362 (N_17362,N_17048,N_17037);
and U17363 (N_17363,N_17077,N_17174);
and U17364 (N_17364,N_17082,N_17054);
nor U17365 (N_17365,N_17076,N_17192);
or U17366 (N_17366,N_17005,N_17010);
and U17367 (N_17367,N_17123,N_17100);
nand U17368 (N_17368,N_17177,N_17166);
or U17369 (N_17369,N_17133,N_17103);
nor U17370 (N_17370,N_17178,N_17021);
and U17371 (N_17371,N_17031,N_17158);
nor U17372 (N_17372,N_17011,N_17017);
or U17373 (N_17373,N_17108,N_17019);
nand U17374 (N_17374,N_17044,N_17097);
nor U17375 (N_17375,N_17092,N_17014);
or U17376 (N_17376,N_17041,N_17100);
xnor U17377 (N_17377,N_17171,N_17034);
and U17378 (N_17378,N_17166,N_17179);
nand U17379 (N_17379,N_17195,N_17133);
or U17380 (N_17380,N_17000,N_17089);
nor U17381 (N_17381,N_17080,N_17098);
or U17382 (N_17382,N_17091,N_17103);
nand U17383 (N_17383,N_17015,N_17017);
or U17384 (N_17384,N_17117,N_17094);
xor U17385 (N_17385,N_17079,N_17033);
xor U17386 (N_17386,N_17166,N_17127);
or U17387 (N_17387,N_17083,N_17189);
or U17388 (N_17388,N_17052,N_17125);
nor U17389 (N_17389,N_17188,N_17066);
and U17390 (N_17390,N_17075,N_17077);
or U17391 (N_17391,N_17071,N_17065);
and U17392 (N_17392,N_17014,N_17011);
nor U17393 (N_17393,N_17157,N_17171);
or U17394 (N_17394,N_17177,N_17043);
and U17395 (N_17395,N_17122,N_17195);
and U17396 (N_17396,N_17038,N_17175);
nor U17397 (N_17397,N_17042,N_17175);
and U17398 (N_17398,N_17119,N_17199);
nand U17399 (N_17399,N_17110,N_17001);
or U17400 (N_17400,N_17200,N_17268);
nand U17401 (N_17401,N_17355,N_17220);
or U17402 (N_17402,N_17300,N_17247);
and U17403 (N_17403,N_17256,N_17258);
nand U17404 (N_17404,N_17282,N_17319);
xnor U17405 (N_17405,N_17295,N_17287);
nand U17406 (N_17406,N_17371,N_17294);
and U17407 (N_17407,N_17390,N_17380);
or U17408 (N_17408,N_17352,N_17350);
xor U17409 (N_17409,N_17316,N_17344);
and U17410 (N_17410,N_17323,N_17237);
and U17411 (N_17411,N_17213,N_17398);
xnor U17412 (N_17412,N_17228,N_17288);
xnor U17413 (N_17413,N_17250,N_17266);
and U17414 (N_17414,N_17364,N_17299);
or U17415 (N_17415,N_17331,N_17212);
or U17416 (N_17416,N_17240,N_17204);
or U17417 (N_17417,N_17328,N_17326);
or U17418 (N_17418,N_17394,N_17243);
nand U17419 (N_17419,N_17313,N_17278);
and U17420 (N_17420,N_17361,N_17310);
nand U17421 (N_17421,N_17233,N_17261);
xnor U17422 (N_17422,N_17297,N_17277);
and U17423 (N_17423,N_17242,N_17231);
nand U17424 (N_17424,N_17248,N_17329);
or U17425 (N_17425,N_17254,N_17321);
xor U17426 (N_17426,N_17357,N_17269);
or U17427 (N_17427,N_17202,N_17345);
or U17428 (N_17428,N_17367,N_17351);
and U17429 (N_17429,N_17301,N_17255);
xor U17430 (N_17430,N_17397,N_17377);
nor U17431 (N_17431,N_17298,N_17211);
nand U17432 (N_17432,N_17284,N_17339);
and U17433 (N_17433,N_17221,N_17388);
or U17434 (N_17434,N_17386,N_17332);
nand U17435 (N_17435,N_17214,N_17385);
and U17436 (N_17436,N_17273,N_17320);
or U17437 (N_17437,N_17311,N_17260);
and U17438 (N_17438,N_17376,N_17285);
xnor U17439 (N_17439,N_17356,N_17263);
nand U17440 (N_17440,N_17370,N_17342);
xnor U17441 (N_17441,N_17252,N_17236);
nor U17442 (N_17442,N_17276,N_17373);
xnor U17443 (N_17443,N_17222,N_17271);
nand U17444 (N_17444,N_17217,N_17234);
nand U17445 (N_17445,N_17381,N_17218);
or U17446 (N_17446,N_17343,N_17379);
and U17447 (N_17447,N_17318,N_17224);
nor U17448 (N_17448,N_17229,N_17389);
nor U17449 (N_17449,N_17306,N_17235);
nand U17450 (N_17450,N_17334,N_17291);
xnor U17451 (N_17451,N_17227,N_17340);
nand U17452 (N_17452,N_17363,N_17374);
and U17453 (N_17453,N_17244,N_17360);
and U17454 (N_17454,N_17383,N_17289);
and U17455 (N_17455,N_17302,N_17286);
nand U17456 (N_17456,N_17265,N_17372);
xor U17457 (N_17457,N_17392,N_17362);
nor U17458 (N_17458,N_17209,N_17207);
or U17459 (N_17459,N_17353,N_17226);
nor U17460 (N_17460,N_17366,N_17293);
xor U17461 (N_17461,N_17270,N_17359);
nor U17462 (N_17462,N_17239,N_17280);
xnor U17463 (N_17463,N_17303,N_17206);
and U17464 (N_17464,N_17253,N_17307);
nand U17465 (N_17465,N_17395,N_17322);
nor U17466 (N_17466,N_17304,N_17230);
nand U17467 (N_17467,N_17232,N_17309);
or U17468 (N_17468,N_17396,N_17296);
nand U17469 (N_17469,N_17347,N_17315);
xor U17470 (N_17470,N_17216,N_17335);
nor U17471 (N_17471,N_17274,N_17384);
nor U17472 (N_17472,N_17382,N_17267);
or U17473 (N_17473,N_17308,N_17275);
xor U17474 (N_17474,N_17245,N_17251);
and U17475 (N_17475,N_17348,N_17333);
and U17476 (N_17476,N_17249,N_17312);
xor U17477 (N_17477,N_17257,N_17281);
nand U17478 (N_17478,N_17219,N_17241);
nand U17479 (N_17479,N_17337,N_17279);
and U17480 (N_17480,N_17349,N_17259);
nand U17481 (N_17481,N_17210,N_17246);
nand U17482 (N_17482,N_17292,N_17205);
or U17483 (N_17483,N_17324,N_17264);
nand U17484 (N_17484,N_17375,N_17201);
nand U17485 (N_17485,N_17223,N_17391);
or U17486 (N_17486,N_17225,N_17262);
or U17487 (N_17487,N_17365,N_17325);
nand U17488 (N_17488,N_17238,N_17354);
and U17489 (N_17489,N_17378,N_17341);
nor U17490 (N_17490,N_17290,N_17327);
xor U17491 (N_17491,N_17305,N_17393);
nand U17492 (N_17492,N_17358,N_17387);
nand U17493 (N_17493,N_17336,N_17330);
xnor U17494 (N_17494,N_17399,N_17208);
and U17495 (N_17495,N_17338,N_17203);
nand U17496 (N_17496,N_17314,N_17317);
and U17497 (N_17497,N_17283,N_17346);
and U17498 (N_17498,N_17215,N_17368);
xnor U17499 (N_17499,N_17272,N_17369);
nor U17500 (N_17500,N_17236,N_17243);
and U17501 (N_17501,N_17396,N_17387);
nand U17502 (N_17502,N_17366,N_17327);
nor U17503 (N_17503,N_17354,N_17386);
xor U17504 (N_17504,N_17252,N_17235);
or U17505 (N_17505,N_17242,N_17338);
and U17506 (N_17506,N_17397,N_17294);
xor U17507 (N_17507,N_17311,N_17392);
nor U17508 (N_17508,N_17291,N_17363);
nand U17509 (N_17509,N_17296,N_17222);
and U17510 (N_17510,N_17204,N_17252);
xnor U17511 (N_17511,N_17357,N_17264);
and U17512 (N_17512,N_17341,N_17229);
nand U17513 (N_17513,N_17361,N_17291);
or U17514 (N_17514,N_17237,N_17324);
nand U17515 (N_17515,N_17287,N_17274);
xor U17516 (N_17516,N_17221,N_17356);
and U17517 (N_17517,N_17387,N_17371);
nor U17518 (N_17518,N_17260,N_17274);
nor U17519 (N_17519,N_17256,N_17292);
xor U17520 (N_17520,N_17377,N_17360);
nand U17521 (N_17521,N_17355,N_17239);
nor U17522 (N_17522,N_17202,N_17379);
or U17523 (N_17523,N_17333,N_17241);
or U17524 (N_17524,N_17293,N_17290);
and U17525 (N_17525,N_17321,N_17206);
or U17526 (N_17526,N_17384,N_17254);
nand U17527 (N_17527,N_17303,N_17324);
and U17528 (N_17528,N_17323,N_17218);
xnor U17529 (N_17529,N_17338,N_17356);
nor U17530 (N_17530,N_17259,N_17276);
or U17531 (N_17531,N_17304,N_17275);
nor U17532 (N_17532,N_17318,N_17217);
nand U17533 (N_17533,N_17378,N_17352);
and U17534 (N_17534,N_17312,N_17215);
nand U17535 (N_17535,N_17293,N_17244);
or U17536 (N_17536,N_17375,N_17379);
nor U17537 (N_17537,N_17231,N_17264);
nand U17538 (N_17538,N_17378,N_17327);
nor U17539 (N_17539,N_17378,N_17214);
or U17540 (N_17540,N_17277,N_17233);
nand U17541 (N_17541,N_17282,N_17217);
and U17542 (N_17542,N_17360,N_17205);
nand U17543 (N_17543,N_17209,N_17277);
and U17544 (N_17544,N_17346,N_17262);
xnor U17545 (N_17545,N_17339,N_17241);
xor U17546 (N_17546,N_17222,N_17294);
xor U17547 (N_17547,N_17399,N_17312);
and U17548 (N_17548,N_17338,N_17272);
and U17549 (N_17549,N_17371,N_17245);
nand U17550 (N_17550,N_17300,N_17329);
nor U17551 (N_17551,N_17371,N_17287);
xnor U17552 (N_17552,N_17368,N_17231);
and U17553 (N_17553,N_17361,N_17255);
or U17554 (N_17554,N_17346,N_17317);
and U17555 (N_17555,N_17381,N_17281);
xor U17556 (N_17556,N_17323,N_17330);
or U17557 (N_17557,N_17256,N_17398);
nor U17558 (N_17558,N_17335,N_17219);
or U17559 (N_17559,N_17317,N_17393);
nand U17560 (N_17560,N_17207,N_17308);
nand U17561 (N_17561,N_17393,N_17352);
nand U17562 (N_17562,N_17399,N_17382);
xnor U17563 (N_17563,N_17318,N_17322);
or U17564 (N_17564,N_17224,N_17286);
or U17565 (N_17565,N_17330,N_17296);
nand U17566 (N_17566,N_17224,N_17337);
nand U17567 (N_17567,N_17307,N_17382);
nand U17568 (N_17568,N_17362,N_17248);
nor U17569 (N_17569,N_17366,N_17302);
xnor U17570 (N_17570,N_17327,N_17265);
nand U17571 (N_17571,N_17395,N_17380);
xor U17572 (N_17572,N_17278,N_17355);
or U17573 (N_17573,N_17354,N_17206);
and U17574 (N_17574,N_17396,N_17313);
and U17575 (N_17575,N_17340,N_17294);
xor U17576 (N_17576,N_17245,N_17289);
and U17577 (N_17577,N_17255,N_17351);
xnor U17578 (N_17578,N_17374,N_17383);
or U17579 (N_17579,N_17361,N_17228);
xor U17580 (N_17580,N_17388,N_17328);
or U17581 (N_17581,N_17328,N_17217);
and U17582 (N_17582,N_17328,N_17255);
and U17583 (N_17583,N_17312,N_17390);
nor U17584 (N_17584,N_17246,N_17216);
and U17585 (N_17585,N_17362,N_17379);
nor U17586 (N_17586,N_17230,N_17211);
nand U17587 (N_17587,N_17347,N_17397);
xnor U17588 (N_17588,N_17266,N_17292);
xnor U17589 (N_17589,N_17265,N_17248);
nand U17590 (N_17590,N_17290,N_17266);
or U17591 (N_17591,N_17270,N_17253);
and U17592 (N_17592,N_17291,N_17336);
or U17593 (N_17593,N_17205,N_17283);
or U17594 (N_17594,N_17203,N_17328);
xnor U17595 (N_17595,N_17351,N_17370);
and U17596 (N_17596,N_17233,N_17367);
nand U17597 (N_17597,N_17340,N_17375);
nor U17598 (N_17598,N_17367,N_17210);
xor U17599 (N_17599,N_17283,N_17213);
xnor U17600 (N_17600,N_17413,N_17511);
nand U17601 (N_17601,N_17429,N_17463);
nand U17602 (N_17602,N_17566,N_17575);
nand U17603 (N_17603,N_17504,N_17508);
or U17604 (N_17604,N_17527,N_17441);
nand U17605 (N_17605,N_17414,N_17408);
and U17606 (N_17606,N_17590,N_17598);
nand U17607 (N_17607,N_17516,N_17451);
nand U17608 (N_17608,N_17595,N_17412);
xor U17609 (N_17609,N_17453,N_17418);
nand U17610 (N_17610,N_17407,N_17502);
nor U17611 (N_17611,N_17557,N_17553);
or U17612 (N_17612,N_17594,N_17515);
nor U17613 (N_17613,N_17548,N_17454);
nand U17614 (N_17614,N_17427,N_17499);
xnor U17615 (N_17615,N_17417,N_17443);
nor U17616 (N_17616,N_17561,N_17425);
nand U17617 (N_17617,N_17467,N_17474);
and U17618 (N_17618,N_17599,N_17529);
or U17619 (N_17619,N_17477,N_17591);
xnor U17620 (N_17620,N_17445,N_17531);
xnor U17621 (N_17621,N_17596,N_17469);
and U17622 (N_17622,N_17587,N_17448);
and U17623 (N_17623,N_17568,N_17593);
and U17624 (N_17624,N_17488,N_17479);
or U17625 (N_17625,N_17585,N_17570);
nor U17626 (N_17626,N_17549,N_17422);
nor U17627 (N_17627,N_17440,N_17567);
and U17628 (N_17628,N_17428,N_17468);
nor U17629 (N_17629,N_17520,N_17559);
xnor U17630 (N_17630,N_17457,N_17480);
nand U17631 (N_17631,N_17586,N_17489);
xor U17632 (N_17632,N_17524,N_17534);
and U17633 (N_17633,N_17547,N_17551);
or U17634 (N_17634,N_17470,N_17552);
or U17635 (N_17635,N_17404,N_17563);
nand U17636 (N_17636,N_17434,N_17496);
and U17637 (N_17637,N_17526,N_17461);
nand U17638 (N_17638,N_17406,N_17577);
xor U17639 (N_17639,N_17439,N_17485);
and U17640 (N_17640,N_17539,N_17487);
and U17641 (N_17641,N_17535,N_17426);
nand U17642 (N_17642,N_17532,N_17554);
nand U17643 (N_17643,N_17583,N_17494);
nor U17644 (N_17644,N_17490,N_17458);
nand U17645 (N_17645,N_17546,N_17576);
nand U17646 (N_17646,N_17436,N_17400);
or U17647 (N_17647,N_17541,N_17538);
nand U17648 (N_17648,N_17403,N_17522);
and U17649 (N_17649,N_17423,N_17543);
nand U17650 (N_17650,N_17491,N_17537);
and U17651 (N_17651,N_17518,N_17588);
nor U17652 (N_17652,N_17475,N_17495);
xor U17653 (N_17653,N_17493,N_17444);
or U17654 (N_17654,N_17478,N_17500);
nor U17655 (N_17655,N_17517,N_17424);
or U17656 (N_17656,N_17569,N_17416);
and U17657 (N_17657,N_17510,N_17571);
nand U17658 (N_17658,N_17497,N_17545);
nand U17659 (N_17659,N_17462,N_17579);
nor U17660 (N_17660,N_17580,N_17581);
xor U17661 (N_17661,N_17564,N_17523);
nor U17662 (N_17662,N_17574,N_17466);
xnor U17663 (N_17663,N_17556,N_17481);
xor U17664 (N_17664,N_17438,N_17558);
nand U17665 (N_17665,N_17452,N_17456);
xnor U17666 (N_17666,N_17512,N_17446);
and U17667 (N_17667,N_17437,N_17505);
or U17668 (N_17668,N_17533,N_17540);
or U17669 (N_17669,N_17514,N_17459);
and U17670 (N_17670,N_17447,N_17435);
nand U17671 (N_17671,N_17582,N_17509);
nor U17672 (N_17672,N_17433,N_17460);
and U17673 (N_17673,N_17419,N_17550);
or U17674 (N_17674,N_17415,N_17430);
and U17675 (N_17675,N_17409,N_17420);
and U17676 (N_17676,N_17401,N_17483);
nand U17677 (N_17677,N_17410,N_17486);
nand U17678 (N_17678,N_17449,N_17544);
xor U17679 (N_17679,N_17542,N_17572);
and U17680 (N_17680,N_17562,N_17578);
or U17681 (N_17681,N_17492,N_17536);
or U17682 (N_17682,N_17521,N_17464);
or U17683 (N_17683,N_17455,N_17501);
or U17684 (N_17684,N_17506,N_17589);
and U17685 (N_17685,N_17473,N_17573);
xnor U17686 (N_17686,N_17476,N_17482);
and U17687 (N_17687,N_17472,N_17565);
nand U17688 (N_17688,N_17442,N_17530);
nor U17689 (N_17689,N_17513,N_17411);
or U17690 (N_17690,N_17484,N_17405);
or U17691 (N_17691,N_17432,N_17592);
nor U17692 (N_17692,N_17431,N_17555);
nand U17693 (N_17693,N_17525,N_17507);
or U17694 (N_17694,N_17498,N_17471);
and U17695 (N_17695,N_17560,N_17465);
or U17696 (N_17696,N_17503,N_17519);
or U17697 (N_17697,N_17597,N_17421);
or U17698 (N_17698,N_17402,N_17450);
nand U17699 (N_17699,N_17528,N_17584);
and U17700 (N_17700,N_17450,N_17425);
nor U17701 (N_17701,N_17540,N_17591);
nand U17702 (N_17702,N_17592,N_17403);
nand U17703 (N_17703,N_17434,N_17506);
or U17704 (N_17704,N_17482,N_17544);
and U17705 (N_17705,N_17452,N_17435);
or U17706 (N_17706,N_17514,N_17544);
xnor U17707 (N_17707,N_17489,N_17526);
xnor U17708 (N_17708,N_17422,N_17535);
and U17709 (N_17709,N_17438,N_17423);
or U17710 (N_17710,N_17567,N_17570);
or U17711 (N_17711,N_17514,N_17467);
nor U17712 (N_17712,N_17480,N_17463);
xnor U17713 (N_17713,N_17432,N_17405);
nand U17714 (N_17714,N_17487,N_17409);
xnor U17715 (N_17715,N_17459,N_17531);
nor U17716 (N_17716,N_17417,N_17482);
xnor U17717 (N_17717,N_17539,N_17594);
xnor U17718 (N_17718,N_17487,N_17576);
nor U17719 (N_17719,N_17563,N_17497);
and U17720 (N_17720,N_17442,N_17555);
or U17721 (N_17721,N_17568,N_17566);
and U17722 (N_17722,N_17407,N_17448);
nor U17723 (N_17723,N_17431,N_17567);
nand U17724 (N_17724,N_17461,N_17587);
nor U17725 (N_17725,N_17414,N_17505);
nand U17726 (N_17726,N_17477,N_17516);
and U17727 (N_17727,N_17580,N_17459);
or U17728 (N_17728,N_17599,N_17531);
xor U17729 (N_17729,N_17402,N_17574);
nor U17730 (N_17730,N_17483,N_17428);
and U17731 (N_17731,N_17438,N_17569);
nand U17732 (N_17732,N_17454,N_17587);
nand U17733 (N_17733,N_17549,N_17421);
nor U17734 (N_17734,N_17505,N_17554);
nand U17735 (N_17735,N_17499,N_17432);
nor U17736 (N_17736,N_17487,N_17462);
nor U17737 (N_17737,N_17430,N_17472);
xnor U17738 (N_17738,N_17426,N_17561);
nand U17739 (N_17739,N_17535,N_17471);
or U17740 (N_17740,N_17455,N_17497);
nor U17741 (N_17741,N_17470,N_17426);
xnor U17742 (N_17742,N_17595,N_17504);
nor U17743 (N_17743,N_17435,N_17464);
nor U17744 (N_17744,N_17582,N_17566);
and U17745 (N_17745,N_17475,N_17449);
nor U17746 (N_17746,N_17546,N_17406);
nand U17747 (N_17747,N_17546,N_17543);
and U17748 (N_17748,N_17484,N_17582);
nor U17749 (N_17749,N_17523,N_17528);
xor U17750 (N_17750,N_17506,N_17494);
nor U17751 (N_17751,N_17479,N_17590);
nand U17752 (N_17752,N_17420,N_17414);
nor U17753 (N_17753,N_17449,N_17560);
nand U17754 (N_17754,N_17504,N_17459);
or U17755 (N_17755,N_17536,N_17500);
nand U17756 (N_17756,N_17534,N_17434);
nand U17757 (N_17757,N_17485,N_17476);
xor U17758 (N_17758,N_17559,N_17529);
xnor U17759 (N_17759,N_17482,N_17572);
nand U17760 (N_17760,N_17526,N_17495);
nand U17761 (N_17761,N_17599,N_17501);
nor U17762 (N_17762,N_17429,N_17510);
xnor U17763 (N_17763,N_17560,N_17553);
or U17764 (N_17764,N_17492,N_17495);
xnor U17765 (N_17765,N_17419,N_17417);
xor U17766 (N_17766,N_17433,N_17409);
and U17767 (N_17767,N_17523,N_17426);
and U17768 (N_17768,N_17442,N_17554);
and U17769 (N_17769,N_17473,N_17458);
nand U17770 (N_17770,N_17553,N_17498);
or U17771 (N_17771,N_17512,N_17485);
or U17772 (N_17772,N_17475,N_17567);
and U17773 (N_17773,N_17420,N_17416);
nand U17774 (N_17774,N_17564,N_17596);
nand U17775 (N_17775,N_17408,N_17485);
and U17776 (N_17776,N_17538,N_17510);
xnor U17777 (N_17777,N_17410,N_17546);
or U17778 (N_17778,N_17455,N_17464);
nand U17779 (N_17779,N_17542,N_17465);
nor U17780 (N_17780,N_17500,N_17485);
xnor U17781 (N_17781,N_17474,N_17447);
or U17782 (N_17782,N_17428,N_17436);
or U17783 (N_17783,N_17469,N_17498);
nand U17784 (N_17784,N_17472,N_17489);
nor U17785 (N_17785,N_17592,N_17439);
nor U17786 (N_17786,N_17490,N_17410);
nor U17787 (N_17787,N_17554,N_17451);
xnor U17788 (N_17788,N_17560,N_17502);
or U17789 (N_17789,N_17502,N_17426);
or U17790 (N_17790,N_17555,N_17529);
xnor U17791 (N_17791,N_17466,N_17544);
xnor U17792 (N_17792,N_17442,N_17583);
xnor U17793 (N_17793,N_17501,N_17572);
xnor U17794 (N_17794,N_17470,N_17436);
nor U17795 (N_17795,N_17581,N_17432);
nor U17796 (N_17796,N_17553,N_17484);
xnor U17797 (N_17797,N_17409,N_17504);
or U17798 (N_17798,N_17504,N_17441);
xnor U17799 (N_17799,N_17556,N_17540);
or U17800 (N_17800,N_17632,N_17664);
nor U17801 (N_17801,N_17657,N_17637);
and U17802 (N_17802,N_17652,N_17715);
nor U17803 (N_17803,N_17734,N_17675);
nor U17804 (N_17804,N_17741,N_17693);
and U17805 (N_17805,N_17682,N_17759);
or U17806 (N_17806,N_17781,N_17604);
and U17807 (N_17807,N_17721,N_17718);
nand U17808 (N_17808,N_17736,N_17738);
or U17809 (N_17809,N_17614,N_17622);
or U17810 (N_17810,N_17719,N_17671);
nand U17811 (N_17811,N_17737,N_17603);
or U17812 (N_17812,N_17793,N_17768);
nor U17813 (N_17813,N_17717,N_17624);
xnor U17814 (N_17814,N_17635,N_17654);
xor U17815 (N_17815,N_17771,N_17679);
xor U17816 (N_17816,N_17714,N_17748);
and U17817 (N_17817,N_17611,N_17758);
and U17818 (N_17818,N_17647,N_17623);
nor U17819 (N_17819,N_17764,N_17602);
nor U17820 (N_17820,N_17687,N_17605);
or U17821 (N_17821,N_17750,N_17754);
or U17822 (N_17822,N_17711,N_17673);
and U17823 (N_17823,N_17629,N_17615);
and U17824 (N_17824,N_17722,N_17643);
nand U17825 (N_17825,N_17767,N_17696);
or U17826 (N_17826,N_17630,N_17704);
nand U17827 (N_17827,N_17731,N_17742);
and U17828 (N_17828,N_17695,N_17620);
xnor U17829 (N_17829,N_17668,N_17601);
xnor U17830 (N_17830,N_17728,N_17653);
or U17831 (N_17831,N_17669,N_17778);
and U17832 (N_17832,N_17708,N_17600);
or U17833 (N_17833,N_17660,N_17612);
and U17834 (N_17834,N_17785,N_17766);
and U17835 (N_17835,N_17650,N_17729);
nand U17836 (N_17836,N_17656,N_17783);
xor U17837 (N_17837,N_17712,N_17709);
xor U17838 (N_17838,N_17747,N_17658);
nor U17839 (N_17839,N_17792,N_17757);
or U17840 (N_17840,N_17752,N_17725);
nor U17841 (N_17841,N_17774,N_17617);
or U17842 (N_17842,N_17649,N_17703);
nor U17843 (N_17843,N_17723,N_17716);
and U17844 (N_17844,N_17796,N_17616);
or U17845 (N_17845,N_17706,N_17610);
nand U17846 (N_17846,N_17694,N_17772);
or U17847 (N_17847,N_17638,N_17628);
or U17848 (N_17848,N_17676,N_17730);
nand U17849 (N_17849,N_17626,N_17769);
nand U17850 (N_17850,N_17776,N_17689);
nand U17851 (N_17851,N_17684,N_17797);
xor U17852 (N_17852,N_17688,N_17681);
and U17853 (N_17853,N_17698,N_17640);
or U17854 (N_17854,N_17782,N_17756);
xnor U17855 (N_17855,N_17697,N_17621);
or U17856 (N_17856,N_17701,N_17775);
nand U17857 (N_17857,N_17740,N_17609);
and U17858 (N_17858,N_17700,N_17753);
and U17859 (N_17859,N_17791,N_17648);
nand U17860 (N_17860,N_17780,N_17606);
or U17861 (N_17861,N_17659,N_17705);
xnor U17862 (N_17862,N_17674,N_17779);
xnor U17863 (N_17863,N_17618,N_17642);
and U17864 (N_17864,N_17627,N_17651);
nand U17865 (N_17865,N_17670,N_17678);
nand U17866 (N_17866,N_17765,N_17777);
nand U17867 (N_17867,N_17744,N_17631);
or U17868 (N_17868,N_17644,N_17691);
xor U17869 (N_17869,N_17661,N_17667);
nand U17870 (N_17870,N_17639,N_17686);
nor U17871 (N_17871,N_17794,N_17733);
or U17872 (N_17872,N_17608,N_17655);
and U17873 (N_17873,N_17607,N_17746);
nor U17874 (N_17874,N_17690,N_17795);
nor U17875 (N_17875,N_17636,N_17773);
nor U17876 (N_17876,N_17641,N_17786);
or U17877 (N_17877,N_17770,N_17634);
xnor U17878 (N_17878,N_17645,N_17788);
xor U17879 (N_17879,N_17613,N_17713);
or U17880 (N_17880,N_17683,N_17727);
and U17881 (N_17881,N_17665,N_17710);
nor U17882 (N_17882,N_17685,N_17662);
and U17883 (N_17883,N_17789,N_17735);
xnor U17884 (N_17884,N_17672,N_17761);
nor U17885 (N_17885,N_17625,N_17760);
nand U17886 (N_17886,N_17646,N_17751);
or U17887 (N_17887,N_17745,N_17762);
and U17888 (N_17888,N_17724,N_17663);
nor U17889 (N_17889,N_17666,N_17749);
nor U17890 (N_17890,N_17692,N_17707);
xnor U17891 (N_17891,N_17763,N_17680);
and U17892 (N_17892,N_17799,N_17619);
nor U17893 (N_17893,N_17798,N_17784);
or U17894 (N_17894,N_17787,N_17790);
or U17895 (N_17895,N_17732,N_17677);
nand U17896 (N_17896,N_17699,N_17702);
nor U17897 (N_17897,N_17739,N_17743);
and U17898 (N_17898,N_17726,N_17633);
nor U17899 (N_17899,N_17720,N_17755);
nand U17900 (N_17900,N_17715,N_17700);
or U17901 (N_17901,N_17733,N_17611);
nor U17902 (N_17902,N_17787,N_17621);
nand U17903 (N_17903,N_17709,N_17757);
or U17904 (N_17904,N_17660,N_17642);
or U17905 (N_17905,N_17769,N_17630);
nor U17906 (N_17906,N_17727,N_17716);
or U17907 (N_17907,N_17698,N_17712);
or U17908 (N_17908,N_17783,N_17620);
xor U17909 (N_17909,N_17650,N_17661);
xor U17910 (N_17910,N_17738,N_17789);
or U17911 (N_17911,N_17609,N_17679);
or U17912 (N_17912,N_17743,N_17648);
nand U17913 (N_17913,N_17680,N_17720);
xor U17914 (N_17914,N_17687,N_17713);
nor U17915 (N_17915,N_17681,N_17725);
nor U17916 (N_17916,N_17681,N_17621);
nor U17917 (N_17917,N_17623,N_17769);
nor U17918 (N_17918,N_17688,N_17632);
xnor U17919 (N_17919,N_17690,N_17695);
nor U17920 (N_17920,N_17788,N_17652);
nand U17921 (N_17921,N_17612,N_17713);
and U17922 (N_17922,N_17613,N_17666);
and U17923 (N_17923,N_17617,N_17728);
xnor U17924 (N_17924,N_17721,N_17629);
or U17925 (N_17925,N_17710,N_17733);
xnor U17926 (N_17926,N_17738,N_17700);
xnor U17927 (N_17927,N_17637,N_17703);
xnor U17928 (N_17928,N_17783,N_17674);
nor U17929 (N_17929,N_17715,N_17795);
nand U17930 (N_17930,N_17715,N_17638);
nand U17931 (N_17931,N_17724,N_17767);
nand U17932 (N_17932,N_17797,N_17667);
or U17933 (N_17933,N_17638,N_17772);
or U17934 (N_17934,N_17684,N_17743);
nor U17935 (N_17935,N_17631,N_17638);
nand U17936 (N_17936,N_17607,N_17764);
xor U17937 (N_17937,N_17650,N_17630);
nor U17938 (N_17938,N_17637,N_17613);
xor U17939 (N_17939,N_17784,N_17686);
and U17940 (N_17940,N_17670,N_17677);
nand U17941 (N_17941,N_17751,N_17672);
nor U17942 (N_17942,N_17721,N_17604);
or U17943 (N_17943,N_17622,N_17668);
xnor U17944 (N_17944,N_17725,N_17754);
or U17945 (N_17945,N_17671,N_17644);
or U17946 (N_17946,N_17680,N_17664);
nand U17947 (N_17947,N_17728,N_17688);
or U17948 (N_17948,N_17659,N_17710);
or U17949 (N_17949,N_17778,N_17675);
nand U17950 (N_17950,N_17769,N_17771);
xor U17951 (N_17951,N_17628,N_17742);
nor U17952 (N_17952,N_17681,N_17693);
nor U17953 (N_17953,N_17647,N_17732);
or U17954 (N_17954,N_17607,N_17751);
nor U17955 (N_17955,N_17614,N_17624);
xnor U17956 (N_17956,N_17620,N_17688);
and U17957 (N_17957,N_17636,N_17654);
nor U17958 (N_17958,N_17718,N_17681);
nand U17959 (N_17959,N_17761,N_17676);
xnor U17960 (N_17960,N_17606,N_17705);
xor U17961 (N_17961,N_17756,N_17633);
or U17962 (N_17962,N_17641,N_17705);
xnor U17963 (N_17963,N_17752,N_17658);
nand U17964 (N_17964,N_17638,N_17786);
xnor U17965 (N_17965,N_17773,N_17741);
and U17966 (N_17966,N_17621,N_17667);
xor U17967 (N_17967,N_17607,N_17693);
nand U17968 (N_17968,N_17743,N_17722);
xor U17969 (N_17969,N_17777,N_17796);
nand U17970 (N_17970,N_17778,N_17792);
nor U17971 (N_17971,N_17685,N_17675);
nor U17972 (N_17972,N_17723,N_17667);
nand U17973 (N_17973,N_17739,N_17746);
nand U17974 (N_17974,N_17641,N_17719);
nand U17975 (N_17975,N_17782,N_17691);
xnor U17976 (N_17976,N_17612,N_17608);
nand U17977 (N_17977,N_17679,N_17715);
xnor U17978 (N_17978,N_17696,N_17718);
nor U17979 (N_17979,N_17664,N_17699);
xor U17980 (N_17980,N_17678,N_17749);
nor U17981 (N_17981,N_17640,N_17775);
nand U17982 (N_17982,N_17763,N_17725);
and U17983 (N_17983,N_17609,N_17783);
nand U17984 (N_17984,N_17721,N_17684);
xnor U17985 (N_17985,N_17794,N_17729);
and U17986 (N_17986,N_17615,N_17656);
or U17987 (N_17987,N_17618,N_17710);
and U17988 (N_17988,N_17769,N_17775);
xnor U17989 (N_17989,N_17705,N_17622);
and U17990 (N_17990,N_17641,N_17608);
nor U17991 (N_17991,N_17614,N_17670);
nor U17992 (N_17992,N_17608,N_17616);
xnor U17993 (N_17993,N_17784,N_17682);
and U17994 (N_17994,N_17659,N_17767);
and U17995 (N_17995,N_17701,N_17640);
nor U17996 (N_17996,N_17685,N_17621);
xnor U17997 (N_17997,N_17603,N_17681);
and U17998 (N_17998,N_17639,N_17668);
or U17999 (N_17999,N_17638,N_17778);
or U18000 (N_18000,N_17863,N_17821);
nand U18001 (N_18001,N_17910,N_17842);
nor U18002 (N_18002,N_17894,N_17960);
nand U18003 (N_18003,N_17984,N_17986);
and U18004 (N_18004,N_17869,N_17962);
xnor U18005 (N_18005,N_17889,N_17811);
nand U18006 (N_18006,N_17857,N_17921);
and U18007 (N_18007,N_17911,N_17899);
xnor U18008 (N_18008,N_17951,N_17848);
nor U18009 (N_18009,N_17812,N_17939);
xor U18010 (N_18010,N_17994,N_17856);
nor U18011 (N_18011,N_17950,N_17844);
nand U18012 (N_18012,N_17928,N_17849);
and U18013 (N_18013,N_17886,N_17909);
and U18014 (N_18014,N_17813,N_17904);
nand U18015 (N_18015,N_17829,N_17888);
xor U18016 (N_18016,N_17968,N_17961);
nor U18017 (N_18017,N_17884,N_17837);
xnor U18018 (N_18018,N_17808,N_17882);
or U18019 (N_18019,N_17998,N_17891);
xor U18020 (N_18020,N_17864,N_17877);
nor U18021 (N_18021,N_17918,N_17847);
nand U18022 (N_18022,N_17955,N_17983);
xor U18023 (N_18023,N_17903,N_17875);
or U18024 (N_18024,N_17896,N_17982);
xnor U18025 (N_18025,N_17971,N_17820);
nand U18026 (N_18026,N_17803,N_17947);
nand U18027 (N_18027,N_17948,N_17809);
or U18028 (N_18028,N_17810,N_17956);
or U18029 (N_18029,N_17926,N_17940);
nor U18030 (N_18030,N_17807,N_17925);
xor U18031 (N_18031,N_17854,N_17945);
xor U18032 (N_18032,N_17908,N_17852);
nand U18033 (N_18033,N_17885,N_17816);
nor U18034 (N_18034,N_17938,N_17805);
nand U18035 (N_18035,N_17929,N_17941);
or U18036 (N_18036,N_17953,N_17907);
xnor U18037 (N_18037,N_17978,N_17912);
nand U18038 (N_18038,N_17972,N_17963);
and U18039 (N_18039,N_17976,N_17828);
nand U18040 (N_18040,N_17826,N_17917);
nor U18041 (N_18041,N_17817,N_17897);
nor U18042 (N_18042,N_17834,N_17924);
xor U18043 (N_18043,N_17952,N_17946);
nor U18044 (N_18044,N_17870,N_17898);
xor U18045 (N_18045,N_17943,N_17937);
or U18046 (N_18046,N_17914,N_17954);
xor U18047 (N_18047,N_17977,N_17999);
or U18048 (N_18048,N_17985,N_17900);
and U18049 (N_18049,N_17964,N_17873);
nor U18050 (N_18050,N_17927,N_17892);
and U18051 (N_18051,N_17975,N_17804);
nand U18052 (N_18052,N_17931,N_17836);
or U18053 (N_18053,N_17843,N_17930);
nor U18054 (N_18054,N_17922,N_17936);
and U18055 (N_18055,N_17887,N_17860);
xnor U18056 (N_18056,N_17989,N_17965);
nor U18057 (N_18057,N_17916,N_17827);
xnor U18058 (N_18058,N_17851,N_17823);
or U18059 (N_18059,N_17876,N_17967);
nand U18060 (N_18060,N_17872,N_17979);
xor U18061 (N_18061,N_17833,N_17988);
nor U18062 (N_18062,N_17981,N_17919);
and U18063 (N_18063,N_17880,N_17881);
or U18064 (N_18064,N_17966,N_17987);
xnor U18065 (N_18065,N_17831,N_17825);
xnor U18066 (N_18066,N_17934,N_17871);
or U18067 (N_18067,N_17932,N_17846);
xor U18068 (N_18068,N_17902,N_17832);
nand U18069 (N_18069,N_17895,N_17942);
and U18070 (N_18070,N_17997,N_17862);
nor U18071 (N_18071,N_17815,N_17801);
nor U18072 (N_18072,N_17970,N_17993);
or U18073 (N_18073,N_17915,N_17830);
or U18074 (N_18074,N_17806,N_17850);
and U18075 (N_18075,N_17890,N_17974);
nand U18076 (N_18076,N_17845,N_17883);
nand U18077 (N_18077,N_17969,N_17992);
or U18078 (N_18078,N_17861,N_17944);
or U18079 (N_18079,N_17995,N_17841);
xor U18080 (N_18080,N_17822,N_17959);
nor U18081 (N_18081,N_17980,N_17853);
or U18082 (N_18082,N_17865,N_17866);
or U18083 (N_18083,N_17905,N_17835);
and U18084 (N_18084,N_17859,N_17858);
nand U18085 (N_18085,N_17893,N_17906);
nor U18086 (N_18086,N_17991,N_17824);
nand U18087 (N_18087,N_17838,N_17878);
xor U18088 (N_18088,N_17935,N_17990);
or U18089 (N_18089,N_17933,N_17949);
nor U18090 (N_18090,N_17913,N_17920);
nand U18091 (N_18091,N_17839,N_17819);
or U18092 (N_18092,N_17800,N_17923);
and U18093 (N_18093,N_17868,N_17840);
nor U18094 (N_18094,N_17901,N_17855);
xnor U18095 (N_18095,N_17814,N_17818);
or U18096 (N_18096,N_17996,N_17958);
or U18097 (N_18097,N_17973,N_17879);
or U18098 (N_18098,N_17802,N_17874);
or U18099 (N_18099,N_17867,N_17957);
nor U18100 (N_18100,N_17841,N_17896);
or U18101 (N_18101,N_17874,N_17808);
nor U18102 (N_18102,N_17921,N_17813);
or U18103 (N_18103,N_17908,N_17869);
nand U18104 (N_18104,N_17827,N_17848);
nand U18105 (N_18105,N_17908,N_17820);
or U18106 (N_18106,N_17822,N_17839);
and U18107 (N_18107,N_17991,N_17878);
nand U18108 (N_18108,N_17993,N_17918);
nand U18109 (N_18109,N_17814,N_17934);
nor U18110 (N_18110,N_17921,N_17917);
nand U18111 (N_18111,N_17923,N_17946);
nand U18112 (N_18112,N_17911,N_17955);
nor U18113 (N_18113,N_17873,N_17978);
nand U18114 (N_18114,N_17856,N_17887);
nor U18115 (N_18115,N_17810,N_17841);
nor U18116 (N_18116,N_17950,N_17963);
nor U18117 (N_18117,N_17947,N_17876);
and U18118 (N_18118,N_17803,N_17913);
nand U18119 (N_18119,N_17877,N_17951);
and U18120 (N_18120,N_17991,N_17915);
nand U18121 (N_18121,N_17904,N_17888);
or U18122 (N_18122,N_17972,N_17825);
nand U18123 (N_18123,N_17847,N_17842);
and U18124 (N_18124,N_17976,N_17950);
or U18125 (N_18125,N_17984,N_17807);
and U18126 (N_18126,N_17948,N_17912);
nand U18127 (N_18127,N_17863,N_17908);
or U18128 (N_18128,N_17801,N_17959);
xor U18129 (N_18129,N_17834,N_17837);
or U18130 (N_18130,N_17844,N_17887);
nand U18131 (N_18131,N_17972,N_17863);
nor U18132 (N_18132,N_17937,N_17963);
nand U18133 (N_18133,N_17844,N_17929);
nor U18134 (N_18134,N_17982,N_17842);
xnor U18135 (N_18135,N_17817,N_17824);
or U18136 (N_18136,N_17876,N_17950);
nor U18137 (N_18137,N_17828,N_17953);
and U18138 (N_18138,N_17906,N_17857);
xnor U18139 (N_18139,N_17916,N_17853);
nand U18140 (N_18140,N_17998,N_17867);
nor U18141 (N_18141,N_17835,N_17963);
nor U18142 (N_18142,N_17871,N_17979);
and U18143 (N_18143,N_17801,N_17927);
nor U18144 (N_18144,N_17810,N_17940);
nor U18145 (N_18145,N_17836,N_17919);
nand U18146 (N_18146,N_17932,N_17861);
or U18147 (N_18147,N_17965,N_17893);
and U18148 (N_18148,N_17916,N_17850);
or U18149 (N_18149,N_17810,N_17947);
nand U18150 (N_18150,N_17847,N_17923);
xnor U18151 (N_18151,N_17875,N_17890);
and U18152 (N_18152,N_17856,N_17884);
xnor U18153 (N_18153,N_17881,N_17910);
nand U18154 (N_18154,N_17962,N_17845);
nand U18155 (N_18155,N_17897,N_17862);
and U18156 (N_18156,N_17922,N_17886);
and U18157 (N_18157,N_17978,N_17871);
or U18158 (N_18158,N_17823,N_17894);
nor U18159 (N_18159,N_17907,N_17961);
nor U18160 (N_18160,N_17863,N_17852);
nor U18161 (N_18161,N_17942,N_17976);
xor U18162 (N_18162,N_17876,N_17847);
or U18163 (N_18163,N_17954,N_17823);
nand U18164 (N_18164,N_17967,N_17846);
nand U18165 (N_18165,N_17970,N_17871);
nor U18166 (N_18166,N_17887,N_17922);
or U18167 (N_18167,N_17932,N_17999);
xnor U18168 (N_18168,N_17937,N_17926);
and U18169 (N_18169,N_17974,N_17897);
nand U18170 (N_18170,N_17976,N_17915);
nor U18171 (N_18171,N_17808,N_17988);
nor U18172 (N_18172,N_17881,N_17844);
and U18173 (N_18173,N_17866,N_17847);
nor U18174 (N_18174,N_17990,N_17962);
nand U18175 (N_18175,N_17801,N_17973);
nand U18176 (N_18176,N_17833,N_17970);
or U18177 (N_18177,N_17896,N_17807);
nor U18178 (N_18178,N_17982,N_17989);
xor U18179 (N_18179,N_17928,N_17829);
nor U18180 (N_18180,N_17843,N_17826);
and U18181 (N_18181,N_17806,N_17966);
nand U18182 (N_18182,N_17823,N_17914);
and U18183 (N_18183,N_17908,N_17975);
nor U18184 (N_18184,N_17891,N_17900);
xnor U18185 (N_18185,N_17979,N_17853);
and U18186 (N_18186,N_17870,N_17955);
nor U18187 (N_18187,N_17975,N_17993);
xnor U18188 (N_18188,N_17908,N_17946);
or U18189 (N_18189,N_17954,N_17934);
or U18190 (N_18190,N_17815,N_17990);
or U18191 (N_18191,N_17930,N_17942);
xor U18192 (N_18192,N_17850,N_17995);
xnor U18193 (N_18193,N_17858,N_17991);
xnor U18194 (N_18194,N_17956,N_17840);
nor U18195 (N_18195,N_17986,N_17969);
and U18196 (N_18196,N_17883,N_17825);
nand U18197 (N_18197,N_17808,N_17913);
nand U18198 (N_18198,N_17807,N_17880);
or U18199 (N_18199,N_17953,N_17813);
or U18200 (N_18200,N_18146,N_18129);
or U18201 (N_18201,N_18157,N_18030);
nor U18202 (N_18202,N_18118,N_18028);
or U18203 (N_18203,N_18098,N_18102);
or U18204 (N_18204,N_18005,N_18168);
nor U18205 (N_18205,N_18127,N_18064);
or U18206 (N_18206,N_18128,N_18160);
nand U18207 (N_18207,N_18023,N_18036);
xnor U18208 (N_18208,N_18143,N_18070);
nand U18209 (N_18209,N_18130,N_18039);
nor U18210 (N_18210,N_18014,N_18029);
and U18211 (N_18211,N_18046,N_18117);
or U18212 (N_18212,N_18096,N_18162);
and U18213 (N_18213,N_18188,N_18078);
and U18214 (N_18214,N_18182,N_18183);
and U18215 (N_18215,N_18038,N_18075);
and U18216 (N_18216,N_18055,N_18185);
nand U18217 (N_18217,N_18139,N_18024);
nor U18218 (N_18218,N_18158,N_18174);
xnor U18219 (N_18219,N_18135,N_18093);
nor U18220 (N_18220,N_18044,N_18140);
or U18221 (N_18221,N_18145,N_18058);
nor U18222 (N_18222,N_18103,N_18091);
or U18223 (N_18223,N_18152,N_18155);
or U18224 (N_18224,N_18047,N_18032);
nor U18225 (N_18225,N_18089,N_18006);
or U18226 (N_18226,N_18052,N_18010);
or U18227 (N_18227,N_18149,N_18009);
nor U18228 (N_18228,N_18177,N_18186);
and U18229 (N_18229,N_18119,N_18048);
nand U18230 (N_18230,N_18147,N_18124);
and U18231 (N_18231,N_18088,N_18082);
and U18232 (N_18232,N_18144,N_18167);
and U18233 (N_18233,N_18198,N_18085);
nor U18234 (N_18234,N_18132,N_18106);
nand U18235 (N_18235,N_18173,N_18115);
and U18236 (N_18236,N_18042,N_18081);
xor U18237 (N_18237,N_18138,N_18123);
xor U18238 (N_18238,N_18142,N_18056);
and U18239 (N_18239,N_18192,N_18193);
and U18240 (N_18240,N_18086,N_18134);
nor U18241 (N_18241,N_18136,N_18197);
nor U18242 (N_18242,N_18092,N_18045);
nor U18243 (N_18243,N_18073,N_18033);
nor U18244 (N_18244,N_18074,N_18060);
xor U18245 (N_18245,N_18097,N_18004);
xor U18246 (N_18246,N_18002,N_18170);
or U18247 (N_18247,N_18012,N_18001);
xnor U18248 (N_18248,N_18099,N_18189);
or U18249 (N_18249,N_18020,N_18125);
xnor U18250 (N_18250,N_18062,N_18007);
nor U18251 (N_18251,N_18069,N_18126);
or U18252 (N_18252,N_18133,N_18013);
xnor U18253 (N_18253,N_18026,N_18066);
nand U18254 (N_18254,N_18008,N_18034);
and U18255 (N_18255,N_18151,N_18153);
nand U18256 (N_18256,N_18181,N_18179);
nand U18257 (N_18257,N_18003,N_18101);
xnor U18258 (N_18258,N_18111,N_18022);
or U18259 (N_18259,N_18037,N_18015);
xnor U18260 (N_18260,N_18080,N_18190);
or U18261 (N_18261,N_18159,N_18107);
nor U18262 (N_18262,N_18108,N_18172);
nand U18263 (N_18263,N_18011,N_18049);
and U18264 (N_18264,N_18137,N_18112);
or U18265 (N_18265,N_18027,N_18169);
or U18266 (N_18266,N_18072,N_18031);
or U18267 (N_18267,N_18154,N_18122);
or U18268 (N_18268,N_18063,N_18017);
nand U18269 (N_18269,N_18116,N_18150);
and U18270 (N_18270,N_18016,N_18121);
or U18271 (N_18271,N_18110,N_18051);
nor U18272 (N_18272,N_18071,N_18041);
xor U18273 (N_18273,N_18035,N_18065);
nor U18274 (N_18274,N_18161,N_18180);
or U18275 (N_18275,N_18131,N_18053);
and U18276 (N_18276,N_18067,N_18120);
and U18277 (N_18277,N_18148,N_18076);
xor U18278 (N_18278,N_18057,N_18090);
nand U18279 (N_18279,N_18019,N_18021);
nand U18280 (N_18280,N_18175,N_18084);
and U18281 (N_18281,N_18194,N_18100);
and U18282 (N_18282,N_18083,N_18050);
nor U18283 (N_18283,N_18077,N_18109);
and U18284 (N_18284,N_18195,N_18059);
xor U18285 (N_18285,N_18156,N_18165);
nand U18286 (N_18286,N_18163,N_18061);
and U18287 (N_18287,N_18025,N_18164);
and U18288 (N_18288,N_18054,N_18176);
or U18289 (N_18289,N_18196,N_18171);
xnor U18290 (N_18290,N_18191,N_18094);
nor U18291 (N_18291,N_18178,N_18104);
xnor U18292 (N_18292,N_18199,N_18018);
nand U18293 (N_18293,N_18105,N_18166);
and U18294 (N_18294,N_18114,N_18187);
xnor U18295 (N_18295,N_18087,N_18043);
xnor U18296 (N_18296,N_18040,N_18184);
nand U18297 (N_18297,N_18079,N_18068);
nand U18298 (N_18298,N_18000,N_18095);
nand U18299 (N_18299,N_18141,N_18113);
nor U18300 (N_18300,N_18110,N_18194);
and U18301 (N_18301,N_18177,N_18114);
nand U18302 (N_18302,N_18190,N_18116);
or U18303 (N_18303,N_18044,N_18118);
and U18304 (N_18304,N_18030,N_18155);
or U18305 (N_18305,N_18129,N_18126);
xnor U18306 (N_18306,N_18104,N_18036);
xor U18307 (N_18307,N_18078,N_18027);
nand U18308 (N_18308,N_18117,N_18012);
nand U18309 (N_18309,N_18124,N_18010);
and U18310 (N_18310,N_18126,N_18145);
or U18311 (N_18311,N_18133,N_18187);
xor U18312 (N_18312,N_18024,N_18010);
or U18313 (N_18313,N_18127,N_18136);
and U18314 (N_18314,N_18022,N_18156);
xnor U18315 (N_18315,N_18181,N_18145);
or U18316 (N_18316,N_18089,N_18192);
nor U18317 (N_18317,N_18065,N_18166);
and U18318 (N_18318,N_18175,N_18023);
nand U18319 (N_18319,N_18163,N_18083);
and U18320 (N_18320,N_18094,N_18070);
or U18321 (N_18321,N_18072,N_18197);
nand U18322 (N_18322,N_18082,N_18003);
and U18323 (N_18323,N_18013,N_18085);
nand U18324 (N_18324,N_18076,N_18119);
nand U18325 (N_18325,N_18089,N_18175);
nor U18326 (N_18326,N_18143,N_18062);
nand U18327 (N_18327,N_18099,N_18079);
nand U18328 (N_18328,N_18074,N_18036);
xor U18329 (N_18329,N_18143,N_18105);
nand U18330 (N_18330,N_18087,N_18144);
xnor U18331 (N_18331,N_18075,N_18077);
nand U18332 (N_18332,N_18087,N_18184);
or U18333 (N_18333,N_18066,N_18151);
nand U18334 (N_18334,N_18160,N_18148);
nand U18335 (N_18335,N_18128,N_18007);
xnor U18336 (N_18336,N_18199,N_18022);
or U18337 (N_18337,N_18008,N_18181);
nor U18338 (N_18338,N_18159,N_18016);
nand U18339 (N_18339,N_18079,N_18127);
xnor U18340 (N_18340,N_18035,N_18007);
or U18341 (N_18341,N_18034,N_18167);
nand U18342 (N_18342,N_18176,N_18127);
nor U18343 (N_18343,N_18086,N_18061);
or U18344 (N_18344,N_18192,N_18125);
or U18345 (N_18345,N_18172,N_18050);
or U18346 (N_18346,N_18120,N_18072);
or U18347 (N_18347,N_18184,N_18165);
and U18348 (N_18348,N_18036,N_18018);
nor U18349 (N_18349,N_18000,N_18131);
or U18350 (N_18350,N_18057,N_18052);
or U18351 (N_18351,N_18078,N_18064);
nand U18352 (N_18352,N_18160,N_18031);
or U18353 (N_18353,N_18166,N_18196);
xnor U18354 (N_18354,N_18097,N_18163);
and U18355 (N_18355,N_18141,N_18053);
or U18356 (N_18356,N_18132,N_18028);
nand U18357 (N_18357,N_18026,N_18044);
nor U18358 (N_18358,N_18096,N_18000);
nor U18359 (N_18359,N_18073,N_18172);
and U18360 (N_18360,N_18017,N_18072);
or U18361 (N_18361,N_18134,N_18026);
and U18362 (N_18362,N_18146,N_18112);
nand U18363 (N_18363,N_18159,N_18139);
nor U18364 (N_18364,N_18059,N_18058);
nor U18365 (N_18365,N_18140,N_18159);
or U18366 (N_18366,N_18171,N_18121);
and U18367 (N_18367,N_18125,N_18163);
nand U18368 (N_18368,N_18021,N_18109);
or U18369 (N_18369,N_18029,N_18107);
or U18370 (N_18370,N_18181,N_18185);
and U18371 (N_18371,N_18083,N_18033);
or U18372 (N_18372,N_18169,N_18152);
or U18373 (N_18373,N_18044,N_18149);
or U18374 (N_18374,N_18080,N_18036);
xor U18375 (N_18375,N_18199,N_18128);
and U18376 (N_18376,N_18152,N_18198);
and U18377 (N_18377,N_18161,N_18024);
nor U18378 (N_18378,N_18005,N_18127);
and U18379 (N_18379,N_18035,N_18068);
or U18380 (N_18380,N_18029,N_18088);
xor U18381 (N_18381,N_18003,N_18199);
or U18382 (N_18382,N_18034,N_18126);
or U18383 (N_18383,N_18189,N_18175);
nand U18384 (N_18384,N_18022,N_18061);
nand U18385 (N_18385,N_18190,N_18099);
and U18386 (N_18386,N_18129,N_18054);
nor U18387 (N_18387,N_18129,N_18177);
nand U18388 (N_18388,N_18014,N_18145);
and U18389 (N_18389,N_18016,N_18143);
and U18390 (N_18390,N_18158,N_18062);
xor U18391 (N_18391,N_18153,N_18055);
or U18392 (N_18392,N_18054,N_18007);
nand U18393 (N_18393,N_18039,N_18102);
xnor U18394 (N_18394,N_18015,N_18070);
nand U18395 (N_18395,N_18188,N_18051);
and U18396 (N_18396,N_18179,N_18166);
xnor U18397 (N_18397,N_18107,N_18146);
xnor U18398 (N_18398,N_18170,N_18000);
nor U18399 (N_18399,N_18175,N_18123);
nor U18400 (N_18400,N_18363,N_18264);
nor U18401 (N_18401,N_18327,N_18318);
or U18402 (N_18402,N_18307,N_18222);
xor U18403 (N_18403,N_18393,N_18238);
xnor U18404 (N_18404,N_18232,N_18287);
and U18405 (N_18405,N_18276,N_18252);
or U18406 (N_18406,N_18220,N_18314);
or U18407 (N_18407,N_18227,N_18371);
xor U18408 (N_18408,N_18369,N_18310);
xor U18409 (N_18409,N_18272,N_18376);
or U18410 (N_18410,N_18315,N_18263);
nor U18411 (N_18411,N_18253,N_18245);
and U18412 (N_18412,N_18381,N_18229);
and U18413 (N_18413,N_18350,N_18321);
and U18414 (N_18414,N_18281,N_18250);
and U18415 (N_18415,N_18390,N_18334);
or U18416 (N_18416,N_18361,N_18308);
nand U18417 (N_18417,N_18243,N_18246);
and U18418 (N_18418,N_18269,N_18370);
and U18419 (N_18419,N_18212,N_18348);
xnor U18420 (N_18420,N_18224,N_18251);
xnor U18421 (N_18421,N_18386,N_18219);
nand U18422 (N_18422,N_18274,N_18324);
xor U18423 (N_18423,N_18268,N_18210);
and U18424 (N_18424,N_18280,N_18313);
and U18425 (N_18425,N_18275,N_18207);
xnor U18426 (N_18426,N_18378,N_18312);
or U18427 (N_18427,N_18316,N_18328);
and U18428 (N_18428,N_18330,N_18325);
or U18429 (N_18429,N_18341,N_18225);
xnor U18430 (N_18430,N_18244,N_18297);
and U18431 (N_18431,N_18266,N_18217);
nor U18432 (N_18432,N_18296,N_18366);
or U18433 (N_18433,N_18346,N_18392);
nor U18434 (N_18434,N_18391,N_18396);
xnor U18435 (N_18435,N_18382,N_18367);
or U18436 (N_18436,N_18323,N_18206);
xnor U18437 (N_18437,N_18331,N_18213);
or U18438 (N_18438,N_18344,N_18298);
or U18439 (N_18439,N_18231,N_18306);
nor U18440 (N_18440,N_18211,N_18322);
or U18441 (N_18441,N_18230,N_18291);
xnor U18442 (N_18442,N_18236,N_18277);
and U18443 (N_18443,N_18387,N_18290);
and U18444 (N_18444,N_18205,N_18248);
and U18445 (N_18445,N_18258,N_18304);
nor U18446 (N_18446,N_18289,N_18311);
xor U18447 (N_18447,N_18240,N_18309);
nand U18448 (N_18448,N_18265,N_18254);
nand U18449 (N_18449,N_18388,N_18237);
nand U18450 (N_18450,N_18302,N_18273);
xor U18451 (N_18451,N_18215,N_18288);
and U18452 (N_18452,N_18226,N_18295);
xnor U18453 (N_18453,N_18345,N_18299);
xor U18454 (N_18454,N_18365,N_18214);
xnor U18455 (N_18455,N_18383,N_18200);
xor U18456 (N_18456,N_18317,N_18239);
nand U18457 (N_18457,N_18270,N_18209);
nor U18458 (N_18458,N_18249,N_18373);
and U18459 (N_18459,N_18357,N_18358);
xnor U18460 (N_18460,N_18362,N_18257);
nand U18461 (N_18461,N_18300,N_18329);
xor U18462 (N_18462,N_18359,N_18292);
nand U18463 (N_18463,N_18336,N_18395);
or U18464 (N_18464,N_18377,N_18216);
nand U18465 (N_18465,N_18305,N_18398);
and U18466 (N_18466,N_18221,N_18279);
or U18467 (N_18467,N_18202,N_18352);
nand U18468 (N_18468,N_18389,N_18267);
or U18469 (N_18469,N_18260,N_18333);
nand U18470 (N_18470,N_18354,N_18301);
xor U18471 (N_18471,N_18203,N_18338);
or U18472 (N_18472,N_18343,N_18241);
and U18473 (N_18473,N_18271,N_18326);
or U18474 (N_18474,N_18286,N_18247);
xnor U18475 (N_18475,N_18351,N_18394);
nor U18476 (N_18476,N_18355,N_18397);
nand U18477 (N_18477,N_18278,N_18375);
xnor U18478 (N_18478,N_18261,N_18259);
nor U18479 (N_18479,N_18335,N_18204);
nand U18480 (N_18480,N_18340,N_18360);
xor U18481 (N_18481,N_18235,N_18201);
or U18482 (N_18482,N_18208,N_18342);
xor U18483 (N_18483,N_18282,N_18255);
and U18484 (N_18484,N_18399,N_18349);
and U18485 (N_18485,N_18339,N_18337);
xnor U18486 (N_18486,N_18293,N_18223);
and U18487 (N_18487,N_18303,N_18233);
xnor U18488 (N_18488,N_18228,N_18374);
nor U18489 (N_18489,N_18256,N_18379);
and U18490 (N_18490,N_18262,N_18319);
xor U18491 (N_18491,N_18384,N_18285);
nand U18492 (N_18492,N_18294,N_18372);
or U18493 (N_18493,N_18347,N_18218);
and U18494 (N_18494,N_18284,N_18234);
nand U18495 (N_18495,N_18283,N_18385);
or U18496 (N_18496,N_18320,N_18368);
nor U18497 (N_18497,N_18332,N_18353);
or U18498 (N_18498,N_18356,N_18380);
nor U18499 (N_18499,N_18242,N_18364);
nand U18500 (N_18500,N_18367,N_18309);
or U18501 (N_18501,N_18304,N_18265);
xnor U18502 (N_18502,N_18383,N_18375);
nor U18503 (N_18503,N_18292,N_18352);
xnor U18504 (N_18504,N_18210,N_18238);
nor U18505 (N_18505,N_18325,N_18392);
nor U18506 (N_18506,N_18274,N_18322);
nand U18507 (N_18507,N_18317,N_18338);
nand U18508 (N_18508,N_18280,N_18386);
or U18509 (N_18509,N_18246,N_18210);
nor U18510 (N_18510,N_18364,N_18266);
or U18511 (N_18511,N_18334,N_18344);
nor U18512 (N_18512,N_18279,N_18208);
nor U18513 (N_18513,N_18220,N_18276);
and U18514 (N_18514,N_18330,N_18371);
and U18515 (N_18515,N_18352,N_18256);
xnor U18516 (N_18516,N_18241,N_18355);
and U18517 (N_18517,N_18228,N_18217);
nand U18518 (N_18518,N_18267,N_18273);
nand U18519 (N_18519,N_18371,N_18269);
nand U18520 (N_18520,N_18305,N_18235);
or U18521 (N_18521,N_18364,N_18346);
and U18522 (N_18522,N_18207,N_18267);
or U18523 (N_18523,N_18248,N_18331);
or U18524 (N_18524,N_18298,N_18266);
xor U18525 (N_18525,N_18361,N_18397);
or U18526 (N_18526,N_18307,N_18211);
nor U18527 (N_18527,N_18242,N_18283);
xnor U18528 (N_18528,N_18325,N_18275);
or U18529 (N_18529,N_18381,N_18382);
and U18530 (N_18530,N_18217,N_18308);
nor U18531 (N_18531,N_18316,N_18322);
nor U18532 (N_18532,N_18259,N_18227);
or U18533 (N_18533,N_18215,N_18213);
or U18534 (N_18534,N_18387,N_18234);
xnor U18535 (N_18535,N_18349,N_18317);
nand U18536 (N_18536,N_18286,N_18380);
xnor U18537 (N_18537,N_18348,N_18235);
nor U18538 (N_18538,N_18328,N_18344);
xnor U18539 (N_18539,N_18315,N_18203);
nor U18540 (N_18540,N_18335,N_18322);
and U18541 (N_18541,N_18303,N_18284);
and U18542 (N_18542,N_18398,N_18219);
nand U18543 (N_18543,N_18234,N_18230);
and U18544 (N_18544,N_18244,N_18368);
or U18545 (N_18545,N_18347,N_18385);
xnor U18546 (N_18546,N_18347,N_18374);
or U18547 (N_18547,N_18215,N_18308);
nor U18548 (N_18548,N_18331,N_18307);
nor U18549 (N_18549,N_18337,N_18241);
and U18550 (N_18550,N_18310,N_18243);
nor U18551 (N_18551,N_18260,N_18254);
and U18552 (N_18552,N_18314,N_18384);
or U18553 (N_18553,N_18318,N_18309);
xnor U18554 (N_18554,N_18203,N_18207);
nand U18555 (N_18555,N_18246,N_18363);
or U18556 (N_18556,N_18345,N_18373);
xor U18557 (N_18557,N_18397,N_18247);
nand U18558 (N_18558,N_18397,N_18296);
nand U18559 (N_18559,N_18373,N_18321);
nor U18560 (N_18560,N_18245,N_18363);
xor U18561 (N_18561,N_18366,N_18363);
nor U18562 (N_18562,N_18299,N_18373);
or U18563 (N_18563,N_18257,N_18297);
nor U18564 (N_18564,N_18377,N_18345);
nand U18565 (N_18565,N_18344,N_18256);
xnor U18566 (N_18566,N_18277,N_18353);
nand U18567 (N_18567,N_18386,N_18354);
nand U18568 (N_18568,N_18329,N_18243);
and U18569 (N_18569,N_18387,N_18339);
nand U18570 (N_18570,N_18270,N_18306);
nor U18571 (N_18571,N_18337,N_18218);
and U18572 (N_18572,N_18359,N_18289);
and U18573 (N_18573,N_18393,N_18364);
and U18574 (N_18574,N_18291,N_18312);
xnor U18575 (N_18575,N_18291,N_18260);
nand U18576 (N_18576,N_18396,N_18367);
xor U18577 (N_18577,N_18230,N_18288);
and U18578 (N_18578,N_18265,N_18283);
or U18579 (N_18579,N_18323,N_18223);
xnor U18580 (N_18580,N_18221,N_18213);
nor U18581 (N_18581,N_18299,N_18320);
or U18582 (N_18582,N_18244,N_18286);
nand U18583 (N_18583,N_18254,N_18225);
and U18584 (N_18584,N_18264,N_18370);
nor U18585 (N_18585,N_18267,N_18363);
and U18586 (N_18586,N_18211,N_18342);
and U18587 (N_18587,N_18347,N_18291);
xnor U18588 (N_18588,N_18339,N_18203);
and U18589 (N_18589,N_18304,N_18395);
xnor U18590 (N_18590,N_18345,N_18336);
or U18591 (N_18591,N_18348,N_18243);
nor U18592 (N_18592,N_18388,N_18205);
xnor U18593 (N_18593,N_18378,N_18264);
nor U18594 (N_18594,N_18322,N_18229);
or U18595 (N_18595,N_18252,N_18272);
and U18596 (N_18596,N_18310,N_18256);
and U18597 (N_18597,N_18242,N_18333);
and U18598 (N_18598,N_18219,N_18233);
nand U18599 (N_18599,N_18338,N_18314);
nor U18600 (N_18600,N_18543,N_18456);
nand U18601 (N_18601,N_18493,N_18558);
or U18602 (N_18602,N_18473,N_18494);
xnor U18603 (N_18603,N_18461,N_18564);
and U18604 (N_18604,N_18414,N_18472);
xor U18605 (N_18605,N_18512,N_18492);
nor U18606 (N_18606,N_18572,N_18406);
xor U18607 (N_18607,N_18412,N_18486);
nand U18608 (N_18608,N_18415,N_18591);
nor U18609 (N_18609,N_18556,N_18560);
or U18610 (N_18610,N_18573,N_18477);
nand U18611 (N_18611,N_18580,N_18554);
nor U18612 (N_18612,N_18459,N_18559);
nand U18613 (N_18613,N_18531,N_18557);
nor U18614 (N_18614,N_18429,N_18498);
xor U18615 (N_18615,N_18575,N_18444);
nand U18616 (N_18616,N_18588,N_18402);
nand U18617 (N_18617,N_18578,N_18535);
and U18618 (N_18618,N_18469,N_18586);
or U18619 (N_18619,N_18446,N_18458);
nand U18620 (N_18620,N_18421,N_18448);
xor U18621 (N_18621,N_18404,N_18562);
or U18622 (N_18622,N_18519,N_18409);
or U18623 (N_18623,N_18481,N_18538);
nand U18624 (N_18624,N_18569,N_18540);
and U18625 (N_18625,N_18521,N_18438);
or U18626 (N_18626,N_18565,N_18434);
nand U18627 (N_18627,N_18593,N_18435);
xnor U18628 (N_18628,N_18561,N_18507);
and U18629 (N_18629,N_18466,N_18515);
and U18630 (N_18630,N_18453,N_18550);
and U18631 (N_18631,N_18584,N_18528);
and U18632 (N_18632,N_18529,N_18503);
or U18633 (N_18633,N_18518,N_18549);
nor U18634 (N_18634,N_18483,N_18442);
nand U18635 (N_18635,N_18548,N_18506);
or U18636 (N_18636,N_18451,N_18596);
xor U18637 (N_18637,N_18537,N_18581);
or U18638 (N_18638,N_18422,N_18430);
nor U18639 (N_18639,N_18460,N_18485);
or U18640 (N_18640,N_18418,N_18502);
and U18641 (N_18641,N_18497,N_18536);
and U18642 (N_18642,N_18568,N_18504);
nand U18643 (N_18643,N_18416,N_18525);
xnor U18644 (N_18644,N_18488,N_18545);
nand U18645 (N_18645,N_18441,N_18479);
nor U18646 (N_18646,N_18455,N_18595);
or U18647 (N_18647,N_18501,N_18583);
xnor U18648 (N_18648,N_18594,N_18571);
nor U18649 (N_18649,N_18547,N_18495);
nor U18650 (N_18650,N_18433,N_18457);
nor U18651 (N_18651,N_18410,N_18443);
nand U18652 (N_18652,N_18424,N_18514);
xnor U18653 (N_18653,N_18475,N_18567);
or U18654 (N_18654,N_18474,N_18432);
nand U18655 (N_18655,N_18577,N_18464);
nand U18656 (N_18656,N_18419,N_18417);
nand U18657 (N_18657,N_18534,N_18449);
or U18658 (N_18658,N_18478,N_18517);
and U18659 (N_18659,N_18511,N_18582);
nor U18660 (N_18660,N_18484,N_18425);
nand U18661 (N_18661,N_18516,N_18403);
and U18662 (N_18662,N_18445,N_18551);
nand U18663 (N_18663,N_18522,N_18462);
xnor U18664 (N_18664,N_18589,N_18599);
nor U18665 (N_18665,N_18541,N_18463);
and U18666 (N_18666,N_18482,N_18408);
nand U18667 (N_18667,N_18590,N_18597);
and U18668 (N_18668,N_18407,N_18454);
or U18669 (N_18669,N_18546,N_18440);
nor U18670 (N_18670,N_18489,N_18539);
nor U18671 (N_18671,N_18476,N_18527);
nor U18672 (N_18672,N_18552,N_18523);
or U18673 (N_18673,N_18431,N_18420);
nand U18674 (N_18674,N_18426,N_18470);
and U18675 (N_18675,N_18505,N_18563);
and U18676 (N_18676,N_18437,N_18592);
nand U18677 (N_18677,N_18530,N_18465);
nor U18678 (N_18678,N_18500,N_18579);
and U18679 (N_18679,N_18428,N_18439);
or U18680 (N_18680,N_18544,N_18587);
or U18681 (N_18681,N_18487,N_18405);
and U18682 (N_18682,N_18598,N_18496);
nand U18683 (N_18683,N_18400,N_18452);
or U18684 (N_18684,N_18468,N_18526);
or U18685 (N_18685,N_18533,N_18427);
xor U18686 (N_18686,N_18423,N_18411);
or U18687 (N_18687,N_18524,N_18520);
and U18688 (N_18688,N_18447,N_18574);
nor U18689 (N_18689,N_18566,N_18436);
xnor U18690 (N_18690,N_18570,N_18471);
and U18691 (N_18691,N_18509,N_18480);
or U18692 (N_18692,N_18576,N_18450);
nor U18693 (N_18693,N_18542,N_18467);
xor U18694 (N_18694,N_18491,N_18585);
or U18695 (N_18695,N_18513,N_18401);
or U18696 (N_18696,N_18490,N_18532);
and U18697 (N_18697,N_18555,N_18508);
nand U18698 (N_18698,N_18413,N_18510);
and U18699 (N_18699,N_18499,N_18553);
xor U18700 (N_18700,N_18557,N_18407);
xor U18701 (N_18701,N_18582,N_18462);
or U18702 (N_18702,N_18441,N_18531);
nor U18703 (N_18703,N_18593,N_18563);
nor U18704 (N_18704,N_18599,N_18466);
xnor U18705 (N_18705,N_18442,N_18596);
and U18706 (N_18706,N_18540,N_18590);
xnor U18707 (N_18707,N_18467,N_18455);
nand U18708 (N_18708,N_18491,N_18440);
or U18709 (N_18709,N_18540,N_18465);
nand U18710 (N_18710,N_18506,N_18427);
nor U18711 (N_18711,N_18434,N_18517);
nor U18712 (N_18712,N_18491,N_18501);
or U18713 (N_18713,N_18420,N_18533);
nand U18714 (N_18714,N_18480,N_18599);
and U18715 (N_18715,N_18503,N_18515);
nor U18716 (N_18716,N_18462,N_18516);
or U18717 (N_18717,N_18437,N_18402);
nand U18718 (N_18718,N_18497,N_18461);
and U18719 (N_18719,N_18438,N_18462);
nand U18720 (N_18720,N_18570,N_18517);
or U18721 (N_18721,N_18599,N_18418);
nand U18722 (N_18722,N_18466,N_18429);
or U18723 (N_18723,N_18478,N_18599);
nor U18724 (N_18724,N_18567,N_18525);
nor U18725 (N_18725,N_18537,N_18499);
xor U18726 (N_18726,N_18421,N_18404);
nand U18727 (N_18727,N_18485,N_18449);
xnor U18728 (N_18728,N_18555,N_18459);
xnor U18729 (N_18729,N_18419,N_18444);
xnor U18730 (N_18730,N_18548,N_18462);
nor U18731 (N_18731,N_18533,N_18464);
and U18732 (N_18732,N_18495,N_18404);
or U18733 (N_18733,N_18573,N_18484);
xor U18734 (N_18734,N_18438,N_18560);
nand U18735 (N_18735,N_18539,N_18474);
or U18736 (N_18736,N_18443,N_18446);
nor U18737 (N_18737,N_18501,N_18474);
and U18738 (N_18738,N_18438,N_18593);
xnor U18739 (N_18739,N_18590,N_18519);
or U18740 (N_18740,N_18400,N_18435);
nor U18741 (N_18741,N_18469,N_18529);
nor U18742 (N_18742,N_18411,N_18589);
nor U18743 (N_18743,N_18555,N_18594);
nor U18744 (N_18744,N_18472,N_18418);
nand U18745 (N_18745,N_18508,N_18527);
or U18746 (N_18746,N_18453,N_18440);
nor U18747 (N_18747,N_18508,N_18452);
nand U18748 (N_18748,N_18425,N_18560);
nor U18749 (N_18749,N_18435,N_18562);
nor U18750 (N_18750,N_18416,N_18517);
or U18751 (N_18751,N_18565,N_18442);
nor U18752 (N_18752,N_18550,N_18591);
and U18753 (N_18753,N_18578,N_18539);
or U18754 (N_18754,N_18492,N_18455);
and U18755 (N_18755,N_18428,N_18440);
or U18756 (N_18756,N_18414,N_18464);
nand U18757 (N_18757,N_18595,N_18501);
nand U18758 (N_18758,N_18450,N_18570);
nor U18759 (N_18759,N_18570,N_18403);
and U18760 (N_18760,N_18567,N_18442);
nand U18761 (N_18761,N_18497,N_18425);
xor U18762 (N_18762,N_18513,N_18550);
nor U18763 (N_18763,N_18540,N_18534);
nand U18764 (N_18764,N_18542,N_18478);
or U18765 (N_18765,N_18416,N_18557);
or U18766 (N_18766,N_18403,N_18586);
nor U18767 (N_18767,N_18483,N_18486);
xnor U18768 (N_18768,N_18536,N_18494);
and U18769 (N_18769,N_18590,N_18412);
xnor U18770 (N_18770,N_18506,N_18416);
nor U18771 (N_18771,N_18469,N_18420);
xnor U18772 (N_18772,N_18441,N_18530);
and U18773 (N_18773,N_18597,N_18460);
nor U18774 (N_18774,N_18492,N_18441);
and U18775 (N_18775,N_18439,N_18450);
nor U18776 (N_18776,N_18570,N_18584);
or U18777 (N_18777,N_18571,N_18421);
and U18778 (N_18778,N_18465,N_18502);
nand U18779 (N_18779,N_18516,N_18460);
nand U18780 (N_18780,N_18429,N_18583);
or U18781 (N_18781,N_18496,N_18439);
nor U18782 (N_18782,N_18511,N_18430);
xnor U18783 (N_18783,N_18417,N_18445);
nor U18784 (N_18784,N_18506,N_18535);
nor U18785 (N_18785,N_18438,N_18474);
xnor U18786 (N_18786,N_18432,N_18492);
nor U18787 (N_18787,N_18531,N_18437);
nor U18788 (N_18788,N_18454,N_18537);
xor U18789 (N_18789,N_18487,N_18565);
or U18790 (N_18790,N_18421,N_18575);
and U18791 (N_18791,N_18506,N_18408);
nand U18792 (N_18792,N_18528,N_18482);
nor U18793 (N_18793,N_18489,N_18547);
and U18794 (N_18794,N_18527,N_18544);
or U18795 (N_18795,N_18477,N_18442);
nor U18796 (N_18796,N_18584,N_18408);
nor U18797 (N_18797,N_18453,N_18598);
xnor U18798 (N_18798,N_18434,N_18401);
xnor U18799 (N_18799,N_18579,N_18546);
or U18800 (N_18800,N_18603,N_18632);
xnor U18801 (N_18801,N_18738,N_18754);
nor U18802 (N_18802,N_18623,N_18732);
xnor U18803 (N_18803,N_18651,N_18712);
xor U18804 (N_18804,N_18766,N_18608);
or U18805 (N_18805,N_18745,N_18677);
nor U18806 (N_18806,N_18678,N_18740);
xnor U18807 (N_18807,N_18760,N_18767);
xor U18808 (N_18808,N_18601,N_18799);
or U18809 (N_18809,N_18641,N_18634);
nand U18810 (N_18810,N_18693,N_18646);
nor U18811 (N_18811,N_18764,N_18749);
or U18812 (N_18812,N_18727,N_18700);
xor U18813 (N_18813,N_18779,N_18705);
nand U18814 (N_18814,N_18728,N_18658);
nor U18815 (N_18815,N_18718,N_18605);
nor U18816 (N_18816,N_18751,N_18633);
and U18817 (N_18817,N_18798,N_18719);
xor U18818 (N_18818,N_18609,N_18723);
nand U18819 (N_18819,N_18682,N_18604);
nand U18820 (N_18820,N_18681,N_18781);
nand U18821 (N_18821,N_18787,N_18638);
nand U18822 (N_18822,N_18743,N_18716);
xnor U18823 (N_18823,N_18683,N_18611);
xnor U18824 (N_18824,N_18676,N_18769);
or U18825 (N_18825,N_18635,N_18748);
nor U18826 (N_18826,N_18672,N_18600);
and U18827 (N_18827,N_18697,N_18689);
nor U18828 (N_18828,N_18688,N_18667);
nand U18829 (N_18829,N_18765,N_18655);
xnor U18830 (N_18830,N_18675,N_18643);
nand U18831 (N_18831,N_18660,N_18742);
or U18832 (N_18832,N_18726,N_18797);
or U18833 (N_18833,N_18747,N_18702);
or U18834 (N_18834,N_18791,N_18795);
xnor U18835 (N_18835,N_18616,N_18717);
and U18836 (N_18836,N_18636,N_18701);
and U18837 (N_18837,N_18714,N_18614);
and U18838 (N_18838,N_18656,N_18670);
or U18839 (N_18839,N_18648,N_18731);
xnor U18840 (N_18840,N_18639,N_18708);
nor U18841 (N_18841,N_18711,N_18789);
and U18842 (N_18842,N_18730,N_18673);
or U18843 (N_18843,N_18724,N_18761);
xnor U18844 (N_18844,N_18773,N_18715);
and U18845 (N_18845,N_18763,N_18615);
xnor U18846 (N_18846,N_18704,N_18734);
xnor U18847 (N_18847,N_18628,N_18680);
and U18848 (N_18848,N_18780,N_18692);
or U18849 (N_18849,N_18630,N_18737);
xor U18850 (N_18850,N_18694,N_18721);
or U18851 (N_18851,N_18733,N_18776);
and U18852 (N_18852,N_18669,N_18750);
and U18853 (N_18853,N_18624,N_18720);
xnor U18854 (N_18854,N_18713,N_18674);
or U18855 (N_18855,N_18777,N_18653);
or U18856 (N_18856,N_18663,N_18629);
nand U18857 (N_18857,N_18659,N_18735);
or U18858 (N_18858,N_18758,N_18622);
nand U18859 (N_18859,N_18759,N_18690);
xor U18860 (N_18860,N_18770,N_18796);
and U18861 (N_18861,N_18647,N_18661);
and U18862 (N_18862,N_18752,N_18640);
nand U18863 (N_18863,N_18685,N_18666);
xnor U18864 (N_18864,N_18771,N_18775);
xor U18865 (N_18865,N_18652,N_18772);
and U18866 (N_18866,N_18606,N_18783);
nor U18867 (N_18867,N_18785,N_18644);
xor U18868 (N_18868,N_18613,N_18756);
xnor U18869 (N_18869,N_18665,N_18790);
or U18870 (N_18870,N_18679,N_18662);
nand U18871 (N_18871,N_18645,N_18698);
or U18872 (N_18872,N_18710,N_18602);
and U18873 (N_18873,N_18687,N_18620);
nor U18874 (N_18874,N_18784,N_18631);
nor U18875 (N_18875,N_18755,N_18707);
and U18876 (N_18876,N_18699,N_18691);
nor U18877 (N_18877,N_18654,N_18774);
xnor U18878 (N_18878,N_18684,N_18762);
nand U18879 (N_18879,N_18768,N_18664);
or U18880 (N_18880,N_18722,N_18794);
nand U18881 (N_18881,N_18736,N_18782);
xnor U18882 (N_18882,N_18650,N_18642);
xnor U18883 (N_18883,N_18786,N_18637);
xnor U18884 (N_18884,N_18746,N_18696);
nor U18885 (N_18885,N_18668,N_18778);
and U18886 (N_18886,N_18744,N_18627);
nand U18887 (N_18887,N_18706,N_18657);
and U18888 (N_18888,N_18792,N_18695);
and U18889 (N_18889,N_18625,N_18686);
xnor U18890 (N_18890,N_18709,N_18617);
or U18891 (N_18891,N_18607,N_18753);
xnor U18892 (N_18892,N_18793,N_18610);
or U18893 (N_18893,N_18612,N_18739);
xnor U18894 (N_18894,N_18788,N_18619);
and U18895 (N_18895,N_18618,N_18626);
nor U18896 (N_18896,N_18621,N_18725);
xor U18897 (N_18897,N_18649,N_18671);
xnor U18898 (N_18898,N_18757,N_18741);
and U18899 (N_18899,N_18703,N_18729);
and U18900 (N_18900,N_18746,N_18712);
or U18901 (N_18901,N_18675,N_18653);
or U18902 (N_18902,N_18742,N_18605);
xnor U18903 (N_18903,N_18670,N_18744);
nand U18904 (N_18904,N_18641,N_18645);
xor U18905 (N_18905,N_18643,N_18664);
nand U18906 (N_18906,N_18728,N_18768);
xnor U18907 (N_18907,N_18671,N_18772);
xnor U18908 (N_18908,N_18703,N_18649);
nand U18909 (N_18909,N_18694,N_18753);
or U18910 (N_18910,N_18638,N_18748);
and U18911 (N_18911,N_18635,N_18752);
or U18912 (N_18912,N_18728,N_18606);
xnor U18913 (N_18913,N_18791,N_18615);
nor U18914 (N_18914,N_18786,N_18799);
and U18915 (N_18915,N_18629,N_18681);
nand U18916 (N_18916,N_18676,N_18610);
nor U18917 (N_18917,N_18673,N_18614);
or U18918 (N_18918,N_18707,N_18747);
nand U18919 (N_18919,N_18606,N_18757);
nand U18920 (N_18920,N_18622,N_18683);
nand U18921 (N_18921,N_18673,N_18702);
or U18922 (N_18922,N_18618,N_18735);
nand U18923 (N_18923,N_18686,N_18731);
xor U18924 (N_18924,N_18675,N_18637);
nor U18925 (N_18925,N_18767,N_18629);
and U18926 (N_18926,N_18760,N_18746);
and U18927 (N_18927,N_18670,N_18620);
xor U18928 (N_18928,N_18653,N_18669);
nor U18929 (N_18929,N_18624,N_18742);
and U18930 (N_18930,N_18656,N_18768);
or U18931 (N_18931,N_18675,N_18693);
nor U18932 (N_18932,N_18633,N_18780);
nor U18933 (N_18933,N_18737,N_18716);
xor U18934 (N_18934,N_18797,N_18694);
nor U18935 (N_18935,N_18689,N_18705);
and U18936 (N_18936,N_18635,N_18608);
or U18937 (N_18937,N_18796,N_18736);
nand U18938 (N_18938,N_18671,N_18793);
or U18939 (N_18939,N_18714,N_18766);
or U18940 (N_18940,N_18797,N_18616);
or U18941 (N_18941,N_18608,N_18778);
or U18942 (N_18942,N_18772,N_18796);
nor U18943 (N_18943,N_18614,N_18631);
or U18944 (N_18944,N_18607,N_18605);
or U18945 (N_18945,N_18652,N_18692);
or U18946 (N_18946,N_18713,N_18699);
or U18947 (N_18947,N_18664,N_18698);
nor U18948 (N_18948,N_18749,N_18712);
and U18949 (N_18949,N_18610,N_18777);
or U18950 (N_18950,N_18774,N_18619);
xor U18951 (N_18951,N_18645,N_18705);
or U18952 (N_18952,N_18687,N_18689);
xor U18953 (N_18953,N_18639,N_18635);
xnor U18954 (N_18954,N_18748,N_18707);
and U18955 (N_18955,N_18627,N_18720);
and U18956 (N_18956,N_18609,N_18657);
xor U18957 (N_18957,N_18791,N_18712);
or U18958 (N_18958,N_18640,N_18798);
nor U18959 (N_18959,N_18758,N_18740);
nand U18960 (N_18960,N_18730,N_18691);
xnor U18961 (N_18961,N_18648,N_18735);
nand U18962 (N_18962,N_18747,N_18663);
nor U18963 (N_18963,N_18641,N_18669);
nand U18964 (N_18964,N_18625,N_18621);
nor U18965 (N_18965,N_18784,N_18650);
xnor U18966 (N_18966,N_18730,N_18764);
xnor U18967 (N_18967,N_18785,N_18690);
xnor U18968 (N_18968,N_18778,N_18631);
or U18969 (N_18969,N_18721,N_18653);
and U18970 (N_18970,N_18704,N_18647);
xor U18971 (N_18971,N_18630,N_18739);
and U18972 (N_18972,N_18692,N_18722);
xnor U18973 (N_18973,N_18790,N_18616);
nand U18974 (N_18974,N_18617,N_18764);
nand U18975 (N_18975,N_18797,N_18671);
or U18976 (N_18976,N_18658,N_18760);
xnor U18977 (N_18977,N_18738,N_18785);
nand U18978 (N_18978,N_18751,N_18604);
nand U18979 (N_18979,N_18778,N_18615);
nor U18980 (N_18980,N_18735,N_18734);
or U18981 (N_18981,N_18760,N_18689);
and U18982 (N_18982,N_18772,N_18691);
and U18983 (N_18983,N_18606,N_18741);
nor U18984 (N_18984,N_18667,N_18687);
nor U18985 (N_18985,N_18668,N_18700);
nand U18986 (N_18986,N_18601,N_18636);
xnor U18987 (N_18987,N_18730,N_18652);
nor U18988 (N_18988,N_18638,N_18635);
nor U18989 (N_18989,N_18709,N_18685);
nand U18990 (N_18990,N_18604,N_18684);
and U18991 (N_18991,N_18699,N_18798);
nand U18992 (N_18992,N_18640,N_18695);
or U18993 (N_18993,N_18639,N_18742);
nand U18994 (N_18994,N_18753,N_18742);
nor U18995 (N_18995,N_18747,N_18750);
or U18996 (N_18996,N_18757,N_18701);
and U18997 (N_18997,N_18621,N_18622);
xnor U18998 (N_18998,N_18640,N_18783);
and U18999 (N_18999,N_18751,N_18782);
and U19000 (N_19000,N_18918,N_18838);
nor U19001 (N_19001,N_18863,N_18980);
and U19002 (N_19002,N_18801,N_18826);
nor U19003 (N_19003,N_18875,N_18988);
and U19004 (N_19004,N_18845,N_18902);
xnor U19005 (N_19005,N_18944,N_18858);
nand U19006 (N_19006,N_18962,N_18813);
nand U19007 (N_19007,N_18814,N_18898);
nand U19008 (N_19008,N_18879,N_18954);
or U19009 (N_19009,N_18904,N_18855);
xnor U19010 (N_19010,N_18862,N_18880);
and U19011 (N_19011,N_18846,N_18803);
and U19012 (N_19012,N_18854,N_18874);
nor U19013 (N_19013,N_18828,N_18866);
or U19014 (N_19014,N_18834,N_18892);
nor U19015 (N_19015,N_18885,N_18881);
nand U19016 (N_19016,N_18946,N_18939);
xor U19017 (N_19017,N_18850,N_18809);
xor U19018 (N_19018,N_18975,N_18965);
xnor U19019 (N_19019,N_18808,N_18891);
and U19020 (N_19020,N_18893,N_18934);
nor U19021 (N_19021,N_18938,N_18847);
and U19022 (N_19022,N_18958,N_18986);
nand U19023 (N_19023,N_18802,N_18851);
nor U19024 (N_19024,N_18816,N_18922);
or U19025 (N_19025,N_18833,N_18848);
or U19026 (N_19026,N_18910,N_18900);
nor U19027 (N_19027,N_18835,N_18890);
nand U19028 (N_19028,N_18953,N_18989);
and U19029 (N_19029,N_18811,N_18932);
or U19030 (N_19030,N_18925,N_18987);
nand U19031 (N_19031,N_18810,N_18842);
xor U19032 (N_19032,N_18991,N_18873);
nand U19033 (N_19033,N_18889,N_18996);
nand U19034 (N_19034,N_18903,N_18919);
or U19035 (N_19035,N_18959,N_18941);
nand U19036 (N_19036,N_18815,N_18940);
or U19037 (N_19037,N_18859,N_18994);
or U19038 (N_19038,N_18955,N_18995);
and U19039 (N_19039,N_18818,N_18857);
or U19040 (N_19040,N_18886,N_18830);
and U19041 (N_19041,N_18884,N_18990);
nand U19042 (N_19042,N_18856,N_18906);
and U19043 (N_19043,N_18945,N_18908);
or U19044 (N_19044,N_18947,N_18825);
nor U19045 (N_19045,N_18817,N_18853);
xor U19046 (N_19046,N_18912,N_18871);
nor U19047 (N_19047,N_18951,N_18914);
xor U19048 (N_19048,N_18878,N_18992);
or U19049 (N_19049,N_18957,N_18887);
xnor U19050 (N_19050,N_18829,N_18819);
nand U19051 (N_19051,N_18942,N_18971);
or U19052 (N_19052,N_18870,N_18868);
nor U19053 (N_19053,N_18909,N_18901);
or U19054 (N_19054,N_18981,N_18929);
nor U19055 (N_19055,N_18974,N_18841);
xor U19056 (N_19056,N_18812,N_18832);
or U19057 (N_19057,N_18831,N_18923);
or U19058 (N_19058,N_18800,N_18948);
nor U19059 (N_19059,N_18964,N_18979);
or U19060 (N_19060,N_18935,N_18915);
nor U19061 (N_19061,N_18933,N_18877);
nor U19062 (N_19062,N_18961,N_18894);
and U19063 (N_19063,N_18930,N_18843);
nor U19064 (N_19064,N_18888,N_18982);
or U19065 (N_19065,N_18949,N_18907);
and U19066 (N_19066,N_18997,N_18849);
xor U19067 (N_19067,N_18916,N_18928);
and U19068 (N_19068,N_18911,N_18896);
nor U19069 (N_19069,N_18865,N_18805);
or U19070 (N_19070,N_18973,N_18924);
nor U19071 (N_19071,N_18876,N_18984);
nand U19072 (N_19072,N_18899,N_18972);
and U19073 (N_19073,N_18998,N_18883);
or U19074 (N_19074,N_18860,N_18993);
xor U19075 (N_19075,N_18852,N_18963);
nand U19076 (N_19076,N_18966,N_18927);
xor U19077 (N_19077,N_18960,N_18806);
nand U19078 (N_19078,N_18917,N_18823);
or U19079 (N_19079,N_18869,N_18839);
or U19080 (N_19080,N_18967,N_18985);
nor U19081 (N_19081,N_18836,N_18837);
or U19082 (N_19082,N_18920,N_18978);
xor U19083 (N_19083,N_18844,N_18872);
nor U19084 (N_19084,N_18937,N_18820);
and U19085 (N_19085,N_18950,N_18824);
xnor U19086 (N_19086,N_18807,N_18827);
nand U19087 (N_19087,N_18895,N_18921);
nor U19088 (N_19088,N_18861,N_18968);
nand U19089 (N_19089,N_18822,N_18905);
and U19090 (N_19090,N_18840,N_18999);
nor U19091 (N_19091,N_18926,N_18977);
nor U19092 (N_19092,N_18864,N_18882);
and U19093 (N_19093,N_18943,N_18897);
nor U19094 (N_19094,N_18913,N_18976);
or U19095 (N_19095,N_18983,N_18804);
nand U19096 (N_19096,N_18970,N_18952);
nand U19097 (N_19097,N_18821,N_18867);
nand U19098 (N_19098,N_18936,N_18956);
nand U19099 (N_19099,N_18969,N_18931);
nand U19100 (N_19100,N_18825,N_18844);
xnor U19101 (N_19101,N_18857,N_18934);
and U19102 (N_19102,N_18803,N_18917);
nand U19103 (N_19103,N_18937,N_18911);
nand U19104 (N_19104,N_18879,N_18822);
and U19105 (N_19105,N_18877,N_18847);
xnor U19106 (N_19106,N_18863,N_18930);
and U19107 (N_19107,N_18825,N_18848);
or U19108 (N_19108,N_18857,N_18991);
nor U19109 (N_19109,N_18908,N_18971);
or U19110 (N_19110,N_18998,N_18929);
or U19111 (N_19111,N_18951,N_18893);
nand U19112 (N_19112,N_18811,N_18995);
xnor U19113 (N_19113,N_18951,N_18864);
and U19114 (N_19114,N_18850,N_18866);
xor U19115 (N_19115,N_18854,N_18969);
or U19116 (N_19116,N_18840,N_18998);
nand U19117 (N_19117,N_18948,N_18936);
and U19118 (N_19118,N_18934,N_18881);
nor U19119 (N_19119,N_18927,N_18855);
and U19120 (N_19120,N_18971,N_18800);
or U19121 (N_19121,N_18938,N_18865);
nand U19122 (N_19122,N_18866,N_18827);
nand U19123 (N_19123,N_18997,N_18859);
or U19124 (N_19124,N_18987,N_18902);
and U19125 (N_19125,N_18808,N_18965);
and U19126 (N_19126,N_18809,N_18973);
nor U19127 (N_19127,N_18914,N_18956);
nor U19128 (N_19128,N_18973,N_18964);
nand U19129 (N_19129,N_18957,N_18988);
or U19130 (N_19130,N_18899,N_18893);
xnor U19131 (N_19131,N_18931,N_18820);
nor U19132 (N_19132,N_18851,N_18889);
and U19133 (N_19133,N_18871,N_18850);
xnor U19134 (N_19134,N_18870,N_18924);
and U19135 (N_19135,N_18864,N_18806);
nand U19136 (N_19136,N_18919,N_18815);
nor U19137 (N_19137,N_18972,N_18974);
and U19138 (N_19138,N_18939,N_18907);
nand U19139 (N_19139,N_18913,N_18876);
or U19140 (N_19140,N_18974,N_18954);
nand U19141 (N_19141,N_18992,N_18997);
xor U19142 (N_19142,N_18810,N_18899);
nand U19143 (N_19143,N_18993,N_18895);
or U19144 (N_19144,N_18915,N_18830);
and U19145 (N_19145,N_18977,N_18858);
nor U19146 (N_19146,N_18802,N_18955);
and U19147 (N_19147,N_18868,N_18969);
xnor U19148 (N_19148,N_18876,N_18851);
nand U19149 (N_19149,N_18991,N_18980);
or U19150 (N_19150,N_18925,N_18914);
or U19151 (N_19151,N_18926,N_18985);
nand U19152 (N_19152,N_18874,N_18824);
nand U19153 (N_19153,N_18930,N_18911);
and U19154 (N_19154,N_18833,N_18901);
and U19155 (N_19155,N_18966,N_18881);
nand U19156 (N_19156,N_18968,N_18850);
and U19157 (N_19157,N_18984,N_18990);
nand U19158 (N_19158,N_18986,N_18916);
nand U19159 (N_19159,N_18874,N_18977);
and U19160 (N_19160,N_18949,N_18909);
and U19161 (N_19161,N_18811,N_18891);
xor U19162 (N_19162,N_18807,N_18873);
and U19163 (N_19163,N_18947,N_18816);
nor U19164 (N_19164,N_18946,N_18950);
xor U19165 (N_19165,N_18861,N_18837);
or U19166 (N_19166,N_18908,N_18977);
or U19167 (N_19167,N_18900,N_18840);
nor U19168 (N_19168,N_18879,N_18889);
or U19169 (N_19169,N_18811,N_18910);
nor U19170 (N_19170,N_18958,N_18909);
nand U19171 (N_19171,N_18915,N_18837);
xor U19172 (N_19172,N_18841,N_18858);
xnor U19173 (N_19173,N_18959,N_18944);
xnor U19174 (N_19174,N_18803,N_18808);
and U19175 (N_19175,N_18943,N_18948);
and U19176 (N_19176,N_18890,N_18947);
nand U19177 (N_19177,N_18961,N_18916);
xnor U19178 (N_19178,N_18848,N_18957);
nand U19179 (N_19179,N_18918,N_18828);
nor U19180 (N_19180,N_18930,N_18912);
and U19181 (N_19181,N_18882,N_18878);
xnor U19182 (N_19182,N_18861,N_18886);
and U19183 (N_19183,N_18824,N_18923);
xnor U19184 (N_19184,N_18948,N_18996);
nor U19185 (N_19185,N_18842,N_18863);
and U19186 (N_19186,N_18873,N_18906);
xnor U19187 (N_19187,N_18985,N_18957);
nor U19188 (N_19188,N_18904,N_18996);
nor U19189 (N_19189,N_18903,N_18962);
xor U19190 (N_19190,N_18955,N_18810);
nor U19191 (N_19191,N_18913,N_18820);
nor U19192 (N_19192,N_18975,N_18802);
nand U19193 (N_19193,N_18926,N_18933);
nor U19194 (N_19194,N_18994,N_18983);
nand U19195 (N_19195,N_18978,N_18953);
or U19196 (N_19196,N_18833,N_18978);
nand U19197 (N_19197,N_18862,N_18911);
and U19198 (N_19198,N_18962,N_18865);
nor U19199 (N_19199,N_18806,N_18814);
nor U19200 (N_19200,N_19187,N_19022);
nand U19201 (N_19201,N_19100,N_19003);
xnor U19202 (N_19202,N_19058,N_19101);
or U19203 (N_19203,N_19031,N_19122);
xor U19204 (N_19204,N_19070,N_19159);
and U19205 (N_19205,N_19179,N_19150);
or U19206 (N_19206,N_19000,N_19098);
and U19207 (N_19207,N_19182,N_19132);
xor U19208 (N_19208,N_19171,N_19020);
and U19209 (N_19209,N_19166,N_19034);
xnor U19210 (N_19210,N_19117,N_19118);
nand U19211 (N_19211,N_19040,N_19078);
nor U19212 (N_19212,N_19061,N_19199);
xor U19213 (N_19213,N_19093,N_19069);
or U19214 (N_19214,N_19115,N_19110);
nand U19215 (N_19215,N_19194,N_19006);
nand U19216 (N_19216,N_19081,N_19095);
xor U19217 (N_19217,N_19025,N_19176);
or U19218 (N_19218,N_19116,N_19133);
and U19219 (N_19219,N_19195,N_19173);
and U19220 (N_19220,N_19074,N_19027);
nand U19221 (N_19221,N_19043,N_19083);
xnor U19222 (N_19222,N_19044,N_19155);
nand U19223 (N_19223,N_19036,N_19158);
nor U19224 (N_19224,N_19143,N_19090);
nor U19225 (N_19225,N_19151,N_19029);
xnor U19226 (N_19226,N_19005,N_19124);
nor U19227 (N_19227,N_19128,N_19041);
nand U19228 (N_19228,N_19059,N_19190);
xor U19229 (N_19229,N_19014,N_19053);
nand U19230 (N_19230,N_19008,N_19102);
xnor U19231 (N_19231,N_19096,N_19156);
nand U19232 (N_19232,N_19112,N_19021);
xor U19233 (N_19233,N_19170,N_19120);
nand U19234 (N_19234,N_19049,N_19088);
nor U19235 (N_19235,N_19015,N_19048);
nand U19236 (N_19236,N_19001,N_19146);
nor U19237 (N_19237,N_19172,N_19052);
and U19238 (N_19238,N_19032,N_19189);
and U19239 (N_19239,N_19129,N_19063);
nand U19240 (N_19240,N_19094,N_19138);
or U19241 (N_19241,N_19144,N_19186);
or U19242 (N_19242,N_19039,N_19180);
xnor U19243 (N_19243,N_19157,N_19033);
or U19244 (N_19244,N_19071,N_19068);
xnor U19245 (N_19245,N_19177,N_19099);
nand U19246 (N_19246,N_19026,N_19178);
nor U19247 (N_19247,N_19185,N_19057);
and U19248 (N_19248,N_19079,N_19136);
and U19249 (N_19249,N_19114,N_19105);
nor U19250 (N_19250,N_19097,N_19089);
nand U19251 (N_19251,N_19140,N_19017);
xnor U19252 (N_19252,N_19051,N_19073);
nor U19253 (N_19253,N_19012,N_19145);
and U19254 (N_19254,N_19137,N_19126);
nand U19255 (N_19255,N_19060,N_19160);
and U19256 (N_19256,N_19056,N_19169);
and U19257 (N_19257,N_19107,N_19084);
and U19258 (N_19258,N_19002,N_19154);
nor U19259 (N_19259,N_19113,N_19062);
xor U19260 (N_19260,N_19192,N_19103);
nor U19261 (N_19261,N_19024,N_19065);
nand U19262 (N_19262,N_19050,N_19141);
xnor U19263 (N_19263,N_19193,N_19086);
nor U19264 (N_19264,N_19127,N_19064);
nor U19265 (N_19265,N_19168,N_19191);
or U19266 (N_19266,N_19010,N_19167);
and U19267 (N_19267,N_19184,N_19131);
or U19268 (N_19268,N_19121,N_19066);
nor U19269 (N_19269,N_19018,N_19130);
or U19270 (N_19270,N_19030,N_19123);
nor U19271 (N_19271,N_19004,N_19152);
and U19272 (N_19272,N_19109,N_19135);
and U19273 (N_19273,N_19111,N_19082);
xor U19274 (N_19274,N_19188,N_19075);
nor U19275 (N_19275,N_19077,N_19148);
nor U19276 (N_19276,N_19067,N_19009);
or U19277 (N_19277,N_19104,N_19119);
nand U19278 (N_19278,N_19019,N_19161);
and U19279 (N_19279,N_19055,N_19028);
nand U19280 (N_19280,N_19080,N_19016);
or U19281 (N_19281,N_19037,N_19134);
nor U19282 (N_19282,N_19147,N_19042);
and U19283 (N_19283,N_19035,N_19164);
and U19284 (N_19284,N_19085,N_19038);
nor U19285 (N_19285,N_19023,N_19087);
nor U19286 (N_19286,N_19139,N_19142);
nand U19287 (N_19287,N_19197,N_19007);
or U19288 (N_19288,N_19092,N_19054);
or U19289 (N_19289,N_19163,N_19125);
nand U19290 (N_19290,N_19013,N_19198);
xor U19291 (N_19291,N_19091,N_19076);
and U19292 (N_19292,N_19165,N_19181);
and U19293 (N_19293,N_19047,N_19011);
and U19294 (N_19294,N_19174,N_19196);
nand U19295 (N_19295,N_19045,N_19183);
xor U19296 (N_19296,N_19149,N_19046);
nor U19297 (N_19297,N_19162,N_19108);
or U19298 (N_19298,N_19106,N_19072);
or U19299 (N_19299,N_19175,N_19153);
and U19300 (N_19300,N_19123,N_19018);
xnor U19301 (N_19301,N_19053,N_19013);
and U19302 (N_19302,N_19117,N_19080);
or U19303 (N_19303,N_19180,N_19174);
or U19304 (N_19304,N_19016,N_19107);
and U19305 (N_19305,N_19022,N_19169);
and U19306 (N_19306,N_19109,N_19129);
nor U19307 (N_19307,N_19131,N_19194);
xnor U19308 (N_19308,N_19193,N_19151);
or U19309 (N_19309,N_19048,N_19120);
and U19310 (N_19310,N_19093,N_19156);
nor U19311 (N_19311,N_19127,N_19034);
xor U19312 (N_19312,N_19147,N_19027);
nand U19313 (N_19313,N_19081,N_19053);
xor U19314 (N_19314,N_19053,N_19168);
nand U19315 (N_19315,N_19064,N_19088);
nor U19316 (N_19316,N_19089,N_19178);
and U19317 (N_19317,N_19068,N_19187);
nand U19318 (N_19318,N_19039,N_19018);
or U19319 (N_19319,N_19187,N_19040);
or U19320 (N_19320,N_19028,N_19141);
and U19321 (N_19321,N_19045,N_19153);
xor U19322 (N_19322,N_19149,N_19120);
nand U19323 (N_19323,N_19025,N_19012);
nor U19324 (N_19324,N_19064,N_19130);
and U19325 (N_19325,N_19144,N_19165);
xor U19326 (N_19326,N_19199,N_19119);
nand U19327 (N_19327,N_19027,N_19107);
nor U19328 (N_19328,N_19133,N_19058);
nor U19329 (N_19329,N_19132,N_19151);
or U19330 (N_19330,N_19190,N_19057);
nand U19331 (N_19331,N_19013,N_19107);
xnor U19332 (N_19332,N_19049,N_19033);
xnor U19333 (N_19333,N_19116,N_19026);
nor U19334 (N_19334,N_19098,N_19117);
nand U19335 (N_19335,N_19014,N_19161);
nor U19336 (N_19336,N_19005,N_19019);
xnor U19337 (N_19337,N_19056,N_19064);
xor U19338 (N_19338,N_19137,N_19169);
nor U19339 (N_19339,N_19141,N_19191);
and U19340 (N_19340,N_19086,N_19143);
and U19341 (N_19341,N_19129,N_19074);
nand U19342 (N_19342,N_19128,N_19053);
nand U19343 (N_19343,N_19009,N_19107);
xnor U19344 (N_19344,N_19044,N_19132);
nor U19345 (N_19345,N_19178,N_19030);
xor U19346 (N_19346,N_19133,N_19046);
and U19347 (N_19347,N_19138,N_19022);
nand U19348 (N_19348,N_19090,N_19157);
nand U19349 (N_19349,N_19195,N_19104);
nand U19350 (N_19350,N_19191,N_19131);
nand U19351 (N_19351,N_19063,N_19013);
nor U19352 (N_19352,N_19190,N_19199);
nor U19353 (N_19353,N_19105,N_19165);
nand U19354 (N_19354,N_19034,N_19191);
xor U19355 (N_19355,N_19130,N_19183);
nand U19356 (N_19356,N_19005,N_19196);
and U19357 (N_19357,N_19166,N_19194);
or U19358 (N_19358,N_19108,N_19177);
nand U19359 (N_19359,N_19132,N_19168);
or U19360 (N_19360,N_19037,N_19062);
and U19361 (N_19361,N_19034,N_19063);
nor U19362 (N_19362,N_19129,N_19100);
and U19363 (N_19363,N_19197,N_19130);
nor U19364 (N_19364,N_19080,N_19038);
nor U19365 (N_19365,N_19089,N_19052);
or U19366 (N_19366,N_19199,N_19002);
or U19367 (N_19367,N_19195,N_19189);
and U19368 (N_19368,N_19150,N_19012);
nor U19369 (N_19369,N_19050,N_19045);
or U19370 (N_19370,N_19112,N_19000);
xnor U19371 (N_19371,N_19077,N_19146);
nand U19372 (N_19372,N_19087,N_19187);
nand U19373 (N_19373,N_19084,N_19092);
xor U19374 (N_19374,N_19148,N_19199);
and U19375 (N_19375,N_19040,N_19185);
nor U19376 (N_19376,N_19095,N_19004);
nand U19377 (N_19377,N_19034,N_19098);
or U19378 (N_19378,N_19056,N_19011);
nor U19379 (N_19379,N_19188,N_19162);
nand U19380 (N_19380,N_19015,N_19068);
nor U19381 (N_19381,N_19162,N_19040);
nand U19382 (N_19382,N_19073,N_19002);
and U19383 (N_19383,N_19066,N_19135);
and U19384 (N_19384,N_19045,N_19068);
xnor U19385 (N_19385,N_19150,N_19142);
nor U19386 (N_19386,N_19097,N_19057);
xnor U19387 (N_19387,N_19057,N_19077);
nor U19388 (N_19388,N_19119,N_19175);
or U19389 (N_19389,N_19014,N_19091);
xor U19390 (N_19390,N_19075,N_19162);
nand U19391 (N_19391,N_19183,N_19017);
nor U19392 (N_19392,N_19039,N_19058);
nor U19393 (N_19393,N_19030,N_19075);
or U19394 (N_19394,N_19144,N_19057);
xor U19395 (N_19395,N_19008,N_19186);
and U19396 (N_19396,N_19136,N_19151);
nand U19397 (N_19397,N_19190,N_19143);
xor U19398 (N_19398,N_19118,N_19141);
xnor U19399 (N_19399,N_19171,N_19128);
or U19400 (N_19400,N_19295,N_19333);
nor U19401 (N_19401,N_19278,N_19228);
or U19402 (N_19402,N_19214,N_19327);
nor U19403 (N_19403,N_19218,N_19282);
or U19404 (N_19404,N_19202,N_19280);
nand U19405 (N_19405,N_19323,N_19245);
nand U19406 (N_19406,N_19331,N_19366);
or U19407 (N_19407,N_19240,N_19233);
nor U19408 (N_19408,N_19312,N_19258);
nor U19409 (N_19409,N_19390,N_19203);
and U19410 (N_19410,N_19296,N_19384);
nand U19411 (N_19411,N_19306,N_19330);
nor U19412 (N_19412,N_19362,N_19342);
or U19413 (N_19413,N_19381,N_19298);
nand U19414 (N_19414,N_19205,N_19287);
nor U19415 (N_19415,N_19346,N_19399);
and U19416 (N_19416,N_19373,N_19253);
and U19417 (N_19417,N_19397,N_19372);
xnor U19418 (N_19418,N_19355,N_19208);
nand U19419 (N_19419,N_19246,N_19269);
xor U19420 (N_19420,N_19250,N_19315);
or U19421 (N_19421,N_19222,N_19207);
and U19422 (N_19422,N_19386,N_19236);
xor U19423 (N_19423,N_19304,N_19393);
nand U19424 (N_19424,N_19337,N_19395);
xnor U19425 (N_19425,N_19396,N_19279);
or U19426 (N_19426,N_19369,N_19285);
nand U19427 (N_19427,N_19284,N_19271);
nand U19428 (N_19428,N_19272,N_19345);
xor U19429 (N_19429,N_19297,N_19326);
xnor U19430 (N_19430,N_19354,N_19379);
xnor U19431 (N_19431,N_19352,N_19394);
or U19432 (N_19432,N_19343,N_19249);
nand U19433 (N_19433,N_19252,N_19398);
and U19434 (N_19434,N_19367,N_19294);
and U19435 (N_19435,N_19350,N_19229);
nand U19436 (N_19436,N_19359,N_19365);
xor U19437 (N_19437,N_19358,N_19314);
nor U19438 (N_19438,N_19225,N_19257);
nor U19439 (N_19439,N_19310,N_19389);
xor U19440 (N_19440,N_19235,N_19300);
and U19441 (N_19441,N_19264,N_19290);
and U19442 (N_19442,N_19319,N_19200);
or U19443 (N_19443,N_19232,N_19204);
and U19444 (N_19444,N_19242,N_19224);
nand U19445 (N_19445,N_19237,N_19274);
or U19446 (N_19446,N_19288,N_19316);
nand U19447 (N_19447,N_19324,N_19217);
nor U19448 (N_19448,N_19338,N_19223);
xor U19449 (N_19449,N_19378,N_19388);
nand U19450 (N_19450,N_19201,N_19351);
xnor U19451 (N_19451,N_19244,N_19377);
or U19452 (N_19452,N_19347,N_19322);
or U19453 (N_19453,N_19344,N_19227);
xnor U19454 (N_19454,N_19230,N_19241);
and U19455 (N_19455,N_19275,N_19387);
and U19456 (N_19456,N_19318,N_19270);
or U19457 (N_19457,N_19339,N_19392);
xnor U19458 (N_19458,N_19260,N_19216);
nor U19459 (N_19459,N_19238,N_19317);
nand U19460 (N_19460,N_19231,N_19305);
nor U19461 (N_19461,N_19311,N_19265);
nand U19462 (N_19462,N_19353,N_19239);
nand U19463 (N_19463,N_19206,N_19209);
and U19464 (N_19464,N_19375,N_19283);
or U19465 (N_19465,N_19266,N_19334);
nor U19466 (N_19466,N_19307,N_19289);
nand U19467 (N_19467,N_19325,N_19301);
nand U19468 (N_19468,N_19226,N_19374);
or U19469 (N_19469,N_19340,N_19267);
and U19470 (N_19470,N_19368,N_19313);
or U19471 (N_19471,N_19210,N_19255);
nand U19472 (N_19472,N_19309,N_19211);
nor U19473 (N_19473,N_19251,N_19268);
nand U19474 (N_19474,N_19286,N_19360);
nand U19475 (N_19475,N_19302,N_19341);
or U19476 (N_19476,N_19361,N_19221);
xor U19477 (N_19477,N_19248,N_19263);
nand U19478 (N_19478,N_19380,N_19215);
and U19479 (N_19479,N_19308,N_19219);
or U19480 (N_19480,N_19371,N_19370);
nor U19481 (N_19481,N_19303,N_19328);
or U19482 (N_19482,N_19321,N_19348);
xor U19483 (N_19483,N_19234,N_19243);
or U19484 (N_19484,N_19254,N_19281);
and U19485 (N_19485,N_19292,N_19276);
nand U19486 (N_19486,N_19364,N_19261);
nor U19487 (N_19487,N_19256,N_19220);
xnor U19488 (N_19488,N_19320,N_19363);
and U19489 (N_19489,N_19293,N_19391);
or U19490 (N_19490,N_19262,N_19329);
nor U19491 (N_19491,N_19299,N_19356);
and U19492 (N_19492,N_19357,N_19291);
or U19493 (N_19493,N_19383,N_19247);
nand U19494 (N_19494,N_19376,N_19212);
nand U19495 (N_19495,N_19349,N_19385);
xor U19496 (N_19496,N_19336,N_19213);
xnor U19497 (N_19497,N_19273,N_19335);
nand U19498 (N_19498,N_19382,N_19332);
xnor U19499 (N_19499,N_19277,N_19259);
and U19500 (N_19500,N_19367,N_19389);
or U19501 (N_19501,N_19241,N_19279);
or U19502 (N_19502,N_19283,N_19357);
and U19503 (N_19503,N_19346,N_19203);
nand U19504 (N_19504,N_19356,N_19219);
nor U19505 (N_19505,N_19300,N_19323);
and U19506 (N_19506,N_19350,N_19283);
or U19507 (N_19507,N_19358,N_19268);
xnor U19508 (N_19508,N_19388,N_19348);
nor U19509 (N_19509,N_19207,N_19297);
nand U19510 (N_19510,N_19334,N_19274);
nand U19511 (N_19511,N_19251,N_19357);
xor U19512 (N_19512,N_19235,N_19306);
nor U19513 (N_19513,N_19365,N_19229);
and U19514 (N_19514,N_19380,N_19245);
xor U19515 (N_19515,N_19358,N_19322);
nor U19516 (N_19516,N_19373,N_19387);
xor U19517 (N_19517,N_19357,N_19332);
nor U19518 (N_19518,N_19240,N_19289);
xnor U19519 (N_19519,N_19248,N_19284);
nor U19520 (N_19520,N_19274,N_19295);
nand U19521 (N_19521,N_19365,N_19249);
nand U19522 (N_19522,N_19314,N_19345);
nor U19523 (N_19523,N_19395,N_19306);
nand U19524 (N_19524,N_19287,N_19261);
or U19525 (N_19525,N_19271,N_19268);
nor U19526 (N_19526,N_19392,N_19241);
and U19527 (N_19527,N_19303,N_19278);
or U19528 (N_19528,N_19225,N_19337);
nor U19529 (N_19529,N_19381,N_19274);
xnor U19530 (N_19530,N_19330,N_19230);
nand U19531 (N_19531,N_19373,N_19318);
nand U19532 (N_19532,N_19302,N_19262);
nor U19533 (N_19533,N_19210,N_19281);
and U19534 (N_19534,N_19228,N_19260);
or U19535 (N_19535,N_19293,N_19312);
nand U19536 (N_19536,N_19308,N_19326);
nand U19537 (N_19537,N_19298,N_19263);
or U19538 (N_19538,N_19279,N_19216);
xnor U19539 (N_19539,N_19287,N_19202);
nand U19540 (N_19540,N_19242,N_19249);
and U19541 (N_19541,N_19269,N_19313);
and U19542 (N_19542,N_19345,N_19201);
and U19543 (N_19543,N_19251,N_19299);
and U19544 (N_19544,N_19310,N_19247);
or U19545 (N_19545,N_19208,N_19360);
nand U19546 (N_19546,N_19244,N_19253);
or U19547 (N_19547,N_19383,N_19202);
or U19548 (N_19548,N_19238,N_19369);
xor U19549 (N_19549,N_19308,N_19234);
nand U19550 (N_19550,N_19255,N_19247);
nor U19551 (N_19551,N_19281,N_19332);
or U19552 (N_19552,N_19349,N_19222);
or U19553 (N_19553,N_19336,N_19310);
nor U19554 (N_19554,N_19230,N_19240);
nand U19555 (N_19555,N_19335,N_19321);
and U19556 (N_19556,N_19221,N_19385);
or U19557 (N_19557,N_19356,N_19313);
nand U19558 (N_19558,N_19327,N_19235);
nand U19559 (N_19559,N_19201,N_19354);
nor U19560 (N_19560,N_19223,N_19265);
nor U19561 (N_19561,N_19205,N_19322);
nand U19562 (N_19562,N_19223,N_19230);
and U19563 (N_19563,N_19360,N_19328);
and U19564 (N_19564,N_19281,N_19374);
xor U19565 (N_19565,N_19257,N_19277);
xnor U19566 (N_19566,N_19285,N_19257);
nor U19567 (N_19567,N_19303,N_19333);
or U19568 (N_19568,N_19233,N_19345);
nand U19569 (N_19569,N_19355,N_19271);
nand U19570 (N_19570,N_19291,N_19379);
xnor U19571 (N_19571,N_19213,N_19247);
xor U19572 (N_19572,N_19291,N_19228);
xnor U19573 (N_19573,N_19279,N_19219);
or U19574 (N_19574,N_19394,N_19248);
nand U19575 (N_19575,N_19229,N_19294);
nor U19576 (N_19576,N_19225,N_19325);
nand U19577 (N_19577,N_19281,N_19379);
nor U19578 (N_19578,N_19374,N_19390);
xnor U19579 (N_19579,N_19232,N_19292);
xor U19580 (N_19580,N_19391,N_19247);
and U19581 (N_19581,N_19231,N_19394);
xor U19582 (N_19582,N_19368,N_19231);
and U19583 (N_19583,N_19380,N_19325);
nand U19584 (N_19584,N_19275,N_19318);
and U19585 (N_19585,N_19214,N_19312);
or U19586 (N_19586,N_19362,N_19350);
nand U19587 (N_19587,N_19266,N_19224);
nor U19588 (N_19588,N_19326,N_19388);
or U19589 (N_19589,N_19392,N_19396);
and U19590 (N_19590,N_19234,N_19281);
xor U19591 (N_19591,N_19276,N_19398);
and U19592 (N_19592,N_19357,N_19364);
nor U19593 (N_19593,N_19229,N_19353);
xor U19594 (N_19594,N_19373,N_19314);
nand U19595 (N_19595,N_19242,N_19339);
xor U19596 (N_19596,N_19319,N_19230);
nor U19597 (N_19597,N_19324,N_19244);
xnor U19598 (N_19598,N_19387,N_19344);
or U19599 (N_19599,N_19350,N_19393);
xor U19600 (N_19600,N_19520,N_19427);
xnor U19601 (N_19601,N_19508,N_19476);
or U19602 (N_19602,N_19527,N_19409);
or U19603 (N_19603,N_19578,N_19471);
nand U19604 (N_19604,N_19441,N_19473);
nand U19605 (N_19605,N_19599,N_19587);
nor U19606 (N_19606,N_19522,N_19435);
nand U19607 (N_19607,N_19431,N_19541);
and U19608 (N_19608,N_19536,N_19547);
and U19609 (N_19609,N_19448,N_19417);
xor U19610 (N_19610,N_19425,N_19485);
or U19611 (N_19611,N_19489,N_19436);
xor U19612 (N_19612,N_19492,N_19424);
nand U19613 (N_19613,N_19418,N_19574);
and U19614 (N_19614,N_19475,N_19458);
nor U19615 (N_19615,N_19483,N_19468);
nand U19616 (N_19616,N_19437,N_19443);
or U19617 (N_19617,N_19429,N_19538);
nor U19618 (N_19618,N_19400,N_19558);
or U19619 (N_19619,N_19432,N_19446);
or U19620 (N_19620,N_19430,N_19519);
or U19621 (N_19621,N_19466,N_19533);
or U19622 (N_19622,N_19516,N_19420);
nand U19623 (N_19623,N_19551,N_19532);
xor U19624 (N_19624,N_19449,N_19535);
xnor U19625 (N_19625,N_19543,N_19445);
xnor U19626 (N_19626,N_19524,N_19579);
or U19627 (N_19627,N_19404,N_19534);
or U19628 (N_19628,N_19461,N_19539);
nand U19629 (N_19629,N_19518,N_19593);
nand U19630 (N_19630,N_19584,N_19564);
and U19631 (N_19631,N_19572,N_19464);
nor U19632 (N_19632,N_19488,N_19598);
nand U19633 (N_19633,N_19451,N_19414);
or U19634 (N_19634,N_19582,N_19523);
or U19635 (N_19635,N_19470,N_19456);
and U19636 (N_19636,N_19490,N_19503);
nor U19637 (N_19637,N_19560,N_19462);
nor U19638 (N_19638,N_19549,N_19511);
nand U19639 (N_19639,N_19561,N_19596);
nor U19640 (N_19640,N_19563,N_19428);
nand U19641 (N_19641,N_19531,N_19416);
nor U19642 (N_19642,N_19559,N_19502);
xnor U19643 (N_19643,N_19433,N_19467);
and U19644 (N_19644,N_19506,N_19548);
xnor U19645 (N_19645,N_19501,N_19542);
xnor U19646 (N_19646,N_19465,N_19412);
nor U19647 (N_19647,N_19410,N_19591);
nand U19648 (N_19648,N_19571,N_19480);
nor U19649 (N_19649,N_19590,N_19546);
nand U19650 (N_19650,N_19455,N_19460);
or U19651 (N_19651,N_19595,N_19529);
nor U19652 (N_19652,N_19512,N_19528);
xor U19653 (N_19653,N_19500,N_19576);
and U19654 (N_19654,N_19413,N_19555);
or U19655 (N_19655,N_19575,N_19509);
xnor U19656 (N_19656,N_19459,N_19469);
xnor U19657 (N_19657,N_19521,N_19567);
nor U19658 (N_19658,N_19497,N_19550);
xor U19659 (N_19659,N_19517,N_19401);
and U19660 (N_19660,N_19407,N_19440);
nand U19661 (N_19661,N_19592,N_19566);
xor U19662 (N_19662,N_19447,N_19487);
xnor U19663 (N_19663,N_19463,N_19577);
xor U19664 (N_19664,N_19453,N_19484);
xnor U19665 (N_19665,N_19589,N_19588);
and U19666 (N_19666,N_19457,N_19408);
nand U19667 (N_19667,N_19477,N_19526);
and U19668 (N_19668,N_19495,N_19586);
or U19669 (N_19669,N_19537,N_19553);
xor U19670 (N_19670,N_19405,N_19493);
or U19671 (N_19671,N_19454,N_19507);
xor U19672 (N_19672,N_19434,N_19585);
and U19673 (N_19673,N_19554,N_19411);
xnor U19674 (N_19674,N_19494,N_19499);
or U19675 (N_19675,N_19486,N_19515);
nor U19676 (N_19676,N_19552,N_19530);
nand U19677 (N_19677,N_19573,N_19569);
and U19678 (N_19678,N_19444,N_19479);
nor U19679 (N_19679,N_19556,N_19496);
nand U19680 (N_19680,N_19568,N_19498);
or U19681 (N_19681,N_19422,N_19450);
and U19682 (N_19682,N_19505,N_19474);
and U19683 (N_19683,N_19406,N_19403);
nor U19684 (N_19684,N_19482,N_19557);
nor U19685 (N_19685,N_19580,N_19426);
or U19686 (N_19686,N_19491,N_19510);
and U19687 (N_19687,N_19597,N_19481);
nand U19688 (N_19688,N_19415,N_19525);
or U19689 (N_19689,N_19452,N_19583);
and U19690 (N_19690,N_19423,N_19504);
or U19691 (N_19691,N_19442,N_19565);
xor U19692 (N_19692,N_19419,N_19513);
or U19693 (N_19693,N_19581,N_19472);
or U19694 (N_19694,N_19570,N_19562);
xnor U19695 (N_19695,N_19545,N_19438);
xor U19696 (N_19696,N_19421,N_19540);
and U19697 (N_19697,N_19402,N_19439);
xor U19698 (N_19698,N_19514,N_19594);
nand U19699 (N_19699,N_19478,N_19544);
or U19700 (N_19700,N_19557,N_19599);
nand U19701 (N_19701,N_19400,N_19480);
or U19702 (N_19702,N_19545,N_19515);
nand U19703 (N_19703,N_19404,N_19523);
nor U19704 (N_19704,N_19569,N_19426);
xnor U19705 (N_19705,N_19580,N_19468);
nor U19706 (N_19706,N_19426,N_19535);
and U19707 (N_19707,N_19445,N_19435);
or U19708 (N_19708,N_19530,N_19589);
xor U19709 (N_19709,N_19527,N_19431);
or U19710 (N_19710,N_19552,N_19494);
nand U19711 (N_19711,N_19407,N_19405);
or U19712 (N_19712,N_19441,N_19485);
nor U19713 (N_19713,N_19469,N_19525);
xor U19714 (N_19714,N_19497,N_19553);
or U19715 (N_19715,N_19526,N_19432);
and U19716 (N_19716,N_19537,N_19412);
or U19717 (N_19717,N_19554,N_19493);
and U19718 (N_19718,N_19543,N_19457);
and U19719 (N_19719,N_19514,N_19436);
and U19720 (N_19720,N_19528,N_19542);
nand U19721 (N_19721,N_19503,N_19537);
xor U19722 (N_19722,N_19558,N_19564);
and U19723 (N_19723,N_19470,N_19573);
nor U19724 (N_19724,N_19553,N_19556);
nand U19725 (N_19725,N_19427,N_19449);
and U19726 (N_19726,N_19426,N_19443);
xnor U19727 (N_19727,N_19415,N_19421);
or U19728 (N_19728,N_19417,N_19425);
and U19729 (N_19729,N_19583,N_19430);
nor U19730 (N_19730,N_19419,N_19416);
nand U19731 (N_19731,N_19489,N_19587);
nor U19732 (N_19732,N_19570,N_19446);
and U19733 (N_19733,N_19425,N_19520);
xnor U19734 (N_19734,N_19537,N_19527);
xnor U19735 (N_19735,N_19490,N_19459);
and U19736 (N_19736,N_19527,N_19578);
or U19737 (N_19737,N_19413,N_19401);
xnor U19738 (N_19738,N_19473,N_19552);
nand U19739 (N_19739,N_19414,N_19469);
and U19740 (N_19740,N_19449,N_19471);
and U19741 (N_19741,N_19596,N_19480);
nand U19742 (N_19742,N_19451,N_19501);
or U19743 (N_19743,N_19557,N_19512);
or U19744 (N_19744,N_19499,N_19408);
xnor U19745 (N_19745,N_19419,N_19411);
or U19746 (N_19746,N_19567,N_19441);
nor U19747 (N_19747,N_19449,N_19526);
xor U19748 (N_19748,N_19544,N_19573);
or U19749 (N_19749,N_19463,N_19510);
xnor U19750 (N_19750,N_19587,N_19554);
nor U19751 (N_19751,N_19410,N_19503);
nor U19752 (N_19752,N_19546,N_19545);
nand U19753 (N_19753,N_19576,N_19593);
nand U19754 (N_19754,N_19503,N_19413);
nor U19755 (N_19755,N_19542,N_19445);
and U19756 (N_19756,N_19421,N_19502);
xor U19757 (N_19757,N_19408,N_19537);
nor U19758 (N_19758,N_19425,N_19461);
or U19759 (N_19759,N_19404,N_19580);
nor U19760 (N_19760,N_19532,N_19540);
or U19761 (N_19761,N_19555,N_19574);
or U19762 (N_19762,N_19514,N_19558);
nand U19763 (N_19763,N_19538,N_19456);
and U19764 (N_19764,N_19442,N_19461);
or U19765 (N_19765,N_19538,N_19587);
xor U19766 (N_19766,N_19526,N_19518);
nor U19767 (N_19767,N_19461,N_19560);
or U19768 (N_19768,N_19425,N_19458);
nor U19769 (N_19769,N_19428,N_19425);
and U19770 (N_19770,N_19512,N_19580);
and U19771 (N_19771,N_19571,N_19411);
nand U19772 (N_19772,N_19423,N_19566);
nor U19773 (N_19773,N_19533,N_19447);
xor U19774 (N_19774,N_19494,N_19572);
xor U19775 (N_19775,N_19545,N_19535);
or U19776 (N_19776,N_19586,N_19468);
nand U19777 (N_19777,N_19418,N_19408);
or U19778 (N_19778,N_19443,N_19477);
nor U19779 (N_19779,N_19546,N_19544);
nor U19780 (N_19780,N_19451,N_19496);
xnor U19781 (N_19781,N_19423,N_19544);
xor U19782 (N_19782,N_19467,N_19441);
nand U19783 (N_19783,N_19531,N_19499);
xnor U19784 (N_19784,N_19533,N_19535);
nand U19785 (N_19785,N_19487,N_19512);
xor U19786 (N_19786,N_19586,N_19430);
or U19787 (N_19787,N_19597,N_19406);
xnor U19788 (N_19788,N_19596,N_19440);
nor U19789 (N_19789,N_19486,N_19410);
xor U19790 (N_19790,N_19448,N_19583);
nor U19791 (N_19791,N_19456,N_19406);
nor U19792 (N_19792,N_19518,N_19564);
and U19793 (N_19793,N_19572,N_19581);
nand U19794 (N_19794,N_19561,N_19568);
or U19795 (N_19795,N_19544,N_19489);
or U19796 (N_19796,N_19595,N_19511);
and U19797 (N_19797,N_19477,N_19582);
xor U19798 (N_19798,N_19506,N_19520);
nand U19799 (N_19799,N_19469,N_19504);
xor U19800 (N_19800,N_19720,N_19612);
nor U19801 (N_19801,N_19771,N_19774);
nor U19802 (N_19802,N_19687,N_19668);
nor U19803 (N_19803,N_19615,N_19752);
nand U19804 (N_19804,N_19766,N_19762);
and U19805 (N_19805,N_19734,N_19730);
nor U19806 (N_19806,N_19627,N_19735);
or U19807 (N_19807,N_19650,N_19791);
and U19808 (N_19808,N_19649,N_19754);
or U19809 (N_19809,N_19708,N_19608);
xor U19810 (N_19810,N_19672,N_19736);
or U19811 (N_19811,N_19661,N_19698);
nor U19812 (N_19812,N_19799,N_19633);
nor U19813 (N_19813,N_19757,N_19782);
nand U19814 (N_19814,N_19689,N_19658);
xor U19815 (N_19815,N_19677,N_19636);
or U19816 (N_19816,N_19699,N_19745);
nor U19817 (N_19817,N_19613,N_19713);
and U19818 (N_19818,N_19670,N_19755);
nor U19819 (N_19819,N_19690,N_19739);
nor U19820 (N_19820,N_19751,N_19606);
nor U19821 (N_19821,N_19785,N_19674);
or U19822 (N_19822,N_19623,N_19767);
xor U19823 (N_19823,N_19628,N_19645);
or U19824 (N_19824,N_19748,N_19728);
xor U19825 (N_19825,N_19700,N_19776);
nand U19826 (N_19826,N_19692,N_19789);
or U19827 (N_19827,N_19760,N_19753);
xor U19828 (N_19828,N_19683,N_19669);
nor U19829 (N_19829,N_19733,N_19746);
and U19830 (N_19830,N_19644,N_19701);
xor U19831 (N_19831,N_19702,N_19775);
and U19832 (N_19832,N_19703,N_19626);
or U19833 (N_19833,N_19717,N_19664);
xor U19834 (N_19834,N_19639,N_19707);
nand U19835 (N_19835,N_19617,N_19679);
and U19836 (N_19836,N_19647,N_19779);
or U19837 (N_19837,N_19624,N_19662);
nand U19838 (N_19838,N_19678,N_19769);
or U19839 (N_19839,N_19686,N_19709);
nand U19840 (N_19840,N_19660,N_19749);
xor U19841 (N_19841,N_19625,N_19609);
or U19842 (N_19842,N_19648,N_19607);
xnor U19843 (N_19843,N_19667,N_19721);
nand U19844 (N_19844,N_19693,N_19764);
xnor U19845 (N_19845,N_19632,N_19792);
and U19846 (N_19846,N_19696,N_19705);
and U19847 (N_19847,N_19656,N_19605);
nor U19848 (N_19848,N_19681,N_19742);
xor U19849 (N_19849,N_19768,N_19653);
and U19850 (N_19850,N_19604,N_19714);
and U19851 (N_19851,N_19795,N_19652);
xnor U19852 (N_19852,N_19716,N_19727);
or U19853 (N_19853,N_19732,N_19726);
xor U19854 (N_19854,N_19706,N_19618);
xor U19855 (N_19855,N_19747,N_19646);
nor U19856 (N_19856,N_19603,N_19614);
nor U19857 (N_19857,N_19723,N_19621);
xnor U19858 (N_19858,N_19600,N_19725);
nor U19859 (N_19859,N_19655,N_19796);
nor U19860 (N_19860,N_19622,N_19790);
nor U19861 (N_19861,N_19759,N_19772);
nor U19862 (N_19862,N_19629,N_19634);
or U19863 (N_19863,N_19631,N_19688);
xnor U19864 (N_19864,N_19610,N_19680);
or U19865 (N_19865,N_19654,N_19763);
nand U19866 (N_19866,N_19743,N_19740);
xor U19867 (N_19867,N_19694,N_19741);
and U19868 (N_19868,N_19616,N_19640);
and U19869 (N_19869,N_19673,N_19781);
nand U19870 (N_19870,N_19750,N_19601);
and U19871 (N_19871,N_19758,N_19697);
and U19872 (N_19872,N_19710,N_19641);
xor U19873 (N_19873,N_19620,N_19780);
xor U19874 (N_19874,N_19685,N_19676);
and U19875 (N_19875,N_19611,N_19637);
nand U19876 (N_19876,N_19793,N_19675);
or U19877 (N_19877,N_19798,N_19719);
nand U19878 (N_19878,N_19712,N_19715);
nor U19879 (N_19879,N_19756,N_19704);
and U19880 (N_19880,N_19695,N_19744);
or U19881 (N_19881,N_19738,N_19643);
nor U19882 (N_19882,N_19729,N_19666);
nand U19883 (N_19883,N_19665,N_19671);
nor U19884 (N_19884,N_19635,N_19619);
and U19885 (N_19885,N_19602,N_19737);
xnor U19886 (N_19886,N_19783,N_19794);
xnor U19887 (N_19887,N_19651,N_19797);
xor U19888 (N_19888,N_19765,N_19638);
xnor U19889 (N_19889,N_19787,N_19691);
xnor U19890 (N_19890,N_19684,N_19663);
xor U19891 (N_19891,N_19770,N_19724);
nand U19892 (N_19892,N_19682,N_19761);
and U19893 (N_19893,N_19642,N_19788);
or U19894 (N_19894,N_19786,N_19777);
and U19895 (N_19895,N_19718,N_19778);
nand U19896 (N_19896,N_19773,N_19711);
nand U19897 (N_19897,N_19722,N_19784);
nor U19898 (N_19898,N_19657,N_19630);
xnor U19899 (N_19899,N_19731,N_19659);
and U19900 (N_19900,N_19738,N_19663);
nor U19901 (N_19901,N_19720,N_19799);
and U19902 (N_19902,N_19698,N_19766);
nor U19903 (N_19903,N_19685,N_19657);
nand U19904 (N_19904,N_19719,N_19753);
or U19905 (N_19905,N_19766,N_19785);
or U19906 (N_19906,N_19716,N_19785);
nor U19907 (N_19907,N_19727,N_19693);
nor U19908 (N_19908,N_19761,N_19789);
or U19909 (N_19909,N_19763,N_19674);
nand U19910 (N_19910,N_19784,N_19707);
nand U19911 (N_19911,N_19760,N_19722);
xor U19912 (N_19912,N_19701,N_19721);
nand U19913 (N_19913,N_19793,N_19677);
and U19914 (N_19914,N_19746,N_19625);
xor U19915 (N_19915,N_19654,N_19749);
xnor U19916 (N_19916,N_19738,N_19677);
or U19917 (N_19917,N_19721,N_19634);
and U19918 (N_19918,N_19796,N_19725);
or U19919 (N_19919,N_19668,N_19767);
or U19920 (N_19920,N_19695,N_19678);
or U19921 (N_19921,N_19721,N_19734);
or U19922 (N_19922,N_19693,N_19766);
nor U19923 (N_19923,N_19774,N_19659);
and U19924 (N_19924,N_19624,N_19775);
nand U19925 (N_19925,N_19634,N_19786);
nand U19926 (N_19926,N_19600,N_19620);
or U19927 (N_19927,N_19626,N_19639);
nor U19928 (N_19928,N_19798,N_19641);
and U19929 (N_19929,N_19770,N_19756);
xnor U19930 (N_19930,N_19700,N_19748);
nor U19931 (N_19931,N_19714,N_19757);
xor U19932 (N_19932,N_19759,N_19793);
xor U19933 (N_19933,N_19643,N_19765);
nor U19934 (N_19934,N_19693,N_19714);
nand U19935 (N_19935,N_19788,N_19612);
nand U19936 (N_19936,N_19607,N_19714);
nor U19937 (N_19937,N_19790,N_19682);
xnor U19938 (N_19938,N_19636,N_19769);
and U19939 (N_19939,N_19797,N_19643);
and U19940 (N_19940,N_19624,N_19633);
or U19941 (N_19941,N_19621,N_19781);
nand U19942 (N_19942,N_19751,N_19735);
nor U19943 (N_19943,N_19791,N_19738);
or U19944 (N_19944,N_19750,N_19735);
and U19945 (N_19945,N_19636,N_19737);
nor U19946 (N_19946,N_19723,N_19636);
and U19947 (N_19947,N_19751,N_19628);
and U19948 (N_19948,N_19668,N_19729);
nand U19949 (N_19949,N_19689,N_19757);
xnor U19950 (N_19950,N_19784,N_19666);
xnor U19951 (N_19951,N_19769,N_19726);
and U19952 (N_19952,N_19647,N_19778);
nor U19953 (N_19953,N_19628,N_19650);
nand U19954 (N_19954,N_19628,N_19648);
nand U19955 (N_19955,N_19641,N_19605);
xor U19956 (N_19956,N_19695,N_19729);
nor U19957 (N_19957,N_19799,N_19628);
and U19958 (N_19958,N_19772,N_19760);
or U19959 (N_19959,N_19619,N_19674);
xnor U19960 (N_19960,N_19627,N_19652);
nand U19961 (N_19961,N_19792,N_19768);
xor U19962 (N_19962,N_19656,N_19706);
nand U19963 (N_19963,N_19720,N_19735);
nor U19964 (N_19964,N_19662,N_19777);
or U19965 (N_19965,N_19771,N_19660);
nor U19966 (N_19966,N_19629,N_19616);
nand U19967 (N_19967,N_19645,N_19618);
xnor U19968 (N_19968,N_19659,N_19623);
or U19969 (N_19969,N_19673,N_19625);
nand U19970 (N_19970,N_19741,N_19783);
nand U19971 (N_19971,N_19641,N_19655);
nand U19972 (N_19972,N_19612,N_19658);
nor U19973 (N_19973,N_19737,N_19616);
nand U19974 (N_19974,N_19629,N_19619);
nor U19975 (N_19975,N_19678,N_19720);
nand U19976 (N_19976,N_19622,N_19672);
xnor U19977 (N_19977,N_19789,N_19626);
nor U19978 (N_19978,N_19781,N_19717);
xor U19979 (N_19979,N_19761,N_19700);
nand U19980 (N_19980,N_19718,N_19688);
or U19981 (N_19981,N_19680,N_19712);
and U19982 (N_19982,N_19606,N_19798);
nand U19983 (N_19983,N_19747,N_19749);
nor U19984 (N_19984,N_19793,N_19734);
nor U19985 (N_19985,N_19642,N_19706);
nor U19986 (N_19986,N_19617,N_19621);
or U19987 (N_19987,N_19732,N_19784);
xor U19988 (N_19988,N_19652,N_19770);
nor U19989 (N_19989,N_19761,N_19777);
nand U19990 (N_19990,N_19613,N_19629);
nor U19991 (N_19991,N_19732,N_19671);
xnor U19992 (N_19992,N_19793,N_19624);
or U19993 (N_19993,N_19645,N_19663);
or U19994 (N_19994,N_19610,N_19769);
nor U19995 (N_19995,N_19779,N_19615);
nand U19996 (N_19996,N_19790,N_19799);
nand U19997 (N_19997,N_19665,N_19703);
or U19998 (N_19998,N_19612,N_19764);
and U19999 (N_19999,N_19642,N_19777);
xor U20000 (N_20000,N_19931,N_19918);
nor U20001 (N_20001,N_19827,N_19988);
xnor U20002 (N_20002,N_19881,N_19889);
nand U20003 (N_20003,N_19924,N_19857);
and U20004 (N_20004,N_19993,N_19958);
nor U20005 (N_20005,N_19899,N_19966);
nor U20006 (N_20006,N_19987,N_19840);
nand U20007 (N_20007,N_19922,N_19850);
xnor U20008 (N_20008,N_19878,N_19858);
nand U20009 (N_20009,N_19900,N_19983);
xnor U20010 (N_20010,N_19872,N_19930);
nand U20011 (N_20011,N_19933,N_19945);
nand U20012 (N_20012,N_19898,N_19928);
xor U20013 (N_20013,N_19916,N_19940);
xor U20014 (N_20014,N_19822,N_19883);
xnor U20015 (N_20015,N_19960,N_19825);
nor U20016 (N_20016,N_19910,N_19861);
nand U20017 (N_20017,N_19819,N_19909);
xnor U20018 (N_20018,N_19920,N_19813);
and U20019 (N_20019,N_19886,N_19999);
or U20020 (N_20020,N_19882,N_19994);
nand U20021 (N_20021,N_19908,N_19978);
nand U20022 (N_20022,N_19851,N_19831);
and U20023 (N_20023,N_19811,N_19856);
or U20024 (N_20024,N_19895,N_19890);
or U20025 (N_20025,N_19997,N_19874);
xor U20026 (N_20026,N_19863,N_19849);
and U20027 (N_20027,N_19996,N_19842);
nand U20028 (N_20028,N_19864,N_19961);
xnor U20029 (N_20029,N_19954,N_19912);
and U20030 (N_20030,N_19968,N_19855);
and U20031 (N_20031,N_19880,N_19963);
nand U20032 (N_20032,N_19977,N_19824);
nand U20033 (N_20033,N_19917,N_19875);
nor U20034 (N_20034,N_19845,N_19816);
xor U20035 (N_20035,N_19995,N_19852);
and U20036 (N_20036,N_19873,N_19906);
xor U20037 (N_20037,N_19932,N_19943);
and U20038 (N_20038,N_19990,N_19938);
and U20039 (N_20039,N_19870,N_19967);
or U20040 (N_20040,N_19979,N_19893);
nand U20041 (N_20041,N_19804,N_19809);
nor U20042 (N_20042,N_19927,N_19843);
and U20043 (N_20043,N_19803,N_19826);
xnor U20044 (N_20044,N_19936,N_19948);
and U20045 (N_20045,N_19903,N_19876);
xor U20046 (N_20046,N_19833,N_19911);
and U20047 (N_20047,N_19934,N_19965);
or U20048 (N_20048,N_19981,N_19853);
nand U20049 (N_20049,N_19854,N_19986);
nand U20050 (N_20050,N_19865,N_19859);
nand U20051 (N_20051,N_19946,N_19836);
nand U20052 (N_20052,N_19925,N_19947);
and U20053 (N_20053,N_19941,N_19835);
nand U20054 (N_20054,N_19974,N_19976);
nand U20055 (N_20055,N_19829,N_19952);
or U20056 (N_20056,N_19959,N_19964);
xor U20057 (N_20057,N_19805,N_19820);
nor U20058 (N_20058,N_19888,N_19926);
or U20059 (N_20059,N_19894,N_19998);
and U20060 (N_20060,N_19973,N_19862);
xor U20061 (N_20061,N_19812,N_19923);
and U20062 (N_20062,N_19807,N_19884);
and U20063 (N_20063,N_19935,N_19839);
nand U20064 (N_20064,N_19971,N_19985);
xor U20065 (N_20065,N_19972,N_19830);
xor U20066 (N_20066,N_19866,N_19837);
or U20067 (N_20067,N_19919,N_19846);
and U20068 (N_20068,N_19953,N_19885);
or U20069 (N_20069,N_19950,N_19848);
or U20070 (N_20070,N_19970,N_19817);
xor U20071 (N_20071,N_19834,N_19991);
nor U20072 (N_20072,N_19832,N_19907);
xor U20073 (N_20073,N_19871,N_19942);
or U20074 (N_20074,N_19868,N_19828);
nand U20075 (N_20075,N_19821,N_19955);
and U20076 (N_20076,N_19867,N_19980);
xnor U20077 (N_20077,N_19975,N_19914);
nand U20078 (N_20078,N_19841,N_19808);
nor U20079 (N_20079,N_19891,N_19814);
nand U20080 (N_20080,N_19929,N_19844);
xor U20081 (N_20081,N_19962,N_19957);
or U20082 (N_20082,N_19984,N_19887);
nor U20083 (N_20083,N_19800,N_19847);
and U20084 (N_20084,N_19921,N_19823);
xor U20085 (N_20085,N_19806,N_19897);
nor U20086 (N_20086,N_19869,N_19892);
and U20087 (N_20087,N_19810,N_19838);
nor U20088 (N_20088,N_19901,N_19905);
or U20089 (N_20089,N_19818,N_19877);
nand U20090 (N_20090,N_19802,N_19815);
nor U20091 (N_20091,N_19939,N_19915);
nand U20092 (N_20092,N_19937,N_19904);
and U20093 (N_20093,N_19913,N_19896);
nor U20094 (N_20094,N_19860,N_19879);
and U20095 (N_20095,N_19956,N_19982);
nand U20096 (N_20096,N_19801,N_19992);
and U20097 (N_20097,N_19902,N_19969);
nand U20098 (N_20098,N_19944,N_19989);
xnor U20099 (N_20099,N_19951,N_19949);
nor U20100 (N_20100,N_19872,N_19808);
and U20101 (N_20101,N_19832,N_19838);
nor U20102 (N_20102,N_19937,N_19944);
and U20103 (N_20103,N_19947,N_19866);
or U20104 (N_20104,N_19894,N_19831);
nor U20105 (N_20105,N_19810,N_19931);
nor U20106 (N_20106,N_19980,N_19834);
nand U20107 (N_20107,N_19992,N_19943);
xnor U20108 (N_20108,N_19830,N_19856);
xnor U20109 (N_20109,N_19904,N_19983);
or U20110 (N_20110,N_19926,N_19965);
nand U20111 (N_20111,N_19839,N_19921);
nand U20112 (N_20112,N_19954,N_19902);
and U20113 (N_20113,N_19892,N_19896);
or U20114 (N_20114,N_19835,N_19977);
or U20115 (N_20115,N_19944,N_19951);
or U20116 (N_20116,N_19820,N_19899);
xor U20117 (N_20117,N_19963,N_19855);
or U20118 (N_20118,N_19837,N_19889);
nand U20119 (N_20119,N_19844,N_19912);
and U20120 (N_20120,N_19994,N_19988);
and U20121 (N_20121,N_19990,N_19953);
nand U20122 (N_20122,N_19913,N_19828);
nand U20123 (N_20123,N_19862,N_19923);
xor U20124 (N_20124,N_19837,N_19924);
and U20125 (N_20125,N_19954,N_19932);
nand U20126 (N_20126,N_19930,N_19960);
or U20127 (N_20127,N_19834,N_19921);
nand U20128 (N_20128,N_19927,N_19813);
nand U20129 (N_20129,N_19910,N_19813);
and U20130 (N_20130,N_19975,N_19953);
xor U20131 (N_20131,N_19864,N_19804);
nor U20132 (N_20132,N_19979,N_19904);
nand U20133 (N_20133,N_19952,N_19813);
nand U20134 (N_20134,N_19856,N_19916);
or U20135 (N_20135,N_19800,N_19877);
xor U20136 (N_20136,N_19978,N_19940);
and U20137 (N_20137,N_19825,N_19964);
or U20138 (N_20138,N_19834,N_19955);
nor U20139 (N_20139,N_19999,N_19900);
nand U20140 (N_20140,N_19937,N_19905);
xor U20141 (N_20141,N_19983,N_19909);
nand U20142 (N_20142,N_19940,N_19855);
nor U20143 (N_20143,N_19918,N_19925);
nor U20144 (N_20144,N_19863,N_19941);
nor U20145 (N_20145,N_19955,N_19861);
nor U20146 (N_20146,N_19806,N_19939);
xor U20147 (N_20147,N_19804,N_19922);
nand U20148 (N_20148,N_19905,N_19875);
or U20149 (N_20149,N_19948,N_19898);
nor U20150 (N_20150,N_19912,N_19998);
and U20151 (N_20151,N_19950,N_19826);
xnor U20152 (N_20152,N_19808,N_19925);
xor U20153 (N_20153,N_19870,N_19950);
nand U20154 (N_20154,N_19848,N_19836);
nand U20155 (N_20155,N_19803,N_19938);
and U20156 (N_20156,N_19983,N_19994);
nor U20157 (N_20157,N_19885,N_19987);
nor U20158 (N_20158,N_19865,N_19839);
and U20159 (N_20159,N_19846,N_19885);
xnor U20160 (N_20160,N_19933,N_19904);
xor U20161 (N_20161,N_19829,N_19854);
nand U20162 (N_20162,N_19867,N_19943);
nand U20163 (N_20163,N_19916,N_19997);
or U20164 (N_20164,N_19812,N_19927);
or U20165 (N_20165,N_19969,N_19813);
and U20166 (N_20166,N_19924,N_19960);
nor U20167 (N_20167,N_19895,N_19910);
nand U20168 (N_20168,N_19900,N_19923);
nand U20169 (N_20169,N_19912,N_19934);
and U20170 (N_20170,N_19884,N_19816);
and U20171 (N_20171,N_19910,N_19950);
and U20172 (N_20172,N_19995,N_19991);
xnor U20173 (N_20173,N_19800,N_19911);
and U20174 (N_20174,N_19853,N_19885);
xor U20175 (N_20175,N_19985,N_19855);
nand U20176 (N_20176,N_19924,N_19885);
nand U20177 (N_20177,N_19949,N_19987);
nor U20178 (N_20178,N_19861,N_19984);
nor U20179 (N_20179,N_19973,N_19883);
nor U20180 (N_20180,N_19973,N_19801);
or U20181 (N_20181,N_19898,N_19945);
and U20182 (N_20182,N_19984,N_19802);
and U20183 (N_20183,N_19926,N_19951);
xnor U20184 (N_20184,N_19858,N_19819);
and U20185 (N_20185,N_19908,N_19897);
or U20186 (N_20186,N_19989,N_19859);
or U20187 (N_20187,N_19807,N_19804);
nand U20188 (N_20188,N_19998,N_19989);
xor U20189 (N_20189,N_19860,N_19943);
nor U20190 (N_20190,N_19975,N_19847);
xnor U20191 (N_20191,N_19902,N_19997);
or U20192 (N_20192,N_19872,N_19800);
or U20193 (N_20193,N_19943,N_19895);
and U20194 (N_20194,N_19913,N_19916);
nand U20195 (N_20195,N_19824,N_19949);
nor U20196 (N_20196,N_19955,N_19971);
xnor U20197 (N_20197,N_19802,N_19857);
nand U20198 (N_20198,N_19869,N_19807);
xnor U20199 (N_20199,N_19982,N_19822);
and U20200 (N_20200,N_20162,N_20038);
nor U20201 (N_20201,N_20022,N_20139);
or U20202 (N_20202,N_20175,N_20024);
or U20203 (N_20203,N_20133,N_20153);
xnor U20204 (N_20204,N_20183,N_20116);
or U20205 (N_20205,N_20036,N_20051);
xnor U20206 (N_20206,N_20002,N_20121);
nand U20207 (N_20207,N_20098,N_20012);
nand U20208 (N_20208,N_20145,N_20006);
nand U20209 (N_20209,N_20196,N_20021);
nor U20210 (N_20210,N_20168,N_20041);
or U20211 (N_20211,N_20099,N_20026);
or U20212 (N_20212,N_20135,N_20105);
nor U20213 (N_20213,N_20078,N_20046);
xnor U20214 (N_20214,N_20010,N_20195);
and U20215 (N_20215,N_20123,N_20074);
and U20216 (N_20216,N_20190,N_20072);
or U20217 (N_20217,N_20114,N_20065);
and U20218 (N_20218,N_20048,N_20068);
nand U20219 (N_20219,N_20113,N_20148);
or U20220 (N_20220,N_20188,N_20060);
nand U20221 (N_20221,N_20025,N_20126);
or U20222 (N_20222,N_20134,N_20193);
nor U20223 (N_20223,N_20144,N_20140);
xor U20224 (N_20224,N_20111,N_20043);
and U20225 (N_20225,N_20035,N_20191);
or U20226 (N_20226,N_20198,N_20131);
nor U20227 (N_20227,N_20056,N_20174);
xor U20228 (N_20228,N_20164,N_20054);
xor U20229 (N_20229,N_20128,N_20080);
or U20230 (N_20230,N_20184,N_20057);
and U20231 (N_20231,N_20094,N_20152);
or U20232 (N_20232,N_20015,N_20163);
xnor U20233 (N_20233,N_20138,N_20008);
nor U20234 (N_20234,N_20049,N_20085);
nand U20235 (N_20235,N_20079,N_20023);
or U20236 (N_20236,N_20030,N_20161);
xor U20237 (N_20237,N_20101,N_20180);
nor U20238 (N_20238,N_20125,N_20004);
nor U20239 (N_20239,N_20115,N_20013);
nor U20240 (N_20240,N_20171,N_20141);
xnor U20241 (N_20241,N_20118,N_20100);
nand U20242 (N_20242,N_20042,N_20146);
or U20243 (N_20243,N_20084,N_20058);
nand U20244 (N_20244,N_20076,N_20073);
nor U20245 (N_20245,N_20071,N_20095);
nor U20246 (N_20246,N_20097,N_20005);
nor U20247 (N_20247,N_20032,N_20077);
and U20248 (N_20248,N_20062,N_20155);
and U20249 (N_20249,N_20143,N_20092);
and U20250 (N_20250,N_20103,N_20039);
xnor U20251 (N_20251,N_20102,N_20189);
nor U20252 (N_20252,N_20093,N_20044);
nor U20253 (N_20253,N_20059,N_20127);
and U20254 (N_20254,N_20052,N_20082);
nor U20255 (N_20255,N_20187,N_20086);
or U20256 (N_20256,N_20173,N_20063);
nand U20257 (N_20257,N_20177,N_20176);
or U20258 (N_20258,N_20090,N_20003);
and U20259 (N_20259,N_20107,N_20083);
xor U20260 (N_20260,N_20050,N_20147);
or U20261 (N_20261,N_20066,N_20150);
nand U20262 (N_20262,N_20064,N_20170);
nand U20263 (N_20263,N_20027,N_20061);
or U20264 (N_20264,N_20199,N_20165);
or U20265 (N_20265,N_20089,N_20047);
nand U20266 (N_20266,N_20104,N_20166);
and U20267 (N_20267,N_20034,N_20136);
or U20268 (N_20268,N_20108,N_20186);
and U20269 (N_20269,N_20182,N_20001);
xor U20270 (N_20270,N_20017,N_20132);
nor U20271 (N_20271,N_20055,N_20167);
xnor U20272 (N_20272,N_20122,N_20124);
nor U20273 (N_20273,N_20119,N_20037);
or U20274 (N_20274,N_20053,N_20181);
xnor U20275 (N_20275,N_20007,N_20009);
nor U20276 (N_20276,N_20197,N_20075);
nand U20277 (N_20277,N_20019,N_20045);
and U20278 (N_20278,N_20156,N_20172);
and U20279 (N_20279,N_20011,N_20129);
or U20280 (N_20280,N_20154,N_20081);
or U20281 (N_20281,N_20142,N_20106);
or U20282 (N_20282,N_20033,N_20110);
nor U20283 (N_20283,N_20028,N_20149);
nor U20284 (N_20284,N_20020,N_20088);
nor U20285 (N_20285,N_20159,N_20117);
xor U20286 (N_20286,N_20169,N_20137);
or U20287 (N_20287,N_20109,N_20112);
xor U20288 (N_20288,N_20192,N_20178);
xor U20289 (N_20289,N_20018,N_20070);
nand U20290 (N_20290,N_20069,N_20091);
nor U20291 (N_20291,N_20087,N_20157);
or U20292 (N_20292,N_20096,N_20185);
nor U20293 (N_20293,N_20130,N_20194);
nor U20294 (N_20294,N_20151,N_20016);
or U20295 (N_20295,N_20160,N_20031);
and U20296 (N_20296,N_20029,N_20120);
xnor U20297 (N_20297,N_20067,N_20179);
and U20298 (N_20298,N_20158,N_20000);
nand U20299 (N_20299,N_20040,N_20014);
and U20300 (N_20300,N_20076,N_20149);
nor U20301 (N_20301,N_20022,N_20151);
nor U20302 (N_20302,N_20163,N_20012);
xor U20303 (N_20303,N_20013,N_20153);
nand U20304 (N_20304,N_20124,N_20048);
xor U20305 (N_20305,N_20006,N_20128);
and U20306 (N_20306,N_20142,N_20140);
nand U20307 (N_20307,N_20002,N_20184);
and U20308 (N_20308,N_20157,N_20163);
or U20309 (N_20309,N_20157,N_20068);
nand U20310 (N_20310,N_20076,N_20140);
and U20311 (N_20311,N_20048,N_20163);
xor U20312 (N_20312,N_20133,N_20080);
and U20313 (N_20313,N_20111,N_20085);
and U20314 (N_20314,N_20019,N_20173);
nor U20315 (N_20315,N_20099,N_20100);
nand U20316 (N_20316,N_20019,N_20050);
nor U20317 (N_20317,N_20083,N_20044);
and U20318 (N_20318,N_20077,N_20028);
nand U20319 (N_20319,N_20197,N_20172);
nor U20320 (N_20320,N_20006,N_20001);
nand U20321 (N_20321,N_20034,N_20029);
xnor U20322 (N_20322,N_20023,N_20085);
xor U20323 (N_20323,N_20186,N_20085);
and U20324 (N_20324,N_20027,N_20170);
and U20325 (N_20325,N_20149,N_20163);
xor U20326 (N_20326,N_20068,N_20152);
or U20327 (N_20327,N_20066,N_20181);
and U20328 (N_20328,N_20091,N_20186);
nor U20329 (N_20329,N_20037,N_20065);
and U20330 (N_20330,N_20082,N_20019);
and U20331 (N_20331,N_20149,N_20009);
nand U20332 (N_20332,N_20172,N_20127);
nor U20333 (N_20333,N_20051,N_20184);
and U20334 (N_20334,N_20025,N_20006);
and U20335 (N_20335,N_20087,N_20053);
nor U20336 (N_20336,N_20188,N_20028);
nor U20337 (N_20337,N_20140,N_20064);
nand U20338 (N_20338,N_20073,N_20006);
nor U20339 (N_20339,N_20103,N_20159);
xnor U20340 (N_20340,N_20121,N_20014);
or U20341 (N_20341,N_20104,N_20193);
and U20342 (N_20342,N_20065,N_20144);
nand U20343 (N_20343,N_20196,N_20045);
nand U20344 (N_20344,N_20150,N_20031);
and U20345 (N_20345,N_20091,N_20183);
and U20346 (N_20346,N_20130,N_20084);
or U20347 (N_20347,N_20077,N_20064);
or U20348 (N_20348,N_20176,N_20025);
nor U20349 (N_20349,N_20155,N_20160);
xor U20350 (N_20350,N_20070,N_20040);
nand U20351 (N_20351,N_20060,N_20117);
and U20352 (N_20352,N_20113,N_20098);
and U20353 (N_20353,N_20158,N_20098);
or U20354 (N_20354,N_20106,N_20144);
and U20355 (N_20355,N_20061,N_20197);
xnor U20356 (N_20356,N_20164,N_20038);
nor U20357 (N_20357,N_20071,N_20058);
and U20358 (N_20358,N_20138,N_20130);
nand U20359 (N_20359,N_20145,N_20012);
and U20360 (N_20360,N_20162,N_20087);
and U20361 (N_20361,N_20049,N_20061);
nand U20362 (N_20362,N_20187,N_20001);
xnor U20363 (N_20363,N_20110,N_20159);
xnor U20364 (N_20364,N_20117,N_20004);
nand U20365 (N_20365,N_20042,N_20029);
xor U20366 (N_20366,N_20177,N_20088);
nor U20367 (N_20367,N_20104,N_20027);
nand U20368 (N_20368,N_20091,N_20198);
nor U20369 (N_20369,N_20129,N_20022);
xnor U20370 (N_20370,N_20020,N_20028);
xnor U20371 (N_20371,N_20025,N_20197);
and U20372 (N_20372,N_20157,N_20135);
or U20373 (N_20373,N_20146,N_20128);
xnor U20374 (N_20374,N_20140,N_20039);
xor U20375 (N_20375,N_20151,N_20057);
or U20376 (N_20376,N_20159,N_20154);
and U20377 (N_20377,N_20171,N_20056);
xor U20378 (N_20378,N_20033,N_20060);
and U20379 (N_20379,N_20141,N_20172);
or U20380 (N_20380,N_20144,N_20043);
xor U20381 (N_20381,N_20130,N_20142);
nor U20382 (N_20382,N_20080,N_20091);
nor U20383 (N_20383,N_20111,N_20185);
or U20384 (N_20384,N_20196,N_20126);
xnor U20385 (N_20385,N_20130,N_20105);
nor U20386 (N_20386,N_20136,N_20006);
nand U20387 (N_20387,N_20011,N_20137);
nor U20388 (N_20388,N_20103,N_20109);
xor U20389 (N_20389,N_20047,N_20022);
and U20390 (N_20390,N_20075,N_20010);
nand U20391 (N_20391,N_20114,N_20075);
xor U20392 (N_20392,N_20015,N_20121);
nor U20393 (N_20393,N_20122,N_20085);
and U20394 (N_20394,N_20086,N_20135);
and U20395 (N_20395,N_20132,N_20099);
xor U20396 (N_20396,N_20106,N_20019);
or U20397 (N_20397,N_20169,N_20016);
and U20398 (N_20398,N_20120,N_20146);
or U20399 (N_20399,N_20127,N_20179);
and U20400 (N_20400,N_20369,N_20312);
nand U20401 (N_20401,N_20387,N_20364);
and U20402 (N_20402,N_20357,N_20338);
xnor U20403 (N_20403,N_20230,N_20318);
nand U20404 (N_20404,N_20297,N_20212);
or U20405 (N_20405,N_20295,N_20215);
or U20406 (N_20406,N_20375,N_20384);
or U20407 (N_20407,N_20213,N_20388);
nand U20408 (N_20408,N_20315,N_20352);
or U20409 (N_20409,N_20272,N_20285);
and U20410 (N_20410,N_20282,N_20235);
or U20411 (N_20411,N_20380,N_20217);
nor U20412 (N_20412,N_20370,N_20311);
nand U20413 (N_20413,N_20309,N_20374);
xor U20414 (N_20414,N_20392,N_20216);
or U20415 (N_20415,N_20344,N_20314);
xnor U20416 (N_20416,N_20317,N_20365);
xnor U20417 (N_20417,N_20367,N_20274);
and U20418 (N_20418,N_20305,N_20381);
or U20419 (N_20419,N_20225,N_20292);
xnor U20420 (N_20420,N_20332,N_20334);
xor U20421 (N_20421,N_20356,N_20228);
nor U20422 (N_20422,N_20277,N_20345);
or U20423 (N_20423,N_20249,N_20383);
nand U20424 (N_20424,N_20267,N_20266);
nor U20425 (N_20425,N_20320,N_20244);
nand U20426 (N_20426,N_20296,N_20303);
or U20427 (N_20427,N_20399,N_20385);
or U20428 (N_20428,N_20302,N_20233);
and U20429 (N_20429,N_20218,N_20358);
nor U20430 (N_20430,N_20264,N_20382);
and U20431 (N_20431,N_20286,N_20354);
and U20432 (N_20432,N_20340,N_20263);
or U20433 (N_20433,N_20265,N_20372);
xor U20434 (N_20434,N_20227,N_20321);
nor U20435 (N_20435,N_20278,N_20214);
and U20436 (N_20436,N_20223,N_20243);
and U20437 (N_20437,N_20280,N_20211);
xor U20438 (N_20438,N_20323,N_20289);
nor U20439 (N_20439,N_20329,N_20205);
and U20440 (N_20440,N_20240,N_20396);
xnor U20441 (N_20441,N_20208,N_20248);
xnor U20442 (N_20442,N_20262,N_20234);
nor U20443 (N_20443,N_20333,N_20341);
nor U20444 (N_20444,N_20390,N_20226);
or U20445 (N_20445,N_20232,N_20336);
nor U20446 (N_20446,N_20253,N_20347);
xor U20447 (N_20447,N_20252,N_20238);
xor U20448 (N_20448,N_20247,N_20306);
nor U20449 (N_20449,N_20319,N_20326);
and U20450 (N_20450,N_20255,N_20281);
nor U20451 (N_20451,N_20254,N_20207);
xor U20452 (N_20452,N_20299,N_20220);
nor U20453 (N_20453,N_20209,N_20376);
xor U20454 (N_20454,N_20201,N_20391);
or U20455 (N_20455,N_20346,N_20276);
and U20456 (N_20456,N_20393,N_20293);
nor U20457 (N_20457,N_20246,N_20337);
or U20458 (N_20458,N_20298,N_20219);
and U20459 (N_20459,N_20342,N_20222);
nor U20460 (N_20460,N_20327,N_20386);
nand U20461 (N_20461,N_20398,N_20287);
nand U20462 (N_20462,N_20202,N_20245);
nand U20463 (N_20463,N_20324,N_20339);
or U20464 (N_20464,N_20310,N_20283);
xor U20465 (N_20465,N_20368,N_20394);
nor U20466 (N_20466,N_20268,N_20275);
nand U20467 (N_20467,N_20269,N_20322);
nand U20468 (N_20468,N_20359,N_20273);
nand U20469 (N_20469,N_20229,N_20343);
or U20470 (N_20470,N_20378,N_20325);
or U20471 (N_20471,N_20236,N_20397);
or U20472 (N_20472,N_20328,N_20373);
or U20473 (N_20473,N_20256,N_20294);
or U20474 (N_20474,N_20350,N_20271);
or U20475 (N_20475,N_20361,N_20284);
and U20476 (N_20476,N_20379,N_20316);
xnor U20477 (N_20477,N_20308,N_20251);
nand U20478 (N_20478,N_20362,N_20301);
xnor U20479 (N_20479,N_20389,N_20363);
nand U20480 (N_20480,N_20291,N_20313);
or U20481 (N_20481,N_20204,N_20351);
nor U20482 (N_20482,N_20250,N_20237);
and U20483 (N_20483,N_20259,N_20331);
xor U20484 (N_20484,N_20206,N_20371);
or U20485 (N_20485,N_20258,N_20221);
nand U20486 (N_20486,N_20360,N_20231);
nor U20487 (N_20487,N_20366,N_20307);
xor U20488 (N_20488,N_20348,N_20239);
nor U20489 (N_20489,N_20290,N_20300);
nand U20490 (N_20490,N_20353,N_20279);
nor U20491 (N_20491,N_20200,N_20210);
and U20492 (N_20492,N_20288,N_20261);
xor U20493 (N_20493,N_20203,N_20377);
nand U20494 (N_20494,N_20260,N_20395);
nor U20495 (N_20495,N_20224,N_20257);
xor U20496 (N_20496,N_20349,N_20242);
and U20497 (N_20497,N_20304,N_20330);
nand U20498 (N_20498,N_20270,N_20355);
and U20499 (N_20499,N_20241,N_20335);
nor U20500 (N_20500,N_20357,N_20255);
or U20501 (N_20501,N_20235,N_20391);
or U20502 (N_20502,N_20371,N_20351);
xor U20503 (N_20503,N_20234,N_20212);
nand U20504 (N_20504,N_20387,N_20305);
or U20505 (N_20505,N_20307,N_20355);
or U20506 (N_20506,N_20246,N_20308);
nor U20507 (N_20507,N_20384,N_20323);
xnor U20508 (N_20508,N_20232,N_20321);
or U20509 (N_20509,N_20325,N_20327);
or U20510 (N_20510,N_20249,N_20206);
xnor U20511 (N_20511,N_20227,N_20223);
and U20512 (N_20512,N_20206,N_20334);
and U20513 (N_20513,N_20337,N_20210);
or U20514 (N_20514,N_20318,N_20242);
or U20515 (N_20515,N_20246,N_20398);
xnor U20516 (N_20516,N_20348,N_20396);
and U20517 (N_20517,N_20206,N_20388);
xor U20518 (N_20518,N_20269,N_20290);
and U20519 (N_20519,N_20322,N_20357);
xnor U20520 (N_20520,N_20395,N_20333);
xnor U20521 (N_20521,N_20285,N_20344);
nand U20522 (N_20522,N_20212,N_20364);
or U20523 (N_20523,N_20306,N_20397);
xnor U20524 (N_20524,N_20302,N_20242);
and U20525 (N_20525,N_20269,N_20260);
and U20526 (N_20526,N_20262,N_20387);
xnor U20527 (N_20527,N_20318,N_20330);
nor U20528 (N_20528,N_20201,N_20226);
or U20529 (N_20529,N_20399,N_20204);
and U20530 (N_20530,N_20340,N_20352);
or U20531 (N_20531,N_20375,N_20224);
nand U20532 (N_20532,N_20337,N_20302);
nor U20533 (N_20533,N_20360,N_20268);
nand U20534 (N_20534,N_20349,N_20272);
nor U20535 (N_20535,N_20379,N_20372);
or U20536 (N_20536,N_20229,N_20277);
or U20537 (N_20537,N_20209,N_20297);
xnor U20538 (N_20538,N_20221,N_20369);
nor U20539 (N_20539,N_20226,N_20205);
xnor U20540 (N_20540,N_20262,N_20252);
nor U20541 (N_20541,N_20346,N_20371);
nor U20542 (N_20542,N_20240,N_20378);
and U20543 (N_20543,N_20374,N_20338);
or U20544 (N_20544,N_20349,N_20231);
and U20545 (N_20545,N_20307,N_20372);
and U20546 (N_20546,N_20371,N_20251);
or U20547 (N_20547,N_20251,N_20204);
and U20548 (N_20548,N_20279,N_20349);
or U20549 (N_20549,N_20326,N_20395);
and U20550 (N_20550,N_20218,N_20319);
nand U20551 (N_20551,N_20235,N_20327);
or U20552 (N_20552,N_20389,N_20314);
or U20553 (N_20553,N_20208,N_20225);
nor U20554 (N_20554,N_20211,N_20372);
nor U20555 (N_20555,N_20353,N_20262);
nor U20556 (N_20556,N_20334,N_20282);
xnor U20557 (N_20557,N_20320,N_20310);
or U20558 (N_20558,N_20323,N_20264);
and U20559 (N_20559,N_20233,N_20397);
or U20560 (N_20560,N_20348,N_20377);
and U20561 (N_20561,N_20217,N_20362);
nor U20562 (N_20562,N_20397,N_20280);
nand U20563 (N_20563,N_20207,N_20296);
or U20564 (N_20564,N_20249,N_20377);
or U20565 (N_20565,N_20272,N_20322);
or U20566 (N_20566,N_20342,N_20316);
nor U20567 (N_20567,N_20336,N_20262);
or U20568 (N_20568,N_20332,N_20221);
xor U20569 (N_20569,N_20257,N_20251);
nor U20570 (N_20570,N_20269,N_20238);
nand U20571 (N_20571,N_20378,N_20364);
nand U20572 (N_20572,N_20317,N_20378);
nor U20573 (N_20573,N_20215,N_20270);
nand U20574 (N_20574,N_20302,N_20235);
xnor U20575 (N_20575,N_20292,N_20224);
nand U20576 (N_20576,N_20318,N_20324);
nor U20577 (N_20577,N_20241,N_20216);
xor U20578 (N_20578,N_20288,N_20354);
or U20579 (N_20579,N_20212,N_20320);
or U20580 (N_20580,N_20326,N_20329);
xnor U20581 (N_20581,N_20229,N_20348);
and U20582 (N_20582,N_20373,N_20244);
xor U20583 (N_20583,N_20217,N_20309);
and U20584 (N_20584,N_20263,N_20205);
nand U20585 (N_20585,N_20249,N_20354);
nand U20586 (N_20586,N_20296,N_20287);
and U20587 (N_20587,N_20259,N_20205);
xnor U20588 (N_20588,N_20367,N_20331);
nand U20589 (N_20589,N_20310,N_20220);
and U20590 (N_20590,N_20272,N_20371);
xor U20591 (N_20591,N_20229,N_20241);
and U20592 (N_20592,N_20341,N_20205);
nand U20593 (N_20593,N_20339,N_20207);
nand U20594 (N_20594,N_20257,N_20394);
nand U20595 (N_20595,N_20286,N_20323);
and U20596 (N_20596,N_20359,N_20350);
xor U20597 (N_20597,N_20240,N_20386);
and U20598 (N_20598,N_20315,N_20259);
and U20599 (N_20599,N_20207,N_20242);
nand U20600 (N_20600,N_20494,N_20544);
nor U20601 (N_20601,N_20422,N_20512);
xor U20602 (N_20602,N_20489,N_20576);
nand U20603 (N_20603,N_20431,N_20595);
and U20604 (N_20604,N_20403,N_20402);
and U20605 (N_20605,N_20547,N_20421);
or U20606 (N_20606,N_20507,N_20492);
or U20607 (N_20607,N_20480,N_20574);
or U20608 (N_20608,N_20486,N_20482);
nor U20609 (N_20609,N_20521,N_20520);
xnor U20610 (N_20610,N_20585,N_20542);
nor U20611 (N_20611,N_20589,N_20514);
or U20612 (N_20612,N_20597,N_20581);
nor U20613 (N_20613,N_20473,N_20546);
xor U20614 (N_20614,N_20466,N_20543);
nor U20615 (N_20615,N_20592,N_20506);
nand U20616 (N_20616,N_20508,N_20411);
or U20617 (N_20617,N_20439,N_20485);
xnor U20618 (N_20618,N_20457,N_20529);
or U20619 (N_20619,N_20530,N_20562);
nand U20620 (N_20620,N_20469,N_20515);
xor U20621 (N_20621,N_20594,N_20598);
nand U20622 (N_20622,N_20596,N_20573);
and U20623 (N_20623,N_20458,N_20407);
nor U20624 (N_20624,N_20417,N_20541);
nor U20625 (N_20625,N_20495,N_20432);
nand U20626 (N_20626,N_20410,N_20519);
or U20627 (N_20627,N_20447,N_20516);
nor U20628 (N_20628,N_20496,N_20559);
and U20629 (N_20629,N_20577,N_20591);
or U20630 (N_20630,N_20548,N_20501);
nor U20631 (N_20631,N_20517,N_20582);
and U20632 (N_20632,N_20537,N_20586);
and U20633 (N_20633,N_20572,N_20427);
or U20634 (N_20634,N_20455,N_20483);
or U20635 (N_20635,N_20430,N_20563);
or U20636 (N_20636,N_20500,N_20535);
nand U20637 (N_20637,N_20477,N_20404);
nor U20638 (N_20638,N_20570,N_20524);
xor U20639 (N_20639,N_20545,N_20536);
and U20640 (N_20640,N_20493,N_20476);
xnor U20641 (N_20641,N_20557,N_20522);
or U20642 (N_20642,N_20461,N_20532);
nand U20643 (N_20643,N_20479,N_20564);
nor U20644 (N_20644,N_20587,N_20565);
xnor U20645 (N_20645,N_20440,N_20425);
nand U20646 (N_20646,N_20510,N_20567);
nor U20647 (N_20647,N_20504,N_20499);
nor U20648 (N_20648,N_20491,N_20505);
xnor U20649 (N_20649,N_20540,N_20405);
and U20650 (N_20650,N_20571,N_20468);
and U20651 (N_20651,N_20481,N_20451);
or U20652 (N_20652,N_20400,N_20470);
nor U20653 (N_20653,N_20560,N_20549);
nand U20654 (N_20654,N_20533,N_20472);
nand U20655 (N_20655,N_20462,N_20438);
nor U20656 (N_20656,N_20453,N_20450);
and U20657 (N_20657,N_20416,N_20478);
nor U20658 (N_20658,N_20456,N_20471);
xnor U20659 (N_20659,N_20434,N_20558);
nand U20660 (N_20660,N_20409,N_20490);
nor U20661 (N_20661,N_20525,N_20413);
nand U20662 (N_20662,N_20467,N_20474);
and U20663 (N_20663,N_20454,N_20502);
xnor U20664 (N_20664,N_20415,N_20555);
or U20665 (N_20665,N_20452,N_20408);
or U20666 (N_20666,N_20518,N_20578);
nand U20667 (N_20667,N_20513,N_20406);
nor U20668 (N_20668,N_20448,N_20412);
nand U20669 (N_20669,N_20449,N_20561);
nand U20670 (N_20670,N_20437,N_20556);
nand U20671 (N_20671,N_20534,N_20464);
nand U20672 (N_20672,N_20429,N_20484);
nor U20673 (N_20673,N_20488,N_20418);
nor U20674 (N_20674,N_20487,N_20580);
or U20675 (N_20675,N_20419,N_20593);
and U20676 (N_20676,N_20568,N_20414);
and U20677 (N_20677,N_20433,N_20551);
nand U20678 (N_20678,N_20511,N_20445);
or U20679 (N_20679,N_20401,N_20460);
and U20680 (N_20680,N_20441,N_20575);
nand U20681 (N_20681,N_20435,N_20554);
nand U20682 (N_20682,N_20509,N_20539);
nand U20683 (N_20683,N_20446,N_20526);
xnor U20684 (N_20684,N_20444,N_20590);
nand U20685 (N_20685,N_20503,N_20420);
and U20686 (N_20686,N_20423,N_20550);
nand U20687 (N_20687,N_20428,N_20465);
and U20688 (N_20688,N_20424,N_20436);
nor U20689 (N_20689,N_20531,N_20523);
nand U20690 (N_20690,N_20442,N_20553);
or U20691 (N_20691,N_20599,N_20569);
and U20692 (N_20692,N_20426,N_20527);
xnor U20693 (N_20693,N_20443,N_20538);
nand U20694 (N_20694,N_20588,N_20583);
or U20695 (N_20695,N_20566,N_20463);
or U20696 (N_20696,N_20579,N_20475);
xnor U20697 (N_20697,N_20497,N_20498);
nor U20698 (N_20698,N_20528,N_20584);
xnor U20699 (N_20699,N_20459,N_20552);
xor U20700 (N_20700,N_20433,N_20441);
and U20701 (N_20701,N_20401,N_20503);
xnor U20702 (N_20702,N_20506,N_20423);
or U20703 (N_20703,N_20435,N_20406);
xor U20704 (N_20704,N_20534,N_20515);
or U20705 (N_20705,N_20408,N_20519);
or U20706 (N_20706,N_20469,N_20445);
xor U20707 (N_20707,N_20541,N_20517);
nor U20708 (N_20708,N_20440,N_20555);
and U20709 (N_20709,N_20526,N_20452);
nor U20710 (N_20710,N_20443,N_20492);
or U20711 (N_20711,N_20570,N_20419);
and U20712 (N_20712,N_20576,N_20416);
nand U20713 (N_20713,N_20445,N_20401);
xnor U20714 (N_20714,N_20516,N_20509);
nand U20715 (N_20715,N_20446,N_20439);
nor U20716 (N_20716,N_20587,N_20437);
or U20717 (N_20717,N_20486,N_20565);
and U20718 (N_20718,N_20471,N_20494);
nand U20719 (N_20719,N_20464,N_20422);
nor U20720 (N_20720,N_20504,N_20481);
nor U20721 (N_20721,N_20570,N_20587);
nor U20722 (N_20722,N_20463,N_20464);
xnor U20723 (N_20723,N_20508,N_20585);
and U20724 (N_20724,N_20531,N_20428);
or U20725 (N_20725,N_20526,N_20531);
nand U20726 (N_20726,N_20521,N_20583);
nand U20727 (N_20727,N_20501,N_20473);
and U20728 (N_20728,N_20540,N_20567);
or U20729 (N_20729,N_20486,N_20557);
nand U20730 (N_20730,N_20587,N_20446);
or U20731 (N_20731,N_20544,N_20469);
or U20732 (N_20732,N_20482,N_20461);
xor U20733 (N_20733,N_20567,N_20582);
nand U20734 (N_20734,N_20487,N_20416);
xor U20735 (N_20735,N_20530,N_20501);
or U20736 (N_20736,N_20598,N_20567);
xnor U20737 (N_20737,N_20572,N_20492);
nand U20738 (N_20738,N_20408,N_20470);
nor U20739 (N_20739,N_20410,N_20413);
nand U20740 (N_20740,N_20536,N_20594);
or U20741 (N_20741,N_20540,N_20560);
nand U20742 (N_20742,N_20419,N_20468);
nand U20743 (N_20743,N_20417,N_20486);
and U20744 (N_20744,N_20567,N_20492);
xnor U20745 (N_20745,N_20512,N_20485);
or U20746 (N_20746,N_20434,N_20476);
nor U20747 (N_20747,N_20494,N_20441);
and U20748 (N_20748,N_20455,N_20440);
xnor U20749 (N_20749,N_20532,N_20550);
nand U20750 (N_20750,N_20573,N_20405);
nand U20751 (N_20751,N_20548,N_20405);
nor U20752 (N_20752,N_20477,N_20582);
and U20753 (N_20753,N_20462,N_20414);
or U20754 (N_20754,N_20582,N_20596);
nor U20755 (N_20755,N_20479,N_20582);
nand U20756 (N_20756,N_20579,N_20436);
nor U20757 (N_20757,N_20446,N_20469);
nor U20758 (N_20758,N_20459,N_20589);
and U20759 (N_20759,N_20478,N_20473);
nor U20760 (N_20760,N_20588,N_20519);
and U20761 (N_20761,N_20582,N_20572);
nor U20762 (N_20762,N_20490,N_20460);
nand U20763 (N_20763,N_20552,N_20423);
nor U20764 (N_20764,N_20570,N_20445);
nand U20765 (N_20765,N_20506,N_20500);
nor U20766 (N_20766,N_20589,N_20574);
nor U20767 (N_20767,N_20591,N_20426);
nor U20768 (N_20768,N_20575,N_20549);
nor U20769 (N_20769,N_20422,N_20504);
or U20770 (N_20770,N_20492,N_20403);
nand U20771 (N_20771,N_20548,N_20518);
nand U20772 (N_20772,N_20462,N_20456);
xnor U20773 (N_20773,N_20581,N_20409);
nor U20774 (N_20774,N_20407,N_20537);
nand U20775 (N_20775,N_20465,N_20527);
nor U20776 (N_20776,N_20565,N_20582);
nor U20777 (N_20777,N_20560,N_20529);
nand U20778 (N_20778,N_20434,N_20451);
nand U20779 (N_20779,N_20443,N_20540);
or U20780 (N_20780,N_20404,N_20432);
or U20781 (N_20781,N_20507,N_20475);
xor U20782 (N_20782,N_20480,N_20504);
or U20783 (N_20783,N_20497,N_20588);
or U20784 (N_20784,N_20547,N_20540);
and U20785 (N_20785,N_20415,N_20518);
nand U20786 (N_20786,N_20475,N_20421);
or U20787 (N_20787,N_20553,N_20573);
nor U20788 (N_20788,N_20401,N_20492);
and U20789 (N_20789,N_20523,N_20509);
xor U20790 (N_20790,N_20548,N_20577);
and U20791 (N_20791,N_20560,N_20495);
or U20792 (N_20792,N_20513,N_20568);
nand U20793 (N_20793,N_20586,N_20489);
or U20794 (N_20794,N_20588,N_20477);
xnor U20795 (N_20795,N_20455,N_20565);
xor U20796 (N_20796,N_20448,N_20498);
and U20797 (N_20797,N_20503,N_20484);
nor U20798 (N_20798,N_20423,N_20417);
or U20799 (N_20799,N_20414,N_20400);
nor U20800 (N_20800,N_20717,N_20727);
nor U20801 (N_20801,N_20651,N_20737);
nand U20802 (N_20802,N_20794,N_20626);
or U20803 (N_20803,N_20674,N_20754);
xor U20804 (N_20804,N_20732,N_20616);
and U20805 (N_20805,N_20612,N_20729);
xor U20806 (N_20806,N_20765,N_20780);
and U20807 (N_20807,N_20630,N_20688);
and U20808 (N_20808,N_20639,N_20681);
and U20809 (N_20809,N_20691,N_20698);
nand U20810 (N_20810,N_20778,N_20654);
and U20811 (N_20811,N_20624,N_20632);
or U20812 (N_20812,N_20665,N_20606);
or U20813 (N_20813,N_20693,N_20713);
and U20814 (N_20814,N_20670,N_20694);
nand U20815 (N_20815,N_20603,N_20657);
and U20816 (N_20816,N_20753,N_20623);
nor U20817 (N_20817,N_20745,N_20772);
xor U20818 (N_20818,N_20705,N_20748);
xor U20819 (N_20819,N_20667,N_20782);
or U20820 (N_20820,N_20704,N_20611);
xnor U20821 (N_20821,N_20669,N_20786);
or U20822 (N_20822,N_20712,N_20771);
nand U20823 (N_20823,N_20796,N_20615);
xor U20824 (N_20824,N_20672,N_20768);
or U20825 (N_20825,N_20760,N_20677);
xor U20826 (N_20826,N_20610,N_20730);
and U20827 (N_20827,N_20661,N_20638);
nor U20828 (N_20828,N_20758,N_20660);
xnor U20829 (N_20829,N_20620,N_20631);
xor U20830 (N_20830,N_20707,N_20618);
nor U20831 (N_20831,N_20696,N_20723);
nor U20832 (N_20832,N_20656,N_20766);
nor U20833 (N_20833,N_20637,N_20684);
nand U20834 (N_20834,N_20728,N_20678);
or U20835 (N_20835,N_20746,N_20605);
xnor U20836 (N_20836,N_20608,N_20602);
nand U20837 (N_20837,N_20719,N_20708);
or U20838 (N_20838,N_20726,N_20617);
nor U20839 (N_20839,N_20613,N_20761);
or U20840 (N_20840,N_20734,N_20756);
or U20841 (N_20841,N_20647,N_20784);
nor U20842 (N_20842,N_20648,N_20663);
nand U20843 (N_20843,N_20673,N_20783);
or U20844 (N_20844,N_20628,N_20750);
or U20845 (N_20845,N_20742,N_20664);
xnor U20846 (N_20846,N_20722,N_20706);
xnor U20847 (N_20847,N_20655,N_20682);
and U20848 (N_20848,N_20791,N_20721);
nand U20849 (N_20849,N_20697,N_20738);
nand U20850 (N_20850,N_20741,N_20650);
xor U20851 (N_20851,N_20767,N_20755);
or U20852 (N_20852,N_20649,N_20646);
nand U20853 (N_20853,N_20675,N_20720);
and U20854 (N_20854,N_20621,N_20716);
or U20855 (N_20855,N_20652,N_20793);
nand U20856 (N_20856,N_20788,N_20799);
nand U20857 (N_20857,N_20789,N_20659);
nand U20858 (N_20858,N_20744,N_20636);
and U20859 (N_20859,N_20773,N_20690);
xor U20860 (N_20860,N_20770,N_20736);
xnor U20861 (N_20861,N_20640,N_20635);
and U20862 (N_20862,N_20774,N_20790);
or U20863 (N_20863,N_20699,N_20743);
xor U20864 (N_20864,N_20625,N_20781);
nand U20865 (N_20865,N_20622,N_20683);
xor U20866 (N_20866,N_20762,N_20700);
nor U20867 (N_20867,N_20757,N_20763);
and U20868 (N_20868,N_20644,N_20797);
nand U20869 (N_20869,N_20614,N_20785);
and U20870 (N_20870,N_20792,N_20666);
or U20871 (N_20871,N_20619,N_20662);
nor U20872 (N_20872,N_20658,N_20779);
nor U20873 (N_20873,N_20714,N_20679);
nand U20874 (N_20874,N_20687,N_20642);
and U20875 (N_20875,N_20747,N_20749);
nand U20876 (N_20876,N_20725,N_20703);
and U20877 (N_20877,N_20604,N_20701);
or U20878 (N_20878,N_20692,N_20752);
nand U20879 (N_20879,N_20634,N_20739);
or U20880 (N_20880,N_20653,N_20641);
nand U20881 (N_20881,N_20718,N_20607);
xnor U20882 (N_20882,N_20685,N_20764);
or U20883 (N_20883,N_20724,N_20686);
nand U20884 (N_20884,N_20643,N_20740);
xnor U20885 (N_20885,N_20798,N_20769);
and U20886 (N_20886,N_20731,N_20633);
nand U20887 (N_20887,N_20759,N_20709);
xnor U20888 (N_20888,N_20689,N_20735);
or U20889 (N_20889,N_20777,N_20600);
or U20890 (N_20890,N_20751,N_20795);
xor U20891 (N_20891,N_20629,N_20695);
or U20892 (N_20892,N_20668,N_20676);
nand U20893 (N_20893,N_20601,N_20627);
and U20894 (N_20894,N_20733,N_20776);
and U20895 (N_20895,N_20715,N_20775);
nor U20896 (N_20896,N_20702,N_20787);
nor U20897 (N_20897,N_20710,N_20711);
xor U20898 (N_20898,N_20680,N_20609);
nand U20899 (N_20899,N_20645,N_20671);
xor U20900 (N_20900,N_20639,N_20712);
and U20901 (N_20901,N_20691,N_20766);
xnor U20902 (N_20902,N_20730,N_20665);
nor U20903 (N_20903,N_20654,N_20797);
nor U20904 (N_20904,N_20693,N_20701);
nand U20905 (N_20905,N_20690,N_20697);
and U20906 (N_20906,N_20623,N_20769);
or U20907 (N_20907,N_20773,N_20696);
and U20908 (N_20908,N_20782,N_20763);
and U20909 (N_20909,N_20708,N_20650);
xnor U20910 (N_20910,N_20754,N_20647);
xor U20911 (N_20911,N_20795,N_20689);
xor U20912 (N_20912,N_20668,N_20763);
and U20913 (N_20913,N_20671,N_20647);
and U20914 (N_20914,N_20639,N_20671);
or U20915 (N_20915,N_20667,N_20727);
xor U20916 (N_20916,N_20798,N_20782);
and U20917 (N_20917,N_20652,N_20644);
xnor U20918 (N_20918,N_20692,N_20633);
or U20919 (N_20919,N_20663,N_20662);
xor U20920 (N_20920,N_20794,N_20744);
and U20921 (N_20921,N_20646,N_20789);
nor U20922 (N_20922,N_20780,N_20648);
or U20923 (N_20923,N_20751,N_20603);
or U20924 (N_20924,N_20785,N_20781);
xnor U20925 (N_20925,N_20643,N_20728);
nor U20926 (N_20926,N_20645,N_20639);
xor U20927 (N_20927,N_20640,N_20782);
and U20928 (N_20928,N_20640,N_20626);
xor U20929 (N_20929,N_20765,N_20664);
and U20930 (N_20930,N_20633,N_20652);
nor U20931 (N_20931,N_20739,N_20631);
or U20932 (N_20932,N_20712,N_20740);
nand U20933 (N_20933,N_20765,N_20752);
or U20934 (N_20934,N_20629,N_20703);
nand U20935 (N_20935,N_20727,N_20787);
or U20936 (N_20936,N_20774,N_20755);
nand U20937 (N_20937,N_20616,N_20776);
xnor U20938 (N_20938,N_20725,N_20668);
nor U20939 (N_20939,N_20673,N_20600);
nand U20940 (N_20940,N_20734,N_20608);
nand U20941 (N_20941,N_20776,N_20767);
nand U20942 (N_20942,N_20675,N_20603);
and U20943 (N_20943,N_20631,N_20738);
and U20944 (N_20944,N_20774,N_20775);
nor U20945 (N_20945,N_20613,N_20757);
nor U20946 (N_20946,N_20660,N_20782);
and U20947 (N_20947,N_20667,N_20680);
or U20948 (N_20948,N_20734,N_20708);
nor U20949 (N_20949,N_20795,N_20755);
xor U20950 (N_20950,N_20745,N_20761);
and U20951 (N_20951,N_20754,N_20780);
nor U20952 (N_20952,N_20796,N_20720);
nand U20953 (N_20953,N_20634,N_20655);
or U20954 (N_20954,N_20641,N_20722);
nand U20955 (N_20955,N_20739,N_20754);
and U20956 (N_20956,N_20666,N_20754);
xnor U20957 (N_20957,N_20652,N_20744);
nor U20958 (N_20958,N_20688,N_20770);
nand U20959 (N_20959,N_20662,N_20697);
nor U20960 (N_20960,N_20693,N_20639);
nand U20961 (N_20961,N_20745,N_20795);
and U20962 (N_20962,N_20682,N_20722);
nor U20963 (N_20963,N_20626,N_20718);
xor U20964 (N_20964,N_20623,N_20732);
nand U20965 (N_20965,N_20660,N_20632);
and U20966 (N_20966,N_20614,N_20685);
or U20967 (N_20967,N_20792,N_20778);
and U20968 (N_20968,N_20688,N_20746);
and U20969 (N_20969,N_20771,N_20674);
or U20970 (N_20970,N_20721,N_20644);
or U20971 (N_20971,N_20776,N_20720);
or U20972 (N_20972,N_20635,N_20753);
xnor U20973 (N_20973,N_20798,N_20688);
nor U20974 (N_20974,N_20776,N_20653);
and U20975 (N_20975,N_20707,N_20623);
nor U20976 (N_20976,N_20704,N_20687);
nand U20977 (N_20977,N_20702,N_20606);
xor U20978 (N_20978,N_20605,N_20651);
xor U20979 (N_20979,N_20737,N_20725);
xor U20980 (N_20980,N_20744,N_20625);
xnor U20981 (N_20981,N_20650,N_20756);
and U20982 (N_20982,N_20674,N_20648);
xor U20983 (N_20983,N_20797,N_20737);
and U20984 (N_20984,N_20768,N_20653);
nor U20985 (N_20985,N_20730,N_20759);
xor U20986 (N_20986,N_20767,N_20789);
and U20987 (N_20987,N_20665,N_20644);
xnor U20988 (N_20988,N_20649,N_20604);
nor U20989 (N_20989,N_20721,N_20797);
nor U20990 (N_20990,N_20657,N_20616);
nand U20991 (N_20991,N_20765,N_20631);
xor U20992 (N_20992,N_20666,N_20678);
nor U20993 (N_20993,N_20645,N_20782);
or U20994 (N_20994,N_20763,N_20729);
nor U20995 (N_20995,N_20692,N_20718);
and U20996 (N_20996,N_20737,N_20768);
nor U20997 (N_20997,N_20760,N_20724);
xor U20998 (N_20998,N_20656,N_20689);
nand U20999 (N_20999,N_20778,N_20776);
and U21000 (N_21000,N_20852,N_20840);
xor U21001 (N_21001,N_20981,N_20999);
and U21002 (N_21002,N_20837,N_20950);
and U21003 (N_21003,N_20888,N_20801);
or U21004 (N_21004,N_20823,N_20929);
nor U21005 (N_21005,N_20937,N_20897);
nor U21006 (N_21006,N_20844,N_20831);
nor U21007 (N_21007,N_20945,N_20963);
or U21008 (N_21008,N_20836,N_20901);
nor U21009 (N_21009,N_20900,N_20804);
and U21010 (N_21010,N_20848,N_20931);
nor U21011 (N_21011,N_20946,N_20940);
xor U21012 (N_21012,N_20994,N_20984);
xnor U21013 (N_21013,N_20976,N_20975);
nand U21014 (N_21014,N_20849,N_20908);
or U21015 (N_21015,N_20991,N_20838);
or U21016 (N_21016,N_20827,N_20828);
nor U21017 (N_21017,N_20830,N_20839);
and U21018 (N_21018,N_20814,N_20986);
xnor U21019 (N_21019,N_20859,N_20921);
or U21020 (N_21020,N_20861,N_20802);
and U21021 (N_21021,N_20974,N_20807);
xnor U21022 (N_21022,N_20817,N_20925);
and U21023 (N_21023,N_20887,N_20961);
xor U21024 (N_21024,N_20924,N_20906);
and U21025 (N_21025,N_20987,N_20850);
and U21026 (N_21026,N_20959,N_20870);
or U21027 (N_21027,N_20862,N_20882);
nand U21028 (N_21028,N_20926,N_20892);
or U21029 (N_21029,N_20853,N_20810);
nor U21030 (N_21030,N_20867,N_20915);
or U21031 (N_21031,N_20927,N_20938);
xnor U21032 (N_21032,N_20889,N_20972);
xor U21033 (N_21033,N_20910,N_20868);
xor U21034 (N_21034,N_20983,N_20812);
and U21035 (N_21035,N_20876,N_20829);
nand U21036 (N_21036,N_20855,N_20835);
nor U21037 (N_21037,N_20824,N_20885);
xor U21038 (N_21038,N_20898,N_20942);
xnor U21039 (N_21039,N_20922,N_20866);
xnor U21040 (N_21040,N_20894,N_20904);
xor U21041 (N_21041,N_20988,N_20952);
xor U21042 (N_21042,N_20919,N_20934);
nand U21043 (N_21043,N_20913,N_20822);
nor U21044 (N_21044,N_20857,N_20944);
or U21045 (N_21045,N_20834,N_20912);
nor U21046 (N_21046,N_20815,N_20821);
nor U21047 (N_21047,N_20808,N_20918);
nand U21048 (N_21048,N_20960,N_20930);
nor U21049 (N_21049,N_20956,N_20971);
nor U21050 (N_21050,N_20943,N_20879);
xnor U21051 (N_21051,N_20955,N_20949);
and U21052 (N_21052,N_20869,N_20905);
xnor U21053 (N_21053,N_20966,N_20883);
or U21054 (N_21054,N_20874,N_20809);
or U21055 (N_21055,N_20967,N_20843);
nor U21056 (N_21056,N_20872,N_20928);
and U21057 (N_21057,N_20978,N_20841);
nand U21058 (N_21058,N_20902,N_20800);
nor U21059 (N_21059,N_20951,N_20997);
nor U21060 (N_21060,N_20858,N_20965);
nand U21061 (N_21061,N_20935,N_20939);
nand U21062 (N_21062,N_20881,N_20958);
xor U21063 (N_21063,N_20811,N_20825);
or U21064 (N_21064,N_20989,N_20911);
xnor U21065 (N_21065,N_20886,N_20819);
xnor U21066 (N_21066,N_20923,N_20964);
nand U21067 (N_21067,N_20968,N_20877);
xor U21068 (N_21068,N_20969,N_20973);
nand U21069 (N_21069,N_20863,N_20820);
nor U21070 (N_21070,N_20995,N_20860);
or U21071 (N_21071,N_20899,N_20982);
nand U21072 (N_21072,N_20846,N_20980);
and U21073 (N_21073,N_20832,N_20909);
or U21074 (N_21074,N_20979,N_20948);
xor U21075 (N_21075,N_20992,N_20920);
xor U21076 (N_21076,N_20970,N_20917);
xnor U21077 (N_21077,N_20953,N_20896);
nor U21078 (N_21078,N_20936,N_20842);
nor U21079 (N_21079,N_20916,N_20954);
and U21080 (N_21080,N_20977,N_20998);
xor U21081 (N_21081,N_20884,N_20833);
nor U21082 (N_21082,N_20845,N_20893);
nor U21083 (N_21083,N_20985,N_20865);
and U21084 (N_21084,N_20854,N_20907);
or U21085 (N_21085,N_20895,N_20826);
nand U21086 (N_21086,N_20880,N_20890);
or U21087 (N_21087,N_20864,N_20947);
or U21088 (N_21088,N_20993,N_20818);
and U21089 (N_21089,N_20856,N_20941);
xnor U21090 (N_21090,N_20806,N_20851);
or U21091 (N_21091,N_20875,N_20878);
or U21092 (N_21092,N_20805,N_20990);
and U21093 (N_21093,N_20914,N_20871);
nand U21094 (N_21094,N_20813,N_20933);
or U21095 (N_21095,N_20957,N_20873);
nor U21096 (N_21096,N_20847,N_20816);
and U21097 (N_21097,N_20996,N_20932);
or U21098 (N_21098,N_20803,N_20891);
nand U21099 (N_21099,N_20903,N_20962);
or U21100 (N_21100,N_20803,N_20839);
nand U21101 (N_21101,N_20892,N_20836);
xor U21102 (N_21102,N_20979,N_20915);
nand U21103 (N_21103,N_20919,N_20840);
or U21104 (N_21104,N_20855,N_20949);
xnor U21105 (N_21105,N_20925,N_20916);
nand U21106 (N_21106,N_20947,N_20901);
nand U21107 (N_21107,N_20985,N_20888);
nand U21108 (N_21108,N_20860,N_20879);
and U21109 (N_21109,N_20920,N_20844);
or U21110 (N_21110,N_20908,N_20866);
xnor U21111 (N_21111,N_20877,N_20983);
nand U21112 (N_21112,N_20951,N_20868);
nand U21113 (N_21113,N_20946,N_20820);
nor U21114 (N_21114,N_20804,N_20974);
nor U21115 (N_21115,N_20970,N_20916);
xor U21116 (N_21116,N_20951,N_20958);
nor U21117 (N_21117,N_20862,N_20867);
xnor U21118 (N_21118,N_20993,N_20938);
or U21119 (N_21119,N_20945,N_20990);
or U21120 (N_21120,N_20942,N_20937);
nand U21121 (N_21121,N_20815,N_20800);
nand U21122 (N_21122,N_20859,N_20963);
nand U21123 (N_21123,N_20927,N_20891);
nand U21124 (N_21124,N_20961,N_20877);
xnor U21125 (N_21125,N_20927,N_20951);
or U21126 (N_21126,N_20831,N_20910);
and U21127 (N_21127,N_20901,N_20940);
xor U21128 (N_21128,N_20852,N_20945);
xor U21129 (N_21129,N_20903,N_20847);
and U21130 (N_21130,N_20975,N_20838);
or U21131 (N_21131,N_20878,N_20965);
or U21132 (N_21132,N_20974,N_20970);
xor U21133 (N_21133,N_20949,N_20998);
nor U21134 (N_21134,N_20890,N_20851);
or U21135 (N_21135,N_20827,N_20810);
xor U21136 (N_21136,N_20810,N_20905);
xnor U21137 (N_21137,N_20848,N_20811);
and U21138 (N_21138,N_20987,N_20869);
nor U21139 (N_21139,N_20871,N_20873);
nand U21140 (N_21140,N_20992,N_20995);
or U21141 (N_21141,N_20808,N_20860);
nor U21142 (N_21142,N_20872,N_20977);
xnor U21143 (N_21143,N_20855,N_20817);
xor U21144 (N_21144,N_20863,N_20926);
or U21145 (N_21145,N_20982,N_20988);
xnor U21146 (N_21146,N_20908,N_20865);
nor U21147 (N_21147,N_20877,N_20959);
and U21148 (N_21148,N_20984,N_20852);
nand U21149 (N_21149,N_20964,N_20853);
or U21150 (N_21150,N_20877,N_20990);
and U21151 (N_21151,N_20820,N_20961);
or U21152 (N_21152,N_20847,N_20936);
and U21153 (N_21153,N_20961,N_20900);
nor U21154 (N_21154,N_20836,N_20810);
nand U21155 (N_21155,N_20978,N_20866);
nor U21156 (N_21156,N_20970,N_20939);
xor U21157 (N_21157,N_20885,N_20869);
nor U21158 (N_21158,N_20946,N_20913);
nand U21159 (N_21159,N_20851,N_20887);
or U21160 (N_21160,N_20925,N_20991);
xor U21161 (N_21161,N_20926,N_20972);
xnor U21162 (N_21162,N_20943,N_20989);
xnor U21163 (N_21163,N_20800,N_20976);
xnor U21164 (N_21164,N_20862,N_20884);
or U21165 (N_21165,N_20822,N_20953);
xor U21166 (N_21166,N_20817,N_20825);
xor U21167 (N_21167,N_20886,N_20805);
nor U21168 (N_21168,N_20825,N_20840);
nand U21169 (N_21169,N_20906,N_20812);
xor U21170 (N_21170,N_20959,N_20840);
nand U21171 (N_21171,N_20971,N_20843);
or U21172 (N_21172,N_20877,N_20962);
and U21173 (N_21173,N_20900,N_20923);
xor U21174 (N_21174,N_20965,N_20807);
and U21175 (N_21175,N_20870,N_20967);
nand U21176 (N_21176,N_20880,N_20947);
nor U21177 (N_21177,N_20951,N_20812);
nor U21178 (N_21178,N_20922,N_20893);
or U21179 (N_21179,N_20924,N_20895);
nor U21180 (N_21180,N_20819,N_20869);
xnor U21181 (N_21181,N_20849,N_20957);
and U21182 (N_21182,N_20995,N_20953);
and U21183 (N_21183,N_20802,N_20925);
nor U21184 (N_21184,N_20851,N_20965);
xnor U21185 (N_21185,N_20971,N_20961);
or U21186 (N_21186,N_20931,N_20951);
nor U21187 (N_21187,N_20921,N_20820);
and U21188 (N_21188,N_20964,N_20954);
nor U21189 (N_21189,N_20916,N_20906);
xnor U21190 (N_21190,N_20968,N_20996);
or U21191 (N_21191,N_20875,N_20856);
and U21192 (N_21192,N_20905,N_20899);
xnor U21193 (N_21193,N_20828,N_20936);
or U21194 (N_21194,N_20879,N_20948);
xor U21195 (N_21195,N_20857,N_20917);
and U21196 (N_21196,N_20811,N_20957);
or U21197 (N_21197,N_20828,N_20846);
xnor U21198 (N_21198,N_20825,N_20959);
and U21199 (N_21199,N_20970,N_20954);
and U21200 (N_21200,N_21004,N_21022);
nand U21201 (N_21201,N_21170,N_21007);
xor U21202 (N_21202,N_21072,N_21058);
and U21203 (N_21203,N_21136,N_21037);
and U21204 (N_21204,N_21156,N_21149);
or U21205 (N_21205,N_21084,N_21100);
xnor U21206 (N_21206,N_21083,N_21002);
nor U21207 (N_21207,N_21173,N_21109);
nor U21208 (N_21208,N_21044,N_21011);
nand U21209 (N_21209,N_21154,N_21014);
nand U21210 (N_21210,N_21023,N_21094);
nand U21211 (N_21211,N_21157,N_21150);
or U21212 (N_21212,N_21138,N_21021);
and U21213 (N_21213,N_21195,N_21045);
nand U21214 (N_21214,N_21118,N_21019);
or U21215 (N_21215,N_21175,N_21171);
xnor U21216 (N_21216,N_21038,N_21028);
xnor U21217 (N_21217,N_21061,N_21114);
or U21218 (N_21218,N_21165,N_21142);
nor U21219 (N_21219,N_21132,N_21107);
and U21220 (N_21220,N_21128,N_21112);
xor U21221 (N_21221,N_21148,N_21020);
or U21222 (N_21222,N_21184,N_21013);
and U21223 (N_21223,N_21090,N_21104);
xnor U21224 (N_21224,N_21127,N_21026);
xor U21225 (N_21225,N_21032,N_21027);
nand U21226 (N_21226,N_21144,N_21135);
nand U21227 (N_21227,N_21160,N_21041);
xor U21228 (N_21228,N_21187,N_21024);
or U21229 (N_21229,N_21102,N_21034);
nor U21230 (N_21230,N_21054,N_21015);
nor U21231 (N_21231,N_21153,N_21003);
or U21232 (N_21232,N_21191,N_21111);
and U21233 (N_21233,N_21120,N_21182);
nor U21234 (N_21234,N_21080,N_21008);
or U21235 (N_21235,N_21172,N_21155);
nand U21236 (N_21236,N_21091,N_21099);
nand U21237 (N_21237,N_21039,N_21159);
nor U21238 (N_21238,N_21001,N_21093);
or U21239 (N_21239,N_21052,N_21035);
xor U21240 (N_21240,N_21095,N_21079);
or U21241 (N_21241,N_21197,N_21167);
nand U21242 (N_21242,N_21030,N_21193);
nor U21243 (N_21243,N_21125,N_21049);
xnor U21244 (N_21244,N_21115,N_21189);
or U21245 (N_21245,N_21117,N_21124);
and U21246 (N_21246,N_21075,N_21178);
or U21247 (N_21247,N_21000,N_21055);
nor U21248 (N_21248,N_21169,N_21101);
xnor U21249 (N_21249,N_21057,N_21063);
nand U21250 (N_21250,N_21005,N_21121);
nand U21251 (N_21251,N_21183,N_21050);
nor U21252 (N_21252,N_21053,N_21110);
nand U21253 (N_21253,N_21129,N_21033);
or U21254 (N_21254,N_21017,N_21056);
nor U21255 (N_21255,N_21010,N_21087);
or U21256 (N_21256,N_21076,N_21194);
nand U21257 (N_21257,N_21163,N_21036);
nor U21258 (N_21258,N_21152,N_21066);
and U21259 (N_21259,N_21126,N_21164);
xor U21260 (N_21260,N_21180,N_21070);
nor U21261 (N_21261,N_21025,N_21143);
or U21262 (N_21262,N_21016,N_21151);
and U21263 (N_21263,N_21166,N_21198);
or U21264 (N_21264,N_21074,N_21012);
nand U21265 (N_21265,N_21051,N_21060);
and U21266 (N_21266,N_21068,N_21062);
xor U21267 (N_21267,N_21131,N_21098);
or U21268 (N_21268,N_21179,N_21134);
xor U21269 (N_21269,N_21031,N_21123);
nand U21270 (N_21270,N_21168,N_21082);
nand U21271 (N_21271,N_21119,N_21130);
and U21272 (N_21272,N_21089,N_21185);
xnor U21273 (N_21273,N_21181,N_21047);
nand U21274 (N_21274,N_21065,N_21078);
nor U21275 (N_21275,N_21137,N_21199);
xnor U21276 (N_21276,N_21177,N_21158);
or U21277 (N_21277,N_21188,N_21140);
nor U21278 (N_21278,N_21106,N_21162);
nand U21279 (N_21279,N_21029,N_21145);
and U21280 (N_21280,N_21071,N_21146);
and U21281 (N_21281,N_21018,N_21122);
or U21282 (N_21282,N_21174,N_21141);
and U21283 (N_21283,N_21176,N_21086);
nand U21284 (N_21284,N_21009,N_21059);
and U21285 (N_21285,N_21046,N_21092);
nor U21286 (N_21286,N_21069,N_21108);
and U21287 (N_21287,N_21043,N_21192);
nor U21288 (N_21288,N_21042,N_21088);
nor U21289 (N_21289,N_21105,N_21186);
or U21290 (N_21290,N_21097,N_21133);
nor U21291 (N_21291,N_21139,N_21113);
xor U21292 (N_21292,N_21077,N_21116);
and U21293 (N_21293,N_21161,N_21064);
nor U21294 (N_21294,N_21196,N_21040);
and U21295 (N_21295,N_21190,N_21048);
and U21296 (N_21296,N_21096,N_21103);
xor U21297 (N_21297,N_21081,N_21073);
nor U21298 (N_21298,N_21006,N_21067);
nor U21299 (N_21299,N_21085,N_21147);
and U21300 (N_21300,N_21028,N_21067);
nand U21301 (N_21301,N_21175,N_21020);
and U21302 (N_21302,N_21051,N_21167);
xnor U21303 (N_21303,N_21077,N_21167);
or U21304 (N_21304,N_21026,N_21071);
and U21305 (N_21305,N_21033,N_21174);
and U21306 (N_21306,N_21146,N_21102);
nor U21307 (N_21307,N_21031,N_21167);
xnor U21308 (N_21308,N_21137,N_21177);
nand U21309 (N_21309,N_21110,N_21090);
nand U21310 (N_21310,N_21081,N_21070);
nor U21311 (N_21311,N_21061,N_21081);
or U21312 (N_21312,N_21153,N_21140);
xnor U21313 (N_21313,N_21033,N_21085);
nor U21314 (N_21314,N_21183,N_21103);
and U21315 (N_21315,N_21165,N_21155);
or U21316 (N_21316,N_21108,N_21039);
nand U21317 (N_21317,N_21125,N_21045);
nand U21318 (N_21318,N_21079,N_21076);
xor U21319 (N_21319,N_21029,N_21082);
or U21320 (N_21320,N_21093,N_21018);
or U21321 (N_21321,N_21092,N_21182);
nor U21322 (N_21322,N_21020,N_21100);
and U21323 (N_21323,N_21006,N_21032);
and U21324 (N_21324,N_21138,N_21023);
nand U21325 (N_21325,N_21075,N_21103);
and U21326 (N_21326,N_21167,N_21199);
or U21327 (N_21327,N_21002,N_21183);
xnor U21328 (N_21328,N_21171,N_21008);
nor U21329 (N_21329,N_21084,N_21184);
nor U21330 (N_21330,N_21125,N_21003);
nor U21331 (N_21331,N_21034,N_21070);
and U21332 (N_21332,N_21170,N_21117);
nand U21333 (N_21333,N_21068,N_21126);
xor U21334 (N_21334,N_21044,N_21025);
nand U21335 (N_21335,N_21009,N_21191);
nand U21336 (N_21336,N_21019,N_21002);
and U21337 (N_21337,N_21041,N_21170);
nand U21338 (N_21338,N_21039,N_21014);
nand U21339 (N_21339,N_21191,N_21103);
nand U21340 (N_21340,N_21083,N_21162);
xnor U21341 (N_21341,N_21016,N_21199);
nor U21342 (N_21342,N_21168,N_21036);
xnor U21343 (N_21343,N_21138,N_21030);
xor U21344 (N_21344,N_21061,N_21084);
xor U21345 (N_21345,N_21193,N_21116);
and U21346 (N_21346,N_21139,N_21065);
or U21347 (N_21347,N_21067,N_21114);
or U21348 (N_21348,N_21131,N_21049);
nor U21349 (N_21349,N_21110,N_21169);
xor U21350 (N_21350,N_21088,N_21087);
and U21351 (N_21351,N_21087,N_21044);
nor U21352 (N_21352,N_21005,N_21013);
nor U21353 (N_21353,N_21042,N_21177);
and U21354 (N_21354,N_21070,N_21162);
and U21355 (N_21355,N_21115,N_21017);
or U21356 (N_21356,N_21032,N_21149);
or U21357 (N_21357,N_21149,N_21192);
and U21358 (N_21358,N_21042,N_21072);
nor U21359 (N_21359,N_21084,N_21122);
or U21360 (N_21360,N_21174,N_21112);
nand U21361 (N_21361,N_21054,N_21065);
and U21362 (N_21362,N_21065,N_21109);
and U21363 (N_21363,N_21052,N_21017);
nand U21364 (N_21364,N_21042,N_21089);
xor U21365 (N_21365,N_21090,N_21199);
nand U21366 (N_21366,N_21023,N_21022);
and U21367 (N_21367,N_21048,N_21032);
nor U21368 (N_21368,N_21145,N_21024);
nor U21369 (N_21369,N_21176,N_21050);
xnor U21370 (N_21370,N_21102,N_21127);
nor U21371 (N_21371,N_21148,N_21185);
nor U21372 (N_21372,N_21105,N_21133);
nor U21373 (N_21373,N_21149,N_21166);
xnor U21374 (N_21374,N_21172,N_21104);
or U21375 (N_21375,N_21130,N_21088);
nand U21376 (N_21376,N_21125,N_21185);
nand U21377 (N_21377,N_21110,N_21179);
nor U21378 (N_21378,N_21095,N_21014);
nand U21379 (N_21379,N_21180,N_21014);
and U21380 (N_21380,N_21168,N_21130);
or U21381 (N_21381,N_21006,N_21082);
or U21382 (N_21382,N_21012,N_21009);
and U21383 (N_21383,N_21178,N_21189);
nor U21384 (N_21384,N_21192,N_21122);
and U21385 (N_21385,N_21108,N_21195);
nor U21386 (N_21386,N_21063,N_21191);
or U21387 (N_21387,N_21011,N_21173);
and U21388 (N_21388,N_21039,N_21017);
nor U21389 (N_21389,N_21048,N_21057);
or U21390 (N_21390,N_21044,N_21148);
nand U21391 (N_21391,N_21071,N_21142);
nor U21392 (N_21392,N_21003,N_21031);
nor U21393 (N_21393,N_21190,N_21020);
nand U21394 (N_21394,N_21024,N_21031);
and U21395 (N_21395,N_21043,N_21190);
or U21396 (N_21396,N_21139,N_21010);
nor U21397 (N_21397,N_21003,N_21099);
or U21398 (N_21398,N_21175,N_21069);
and U21399 (N_21399,N_21064,N_21106);
nor U21400 (N_21400,N_21296,N_21242);
or U21401 (N_21401,N_21340,N_21358);
xnor U21402 (N_21402,N_21353,N_21321);
nor U21403 (N_21403,N_21378,N_21273);
nand U21404 (N_21404,N_21349,N_21337);
nor U21405 (N_21405,N_21259,N_21260);
and U21406 (N_21406,N_21372,N_21308);
nand U21407 (N_21407,N_21280,N_21215);
or U21408 (N_21408,N_21394,N_21342);
nand U21409 (N_21409,N_21395,N_21346);
nand U21410 (N_21410,N_21294,N_21206);
or U21411 (N_21411,N_21329,N_21210);
or U21412 (N_21412,N_21276,N_21275);
nand U21413 (N_21413,N_21355,N_21331);
nand U21414 (N_21414,N_21257,N_21357);
xnor U21415 (N_21415,N_21200,N_21309);
nand U21416 (N_21416,N_21343,N_21222);
or U21417 (N_21417,N_21283,N_21364);
nand U21418 (N_21418,N_21333,N_21396);
nand U21419 (N_21419,N_21310,N_21356);
and U21420 (N_21420,N_21214,N_21319);
xnor U21421 (N_21421,N_21362,N_21313);
or U21422 (N_21422,N_21256,N_21204);
or U21423 (N_21423,N_21387,N_21376);
xor U21424 (N_21424,N_21380,N_21374);
xor U21425 (N_21425,N_21315,N_21347);
nor U21426 (N_21426,N_21390,N_21295);
nor U21427 (N_21427,N_21251,N_21237);
or U21428 (N_21428,N_21258,N_21377);
nor U21429 (N_21429,N_21304,N_21207);
or U21430 (N_21430,N_21216,N_21320);
nor U21431 (N_21431,N_21359,N_21263);
or U21432 (N_21432,N_21290,N_21203);
xnor U21433 (N_21433,N_21219,N_21384);
nand U21434 (N_21434,N_21370,N_21247);
nand U21435 (N_21435,N_21250,N_21234);
nor U21436 (N_21436,N_21239,N_21299);
xor U21437 (N_21437,N_21391,N_21350);
nand U21438 (N_21438,N_21375,N_21270);
or U21439 (N_21439,N_21326,N_21245);
nor U21440 (N_21440,N_21332,N_21302);
and U21441 (N_21441,N_21262,N_21318);
or U21442 (N_21442,N_21352,N_21316);
nor U21443 (N_21443,N_21366,N_21334);
nor U21444 (N_21444,N_21365,N_21348);
or U21445 (N_21445,N_21341,N_21360);
and U21446 (N_21446,N_21286,N_21227);
nor U21447 (N_21447,N_21211,N_21393);
nand U21448 (N_21448,N_21323,N_21240);
xor U21449 (N_21449,N_21314,N_21264);
and U21450 (N_21450,N_21266,N_21298);
or U21451 (N_21451,N_21361,N_21363);
nor U21452 (N_21452,N_21297,N_21307);
xnor U21453 (N_21453,N_21399,N_21312);
and U21454 (N_21454,N_21383,N_21287);
xnor U21455 (N_21455,N_21382,N_21261);
nor U21456 (N_21456,N_21324,N_21351);
or U21457 (N_21457,N_21209,N_21202);
xor U21458 (N_21458,N_21249,N_21267);
or U21459 (N_21459,N_21278,N_21208);
or U21460 (N_21460,N_21281,N_21201);
nand U21461 (N_21461,N_21241,N_21229);
nor U21462 (N_21462,N_21389,N_21205);
and U21463 (N_21463,N_21371,N_21230);
xnor U21464 (N_21464,N_21272,N_21379);
or U21465 (N_21465,N_21292,N_21367);
nor U21466 (N_21466,N_21328,N_21255);
and U21467 (N_21467,N_21388,N_21235);
nor U21468 (N_21468,N_21311,N_21269);
and U21469 (N_21469,N_21265,N_21327);
xor U21470 (N_21470,N_21226,N_21212);
xnor U21471 (N_21471,N_21243,N_21386);
or U21472 (N_21472,N_21248,N_21232);
or U21473 (N_21473,N_21373,N_21252);
or U21474 (N_21474,N_21274,N_21224);
xor U21475 (N_21475,N_21368,N_21220);
nand U21476 (N_21476,N_21285,N_21322);
and U21477 (N_21477,N_21268,N_21392);
and U21478 (N_21478,N_21284,N_21335);
nor U21479 (N_21479,N_21325,N_21217);
and U21480 (N_21480,N_21225,N_21385);
or U21481 (N_21481,N_21330,N_21253);
nor U21482 (N_21482,N_21221,N_21303);
nand U21483 (N_21483,N_21291,N_21279);
and U21484 (N_21484,N_21271,N_21233);
or U21485 (N_21485,N_21398,N_21254);
nand U21486 (N_21486,N_21339,N_21354);
and U21487 (N_21487,N_21228,N_21218);
nand U21488 (N_21488,N_21369,N_21213);
xor U21489 (N_21489,N_21236,N_21397);
or U21490 (N_21490,N_21246,N_21238);
xnor U21491 (N_21491,N_21344,N_21300);
xnor U21492 (N_21492,N_21231,N_21289);
and U21493 (N_21493,N_21305,N_21277);
nand U21494 (N_21494,N_21223,N_21381);
or U21495 (N_21495,N_21293,N_21336);
xor U21496 (N_21496,N_21306,N_21345);
nand U21497 (N_21497,N_21301,N_21288);
xor U21498 (N_21498,N_21338,N_21244);
or U21499 (N_21499,N_21317,N_21282);
or U21500 (N_21500,N_21230,N_21296);
and U21501 (N_21501,N_21226,N_21306);
xnor U21502 (N_21502,N_21323,N_21395);
and U21503 (N_21503,N_21234,N_21225);
nand U21504 (N_21504,N_21376,N_21247);
and U21505 (N_21505,N_21311,N_21358);
nand U21506 (N_21506,N_21370,N_21390);
nand U21507 (N_21507,N_21204,N_21238);
and U21508 (N_21508,N_21247,N_21256);
nor U21509 (N_21509,N_21365,N_21305);
or U21510 (N_21510,N_21230,N_21379);
and U21511 (N_21511,N_21278,N_21204);
and U21512 (N_21512,N_21337,N_21344);
and U21513 (N_21513,N_21247,N_21344);
nor U21514 (N_21514,N_21348,N_21261);
nor U21515 (N_21515,N_21260,N_21265);
xnor U21516 (N_21516,N_21331,N_21291);
and U21517 (N_21517,N_21362,N_21386);
nor U21518 (N_21518,N_21317,N_21256);
nor U21519 (N_21519,N_21305,N_21383);
nand U21520 (N_21520,N_21369,N_21309);
nand U21521 (N_21521,N_21273,N_21397);
nor U21522 (N_21522,N_21399,N_21279);
nand U21523 (N_21523,N_21351,N_21282);
nand U21524 (N_21524,N_21355,N_21371);
and U21525 (N_21525,N_21305,N_21282);
or U21526 (N_21526,N_21240,N_21388);
and U21527 (N_21527,N_21349,N_21306);
nand U21528 (N_21528,N_21272,N_21314);
xor U21529 (N_21529,N_21326,N_21313);
nand U21530 (N_21530,N_21251,N_21335);
and U21531 (N_21531,N_21211,N_21274);
nand U21532 (N_21532,N_21296,N_21250);
nor U21533 (N_21533,N_21327,N_21303);
nor U21534 (N_21534,N_21302,N_21320);
and U21535 (N_21535,N_21209,N_21253);
or U21536 (N_21536,N_21257,N_21306);
xor U21537 (N_21537,N_21277,N_21246);
xor U21538 (N_21538,N_21215,N_21313);
or U21539 (N_21539,N_21295,N_21371);
nand U21540 (N_21540,N_21311,N_21281);
xor U21541 (N_21541,N_21399,N_21221);
xor U21542 (N_21542,N_21343,N_21368);
xnor U21543 (N_21543,N_21326,N_21395);
nand U21544 (N_21544,N_21365,N_21319);
or U21545 (N_21545,N_21222,N_21281);
or U21546 (N_21546,N_21281,N_21275);
nand U21547 (N_21547,N_21252,N_21345);
nand U21548 (N_21548,N_21281,N_21241);
and U21549 (N_21549,N_21210,N_21312);
nor U21550 (N_21550,N_21210,N_21217);
xnor U21551 (N_21551,N_21356,N_21396);
or U21552 (N_21552,N_21213,N_21291);
nand U21553 (N_21553,N_21307,N_21279);
and U21554 (N_21554,N_21286,N_21280);
and U21555 (N_21555,N_21324,N_21207);
xnor U21556 (N_21556,N_21278,N_21247);
or U21557 (N_21557,N_21254,N_21395);
nor U21558 (N_21558,N_21267,N_21387);
and U21559 (N_21559,N_21224,N_21360);
nor U21560 (N_21560,N_21324,N_21339);
nor U21561 (N_21561,N_21324,N_21316);
and U21562 (N_21562,N_21294,N_21370);
nand U21563 (N_21563,N_21374,N_21381);
nor U21564 (N_21564,N_21350,N_21206);
xnor U21565 (N_21565,N_21358,N_21370);
xor U21566 (N_21566,N_21300,N_21380);
xor U21567 (N_21567,N_21230,N_21251);
and U21568 (N_21568,N_21242,N_21341);
and U21569 (N_21569,N_21279,N_21244);
xnor U21570 (N_21570,N_21275,N_21289);
nand U21571 (N_21571,N_21239,N_21338);
nor U21572 (N_21572,N_21370,N_21253);
nand U21573 (N_21573,N_21207,N_21325);
or U21574 (N_21574,N_21242,N_21262);
or U21575 (N_21575,N_21233,N_21320);
or U21576 (N_21576,N_21366,N_21259);
or U21577 (N_21577,N_21313,N_21353);
xor U21578 (N_21578,N_21217,N_21264);
nand U21579 (N_21579,N_21351,N_21376);
nand U21580 (N_21580,N_21391,N_21273);
nor U21581 (N_21581,N_21294,N_21306);
nor U21582 (N_21582,N_21303,N_21237);
and U21583 (N_21583,N_21349,N_21327);
xor U21584 (N_21584,N_21242,N_21240);
nor U21585 (N_21585,N_21301,N_21370);
and U21586 (N_21586,N_21260,N_21300);
and U21587 (N_21587,N_21217,N_21361);
xor U21588 (N_21588,N_21330,N_21236);
nor U21589 (N_21589,N_21279,N_21380);
or U21590 (N_21590,N_21315,N_21313);
nor U21591 (N_21591,N_21251,N_21284);
or U21592 (N_21592,N_21274,N_21245);
and U21593 (N_21593,N_21309,N_21273);
nor U21594 (N_21594,N_21350,N_21327);
nor U21595 (N_21595,N_21359,N_21277);
nor U21596 (N_21596,N_21276,N_21234);
nand U21597 (N_21597,N_21316,N_21361);
xnor U21598 (N_21598,N_21338,N_21291);
nor U21599 (N_21599,N_21342,N_21378);
nand U21600 (N_21600,N_21530,N_21542);
nand U21601 (N_21601,N_21484,N_21446);
nor U21602 (N_21602,N_21409,N_21463);
or U21603 (N_21603,N_21493,N_21414);
nand U21604 (N_21604,N_21568,N_21522);
xor U21605 (N_21605,N_21574,N_21471);
nand U21606 (N_21606,N_21591,N_21475);
or U21607 (N_21607,N_21564,N_21435);
xnor U21608 (N_21608,N_21427,N_21528);
nand U21609 (N_21609,N_21527,N_21506);
nor U21610 (N_21610,N_21592,N_21407);
nand U21611 (N_21611,N_21533,N_21408);
or U21612 (N_21612,N_21469,N_21425);
nand U21613 (N_21613,N_21400,N_21460);
and U21614 (N_21614,N_21500,N_21501);
and U21615 (N_21615,N_21468,N_21454);
or U21616 (N_21616,N_21441,N_21518);
xnor U21617 (N_21617,N_21562,N_21520);
and U21618 (N_21618,N_21431,N_21481);
and U21619 (N_21619,N_21554,N_21413);
xor U21620 (N_21620,N_21491,N_21442);
nor U21621 (N_21621,N_21581,N_21443);
and U21622 (N_21622,N_21423,N_21496);
xnor U21623 (N_21623,N_21585,N_21565);
and U21624 (N_21624,N_21590,N_21444);
and U21625 (N_21625,N_21464,N_21438);
and U21626 (N_21626,N_21452,N_21473);
xor U21627 (N_21627,N_21434,N_21449);
xor U21628 (N_21628,N_21466,N_21429);
nor U21629 (N_21629,N_21428,N_21558);
nor U21630 (N_21630,N_21453,N_21439);
xnor U21631 (N_21631,N_21432,N_21509);
and U21632 (N_21632,N_21461,N_21476);
nor U21633 (N_21633,N_21552,N_21597);
xnor U21634 (N_21634,N_21417,N_21508);
or U21635 (N_21635,N_21456,N_21516);
nor U21636 (N_21636,N_21436,N_21477);
nor U21637 (N_21637,N_21594,N_21513);
xor U21638 (N_21638,N_21497,N_21563);
nor U21639 (N_21639,N_21521,N_21448);
xor U21640 (N_21640,N_21503,N_21412);
nor U21641 (N_21641,N_21499,N_21487);
or U21642 (N_21642,N_21517,N_21437);
nor U21643 (N_21643,N_21587,N_21515);
or U21644 (N_21644,N_21571,N_21538);
and U21645 (N_21645,N_21405,N_21485);
nand U21646 (N_21646,N_21573,N_21422);
and U21647 (N_21647,N_21512,N_21575);
xor U21648 (N_21648,N_21589,N_21459);
or U21649 (N_21649,N_21539,N_21540);
nand U21650 (N_21650,N_21507,N_21545);
xnor U21651 (N_21651,N_21553,N_21596);
or U21652 (N_21652,N_21483,N_21572);
nand U21653 (N_21653,N_21451,N_21566);
nand U21654 (N_21654,N_21495,N_21544);
xnor U21655 (N_21655,N_21482,N_21547);
xor U21656 (N_21656,N_21549,N_21465);
xor U21657 (N_21657,N_21579,N_21582);
and U21658 (N_21658,N_21599,N_21535);
nand U21659 (N_21659,N_21467,N_21598);
and U21660 (N_21660,N_21430,N_21494);
nor U21661 (N_21661,N_21505,N_21531);
and U21662 (N_21662,N_21593,N_21424);
nor U21663 (N_21663,N_21404,N_21478);
nor U21664 (N_21664,N_21526,N_21498);
nand U21665 (N_21665,N_21480,N_21567);
nand U21666 (N_21666,N_21523,N_21474);
nand U21667 (N_21667,N_21541,N_21457);
xnor U21668 (N_21668,N_21559,N_21455);
or U21669 (N_21669,N_21570,N_21411);
xnor U21670 (N_21670,N_21536,N_21557);
xnor U21671 (N_21671,N_21556,N_21504);
xor U21672 (N_21672,N_21534,N_21458);
xor U21673 (N_21673,N_21402,N_21489);
nand U21674 (N_21674,N_21578,N_21595);
or U21675 (N_21675,N_21514,N_21421);
and U21676 (N_21676,N_21416,N_21445);
nand U21677 (N_21677,N_21492,N_21401);
nor U21678 (N_21678,N_21410,N_21486);
and U21679 (N_21679,N_21546,N_21418);
nand U21680 (N_21680,N_21551,N_21488);
nor U21681 (N_21681,N_21519,N_21586);
nor U21682 (N_21682,N_21555,N_21502);
nor U21683 (N_21683,N_21433,N_21550);
or U21684 (N_21684,N_21525,N_21450);
xor U21685 (N_21685,N_21560,N_21537);
nor U21686 (N_21686,N_21548,N_21584);
nor U21687 (N_21687,N_21561,N_21415);
nand U21688 (N_21688,N_21470,N_21576);
or U21689 (N_21689,N_21583,N_21577);
xnor U21690 (N_21690,N_21472,N_21479);
xnor U21691 (N_21691,N_21580,N_21543);
nand U21692 (N_21692,N_21426,N_21462);
nand U21693 (N_21693,N_21529,N_21569);
nand U21694 (N_21694,N_21490,N_21511);
and U21695 (N_21695,N_21524,N_21588);
xor U21696 (N_21696,N_21420,N_21510);
nor U21697 (N_21697,N_21419,N_21403);
nor U21698 (N_21698,N_21532,N_21440);
or U21699 (N_21699,N_21406,N_21447);
and U21700 (N_21700,N_21587,N_21460);
nor U21701 (N_21701,N_21584,N_21439);
nand U21702 (N_21702,N_21506,N_21541);
nor U21703 (N_21703,N_21432,N_21507);
nand U21704 (N_21704,N_21403,N_21522);
and U21705 (N_21705,N_21551,N_21425);
and U21706 (N_21706,N_21524,N_21557);
and U21707 (N_21707,N_21465,N_21408);
and U21708 (N_21708,N_21469,N_21507);
xnor U21709 (N_21709,N_21543,N_21526);
and U21710 (N_21710,N_21595,N_21570);
nand U21711 (N_21711,N_21454,N_21490);
or U21712 (N_21712,N_21501,N_21464);
and U21713 (N_21713,N_21529,N_21450);
nand U21714 (N_21714,N_21433,N_21551);
or U21715 (N_21715,N_21511,N_21432);
xor U21716 (N_21716,N_21413,N_21522);
nor U21717 (N_21717,N_21519,N_21427);
nand U21718 (N_21718,N_21505,N_21526);
and U21719 (N_21719,N_21489,N_21407);
and U21720 (N_21720,N_21583,N_21402);
nand U21721 (N_21721,N_21481,N_21496);
nand U21722 (N_21722,N_21538,N_21455);
and U21723 (N_21723,N_21428,N_21555);
nor U21724 (N_21724,N_21598,N_21419);
or U21725 (N_21725,N_21415,N_21457);
or U21726 (N_21726,N_21597,N_21541);
nand U21727 (N_21727,N_21422,N_21458);
and U21728 (N_21728,N_21589,N_21576);
xnor U21729 (N_21729,N_21512,N_21592);
and U21730 (N_21730,N_21510,N_21498);
nand U21731 (N_21731,N_21402,N_21500);
nor U21732 (N_21732,N_21477,N_21467);
xor U21733 (N_21733,N_21521,N_21400);
nand U21734 (N_21734,N_21530,N_21441);
xor U21735 (N_21735,N_21507,N_21557);
xnor U21736 (N_21736,N_21515,N_21534);
xnor U21737 (N_21737,N_21484,N_21562);
nand U21738 (N_21738,N_21512,N_21591);
or U21739 (N_21739,N_21500,N_21533);
nand U21740 (N_21740,N_21554,N_21572);
nor U21741 (N_21741,N_21435,N_21566);
nor U21742 (N_21742,N_21420,N_21583);
and U21743 (N_21743,N_21583,N_21460);
xnor U21744 (N_21744,N_21454,N_21558);
xnor U21745 (N_21745,N_21436,N_21509);
nor U21746 (N_21746,N_21407,N_21515);
xor U21747 (N_21747,N_21455,N_21415);
xnor U21748 (N_21748,N_21417,N_21585);
nand U21749 (N_21749,N_21446,N_21452);
nand U21750 (N_21750,N_21540,N_21417);
and U21751 (N_21751,N_21567,N_21505);
nand U21752 (N_21752,N_21417,N_21526);
or U21753 (N_21753,N_21592,N_21588);
nand U21754 (N_21754,N_21482,N_21422);
xor U21755 (N_21755,N_21436,N_21478);
or U21756 (N_21756,N_21517,N_21483);
and U21757 (N_21757,N_21550,N_21458);
nor U21758 (N_21758,N_21532,N_21448);
xor U21759 (N_21759,N_21598,N_21402);
xnor U21760 (N_21760,N_21503,N_21599);
nor U21761 (N_21761,N_21562,N_21501);
nand U21762 (N_21762,N_21585,N_21562);
nor U21763 (N_21763,N_21461,N_21406);
nor U21764 (N_21764,N_21539,N_21551);
or U21765 (N_21765,N_21599,N_21545);
or U21766 (N_21766,N_21420,N_21449);
and U21767 (N_21767,N_21542,N_21502);
and U21768 (N_21768,N_21590,N_21439);
or U21769 (N_21769,N_21468,N_21475);
nand U21770 (N_21770,N_21558,N_21484);
and U21771 (N_21771,N_21572,N_21509);
xor U21772 (N_21772,N_21404,N_21447);
or U21773 (N_21773,N_21412,N_21508);
and U21774 (N_21774,N_21401,N_21402);
xnor U21775 (N_21775,N_21442,N_21426);
xnor U21776 (N_21776,N_21549,N_21474);
nand U21777 (N_21777,N_21593,N_21586);
nand U21778 (N_21778,N_21529,N_21444);
or U21779 (N_21779,N_21468,N_21446);
nor U21780 (N_21780,N_21556,N_21552);
and U21781 (N_21781,N_21569,N_21599);
xnor U21782 (N_21782,N_21458,N_21568);
nor U21783 (N_21783,N_21463,N_21579);
nand U21784 (N_21784,N_21501,N_21549);
xor U21785 (N_21785,N_21456,N_21503);
xnor U21786 (N_21786,N_21569,N_21575);
xnor U21787 (N_21787,N_21561,N_21548);
or U21788 (N_21788,N_21525,N_21434);
nand U21789 (N_21789,N_21534,N_21504);
xnor U21790 (N_21790,N_21589,N_21429);
nand U21791 (N_21791,N_21561,N_21517);
xor U21792 (N_21792,N_21495,N_21498);
nor U21793 (N_21793,N_21482,N_21584);
xnor U21794 (N_21794,N_21528,N_21592);
nor U21795 (N_21795,N_21467,N_21504);
or U21796 (N_21796,N_21500,N_21448);
xnor U21797 (N_21797,N_21435,N_21538);
nor U21798 (N_21798,N_21462,N_21418);
and U21799 (N_21799,N_21441,N_21468);
nand U21800 (N_21800,N_21777,N_21792);
and U21801 (N_21801,N_21674,N_21708);
nor U21802 (N_21802,N_21681,N_21783);
nand U21803 (N_21803,N_21725,N_21680);
nand U21804 (N_21804,N_21616,N_21627);
nor U21805 (N_21805,N_21633,N_21671);
nand U21806 (N_21806,N_21658,N_21799);
or U21807 (N_21807,N_21669,N_21763);
nor U21808 (N_21808,N_21682,N_21751);
nand U21809 (N_21809,N_21702,N_21698);
or U21810 (N_21810,N_21764,N_21768);
and U21811 (N_21811,N_21743,N_21664);
nand U21812 (N_21812,N_21793,N_21614);
or U21813 (N_21813,N_21735,N_21677);
xor U21814 (N_21814,N_21619,N_21626);
and U21815 (N_21815,N_21731,N_21718);
nor U21816 (N_21816,N_21608,N_21625);
nor U21817 (N_21817,N_21646,N_21772);
nor U21818 (N_21818,N_21696,N_21632);
or U21819 (N_21819,N_21700,N_21752);
and U21820 (N_21820,N_21756,N_21606);
xnor U21821 (N_21821,N_21791,N_21683);
and U21822 (N_21822,N_21761,N_21788);
and U21823 (N_21823,N_21732,N_21612);
and U21824 (N_21824,N_21733,N_21621);
nand U21825 (N_21825,N_21607,N_21659);
or U21826 (N_21826,N_21650,N_21631);
xnor U21827 (N_21827,N_21609,N_21647);
or U21828 (N_21828,N_21666,N_21766);
and U21829 (N_21829,N_21762,N_21712);
nand U21830 (N_21830,N_21637,N_21635);
or U21831 (N_21831,N_21667,N_21651);
and U21832 (N_21832,N_21736,N_21748);
nor U21833 (N_21833,N_21789,N_21711);
nand U21834 (N_21834,N_21796,N_21781);
and U21835 (N_21835,N_21740,N_21717);
nand U21836 (N_21836,N_21730,N_21727);
xnor U21837 (N_21837,N_21604,N_21729);
nand U21838 (N_21838,N_21737,N_21794);
nand U21839 (N_21839,N_21774,N_21655);
xnor U21840 (N_21840,N_21678,N_21784);
nor U21841 (N_21841,N_21689,N_21685);
or U21842 (N_21842,N_21780,N_21779);
nor U21843 (N_21843,N_21746,N_21786);
or U21844 (N_21844,N_21684,N_21721);
xor U21845 (N_21845,N_21744,N_21640);
nand U21846 (N_21846,N_21691,N_21798);
and U21847 (N_21847,N_21723,N_21636);
xor U21848 (N_21848,N_21770,N_21715);
or U21849 (N_21849,N_21672,N_21716);
nand U21850 (N_21850,N_21734,N_21634);
xor U21851 (N_21851,N_21600,N_21755);
nor U21852 (N_21852,N_21645,N_21617);
and U21853 (N_21853,N_21653,N_21676);
nand U21854 (N_21854,N_21693,N_21639);
nor U21855 (N_21855,N_21710,N_21760);
xor U21856 (N_21856,N_21648,N_21652);
or U21857 (N_21857,N_21785,N_21724);
and U21858 (N_21858,N_21765,N_21690);
xnor U21859 (N_21859,N_21704,N_21714);
xor U21860 (N_21860,N_21782,N_21787);
or U21861 (N_21861,N_21602,N_21668);
and U21862 (N_21862,N_21726,N_21750);
or U21863 (N_21863,N_21643,N_21638);
nor U21864 (N_21864,N_21699,N_21620);
nor U21865 (N_21865,N_21670,N_21661);
nor U21866 (N_21866,N_21739,N_21757);
or U21867 (N_21867,N_21679,N_21611);
and U21868 (N_21868,N_21613,N_21697);
nand U21869 (N_21869,N_21623,N_21665);
or U21870 (N_21870,N_21622,N_21705);
or U21871 (N_21871,N_21642,N_21759);
nand U21872 (N_21872,N_21618,N_21707);
nand U21873 (N_21873,N_21713,N_21722);
nand U21874 (N_21874,N_21629,N_21728);
or U21875 (N_21875,N_21686,N_21641);
and U21876 (N_21876,N_21797,N_21701);
xor U21877 (N_21877,N_21706,N_21654);
nor U21878 (N_21878,N_21790,N_21601);
or U21879 (N_21879,N_21719,N_21758);
or U21880 (N_21880,N_21741,N_21773);
nor U21881 (N_21881,N_21742,N_21695);
or U21882 (N_21882,N_21687,N_21775);
nand U21883 (N_21883,N_21610,N_21747);
nor U21884 (N_21884,N_21660,N_21778);
xnor U21885 (N_21885,N_21603,N_21624);
xor U21886 (N_21886,N_21605,N_21649);
xor U21887 (N_21887,N_21656,N_21795);
nor U21888 (N_21888,N_21771,N_21630);
nand U21889 (N_21889,N_21754,N_21753);
nand U21890 (N_21890,N_21662,N_21692);
or U21891 (N_21891,N_21769,N_21657);
and U21892 (N_21892,N_21628,N_21644);
and U21893 (N_21893,N_21703,N_21767);
xnor U21894 (N_21894,N_21663,N_21749);
nand U21895 (N_21895,N_21688,N_21738);
nor U21896 (N_21896,N_21720,N_21673);
and U21897 (N_21897,N_21675,N_21694);
or U21898 (N_21898,N_21615,N_21776);
nand U21899 (N_21899,N_21745,N_21709);
nand U21900 (N_21900,N_21699,N_21704);
nor U21901 (N_21901,N_21651,N_21677);
or U21902 (N_21902,N_21648,N_21732);
nor U21903 (N_21903,N_21717,N_21612);
xnor U21904 (N_21904,N_21602,N_21681);
xnor U21905 (N_21905,N_21678,N_21642);
nand U21906 (N_21906,N_21790,N_21692);
xnor U21907 (N_21907,N_21633,N_21772);
or U21908 (N_21908,N_21621,N_21680);
nand U21909 (N_21909,N_21776,N_21693);
nand U21910 (N_21910,N_21769,N_21641);
nand U21911 (N_21911,N_21626,N_21709);
and U21912 (N_21912,N_21612,N_21727);
nor U21913 (N_21913,N_21715,N_21603);
nor U21914 (N_21914,N_21646,N_21667);
nand U21915 (N_21915,N_21771,N_21753);
xnor U21916 (N_21916,N_21669,N_21648);
and U21917 (N_21917,N_21627,N_21677);
xor U21918 (N_21918,N_21690,N_21643);
xnor U21919 (N_21919,N_21757,N_21600);
and U21920 (N_21920,N_21706,N_21761);
xnor U21921 (N_21921,N_21728,N_21666);
or U21922 (N_21922,N_21652,N_21604);
nand U21923 (N_21923,N_21746,N_21690);
or U21924 (N_21924,N_21740,N_21746);
nand U21925 (N_21925,N_21759,N_21790);
and U21926 (N_21926,N_21677,N_21699);
and U21927 (N_21927,N_21624,N_21658);
and U21928 (N_21928,N_21679,N_21730);
nor U21929 (N_21929,N_21719,N_21745);
nor U21930 (N_21930,N_21681,N_21791);
and U21931 (N_21931,N_21683,N_21787);
xor U21932 (N_21932,N_21625,N_21696);
or U21933 (N_21933,N_21634,N_21610);
nor U21934 (N_21934,N_21706,N_21638);
nand U21935 (N_21935,N_21622,N_21759);
and U21936 (N_21936,N_21668,N_21784);
xnor U21937 (N_21937,N_21795,N_21652);
nand U21938 (N_21938,N_21631,N_21673);
and U21939 (N_21939,N_21708,N_21794);
or U21940 (N_21940,N_21757,N_21688);
or U21941 (N_21941,N_21716,N_21665);
xnor U21942 (N_21942,N_21643,N_21601);
or U21943 (N_21943,N_21776,N_21744);
xor U21944 (N_21944,N_21718,N_21682);
and U21945 (N_21945,N_21641,N_21709);
nand U21946 (N_21946,N_21606,N_21711);
nand U21947 (N_21947,N_21754,N_21792);
or U21948 (N_21948,N_21722,N_21689);
and U21949 (N_21949,N_21670,N_21608);
or U21950 (N_21950,N_21710,N_21661);
xnor U21951 (N_21951,N_21676,N_21679);
nor U21952 (N_21952,N_21679,N_21708);
and U21953 (N_21953,N_21675,N_21624);
xnor U21954 (N_21954,N_21725,N_21677);
nand U21955 (N_21955,N_21669,N_21673);
nor U21956 (N_21956,N_21627,N_21776);
xnor U21957 (N_21957,N_21732,N_21708);
xor U21958 (N_21958,N_21718,N_21708);
and U21959 (N_21959,N_21758,N_21783);
nor U21960 (N_21960,N_21770,N_21677);
xor U21961 (N_21961,N_21700,N_21638);
and U21962 (N_21962,N_21677,N_21784);
or U21963 (N_21963,N_21749,N_21672);
nand U21964 (N_21964,N_21753,N_21745);
xnor U21965 (N_21965,N_21700,N_21602);
and U21966 (N_21966,N_21728,N_21770);
xnor U21967 (N_21967,N_21675,N_21644);
and U21968 (N_21968,N_21753,N_21709);
nor U21969 (N_21969,N_21764,N_21660);
nand U21970 (N_21970,N_21766,N_21742);
and U21971 (N_21971,N_21600,N_21659);
or U21972 (N_21972,N_21764,N_21676);
or U21973 (N_21973,N_21626,N_21706);
xnor U21974 (N_21974,N_21659,N_21644);
or U21975 (N_21975,N_21770,N_21650);
nand U21976 (N_21976,N_21611,N_21797);
nor U21977 (N_21977,N_21634,N_21649);
xor U21978 (N_21978,N_21619,N_21647);
nand U21979 (N_21979,N_21669,N_21732);
nor U21980 (N_21980,N_21690,N_21787);
xor U21981 (N_21981,N_21781,N_21685);
and U21982 (N_21982,N_21749,N_21658);
or U21983 (N_21983,N_21743,N_21643);
xor U21984 (N_21984,N_21721,N_21639);
nand U21985 (N_21985,N_21681,N_21773);
and U21986 (N_21986,N_21619,N_21705);
nand U21987 (N_21987,N_21652,N_21655);
xor U21988 (N_21988,N_21768,N_21671);
nor U21989 (N_21989,N_21627,N_21610);
xor U21990 (N_21990,N_21793,N_21692);
nand U21991 (N_21991,N_21643,N_21798);
nor U21992 (N_21992,N_21644,N_21714);
and U21993 (N_21993,N_21757,N_21710);
nor U21994 (N_21994,N_21735,N_21616);
nand U21995 (N_21995,N_21707,N_21639);
nand U21996 (N_21996,N_21713,N_21671);
or U21997 (N_21997,N_21786,N_21764);
xor U21998 (N_21998,N_21624,N_21742);
nand U21999 (N_21999,N_21795,N_21629);
nor U22000 (N_22000,N_21838,N_21897);
nor U22001 (N_22001,N_21855,N_21818);
or U22002 (N_22002,N_21957,N_21839);
or U22003 (N_22003,N_21862,N_21975);
nand U22004 (N_22004,N_21984,N_21942);
or U22005 (N_22005,N_21845,N_21896);
or U22006 (N_22006,N_21907,N_21873);
xor U22007 (N_22007,N_21870,N_21884);
xnor U22008 (N_22008,N_21894,N_21969);
nor U22009 (N_22009,N_21997,N_21835);
nand U22010 (N_22010,N_21893,N_21949);
xnor U22011 (N_22011,N_21970,N_21808);
and U22012 (N_22012,N_21937,N_21848);
and U22013 (N_22013,N_21974,N_21943);
xor U22014 (N_22014,N_21982,N_21924);
xnor U22015 (N_22015,N_21928,N_21864);
nand U22016 (N_22016,N_21918,N_21929);
nor U22017 (N_22017,N_21917,N_21901);
xor U22018 (N_22018,N_21846,N_21995);
xnor U22019 (N_22019,N_21939,N_21851);
or U22020 (N_22020,N_21804,N_21826);
and U22021 (N_22021,N_21944,N_21978);
nor U22022 (N_22022,N_21852,N_21932);
or U22023 (N_22023,N_21867,N_21954);
xnor U22024 (N_22024,N_21821,N_21996);
and U22025 (N_22025,N_21966,N_21948);
nor U22026 (N_22026,N_21993,N_21859);
nand U22027 (N_22027,N_21908,N_21813);
nand U22028 (N_22028,N_21880,N_21881);
xor U22029 (N_22029,N_21865,N_21874);
nor U22030 (N_22030,N_21815,N_21910);
nand U22031 (N_22031,N_21999,N_21895);
and U22032 (N_22032,N_21827,N_21951);
xnor U22033 (N_22033,N_21931,N_21946);
nor U22034 (N_22034,N_21922,N_21983);
or U22035 (N_22035,N_21915,N_21926);
xor U22036 (N_22036,N_21806,N_21869);
and U22037 (N_22037,N_21913,N_21909);
or U22038 (N_22038,N_21930,N_21921);
and U22039 (N_22039,N_21860,N_21812);
and U22040 (N_22040,N_21847,N_21967);
or U22041 (N_22041,N_21986,N_21803);
or U22042 (N_22042,N_21875,N_21866);
nand U22043 (N_22043,N_21971,N_21998);
xnor U22044 (N_22044,N_21950,N_21962);
nor U22045 (N_22045,N_21833,N_21842);
or U22046 (N_22046,N_21817,N_21941);
nand U22047 (N_22047,N_21994,N_21871);
or U22048 (N_22048,N_21912,N_21976);
nor U22049 (N_22049,N_21840,N_21952);
or U22050 (N_22050,N_21800,N_21883);
or U22051 (N_22051,N_21919,N_21816);
nand U22052 (N_22052,N_21825,N_21843);
nor U22053 (N_22053,N_21853,N_21927);
nand U22054 (N_22054,N_21953,N_21963);
xnor U22055 (N_22055,N_21824,N_21923);
or U22056 (N_22056,N_21981,N_21837);
xnor U22057 (N_22057,N_21876,N_21899);
nor U22058 (N_22058,N_21872,N_21977);
nor U22059 (N_22059,N_21905,N_21955);
nor U22060 (N_22060,N_21900,N_21947);
xor U22061 (N_22061,N_21904,N_21965);
or U22062 (N_22062,N_21925,N_21933);
nor U22063 (N_22063,N_21885,N_21911);
xnor U22064 (N_22064,N_21903,N_21809);
and U22065 (N_22065,N_21822,N_21879);
or U22066 (N_22066,N_21914,N_21811);
xor U22067 (N_22067,N_21814,N_21945);
xor U22068 (N_22068,N_21834,N_21830);
and U22069 (N_22069,N_21841,N_21861);
nor U22070 (N_22070,N_21958,N_21831);
xor U22071 (N_22071,N_21819,N_21979);
or U22072 (N_22072,N_21857,N_21989);
nor U22073 (N_22073,N_21844,N_21888);
and U22074 (N_22074,N_21940,N_21985);
and U22075 (N_22075,N_21882,N_21935);
and U22076 (N_22076,N_21906,N_21936);
and U22077 (N_22077,N_21902,N_21877);
or U22078 (N_22078,N_21990,N_21887);
nor U22079 (N_22079,N_21898,N_21991);
nor U22080 (N_22080,N_21972,N_21956);
nor U22081 (N_22081,N_21889,N_21805);
or U22082 (N_22082,N_21987,N_21802);
or U22083 (N_22083,N_21938,N_21964);
nand U22084 (N_22084,N_21832,N_21858);
or U22085 (N_22085,N_21836,N_21916);
and U22086 (N_22086,N_21828,N_21934);
nor U22087 (N_22087,N_21988,N_21890);
xnor U22088 (N_22088,N_21920,N_21968);
and U22089 (N_22089,N_21820,N_21807);
xnor U22090 (N_22090,N_21961,N_21992);
xor U22091 (N_22091,N_21854,N_21886);
xor U22092 (N_22092,N_21980,N_21850);
nor U22093 (N_22093,N_21878,N_21849);
nand U22094 (N_22094,N_21892,N_21863);
and U22095 (N_22095,N_21973,N_21891);
nor U22096 (N_22096,N_21959,N_21829);
nand U22097 (N_22097,N_21960,N_21801);
or U22098 (N_22098,N_21810,N_21868);
nand U22099 (N_22099,N_21823,N_21856);
nor U22100 (N_22100,N_21907,N_21830);
nor U22101 (N_22101,N_21890,N_21977);
xnor U22102 (N_22102,N_21925,N_21960);
or U22103 (N_22103,N_21987,N_21963);
or U22104 (N_22104,N_21973,N_21932);
nor U22105 (N_22105,N_21818,N_21805);
xor U22106 (N_22106,N_21928,N_21917);
and U22107 (N_22107,N_21869,N_21909);
nor U22108 (N_22108,N_21930,N_21886);
xor U22109 (N_22109,N_21925,N_21929);
or U22110 (N_22110,N_21953,N_21904);
xnor U22111 (N_22111,N_21891,N_21944);
nand U22112 (N_22112,N_21974,N_21912);
or U22113 (N_22113,N_21831,N_21972);
nor U22114 (N_22114,N_21846,N_21871);
nand U22115 (N_22115,N_21924,N_21995);
xnor U22116 (N_22116,N_21838,N_21922);
nor U22117 (N_22117,N_21951,N_21965);
xnor U22118 (N_22118,N_21964,N_21994);
or U22119 (N_22119,N_21861,N_21947);
or U22120 (N_22120,N_21963,N_21831);
or U22121 (N_22121,N_21826,N_21825);
or U22122 (N_22122,N_21817,N_21925);
nand U22123 (N_22123,N_21870,N_21914);
nand U22124 (N_22124,N_21877,N_21903);
xnor U22125 (N_22125,N_21898,N_21966);
nand U22126 (N_22126,N_21992,N_21901);
and U22127 (N_22127,N_21959,N_21802);
and U22128 (N_22128,N_21976,N_21911);
xor U22129 (N_22129,N_21807,N_21981);
or U22130 (N_22130,N_21814,N_21834);
or U22131 (N_22131,N_21971,N_21987);
nor U22132 (N_22132,N_21959,N_21826);
or U22133 (N_22133,N_21998,N_21837);
or U22134 (N_22134,N_21877,N_21929);
nor U22135 (N_22135,N_21874,N_21824);
and U22136 (N_22136,N_21926,N_21869);
xnor U22137 (N_22137,N_21986,N_21907);
nor U22138 (N_22138,N_21975,N_21994);
nand U22139 (N_22139,N_21805,N_21918);
and U22140 (N_22140,N_21946,N_21877);
nand U22141 (N_22141,N_21989,N_21860);
and U22142 (N_22142,N_21967,N_21839);
or U22143 (N_22143,N_21988,N_21832);
or U22144 (N_22144,N_21921,N_21873);
or U22145 (N_22145,N_21876,N_21854);
and U22146 (N_22146,N_21823,N_21929);
or U22147 (N_22147,N_21939,N_21856);
xnor U22148 (N_22148,N_21871,N_21875);
xnor U22149 (N_22149,N_21877,N_21879);
or U22150 (N_22150,N_21962,N_21889);
or U22151 (N_22151,N_21959,N_21992);
or U22152 (N_22152,N_21996,N_21973);
or U22153 (N_22153,N_21896,N_21952);
and U22154 (N_22154,N_21952,N_21875);
and U22155 (N_22155,N_21879,N_21973);
nand U22156 (N_22156,N_21865,N_21875);
xnor U22157 (N_22157,N_21950,N_21837);
or U22158 (N_22158,N_21933,N_21916);
and U22159 (N_22159,N_21865,N_21919);
nand U22160 (N_22160,N_21865,N_21904);
or U22161 (N_22161,N_21878,N_21918);
nor U22162 (N_22162,N_21859,N_21963);
and U22163 (N_22163,N_21952,N_21941);
nand U22164 (N_22164,N_21873,N_21895);
xnor U22165 (N_22165,N_21845,N_21970);
nor U22166 (N_22166,N_21928,N_21838);
nand U22167 (N_22167,N_21985,N_21832);
xor U22168 (N_22168,N_21873,N_21981);
and U22169 (N_22169,N_21937,N_21813);
nand U22170 (N_22170,N_21810,N_21877);
nand U22171 (N_22171,N_21982,N_21899);
xor U22172 (N_22172,N_21941,N_21842);
xor U22173 (N_22173,N_21947,N_21939);
xnor U22174 (N_22174,N_21873,N_21968);
and U22175 (N_22175,N_21863,N_21826);
xor U22176 (N_22176,N_21988,N_21894);
nand U22177 (N_22177,N_21953,N_21946);
xnor U22178 (N_22178,N_21855,N_21883);
or U22179 (N_22179,N_21852,N_21925);
nand U22180 (N_22180,N_21835,N_21940);
nand U22181 (N_22181,N_21999,N_21855);
and U22182 (N_22182,N_21982,N_21846);
and U22183 (N_22183,N_21934,N_21992);
nor U22184 (N_22184,N_21951,N_21881);
nand U22185 (N_22185,N_21878,N_21827);
and U22186 (N_22186,N_21808,N_21899);
and U22187 (N_22187,N_21810,N_21997);
nor U22188 (N_22188,N_21993,N_21818);
nand U22189 (N_22189,N_21823,N_21858);
or U22190 (N_22190,N_21855,N_21895);
nor U22191 (N_22191,N_21961,N_21911);
nand U22192 (N_22192,N_21971,N_21852);
or U22193 (N_22193,N_21979,N_21959);
or U22194 (N_22194,N_21856,N_21990);
or U22195 (N_22195,N_21918,N_21864);
or U22196 (N_22196,N_21869,N_21920);
or U22197 (N_22197,N_21924,N_21805);
xnor U22198 (N_22198,N_21902,N_21856);
or U22199 (N_22199,N_21876,N_21892);
xnor U22200 (N_22200,N_22179,N_22050);
xnor U22201 (N_22201,N_22017,N_22058);
nand U22202 (N_22202,N_22014,N_22121);
xor U22203 (N_22203,N_22194,N_22141);
xor U22204 (N_22204,N_22146,N_22186);
nor U22205 (N_22205,N_22090,N_22076);
nor U22206 (N_22206,N_22159,N_22052);
xor U22207 (N_22207,N_22118,N_22087);
and U22208 (N_22208,N_22197,N_22022);
nand U22209 (N_22209,N_22130,N_22075);
or U22210 (N_22210,N_22184,N_22077);
or U22211 (N_22211,N_22104,N_22199);
and U22212 (N_22212,N_22092,N_22117);
nand U22213 (N_22213,N_22019,N_22166);
or U22214 (N_22214,N_22127,N_22085);
nor U22215 (N_22215,N_22115,N_22031);
and U22216 (N_22216,N_22078,N_22182);
or U22217 (N_22217,N_22148,N_22057);
xor U22218 (N_22218,N_22047,N_22142);
xor U22219 (N_22219,N_22154,N_22097);
or U22220 (N_22220,N_22125,N_22151);
nor U22221 (N_22221,N_22028,N_22086);
and U22222 (N_22222,N_22144,N_22176);
or U22223 (N_22223,N_22089,N_22059);
nor U22224 (N_22224,N_22039,N_22070);
nor U22225 (N_22225,N_22023,N_22114);
nand U22226 (N_22226,N_22049,N_22034);
or U22227 (N_22227,N_22063,N_22064);
or U22228 (N_22228,N_22020,N_22160);
and U22229 (N_22229,N_22068,N_22080);
nand U22230 (N_22230,N_22196,N_22084);
nor U22231 (N_22231,N_22046,N_22177);
xnor U22232 (N_22232,N_22113,N_22012);
xnor U22233 (N_22233,N_22072,N_22171);
or U22234 (N_22234,N_22073,N_22140);
nand U22235 (N_22235,N_22133,N_22003);
and U22236 (N_22236,N_22095,N_22139);
xnor U22237 (N_22237,N_22183,N_22067);
or U22238 (N_22238,N_22054,N_22102);
xor U22239 (N_22239,N_22172,N_22103);
nand U22240 (N_22240,N_22007,N_22198);
nand U22241 (N_22241,N_22093,N_22165);
nor U22242 (N_22242,N_22045,N_22018);
xnor U22243 (N_22243,N_22116,N_22147);
and U22244 (N_22244,N_22101,N_22191);
xnor U22245 (N_22245,N_22035,N_22037);
or U22246 (N_22246,N_22106,N_22026);
nor U22247 (N_22247,N_22163,N_22021);
or U22248 (N_22248,N_22002,N_22053);
and U22249 (N_22249,N_22061,N_22043);
xnor U22250 (N_22250,N_22190,N_22074);
or U22251 (N_22251,N_22000,N_22156);
nand U22252 (N_22252,N_22005,N_22162);
or U22253 (N_22253,N_22155,N_22025);
or U22254 (N_22254,N_22110,N_22055);
nor U22255 (N_22255,N_22042,N_22016);
nand U22256 (N_22256,N_22189,N_22030);
nor U22257 (N_22257,N_22149,N_22187);
nor U22258 (N_22258,N_22137,N_22013);
or U22259 (N_22259,N_22044,N_22006);
or U22260 (N_22260,N_22066,N_22181);
and U22261 (N_22261,N_22145,N_22100);
or U22262 (N_22262,N_22071,N_22004);
xnor U22263 (N_22263,N_22107,N_22131);
xor U22264 (N_22264,N_22065,N_22040);
nor U22265 (N_22265,N_22123,N_22112);
and U22266 (N_22266,N_22193,N_22134);
nor U22267 (N_22267,N_22029,N_22136);
nor U22268 (N_22268,N_22094,N_22081);
and U22269 (N_22269,N_22024,N_22119);
nand U22270 (N_22270,N_22188,N_22180);
and U22271 (N_22271,N_22011,N_22041);
xor U22272 (N_22272,N_22169,N_22082);
xnor U22273 (N_22273,N_22056,N_22175);
nor U22274 (N_22274,N_22124,N_22109);
nor U22275 (N_22275,N_22126,N_22108);
and U22276 (N_22276,N_22143,N_22069);
xor U22277 (N_22277,N_22174,N_22150);
or U22278 (N_22278,N_22164,N_22008);
and U22279 (N_22279,N_22091,N_22051);
nor U22280 (N_22280,N_22083,N_22168);
xor U22281 (N_22281,N_22079,N_22048);
xor U22282 (N_22282,N_22132,N_22122);
xor U22283 (N_22283,N_22157,N_22105);
nor U22284 (N_22284,N_22001,N_22096);
nor U22285 (N_22285,N_22170,N_22027);
nor U22286 (N_22286,N_22161,N_22088);
and U22287 (N_22287,N_22060,N_22135);
or U22288 (N_22288,N_22192,N_22167);
nand U22289 (N_22289,N_22153,N_22032);
nand U22290 (N_22290,N_22010,N_22158);
or U22291 (N_22291,N_22036,N_22098);
nor U22292 (N_22292,N_22015,N_22120);
nand U22293 (N_22293,N_22033,N_22099);
nor U22294 (N_22294,N_22111,N_22128);
or U22295 (N_22295,N_22038,N_22173);
and U22296 (N_22296,N_22138,N_22009);
xor U22297 (N_22297,N_22178,N_22152);
and U22298 (N_22298,N_22195,N_22062);
nand U22299 (N_22299,N_22185,N_22129);
nand U22300 (N_22300,N_22133,N_22013);
nor U22301 (N_22301,N_22010,N_22022);
nor U22302 (N_22302,N_22105,N_22037);
nand U22303 (N_22303,N_22016,N_22084);
nand U22304 (N_22304,N_22175,N_22017);
and U22305 (N_22305,N_22009,N_22070);
xnor U22306 (N_22306,N_22138,N_22010);
xor U22307 (N_22307,N_22121,N_22126);
xnor U22308 (N_22308,N_22194,N_22094);
xnor U22309 (N_22309,N_22092,N_22109);
nand U22310 (N_22310,N_22198,N_22005);
or U22311 (N_22311,N_22155,N_22068);
or U22312 (N_22312,N_22107,N_22095);
and U22313 (N_22313,N_22055,N_22018);
or U22314 (N_22314,N_22085,N_22163);
or U22315 (N_22315,N_22140,N_22107);
nand U22316 (N_22316,N_22138,N_22153);
or U22317 (N_22317,N_22143,N_22053);
nor U22318 (N_22318,N_22078,N_22159);
nand U22319 (N_22319,N_22052,N_22042);
nor U22320 (N_22320,N_22039,N_22151);
nor U22321 (N_22321,N_22066,N_22012);
and U22322 (N_22322,N_22095,N_22068);
xor U22323 (N_22323,N_22017,N_22116);
and U22324 (N_22324,N_22007,N_22183);
xnor U22325 (N_22325,N_22049,N_22024);
nand U22326 (N_22326,N_22031,N_22020);
nor U22327 (N_22327,N_22103,N_22068);
and U22328 (N_22328,N_22001,N_22199);
xor U22329 (N_22329,N_22045,N_22003);
or U22330 (N_22330,N_22127,N_22170);
or U22331 (N_22331,N_22131,N_22137);
nor U22332 (N_22332,N_22140,N_22118);
or U22333 (N_22333,N_22164,N_22144);
or U22334 (N_22334,N_22190,N_22162);
xor U22335 (N_22335,N_22044,N_22117);
and U22336 (N_22336,N_22104,N_22021);
and U22337 (N_22337,N_22031,N_22196);
xnor U22338 (N_22338,N_22017,N_22077);
and U22339 (N_22339,N_22057,N_22152);
xor U22340 (N_22340,N_22012,N_22044);
xor U22341 (N_22341,N_22083,N_22107);
nand U22342 (N_22342,N_22085,N_22157);
and U22343 (N_22343,N_22145,N_22069);
nor U22344 (N_22344,N_22025,N_22159);
nand U22345 (N_22345,N_22125,N_22163);
xnor U22346 (N_22346,N_22065,N_22057);
nand U22347 (N_22347,N_22103,N_22127);
or U22348 (N_22348,N_22074,N_22081);
or U22349 (N_22349,N_22122,N_22049);
nor U22350 (N_22350,N_22165,N_22109);
or U22351 (N_22351,N_22053,N_22057);
xnor U22352 (N_22352,N_22026,N_22014);
or U22353 (N_22353,N_22048,N_22158);
xnor U22354 (N_22354,N_22114,N_22037);
or U22355 (N_22355,N_22055,N_22080);
or U22356 (N_22356,N_22047,N_22119);
and U22357 (N_22357,N_22046,N_22161);
and U22358 (N_22358,N_22146,N_22024);
and U22359 (N_22359,N_22031,N_22093);
or U22360 (N_22360,N_22184,N_22130);
or U22361 (N_22361,N_22144,N_22110);
nor U22362 (N_22362,N_22057,N_22039);
nor U22363 (N_22363,N_22017,N_22041);
or U22364 (N_22364,N_22093,N_22189);
nor U22365 (N_22365,N_22128,N_22065);
nand U22366 (N_22366,N_22078,N_22154);
xnor U22367 (N_22367,N_22013,N_22141);
and U22368 (N_22368,N_22100,N_22133);
xor U22369 (N_22369,N_22104,N_22043);
nand U22370 (N_22370,N_22023,N_22144);
nand U22371 (N_22371,N_22125,N_22033);
nand U22372 (N_22372,N_22089,N_22113);
xnor U22373 (N_22373,N_22189,N_22193);
and U22374 (N_22374,N_22044,N_22098);
and U22375 (N_22375,N_22040,N_22123);
nand U22376 (N_22376,N_22127,N_22158);
nor U22377 (N_22377,N_22065,N_22041);
and U22378 (N_22378,N_22000,N_22153);
nor U22379 (N_22379,N_22008,N_22044);
xor U22380 (N_22380,N_22121,N_22136);
nor U22381 (N_22381,N_22060,N_22163);
nand U22382 (N_22382,N_22162,N_22067);
nand U22383 (N_22383,N_22137,N_22035);
nand U22384 (N_22384,N_22194,N_22041);
or U22385 (N_22385,N_22090,N_22034);
nand U22386 (N_22386,N_22072,N_22019);
or U22387 (N_22387,N_22095,N_22010);
xnor U22388 (N_22388,N_22141,N_22058);
and U22389 (N_22389,N_22081,N_22018);
nor U22390 (N_22390,N_22180,N_22004);
nand U22391 (N_22391,N_22065,N_22011);
or U22392 (N_22392,N_22170,N_22062);
xor U22393 (N_22393,N_22010,N_22058);
nor U22394 (N_22394,N_22099,N_22019);
and U22395 (N_22395,N_22008,N_22165);
nand U22396 (N_22396,N_22111,N_22030);
nand U22397 (N_22397,N_22184,N_22135);
nand U22398 (N_22398,N_22148,N_22091);
and U22399 (N_22399,N_22032,N_22011);
and U22400 (N_22400,N_22233,N_22356);
or U22401 (N_22401,N_22282,N_22371);
and U22402 (N_22402,N_22340,N_22226);
nand U22403 (N_22403,N_22230,N_22345);
nor U22404 (N_22404,N_22241,N_22310);
nor U22405 (N_22405,N_22318,N_22325);
and U22406 (N_22406,N_22301,N_22288);
nand U22407 (N_22407,N_22245,N_22341);
nand U22408 (N_22408,N_22270,N_22374);
nor U22409 (N_22409,N_22332,N_22229);
xnor U22410 (N_22410,N_22266,N_22331);
nor U22411 (N_22411,N_22242,N_22315);
nor U22412 (N_22412,N_22367,N_22231);
xnor U22413 (N_22413,N_22394,N_22292);
and U22414 (N_22414,N_22380,N_22295);
or U22415 (N_22415,N_22364,N_22204);
or U22416 (N_22416,N_22283,N_22333);
or U22417 (N_22417,N_22389,N_22207);
or U22418 (N_22418,N_22381,N_22272);
or U22419 (N_22419,N_22335,N_22323);
and U22420 (N_22420,N_22312,N_22299);
nor U22421 (N_22421,N_22317,N_22251);
nand U22422 (N_22422,N_22281,N_22308);
xnor U22423 (N_22423,N_22214,N_22348);
xor U22424 (N_22424,N_22327,N_22240);
and U22425 (N_22425,N_22361,N_22338);
xnor U22426 (N_22426,N_22238,N_22225);
nand U22427 (N_22427,N_22239,N_22391);
xor U22428 (N_22428,N_22213,N_22291);
xnor U22429 (N_22429,N_22290,N_22390);
nand U22430 (N_22430,N_22396,N_22215);
or U22431 (N_22431,N_22309,N_22393);
nand U22432 (N_22432,N_22320,N_22379);
xnor U22433 (N_22433,N_22383,N_22307);
nor U22434 (N_22434,N_22398,N_22293);
nand U22435 (N_22435,N_22277,N_22205);
and U22436 (N_22436,N_22336,N_22275);
or U22437 (N_22437,N_22375,N_22246);
nand U22438 (N_22438,N_22206,N_22313);
or U22439 (N_22439,N_22280,N_22399);
or U22440 (N_22440,N_22321,N_22286);
or U22441 (N_22441,N_22250,N_22287);
xor U22442 (N_22442,N_22300,N_22330);
nor U22443 (N_22443,N_22339,N_22324);
and U22444 (N_22444,N_22319,N_22284);
xor U22445 (N_22445,N_22358,N_22261);
and U22446 (N_22446,N_22202,N_22349);
xor U22447 (N_22447,N_22237,N_22328);
nor U22448 (N_22448,N_22298,N_22397);
and U22449 (N_22449,N_22216,N_22264);
nand U22450 (N_22450,N_22259,N_22350);
and U22451 (N_22451,N_22297,N_22363);
and U22452 (N_22452,N_22279,N_22235);
nor U22453 (N_22453,N_22218,N_22201);
and U22454 (N_22454,N_22278,N_22354);
xor U22455 (N_22455,N_22377,N_22252);
nand U22456 (N_22456,N_22342,N_22247);
or U22457 (N_22457,N_22285,N_22343);
or U22458 (N_22458,N_22228,N_22269);
nand U22459 (N_22459,N_22256,N_22362);
or U22460 (N_22460,N_22337,N_22200);
nand U22461 (N_22461,N_22232,N_22357);
and U22462 (N_22462,N_22257,N_22376);
nor U22463 (N_22463,N_22373,N_22388);
nor U22464 (N_22464,N_22360,N_22227);
xor U22465 (N_22465,N_22211,N_22347);
or U22466 (N_22466,N_22344,N_22271);
or U22467 (N_22467,N_22289,N_22255);
nor U22468 (N_22468,N_22276,N_22316);
and U22469 (N_22469,N_22346,N_22222);
xnor U22470 (N_22470,N_22334,N_22209);
xor U22471 (N_22471,N_22365,N_22359);
nand U22472 (N_22472,N_22258,N_22387);
nor U22473 (N_22473,N_22305,N_22273);
or U22474 (N_22474,N_22248,N_22352);
xor U22475 (N_22475,N_22224,N_22234);
and U22476 (N_22476,N_22385,N_22355);
nand U22477 (N_22477,N_22386,N_22217);
xor U22478 (N_22478,N_22203,N_22384);
nand U22479 (N_22479,N_22351,N_22296);
nand U22480 (N_22480,N_22260,N_22210);
xor U22481 (N_22481,N_22268,N_22306);
xnor U22482 (N_22482,N_22326,N_22294);
or U22483 (N_22483,N_22353,N_22303);
or U22484 (N_22484,N_22372,N_22265);
nor U22485 (N_22485,N_22236,N_22223);
nand U22486 (N_22486,N_22302,N_22322);
and U22487 (N_22487,N_22311,N_22378);
nor U22488 (N_22488,N_22244,N_22382);
or U22489 (N_22489,N_22263,N_22314);
xnor U22490 (N_22490,N_22274,N_22220);
nor U22491 (N_22491,N_22243,N_22329);
and U22492 (N_22492,N_22370,N_22249);
nor U22493 (N_22493,N_22221,N_22254);
nand U22494 (N_22494,N_22219,N_22253);
nor U22495 (N_22495,N_22366,N_22304);
and U22496 (N_22496,N_22212,N_22369);
or U22497 (N_22497,N_22368,N_22208);
nand U22498 (N_22498,N_22395,N_22262);
xnor U22499 (N_22499,N_22267,N_22392);
xor U22500 (N_22500,N_22348,N_22221);
xor U22501 (N_22501,N_22224,N_22265);
or U22502 (N_22502,N_22217,N_22343);
and U22503 (N_22503,N_22247,N_22290);
and U22504 (N_22504,N_22313,N_22285);
xnor U22505 (N_22505,N_22274,N_22378);
or U22506 (N_22506,N_22357,N_22217);
xor U22507 (N_22507,N_22334,N_22236);
or U22508 (N_22508,N_22200,N_22348);
nand U22509 (N_22509,N_22389,N_22205);
and U22510 (N_22510,N_22260,N_22369);
or U22511 (N_22511,N_22361,N_22354);
xnor U22512 (N_22512,N_22382,N_22329);
nor U22513 (N_22513,N_22340,N_22385);
and U22514 (N_22514,N_22274,N_22221);
nand U22515 (N_22515,N_22260,N_22285);
nand U22516 (N_22516,N_22209,N_22213);
xnor U22517 (N_22517,N_22249,N_22269);
nor U22518 (N_22518,N_22333,N_22358);
or U22519 (N_22519,N_22358,N_22235);
and U22520 (N_22520,N_22355,N_22248);
nor U22521 (N_22521,N_22337,N_22225);
nand U22522 (N_22522,N_22265,N_22368);
and U22523 (N_22523,N_22235,N_22334);
nor U22524 (N_22524,N_22355,N_22329);
nor U22525 (N_22525,N_22378,N_22310);
xnor U22526 (N_22526,N_22335,N_22375);
xnor U22527 (N_22527,N_22330,N_22251);
and U22528 (N_22528,N_22213,N_22271);
or U22529 (N_22529,N_22379,N_22301);
or U22530 (N_22530,N_22357,N_22261);
or U22531 (N_22531,N_22298,N_22384);
nor U22532 (N_22532,N_22278,N_22211);
xnor U22533 (N_22533,N_22304,N_22210);
nor U22534 (N_22534,N_22327,N_22377);
xor U22535 (N_22535,N_22377,N_22259);
nor U22536 (N_22536,N_22298,N_22379);
nor U22537 (N_22537,N_22286,N_22381);
nand U22538 (N_22538,N_22344,N_22379);
nand U22539 (N_22539,N_22336,N_22364);
xor U22540 (N_22540,N_22278,N_22341);
nor U22541 (N_22541,N_22256,N_22346);
nand U22542 (N_22542,N_22238,N_22385);
nor U22543 (N_22543,N_22312,N_22258);
xnor U22544 (N_22544,N_22370,N_22341);
or U22545 (N_22545,N_22354,N_22258);
nor U22546 (N_22546,N_22267,N_22398);
nor U22547 (N_22547,N_22303,N_22237);
xor U22548 (N_22548,N_22264,N_22395);
nand U22549 (N_22549,N_22355,N_22226);
nand U22550 (N_22550,N_22347,N_22275);
xnor U22551 (N_22551,N_22222,N_22305);
xnor U22552 (N_22552,N_22212,N_22221);
nor U22553 (N_22553,N_22329,N_22376);
nand U22554 (N_22554,N_22365,N_22228);
nor U22555 (N_22555,N_22210,N_22366);
nor U22556 (N_22556,N_22204,N_22335);
nand U22557 (N_22557,N_22289,N_22332);
and U22558 (N_22558,N_22218,N_22318);
and U22559 (N_22559,N_22361,N_22283);
xnor U22560 (N_22560,N_22329,N_22212);
or U22561 (N_22561,N_22333,N_22234);
nor U22562 (N_22562,N_22228,N_22319);
and U22563 (N_22563,N_22300,N_22253);
xnor U22564 (N_22564,N_22243,N_22316);
and U22565 (N_22565,N_22325,N_22300);
and U22566 (N_22566,N_22224,N_22387);
xor U22567 (N_22567,N_22313,N_22376);
and U22568 (N_22568,N_22314,N_22267);
nor U22569 (N_22569,N_22387,N_22209);
nand U22570 (N_22570,N_22373,N_22263);
nor U22571 (N_22571,N_22308,N_22234);
nor U22572 (N_22572,N_22263,N_22326);
nor U22573 (N_22573,N_22341,N_22354);
nor U22574 (N_22574,N_22338,N_22259);
xnor U22575 (N_22575,N_22241,N_22228);
or U22576 (N_22576,N_22242,N_22327);
nor U22577 (N_22577,N_22314,N_22309);
and U22578 (N_22578,N_22256,N_22211);
and U22579 (N_22579,N_22298,N_22372);
nand U22580 (N_22580,N_22241,N_22247);
xnor U22581 (N_22581,N_22211,N_22356);
and U22582 (N_22582,N_22385,N_22229);
nor U22583 (N_22583,N_22308,N_22337);
nand U22584 (N_22584,N_22205,N_22292);
xnor U22585 (N_22585,N_22222,N_22351);
or U22586 (N_22586,N_22292,N_22354);
nand U22587 (N_22587,N_22266,N_22304);
nand U22588 (N_22588,N_22265,N_22211);
and U22589 (N_22589,N_22322,N_22258);
xnor U22590 (N_22590,N_22276,N_22248);
nor U22591 (N_22591,N_22207,N_22353);
xnor U22592 (N_22592,N_22348,N_22366);
nand U22593 (N_22593,N_22310,N_22291);
nor U22594 (N_22594,N_22274,N_22364);
and U22595 (N_22595,N_22285,N_22252);
or U22596 (N_22596,N_22285,N_22361);
or U22597 (N_22597,N_22226,N_22313);
and U22598 (N_22598,N_22287,N_22268);
nand U22599 (N_22599,N_22383,N_22247);
nand U22600 (N_22600,N_22487,N_22552);
xnor U22601 (N_22601,N_22475,N_22402);
and U22602 (N_22602,N_22417,N_22509);
xnor U22603 (N_22603,N_22459,N_22473);
xor U22604 (N_22604,N_22478,N_22565);
nand U22605 (N_22605,N_22585,N_22546);
xor U22606 (N_22606,N_22582,N_22500);
or U22607 (N_22607,N_22533,N_22465);
or U22608 (N_22608,N_22492,N_22597);
nand U22609 (N_22609,N_22470,N_22522);
nand U22610 (N_22610,N_22404,N_22513);
or U22611 (N_22611,N_22457,N_22499);
xnor U22612 (N_22612,N_22434,N_22431);
nand U22613 (N_22613,N_22575,N_22535);
nand U22614 (N_22614,N_22550,N_22577);
xnor U22615 (N_22615,N_22409,N_22527);
nor U22616 (N_22616,N_22521,N_22598);
nand U22617 (N_22617,N_22589,N_22541);
and U22618 (N_22618,N_22496,N_22490);
or U22619 (N_22619,N_22573,N_22440);
or U22620 (N_22620,N_22551,N_22429);
nand U22621 (N_22621,N_22588,N_22427);
xnor U22622 (N_22622,N_22566,N_22558);
and U22623 (N_22623,N_22413,N_22471);
nor U22624 (N_22624,N_22415,N_22572);
nand U22625 (N_22625,N_22532,N_22439);
xor U22626 (N_22626,N_22591,N_22469);
nor U22627 (N_22627,N_22489,N_22537);
or U22628 (N_22628,N_22435,N_22481);
xor U22629 (N_22629,N_22548,N_22514);
nor U22630 (N_22630,N_22557,N_22410);
or U22631 (N_22631,N_22425,N_22512);
xor U22632 (N_22632,N_22599,N_22594);
nand U22633 (N_22633,N_22511,N_22505);
nand U22634 (N_22634,N_22460,N_22507);
or U22635 (N_22635,N_22408,N_22424);
nor U22636 (N_22636,N_22556,N_22497);
nand U22637 (N_22637,N_22531,N_22484);
nor U22638 (N_22638,N_22405,N_22559);
nand U22639 (N_22639,N_22420,N_22549);
or U22640 (N_22640,N_22430,N_22596);
or U22641 (N_22641,N_22508,N_22561);
nor U22642 (N_22642,N_22504,N_22567);
xor U22643 (N_22643,N_22547,N_22580);
nor U22644 (N_22644,N_22510,N_22401);
or U22645 (N_22645,N_22526,N_22477);
or U22646 (N_22646,N_22542,N_22432);
and U22647 (N_22647,N_22540,N_22570);
or U22648 (N_22648,N_22563,N_22506);
xnor U22649 (N_22649,N_22555,N_22486);
or U22650 (N_22650,N_22560,N_22441);
or U22651 (N_22651,N_22433,N_22586);
or U22652 (N_22652,N_22450,N_22587);
nand U22653 (N_22653,N_22437,N_22468);
nand U22654 (N_22654,N_22528,N_22464);
and U22655 (N_22655,N_22592,N_22517);
xnor U22656 (N_22656,N_22519,N_22406);
and U22657 (N_22657,N_22480,N_22458);
and U22658 (N_22658,N_22466,N_22423);
nand U22659 (N_22659,N_22456,N_22538);
xor U22660 (N_22660,N_22422,N_22524);
nor U22661 (N_22661,N_22571,N_22447);
or U22662 (N_22662,N_22448,N_22529);
or U22663 (N_22663,N_22523,N_22564);
xor U22664 (N_22664,N_22426,N_22474);
nor U22665 (N_22665,N_22515,N_22462);
nor U22666 (N_22666,N_22530,N_22576);
nor U22667 (N_22667,N_22467,N_22449);
nand U22668 (N_22668,N_22438,N_22562);
or U22669 (N_22669,N_22488,N_22491);
xnor U22670 (N_22670,N_22493,N_22412);
nor U22671 (N_22671,N_22498,N_22442);
xor U22672 (N_22672,N_22483,N_22411);
and U22673 (N_22673,N_22403,N_22502);
or U22674 (N_22674,N_22544,N_22539);
and U22675 (N_22675,N_22578,N_22482);
xor U22676 (N_22676,N_22516,N_22503);
or U22677 (N_22677,N_22501,N_22414);
xnor U22678 (N_22678,N_22461,N_22579);
xnor U22679 (N_22679,N_22543,N_22400);
nor U22680 (N_22680,N_22428,N_22495);
xor U22681 (N_22681,N_22494,N_22581);
nor U22682 (N_22682,N_22463,N_22407);
or U22683 (N_22683,N_22553,N_22590);
xor U22684 (N_22684,N_22453,N_22476);
xnor U22685 (N_22685,N_22593,N_22454);
xnor U22686 (N_22686,N_22451,N_22595);
nor U22687 (N_22687,N_22421,N_22534);
and U22688 (N_22688,N_22583,N_22419);
or U22689 (N_22689,N_22443,N_22479);
or U22690 (N_22690,N_22445,N_22518);
and U22691 (N_22691,N_22554,N_22545);
xnor U22692 (N_22692,N_22455,N_22446);
nor U22693 (N_22693,N_22452,N_22418);
nand U22694 (N_22694,N_22568,N_22485);
xnor U22695 (N_22695,N_22569,N_22416);
or U22696 (N_22696,N_22472,N_22520);
xnor U22697 (N_22697,N_22536,N_22525);
nor U22698 (N_22698,N_22574,N_22584);
and U22699 (N_22699,N_22436,N_22444);
xnor U22700 (N_22700,N_22594,N_22538);
nand U22701 (N_22701,N_22433,N_22423);
nand U22702 (N_22702,N_22476,N_22402);
and U22703 (N_22703,N_22529,N_22538);
and U22704 (N_22704,N_22582,N_22594);
nand U22705 (N_22705,N_22424,N_22526);
nand U22706 (N_22706,N_22460,N_22533);
xnor U22707 (N_22707,N_22510,N_22514);
and U22708 (N_22708,N_22518,N_22594);
and U22709 (N_22709,N_22514,N_22594);
and U22710 (N_22710,N_22438,N_22596);
nand U22711 (N_22711,N_22521,N_22482);
and U22712 (N_22712,N_22536,N_22482);
nand U22713 (N_22713,N_22481,N_22434);
or U22714 (N_22714,N_22427,N_22419);
nand U22715 (N_22715,N_22528,N_22479);
or U22716 (N_22716,N_22472,N_22577);
and U22717 (N_22717,N_22532,N_22556);
nand U22718 (N_22718,N_22504,N_22490);
and U22719 (N_22719,N_22425,N_22562);
nand U22720 (N_22720,N_22519,N_22512);
and U22721 (N_22721,N_22580,N_22491);
or U22722 (N_22722,N_22403,N_22412);
xor U22723 (N_22723,N_22437,N_22593);
or U22724 (N_22724,N_22476,N_22478);
and U22725 (N_22725,N_22488,N_22501);
nor U22726 (N_22726,N_22547,N_22563);
and U22727 (N_22727,N_22593,N_22465);
and U22728 (N_22728,N_22479,N_22518);
xor U22729 (N_22729,N_22569,N_22540);
nand U22730 (N_22730,N_22547,N_22422);
or U22731 (N_22731,N_22414,N_22573);
nor U22732 (N_22732,N_22463,N_22510);
and U22733 (N_22733,N_22418,N_22473);
and U22734 (N_22734,N_22575,N_22522);
or U22735 (N_22735,N_22504,N_22447);
or U22736 (N_22736,N_22587,N_22540);
or U22737 (N_22737,N_22474,N_22594);
and U22738 (N_22738,N_22475,N_22419);
or U22739 (N_22739,N_22401,N_22552);
or U22740 (N_22740,N_22577,N_22529);
nand U22741 (N_22741,N_22586,N_22478);
or U22742 (N_22742,N_22564,N_22510);
nor U22743 (N_22743,N_22417,N_22544);
and U22744 (N_22744,N_22434,N_22401);
nor U22745 (N_22745,N_22463,N_22479);
xor U22746 (N_22746,N_22555,N_22520);
nand U22747 (N_22747,N_22448,N_22429);
nand U22748 (N_22748,N_22495,N_22538);
xnor U22749 (N_22749,N_22511,N_22464);
nor U22750 (N_22750,N_22555,N_22500);
and U22751 (N_22751,N_22586,N_22475);
xor U22752 (N_22752,N_22481,N_22538);
nor U22753 (N_22753,N_22547,N_22405);
and U22754 (N_22754,N_22430,N_22571);
or U22755 (N_22755,N_22491,N_22418);
nand U22756 (N_22756,N_22462,N_22530);
nor U22757 (N_22757,N_22418,N_22434);
and U22758 (N_22758,N_22489,N_22547);
nand U22759 (N_22759,N_22407,N_22521);
nand U22760 (N_22760,N_22506,N_22488);
and U22761 (N_22761,N_22535,N_22407);
nor U22762 (N_22762,N_22582,N_22578);
nor U22763 (N_22763,N_22483,N_22423);
or U22764 (N_22764,N_22476,N_22429);
nand U22765 (N_22765,N_22472,N_22412);
or U22766 (N_22766,N_22575,N_22493);
or U22767 (N_22767,N_22414,N_22599);
nor U22768 (N_22768,N_22514,N_22462);
xor U22769 (N_22769,N_22416,N_22434);
nor U22770 (N_22770,N_22469,N_22548);
or U22771 (N_22771,N_22475,N_22469);
xnor U22772 (N_22772,N_22572,N_22447);
and U22773 (N_22773,N_22437,N_22457);
and U22774 (N_22774,N_22554,N_22494);
and U22775 (N_22775,N_22576,N_22548);
nor U22776 (N_22776,N_22473,N_22485);
nor U22777 (N_22777,N_22552,N_22433);
nor U22778 (N_22778,N_22561,N_22429);
nand U22779 (N_22779,N_22537,N_22516);
nand U22780 (N_22780,N_22415,N_22551);
and U22781 (N_22781,N_22461,N_22594);
nor U22782 (N_22782,N_22553,N_22498);
nor U22783 (N_22783,N_22450,N_22501);
nor U22784 (N_22784,N_22407,N_22576);
and U22785 (N_22785,N_22508,N_22457);
nor U22786 (N_22786,N_22456,N_22540);
and U22787 (N_22787,N_22586,N_22583);
xnor U22788 (N_22788,N_22493,N_22572);
and U22789 (N_22789,N_22495,N_22493);
nor U22790 (N_22790,N_22520,N_22516);
nor U22791 (N_22791,N_22428,N_22403);
nand U22792 (N_22792,N_22505,N_22594);
nand U22793 (N_22793,N_22434,N_22583);
nor U22794 (N_22794,N_22598,N_22506);
and U22795 (N_22795,N_22503,N_22551);
or U22796 (N_22796,N_22521,N_22541);
nor U22797 (N_22797,N_22441,N_22469);
nor U22798 (N_22798,N_22468,N_22446);
nand U22799 (N_22799,N_22576,N_22567);
xor U22800 (N_22800,N_22786,N_22741);
nor U22801 (N_22801,N_22670,N_22742);
or U22802 (N_22802,N_22606,N_22608);
and U22803 (N_22803,N_22623,N_22745);
xnor U22804 (N_22804,N_22733,N_22689);
or U22805 (N_22805,N_22692,N_22641);
or U22806 (N_22806,N_22752,N_22624);
nor U22807 (N_22807,N_22725,N_22798);
nand U22808 (N_22808,N_22613,N_22644);
nand U22809 (N_22809,N_22609,N_22612);
nor U22810 (N_22810,N_22674,N_22764);
xnor U22811 (N_22811,N_22707,N_22796);
nor U22812 (N_22812,N_22767,N_22638);
nand U22813 (N_22813,N_22738,N_22756);
xnor U22814 (N_22814,N_22646,N_22712);
nand U22815 (N_22815,N_22617,N_22761);
xor U22816 (N_22816,N_22797,N_22766);
and U22817 (N_22817,N_22619,N_22622);
nand U22818 (N_22818,N_22732,N_22603);
nor U22819 (N_22819,N_22653,N_22727);
or U22820 (N_22820,N_22634,N_22749);
xnor U22821 (N_22821,N_22677,N_22630);
or U22822 (N_22822,N_22770,N_22691);
xnor U22823 (N_22823,N_22690,N_22649);
xor U22824 (N_22824,N_22771,N_22779);
and U22825 (N_22825,N_22718,N_22753);
nor U22826 (N_22826,N_22668,N_22792);
nand U22827 (N_22827,N_22729,N_22610);
xnor U22828 (N_22828,N_22679,N_22618);
xor U22829 (N_22829,N_22794,N_22743);
and U22830 (N_22830,N_22789,N_22628);
nand U22831 (N_22831,N_22639,N_22751);
and U22832 (N_22832,N_22774,N_22731);
or U22833 (N_22833,N_22775,N_22723);
and U22834 (N_22834,N_22715,N_22784);
nor U22835 (N_22835,N_22680,N_22759);
and U22836 (N_22836,N_22795,N_22714);
or U22837 (N_22837,N_22686,N_22654);
and U22838 (N_22838,N_22720,N_22768);
nor U22839 (N_22839,N_22688,N_22671);
and U22840 (N_22840,N_22744,N_22710);
xor U22841 (N_22841,N_22781,N_22735);
or U22842 (N_22842,N_22746,N_22685);
nor U22843 (N_22843,N_22625,N_22696);
nand U22844 (N_22844,N_22728,N_22650);
or U22845 (N_22845,N_22736,N_22785);
xor U22846 (N_22846,N_22683,N_22621);
or U22847 (N_22847,N_22698,N_22645);
xnor U22848 (N_22848,N_22661,N_22665);
nand U22849 (N_22849,N_22787,N_22701);
and U22850 (N_22850,N_22703,N_22765);
or U22851 (N_22851,N_22694,N_22730);
and U22852 (N_22852,N_22636,N_22758);
or U22853 (N_22853,N_22705,N_22763);
xor U22854 (N_22854,N_22709,N_22687);
and U22855 (N_22855,N_22658,N_22607);
or U22856 (N_22856,N_22600,N_22669);
or U22857 (N_22857,N_22706,N_22783);
nor U22858 (N_22858,N_22776,N_22711);
nor U22859 (N_22859,N_22755,N_22663);
nand U22860 (N_22860,N_22602,N_22791);
and U22861 (N_22861,N_22660,N_22702);
or U22862 (N_22862,N_22635,N_22632);
xnor U22863 (N_22863,N_22793,N_22611);
or U22864 (N_22864,N_22724,N_22722);
and U22865 (N_22865,N_22652,N_22648);
nand U22866 (N_22866,N_22666,N_22762);
nor U22867 (N_22867,N_22633,N_22773);
nand U22868 (N_22868,N_22643,N_22662);
nor U22869 (N_22869,N_22778,N_22748);
or U22870 (N_22870,N_22726,N_22620);
nand U22871 (N_22871,N_22708,N_22676);
or U22872 (N_22872,N_22664,N_22673);
or U22873 (N_22873,N_22626,N_22642);
nor U22874 (N_22874,N_22737,N_22695);
xnor U22875 (N_22875,N_22655,N_22682);
nand U22876 (N_22876,N_22721,N_22769);
and U22877 (N_22877,N_22604,N_22757);
and U22878 (N_22878,N_22647,N_22699);
nor U22879 (N_22879,N_22693,N_22734);
and U22880 (N_22880,N_22713,N_22678);
nand U22881 (N_22881,N_22601,N_22651);
and U22882 (N_22882,N_22799,N_22750);
or U22883 (N_22883,N_22717,N_22790);
or U22884 (N_22884,N_22780,N_22656);
nand U22885 (N_22885,N_22629,N_22747);
and U22886 (N_22886,N_22772,N_22716);
and U22887 (N_22887,N_22631,N_22614);
and U22888 (N_22888,N_22681,N_22616);
nor U22889 (N_22889,N_22627,N_22700);
and U22890 (N_22890,N_22657,N_22605);
and U22891 (N_22891,N_22777,N_22704);
or U22892 (N_22892,N_22684,N_22788);
nor U22893 (N_22893,N_22782,N_22667);
nand U22894 (N_22894,N_22740,N_22697);
xor U22895 (N_22895,N_22640,N_22719);
nand U22896 (N_22896,N_22739,N_22615);
xnor U22897 (N_22897,N_22675,N_22754);
nor U22898 (N_22898,N_22637,N_22659);
nor U22899 (N_22899,N_22760,N_22672);
or U22900 (N_22900,N_22713,N_22673);
nand U22901 (N_22901,N_22615,N_22683);
xnor U22902 (N_22902,N_22613,N_22776);
or U22903 (N_22903,N_22745,N_22757);
or U22904 (N_22904,N_22755,N_22787);
nor U22905 (N_22905,N_22609,N_22765);
and U22906 (N_22906,N_22600,N_22770);
and U22907 (N_22907,N_22678,N_22734);
nand U22908 (N_22908,N_22744,N_22620);
nor U22909 (N_22909,N_22600,N_22711);
xnor U22910 (N_22910,N_22769,N_22713);
nor U22911 (N_22911,N_22649,N_22681);
xnor U22912 (N_22912,N_22778,N_22727);
nor U22913 (N_22913,N_22736,N_22625);
nand U22914 (N_22914,N_22655,N_22683);
xor U22915 (N_22915,N_22706,N_22626);
nor U22916 (N_22916,N_22795,N_22727);
or U22917 (N_22917,N_22734,N_22756);
and U22918 (N_22918,N_22668,N_22756);
or U22919 (N_22919,N_22692,N_22718);
and U22920 (N_22920,N_22661,N_22617);
nor U22921 (N_22921,N_22719,N_22679);
or U22922 (N_22922,N_22735,N_22706);
nand U22923 (N_22923,N_22727,N_22690);
nand U22924 (N_22924,N_22653,N_22613);
or U22925 (N_22925,N_22768,N_22683);
or U22926 (N_22926,N_22673,N_22722);
nor U22927 (N_22927,N_22763,N_22775);
nor U22928 (N_22928,N_22678,N_22656);
and U22929 (N_22929,N_22715,N_22718);
xor U22930 (N_22930,N_22610,N_22697);
xnor U22931 (N_22931,N_22638,N_22705);
nor U22932 (N_22932,N_22774,N_22736);
and U22933 (N_22933,N_22761,N_22647);
nor U22934 (N_22934,N_22633,N_22624);
and U22935 (N_22935,N_22693,N_22703);
or U22936 (N_22936,N_22687,N_22653);
xnor U22937 (N_22937,N_22699,N_22741);
and U22938 (N_22938,N_22641,N_22706);
or U22939 (N_22939,N_22752,N_22702);
or U22940 (N_22940,N_22791,N_22729);
nand U22941 (N_22941,N_22600,N_22609);
and U22942 (N_22942,N_22670,N_22711);
or U22943 (N_22943,N_22791,N_22633);
nor U22944 (N_22944,N_22773,N_22644);
or U22945 (N_22945,N_22754,N_22628);
or U22946 (N_22946,N_22696,N_22773);
xor U22947 (N_22947,N_22695,N_22622);
xnor U22948 (N_22948,N_22683,N_22634);
and U22949 (N_22949,N_22785,N_22702);
and U22950 (N_22950,N_22754,N_22665);
nand U22951 (N_22951,N_22736,N_22661);
xor U22952 (N_22952,N_22628,N_22790);
and U22953 (N_22953,N_22731,N_22749);
xnor U22954 (N_22954,N_22798,N_22740);
and U22955 (N_22955,N_22619,N_22611);
nor U22956 (N_22956,N_22693,N_22765);
and U22957 (N_22957,N_22779,N_22706);
nand U22958 (N_22958,N_22772,N_22621);
nand U22959 (N_22959,N_22614,N_22661);
or U22960 (N_22960,N_22610,N_22630);
xor U22961 (N_22961,N_22780,N_22639);
nand U22962 (N_22962,N_22627,N_22609);
xnor U22963 (N_22963,N_22694,N_22703);
nor U22964 (N_22964,N_22782,N_22656);
nor U22965 (N_22965,N_22736,N_22619);
or U22966 (N_22966,N_22722,N_22615);
and U22967 (N_22967,N_22635,N_22731);
xnor U22968 (N_22968,N_22644,N_22670);
xnor U22969 (N_22969,N_22760,N_22737);
xor U22970 (N_22970,N_22606,N_22760);
nor U22971 (N_22971,N_22712,N_22718);
or U22972 (N_22972,N_22770,N_22613);
nor U22973 (N_22973,N_22675,N_22635);
nor U22974 (N_22974,N_22671,N_22724);
and U22975 (N_22975,N_22664,N_22677);
or U22976 (N_22976,N_22678,N_22788);
and U22977 (N_22977,N_22684,N_22756);
xor U22978 (N_22978,N_22732,N_22654);
and U22979 (N_22979,N_22727,N_22685);
nand U22980 (N_22980,N_22763,N_22758);
nor U22981 (N_22981,N_22795,N_22715);
xor U22982 (N_22982,N_22639,N_22730);
and U22983 (N_22983,N_22677,N_22723);
nor U22984 (N_22984,N_22731,N_22745);
nand U22985 (N_22985,N_22746,N_22671);
xor U22986 (N_22986,N_22609,N_22757);
xor U22987 (N_22987,N_22734,N_22781);
and U22988 (N_22988,N_22698,N_22766);
nor U22989 (N_22989,N_22624,N_22654);
nor U22990 (N_22990,N_22646,N_22735);
nand U22991 (N_22991,N_22739,N_22688);
or U22992 (N_22992,N_22609,N_22701);
nand U22993 (N_22993,N_22630,N_22613);
nand U22994 (N_22994,N_22612,N_22796);
or U22995 (N_22995,N_22764,N_22634);
and U22996 (N_22996,N_22695,N_22751);
and U22997 (N_22997,N_22645,N_22690);
or U22998 (N_22998,N_22763,N_22614);
or U22999 (N_22999,N_22711,N_22648);
nand U23000 (N_23000,N_22928,N_22955);
nand U23001 (N_23001,N_22996,N_22815);
or U23002 (N_23002,N_22857,N_22922);
or U23003 (N_23003,N_22980,N_22887);
xnor U23004 (N_23004,N_22855,N_22945);
nand U23005 (N_23005,N_22822,N_22994);
nand U23006 (N_23006,N_22858,N_22966);
and U23007 (N_23007,N_22910,N_22842);
and U23008 (N_23008,N_22962,N_22856);
xor U23009 (N_23009,N_22847,N_22920);
and U23010 (N_23010,N_22967,N_22901);
xor U23011 (N_23011,N_22986,N_22895);
or U23012 (N_23012,N_22907,N_22829);
xnor U23013 (N_23013,N_22970,N_22894);
and U23014 (N_23014,N_22935,N_22929);
or U23015 (N_23015,N_22978,N_22818);
nor U23016 (N_23016,N_22958,N_22949);
or U23017 (N_23017,N_22806,N_22940);
and U23018 (N_23018,N_22826,N_22937);
nand U23019 (N_23019,N_22892,N_22984);
nand U23020 (N_23020,N_22805,N_22816);
xor U23021 (N_23021,N_22946,N_22942);
nand U23022 (N_23022,N_22943,N_22831);
xnor U23023 (N_23023,N_22999,N_22896);
xnor U23024 (N_23024,N_22953,N_22992);
or U23025 (N_23025,N_22979,N_22851);
xor U23026 (N_23026,N_22990,N_22915);
or U23027 (N_23027,N_22835,N_22860);
xor U23028 (N_23028,N_22874,N_22888);
xor U23029 (N_23029,N_22909,N_22933);
xor U23030 (N_23030,N_22871,N_22832);
xnor U23031 (N_23031,N_22938,N_22982);
and U23032 (N_23032,N_22939,N_22975);
or U23033 (N_23033,N_22801,N_22987);
nor U23034 (N_23034,N_22836,N_22959);
xor U23035 (N_23035,N_22820,N_22930);
and U23036 (N_23036,N_22918,N_22879);
nor U23037 (N_23037,N_22848,N_22828);
nand U23038 (N_23038,N_22889,N_22971);
or U23039 (N_23039,N_22900,N_22886);
nor U23040 (N_23040,N_22866,N_22906);
xnor U23041 (N_23041,N_22878,N_22837);
nand U23042 (N_23042,N_22903,N_22867);
or U23043 (N_23043,N_22988,N_22838);
xor U23044 (N_23044,N_22859,N_22845);
and U23045 (N_23045,N_22808,N_22811);
nand U23046 (N_23046,N_22819,N_22991);
nand U23047 (N_23047,N_22839,N_22948);
xor U23048 (N_23048,N_22985,N_22934);
and U23049 (N_23049,N_22925,N_22824);
nor U23050 (N_23050,N_22983,N_22974);
and U23051 (N_23051,N_22870,N_22981);
and U23052 (N_23052,N_22861,N_22954);
xor U23053 (N_23053,N_22926,N_22905);
nand U23054 (N_23054,N_22969,N_22814);
and U23055 (N_23055,N_22843,N_22872);
xnor U23056 (N_23056,N_22961,N_22912);
nor U23057 (N_23057,N_22883,N_22810);
xor U23058 (N_23058,N_22852,N_22932);
nor U23059 (N_23059,N_22902,N_22825);
nand U23060 (N_23060,N_22927,N_22899);
nor U23061 (N_23061,N_22951,N_22876);
and U23062 (N_23062,N_22908,N_22854);
nand U23063 (N_23063,N_22891,N_22923);
or U23064 (N_23064,N_22997,N_22863);
nand U23065 (N_23065,N_22875,N_22830);
nand U23066 (N_23066,N_22963,N_22881);
and U23067 (N_23067,N_22995,N_22827);
and U23068 (N_23068,N_22873,N_22998);
nand U23069 (N_23069,N_22952,N_22817);
nand U23070 (N_23070,N_22924,N_22917);
or U23071 (N_23071,N_22884,N_22809);
nor U23072 (N_23072,N_22823,N_22804);
xor U23073 (N_23073,N_22893,N_22913);
nand U23074 (N_23074,N_22921,N_22993);
nand U23075 (N_23075,N_22914,N_22897);
nor U23076 (N_23076,N_22841,N_22977);
nor U23077 (N_23077,N_22868,N_22898);
nand U23078 (N_23078,N_22807,N_22973);
or U23079 (N_23079,N_22853,N_22904);
or U23080 (N_23080,N_22821,N_22950);
xor U23081 (N_23081,N_22960,N_22947);
or U23082 (N_23082,N_22840,N_22965);
xor U23083 (N_23083,N_22802,N_22846);
nand U23084 (N_23084,N_22864,N_22882);
and U23085 (N_23085,N_22812,N_22936);
and U23086 (N_23086,N_22890,N_22885);
xnor U23087 (N_23087,N_22944,N_22849);
xor U23088 (N_23088,N_22869,N_22989);
nand U23089 (N_23089,N_22916,N_22862);
and U23090 (N_23090,N_22976,N_22834);
and U23091 (N_23091,N_22956,N_22850);
or U23092 (N_23092,N_22919,N_22813);
nand U23093 (N_23093,N_22844,N_22880);
nor U23094 (N_23094,N_22865,N_22972);
nand U23095 (N_23095,N_22803,N_22833);
nor U23096 (N_23096,N_22957,N_22800);
and U23097 (N_23097,N_22941,N_22931);
or U23098 (N_23098,N_22877,N_22968);
or U23099 (N_23099,N_22911,N_22964);
xor U23100 (N_23100,N_22938,N_22861);
and U23101 (N_23101,N_22865,N_22996);
xor U23102 (N_23102,N_22959,N_22880);
xnor U23103 (N_23103,N_22856,N_22929);
and U23104 (N_23104,N_22808,N_22908);
nor U23105 (N_23105,N_22898,N_22985);
xor U23106 (N_23106,N_22884,N_22870);
nor U23107 (N_23107,N_22906,N_22977);
or U23108 (N_23108,N_22940,N_22889);
nand U23109 (N_23109,N_22891,N_22863);
nor U23110 (N_23110,N_22922,N_22908);
nor U23111 (N_23111,N_22887,N_22858);
nand U23112 (N_23112,N_22885,N_22879);
and U23113 (N_23113,N_22843,N_22827);
nand U23114 (N_23114,N_22886,N_22801);
and U23115 (N_23115,N_22880,N_22877);
nor U23116 (N_23116,N_22991,N_22868);
or U23117 (N_23117,N_22901,N_22887);
and U23118 (N_23118,N_22975,N_22929);
or U23119 (N_23119,N_22949,N_22899);
nor U23120 (N_23120,N_22897,N_22901);
nand U23121 (N_23121,N_22847,N_22866);
nand U23122 (N_23122,N_22933,N_22965);
or U23123 (N_23123,N_22934,N_22962);
nand U23124 (N_23124,N_22858,N_22960);
xnor U23125 (N_23125,N_22942,N_22887);
nand U23126 (N_23126,N_22979,N_22854);
xor U23127 (N_23127,N_22957,N_22968);
nand U23128 (N_23128,N_22959,N_22913);
nand U23129 (N_23129,N_22865,N_22969);
nand U23130 (N_23130,N_22985,N_22908);
nand U23131 (N_23131,N_22917,N_22943);
nor U23132 (N_23132,N_22972,N_22846);
nor U23133 (N_23133,N_22807,N_22965);
or U23134 (N_23134,N_22860,N_22882);
xnor U23135 (N_23135,N_22995,N_22885);
xor U23136 (N_23136,N_22808,N_22834);
and U23137 (N_23137,N_22987,N_22934);
and U23138 (N_23138,N_22851,N_22802);
or U23139 (N_23139,N_22934,N_22900);
and U23140 (N_23140,N_22807,N_22951);
nor U23141 (N_23141,N_22824,N_22997);
or U23142 (N_23142,N_22866,N_22992);
or U23143 (N_23143,N_22954,N_22938);
nand U23144 (N_23144,N_22824,N_22907);
nor U23145 (N_23145,N_22997,N_22994);
xnor U23146 (N_23146,N_22813,N_22982);
or U23147 (N_23147,N_22910,N_22917);
and U23148 (N_23148,N_22908,N_22827);
nor U23149 (N_23149,N_22947,N_22921);
xor U23150 (N_23150,N_22916,N_22993);
xnor U23151 (N_23151,N_22985,N_22988);
xor U23152 (N_23152,N_22852,N_22924);
xnor U23153 (N_23153,N_22837,N_22945);
or U23154 (N_23154,N_22980,N_22854);
and U23155 (N_23155,N_22812,N_22988);
nor U23156 (N_23156,N_22854,N_22803);
xor U23157 (N_23157,N_22968,N_22890);
and U23158 (N_23158,N_22983,N_22950);
nor U23159 (N_23159,N_22924,N_22865);
nor U23160 (N_23160,N_22999,N_22991);
nor U23161 (N_23161,N_22863,N_22876);
nand U23162 (N_23162,N_22867,N_22987);
or U23163 (N_23163,N_22986,N_22983);
and U23164 (N_23164,N_22935,N_22904);
or U23165 (N_23165,N_22800,N_22890);
and U23166 (N_23166,N_22901,N_22818);
and U23167 (N_23167,N_22847,N_22800);
xor U23168 (N_23168,N_22879,N_22836);
xor U23169 (N_23169,N_22923,N_22936);
nand U23170 (N_23170,N_22844,N_22965);
or U23171 (N_23171,N_22823,N_22965);
or U23172 (N_23172,N_22807,N_22975);
nand U23173 (N_23173,N_22807,N_22901);
and U23174 (N_23174,N_22809,N_22918);
nor U23175 (N_23175,N_22925,N_22895);
or U23176 (N_23176,N_22897,N_22966);
nor U23177 (N_23177,N_22878,N_22905);
nor U23178 (N_23178,N_22811,N_22843);
and U23179 (N_23179,N_22802,N_22937);
nand U23180 (N_23180,N_22924,N_22859);
and U23181 (N_23181,N_22875,N_22944);
nand U23182 (N_23182,N_22970,N_22886);
nor U23183 (N_23183,N_22812,N_22849);
nor U23184 (N_23184,N_22927,N_22896);
nand U23185 (N_23185,N_22818,N_22825);
nor U23186 (N_23186,N_22919,N_22985);
and U23187 (N_23187,N_22847,N_22975);
nor U23188 (N_23188,N_22992,N_22854);
xor U23189 (N_23189,N_22874,N_22968);
or U23190 (N_23190,N_22954,N_22929);
or U23191 (N_23191,N_22845,N_22818);
and U23192 (N_23192,N_22914,N_22891);
and U23193 (N_23193,N_22901,N_22981);
or U23194 (N_23194,N_22976,N_22891);
nor U23195 (N_23195,N_22969,N_22916);
nor U23196 (N_23196,N_22922,N_22829);
xor U23197 (N_23197,N_22831,N_22907);
xor U23198 (N_23198,N_22857,N_22898);
or U23199 (N_23199,N_22946,N_22880);
xnor U23200 (N_23200,N_23046,N_23167);
nand U23201 (N_23201,N_23123,N_23192);
and U23202 (N_23202,N_23131,N_23010);
and U23203 (N_23203,N_23011,N_23005);
nand U23204 (N_23204,N_23060,N_23018);
or U23205 (N_23205,N_23121,N_23019);
nor U23206 (N_23206,N_23064,N_23169);
nand U23207 (N_23207,N_23109,N_23154);
and U23208 (N_23208,N_23157,N_23025);
or U23209 (N_23209,N_23139,N_23041);
nor U23210 (N_23210,N_23134,N_23116);
or U23211 (N_23211,N_23016,N_23093);
xor U23212 (N_23212,N_23124,N_23024);
nand U23213 (N_23213,N_23068,N_23120);
and U23214 (N_23214,N_23088,N_23091);
nor U23215 (N_23215,N_23115,N_23017);
nor U23216 (N_23216,N_23113,N_23171);
xor U23217 (N_23217,N_23145,N_23100);
xor U23218 (N_23218,N_23164,N_23193);
nand U23219 (N_23219,N_23151,N_23136);
and U23220 (N_23220,N_23103,N_23057);
and U23221 (N_23221,N_23158,N_23147);
xnor U23222 (N_23222,N_23178,N_23026);
nor U23223 (N_23223,N_23030,N_23022);
and U23224 (N_23224,N_23000,N_23054);
and U23225 (N_23225,N_23190,N_23127);
xor U23226 (N_23226,N_23090,N_23028);
and U23227 (N_23227,N_23066,N_23056);
nand U23228 (N_23228,N_23132,N_23050);
nand U23229 (N_23229,N_23133,N_23085);
nand U23230 (N_23230,N_23189,N_23095);
nor U23231 (N_23231,N_23034,N_23128);
xnor U23232 (N_23232,N_23153,N_23077);
and U23233 (N_23233,N_23089,N_23168);
nand U23234 (N_23234,N_23045,N_23040);
nand U23235 (N_23235,N_23082,N_23078);
nand U23236 (N_23236,N_23180,N_23195);
nand U23237 (N_23237,N_23071,N_23199);
xor U23238 (N_23238,N_23052,N_23062);
and U23239 (N_23239,N_23076,N_23047);
xnor U23240 (N_23240,N_23174,N_23079);
or U23241 (N_23241,N_23179,N_23099);
and U23242 (N_23242,N_23166,N_23013);
xnor U23243 (N_23243,N_23107,N_23141);
or U23244 (N_23244,N_23191,N_23043);
nor U23245 (N_23245,N_23188,N_23058);
or U23246 (N_23246,N_23006,N_23036);
nor U23247 (N_23247,N_23170,N_23014);
and U23248 (N_23248,N_23118,N_23042);
nand U23249 (N_23249,N_23094,N_23027);
nor U23250 (N_23250,N_23106,N_23165);
or U23251 (N_23251,N_23080,N_23098);
or U23252 (N_23252,N_23146,N_23049);
xor U23253 (N_23253,N_23182,N_23149);
and U23254 (N_23254,N_23002,N_23142);
and U23255 (N_23255,N_23184,N_23063);
and U23256 (N_23256,N_23032,N_23159);
and U23257 (N_23257,N_23119,N_23150);
nand U23258 (N_23258,N_23081,N_23087);
or U23259 (N_23259,N_23194,N_23176);
nand U23260 (N_23260,N_23148,N_23023);
xor U23261 (N_23261,N_23117,N_23126);
and U23262 (N_23262,N_23181,N_23055);
or U23263 (N_23263,N_23173,N_23162);
or U23264 (N_23264,N_23075,N_23160);
xor U23265 (N_23265,N_23048,N_23196);
nand U23266 (N_23266,N_23009,N_23156);
nand U23267 (N_23267,N_23001,N_23155);
nor U23268 (N_23268,N_23110,N_23021);
or U23269 (N_23269,N_23163,N_23175);
nor U23270 (N_23270,N_23114,N_23140);
nand U23271 (N_23271,N_23083,N_23074);
and U23272 (N_23272,N_23015,N_23108);
and U23273 (N_23273,N_23172,N_23111);
xnor U23274 (N_23274,N_23073,N_23143);
xnor U23275 (N_23275,N_23051,N_23003);
or U23276 (N_23276,N_23135,N_23187);
nand U23277 (N_23277,N_23101,N_23137);
nor U23278 (N_23278,N_23130,N_23072);
nor U23279 (N_23279,N_23029,N_23129);
nand U23280 (N_23280,N_23008,N_23035);
and U23281 (N_23281,N_23020,N_23037);
xnor U23282 (N_23282,N_23161,N_23061);
xor U23283 (N_23283,N_23092,N_23198);
and U23284 (N_23284,N_23177,N_23044);
nor U23285 (N_23285,N_23039,N_23031);
nand U23286 (N_23286,N_23004,N_23144);
and U23287 (N_23287,N_23097,N_23038);
nand U23288 (N_23288,N_23086,N_23122);
nand U23289 (N_23289,N_23033,N_23102);
nor U23290 (N_23290,N_23112,N_23012);
xnor U23291 (N_23291,N_23152,N_23186);
xor U23292 (N_23292,N_23059,N_23104);
or U23293 (N_23293,N_23069,N_23197);
nor U23294 (N_23294,N_23007,N_23185);
nor U23295 (N_23295,N_23105,N_23125);
nand U23296 (N_23296,N_23096,N_23138);
and U23297 (N_23297,N_23084,N_23067);
nand U23298 (N_23298,N_23183,N_23065);
nand U23299 (N_23299,N_23070,N_23053);
and U23300 (N_23300,N_23104,N_23134);
nand U23301 (N_23301,N_23070,N_23107);
nand U23302 (N_23302,N_23100,N_23115);
nand U23303 (N_23303,N_23084,N_23080);
xor U23304 (N_23304,N_23170,N_23033);
xor U23305 (N_23305,N_23080,N_23179);
nor U23306 (N_23306,N_23023,N_23187);
and U23307 (N_23307,N_23110,N_23083);
and U23308 (N_23308,N_23010,N_23024);
xor U23309 (N_23309,N_23171,N_23046);
or U23310 (N_23310,N_23083,N_23054);
xnor U23311 (N_23311,N_23119,N_23192);
or U23312 (N_23312,N_23001,N_23088);
or U23313 (N_23313,N_23185,N_23010);
and U23314 (N_23314,N_23186,N_23154);
xnor U23315 (N_23315,N_23162,N_23123);
and U23316 (N_23316,N_23099,N_23037);
nor U23317 (N_23317,N_23007,N_23113);
nand U23318 (N_23318,N_23054,N_23069);
nand U23319 (N_23319,N_23063,N_23071);
or U23320 (N_23320,N_23176,N_23091);
xnor U23321 (N_23321,N_23196,N_23154);
xnor U23322 (N_23322,N_23072,N_23096);
or U23323 (N_23323,N_23171,N_23125);
nor U23324 (N_23324,N_23016,N_23114);
nor U23325 (N_23325,N_23092,N_23075);
and U23326 (N_23326,N_23186,N_23189);
nor U23327 (N_23327,N_23110,N_23159);
and U23328 (N_23328,N_23061,N_23119);
nor U23329 (N_23329,N_23184,N_23073);
and U23330 (N_23330,N_23043,N_23021);
and U23331 (N_23331,N_23147,N_23188);
or U23332 (N_23332,N_23163,N_23021);
xnor U23333 (N_23333,N_23149,N_23045);
nand U23334 (N_23334,N_23110,N_23148);
and U23335 (N_23335,N_23138,N_23146);
and U23336 (N_23336,N_23153,N_23004);
nor U23337 (N_23337,N_23175,N_23154);
xnor U23338 (N_23338,N_23075,N_23117);
xor U23339 (N_23339,N_23119,N_23111);
or U23340 (N_23340,N_23150,N_23088);
or U23341 (N_23341,N_23133,N_23058);
or U23342 (N_23342,N_23014,N_23057);
nand U23343 (N_23343,N_23121,N_23160);
and U23344 (N_23344,N_23171,N_23038);
nor U23345 (N_23345,N_23179,N_23041);
nand U23346 (N_23346,N_23007,N_23155);
xnor U23347 (N_23347,N_23140,N_23046);
or U23348 (N_23348,N_23179,N_23004);
nand U23349 (N_23349,N_23072,N_23198);
nor U23350 (N_23350,N_23180,N_23133);
nand U23351 (N_23351,N_23100,N_23135);
and U23352 (N_23352,N_23059,N_23122);
and U23353 (N_23353,N_23136,N_23032);
nand U23354 (N_23354,N_23006,N_23190);
and U23355 (N_23355,N_23194,N_23027);
nor U23356 (N_23356,N_23003,N_23045);
and U23357 (N_23357,N_23060,N_23091);
nor U23358 (N_23358,N_23034,N_23144);
nor U23359 (N_23359,N_23164,N_23020);
nand U23360 (N_23360,N_23020,N_23161);
xnor U23361 (N_23361,N_23094,N_23117);
nor U23362 (N_23362,N_23190,N_23134);
nand U23363 (N_23363,N_23173,N_23097);
nand U23364 (N_23364,N_23098,N_23031);
or U23365 (N_23365,N_23076,N_23107);
and U23366 (N_23366,N_23040,N_23137);
nand U23367 (N_23367,N_23135,N_23040);
nor U23368 (N_23368,N_23066,N_23139);
nor U23369 (N_23369,N_23191,N_23146);
and U23370 (N_23370,N_23101,N_23019);
xnor U23371 (N_23371,N_23117,N_23149);
or U23372 (N_23372,N_23188,N_23014);
or U23373 (N_23373,N_23010,N_23002);
nand U23374 (N_23374,N_23075,N_23175);
nand U23375 (N_23375,N_23099,N_23131);
xor U23376 (N_23376,N_23191,N_23176);
and U23377 (N_23377,N_23198,N_23104);
nand U23378 (N_23378,N_23043,N_23196);
xor U23379 (N_23379,N_23120,N_23151);
and U23380 (N_23380,N_23195,N_23090);
or U23381 (N_23381,N_23032,N_23066);
and U23382 (N_23382,N_23180,N_23000);
or U23383 (N_23383,N_23184,N_23196);
or U23384 (N_23384,N_23179,N_23194);
nand U23385 (N_23385,N_23151,N_23137);
and U23386 (N_23386,N_23099,N_23159);
nor U23387 (N_23387,N_23060,N_23082);
and U23388 (N_23388,N_23076,N_23068);
nor U23389 (N_23389,N_23080,N_23030);
and U23390 (N_23390,N_23025,N_23062);
nand U23391 (N_23391,N_23153,N_23076);
and U23392 (N_23392,N_23170,N_23066);
and U23393 (N_23393,N_23043,N_23136);
nor U23394 (N_23394,N_23199,N_23115);
nor U23395 (N_23395,N_23052,N_23101);
xnor U23396 (N_23396,N_23026,N_23043);
and U23397 (N_23397,N_23199,N_23012);
xnor U23398 (N_23398,N_23198,N_23006);
or U23399 (N_23399,N_23134,N_23181);
and U23400 (N_23400,N_23392,N_23380);
or U23401 (N_23401,N_23345,N_23348);
nand U23402 (N_23402,N_23281,N_23275);
and U23403 (N_23403,N_23235,N_23201);
and U23404 (N_23404,N_23266,N_23312);
and U23405 (N_23405,N_23313,N_23215);
or U23406 (N_23406,N_23340,N_23357);
nand U23407 (N_23407,N_23242,N_23267);
nand U23408 (N_23408,N_23369,N_23301);
nand U23409 (N_23409,N_23280,N_23323);
nand U23410 (N_23410,N_23311,N_23206);
nor U23411 (N_23411,N_23330,N_23337);
nor U23412 (N_23412,N_23287,N_23295);
xor U23413 (N_23413,N_23274,N_23226);
nand U23414 (N_23414,N_23302,N_23253);
nor U23415 (N_23415,N_23254,N_23293);
xnor U23416 (N_23416,N_23391,N_23359);
nand U23417 (N_23417,N_23217,N_23343);
nor U23418 (N_23418,N_23204,N_23265);
nor U23419 (N_23419,N_23374,N_23365);
or U23420 (N_23420,N_23214,N_23223);
xnor U23421 (N_23421,N_23202,N_23211);
or U23422 (N_23422,N_23233,N_23219);
xnor U23423 (N_23423,N_23349,N_23237);
and U23424 (N_23424,N_23218,N_23394);
nor U23425 (N_23425,N_23360,N_23248);
and U23426 (N_23426,N_23342,N_23314);
and U23427 (N_23427,N_23309,N_23396);
and U23428 (N_23428,N_23339,N_23341);
xor U23429 (N_23429,N_23320,N_23382);
nor U23430 (N_23430,N_23353,N_23220);
nand U23431 (N_23431,N_23258,N_23335);
or U23432 (N_23432,N_23378,N_23385);
xor U23433 (N_23433,N_23326,N_23250);
nand U23434 (N_23434,N_23289,N_23328);
or U23435 (N_23435,N_23227,N_23307);
nand U23436 (N_23436,N_23279,N_23208);
nand U23437 (N_23437,N_23388,N_23234);
xor U23438 (N_23438,N_23346,N_23315);
or U23439 (N_23439,N_23232,N_23256);
and U23440 (N_23440,N_23306,N_23207);
nand U23441 (N_23441,N_23246,N_23243);
nor U23442 (N_23442,N_23318,N_23263);
nor U23443 (N_23443,N_23379,N_23308);
nor U23444 (N_23444,N_23347,N_23356);
and U23445 (N_23445,N_23277,N_23244);
or U23446 (N_23446,N_23299,N_23284);
and U23447 (N_23447,N_23310,N_23354);
and U23448 (N_23448,N_23322,N_23352);
nand U23449 (N_23449,N_23331,N_23222);
nand U23450 (N_23450,N_23260,N_23225);
nor U23451 (N_23451,N_23384,N_23325);
xnor U23452 (N_23452,N_23259,N_23247);
nand U23453 (N_23453,N_23355,N_23375);
xnor U23454 (N_23454,N_23350,N_23203);
xnor U23455 (N_23455,N_23252,N_23303);
nand U23456 (N_23456,N_23205,N_23283);
or U23457 (N_23457,N_23268,N_23371);
nand U23458 (N_23458,N_23316,N_23372);
nand U23459 (N_23459,N_23228,N_23393);
nor U23460 (N_23460,N_23200,N_23292);
or U23461 (N_23461,N_23264,N_23398);
nor U23462 (N_23462,N_23294,N_23332);
or U23463 (N_23463,N_23304,N_23209);
xnor U23464 (N_23464,N_23240,N_23224);
or U23465 (N_23465,N_23389,N_23255);
or U23466 (N_23466,N_23364,N_23291);
xor U23467 (N_23467,N_23238,N_23297);
nand U23468 (N_23468,N_23390,N_23361);
nor U23469 (N_23469,N_23338,N_23399);
xnor U23470 (N_23470,N_23285,N_23261);
xor U23471 (N_23471,N_23397,N_23271);
nand U23472 (N_23472,N_23270,N_23288);
nor U23473 (N_23473,N_23377,N_23239);
and U23474 (N_23474,N_23300,N_23276);
nand U23475 (N_23475,N_23298,N_23216);
nand U23476 (N_23476,N_23351,N_23231);
or U23477 (N_23477,N_23273,N_23386);
or U23478 (N_23478,N_23278,N_23395);
nand U23479 (N_23479,N_23262,N_23329);
xnor U23480 (N_23480,N_23290,N_23333);
nand U23481 (N_23481,N_23272,N_23305);
or U23482 (N_23482,N_23221,N_23387);
nor U23483 (N_23483,N_23286,N_23296);
nor U23484 (N_23484,N_23282,N_23327);
xor U23485 (N_23485,N_23251,N_23383);
and U23486 (N_23486,N_23213,N_23269);
and U23487 (N_23487,N_23358,N_23373);
or U23488 (N_23488,N_23376,N_23367);
nand U23489 (N_23489,N_23230,N_23257);
nor U23490 (N_23490,N_23368,N_23241);
or U23491 (N_23491,N_23334,N_23321);
nand U23492 (N_23492,N_23336,N_23317);
nand U23493 (N_23493,N_23249,N_23366);
and U23494 (N_23494,N_23381,N_23324);
and U23495 (N_23495,N_23210,N_23212);
and U23496 (N_23496,N_23319,N_23344);
and U23497 (N_23497,N_23362,N_23229);
nor U23498 (N_23498,N_23236,N_23363);
nand U23499 (N_23499,N_23370,N_23245);
xor U23500 (N_23500,N_23377,N_23337);
nand U23501 (N_23501,N_23238,N_23270);
xnor U23502 (N_23502,N_23221,N_23333);
xor U23503 (N_23503,N_23378,N_23318);
and U23504 (N_23504,N_23374,N_23249);
nand U23505 (N_23505,N_23271,N_23368);
or U23506 (N_23506,N_23283,N_23317);
or U23507 (N_23507,N_23235,N_23374);
nor U23508 (N_23508,N_23260,N_23397);
or U23509 (N_23509,N_23273,N_23216);
xnor U23510 (N_23510,N_23256,N_23286);
and U23511 (N_23511,N_23302,N_23343);
and U23512 (N_23512,N_23363,N_23280);
xnor U23513 (N_23513,N_23377,N_23318);
or U23514 (N_23514,N_23244,N_23290);
or U23515 (N_23515,N_23313,N_23300);
or U23516 (N_23516,N_23237,N_23257);
xor U23517 (N_23517,N_23229,N_23256);
nor U23518 (N_23518,N_23229,N_23344);
nor U23519 (N_23519,N_23383,N_23256);
or U23520 (N_23520,N_23378,N_23274);
nor U23521 (N_23521,N_23305,N_23209);
nand U23522 (N_23522,N_23365,N_23309);
or U23523 (N_23523,N_23337,N_23220);
and U23524 (N_23524,N_23347,N_23274);
nor U23525 (N_23525,N_23396,N_23231);
or U23526 (N_23526,N_23359,N_23345);
xnor U23527 (N_23527,N_23303,N_23391);
nand U23528 (N_23528,N_23260,N_23258);
or U23529 (N_23529,N_23385,N_23260);
nand U23530 (N_23530,N_23328,N_23373);
or U23531 (N_23531,N_23233,N_23260);
and U23532 (N_23532,N_23268,N_23385);
nand U23533 (N_23533,N_23366,N_23388);
nor U23534 (N_23534,N_23357,N_23238);
xnor U23535 (N_23535,N_23303,N_23315);
and U23536 (N_23536,N_23240,N_23370);
nor U23537 (N_23537,N_23215,N_23246);
or U23538 (N_23538,N_23309,N_23246);
or U23539 (N_23539,N_23353,N_23284);
and U23540 (N_23540,N_23272,N_23283);
nor U23541 (N_23541,N_23267,N_23326);
xor U23542 (N_23542,N_23266,N_23349);
nor U23543 (N_23543,N_23363,N_23353);
nor U23544 (N_23544,N_23279,N_23206);
and U23545 (N_23545,N_23205,N_23314);
or U23546 (N_23546,N_23200,N_23257);
xor U23547 (N_23547,N_23228,N_23235);
or U23548 (N_23548,N_23352,N_23237);
and U23549 (N_23549,N_23256,N_23385);
nor U23550 (N_23550,N_23308,N_23369);
xnor U23551 (N_23551,N_23274,N_23348);
nand U23552 (N_23552,N_23256,N_23394);
xor U23553 (N_23553,N_23221,N_23286);
xnor U23554 (N_23554,N_23371,N_23219);
xor U23555 (N_23555,N_23351,N_23306);
nand U23556 (N_23556,N_23232,N_23227);
xnor U23557 (N_23557,N_23337,N_23282);
nor U23558 (N_23558,N_23315,N_23327);
or U23559 (N_23559,N_23306,N_23388);
xnor U23560 (N_23560,N_23354,N_23238);
nand U23561 (N_23561,N_23283,N_23214);
nand U23562 (N_23562,N_23399,N_23361);
or U23563 (N_23563,N_23347,N_23395);
xor U23564 (N_23564,N_23314,N_23316);
or U23565 (N_23565,N_23331,N_23323);
nor U23566 (N_23566,N_23387,N_23378);
xnor U23567 (N_23567,N_23384,N_23299);
nor U23568 (N_23568,N_23368,N_23200);
nand U23569 (N_23569,N_23301,N_23222);
nand U23570 (N_23570,N_23340,N_23295);
xor U23571 (N_23571,N_23215,N_23276);
nor U23572 (N_23572,N_23227,N_23369);
and U23573 (N_23573,N_23311,N_23241);
nor U23574 (N_23574,N_23394,N_23334);
and U23575 (N_23575,N_23291,N_23251);
and U23576 (N_23576,N_23273,N_23335);
nor U23577 (N_23577,N_23382,N_23279);
nand U23578 (N_23578,N_23303,N_23291);
or U23579 (N_23579,N_23274,N_23382);
nor U23580 (N_23580,N_23292,N_23353);
nor U23581 (N_23581,N_23248,N_23290);
nand U23582 (N_23582,N_23232,N_23397);
nor U23583 (N_23583,N_23389,N_23227);
and U23584 (N_23584,N_23344,N_23256);
or U23585 (N_23585,N_23306,N_23383);
and U23586 (N_23586,N_23245,N_23250);
nor U23587 (N_23587,N_23295,N_23257);
nand U23588 (N_23588,N_23204,N_23296);
xnor U23589 (N_23589,N_23369,N_23399);
nor U23590 (N_23590,N_23349,N_23300);
or U23591 (N_23591,N_23241,N_23261);
or U23592 (N_23592,N_23382,N_23216);
xor U23593 (N_23593,N_23343,N_23214);
or U23594 (N_23594,N_23305,N_23396);
or U23595 (N_23595,N_23378,N_23321);
nor U23596 (N_23596,N_23341,N_23365);
xnor U23597 (N_23597,N_23358,N_23377);
nand U23598 (N_23598,N_23242,N_23202);
nor U23599 (N_23599,N_23374,N_23223);
and U23600 (N_23600,N_23545,N_23540);
nand U23601 (N_23601,N_23584,N_23533);
xnor U23602 (N_23602,N_23417,N_23517);
or U23603 (N_23603,N_23420,N_23456);
nand U23604 (N_23604,N_23442,N_23573);
nor U23605 (N_23605,N_23495,N_23422);
nand U23606 (N_23606,N_23571,N_23421);
and U23607 (N_23607,N_23447,N_23550);
nand U23608 (N_23608,N_23561,N_23441);
xor U23609 (N_23609,N_23565,N_23470);
nand U23610 (N_23610,N_23435,N_23488);
nand U23611 (N_23611,N_23536,N_23553);
or U23612 (N_23612,N_23539,N_23411);
nor U23613 (N_23613,N_23446,N_23471);
or U23614 (N_23614,N_23597,N_23588);
and U23615 (N_23615,N_23487,N_23590);
xnor U23616 (N_23616,N_23444,N_23412);
xor U23617 (N_23617,N_23506,N_23521);
nor U23618 (N_23618,N_23496,N_23579);
and U23619 (N_23619,N_23497,N_23523);
nor U23620 (N_23620,N_23459,N_23439);
and U23621 (N_23621,N_23402,N_23480);
and U23622 (N_23622,N_23543,N_23406);
or U23623 (N_23623,N_23587,N_23564);
and U23624 (N_23624,N_23580,N_23449);
or U23625 (N_23625,N_23460,N_23410);
and U23626 (N_23626,N_23489,N_23518);
nand U23627 (N_23627,N_23532,N_23559);
and U23628 (N_23628,N_23551,N_23527);
xnor U23629 (N_23629,N_23596,N_23453);
or U23630 (N_23630,N_23594,N_23486);
or U23631 (N_23631,N_23455,N_23424);
nand U23632 (N_23632,N_23448,N_23567);
nor U23633 (N_23633,N_23552,N_23415);
or U23634 (N_23634,N_23458,N_23546);
and U23635 (N_23635,N_23462,N_23469);
nand U23636 (N_23636,N_23510,N_23520);
nor U23637 (N_23637,N_23478,N_23586);
and U23638 (N_23638,N_23405,N_23475);
xnor U23639 (N_23639,N_23416,N_23537);
nor U23640 (N_23640,N_23400,N_23513);
nor U23641 (N_23641,N_23507,N_23515);
nand U23642 (N_23642,N_23593,N_23472);
and U23643 (N_23643,N_23583,N_23509);
or U23644 (N_23644,N_23554,N_23581);
xor U23645 (N_23645,N_23479,N_23434);
xor U23646 (N_23646,N_23544,N_23485);
nand U23647 (N_23647,N_23503,N_23560);
nand U23648 (N_23648,N_23563,N_23500);
nor U23649 (N_23649,N_23473,N_23401);
nor U23650 (N_23650,N_23505,N_23438);
nor U23651 (N_23651,N_23477,N_23522);
nand U23652 (N_23652,N_23430,N_23548);
xor U23653 (N_23653,N_23493,N_23433);
or U23654 (N_23654,N_23514,N_23598);
and U23655 (N_23655,N_23428,N_23404);
xor U23656 (N_23656,N_23499,N_23512);
xor U23657 (N_23657,N_23490,N_23465);
or U23658 (N_23658,N_23538,N_23595);
nand U23659 (N_23659,N_23549,N_23504);
xnor U23660 (N_23660,N_23556,N_23589);
nor U23661 (N_23661,N_23403,N_23576);
or U23662 (N_23662,N_23592,N_23562);
nor U23663 (N_23663,N_23467,N_23585);
xnor U23664 (N_23664,N_23418,N_23491);
xor U23665 (N_23665,N_23572,N_23461);
xor U23666 (N_23666,N_23457,N_23531);
nand U23667 (N_23667,N_23419,N_23492);
nand U23668 (N_23668,N_23429,N_23569);
xnor U23669 (N_23669,N_23519,N_23466);
or U23670 (N_23670,N_23451,N_23534);
and U23671 (N_23671,N_23599,N_23436);
and U23672 (N_23672,N_23528,N_23570);
nor U23673 (N_23673,N_23566,N_23407);
or U23674 (N_23674,N_23425,N_23511);
xnor U23675 (N_23675,N_23535,N_23577);
xor U23676 (N_23676,N_23431,N_23452);
xnor U23677 (N_23677,N_23474,N_23468);
nand U23678 (N_23678,N_23574,N_23575);
and U23679 (N_23679,N_23423,N_23501);
nand U23680 (N_23680,N_23427,N_23454);
or U23681 (N_23681,N_23445,N_23502);
nand U23682 (N_23682,N_23525,N_23526);
nand U23683 (N_23683,N_23558,N_23413);
nor U23684 (N_23684,N_23481,N_23437);
nor U23685 (N_23685,N_23529,N_23591);
nor U23686 (N_23686,N_23555,N_23450);
and U23687 (N_23687,N_23508,N_23568);
and U23688 (N_23688,N_23483,N_23414);
nand U23689 (N_23689,N_23408,N_23482);
xnor U23690 (N_23690,N_23494,N_23541);
or U23691 (N_23691,N_23498,N_23516);
or U23692 (N_23692,N_23409,N_23578);
or U23693 (N_23693,N_23530,N_23426);
nor U23694 (N_23694,N_23476,N_23440);
nor U23695 (N_23695,N_23464,N_23443);
nor U23696 (N_23696,N_23542,N_23484);
or U23697 (N_23697,N_23582,N_23557);
or U23698 (N_23698,N_23463,N_23432);
and U23699 (N_23699,N_23547,N_23524);
and U23700 (N_23700,N_23557,N_23453);
nand U23701 (N_23701,N_23452,N_23551);
xor U23702 (N_23702,N_23495,N_23522);
or U23703 (N_23703,N_23405,N_23453);
or U23704 (N_23704,N_23404,N_23570);
nand U23705 (N_23705,N_23423,N_23529);
xor U23706 (N_23706,N_23528,N_23535);
xor U23707 (N_23707,N_23437,N_23515);
nor U23708 (N_23708,N_23527,N_23455);
nand U23709 (N_23709,N_23579,N_23535);
nor U23710 (N_23710,N_23557,N_23559);
xnor U23711 (N_23711,N_23568,N_23551);
nand U23712 (N_23712,N_23493,N_23595);
nand U23713 (N_23713,N_23451,N_23597);
nor U23714 (N_23714,N_23573,N_23500);
or U23715 (N_23715,N_23490,N_23498);
xnor U23716 (N_23716,N_23517,N_23565);
nand U23717 (N_23717,N_23410,N_23581);
and U23718 (N_23718,N_23404,N_23490);
nand U23719 (N_23719,N_23427,N_23425);
and U23720 (N_23720,N_23525,N_23576);
or U23721 (N_23721,N_23428,N_23407);
and U23722 (N_23722,N_23517,N_23519);
nor U23723 (N_23723,N_23487,N_23489);
nor U23724 (N_23724,N_23522,N_23530);
xor U23725 (N_23725,N_23447,N_23505);
nand U23726 (N_23726,N_23424,N_23573);
xnor U23727 (N_23727,N_23447,N_23435);
xnor U23728 (N_23728,N_23576,N_23532);
and U23729 (N_23729,N_23592,N_23417);
or U23730 (N_23730,N_23482,N_23493);
nor U23731 (N_23731,N_23545,N_23560);
and U23732 (N_23732,N_23531,N_23555);
nand U23733 (N_23733,N_23555,N_23472);
or U23734 (N_23734,N_23503,N_23592);
nand U23735 (N_23735,N_23498,N_23545);
nor U23736 (N_23736,N_23564,N_23421);
nand U23737 (N_23737,N_23422,N_23559);
or U23738 (N_23738,N_23533,N_23477);
nor U23739 (N_23739,N_23417,N_23551);
nand U23740 (N_23740,N_23426,N_23433);
xnor U23741 (N_23741,N_23586,N_23479);
xnor U23742 (N_23742,N_23440,N_23579);
nand U23743 (N_23743,N_23532,N_23404);
nand U23744 (N_23744,N_23575,N_23587);
xnor U23745 (N_23745,N_23481,N_23483);
nand U23746 (N_23746,N_23564,N_23525);
xor U23747 (N_23747,N_23505,N_23513);
nand U23748 (N_23748,N_23598,N_23577);
and U23749 (N_23749,N_23434,N_23417);
nor U23750 (N_23750,N_23514,N_23543);
nand U23751 (N_23751,N_23411,N_23504);
xor U23752 (N_23752,N_23558,N_23447);
nand U23753 (N_23753,N_23465,N_23561);
xnor U23754 (N_23754,N_23493,N_23598);
xor U23755 (N_23755,N_23563,N_23514);
or U23756 (N_23756,N_23507,N_23445);
nor U23757 (N_23757,N_23411,N_23440);
or U23758 (N_23758,N_23584,N_23568);
nor U23759 (N_23759,N_23562,N_23579);
or U23760 (N_23760,N_23525,N_23567);
nand U23761 (N_23761,N_23511,N_23568);
nor U23762 (N_23762,N_23445,N_23498);
and U23763 (N_23763,N_23430,N_23493);
xor U23764 (N_23764,N_23447,N_23598);
nand U23765 (N_23765,N_23434,N_23408);
nor U23766 (N_23766,N_23429,N_23512);
xnor U23767 (N_23767,N_23494,N_23472);
or U23768 (N_23768,N_23535,N_23561);
nor U23769 (N_23769,N_23421,N_23462);
nor U23770 (N_23770,N_23542,N_23407);
and U23771 (N_23771,N_23516,N_23402);
nand U23772 (N_23772,N_23510,N_23530);
nor U23773 (N_23773,N_23582,N_23570);
and U23774 (N_23774,N_23415,N_23478);
and U23775 (N_23775,N_23598,N_23452);
and U23776 (N_23776,N_23477,N_23572);
nor U23777 (N_23777,N_23479,N_23467);
nor U23778 (N_23778,N_23426,N_23407);
xor U23779 (N_23779,N_23544,N_23486);
and U23780 (N_23780,N_23449,N_23510);
xor U23781 (N_23781,N_23461,N_23542);
nand U23782 (N_23782,N_23478,N_23449);
or U23783 (N_23783,N_23558,N_23535);
and U23784 (N_23784,N_23596,N_23550);
nor U23785 (N_23785,N_23519,N_23530);
or U23786 (N_23786,N_23573,N_23493);
nor U23787 (N_23787,N_23502,N_23536);
or U23788 (N_23788,N_23513,N_23436);
or U23789 (N_23789,N_23542,N_23488);
xnor U23790 (N_23790,N_23583,N_23441);
nand U23791 (N_23791,N_23469,N_23415);
nand U23792 (N_23792,N_23589,N_23457);
xnor U23793 (N_23793,N_23563,N_23562);
nand U23794 (N_23794,N_23446,N_23550);
or U23795 (N_23795,N_23551,N_23469);
and U23796 (N_23796,N_23458,N_23580);
and U23797 (N_23797,N_23524,N_23431);
and U23798 (N_23798,N_23597,N_23418);
nor U23799 (N_23799,N_23585,N_23486);
nor U23800 (N_23800,N_23738,N_23763);
nor U23801 (N_23801,N_23789,N_23795);
nand U23802 (N_23802,N_23764,N_23647);
nand U23803 (N_23803,N_23699,N_23707);
xnor U23804 (N_23804,N_23709,N_23770);
and U23805 (N_23805,N_23618,N_23611);
nor U23806 (N_23806,N_23643,N_23656);
and U23807 (N_23807,N_23775,N_23673);
and U23808 (N_23808,N_23634,N_23632);
xnor U23809 (N_23809,N_23749,N_23743);
and U23810 (N_23810,N_23605,N_23661);
nor U23811 (N_23811,N_23645,N_23724);
xnor U23812 (N_23812,N_23713,N_23607);
nor U23813 (N_23813,N_23682,N_23612);
or U23814 (N_23814,N_23793,N_23625);
and U23815 (N_23815,N_23760,N_23746);
and U23816 (N_23816,N_23765,N_23771);
and U23817 (N_23817,N_23790,N_23762);
or U23818 (N_23818,N_23675,N_23700);
xnor U23819 (N_23819,N_23608,N_23604);
nand U23820 (N_23820,N_23740,N_23722);
nor U23821 (N_23821,N_23719,N_23736);
or U23822 (N_23822,N_23687,N_23704);
or U23823 (N_23823,N_23767,N_23668);
xor U23824 (N_23824,N_23685,N_23626);
or U23825 (N_23825,N_23636,N_23664);
or U23826 (N_23826,N_23737,N_23655);
or U23827 (N_23827,N_23759,N_23774);
and U23828 (N_23828,N_23681,N_23657);
xor U23829 (N_23829,N_23646,N_23603);
nand U23830 (N_23830,N_23637,N_23624);
xor U23831 (N_23831,N_23686,N_23684);
nor U23832 (N_23832,N_23601,N_23698);
nor U23833 (N_23833,N_23797,N_23739);
or U23834 (N_23834,N_23695,N_23691);
xor U23835 (N_23835,N_23742,N_23725);
or U23836 (N_23836,N_23799,N_23796);
or U23837 (N_23837,N_23679,N_23777);
nor U23838 (N_23838,N_23750,N_23702);
nor U23839 (N_23839,N_23641,N_23747);
and U23840 (N_23840,N_23650,N_23613);
and U23841 (N_23841,N_23798,N_23610);
xnor U23842 (N_23842,N_23649,N_23781);
xor U23843 (N_23843,N_23720,N_23628);
xor U23844 (N_23844,N_23776,N_23670);
and U23845 (N_23845,N_23662,N_23680);
nand U23846 (N_23846,N_23640,N_23766);
xnor U23847 (N_23847,N_23727,N_23785);
nor U23848 (N_23848,N_23692,N_23642);
nor U23849 (N_23849,N_23674,N_23755);
and U23850 (N_23850,N_23619,N_23621);
and U23851 (N_23851,N_23653,N_23779);
or U23852 (N_23852,N_23783,N_23614);
xnor U23853 (N_23853,N_23768,N_23609);
xnor U23854 (N_23854,N_23630,N_23689);
xor U23855 (N_23855,N_23748,N_23701);
xor U23856 (N_23856,N_23658,N_23663);
or U23857 (N_23857,N_23620,N_23718);
or U23858 (N_23858,N_23703,N_23758);
and U23859 (N_23859,N_23633,N_23678);
and U23860 (N_23860,N_23710,N_23627);
nand U23861 (N_23861,N_23676,N_23752);
xor U23862 (N_23862,N_23677,N_23696);
xor U23863 (N_23863,N_23683,N_23600);
nand U23864 (N_23864,N_23723,N_23715);
and U23865 (N_23865,N_23741,N_23693);
xnor U23866 (N_23866,N_23669,N_23705);
or U23867 (N_23867,N_23734,N_23792);
nand U23868 (N_23868,N_23623,N_23780);
or U23869 (N_23869,N_23787,N_23757);
xnor U23870 (N_23870,N_23694,N_23730);
nor U23871 (N_23871,N_23617,N_23772);
nor U23872 (N_23872,N_23712,N_23615);
or U23873 (N_23873,N_23606,N_23754);
and U23874 (N_23874,N_23648,N_23671);
or U23875 (N_23875,N_23660,N_23753);
or U23876 (N_23876,N_23773,N_23667);
nor U23877 (N_23877,N_23728,N_23726);
and U23878 (N_23878,N_23659,N_23644);
nand U23879 (N_23879,N_23732,N_23631);
and U23880 (N_23880,N_23788,N_23716);
nor U23881 (N_23881,N_23652,N_23782);
and U23882 (N_23882,N_23666,N_23706);
nand U23883 (N_23883,N_23756,N_23616);
or U23884 (N_23884,N_23769,N_23761);
nor U23885 (N_23885,N_23665,N_23708);
nand U23886 (N_23886,N_23688,N_23744);
xnor U23887 (N_23887,N_23791,N_23711);
nand U23888 (N_23888,N_23651,N_23602);
nor U23889 (N_23889,N_23714,N_23635);
and U23890 (N_23890,N_23784,N_23622);
nor U23891 (N_23891,N_23639,N_23735);
nand U23892 (N_23892,N_23778,N_23672);
or U23893 (N_23893,N_23690,N_23717);
and U23894 (N_23894,N_23751,N_23729);
xor U23895 (N_23895,N_23721,N_23629);
or U23896 (N_23896,N_23731,N_23697);
nand U23897 (N_23897,N_23786,N_23733);
or U23898 (N_23898,N_23638,N_23745);
and U23899 (N_23899,N_23794,N_23654);
and U23900 (N_23900,N_23745,N_23677);
nor U23901 (N_23901,N_23629,N_23613);
nor U23902 (N_23902,N_23785,N_23612);
or U23903 (N_23903,N_23648,N_23652);
nor U23904 (N_23904,N_23703,N_23601);
xor U23905 (N_23905,N_23698,N_23775);
nor U23906 (N_23906,N_23748,N_23650);
nand U23907 (N_23907,N_23677,N_23632);
or U23908 (N_23908,N_23765,N_23613);
nand U23909 (N_23909,N_23768,N_23616);
nor U23910 (N_23910,N_23786,N_23747);
xnor U23911 (N_23911,N_23610,N_23686);
nor U23912 (N_23912,N_23674,N_23614);
nand U23913 (N_23913,N_23652,N_23788);
xnor U23914 (N_23914,N_23645,N_23638);
xnor U23915 (N_23915,N_23791,N_23630);
xor U23916 (N_23916,N_23639,N_23667);
nor U23917 (N_23917,N_23672,N_23745);
nor U23918 (N_23918,N_23689,N_23799);
nand U23919 (N_23919,N_23674,N_23633);
nand U23920 (N_23920,N_23616,N_23627);
nor U23921 (N_23921,N_23792,N_23701);
xnor U23922 (N_23922,N_23678,N_23729);
xor U23923 (N_23923,N_23628,N_23636);
or U23924 (N_23924,N_23713,N_23743);
nor U23925 (N_23925,N_23618,N_23665);
xor U23926 (N_23926,N_23726,N_23707);
nor U23927 (N_23927,N_23627,N_23614);
nor U23928 (N_23928,N_23662,N_23699);
nand U23929 (N_23929,N_23757,N_23769);
xnor U23930 (N_23930,N_23733,N_23756);
and U23931 (N_23931,N_23743,N_23770);
or U23932 (N_23932,N_23647,N_23605);
xor U23933 (N_23933,N_23733,N_23779);
and U23934 (N_23934,N_23701,N_23764);
and U23935 (N_23935,N_23630,N_23619);
xor U23936 (N_23936,N_23729,N_23713);
and U23937 (N_23937,N_23727,N_23758);
nor U23938 (N_23938,N_23600,N_23654);
nand U23939 (N_23939,N_23734,N_23672);
xnor U23940 (N_23940,N_23645,N_23683);
nor U23941 (N_23941,N_23764,N_23620);
nor U23942 (N_23942,N_23702,N_23637);
nand U23943 (N_23943,N_23611,N_23647);
and U23944 (N_23944,N_23636,N_23714);
nand U23945 (N_23945,N_23695,N_23784);
or U23946 (N_23946,N_23739,N_23716);
xor U23947 (N_23947,N_23730,N_23766);
and U23948 (N_23948,N_23695,N_23752);
xor U23949 (N_23949,N_23609,N_23625);
and U23950 (N_23950,N_23675,N_23610);
or U23951 (N_23951,N_23669,N_23657);
nand U23952 (N_23952,N_23691,N_23644);
xnor U23953 (N_23953,N_23636,N_23663);
xor U23954 (N_23954,N_23654,N_23685);
and U23955 (N_23955,N_23722,N_23679);
nand U23956 (N_23956,N_23741,N_23752);
or U23957 (N_23957,N_23747,N_23643);
and U23958 (N_23958,N_23771,N_23656);
xor U23959 (N_23959,N_23678,N_23619);
or U23960 (N_23960,N_23713,N_23700);
nand U23961 (N_23961,N_23772,N_23757);
xnor U23962 (N_23962,N_23745,N_23740);
xor U23963 (N_23963,N_23720,N_23635);
and U23964 (N_23964,N_23675,N_23737);
nor U23965 (N_23965,N_23690,N_23630);
and U23966 (N_23966,N_23679,N_23632);
and U23967 (N_23967,N_23746,N_23622);
or U23968 (N_23968,N_23776,N_23798);
or U23969 (N_23969,N_23673,N_23662);
or U23970 (N_23970,N_23797,N_23721);
and U23971 (N_23971,N_23728,N_23785);
xor U23972 (N_23972,N_23796,N_23700);
xnor U23973 (N_23973,N_23641,N_23738);
xor U23974 (N_23974,N_23689,N_23607);
and U23975 (N_23975,N_23604,N_23709);
and U23976 (N_23976,N_23693,N_23752);
nand U23977 (N_23977,N_23669,N_23662);
or U23978 (N_23978,N_23759,N_23698);
and U23979 (N_23979,N_23736,N_23724);
and U23980 (N_23980,N_23668,N_23677);
and U23981 (N_23981,N_23660,N_23655);
nor U23982 (N_23982,N_23768,N_23648);
xor U23983 (N_23983,N_23628,N_23760);
nor U23984 (N_23984,N_23758,N_23675);
and U23985 (N_23985,N_23630,N_23786);
nand U23986 (N_23986,N_23671,N_23709);
and U23987 (N_23987,N_23612,N_23775);
xor U23988 (N_23988,N_23667,N_23727);
nand U23989 (N_23989,N_23699,N_23757);
nand U23990 (N_23990,N_23639,N_23739);
nor U23991 (N_23991,N_23678,N_23622);
xnor U23992 (N_23992,N_23734,N_23707);
nand U23993 (N_23993,N_23655,N_23762);
xor U23994 (N_23994,N_23744,N_23649);
xor U23995 (N_23995,N_23625,N_23604);
xor U23996 (N_23996,N_23729,N_23620);
or U23997 (N_23997,N_23764,N_23692);
nor U23998 (N_23998,N_23655,N_23779);
and U23999 (N_23999,N_23709,N_23630);
nor U24000 (N_24000,N_23976,N_23863);
or U24001 (N_24001,N_23813,N_23963);
and U24002 (N_24002,N_23859,N_23905);
or U24003 (N_24003,N_23897,N_23808);
nor U24004 (N_24004,N_23869,N_23837);
nor U24005 (N_24005,N_23845,N_23986);
nor U24006 (N_24006,N_23952,N_23853);
and U24007 (N_24007,N_23882,N_23928);
and U24008 (N_24008,N_23877,N_23881);
and U24009 (N_24009,N_23925,N_23930);
nand U24010 (N_24010,N_23997,N_23918);
nand U24011 (N_24011,N_23831,N_23994);
nand U24012 (N_24012,N_23864,N_23811);
nor U24013 (N_24013,N_23923,N_23933);
nor U24014 (N_24014,N_23969,N_23849);
xor U24015 (N_24015,N_23974,N_23807);
or U24016 (N_24016,N_23938,N_23922);
xor U24017 (N_24017,N_23911,N_23862);
xor U24018 (N_24018,N_23815,N_23944);
nand U24019 (N_24019,N_23810,N_23868);
xor U24020 (N_24020,N_23895,N_23800);
xor U24021 (N_24021,N_23945,N_23814);
or U24022 (N_24022,N_23989,N_23840);
nand U24023 (N_24023,N_23872,N_23916);
or U24024 (N_24024,N_23919,N_23826);
or U24025 (N_24025,N_23917,N_23825);
or U24026 (N_24026,N_23817,N_23979);
nand U24027 (N_24027,N_23874,N_23820);
nand U24028 (N_24028,N_23954,N_23931);
or U24029 (N_24029,N_23883,N_23982);
nand U24030 (N_24030,N_23876,N_23962);
and U24031 (N_24031,N_23912,N_23947);
and U24032 (N_24032,N_23865,N_23847);
or U24033 (N_24033,N_23995,N_23898);
nand U24034 (N_24034,N_23926,N_23977);
nand U24035 (N_24035,N_23805,N_23848);
and U24036 (N_24036,N_23892,N_23818);
or U24037 (N_24037,N_23861,N_23824);
or U24038 (N_24038,N_23819,N_23880);
xnor U24039 (N_24039,N_23910,N_23854);
and U24040 (N_24040,N_23834,N_23968);
or U24041 (N_24041,N_23841,N_23955);
nand U24042 (N_24042,N_23970,N_23804);
and U24043 (N_24043,N_23878,N_23851);
xnor U24044 (N_24044,N_23959,N_23875);
or U24045 (N_24045,N_23913,N_23921);
or U24046 (N_24046,N_23915,N_23946);
and U24047 (N_24047,N_23833,N_23873);
nor U24048 (N_24048,N_23980,N_23832);
or U24049 (N_24049,N_23823,N_23920);
and U24050 (N_24050,N_23996,N_23924);
nor U24051 (N_24051,N_23953,N_23827);
and U24052 (N_24052,N_23907,N_23987);
nand U24053 (N_24053,N_23957,N_23900);
xnor U24054 (N_24054,N_23909,N_23879);
nand U24055 (N_24055,N_23850,N_23937);
nor U24056 (N_24056,N_23899,N_23902);
or U24057 (N_24057,N_23958,N_23842);
nor U24058 (N_24058,N_23855,N_23803);
or U24059 (N_24059,N_23992,N_23991);
nand U24060 (N_24060,N_23866,N_23960);
and U24061 (N_24061,N_23836,N_23839);
xnor U24062 (N_24062,N_23889,N_23941);
xnor U24063 (N_24063,N_23870,N_23886);
nor U24064 (N_24064,N_23844,N_23809);
nand U24065 (N_24065,N_23896,N_23943);
nand U24066 (N_24066,N_23829,N_23830);
or U24067 (N_24067,N_23998,N_23965);
xnor U24068 (N_24068,N_23988,N_23906);
xnor U24069 (N_24069,N_23893,N_23971);
or U24070 (N_24070,N_23949,N_23961);
nand U24071 (N_24071,N_23802,N_23951);
and U24072 (N_24072,N_23940,N_23908);
xnor U24073 (N_24073,N_23822,N_23846);
nor U24074 (N_24074,N_23934,N_23948);
xnor U24075 (N_24075,N_23975,N_23867);
and U24076 (N_24076,N_23891,N_23966);
xnor U24077 (N_24077,N_23828,N_23973);
or U24078 (N_24078,N_23821,N_23806);
and U24079 (N_24079,N_23981,N_23812);
nand U24080 (N_24080,N_23993,N_23972);
nand U24081 (N_24081,N_23999,N_23894);
xor U24082 (N_24082,N_23983,N_23942);
and U24083 (N_24083,N_23950,N_23857);
xor U24084 (N_24084,N_23936,N_23860);
and U24085 (N_24085,N_23932,N_23816);
nand U24086 (N_24086,N_23888,N_23885);
or U24087 (N_24087,N_23935,N_23856);
or U24088 (N_24088,N_23871,N_23985);
or U24089 (N_24089,N_23967,N_23978);
and U24090 (N_24090,N_23904,N_23927);
and U24091 (N_24091,N_23939,N_23903);
xor U24092 (N_24092,N_23858,N_23887);
and U24093 (N_24093,N_23801,N_23901);
or U24094 (N_24094,N_23852,N_23929);
nor U24095 (N_24095,N_23990,N_23890);
nand U24096 (N_24096,N_23835,N_23984);
nor U24097 (N_24097,N_23956,N_23914);
xnor U24098 (N_24098,N_23884,N_23964);
nor U24099 (N_24099,N_23838,N_23843);
nor U24100 (N_24100,N_23821,N_23818);
xnor U24101 (N_24101,N_23813,N_23920);
xnor U24102 (N_24102,N_23934,N_23940);
nand U24103 (N_24103,N_23942,N_23982);
or U24104 (N_24104,N_23936,N_23868);
nand U24105 (N_24105,N_23811,N_23940);
and U24106 (N_24106,N_23946,N_23981);
and U24107 (N_24107,N_23807,N_23860);
or U24108 (N_24108,N_23841,N_23965);
nand U24109 (N_24109,N_23909,N_23899);
nor U24110 (N_24110,N_23926,N_23891);
nor U24111 (N_24111,N_23906,N_23851);
nor U24112 (N_24112,N_23962,N_23945);
xnor U24113 (N_24113,N_23851,N_23823);
and U24114 (N_24114,N_23933,N_23994);
nor U24115 (N_24115,N_23801,N_23871);
xor U24116 (N_24116,N_23811,N_23881);
xnor U24117 (N_24117,N_23862,N_23893);
nand U24118 (N_24118,N_23840,N_23969);
or U24119 (N_24119,N_23986,N_23813);
nor U24120 (N_24120,N_23975,N_23958);
or U24121 (N_24121,N_23814,N_23992);
nor U24122 (N_24122,N_23824,N_23991);
nor U24123 (N_24123,N_23944,N_23977);
nor U24124 (N_24124,N_23868,N_23820);
xor U24125 (N_24125,N_23842,N_23848);
and U24126 (N_24126,N_23846,N_23934);
nand U24127 (N_24127,N_23846,N_23907);
nand U24128 (N_24128,N_23852,N_23987);
xnor U24129 (N_24129,N_23922,N_23947);
xnor U24130 (N_24130,N_23951,N_23817);
nor U24131 (N_24131,N_23993,N_23845);
xnor U24132 (N_24132,N_23827,N_23829);
or U24133 (N_24133,N_23928,N_23916);
and U24134 (N_24134,N_23980,N_23897);
nor U24135 (N_24135,N_23977,N_23892);
or U24136 (N_24136,N_23998,N_23891);
or U24137 (N_24137,N_23803,N_23883);
nor U24138 (N_24138,N_23826,N_23873);
nor U24139 (N_24139,N_23987,N_23847);
or U24140 (N_24140,N_23930,N_23921);
and U24141 (N_24141,N_23804,N_23831);
nor U24142 (N_24142,N_23913,N_23880);
xnor U24143 (N_24143,N_23964,N_23802);
nand U24144 (N_24144,N_23810,N_23945);
and U24145 (N_24145,N_23931,N_23966);
and U24146 (N_24146,N_23889,N_23998);
and U24147 (N_24147,N_23907,N_23857);
nor U24148 (N_24148,N_23837,N_23836);
and U24149 (N_24149,N_23934,N_23887);
nor U24150 (N_24150,N_23864,N_23851);
xnor U24151 (N_24151,N_23850,N_23991);
nand U24152 (N_24152,N_23973,N_23883);
xor U24153 (N_24153,N_23955,N_23819);
nor U24154 (N_24154,N_23964,N_23862);
xnor U24155 (N_24155,N_23916,N_23925);
nor U24156 (N_24156,N_23851,N_23976);
and U24157 (N_24157,N_23887,N_23873);
nor U24158 (N_24158,N_23993,N_23981);
nand U24159 (N_24159,N_23980,N_23855);
and U24160 (N_24160,N_23825,N_23800);
and U24161 (N_24161,N_23860,N_23981);
xor U24162 (N_24162,N_23994,N_23911);
nand U24163 (N_24163,N_23943,N_23884);
nand U24164 (N_24164,N_23949,N_23902);
nor U24165 (N_24165,N_23856,N_23994);
and U24166 (N_24166,N_23907,N_23940);
nand U24167 (N_24167,N_23808,N_23838);
or U24168 (N_24168,N_23961,N_23846);
nor U24169 (N_24169,N_23823,N_23815);
and U24170 (N_24170,N_23817,N_23989);
or U24171 (N_24171,N_23869,N_23986);
or U24172 (N_24172,N_23970,N_23928);
or U24173 (N_24173,N_23940,N_23817);
or U24174 (N_24174,N_23847,N_23871);
or U24175 (N_24175,N_23985,N_23942);
nand U24176 (N_24176,N_23912,N_23936);
or U24177 (N_24177,N_23876,N_23929);
or U24178 (N_24178,N_23875,N_23916);
nor U24179 (N_24179,N_23982,N_23823);
nand U24180 (N_24180,N_23849,N_23868);
and U24181 (N_24181,N_23926,N_23983);
nor U24182 (N_24182,N_23991,N_23861);
xnor U24183 (N_24183,N_23815,N_23824);
nand U24184 (N_24184,N_23889,N_23826);
or U24185 (N_24185,N_23885,N_23855);
nand U24186 (N_24186,N_23895,N_23841);
xor U24187 (N_24187,N_23923,N_23899);
nand U24188 (N_24188,N_23812,N_23832);
xor U24189 (N_24189,N_23963,N_23993);
nor U24190 (N_24190,N_23875,N_23828);
nand U24191 (N_24191,N_23900,N_23835);
nand U24192 (N_24192,N_23816,N_23993);
xor U24193 (N_24193,N_23891,N_23988);
nor U24194 (N_24194,N_23949,N_23950);
nand U24195 (N_24195,N_23965,N_23849);
nor U24196 (N_24196,N_23820,N_23850);
xor U24197 (N_24197,N_23857,N_23819);
and U24198 (N_24198,N_23844,N_23842);
or U24199 (N_24199,N_23851,N_23969);
and U24200 (N_24200,N_24078,N_24188);
or U24201 (N_24201,N_24156,N_24172);
nand U24202 (N_24202,N_24042,N_24117);
nand U24203 (N_24203,N_24154,N_24103);
xnor U24204 (N_24204,N_24069,N_24012);
xor U24205 (N_24205,N_24027,N_24127);
nor U24206 (N_24206,N_24085,N_24184);
nor U24207 (N_24207,N_24089,N_24060);
nor U24208 (N_24208,N_24026,N_24025);
or U24209 (N_24209,N_24185,N_24055);
and U24210 (N_24210,N_24120,N_24165);
and U24211 (N_24211,N_24155,N_24008);
xnor U24212 (N_24212,N_24023,N_24097);
or U24213 (N_24213,N_24082,N_24022);
xor U24214 (N_24214,N_24190,N_24086);
nand U24215 (N_24215,N_24095,N_24101);
or U24216 (N_24216,N_24088,N_24031);
xor U24217 (N_24217,N_24092,N_24125);
nand U24218 (N_24218,N_24017,N_24131);
or U24219 (N_24219,N_24080,N_24104);
nor U24220 (N_24220,N_24047,N_24011);
nor U24221 (N_24221,N_24014,N_24112);
nor U24222 (N_24222,N_24074,N_24149);
nand U24223 (N_24223,N_24106,N_24186);
xnor U24224 (N_24224,N_24062,N_24132);
nor U24225 (N_24225,N_24006,N_24063);
nand U24226 (N_24226,N_24122,N_24194);
xnor U24227 (N_24227,N_24076,N_24158);
xor U24228 (N_24228,N_24049,N_24070);
nand U24229 (N_24229,N_24140,N_24151);
nand U24230 (N_24230,N_24032,N_24135);
and U24231 (N_24231,N_24133,N_24065);
xor U24232 (N_24232,N_24142,N_24174);
or U24233 (N_24233,N_24056,N_24040);
or U24234 (N_24234,N_24182,N_24196);
and U24235 (N_24235,N_24020,N_24116);
xnor U24236 (N_24236,N_24183,N_24100);
xor U24237 (N_24237,N_24093,N_24028);
xor U24238 (N_24238,N_24067,N_24004);
xnor U24239 (N_24239,N_24169,N_24128);
xor U24240 (N_24240,N_24146,N_24139);
and U24241 (N_24241,N_24015,N_24197);
nand U24242 (N_24242,N_24123,N_24118);
xor U24243 (N_24243,N_24037,N_24124);
or U24244 (N_24244,N_24199,N_24046);
nand U24245 (N_24245,N_24108,N_24102);
nand U24246 (N_24246,N_24115,N_24129);
nor U24247 (N_24247,N_24144,N_24077);
or U24248 (N_24248,N_24059,N_24036);
and U24249 (N_24249,N_24162,N_24010);
or U24250 (N_24250,N_24180,N_24052);
or U24251 (N_24251,N_24167,N_24000);
or U24252 (N_24252,N_24091,N_24045);
nor U24253 (N_24253,N_24111,N_24003);
xor U24254 (N_24254,N_24176,N_24177);
and U24255 (N_24255,N_24007,N_24002);
nor U24256 (N_24256,N_24050,N_24179);
and U24257 (N_24257,N_24113,N_24141);
xor U24258 (N_24258,N_24198,N_24073);
xnor U24259 (N_24259,N_24134,N_24081);
nand U24260 (N_24260,N_24064,N_24096);
nor U24261 (N_24261,N_24119,N_24137);
nor U24262 (N_24262,N_24173,N_24138);
nor U24263 (N_24263,N_24066,N_24033);
and U24264 (N_24264,N_24009,N_24166);
nand U24265 (N_24265,N_24099,N_24018);
xor U24266 (N_24266,N_24013,N_24121);
nor U24267 (N_24267,N_24126,N_24171);
nor U24268 (N_24268,N_24163,N_24021);
and U24269 (N_24269,N_24043,N_24164);
and U24270 (N_24270,N_24160,N_24035);
or U24271 (N_24271,N_24039,N_24016);
nand U24272 (N_24272,N_24147,N_24072);
and U24273 (N_24273,N_24170,N_24130);
and U24274 (N_24274,N_24153,N_24187);
nor U24275 (N_24275,N_24053,N_24150);
and U24276 (N_24276,N_24054,N_24058);
and U24277 (N_24277,N_24109,N_24114);
and U24278 (N_24278,N_24079,N_24005);
and U24279 (N_24279,N_24191,N_24178);
and U24280 (N_24280,N_24068,N_24061);
or U24281 (N_24281,N_24105,N_24161);
xnor U24282 (N_24282,N_24024,N_24189);
or U24283 (N_24283,N_24098,N_24192);
and U24284 (N_24284,N_24168,N_24083);
xnor U24285 (N_24285,N_24152,N_24030);
xnor U24286 (N_24286,N_24181,N_24107);
and U24287 (N_24287,N_24057,N_24034);
nand U24288 (N_24288,N_24175,N_24195);
nor U24289 (N_24289,N_24136,N_24029);
xor U24290 (N_24290,N_24090,N_24048);
nand U24291 (N_24291,N_24087,N_24075);
nor U24292 (N_24292,N_24148,N_24193);
and U24293 (N_24293,N_24038,N_24019);
xnor U24294 (N_24294,N_24159,N_24094);
xnor U24295 (N_24295,N_24041,N_24110);
nand U24296 (N_24296,N_24143,N_24071);
nor U24297 (N_24297,N_24084,N_24145);
and U24298 (N_24298,N_24157,N_24051);
xor U24299 (N_24299,N_24044,N_24001);
nor U24300 (N_24300,N_24133,N_24115);
xor U24301 (N_24301,N_24017,N_24092);
and U24302 (N_24302,N_24012,N_24051);
nand U24303 (N_24303,N_24180,N_24089);
or U24304 (N_24304,N_24067,N_24084);
nand U24305 (N_24305,N_24010,N_24014);
xor U24306 (N_24306,N_24070,N_24033);
xnor U24307 (N_24307,N_24074,N_24052);
xor U24308 (N_24308,N_24008,N_24187);
xor U24309 (N_24309,N_24074,N_24153);
nor U24310 (N_24310,N_24172,N_24052);
or U24311 (N_24311,N_24123,N_24119);
nor U24312 (N_24312,N_24195,N_24143);
or U24313 (N_24313,N_24030,N_24137);
xnor U24314 (N_24314,N_24154,N_24191);
or U24315 (N_24315,N_24164,N_24133);
or U24316 (N_24316,N_24109,N_24027);
xnor U24317 (N_24317,N_24099,N_24066);
xor U24318 (N_24318,N_24168,N_24171);
xor U24319 (N_24319,N_24129,N_24081);
xnor U24320 (N_24320,N_24058,N_24194);
xor U24321 (N_24321,N_24062,N_24040);
and U24322 (N_24322,N_24108,N_24185);
nor U24323 (N_24323,N_24160,N_24127);
and U24324 (N_24324,N_24034,N_24061);
nand U24325 (N_24325,N_24169,N_24164);
nand U24326 (N_24326,N_24127,N_24120);
or U24327 (N_24327,N_24170,N_24142);
or U24328 (N_24328,N_24048,N_24111);
and U24329 (N_24329,N_24109,N_24010);
and U24330 (N_24330,N_24161,N_24001);
nand U24331 (N_24331,N_24164,N_24111);
or U24332 (N_24332,N_24034,N_24149);
nand U24333 (N_24333,N_24058,N_24076);
and U24334 (N_24334,N_24076,N_24108);
or U24335 (N_24335,N_24075,N_24077);
nor U24336 (N_24336,N_24198,N_24175);
nor U24337 (N_24337,N_24113,N_24001);
xor U24338 (N_24338,N_24039,N_24120);
xor U24339 (N_24339,N_24148,N_24146);
or U24340 (N_24340,N_24182,N_24014);
xor U24341 (N_24341,N_24128,N_24108);
nor U24342 (N_24342,N_24171,N_24102);
nor U24343 (N_24343,N_24090,N_24027);
nand U24344 (N_24344,N_24141,N_24022);
nand U24345 (N_24345,N_24131,N_24146);
nand U24346 (N_24346,N_24093,N_24163);
nor U24347 (N_24347,N_24102,N_24099);
nand U24348 (N_24348,N_24070,N_24039);
nand U24349 (N_24349,N_24073,N_24023);
and U24350 (N_24350,N_24124,N_24083);
nor U24351 (N_24351,N_24109,N_24169);
nor U24352 (N_24352,N_24078,N_24061);
and U24353 (N_24353,N_24175,N_24074);
and U24354 (N_24354,N_24193,N_24188);
or U24355 (N_24355,N_24044,N_24089);
nor U24356 (N_24356,N_24158,N_24108);
xnor U24357 (N_24357,N_24030,N_24043);
and U24358 (N_24358,N_24076,N_24049);
or U24359 (N_24359,N_24126,N_24119);
nor U24360 (N_24360,N_24193,N_24024);
or U24361 (N_24361,N_24021,N_24134);
nor U24362 (N_24362,N_24189,N_24013);
nand U24363 (N_24363,N_24063,N_24170);
nand U24364 (N_24364,N_24089,N_24163);
xor U24365 (N_24365,N_24053,N_24087);
nor U24366 (N_24366,N_24179,N_24144);
or U24367 (N_24367,N_24143,N_24107);
or U24368 (N_24368,N_24141,N_24158);
nand U24369 (N_24369,N_24033,N_24056);
nand U24370 (N_24370,N_24125,N_24027);
or U24371 (N_24371,N_24164,N_24126);
nand U24372 (N_24372,N_24075,N_24167);
xnor U24373 (N_24373,N_24084,N_24197);
nor U24374 (N_24374,N_24024,N_24025);
and U24375 (N_24375,N_24069,N_24140);
and U24376 (N_24376,N_24048,N_24056);
nand U24377 (N_24377,N_24184,N_24071);
or U24378 (N_24378,N_24145,N_24178);
nor U24379 (N_24379,N_24079,N_24053);
or U24380 (N_24380,N_24050,N_24164);
and U24381 (N_24381,N_24029,N_24048);
and U24382 (N_24382,N_24142,N_24178);
nor U24383 (N_24383,N_24103,N_24042);
nand U24384 (N_24384,N_24034,N_24009);
and U24385 (N_24385,N_24038,N_24189);
nor U24386 (N_24386,N_24103,N_24093);
or U24387 (N_24387,N_24098,N_24108);
xor U24388 (N_24388,N_24092,N_24103);
or U24389 (N_24389,N_24003,N_24015);
or U24390 (N_24390,N_24063,N_24135);
xor U24391 (N_24391,N_24185,N_24164);
nor U24392 (N_24392,N_24138,N_24188);
nor U24393 (N_24393,N_24174,N_24157);
or U24394 (N_24394,N_24177,N_24063);
nor U24395 (N_24395,N_24165,N_24020);
xor U24396 (N_24396,N_24190,N_24117);
xor U24397 (N_24397,N_24054,N_24073);
xor U24398 (N_24398,N_24132,N_24016);
nand U24399 (N_24399,N_24034,N_24160);
xor U24400 (N_24400,N_24369,N_24219);
or U24401 (N_24401,N_24233,N_24361);
nor U24402 (N_24402,N_24235,N_24265);
xor U24403 (N_24403,N_24266,N_24240);
nand U24404 (N_24404,N_24318,N_24322);
or U24405 (N_24405,N_24214,N_24356);
nand U24406 (N_24406,N_24383,N_24249);
and U24407 (N_24407,N_24232,N_24252);
nor U24408 (N_24408,N_24342,N_24347);
nand U24409 (N_24409,N_24320,N_24336);
xor U24410 (N_24410,N_24374,N_24377);
nor U24411 (N_24411,N_24255,N_24277);
nor U24412 (N_24412,N_24393,N_24331);
nand U24413 (N_24413,N_24359,N_24310);
xor U24414 (N_24414,N_24243,N_24236);
xnor U24415 (N_24415,N_24313,N_24220);
xor U24416 (N_24416,N_24395,N_24217);
or U24417 (N_24417,N_24341,N_24248);
and U24418 (N_24418,N_24373,N_24376);
nor U24419 (N_24419,N_24215,N_24258);
xnor U24420 (N_24420,N_24271,N_24203);
or U24421 (N_24421,N_24208,N_24365);
nor U24422 (N_24422,N_24293,N_24225);
or U24423 (N_24423,N_24283,N_24273);
and U24424 (N_24424,N_24216,N_24263);
nand U24425 (N_24425,N_24287,N_24382);
and U24426 (N_24426,N_24354,N_24357);
nand U24427 (N_24427,N_24380,N_24372);
nand U24428 (N_24428,N_24275,N_24344);
nor U24429 (N_24429,N_24352,N_24253);
xnor U24430 (N_24430,N_24334,N_24363);
xnor U24431 (N_24431,N_24319,N_24210);
xor U24432 (N_24432,N_24333,N_24229);
nor U24433 (N_24433,N_24228,N_24281);
or U24434 (N_24434,N_24224,N_24389);
and U24435 (N_24435,N_24387,N_24241);
xnor U24436 (N_24436,N_24360,N_24268);
xnor U24437 (N_24437,N_24370,N_24307);
nor U24438 (N_24438,N_24260,N_24378);
xor U24439 (N_24439,N_24392,N_24290);
or U24440 (N_24440,N_24270,N_24304);
and U24441 (N_24441,N_24353,N_24269);
or U24442 (N_24442,N_24244,N_24278);
and U24443 (N_24443,N_24371,N_24238);
nand U24444 (N_24444,N_24251,N_24259);
nor U24445 (N_24445,N_24204,N_24296);
nor U24446 (N_24446,N_24299,N_24300);
nand U24447 (N_24447,N_24398,N_24348);
xor U24448 (N_24448,N_24394,N_24321);
and U24449 (N_24449,N_24303,N_24256);
and U24450 (N_24450,N_24330,N_24335);
nor U24451 (N_24451,N_24221,N_24209);
or U24452 (N_24452,N_24326,N_24350);
or U24453 (N_24453,N_24292,N_24212);
and U24454 (N_24454,N_24323,N_24351);
and U24455 (N_24455,N_24272,N_24230);
xnor U24456 (N_24456,N_24366,N_24329);
xnor U24457 (N_24457,N_24284,N_24332);
xnor U24458 (N_24458,N_24355,N_24302);
nand U24459 (N_24459,N_24367,N_24205);
xnor U24460 (N_24460,N_24305,N_24315);
xnor U24461 (N_24461,N_24309,N_24375);
nor U24462 (N_24462,N_24279,N_24222);
nand U24463 (N_24463,N_24346,N_24379);
or U24464 (N_24464,N_24242,N_24237);
or U24465 (N_24465,N_24286,N_24390);
nor U24466 (N_24466,N_24316,N_24200);
and U24467 (N_24467,N_24223,N_24391);
nand U24468 (N_24468,N_24257,N_24399);
nand U24469 (N_24469,N_24324,N_24246);
nor U24470 (N_24470,N_24280,N_24239);
and U24471 (N_24471,N_24328,N_24338);
nor U24472 (N_24472,N_24254,N_24250);
or U24473 (N_24473,N_24298,N_24314);
nand U24474 (N_24474,N_24261,N_24388);
and U24475 (N_24475,N_24368,N_24337);
nand U24476 (N_24476,N_24226,N_24325);
nor U24477 (N_24477,N_24364,N_24295);
and U24478 (N_24478,N_24306,N_24267);
xnor U24479 (N_24479,N_24297,N_24231);
nor U24480 (N_24480,N_24201,N_24362);
nand U24481 (N_24481,N_24396,N_24386);
nor U24482 (N_24482,N_24285,N_24234);
or U24483 (N_24483,N_24349,N_24227);
or U24484 (N_24484,N_24385,N_24340);
or U24485 (N_24485,N_24308,N_24294);
xor U24486 (N_24486,N_24262,N_24358);
or U24487 (N_24487,N_24282,N_24301);
and U24488 (N_24488,N_24311,N_24207);
nor U24489 (N_24489,N_24206,N_24264);
and U24490 (N_24490,N_24312,N_24245);
or U24491 (N_24491,N_24289,N_24384);
nand U24492 (N_24492,N_24247,N_24381);
xor U24493 (N_24493,N_24339,N_24213);
nor U24494 (N_24494,N_24397,N_24211);
nand U24495 (N_24495,N_24288,N_24202);
or U24496 (N_24496,N_24218,N_24317);
and U24497 (N_24497,N_24345,N_24274);
nor U24498 (N_24498,N_24291,N_24343);
and U24499 (N_24499,N_24327,N_24276);
nand U24500 (N_24500,N_24272,N_24352);
and U24501 (N_24501,N_24318,N_24364);
and U24502 (N_24502,N_24227,N_24263);
nand U24503 (N_24503,N_24324,N_24347);
nor U24504 (N_24504,N_24270,N_24262);
or U24505 (N_24505,N_24303,N_24308);
nand U24506 (N_24506,N_24342,N_24248);
or U24507 (N_24507,N_24394,N_24310);
or U24508 (N_24508,N_24393,N_24266);
and U24509 (N_24509,N_24262,N_24224);
nor U24510 (N_24510,N_24336,N_24380);
xor U24511 (N_24511,N_24258,N_24246);
xor U24512 (N_24512,N_24220,N_24317);
nand U24513 (N_24513,N_24321,N_24387);
or U24514 (N_24514,N_24378,N_24249);
xor U24515 (N_24515,N_24317,N_24248);
xnor U24516 (N_24516,N_24296,N_24361);
xor U24517 (N_24517,N_24257,N_24397);
nor U24518 (N_24518,N_24217,N_24325);
xor U24519 (N_24519,N_24350,N_24339);
nor U24520 (N_24520,N_24257,N_24324);
or U24521 (N_24521,N_24280,N_24251);
nand U24522 (N_24522,N_24306,N_24331);
xnor U24523 (N_24523,N_24234,N_24265);
or U24524 (N_24524,N_24338,N_24276);
nor U24525 (N_24525,N_24231,N_24264);
nand U24526 (N_24526,N_24360,N_24344);
and U24527 (N_24527,N_24337,N_24232);
and U24528 (N_24528,N_24325,N_24328);
nor U24529 (N_24529,N_24320,N_24210);
nand U24530 (N_24530,N_24345,N_24247);
or U24531 (N_24531,N_24274,N_24238);
and U24532 (N_24532,N_24251,N_24377);
and U24533 (N_24533,N_24360,N_24373);
and U24534 (N_24534,N_24302,N_24247);
or U24535 (N_24535,N_24290,N_24269);
nor U24536 (N_24536,N_24272,N_24231);
nor U24537 (N_24537,N_24304,N_24255);
nand U24538 (N_24538,N_24336,N_24348);
or U24539 (N_24539,N_24293,N_24367);
or U24540 (N_24540,N_24229,N_24319);
nand U24541 (N_24541,N_24311,N_24237);
and U24542 (N_24542,N_24243,N_24220);
or U24543 (N_24543,N_24282,N_24276);
and U24544 (N_24544,N_24391,N_24325);
nand U24545 (N_24545,N_24297,N_24331);
nor U24546 (N_24546,N_24297,N_24395);
nand U24547 (N_24547,N_24249,N_24332);
nand U24548 (N_24548,N_24232,N_24248);
or U24549 (N_24549,N_24339,N_24273);
nor U24550 (N_24550,N_24307,N_24301);
xnor U24551 (N_24551,N_24340,N_24341);
nand U24552 (N_24552,N_24284,N_24259);
and U24553 (N_24553,N_24393,N_24276);
xnor U24554 (N_24554,N_24320,N_24303);
and U24555 (N_24555,N_24200,N_24319);
nand U24556 (N_24556,N_24241,N_24303);
xnor U24557 (N_24557,N_24385,N_24363);
nand U24558 (N_24558,N_24202,N_24375);
nor U24559 (N_24559,N_24221,N_24341);
xor U24560 (N_24560,N_24357,N_24335);
xor U24561 (N_24561,N_24229,N_24378);
nand U24562 (N_24562,N_24394,N_24207);
xor U24563 (N_24563,N_24395,N_24287);
xor U24564 (N_24564,N_24311,N_24233);
nand U24565 (N_24565,N_24297,N_24293);
xnor U24566 (N_24566,N_24363,N_24387);
or U24567 (N_24567,N_24219,N_24267);
nand U24568 (N_24568,N_24367,N_24360);
nor U24569 (N_24569,N_24369,N_24287);
nor U24570 (N_24570,N_24243,N_24316);
nand U24571 (N_24571,N_24279,N_24245);
nand U24572 (N_24572,N_24394,N_24324);
xnor U24573 (N_24573,N_24395,N_24385);
and U24574 (N_24574,N_24266,N_24272);
nand U24575 (N_24575,N_24384,N_24233);
xor U24576 (N_24576,N_24258,N_24224);
nand U24577 (N_24577,N_24297,N_24268);
and U24578 (N_24578,N_24231,N_24201);
nor U24579 (N_24579,N_24243,N_24350);
or U24580 (N_24580,N_24283,N_24397);
and U24581 (N_24581,N_24272,N_24386);
nor U24582 (N_24582,N_24362,N_24226);
or U24583 (N_24583,N_24393,N_24356);
and U24584 (N_24584,N_24389,N_24310);
nor U24585 (N_24585,N_24275,N_24218);
xnor U24586 (N_24586,N_24323,N_24379);
xor U24587 (N_24587,N_24274,N_24212);
xor U24588 (N_24588,N_24233,N_24249);
or U24589 (N_24589,N_24356,N_24376);
xor U24590 (N_24590,N_24300,N_24313);
and U24591 (N_24591,N_24262,N_24227);
xnor U24592 (N_24592,N_24301,N_24292);
or U24593 (N_24593,N_24392,N_24208);
xor U24594 (N_24594,N_24384,N_24394);
nor U24595 (N_24595,N_24389,N_24218);
nor U24596 (N_24596,N_24367,N_24374);
xnor U24597 (N_24597,N_24202,N_24214);
nand U24598 (N_24598,N_24350,N_24206);
nand U24599 (N_24599,N_24398,N_24318);
nand U24600 (N_24600,N_24588,N_24468);
and U24601 (N_24601,N_24430,N_24431);
nand U24602 (N_24602,N_24563,N_24577);
or U24603 (N_24603,N_24548,N_24469);
and U24604 (N_24604,N_24457,N_24579);
and U24605 (N_24605,N_24494,N_24446);
nand U24606 (N_24606,N_24454,N_24567);
xor U24607 (N_24607,N_24568,N_24480);
nor U24608 (N_24608,N_24515,N_24594);
nand U24609 (N_24609,N_24412,N_24463);
nor U24610 (N_24610,N_24542,N_24401);
or U24611 (N_24611,N_24429,N_24415);
or U24612 (N_24612,N_24524,N_24532);
nor U24613 (N_24613,N_24426,N_24505);
and U24614 (N_24614,N_24495,N_24525);
xor U24615 (N_24615,N_24417,N_24407);
nand U24616 (N_24616,N_24418,N_24572);
and U24617 (N_24617,N_24547,N_24441);
nand U24618 (N_24618,N_24482,N_24447);
xnor U24619 (N_24619,N_24526,N_24500);
nor U24620 (N_24620,N_24466,N_24599);
or U24621 (N_24621,N_24450,N_24484);
nor U24622 (N_24622,N_24486,N_24491);
and U24623 (N_24623,N_24479,N_24551);
nand U24624 (N_24624,N_24529,N_24459);
nand U24625 (N_24625,N_24522,N_24593);
nor U24626 (N_24626,N_24460,N_24443);
or U24627 (N_24627,N_24513,N_24553);
nor U24628 (N_24628,N_24562,N_24456);
or U24629 (N_24629,N_24424,N_24444);
and U24630 (N_24630,N_24506,N_24597);
and U24631 (N_24631,N_24591,N_24543);
or U24632 (N_24632,N_24538,N_24546);
or U24633 (N_24633,N_24509,N_24467);
and U24634 (N_24634,N_24428,N_24476);
nand U24635 (N_24635,N_24458,N_24590);
nand U24636 (N_24636,N_24580,N_24442);
nand U24637 (N_24637,N_24433,N_24474);
xor U24638 (N_24638,N_24560,N_24583);
or U24639 (N_24639,N_24581,N_24596);
and U24640 (N_24640,N_24473,N_24520);
nor U24641 (N_24641,N_24598,N_24478);
xor U24642 (N_24642,N_24425,N_24549);
nand U24643 (N_24643,N_24409,N_24496);
nand U24644 (N_24644,N_24592,N_24541);
or U24645 (N_24645,N_24406,N_24569);
nor U24646 (N_24646,N_24554,N_24517);
nor U24647 (N_24647,N_24492,N_24565);
xnor U24648 (N_24648,N_24497,N_24503);
nor U24649 (N_24649,N_24545,N_24574);
xor U24650 (N_24650,N_24435,N_24516);
nand U24651 (N_24651,N_24550,N_24576);
nand U24652 (N_24652,N_24531,N_24570);
xor U24653 (N_24653,N_24561,N_24556);
or U24654 (N_24654,N_24405,N_24451);
xor U24655 (N_24655,N_24512,N_24527);
and U24656 (N_24656,N_24534,N_24432);
nand U24657 (N_24657,N_24427,N_24566);
xnor U24658 (N_24658,N_24507,N_24502);
and U24659 (N_24659,N_24488,N_24521);
and U24660 (N_24660,N_24437,N_24552);
and U24661 (N_24661,N_24439,N_24540);
nand U24662 (N_24662,N_24436,N_24438);
nor U24663 (N_24663,N_24499,N_24481);
nor U24664 (N_24664,N_24421,N_24404);
xor U24665 (N_24665,N_24539,N_24575);
and U24666 (N_24666,N_24461,N_24571);
nor U24667 (N_24667,N_24408,N_24477);
xnor U24668 (N_24668,N_24555,N_24490);
xor U24669 (N_24669,N_24402,N_24470);
xnor U24670 (N_24670,N_24595,N_24558);
or U24671 (N_24671,N_24455,N_24519);
nor U24672 (N_24672,N_24416,N_24423);
xor U24673 (N_24673,N_24472,N_24518);
nor U24674 (N_24674,N_24587,N_24420);
or U24675 (N_24675,N_24536,N_24523);
nand U24676 (N_24676,N_24582,N_24448);
xnor U24677 (N_24677,N_24578,N_24535);
and U24678 (N_24678,N_24585,N_24537);
xnor U24679 (N_24679,N_24411,N_24413);
or U24680 (N_24680,N_24498,N_24528);
nand U24681 (N_24681,N_24487,N_24449);
or U24682 (N_24682,N_24564,N_24530);
and U24683 (N_24683,N_24445,N_24400);
or U24684 (N_24684,N_24434,N_24533);
nand U24685 (N_24685,N_24559,N_24464);
and U24686 (N_24686,N_24440,N_24403);
xnor U24687 (N_24687,N_24465,N_24511);
nand U24688 (N_24688,N_24471,N_24504);
nor U24689 (N_24689,N_24493,N_24414);
and U24690 (N_24690,N_24422,N_24489);
or U24691 (N_24691,N_24485,N_24586);
xor U24692 (N_24692,N_24410,N_24589);
nor U24693 (N_24693,N_24452,N_24510);
nand U24694 (N_24694,N_24475,N_24557);
and U24695 (N_24695,N_24419,N_24483);
or U24696 (N_24696,N_24453,N_24584);
or U24697 (N_24697,N_24573,N_24544);
and U24698 (N_24698,N_24514,N_24508);
xor U24699 (N_24699,N_24501,N_24462);
or U24700 (N_24700,N_24503,N_24586);
xnor U24701 (N_24701,N_24430,N_24554);
or U24702 (N_24702,N_24489,N_24412);
or U24703 (N_24703,N_24532,N_24436);
or U24704 (N_24704,N_24516,N_24508);
nand U24705 (N_24705,N_24484,N_24532);
nand U24706 (N_24706,N_24539,N_24595);
nand U24707 (N_24707,N_24425,N_24451);
nand U24708 (N_24708,N_24432,N_24536);
xor U24709 (N_24709,N_24431,N_24570);
or U24710 (N_24710,N_24431,N_24427);
or U24711 (N_24711,N_24539,N_24541);
nand U24712 (N_24712,N_24412,N_24470);
nor U24713 (N_24713,N_24425,N_24493);
and U24714 (N_24714,N_24520,N_24421);
and U24715 (N_24715,N_24548,N_24400);
nand U24716 (N_24716,N_24591,N_24516);
or U24717 (N_24717,N_24583,N_24470);
nor U24718 (N_24718,N_24597,N_24540);
nand U24719 (N_24719,N_24427,N_24476);
xor U24720 (N_24720,N_24401,N_24460);
and U24721 (N_24721,N_24568,N_24584);
nor U24722 (N_24722,N_24528,N_24583);
nor U24723 (N_24723,N_24514,N_24482);
or U24724 (N_24724,N_24476,N_24479);
and U24725 (N_24725,N_24573,N_24437);
or U24726 (N_24726,N_24406,N_24442);
and U24727 (N_24727,N_24518,N_24437);
xor U24728 (N_24728,N_24553,N_24507);
and U24729 (N_24729,N_24588,N_24549);
xnor U24730 (N_24730,N_24428,N_24493);
xnor U24731 (N_24731,N_24404,N_24597);
nand U24732 (N_24732,N_24576,N_24460);
and U24733 (N_24733,N_24408,N_24499);
nor U24734 (N_24734,N_24553,N_24510);
or U24735 (N_24735,N_24412,N_24563);
nor U24736 (N_24736,N_24422,N_24504);
nand U24737 (N_24737,N_24467,N_24457);
xnor U24738 (N_24738,N_24453,N_24527);
and U24739 (N_24739,N_24418,N_24550);
or U24740 (N_24740,N_24470,N_24512);
nor U24741 (N_24741,N_24558,N_24406);
nand U24742 (N_24742,N_24481,N_24574);
xor U24743 (N_24743,N_24502,N_24469);
xor U24744 (N_24744,N_24400,N_24424);
xor U24745 (N_24745,N_24430,N_24517);
nand U24746 (N_24746,N_24562,N_24520);
and U24747 (N_24747,N_24566,N_24523);
or U24748 (N_24748,N_24546,N_24449);
xor U24749 (N_24749,N_24454,N_24461);
nand U24750 (N_24750,N_24404,N_24598);
nor U24751 (N_24751,N_24506,N_24431);
or U24752 (N_24752,N_24472,N_24464);
xor U24753 (N_24753,N_24518,N_24572);
and U24754 (N_24754,N_24522,N_24429);
nor U24755 (N_24755,N_24558,N_24519);
nand U24756 (N_24756,N_24420,N_24433);
nor U24757 (N_24757,N_24402,N_24503);
nor U24758 (N_24758,N_24521,N_24496);
nor U24759 (N_24759,N_24567,N_24468);
nor U24760 (N_24760,N_24405,N_24587);
nor U24761 (N_24761,N_24598,N_24596);
nand U24762 (N_24762,N_24598,N_24491);
or U24763 (N_24763,N_24592,N_24416);
or U24764 (N_24764,N_24492,N_24431);
nand U24765 (N_24765,N_24470,N_24404);
nand U24766 (N_24766,N_24497,N_24523);
nor U24767 (N_24767,N_24541,N_24415);
xor U24768 (N_24768,N_24591,N_24560);
nand U24769 (N_24769,N_24512,N_24490);
xnor U24770 (N_24770,N_24505,N_24454);
nor U24771 (N_24771,N_24453,N_24463);
nor U24772 (N_24772,N_24498,N_24419);
and U24773 (N_24773,N_24419,N_24582);
xor U24774 (N_24774,N_24431,N_24408);
nor U24775 (N_24775,N_24552,N_24402);
and U24776 (N_24776,N_24417,N_24585);
and U24777 (N_24777,N_24580,N_24517);
nand U24778 (N_24778,N_24566,N_24537);
and U24779 (N_24779,N_24438,N_24548);
or U24780 (N_24780,N_24548,N_24573);
xnor U24781 (N_24781,N_24428,N_24466);
xor U24782 (N_24782,N_24506,N_24435);
xor U24783 (N_24783,N_24562,N_24583);
and U24784 (N_24784,N_24525,N_24444);
or U24785 (N_24785,N_24421,N_24438);
or U24786 (N_24786,N_24532,N_24541);
nor U24787 (N_24787,N_24540,N_24454);
xor U24788 (N_24788,N_24563,N_24516);
and U24789 (N_24789,N_24432,N_24550);
or U24790 (N_24790,N_24475,N_24584);
xnor U24791 (N_24791,N_24490,N_24435);
nand U24792 (N_24792,N_24575,N_24560);
nor U24793 (N_24793,N_24423,N_24542);
nor U24794 (N_24794,N_24525,N_24490);
nand U24795 (N_24795,N_24558,N_24464);
and U24796 (N_24796,N_24420,N_24574);
or U24797 (N_24797,N_24445,N_24530);
or U24798 (N_24798,N_24504,N_24501);
or U24799 (N_24799,N_24538,N_24506);
and U24800 (N_24800,N_24725,N_24763);
and U24801 (N_24801,N_24794,N_24607);
or U24802 (N_24802,N_24770,N_24667);
nor U24803 (N_24803,N_24745,N_24751);
nand U24804 (N_24804,N_24603,N_24731);
nor U24805 (N_24805,N_24672,N_24785);
nor U24806 (N_24806,N_24739,N_24711);
nor U24807 (N_24807,N_24764,N_24727);
nand U24808 (N_24808,N_24778,N_24605);
and U24809 (N_24809,N_24722,N_24704);
or U24810 (N_24810,N_24661,N_24736);
nand U24811 (N_24811,N_24760,N_24628);
xor U24812 (N_24812,N_24699,N_24749);
and U24813 (N_24813,N_24693,N_24681);
nor U24814 (N_24814,N_24659,N_24643);
xnor U24815 (N_24815,N_24617,N_24606);
nor U24816 (N_24816,N_24716,N_24653);
nand U24817 (N_24817,N_24608,N_24771);
xor U24818 (N_24818,N_24624,N_24774);
or U24819 (N_24819,N_24791,N_24639);
nor U24820 (N_24820,N_24650,N_24733);
nor U24821 (N_24821,N_24674,N_24756);
xor U24822 (N_24822,N_24720,N_24640);
xor U24823 (N_24823,N_24714,N_24796);
and U24824 (N_24824,N_24767,N_24792);
nor U24825 (N_24825,N_24780,N_24611);
nor U24826 (N_24826,N_24635,N_24743);
and U24827 (N_24827,N_24683,N_24726);
xor U24828 (N_24828,N_24737,N_24670);
nand U24829 (N_24829,N_24758,N_24612);
nor U24830 (N_24830,N_24710,N_24660);
xnor U24831 (N_24831,N_24729,N_24786);
nand U24832 (N_24832,N_24656,N_24684);
nand U24833 (N_24833,N_24676,N_24793);
or U24834 (N_24834,N_24679,N_24795);
xnor U24835 (N_24835,N_24788,N_24754);
nor U24836 (N_24836,N_24621,N_24782);
xor U24837 (N_24837,N_24644,N_24721);
or U24838 (N_24838,N_24610,N_24634);
and U24839 (N_24839,N_24787,N_24799);
nand U24840 (N_24840,N_24741,N_24759);
nor U24841 (N_24841,N_24772,N_24753);
or U24842 (N_24842,N_24709,N_24636);
xor U24843 (N_24843,N_24779,N_24776);
xor U24844 (N_24844,N_24750,N_24678);
xor U24845 (N_24845,N_24713,N_24632);
and U24846 (N_24846,N_24769,N_24789);
nand U24847 (N_24847,N_24762,N_24738);
and U24848 (N_24848,N_24673,N_24744);
or U24849 (N_24849,N_24680,N_24777);
nand U24850 (N_24850,N_24652,N_24641);
or U24851 (N_24851,N_24703,N_24658);
and U24852 (N_24852,N_24685,N_24616);
xor U24853 (N_24853,N_24696,N_24735);
nand U24854 (N_24854,N_24734,N_24798);
xnor U24855 (N_24855,N_24690,N_24651);
nand U24856 (N_24856,N_24723,N_24619);
nand U24857 (N_24857,N_24600,N_24757);
xnor U24858 (N_24858,N_24664,N_24614);
xor U24859 (N_24859,N_24613,N_24662);
nand U24860 (N_24860,N_24645,N_24648);
xor U24861 (N_24861,N_24627,N_24657);
nand U24862 (N_24862,N_24655,N_24626);
nor U24863 (N_24863,N_24695,N_24688);
nand U24864 (N_24864,N_24698,N_24638);
nand U24865 (N_24865,N_24668,N_24687);
xnor U24866 (N_24866,N_24761,N_24781);
and U24867 (N_24867,N_24712,N_24631);
nor U24868 (N_24868,N_24630,N_24748);
xor U24869 (N_24869,N_24718,N_24697);
or U24870 (N_24870,N_24752,N_24665);
xor U24871 (N_24871,N_24790,N_24728);
xor U24872 (N_24872,N_24620,N_24623);
nand U24873 (N_24873,N_24706,N_24675);
and U24874 (N_24874,N_24691,N_24707);
nand U24875 (N_24875,N_24689,N_24633);
nor U24876 (N_24876,N_24602,N_24647);
nor U24877 (N_24877,N_24654,N_24625);
nor U24878 (N_24878,N_24701,N_24646);
nand U24879 (N_24879,N_24717,N_24766);
or U24880 (N_24880,N_24784,N_24773);
nor U24881 (N_24881,N_24677,N_24740);
or U24882 (N_24882,N_24692,N_24666);
xnor U24883 (N_24883,N_24732,N_24629);
and U24884 (N_24884,N_24755,N_24622);
or U24885 (N_24885,N_24797,N_24669);
and U24886 (N_24886,N_24671,N_24747);
or U24887 (N_24887,N_24783,N_24746);
or U24888 (N_24888,N_24642,N_24702);
or U24889 (N_24889,N_24601,N_24708);
nand U24890 (N_24890,N_24686,N_24609);
nand U24891 (N_24891,N_24730,N_24705);
xnor U24892 (N_24892,N_24649,N_24719);
nand U24893 (N_24893,N_24663,N_24694);
and U24894 (N_24894,N_24700,N_24615);
and U24895 (N_24895,N_24724,N_24715);
and U24896 (N_24896,N_24618,N_24637);
or U24897 (N_24897,N_24768,N_24765);
nand U24898 (N_24898,N_24682,N_24775);
nor U24899 (N_24899,N_24604,N_24742);
and U24900 (N_24900,N_24695,N_24634);
and U24901 (N_24901,N_24751,N_24742);
and U24902 (N_24902,N_24655,N_24722);
nor U24903 (N_24903,N_24676,N_24615);
or U24904 (N_24904,N_24678,N_24608);
or U24905 (N_24905,N_24698,N_24658);
and U24906 (N_24906,N_24680,N_24764);
and U24907 (N_24907,N_24698,N_24649);
and U24908 (N_24908,N_24788,N_24637);
nand U24909 (N_24909,N_24606,N_24616);
nor U24910 (N_24910,N_24736,N_24669);
and U24911 (N_24911,N_24668,N_24663);
and U24912 (N_24912,N_24649,N_24633);
and U24913 (N_24913,N_24701,N_24792);
nor U24914 (N_24914,N_24635,N_24702);
nor U24915 (N_24915,N_24649,N_24767);
xor U24916 (N_24916,N_24682,N_24716);
nand U24917 (N_24917,N_24658,N_24788);
nor U24918 (N_24918,N_24744,N_24626);
nor U24919 (N_24919,N_24665,N_24606);
nand U24920 (N_24920,N_24696,N_24668);
or U24921 (N_24921,N_24700,N_24724);
xnor U24922 (N_24922,N_24661,N_24668);
or U24923 (N_24923,N_24722,N_24604);
xnor U24924 (N_24924,N_24666,N_24658);
nand U24925 (N_24925,N_24745,N_24605);
nor U24926 (N_24926,N_24774,N_24735);
or U24927 (N_24927,N_24742,N_24779);
nand U24928 (N_24928,N_24628,N_24658);
and U24929 (N_24929,N_24627,N_24620);
and U24930 (N_24930,N_24725,N_24613);
or U24931 (N_24931,N_24650,N_24631);
xnor U24932 (N_24932,N_24726,N_24730);
nor U24933 (N_24933,N_24618,N_24646);
or U24934 (N_24934,N_24656,N_24766);
nor U24935 (N_24935,N_24611,N_24703);
or U24936 (N_24936,N_24765,N_24675);
nor U24937 (N_24937,N_24793,N_24646);
and U24938 (N_24938,N_24783,N_24623);
or U24939 (N_24939,N_24775,N_24751);
or U24940 (N_24940,N_24760,N_24600);
nor U24941 (N_24941,N_24620,N_24628);
and U24942 (N_24942,N_24679,N_24633);
and U24943 (N_24943,N_24710,N_24772);
nand U24944 (N_24944,N_24721,N_24670);
and U24945 (N_24945,N_24649,N_24781);
nor U24946 (N_24946,N_24698,N_24770);
nand U24947 (N_24947,N_24678,N_24633);
nor U24948 (N_24948,N_24745,N_24711);
xnor U24949 (N_24949,N_24703,N_24705);
xor U24950 (N_24950,N_24741,N_24798);
xnor U24951 (N_24951,N_24684,N_24725);
xor U24952 (N_24952,N_24719,N_24772);
or U24953 (N_24953,N_24743,N_24696);
nor U24954 (N_24954,N_24644,N_24612);
nand U24955 (N_24955,N_24776,N_24667);
and U24956 (N_24956,N_24757,N_24771);
nand U24957 (N_24957,N_24602,N_24638);
xnor U24958 (N_24958,N_24649,N_24710);
or U24959 (N_24959,N_24780,N_24674);
nand U24960 (N_24960,N_24752,N_24720);
or U24961 (N_24961,N_24635,N_24785);
and U24962 (N_24962,N_24764,N_24618);
or U24963 (N_24963,N_24671,N_24721);
nand U24964 (N_24964,N_24658,N_24718);
nand U24965 (N_24965,N_24690,N_24698);
or U24966 (N_24966,N_24656,N_24738);
nor U24967 (N_24967,N_24613,N_24743);
or U24968 (N_24968,N_24747,N_24604);
and U24969 (N_24969,N_24602,N_24691);
xor U24970 (N_24970,N_24647,N_24663);
xnor U24971 (N_24971,N_24719,N_24690);
xnor U24972 (N_24972,N_24612,N_24682);
and U24973 (N_24973,N_24673,N_24727);
nand U24974 (N_24974,N_24657,N_24632);
xnor U24975 (N_24975,N_24736,N_24696);
nand U24976 (N_24976,N_24725,N_24714);
nor U24977 (N_24977,N_24623,N_24686);
nand U24978 (N_24978,N_24749,N_24705);
or U24979 (N_24979,N_24783,N_24727);
nor U24980 (N_24980,N_24780,N_24759);
xnor U24981 (N_24981,N_24698,N_24729);
or U24982 (N_24982,N_24659,N_24692);
or U24983 (N_24983,N_24657,N_24785);
and U24984 (N_24984,N_24688,N_24721);
nor U24985 (N_24985,N_24701,N_24707);
and U24986 (N_24986,N_24659,N_24798);
and U24987 (N_24987,N_24636,N_24610);
nor U24988 (N_24988,N_24650,N_24770);
xor U24989 (N_24989,N_24776,N_24773);
and U24990 (N_24990,N_24640,N_24734);
nor U24991 (N_24991,N_24675,N_24616);
and U24992 (N_24992,N_24667,N_24608);
nor U24993 (N_24993,N_24757,N_24737);
or U24994 (N_24994,N_24704,N_24636);
nand U24995 (N_24995,N_24647,N_24607);
nand U24996 (N_24996,N_24678,N_24644);
nand U24997 (N_24997,N_24744,N_24674);
xor U24998 (N_24998,N_24773,N_24671);
and U24999 (N_24999,N_24661,N_24630);
nand UO_0 (O_0,N_24813,N_24983);
and UO_1 (O_1,N_24911,N_24976);
or UO_2 (O_2,N_24988,N_24935);
xor UO_3 (O_3,N_24898,N_24861);
or UO_4 (O_4,N_24802,N_24975);
nand UO_5 (O_5,N_24932,N_24967);
nor UO_6 (O_6,N_24882,N_24874);
or UO_7 (O_7,N_24917,N_24930);
xor UO_8 (O_8,N_24926,N_24867);
nor UO_9 (O_9,N_24949,N_24998);
or UO_10 (O_10,N_24854,N_24948);
and UO_11 (O_11,N_24810,N_24960);
and UO_12 (O_12,N_24878,N_24916);
and UO_13 (O_13,N_24835,N_24837);
nor UO_14 (O_14,N_24872,N_24952);
and UO_15 (O_15,N_24938,N_24977);
and UO_16 (O_16,N_24929,N_24836);
nand UO_17 (O_17,N_24904,N_24841);
nor UO_18 (O_18,N_24886,N_24939);
nor UO_19 (O_19,N_24927,N_24907);
nand UO_20 (O_20,N_24961,N_24986);
nand UO_21 (O_21,N_24897,N_24857);
xnor UO_22 (O_22,N_24846,N_24879);
or UO_23 (O_23,N_24937,N_24944);
nor UO_24 (O_24,N_24995,N_24807);
xor UO_25 (O_25,N_24824,N_24829);
nand UO_26 (O_26,N_24893,N_24946);
or UO_27 (O_27,N_24808,N_24919);
xor UO_28 (O_28,N_24914,N_24803);
nand UO_29 (O_29,N_24945,N_24962);
or UO_30 (O_30,N_24955,N_24809);
and UO_31 (O_31,N_24902,N_24866);
and UO_32 (O_32,N_24931,N_24870);
nor UO_33 (O_33,N_24827,N_24853);
nand UO_34 (O_34,N_24966,N_24820);
and UO_35 (O_35,N_24964,N_24826);
nor UO_36 (O_36,N_24980,N_24801);
xnor UO_37 (O_37,N_24990,N_24905);
xnor UO_38 (O_38,N_24895,N_24934);
nand UO_39 (O_39,N_24974,N_24942);
or UO_40 (O_40,N_24881,N_24849);
and UO_41 (O_41,N_24873,N_24877);
nor UO_42 (O_42,N_24832,N_24892);
nor UO_43 (O_43,N_24959,N_24847);
and UO_44 (O_44,N_24869,N_24839);
xnor UO_45 (O_45,N_24868,N_24908);
xnor UO_46 (O_46,N_24963,N_24981);
nand UO_47 (O_47,N_24816,N_24830);
and UO_48 (O_48,N_24850,N_24915);
and UO_49 (O_49,N_24834,N_24989);
xnor UO_50 (O_50,N_24985,N_24888);
nand UO_51 (O_51,N_24860,N_24800);
nor UO_52 (O_52,N_24906,N_24936);
nand UO_53 (O_53,N_24855,N_24884);
nor UO_54 (O_54,N_24843,N_24954);
nand UO_55 (O_55,N_24896,N_24819);
and UO_56 (O_56,N_24994,N_24947);
xnor UO_57 (O_57,N_24865,N_24890);
nor UO_58 (O_58,N_24910,N_24970);
xor UO_59 (O_59,N_24968,N_24923);
and UO_60 (O_60,N_24821,N_24903);
nand UO_61 (O_61,N_24838,N_24979);
nand UO_62 (O_62,N_24925,N_24858);
nand UO_63 (O_63,N_24899,N_24871);
nor UO_64 (O_64,N_24842,N_24941);
or UO_65 (O_65,N_24912,N_24924);
xnor UO_66 (O_66,N_24862,N_24894);
nor UO_67 (O_67,N_24956,N_24920);
nand UO_68 (O_68,N_24823,N_24973);
and UO_69 (O_69,N_24805,N_24922);
nor UO_70 (O_70,N_24951,N_24844);
xor UO_71 (O_71,N_24928,N_24804);
nand UO_72 (O_72,N_24993,N_24969);
nand UO_73 (O_73,N_24984,N_24833);
or UO_74 (O_74,N_24814,N_24978);
or UO_75 (O_75,N_24996,N_24999);
and UO_76 (O_76,N_24883,N_24806);
and UO_77 (O_77,N_24933,N_24909);
and UO_78 (O_78,N_24859,N_24876);
or UO_79 (O_79,N_24811,N_24815);
xnor UO_80 (O_80,N_24840,N_24965);
and UO_81 (O_81,N_24953,N_24891);
and UO_82 (O_82,N_24831,N_24921);
xnor UO_83 (O_83,N_24887,N_24943);
or UO_84 (O_84,N_24913,N_24957);
and UO_85 (O_85,N_24987,N_24992);
nor UO_86 (O_86,N_24812,N_24918);
xor UO_87 (O_87,N_24848,N_24958);
xnor UO_88 (O_88,N_24900,N_24852);
or UO_89 (O_89,N_24818,N_24875);
or UO_90 (O_90,N_24822,N_24863);
or UO_91 (O_91,N_24940,N_24971);
nand UO_92 (O_92,N_24991,N_24901);
or UO_93 (O_93,N_24864,N_24817);
xnor UO_94 (O_94,N_24825,N_24982);
or UO_95 (O_95,N_24880,N_24856);
xor UO_96 (O_96,N_24950,N_24851);
nand UO_97 (O_97,N_24828,N_24845);
nor UO_98 (O_98,N_24885,N_24997);
or UO_99 (O_99,N_24972,N_24889);
nor UO_100 (O_100,N_24831,N_24879);
nand UO_101 (O_101,N_24997,N_24964);
nor UO_102 (O_102,N_24912,N_24920);
nand UO_103 (O_103,N_24815,N_24929);
and UO_104 (O_104,N_24987,N_24801);
nor UO_105 (O_105,N_24863,N_24893);
or UO_106 (O_106,N_24891,N_24894);
xnor UO_107 (O_107,N_24814,N_24878);
or UO_108 (O_108,N_24943,N_24882);
or UO_109 (O_109,N_24840,N_24937);
and UO_110 (O_110,N_24986,N_24941);
nand UO_111 (O_111,N_24834,N_24886);
xor UO_112 (O_112,N_24909,N_24869);
or UO_113 (O_113,N_24860,N_24901);
and UO_114 (O_114,N_24987,N_24931);
xnor UO_115 (O_115,N_24878,N_24957);
and UO_116 (O_116,N_24919,N_24874);
nor UO_117 (O_117,N_24885,N_24908);
or UO_118 (O_118,N_24968,N_24969);
nand UO_119 (O_119,N_24871,N_24982);
nor UO_120 (O_120,N_24907,N_24872);
nor UO_121 (O_121,N_24952,N_24839);
xnor UO_122 (O_122,N_24947,N_24859);
xor UO_123 (O_123,N_24814,N_24966);
xor UO_124 (O_124,N_24931,N_24990);
and UO_125 (O_125,N_24840,N_24946);
nor UO_126 (O_126,N_24892,N_24805);
nor UO_127 (O_127,N_24915,N_24815);
or UO_128 (O_128,N_24938,N_24872);
nor UO_129 (O_129,N_24880,N_24828);
nand UO_130 (O_130,N_24938,N_24879);
and UO_131 (O_131,N_24825,N_24894);
or UO_132 (O_132,N_24853,N_24869);
or UO_133 (O_133,N_24926,N_24933);
nor UO_134 (O_134,N_24994,N_24873);
xor UO_135 (O_135,N_24981,N_24872);
nor UO_136 (O_136,N_24912,N_24957);
nand UO_137 (O_137,N_24954,N_24997);
xor UO_138 (O_138,N_24827,N_24880);
nor UO_139 (O_139,N_24865,N_24922);
and UO_140 (O_140,N_24991,N_24804);
xor UO_141 (O_141,N_24879,N_24990);
nor UO_142 (O_142,N_24947,N_24964);
nand UO_143 (O_143,N_24909,N_24834);
xnor UO_144 (O_144,N_24886,N_24859);
nor UO_145 (O_145,N_24928,N_24965);
nor UO_146 (O_146,N_24886,N_24824);
nor UO_147 (O_147,N_24873,N_24820);
nor UO_148 (O_148,N_24992,N_24978);
xor UO_149 (O_149,N_24829,N_24963);
or UO_150 (O_150,N_24971,N_24871);
and UO_151 (O_151,N_24948,N_24873);
nor UO_152 (O_152,N_24852,N_24930);
nor UO_153 (O_153,N_24969,N_24865);
nor UO_154 (O_154,N_24867,N_24915);
nand UO_155 (O_155,N_24956,N_24922);
xor UO_156 (O_156,N_24946,N_24803);
nand UO_157 (O_157,N_24999,N_24887);
xnor UO_158 (O_158,N_24956,N_24840);
nand UO_159 (O_159,N_24821,N_24924);
xnor UO_160 (O_160,N_24985,N_24974);
xor UO_161 (O_161,N_24981,N_24843);
and UO_162 (O_162,N_24901,N_24913);
xnor UO_163 (O_163,N_24876,N_24803);
nand UO_164 (O_164,N_24846,N_24886);
nor UO_165 (O_165,N_24809,N_24913);
nand UO_166 (O_166,N_24972,N_24829);
and UO_167 (O_167,N_24806,N_24915);
nand UO_168 (O_168,N_24821,N_24993);
or UO_169 (O_169,N_24995,N_24808);
nor UO_170 (O_170,N_24998,N_24860);
and UO_171 (O_171,N_24922,N_24924);
or UO_172 (O_172,N_24952,N_24868);
or UO_173 (O_173,N_24832,N_24929);
nor UO_174 (O_174,N_24983,N_24864);
xor UO_175 (O_175,N_24985,N_24820);
nor UO_176 (O_176,N_24907,N_24904);
nor UO_177 (O_177,N_24949,N_24894);
or UO_178 (O_178,N_24990,N_24936);
xor UO_179 (O_179,N_24921,N_24850);
xor UO_180 (O_180,N_24860,N_24890);
and UO_181 (O_181,N_24919,N_24826);
or UO_182 (O_182,N_24848,N_24887);
xor UO_183 (O_183,N_24826,N_24900);
and UO_184 (O_184,N_24993,N_24818);
or UO_185 (O_185,N_24977,N_24901);
nor UO_186 (O_186,N_24906,N_24868);
nand UO_187 (O_187,N_24812,N_24907);
nand UO_188 (O_188,N_24891,N_24876);
and UO_189 (O_189,N_24852,N_24920);
nor UO_190 (O_190,N_24998,N_24842);
or UO_191 (O_191,N_24980,N_24831);
or UO_192 (O_192,N_24849,N_24879);
or UO_193 (O_193,N_24865,N_24914);
nand UO_194 (O_194,N_24895,N_24832);
xnor UO_195 (O_195,N_24979,N_24894);
or UO_196 (O_196,N_24908,N_24970);
and UO_197 (O_197,N_24839,N_24882);
nor UO_198 (O_198,N_24947,N_24980);
and UO_199 (O_199,N_24909,N_24811);
nor UO_200 (O_200,N_24886,N_24927);
and UO_201 (O_201,N_24980,N_24852);
and UO_202 (O_202,N_24943,N_24835);
xnor UO_203 (O_203,N_24948,N_24988);
nand UO_204 (O_204,N_24836,N_24960);
xnor UO_205 (O_205,N_24864,N_24925);
nor UO_206 (O_206,N_24820,N_24989);
nand UO_207 (O_207,N_24802,N_24873);
and UO_208 (O_208,N_24894,N_24842);
nor UO_209 (O_209,N_24980,N_24805);
nor UO_210 (O_210,N_24903,N_24951);
and UO_211 (O_211,N_24868,N_24958);
nand UO_212 (O_212,N_24912,N_24917);
and UO_213 (O_213,N_24915,N_24927);
xnor UO_214 (O_214,N_24857,N_24871);
xnor UO_215 (O_215,N_24922,N_24860);
and UO_216 (O_216,N_24843,N_24828);
or UO_217 (O_217,N_24968,N_24949);
xnor UO_218 (O_218,N_24840,N_24859);
or UO_219 (O_219,N_24883,N_24823);
xor UO_220 (O_220,N_24810,N_24819);
nor UO_221 (O_221,N_24834,N_24918);
xor UO_222 (O_222,N_24982,N_24879);
and UO_223 (O_223,N_24961,N_24982);
or UO_224 (O_224,N_24937,N_24989);
and UO_225 (O_225,N_24812,N_24894);
nor UO_226 (O_226,N_24900,N_24813);
nand UO_227 (O_227,N_24938,N_24953);
xnor UO_228 (O_228,N_24844,N_24804);
or UO_229 (O_229,N_24881,N_24971);
and UO_230 (O_230,N_24971,N_24879);
nand UO_231 (O_231,N_24899,N_24883);
xor UO_232 (O_232,N_24916,N_24906);
and UO_233 (O_233,N_24855,N_24990);
xor UO_234 (O_234,N_24940,N_24892);
nor UO_235 (O_235,N_24981,N_24826);
nand UO_236 (O_236,N_24961,N_24813);
and UO_237 (O_237,N_24907,N_24822);
or UO_238 (O_238,N_24838,N_24972);
or UO_239 (O_239,N_24839,N_24924);
and UO_240 (O_240,N_24815,N_24935);
xor UO_241 (O_241,N_24991,N_24899);
or UO_242 (O_242,N_24884,N_24849);
or UO_243 (O_243,N_24890,N_24972);
or UO_244 (O_244,N_24832,N_24932);
xor UO_245 (O_245,N_24886,N_24949);
nor UO_246 (O_246,N_24921,N_24881);
xor UO_247 (O_247,N_24989,N_24911);
or UO_248 (O_248,N_24847,N_24851);
or UO_249 (O_249,N_24971,N_24894);
and UO_250 (O_250,N_24919,N_24831);
nor UO_251 (O_251,N_24835,N_24869);
xnor UO_252 (O_252,N_24925,N_24936);
nor UO_253 (O_253,N_24957,N_24996);
and UO_254 (O_254,N_24824,N_24937);
and UO_255 (O_255,N_24888,N_24948);
or UO_256 (O_256,N_24808,N_24807);
nor UO_257 (O_257,N_24970,N_24831);
nand UO_258 (O_258,N_24896,N_24836);
or UO_259 (O_259,N_24972,N_24834);
nor UO_260 (O_260,N_24952,N_24834);
nor UO_261 (O_261,N_24977,N_24828);
or UO_262 (O_262,N_24813,N_24876);
and UO_263 (O_263,N_24973,N_24803);
nand UO_264 (O_264,N_24906,N_24819);
xnor UO_265 (O_265,N_24815,N_24870);
nand UO_266 (O_266,N_24832,N_24881);
xnor UO_267 (O_267,N_24933,N_24871);
or UO_268 (O_268,N_24845,N_24968);
nor UO_269 (O_269,N_24845,N_24818);
nor UO_270 (O_270,N_24803,N_24985);
xor UO_271 (O_271,N_24856,N_24816);
nor UO_272 (O_272,N_24896,N_24994);
nor UO_273 (O_273,N_24936,N_24885);
nand UO_274 (O_274,N_24809,N_24946);
and UO_275 (O_275,N_24981,N_24824);
nor UO_276 (O_276,N_24974,N_24891);
and UO_277 (O_277,N_24951,N_24837);
nor UO_278 (O_278,N_24817,N_24870);
or UO_279 (O_279,N_24950,N_24980);
nor UO_280 (O_280,N_24809,N_24885);
xor UO_281 (O_281,N_24949,N_24956);
and UO_282 (O_282,N_24936,N_24913);
nand UO_283 (O_283,N_24965,N_24818);
xnor UO_284 (O_284,N_24801,N_24832);
nor UO_285 (O_285,N_24822,N_24922);
xnor UO_286 (O_286,N_24957,N_24963);
xor UO_287 (O_287,N_24954,N_24973);
xor UO_288 (O_288,N_24834,N_24831);
nand UO_289 (O_289,N_24918,N_24946);
xnor UO_290 (O_290,N_24874,N_24886);
nand UO_291 (O_291,N_24828,N_24969);
and UO_292 (O_292,N_24959,N_24873);
or UO_293 (O_293,N_24965,N_24889);
nor UO_294 (O_294,N_24985,N_24956);
or UO_295 (O_295,N_24971,N_24800);
xor UO_296 (O_296,N_24864,N_24984);
nand UO_297 (O_297,N_24889,N_24895);
and UO_298 (O_298,N_24947,N_24974);
xnor UO_299 (O_299,N_24880,N_24943);
nor UO_300 (O_300,N_24938,N_24802);
xnor UO_301 (O_301,N_24945,N_24938);
or UO_302 (O_302,N_24952,N_24987);
and UO_303 (O_303,N_24847,N_24889);
xor UO_304 (O_304,N_24949,N_24864);
or UO_305 (O_305,N_24988,N_24874);
or UO_306 (O_306,N_24872,N_24848);
nand UO_307 (O_307,N_24916,N_24825);
nor UO_308 (O_308,N_24844,N_24900);
and UO_309 (O_309,N_24940,N_24810);
nor UO_310 (O_310,N_24870,N_24935);
or UO_311 (O_311,N_24864,N_24856);
xor UO_312 (O_312,N_24836,N_24900);
nand UO_313 (O_313,N_24802,N_24960);
nand UO_314 (O_314,N_24938,N_24822);
xnor UO_315 (O_315,N_24842,N_24868);
and UO_316 (O_316,N_24916,N_24943);
nand UO_317 (O_317,N_24975,N_24984);
and UO_318 (O_318,N_24892,N_24842);
xor UO_319 (O_319,N_24915,N_24861);
xor UO_320 (O_320,N_24974,N_24895);
and UO_321 (O_321,N_24862,N_24843);
and UO_322 (O_322,N_24812,N_24953);
and UO_323 (O_323,N_24892,N_24828);
or UO_324 (O_324,N_24884,N_24920);
and UO_325 (O_325,N_24972,N_24825);
and UO_326 (O_326,N_24962,N_24804);
nor UO_327 (O_327,N_24956,N_24882);
nand UO_328 (O_328,N_24920,N_24819);
or UO_329 (O_329,N_24822,N_24976);
nand UO_330 (O_330,N_24891,N_24813);
xnor UO_331 (O_331,N_24890,N_24821);
and UO_332 (O_332,N_24986,N_24805);
nor UO_333 (O_333,N_24900,N_24876);
nor UO_334 (O_334,N_24899,N_24858);
nor UO_335 (O_335,N_24964,N_24887);
or UO_336 (O_336,N_24869,N_24870);
and UO_337 (O_337,N_24948,N_24907);
and UO_338 (O_338,N_24894,N_24885);
and UO_339 (O_339,N_24915,N_24816);
nand UO_340 (O_340,N_24912,N_24835);
and UO_341 (O_341,N_24818,N_24952);
xor UO_342 (O_342,N_24949,N_24876);
xor UO_343 (O_343,N_24813,N_24948);
or UO_344 (O_344,N_24824,N_24920);
xor UO_345 (O_345,N_24815,N_24964);
nand UO_346 (O_346,N_24875,N_24874);
or UO_347 (O_347,N_24969,N_24880);
or UO_348 (O_348,N_24849,N_24957);
xnor UO_349 (O_349,N_24900,N_24984);
xnor UO_350 (O_350,N_24813,N_24916);
or UO_351 (O_351,N_24950,N_24965);
nand UO_352 (O_352,N_24947,N_24917);
and UO_353 (O_353,N_24837,N_24901);
or UO_354 (O_354,N_24852,N_24858);
or UO_355 (O_355,N_24963,N_24806);
xor UO_356 (O_356,N_24993,N_24823);
and UO_357 (O_357,N_24866,N_24817);
nand UO_358 (O_358,N_24845,N_24942);
and UO_359 (O_359,N_24907,N_24831);
nor UO_360 (O_360,N_24889,N_24846);
xor UO_361 (O_361,N_24875,N_24803);
or UO_362 (O_362,N_24974,N_24928);
xor UO_363 (O_363,N_24943,N_24969);
xor UO_364 (O_364,N_24937,N_24807);
or UO_365 (O_365,N_24827,N_24940);
or UO_366 (O_366,N_24846,N_24945);
nor UO_367 (O_367,N_24877,N_24979);
and UO_368 (O_368,N_24813,N_24810);
or UO_369 (O_369,N_24920,N_24903);
or UO_370 (O_370,N_24847,N_24838);
nor UO_371 (O_371,N_24958,N_24814);
and UO_372 (O_372,N_24805,N_24877);
nor UO_373 (O_373,N_24932,N_24876);
xnor UO_374 (O_374,N_24815,N_24980);
and UO_375 (O_375,N_24929,N_24813);
and UO_376 (O_376,N_24829,N_24997);
or UO_377 (O_377,N_24854,N_24913);
nand UO_378 (O_378,N_24821,N_24805);
nand UO_379 (O_379,N_24936,N_24835);
xor UO_380 (O_380,N_24865,N_24887);
or UO_381 (O_381,N_24887,N_24840);
and UO_382 (O_382,N_24925,N_24916);
xor UO_383 (O_383,N_24956,N_24935);
nor UO_384 (O_384,N_24809,N_24923);
nand UO_385 (O_385,N_24921,N_24982);
or UO_386 (O_386,N_24823,N_24884);
and UO_387 (O_387,N_24856,N_24979);
nor UO_388 (O_388,N_24807,N_24875);
or UO_389 (O_389,N_24823,N_24858);
xnor UO_390 (O_390,N_24898,N_24866);
nand UO_391 (O_391,N_24822,N_24960);
or UO_392 (O_392,N_24975,N_24995);
nor UO_393 (O_393,N_24831,N_24869);
nand UO_394 (O_394,N_24818,N_24947);
or UO_395 (O_395,N_24848,N_24806);
or UO_396 (O_396,N_24866,N_24969);
nor UO_397 (O_397,N_24835,N_24816);
or UO_398 (O_398,N_24966,N_24806);
or UO_399 (O_399,N_24811,N_24816);
nand UO_400 (O_400,N_24934,N_24996);
nand UO_401 (O_401,N_24989,N_24983);
or UO_402 (O_402,N_24882,N_24958);
and UO_403 (O_403,N_24961,N_24975);
nor UO_404 (O_404,N_24879,N_24832);
nor UO_405 (O_405,N_24877,N_24941);
and UO_406 (O_406,N_24937,N_24956);
xnor UO_407 (O_407,N_24887,N_24941);
nand UO_408 (O_408,N_24937,N_24899);
nand UO_409 (O_409,N_24990,N_24875);
nor UO_410 (O_410,N_24819,N_24836);
nand UO_411 (O_411,N_24820,N_24907);
xnor UO_412 (O_412,N_24993,N_24953);
or UO_413 (O_413,N_24995,N_24846);
xor UO_414 (O_414,N_24841,N_24840);
nand UO_415 (O_415,N_24837,N_24881);
nor UO_416 (O_416,N_24872,N_24804);
nor UO_417 (O_417,N_24880,N_24906);
and UO_418 (O_418,N_24832,N_24913);
xnor UO_419 (O_419,N_24859,N_24965);
nor UO_420 (O_420,N_24970,N_24842);
and UO_421 (O_421,N_24977,N_24953);
nor UO_422 (O_422,N_24833,N_24811);
or UO_423 (O_423,N_24809,N_24901);
xnor UO_424 (O_424,N_24827,N_24969);
nand UO_425 (O_425,N_24826,N_24897);
nor UO_426 (O_426,N_24959,N_24813);
xnor UO_427 (O_427,N_24938,N_24849);
nand UO_428 (O_428,N_24973,N_24809);
and UO_429 (O_429,N_24874,N_24855);
nand UO_430 (O_430,N_24965,N_24802);
xor UO_431 (O_431,N_24818,N_24995);
nand UO_432 (O_432,N_24989,N_24875);
xor UO_433 (O_433,N_24998,N_24939);
or UO_434 (O_434,N_24984,N_24989);
nand UO_435 (O_435,N_24832,N_24964);
nor UO_436 (O_436,N_24886,N_24814);
nand UO_437 (O_437,N_24820,N_24954);
nor UO_438 (O_438,N_24968,N_24999);
xor UO_439 (O_439,N_24851,N_24906);
nor UO_440 (O_440,N_24930,N_24836);
and UO_441 (O_441,N_24940,N_24847);
or UO_442 (O_442,N_24814,N_24998);
or UO_443 (O_443,N_24867,N_24909);
xnor UO_444 (O_444,N_24967,N_24857);
nor UO_445 (O_445,N_24897,N_24975);
and UO_446 (O_446,N_24949,N_24840);
or UO_447 (O_447,N_24856,N_24804);
nor UO_448 (O_448,N_24948,N_24951);
and UO_449 (O_449,N_24818,N_24847);
or UO_450 (O_450,N_24894,N_24921);
and UO_451 (O_451,N_24830,N_24971);
or UO_452 (O_452,N_24962,N_24864);
xnor UO_453 (O_453,N_24958,N_24970);
xor UO_454 (O_454,N_24956,N_24831);
or UO_455 (O_455,N_24826,N_24899);
and UO_456 (O_456,N_24908,N_24886);
xor UO_457 (O_457,N_24968,N_24988);
nor UO_458 (O_458,N_24953,N_24963);
nand UO_459 (O_459,N_24912,N_24887);
nor UO_460 (O_460,N_24834,N_24868);
nor UO_461 (O_461,N_24899,N_24998);
nor UO_462 (O_462,N_24919,N_24887);
xnor UO_463 (O_463,N_24997,N_24838);
xor UO_464 (O_464,N_24965,N_24845);
nor UO_465 (O_465,N_24846,N_24868);
xnor UO_466 (O_466,N_24903,N_24872);
nand UO_467 (O_467,N_24922,N_24952);
and UO_468 (O_468,N_24838,N_24874);
nand UO_469 (O_469,N_24878,N_24800);
xnor UO_470 (O_470,N_24878,N_24993);
nand UO_471 (O_471,N_24925,N_24904);
or UO_472 (O_472,N_24872,N_24855);
or UO_473 (O_473,N_24806,N_24934);
and UO_474 (O_474,N_24876,N_24968);
or UO_475 (O_475,N_24893,N_24966);
nor UO_476 (O_476,N_24831,N_24855);
or UO_477 (O_477,N_24951,N_24819);
and UO_478 (O_478,N_24828,N_24829);
or UO_479 (O_479,N_24960,N_24940);
nand UO_480 (O_480,N_24931,N_24825);
xnor UO_481 (O_481,N_24986,N_24852);
nand UO_482 (O_482,N_24968,N_24951);
nor UO_483 (O_483,N_24889,N_24906);
xor UO_484 (O_484,N_24960,N_24803);
nand UO_485 (O_485,N_24849,N_24882);
and UO_486 (O_486,N_24968,N_24890);
nor UO_487 (O_487,N_24845,N_24947);
nand UO_488 (O_488,N_24831,N_24849);
xor UO_489 (O_489,N_24800,N_24865);
and UO_490 (O_490,N_24900,N_24818);
and UO_491 (O_491,N_24943,N_24803);
xnor UO_492 (O_492,N_24979,N_24853);
or UO_493 (O_493,N_24952,N_24880);
nor UO_494 (O_494,N_24937,N_24814);
or UO_495 (O_495,N_24817,N_24903);
xnor UO_496 (O_496,N_24808,N_24949);
and UO_497 (O_497,N_24975,N_24905);
xor UO_498 (O_498,N_24968,N_24880);
nand UO_499 (O_499,N_24839,N_24965);
and UO_500 (O_500,N_24925,N_24982);
xor UO_501 (O_501,N_24939,N_24841);
and UO_502 (O_502,N_24974,N_24922);
xnor UO_503 (O_503,N_24940,N_24965);
nand UO_504 (O_504,N_24886,N_24945);
nand UO_505 (O_505,N_24814,N_24902);
nand UO_506 (O_506,N_24878,N_24910);
and UO_507 (O_507,N_24910,N_24815);
nand UO_508 (O_508,N_24895,N_24802);
xnor UO_509 (O_509,N_24870,N_24915);
or UO_510 (O_510,N_24864,N_24990);
nand UO_511 (O_511,N_24885,N_24987);
nor UO_512 (O_512,N_24800,N_24889);
or UO_513 (O_513,N_24858,N_24912);
xnor UO_514 (O_514,N_24995,N_24855);
xnor UO_515 (O_515,N_24979,N_24867);
nor UO_516 (O_516,N_24975,N_24852);
nand UO_517 (O_517,N_24941,N_24894);
nand UO_518 (O_518,N_24901,N_24950);
and UO_519 (O_519,N_24817,N_24824);
nand UO_520 (O_520,N_24894,N_24934);
or UO_521 (O_521,N_24987,N_24975);
xnor UO_522 (O_522,N_24815,N_24966);
xnor UO_523 (O_523,N_24946,N_24884);
and UO_524 (O_524,N_24810,N_24949);
nor UO_525 (O_525,N_24948,N_24916);
and UO_526 (O_526,N_24947,N_24907);
nand UO_527 (O_527,N_24930,N_24956);
xnor UO_528 (O_528,N_24937,N_24971);
nor UO_529 (O_529,N_24852,N_24907);
or UO_530 (O_530,N_24954,N_24926);
and UO_531 (O_531,N_24874,N_24846);
nand UO_532 (O_532,N_24999,N_24826);
or UO_533 (O_533,N_24900,N_24825);
nor UO_534 (O_534,N_24932,N_24923);
xnor UO_535 (O_535,N_24975,N_24922);
xnor UO_536 (O_536,N_24993,N_24961);
or UO_537 (O_537,N_24914,N_24968);
nor UO_538 (O_538,N_24813,N_24868);
nand UO_539 (O_539,N_24936,N_24996);
or UO_540 (O_540,N_24905,N_24878);
nor UO_541 (O_541,N_24807,N_24828);
and UO_542 (O_542,N_24961,N_24879);
or UO_543 (O_543,N_24944,N_24864);
xor UO_544 (O_544,N_24849,N_24878);
and UO_545 (O_545,N_24864,N_24874);
or UO_546 (O_546,N_24862,N_24807);
nand UO_547 (O_547,N_24987,N_24915);
nand UO_548 (O_548,N_24857,N_24822);
nand UO_549 (O_549,N_24852,N_24952);
and UO_550 (O_550,N_24959,N_24915);
xor UO_551 (O_551,N_24909,N_24891);
or UO_552 (O_552,N_24945,N_24892);
or UO_553 (O_553,N_24913,N_24856);
or UO_554 (O_554,N_24902,N_24868);
or UO_555 (O_555,N_24993,N_24813);
nor UO_556 (O_556,N_24819,N_24878);
or UO_557 (O_557,N_24954,N_24862);
nand UO_558 (O_558,N_24944,N_24932);
and UO_559 (O_559,N_24871,N_24855);
nor UO_560 (O_560,N_24946,N_24831);
nand UO_561 (O_561,N_24919,N_24917);
xnor UO_562 (O_562,N_24899,N_24867);
nor UO_563 (O_563,N_24968,N_24871);
or UO_564 (O_564,N_24922,N_24815);
and UO_565 (O_565,N_24983,N_24899);
or UO_566 (O_566,N_24918,N_24861);
and UO_567 (O_567,N_24892,N_24841);
nor UO_568 (O_568,N_24873,N_24945);
nor UO_569 (O_569,N_24922,N_24800);
xor UO_570 (O_570,N_24860,N_24968);
nand UO_571 (O_571,N_24812,N_24961);
and UO_572 (O_572,N_24905,N_24844);
or UO_573 (O_573,N_24821,N_24940);
or UO_574 (O_574,N_24983,N_24849);
xnor UO_575 (O_575,N_24901,N_24850);
xnor UO_576 (O_576,N_24844,N_24908);
nor UO_577 (O_577,N_24906,N_24972);
or UO_578 (O_578,N_24803,N_24904);
and UO_579 (O_579,N_24828,N_24982);
and UO_580 (O_580,N_24880,N_24819);
or UO_581 (O_581,N_24940,N_24942);
nand UO_582 (O_582,N_24987,N_24963);
xnor UO_583 (O_583,N_24900,N_24811);
nor UO_584 (O_584,N_24973,N_24870);
and UO_585 (O_585,N_24854,N_24928);
nand UO_586 (O_586,N_24966,N_24950);
xor UO_587 (O_587,N_24855,N_24964);
and UO_588 (O_588,N_24925,N_24997);
nor UO_589 (O_589,N_24857,N_24983);
xor UO_590 (O_590,N_24800,N_24854);
nand UO_591 (O_591,N_24978,N_24988);
nand UO_592 (O_592,N_24859,N_24853);
nor UO_593 (O_593,N_24832,N_24839);
nand UO_594 (O_594,N_24936,N_24862);
or UO_595 (O_595,N_24953,N_24905);
nor UO_596 (O_596,N_24813,N_24895);
nand UO_597 (O_597,N_24972,N_24806);
or UO_598 (O_598,N_24957,N_24950);
or UO_599 (O_599,N_24913,N_24906);
nand UO_600 (O_600,N_24823,N_24835);
nor UO_601 (O_601,N_24960,N_24821);
nand UO_602 (O_602,N_24988,N_24853);
and UO_603 (O_603,N_24820,N_24963);
nand UO_604 (O_604,N_24961,N_24963);
nor UO_605 (O_605,N_24988,N_24980);
and UO_606 (O_606,N_24929,N_24970);
xor UO_607 (O_607,N_24968,N_24998);
xor UO_608 (O_608,N_24931,N_24866);
nand UO_609 (O_609,N_24943,N_24978);
nand UO_610 (O_610,N_24949,N_24820);
and UO_611 (O_611,N_24995,N_24953);
nor UO_612 (O_612,N_24995,N_24840);
nor UO_613 (O_613,N_24852,N_24985);
nor UO_614 (O_614,N_24958,N_24931);
and UO_615 (O_615,N_24946,N_24923);
nor UO_616 (O_616,N_24812,N_24833);
nand UO_617 (O_617,N_24857,N_24811);
nor UO_618 (O_618,N_24820,N_24919);
and UO_619 (O_619,N_24968,N_24915);
xor UO_620 (O_620,N_24930,N_24921);
and UO_621 (O_621,N_24853,N_24840);
nand UO_622 (O_622,N_24858,N_24875);
or UO_623 (O_623,N_24880,N_24895);
or UO_624 (O_624,N_24833,N_24891);
or UO_625 (O_625,N_24936,N_24952);
and UO_626 (O_626,N_24804,N_24914);
nand UO_627 (O_627,N_24932,N_24945);
nand UO_628 (O_628,N_24866,N_24909);
and UO_629 (O_629,N_24877,N_24848);
nor UO_630 (O_630,N_24855,N_24951);
or UO_631 (O_631,N_24887,N_24895);
nor UO_632 (O_632,N_24827,N_24924);
nand UO_633 (O_633,N_24880,N_24891);
or UO_634 (O_634,N_24831,N_24825);
nand UO_635 (O_635,N_24981,N_24899);
nor UO_636 (O_636,N_24801,N_24842);
and UO_637 (O_637,N_24875,N_24870);
and UO_638 (O_638,N_24820,N_24868);
nor UO_639 (O_639,N_24879,N_24911);
nor UO_640 (O_640,N_24989,N_24885);
and UO_641 (O_641,N_24959,N_24897);
nand UO_642 (O_642,N_24989,N_24916);
nor UO_643 (O_643,N_24958,N_24926);
xor UO_644 (O_644,N_24906,N_24933);
nand UO_645 (O_645,N_24847,N_24874);
nand UO_646 (O_646,N_24926,N_24826);
nand UO_647 (O_647,N_24931,N_24809);
nor UO_648 (O_648,N_24910,N_24902);
xnor UO_649 (O_649,N_24960,N_24847);
or UO_650 (O_650,N_24933,N_24823);
nand UO_651 (O_651,N_24839,N_24855);
nor UO_652 (O_652,N_24869,N_24942);
or UO_653 (O_653,N_24884,N_24877);
nor UO_654 (O_654,N_24931,N_24843);
xnor UO_655 (O_655,N_24950,N_24921);
nor UO_656 (O_656,N_24958,N_24825);
xnor UO_657 (O_657,N_24940,N_24980);
nor UO_658 (O_658,N_24979,N_24957);
nor UO_659 (O_659,N_24833,N_24874);
or UO_660 (O_660,N_24857,N_24851);
and UO_661 (O_661,N_24867,N_24820);
xnor UO_662 (O_662,N_24983,N_24924);
and UO_663 (O_663,N_24898,N_24972);
nor UO_664 (O_664,N_24929,N_24940);
or UO_665 (O_665,N_24839,N_24934);
xnor UO_666 (O_666,N_24819,N_24827);
nand UO_667 (O_667,N_24874,N_24978);
or UO_668 (O_668,N_24942,N_24804);
nand UO_669 (O_669,N_24987,N_24867);
nor UO_670 (O_670,N_24864,N_24821);
or UO_671 (O_671,N_24894,N_24922);
and UO_672 (O_672,N_24820,N_24939);
nor UO_673 (O_673,N_24854,N_24930);
or UO_674 (O_674,N_24832,N_24976);
or UO_675 (O_675,N_24854,N_24992);
nand UO_676 (O_676,N_24807,N_24895);
xor UO_677 (O_677,N_24828,N_24933);
and UO_678 (O_678,N_24903,N_24812);
xnor UO_679 (O_679,N_24856,N_24922);
or UO_680 (O_680,N_24968,N_24863);
or UO_681 (O_681,N_24988,N_24990);
or UO_682 (O_682,N_24800,N_24884);
nand UO_683 (O_683,N_24896,N_24852);
nand UO_684 (O_684,N_24954,N_24992);
xor UO_685 (O_685,N_24913,N_24871);
nor UO_686 (O_686,N_24891,N_24921);
nand UO_687 (O_687,N_24852,N_24892);
or UO_688 (O_688,N_24935,N_24864);
nor UO_689 (O_689,N_24855,N_24894);
xor UO_690 (O_690,N_24828,N_24944);
or UO_691 (O_691,N_24893,N_24905);
and UO_692 (O_692,N_24840,N_24920);
nor UO_693 (O_693,N_24959,N_24921);
nor UO_694 (O_694,N_24924,N_24918);
nor UO_695 (O_695,N_24846,N_24838);
xor UO_696 (O_696,N_24978,N_24829);
xor UO_697 (O_697,N_24891,N_24910);
and UO_698 (O_698,N_24827,N_24985);
xor UO_699 (O_699,N_24981,N_24819);
and UO_700 (O_700,N_24820,N_24999);
xor UO_701 (O_701,N_24810,N_24908);
or UO_702 (O_702,N_24905,N_24804);
nand UO_703 (O_703,N_24879,N_24905);
and UO_704 (O_704,N_24987,N_24802);
nand UO_705 (O_705,N_24905,N_24944);
nand UO_706 (O_706,N_24934,N_24901);
nor UO_707 (O_707,N_24831,N_24824);
xor UO_708 (O_708,N_24876,N_24878);
and UO_709 (O_709,N_24952,N_24884);
or UO_710 (O_710,N_24904,N_24930);
nand UO_711 (O_711,N_24827,N_24972);
xor UO_712 (O_712,N_24838,N_24942);
and UO_713 (O_713,N_24870,N_24981);
nand UO_714 (O_714,N_24870,N_24950);
xor UO_715 (O_715,N_24811,N_24886);
nand UO_716 (O_716,N_24914,N_24948);
xor UO_717 (O_717,N_24892,N_24928);
nand UO_718 (O_718,N_24894,N_24879);
nor UO_719 (O_719,N_24928,N_24815);
nand UO_720 (O_720,N_24833,N_24858);
or UO_721 (O_721,N_24838,N_24920);
or UO_722 (O_722,N_24818,N_24929);
or UO_723 (O_723,N_24992,N_24845);
and UO_724 (O_724,N_24837,N_24962);
and UO_725 (O_725,N_24919,N_24916);
or UO_726 (O_726,N_24921,N_24935);
xor UO_727 (O_727,N_24989,N_24999);
or UO_728 (O_728,N_24902,N_24816);
xnor UO_729 (O_729,N_24933,N_24818);
nor UO_730 (O_730,N_24839,N_24914);
and UO_731 (O_731,N_24921,N_24878);
and UO_732 (O_732,N_24837,N_24842);
and UO_733 (O_733,N_24884,N_24829);
nor UO_734 (O_734,N_24993,N_24867);
or UO_735 (O_735,N_24907,N_24943);
and UO_736 (O_736,N_24961,N_24995);
nor UO_737 (O_737,N_24906,N_24944);
and UO_738 (O_738,N_24800,N_24841);
nand UO_739 (O_739,N_24917,N_24950);
nor UO_740 (O_740,N_24940,N_24922);
or UO_741 (O_741,N_24870,N_24904);
nor UO_742 (O_742,N_24972,N_24864);
xnor UO_743 (O_743,N_24942,N_24832);
nor UO_744 (O_744,N_24990,N_24876);
nor UO_745 (O_745,N_24945,N_24854);
xnor UO_746 (O_746,N_24906,N_24947);
nand UO_747 (O_747,N_24911,N_24832);
nor UO_748 (O_748,N_24972,N_24807);
or UO_749 (O_749,N_24898,N_24821);
or UO_750 (O_750,N_24918,N_24984);
nor UO_751 (O_751,N_24820,N_24840);
xor UO_752 (O_752,N_24982,N_24854);
or UO_753 (O_753,N_24888,N_24806);
nor UO_754 (O_754,N_24990,N_24862);
nor UO_755 (O_755,N_24906,N_24986);
xnor UO_756 (O_756,N_24916,N_24992);
nor UO_757 (O_757,N_24884,N_24832);
or UO_758 (O_758,N_24903,N_24813);
or UO_759 (O_759,N_24904,N_24963);
xnor UO_760 (O_760,N_24851,N_24838);
nand UO_761 (O_761,N_24913,N_24979);
nor UO_762 (O_762,N_24802,N_24890);
xnor UO_763 (O_763,N_24958,N_24831);
or UO_764 (O_764,N_24858,N_24855);
or UO_765 (O_765,N_24971,N_24896);
and UO_766 (O_766,N_24881,N_24835);
or UO_767 (O_767,N_24914,N_24915);
nand UO_768 (O_768,N_24944,N_24860);
and UO_769 (O_769,N_24813,N_24962);
or UO_770 (O_770,N_24856,N_24994);
and UO_771 (O_771,N_24916,N_24966);
and UO_772 (O_772,N_24893,N_24830);
nand UO_773 (O_773,N_24809,N_24974);
and UO_774 (O_774,N_24970,N_24829);
or UO_775 (O_775,N_24955,N_24916);
nand UO_776 (O_776,N_24931,N_24985);
and UO_777 (O_777,N_24941,N_24993);
and UO_778 (O_778,N_24910,N_24845);
nand UO_779 (O_779,N_24861,N_24889);
nand UO_780 (O_780,N_24860,N_24810);
nor UO_781 (O_781,N_24958,N_24817);
nand UO_782 (O_782,N_24968,N_24944);
or UO_783 (O_783,N_24936,N_24945);
and UO_784 (O_784,N_24844,N_24948);
xnor UO_785 (O_785,N_24803,N_24864);
or UO_786 (O_786,N_24935,N_24812);
nor UO_787 (O_787,N_24900,N_24919);
nor UO_788 (O_788,N_24999,N_24952);
xnor UO_789 (O_789,N_24918,N_24840);
nor UO_790 (O_790,N_24923,N_24970);
xnor UO_791 (O_791,N_24877,N_24893);
nor UO_792 (O_792,N_24810,N_24871);
nand UO_793 (O_793,N_24834,N_24835);
xor UO_794 (O_794,N_24811,N_24867);
nand UO_795 (O_795,N_24817,N_24806);
and UO_796 (O_796,N_24811,N_24916);
or UO_797 (O_797,N_24839,N_24803);
nand UO_798 (O_798,N_24986,N_24919);
xor UO_799 (O_799,N_24999,N_24825);
xnor UO_800 (O_800,N_24914,N_24960);
and UO_801 (O_801,N_24908,N_24802);
and UO_802 (O_802,N_24803,N_24993);
nand UO_803 (O_803,N_24928,N_24895);
or UO_804 (O_804,N_24944,N_24985);
xor UO_805 (O_805,N_24811,N_24876);
nand UO_806 (O_806,N_24928,N_24866);
xor UO_807 (O_807,N_24835,N_24870);
and UO_808 (O_808,N_24905,N_24923);
and UO_809 (O_809,N_24871,N_24819);
nand UO_810 (O_810,N_24852,N_24946);
xnor UO_811 (O_811,N_24837,N_24898);
and UO_812 (O_812,N_24917,N_24975);
nor UO_813 (O_813,N_24888,N_24868);
nor UO_814 (O_814,N_24900,N_24966);
and UO_815 (O_815,N_24834,N_24948);
nor UO_816 (O_816,N_24822,N_24974);
nor UO_817 (O_817,N_24842,N_24832);
nor UO_818 (O_818,N_24884,N_24944);
nor UO_819 (O_819,N_24929,N_24833);
xor UO_820 (O_820,N_24961,N_24862);
or UO_821 (O_821,N_24940,N_24862);
nor UO_822 (O_822,N_24856,N_24865);
xor UO_823 (O_823,N_24877,N_24830);
or UO_824 (O_824,N_24939,N_24893);
nor UO_825 (O_825,N_24973,N_24886);
and UO_826 (O_826,N_24925,N_24892);
xnor UO_827 (O_827,N_24849,N_24839);
nand UO_828 (O_828,N_24901,N_24899);
nor UO_829 (O_829,N_24896,N_24895);
nand UO_830 (O_830,N_24868,N_24957);
nor UO_831 (O_831,N_24808,N_24806);
nand UO_832 (O_832,N_24853,N_24882);
and UO_833 (O_833,N_24836,N_24850);
nand UO_834 (O_834,N_24808,N_24865);
or UO_835 (O_835,N_24885,N_24857);
nand UO_836 (O_836,N_24983,N_24945);
nand UO_837 (O_837,N_24823,N_24803);
and UO_838 (O_838,N_24822,N_24862);
nand UO_839 (O_839,N_24832,N_24907);
or UO_840 (O_840,N_24985,N_24884);
xor UO_841 (O_841,N_24897,N_24955);
xnor UO_842 (O_842,N_24893,N_24843);
nor UO_843 (O_843,N_24984,N_24834);
nor UO_844 (O_844,N_24802,N_24945);
or UO_845 (O_845,N_24966,N_24981);
or UO_846 (O_846,N_24828,N_24801);
or UO_847 (O_847,N_24836,N_24925);
nor UO_848 (O_848,N_24874,N_24848);
and UO_849 (O_849,N_24980,N_24937);
nand UO_850 (O_850,N_24900,N_24891);
and UO_851 (O_851,N_24870,N_24947);
and UO_852 (O_852,N_24912,N_24908);
xnor UO_853 (O_853,N_24987,N_24926);
or UO_854 (O_854,N_24843,N_24890);
xor UO_855 (O_855,N_24862,N_24993);
nor UO_856 (O_856,N_24885,N_24827);
and UO_857 (O_857,N_24839,N_24940);
xnor UO_858 (O_858,N_24913,N_24865);
nand UO_859 (O_859,N_24912,N_24867);
or UO_860 (O_860,N_24865,N_24908);
or UO_861 (O_861,N_24991,N_24985);
or UO_862 (O_862,N_24804,N_24881);
xnor UO_863 (O_863,N_24852,N_24808);
nand UO_864 (O_864,N_24905,N_24989);
or UO_865 (O_865,N_24813,N_24901);
nand UO_866 (O_866,N_24881,N_24985);
and UO_867 (O_867,N_24890,N_24928);
xor UO_868 (O_868,N_24948,N_24953);
xnor UO_869 (O_869,N_24814,N_24813);
nand UO_870 (O_870,N_24824,N_24909);
nand UO_871 (O_871,N_24807,N_24932);
xnor UO_872 (O_872,N_24862,N_24888);
nand UO_873 (O_873,N_24878,N_24856);
xnor UO_874 (O_874,N_24933,N_24953);
and UO_875 (O_875,N_24843,N_24891);
xnor UO_876 (O_876,N_24972,N_24940);
or UO_877 (O_877,N_24996,N_24850);
nor UO_878 (O_878,N_24876,N_24828);
nand UO_879 (O_879,N_24926,N_24804);
nand UO_880 (O_880,N_24942,N_24871);
and UO_881 (O_881,N_24826,N_24931);
and UO_882 (O_882,N_24876,N_24874);
nor UO_883 (O_883,N_24844,N_24876);
nand UO_884 (O_884,N_24914,N_24985);
xnor UO_885 (O_885,N_24827,N_24989);
or UO_886 (O_886,N_24852,N_24810);
or UO_887 (O_887,N_24941,N_24878);
nand UO_888 (O_888,N_24903,N_24893);
nand UO_889 (O_889,N_24840,N_24951);
nand UO_890 (O_890,N_24995,N_24819);
xnor UO_891 (O_891,N_24955,N_24847);
nor UO_892 (O_892,N_24837,N_24966);
nand UO_893 (O_893,N_24982,N_24940);
nand UO_894 (O_894,N_24898,N_24962);
and UO_895 (O_895,N_24926,N_24907);
and UO_896 (O_896,N_24930,N_24995);
xnor UO_897 (O_897,N_24857,N_24892);
xor UO_898 (O_898,N_24975,N_24864);
or UO_899 (O_899,N_24807,N_24892);
nand UO_900 (O_900,N_24853,N_24960);
nand UO_901 (O_901,N_24873,N_24965);
nand UO_902 (O_902,N_24981,N_24935);
nand UO_903 (O_903,N_24866,N_24970);
and UO_904 (O_904,N_24989,N_24847);
or UO_905 (O_905,N_24809,N_24857);
or UO_906 (O_906,N_24818,N_24905);
xor UO_907 (O_907,N_24873,N_24885);
nor UO_908 (O_908,N_24946,N_24966);
nand UO_909 (O_909,N_24808,N_24830);
and UO_910 (O_910,N_24819,N_24924);
or UO_911 (O_911,N_24894,N_24806);
nand UO_912 (O_912,N_24992,N_24876);
nor UO_913 (O_913,N_24833,N_24978);
nor UO_914 (O_914,N_24823,N_24862);
and UO_915 (O_915,N_24817,N_24928);
xnor UO_916 (O_916,N_24951,N_24811);
and UO_917 (O_917,N_24952,N_24809);
nand UO_918 (O_918,N_24846,N_24853);
or UO_919 (O_919,N_24975,N_24837);
and UO_920 (O_920,N_24939,N_24977);
nor UO_921 (O_921,N_24866,N_24914);
and UO_922 (O_922,N_24862,N_24919);
xor UO_923 (O_923,N_24985,N_24811);
nor UO_924 (O_924,N_24838,N_24921);
and UO_925 (O_925,N_24875,N_24816);
nor UO_926 (O_926,N_24804,N_24898);
xor UO_927 (O_927,N_24833,N_24821);
nand UO_928 (O_928,N_24835,N_24962);
xor UO_929 (O_929,N_24816,N_24888);
and UO_930 (O_930,N_24878,N_24826);
or UO_931 (O_931,N_24988,N_24954);
xor UO_932 (O_932,N_24898,N_24870);
nand UO_933 (O_933,N_24876,N_24934);
nor UO_934 (O_934,N_24966,N_24917);
and UO_935 (O_935,N_24859,N_24928);
and UO_936 (O_936,N_24980,N_24872);
or UO_937 (O_937,N_24919,N_24939);
or UO_938 (O_938,N_24927,N_24866);
or UO_939 (O_939,N_24996,N_24910);
or UO_940 (O_940,N_24801,N_24804);
and UO_941 (O_941,N_24821,N_24949);
nand UO_942 (O_942,N_24955,N_24926);
xor UO_943 (O_943,N_24833,N_24860);
nand UO_944 (O_944,N_24949,N_24836);
xor UO_945 (O_945,N_24896,N_24891);
xnor UO_946 (O_946,N_24887,N_24934);
and UO_947 (O_947,N_24871,N_24868);
and UO_948 (O_948,N_24985,N_24964);
nand UO_949 (O_949,N_24878,N_24824);
nand UO_950 (O_950,N_24952,N_24866);
or UO_951 (O_951,N_24992,N_24831);
or UO_952 (O_952,N_24872,N_24941);
and UO_953 (O_953,N_24809,N_24884);
or UO_954 (O_954,N_24807,N_24866);
nand UO_955 (O_955,N_24975,N_24821);
and UO_956 (O_956,N_24938,N_24866);
nor UO_957 (O_957,N_24877,N_24938);
or UO_958 (O_958,N_24864,N_24927);
and UO_959 (O_959,N_24882,N_24880);
and UO_960 (O_960,N_24821,N_24989);
and UO_961 (O_961,N_24826,N_24962);
or UO_962 (O_962,N_24865,N_24999);
xor UO_963 (O_963,N_24903,N_24825);
and UO_964 (O_964,N_24967,N_24949);
xnor UO_965 (O_965,N_24903,N_24807);
or UO_966 (O_966,N_24985,N_24949);
xor UO_967 (O_967,N_24869,N_24889);
nand UO_968 (O_968,N_24810,N_24832);
nor UO_969 (O_969,N_24976,N_24876);
nand UO_970 (O_970,N_24948,N_24909);
nand UO_971 (O_971,N_24882,N_24983);
nor UO_972 (O_972,N_24894,N_24961);
nor UO_973 (O_973,N_24822,N_24962);
nor UO_974 (O_974,N_24973,N_24992);
or UO_975 (O_975,N_24982,N_24962);
or UO_976 (O_976,N_24837,N_24856);
or UO_977 (O_977,N_24922,N_24976);
and UO_978 (O_978,N_24917,N_24956);
nor UO_979 (O_979,N_24910,N_24888);
xor UO_980 (O_980,N_24857,N_24913);
and UO_981 (O_981,N_24811,N_24986);
nand UO_982 (O_982,N_24983,N_24808);
nor UO_983 (O_983,N_24994,N_24969);
nor UO_984 (O_984,N_24932,N_24817);
or UO_985 (O_985,N_24955,N_24852);
or UO_986 (O_986,N_24886,N_24845);
and UO_987 (O_987,N_24811,N_24887);
xor UO_988 (O_988,N_24995,N_24914);
nor UO_989 (O_989,N_24830,N_24868);
xnor UO_990 (O_990,N_24839,N_24916);
or UO_991 (O_991,N_24910,N_24955);
or UO_992 (O_992,N_24877,N_24813);
nor UO_993 (O_993,N_24965,N_24952);
and UO_994 (O_994,N_24979,N_24924);
nand UO_995 (O_995,N_24893,N_24991);
nor UO_996 (O_996,N_24968,N_24908);
xnor UO_997 (O_997,N_24901,N_24988);
nand UO_998 (O_998,N_24964,N_24988);
xor UO_999 (O_999,N_24985,N_24934);
or UO_1000 (O_1000,N_24883,N_24808);
xnor UO_1001 (O_1001,N_24882,N_24968);
and UO_1002 (O_1002,N_24957,N_24942);
xnor UO_1003 (O_1003,N_24887,N_24806);
or UO_1004 (O_1004,N_24813,N_24835);
or UO_1005 (O_1005,N_24949,N_24873);
or UO_1006 (O_1006,N_24978,N_24894);
nand UO_1007 (O_1007,N_24805,N_24981);
nand UO_1008 (O_1008,N_24838,N_24869);
xnor UO_1009 (O_1009,N_24886,N_24922);
or UO_1010 (O_1010,N_24881,N_24866);
nand UO_1011 (O_1011,N_24935,N_24915);
nand UO_1012 (O_1012,N_24976,N_24867);
xor UO_1013 (O_1013,N_24878,N_24974);
nand UO_1014 (O_1014,N_24903,N_24834);
nand UO_1015 (O_1015,N_24915,N_24812);
nor UO_1016 (O_1016,N_24871,N_24998);
xor UO_1017 (O_1017,N_24806,N_24843);
nand UO_1018 (O_1018,N_24825,N_24966);
and UO_1019 (O_1019,N_24879,N_24985);
nand UO_1020 (O_1020,N_24891,N_24878);
nand UO_1021 (O_1021,N_24965,N_24820);
or UO_1022 (O_1022,N_24855,N_24934);
or UO_1023 (O_1023,N_24909,N_24829);
and UO_1024 (O_1024,N_24882,N_24810);
nor UO_1025 (O_1025,N_24939,N_24836);
nor UO_1026 (O_1026,N_24854,N_24909);
xnor UO_1027 (O_1027,N_24929,N_24872);
nand UO_1028 (O_1028,N_24905,N_24919);
and UO_1029 (O_1029,N_24983,N_24852);
and UO_1030 (O_1030,N_24897,N_24941);
nor UO_1031 (O_1031,N_24888,N_24974);
and UO_1032 (O_1032,N_24959,N_24931);
xor UO_1033 (O_1033,N_24834,N_24951);
nand UO_1034 (O_1034,N_24964,N_24806);
xnor UO_1035 (O_1035,N_24905,N_24918);
xnor UO_1036 (O_1036,N_24886,N_24931);
or UO_1037 (O_1037,N_24988,N_24906);
nor UO_1038 (O_1038,N_24822,N_24873);
and UO_1039 (O_1039,N_24839,N_24935);
and UO_1040 (O_1040,N_24841,N_24936);
and UO_1041 (O_1041,N_24815,N_24852);
or UO_1042 (O_1042,N_24836,N_24941);
xor UO_1043 (O_1043,N_24822,N_24817);
nand UO_1044 (O_1044,N_24945,N_24800);
and UO_1045 (O_1045,N_24919,N_24971);
nand UO_1046 (O_1046,N_24882,N_24982);
nor UO_1047 (O_1047,N_24914,N_24895);
xor UO_1048 (O_1048,N_24991,N_24826);
and UO_1049 (O_1049,N_24921,N_24848);
or UO_1050 (O_1050,N_24801,N_24946);
and UO_1051 (O_1051,N_24886,N_24817);
xor UO_1052 (O_1052,N_24857,N_24865);
nor UO_1053 (O_1053,N_24821,N_24888);
nand UO_1054 (O_1054,N_24899,N_24808);
or UO_1055 (O_1055,N_24977,N_24945);
xnor UO_1056 (O_1056,N_24937,N_24964);
nand UO_1057 (O_1057,N_24839,N_24861);
or UO_1058 (O_1058,N_24809,N_24904);
xor UO_1059 (O_1059,N_24998,N_24811);
and UO_1060 (O_1060,N_24929,N_24904);
or UO_1061 (O_1061,N_24844,N_24996);
xnor UO_1062 (O_1062,N_24975,N_24883);
and UO_1063 (O_1063,N_24845,N_24854);
nand UO_1064 (O_1064,N_24867,N_24876);
or UO_1065 (O_1065,N_24930,N_24929);
nor UO_1066 (O_1066,N_24820,N_24880);
nor UO_1067 (O_1067,N_24938,N_24851);
nand UO_1068 (O_1068,N_24992,N_24855);
nor UO_1069 (O_1069,N_24849,N_24967);
nor UO_1070 (O_1070,N_24973,N_24891);
xor UO_1071 (O_1071,N_24832,N_24953);
and UO_1072 (O_1072,N_24879,N_24996);
nor UO_1073 (O_1073,N_24805,N_24806);
xor UO_1074 (O_1074,N_24887,N_24946);
nand UO_1075 (O_1075,N_24956,N_24852);
and UO_1076 (O_1076,N_24931,N_24928);
xnor UO_1077 (O_1077,N_24953,N_24874);
nor UO_1078 (O_1078,N_24817,N_24995);
nor UO_1079 (O_1079,N_24952,N_24945);
nand UO_1080 (O_1080,N_24905,N_24908);
and UO_1081 (O_1081,N_24926,N_24978);
nor UO_1082 (O_1082,N_24825,N_24961);
and UO_1083 (O_1083,N_24938,N_24874);
nor UO_1084 (O_1084,N_24991,N_24840);
xor UO_1085 (O_1085,N_24820,N_24851);
or UO_1086 (O_1086,N_24961,N_24968);
or UO_1087 (O_1087,N_24885,N_24836);
and UO_1088 (O_1088,N_24910,N_24834);
and UO_1089 (O_1089,N_24925,N_24970);
nand UO_1090 (O_1090,N_24804,N_24808);
and UO_1091 (O_1091,N_24810,N_24853);
or UO_1092 (O_1092,N_24943,N_24879);
xor UO_1093 (O_1093,N_24972,N_24921);
nor UO_1094 (O_1094,N_24879,N_24862);
nand UO_1095 (O_1095,N_24949,N_24889);
xnor UO_1096 (O_1096,N_24904,N_24882);
and UO_1097 (O_1097,N_24876,N_24936);
and UO_1098 (O_1098,N_24843,N_24902);
nand UO_1099 (O_1099,N_24958,N_24916);
nor UO_1100 (O_1100,N_24863,N_24814);
and UO_1101 (O_1101,N_24839,N_24864);
nand UO_1102 (O_1102,N_24995,N_24900);
xnor UO_1103 (O_1103,N_24831,N_24812);
or UO_1104 (O_1104,N_24811,N_24927);
xnor UO_1105 (O_1105,N_24981,N_24977);
nor UO_1106 (O_1106,N_24856,N_24859);
and UO_1107 (O_1107,N_24978,N_24998);
or UO_1108 (O_1108,N_24938,N_24993);
and UO_1109 (O_1109,N_24835,N_24849);
xor UO_1110 (O_1110,N_24897,N_24839);
or UO_1111 (O_1111,N_24888,N_24972);
and UO_1112 (O_1112,N_24842,N_24846);
nand UO_1113 (O_1113,N_24971,N_24965);
nor UO_1114 (O_1114,N_24951,N_24990);
or UO_1115 (O_1115,N_24919,N_24922);
xnor UO_1116 (O_1116,N_24979,N_24976);
xnor UO_1117 (O_1117,N_24988,N_24909);
and UO_1118 (O_1118,N_24890,N_24957);
and UO_1119 (O_1119,N_24909,N_24973);
xor UO_1120 (O_1120,N_24821,N_24869);
and UO_1121 (O_1121,N_24821,N_24965);
xor UO_1122 (O_1122,N_24810,N_24850);
or UO_1123 (O_1123,N_24936,N_24940);
nor UO_1124 (O_1124,N_24943,N_24829);
nor UO_1125 (O_1125,N_24857,N_24908);
and UO_1126 (O_1126,N_24985,N_24995);
xnor UO_1127 (O_1127,N_24941,N_24998);
xnor UO_1128 (O_1128,N_24828,N_24822);
nor UO_1129 (O_1129,N_24919,N_24813);
and UO_1130 (O_1130,N_24909,N_24857);
nor UO_1131 (O_1131,N_24820,N_24957);
and UO_1132 (O_1132,N_24807,N_24889);
or UO_1133 (O_1133,N_24811,N_24941);
nand UO_1134 (O_1134,N_24837,N_24958);
xor UO_1135 (O_1135,N_24864,N_24950);
xor UO_1136 (O_1136,N_24955,N_24888);
and UO_1137 (O_1137,N_24887,N_24813);
nor UO_1138 (O_1138,N_24901,N_24808);
nor UO_1139 (O_1139,N_24967,N_24982);
and UO_1140 (O_1140,N_24847,N_24999);
or UO_1141 (O_1141,N_24933,N_24853);
or UO_1142 (O_1142,N_24884,N_24995);
nand UO_1143 (O_1143,N_24869,N_24830);
xnor UO_1144 (O_1144,N_24813,N_24989);
nor UO_1145 (O_1145,N_24828,N_24907);
xnor UO_1146 (O_1146,N_24934,N_24884);
nand UO_1147 (O_1147,N_24905,N_24888);
nand UO_1148 (O_1148,N_24839,N_24885);
xnor UO_1149 (O_1149,N_24817,N_24855);
xor UO_1150 (O_1150,N_24879,N_24994);
xnor UO_1151 (O_1151,N_24999,N_24900);
xnor UO_1152 (O_1152,N_24852,N_24909);
xnor UO_1153 (O_1153,N_24920,N_24859);
and UO_1154 (O_1154,N_24919,N_24854);
or UO_1155 (O_1155,N_24869,N_24949);
nand UO_1156 (O_1156,N_24851,N_24899);
or UO_1157 (O_1157,N_24996,N_24894);
or UO_1158 (O_1158,N_24853,N_24901);
xnor UO_1159 (O_1159,N_24809,N_24929);
xnor UO_1160 (O_1160,N_24973,N_24957);
and UO_1161 (O_1161,N_24862,N_24998);
or UO_1162 (O_1162,N_24959,N_24888);
xnor UO_1163 (O_1163,N_24896,N_24927);
and UO_1164 (O_1164,N_24938,N_24834);
and UO_1165 (O_1165,N_24932,N_24857);
xnor UO_1166 (O_1166,N_24949,N_24922);
or UO_1167 (O_1167,N_24991,N_24888);
or UO_1168 (O_1168,N_24998,N_24918);
nor UO_1169 (O_1169,N_24832,N_24818);
and UO_1170 (O_1170,N_24932,N_24809);
nand UO_1171 (O_1171,N_24926,N_24889);
nand UO_1172 (O_1172,N_24917,N_24962);
nor UO_1173 (O_1173,N_24852,N_24961);
or UO_1174 (O_1174,N_24972,N_24885);
nand UO_1175 (O_1175,N_24803,N_24989);
and UO_1176 (O_1176,N_24865,N_24945);
and UO_1177 (O_1177,N_24978,N_24996);
nor UO_1178 (O_1178,N_24923,N_24911);
nand UO_1179 (O_1179,N_24801,N_24827);
nor UO_1180 (O_1180,N_24956,N_24860);
or UO_1181 (O_1181,N_24826,N_24963);
nand UO_1182 (O_1182,N_24993,N_24936);
xnor UO_1183 (O_1183,N_24814,N_24907);
or UO_1184 (O_1184,N_24909,N_24945);
or UO_1185 (O_1185,N_24963,N_24994);
and UO_1186 (O_1186,N_24967,N_24882);
nor UO_1187 (O_1187,N_24831,N_24854);
nand UO_1188 (O_1188,N_24807,N_24805);
nor UO_1189 (O_1189,N_24896,N_24911);
nand UO_1190 (O_1190,N_24865,N_24925);
or UO_1191 (O_1191,N_24958,N_24948);
xnor UO_1192 (O_1192,N_24932,N_24819);
nor UO_1193 (O_1193,N_24929,N_24948);
and UO_1194 (O_1194,N_24983,N_24874);
and UO_1195 (O_1195,N_24852,N_24941);
and UO_1196 (O_1196,N_24931,N_24805);
xor UO_1197 (O_1197,N_24849,N_24952);
nor UO_1198 (O_1198,N_24961,N_24850);
nor UO_1199 (O_1199,N_24811,N_24801);
or UO_1200 (O_1200,N_24854,N_24803);
or UO_1201 (O_1201,N_24879,N_24821);
nand UO_1202 (O_1202,N_24976,N_24875);
and UO_1203 (O_1203,N_24913,N_24883);
xnor UO_1204 (O_1204,N_24901,N_24851);
nand UO_1205 (O_1205,N_24826,N_24986);
nor UO_1206 (O_1206,N_24890,N_24884);
or UO_1207 (O_1207,N_24806,N_24912);
and UO_1208 (O_1208,N_24961,N_24991);
nand UO_1209 (O_1209,N_24855,N_24915);
xnor UO_1210 (O_1210,N_24970,N_24857);
nand UO_1211 (O_1211,N_24959,N_24987);
nand UO_1212 (O_1212,N_24935,N_24879);
nand UO_1213 (O_1213,N_24892,N_24874);
nor UO_1214 (O_1214,N_24917,N_24847);
and UO_1215 (O_1215,N_24957,N_24837);
or UO_1216 (O_1216,N_24820,N_24958);
xnor UO_1217 (O_1217,N_24831,N_24863);
or UO_1218 (O_1218,N_24948,N_24884);
or UO_1219 (O_1219,N_24992,N_24830);
nand UO_1220 (O_1220,N_24851,N_24815);
xor UO_1221 (O_1221,N_24868,N_24924);
and UO_1222 (O_1222,N_24851,N_24852);
nand UO_1223 (O_1223,N_24838,N_24985);
or UO_1224 (O_1224,N_24944,N_24867);
and UO_1225 (O_1225,N_24813,N_24875);
xor UO_1226 (O_1226,N_24959,N_24817);
xor UO_1227 (O_1227,N_24926,N_24896);
or UO_1228 (O_1228,N_24988,N_24908);
nor UO_1229 (O_1229,N_24833,N_24889);
xor UO_1230 (O_1230,N_24997,N_24927);
and UO_1231 (O_1231,N_24871,N_24879);
nor UO_1232 (O_1232,N_24936,N_24811);
xnor UO_1233 (O_1233,N_24968,N_24832);
xnor UO_1234 (O_1234,N_24883,N_24919);
xnor UO_1235 (O_1235,N_24819,N_24857);
nor UO_1236 (O_1236,N_24822,N_24909);
xnor UO_1237 (O_1237,N_24962,N_24814);
xnor UO_1238 (O_1238,N_24871,N_24983);
nand UO_1239 (O_1239,N_24921,N_24834);
and UO_1240 (O_1240,N_24950,N_24928);
and UO_1241 (O_1241,N_24910,N_24838);
xor UO_1242 (O_1242,N_24952,N_24926);
and UO_1243 (O_1243,N_24883,N_24908);
nand UO_1244 (O_1244,N_24899,N_24917);
nor UO_1245 (O_1245,N_24970,N_24961);
nand UO_1246 (O_1246,N_24869,N_24849);
nand UO_1247 (O_1247,N_24894,N_24983);
nor UO_1248 (O_1248,N_24852,N_24992);
xnor UO_1249 (O_1249,N_24897,N_24931);
and UO_1250 (O_1250,N_24915,N_24819);
or UO_1251 (O_1251,N_24928,N_24938);
or UO_1252 (O_1252,N_24899,N_24994);
nor UO_1253 (O_1253,N_24869,N_24986);
or UO_1254 (O_1254,N_24827,N_24823);
or UO_1255 (O_1255,N_24872,N_24970);
or UO_1256 (O_1256,N_24815,N_24819);
and UO_1257 (O_1257,N_24942,N_24884);
nor UO_1258 (O_1258,N_24896,N_24849);
or UO_1259 (O_1259,N_24983,N_24883);
and UO_1260 (O_1260,N_24834,N_24968);
nand UO_1261 (O_1261,N_24864,N_24981);
xnor UO_1262 (O_1262,N_24890,N_24866);
nor UO_1263 (O_1263,N_24924,N_24969);
and UO_1264 (O_1264,N_24928,N_24987);
xnor UO_1265 (O_1265,N_24842,N_24864);
xnor UO_1266 (O_1266,N_24944,N_24832);
nand UO_1267 (O_1267,N_24837,N_24996);
nor UO_1268 (O_1268,N_24863,N_24918);
nand UO_1269 (O_1269,N_24908,N_24987);
nand UO_1270 (O_1270,N_24962,N_24842);
nand UO_1271 (O_1271,N_24890,N_24844);
and UO_1272 (O_1272,N_24862,N_24941);
nand UO_1273 (O_1273,N_24830,N_24875);
or UO_1274 (O_1274,N_24987,N_24887);
or UO_1275 (O_1275,N_24940,N_24860);
nand UO_1276 (O_1276,N_24941,N_24948);
and UO_1277 (O_1277,N_24955,N_24807);
nor UO_1278 (O_1278,N_24914,N_24850);
and UO_1279 (O_1279,N_24914,N_24844);
and UO_1280 (O_1280,N_24812,N_24825);
or UO_1281 (O_1281,N_24855,N_24950);
or UO_1282 (O_1282,N_24986,N_24867);
xor UO_1283 (O_1283,N_24834,N_24883);
nand UO_1284 (O_1284,N_24962,N_24900);
nand UO_1285 (O_1285,N_24977,N_24883);
xnor UO_1286 (O_1286,N_24820,N_24940);
nand UO_1287 (O_1287,N_24893,N_24880);
nor UO_1288 (O_1288,N_24813,N_24985);
or UO_1289 (O_1289,N_24965,N_24972);
or UO_1290 (O_1290,N_24934,N_24831);
nor UO_1291 (O_1291,N_24952,N_24810);
xnor UO_1292 (O_1292,N_24912,N_24885);
nor UO_1293 (O_1293,N_24994,N_24840);
nand UO_1294 (O_1294,N_24868,N_24839);
or UO_1295 (O_1295,N_24875,N_24811);
or UO_1296 (O_1296,N_24921,N_24875);
nor UO_1297 (O_1297,N_24993,N_24929);
nor UO_1298 (O_1298,N_24851,N_24802);
and UO_1299 (O_1299,N_24885,N_24945);
nand UO_1300 (O_1300,N_24950,N_24868);
or UO_1301 (O_1301,N_24999,N_24850);
and UO_1302 (O_1302,N_24914,N_24950);
and UO_1303 (O_1303,N_24941,N_24957);
or UO_1304 (O_1304,N_24953,N_24841);
xnor UO_1305 (O_1305,N_24933,N_24810);
nand UO_1306 (O_1306,N_24959,N_24842);
nor UO_1307 (O_1307,N_24857,N_24838);
and UO_1308 (O_1308,N_24902,N_24917);
and UO_1309 (O_1309,N_24847,N_24945);
nor UO_1310 (O_1310,N_24969,N_24896);
nor UO_1311 (O_1311,N_24996,N_24871);
and UO_1312 (O_1312,N_24855,N_24977);
and UO_1313 (O_1313,N_24980,N_24816);
xor UO_1314 (O_1314,N_24934,N_24910);
and UO_1315 (O_1315,N_24954,N_24887);
and UO_1316 (O_1316,N_24944,N_24967);
and UO_1317 (O_1317,N_24855,N_24865);
nor UO_1318 (O_1318,N_24985,N_24844);
or UO_1319 (O_1319,N_24859,N_24819);
xnor UO_1320 (O_1320,N_24831,N_24940);
or UO_1321 (O_1321,N_24903,N_24928);
xor UO_1322 (O_1322,N_24826,N_24813);
nand UO_1323 (O_1323,N_24836,N_24883);
nand UO_1324 (O_1324,N_24812,N_24942);
nand UO_1325 (O_1325,N_24823,N_24923);
and UO_1326 (O_1326,N_24904,N_24878);
xor UO_1327 (O_1327,N_24970,N_24927);
nand UO_1328 (O_1328,N_24922,N_24901);
or UO_1329 (O_1329,N_24910,N_24881);
xnor UO_1330 (O_1330,N_24910,N_24851);
nand UO_1331 (O_1331,N_24838,N_24954);
and UO_1332 (O_1332,N_24862,N_24836);
nor UO_1333 (O_1333,N_24969,N_24998);
or UO_1334 (O_1334,N_24801,N_24956);
or UO_1335 (O_1335,N_24841,N_24997);
and UO_1336 (O_1336,N_24964,N_24814);
xnor UO_1337 (O_1337,N_24915,N_24916);
or UO_1338 (O_1338,N_24908,N_24984);
nor UO_1339 (O_1339,N_24912,N_24895);
nor UO_1340 (O_1340,N_24972,N_24923);
nand UO_1341 (O_1341,N_24961,N_24959);
nand UO_1342 (O_1342,N_24912,N_24985);
xor UO_1343 (O_1343,N_24928,N_24923);
nand UO_1344 (O_1344,N_24878,N_24932);
nor UO_1345 (O_1345,N_24984,N_24911);
nand UO_1346 (O_1346,N_24841,N_24874);
nor UO_1347 (O_1347,N_24908,N_24992);
xnor UO_1348 (O_1348,N_24825,N_24980);
nor UO_1349 (O_1349,N_24978,N_24808);
or UO_1350 (O_1350,N_24899,N_24835);
and UO_1351 (O_1351,N_24904,N_24933);
nor UO_1352 (O_1352,N_24853,N_24921);
nor UO_1353 (O_1353,N_24923,N_24955);
or UO_1354 (O_1354,N_24981,N_24940);
or UO_1355 (O_1355,N_24829,N_24980);
nand UO_1356 (O_1356,N_24876,N_24857);
or UO_1357 (O_1357,N_24888,N_24988);
nor UO_1358 (O_1358,N_24929,N_24810);
and UO_1359 (O_1359,N_24967,N_24872);
nor UO_1360 (O_1360,N_24804,N_24960);
nor UO_1361 (O_1361,N_24818,N_24890);
and UO_1362 (O_1362,N_24938,N_24972);
nor UO_1363 (O_1363,N_24821,N_24921);
and UO_1364 (O_1364,N_24956,N_24887);
and UO_1365 (O_1365,N_24938,N_24968);
nand UO_1366 (O_1366,N_24806,N_24841);
and UO_1367 (O_1367,N_24960,N_24805);
and UO_1368 (O_1368,N_24917,N_24991);
xor UO_1369 (O_1369,N_24865,N_24882);
nor UO_1370 (O_1370,N_24833,N_24881);
nand UO_1371 (O_1371,N_24800,N_24825);
nor UO_1372 (O_1372,N_24926,N_24827);
nand UO_1373 (O_1373,N_24919,N_24844);
nand UO_1374 (O_1374,N_24973,N_24804);
and UO_1375 (O_1375,N_24888,N_24992);
nand UO_1376 (O_1376,N_24973,N_24846);
xor UO_1377 (O_1377,N_24967,N_24930);
and UO_1378 (O_1378,N_24924,N_24940);
nand UO_1379 (O_1379,N_24815,N_24832);
xor UO_1380 (O_1380,N_24873,N_24888);
xnor UO_1381 (O_1381,N_24803,N_24867);
nor UO_1382 (O_1382,N_24912,N_24976);
nor UO_1383 (O_1383,N_24975,N_24810);
and UO_1384 (O_1384,N_24856,N_24989);
or UO_1385 (O_1385,N_24888,N_24935);
or UO_1386 (O_1386,N_24825,N_24908);
nor UO_1387 (O_1387,N_24873,N_24816);
nor UO_1388 (O_1388,N_24943,N_24960);
nor UO_1389 (O_1389,N_24937,N_24895);
and UO_1390 (O_1390,N_24942,N_24810);
xor UO_1391 (O_1391,N_24853,N_24849);
xor UO_1392 (O_1392,N_24817,N_24960);
nand UO_1393 (O_1393,N_24937,N_24889);
or UO_1394 (O_1394,N_24979,N_24941);
and UO_1395 (O_1395,N_24908,N_24862);
xor UO_1396 (O_1396,N_24947,N_24801);
or UO_1397 (O_1397,N_24868,N_24805);
nor UO_1398 (O_1398,N_24874,N_24967);
nor UO_1399 (O_1399,N_24983,N_24954);
or UO_1400 (O_1400,N_24942,N_24994);
and UO_1401 (O_1401,N_24865,N_24844);
and UO_1402 (O_1402,N_24978,N_24854);
nor UO_1403 (O_1403,N_24846,N_24837);
xor UO_1404 (O_1404,N_24822,N_24920);
nand UO_1405 (O_1405,N_24822,N_24954);
nor UO_1406 (O_1406,N_24900,N_24849);
nand UO_1407 (O_1407,N_24977,N_24891);
xnor UO_1408 (O_1408,N_24975,N_24983);
or UO_1409 (O_1409,N_24889,N_24876);
and UO_1410 (O_1410,N_24828,N_24958);
or UO_1411 (O_1411,N_24986,N_24856);
and UO_1412 (O_1412,N_24975,N_24964);
or UO_1413 (O_1413,N_24924,N_24818);
xnor UO_1414 (O_1414,N_24891,N_24917);
nand UO_1415 (O_1415,N_24958,N_24905);
nand UO_1416 (O_1416,N_24955,N_24990);
or UO_1417 (O_1417,N_24948,N_24833);
or UO_1418 (O_1418,N_24836,N_24849);
and UO_1419 (O_1419,N_24838,N_24955);
nor UO_1420 (O_1420,N_24933,N_24819);
nand UO_1421 (O_1421,N_24917,N_24876);
and UO_1422 (O_1422,N_24978,N_24823);
xnor UO_1423 (O_1423,N_24813,N_24909);
or UO_1424 (O_1424,N_24896,N_24835);
or UO_1425 (O_1425,N_24828,N_24971);
or UO_1426 (O_1426,N_24883,N_24946);
nor UO_1427 (O_1427,N_24992,N_24975);
nor UO_1428 (O_1428,N_24927,N_24945);
xor UO_1429 (O_1429,N_24943,N_24817);
xor UO_1430 (O_1430,N_24870,N_24856);
xnor UO_1431 (O_1431,N_24882,N_24830);
or UO_1432 (O_1432,N_24817,N_24990);
and UO_1433 (O_1433,N_24971,N_24908);
nand UO_1434 (O_1434,N_24963,N_24991);
or UO_1435 (O_1435,N_24994,N_24836);
nand UO_1436 (O_1436,N_24889,N_24920);
or UO_1437 (O_1437,N_24836,N_24871);
or UO_1438 (O_1438,N_24825,N_24829);
and UO_1439 (O_1439,N_24856,N_24861);
nand UO_1440 (O_1440,N_24980,N_24924);
or UO_1441 (O_1441,N_24998,N_24987);
or UO_1442 (O_1442,N_24874,N_24853);
or UO_1443 (O_1443,N_24820,N_24953);
and UO_1444 (O_1444,N_24858,N_24857);
and UO_1445 (O_1445,N_24990,N_24870);
xor UO_1446 (O_1446,N_24917,N_24809);
and UO_1447 (O_1447,N_24923,N_24812);
nor UO_1448 (O_1448,N_24989,N_24949);
and UO_1449 (O_1449,N_24877,N_24901);
and UO_1450 (O_1450,N_24925,N_24894);
nand UO_1451 (O_1451,N_24815,N_24853);
nor UO_1452 (O_1452,N_24971,N_24983);
nor UO_1453 (O_1453,N_24912,N_24894);
xor UO_1454 (O_1454,N_24802,N_24803);
nand UO_1455 (O_1455,N_24901,N_24876);
nor UO_1456 (O_1456,N_24989,N_24859);
or UO_1457 (O_1457,N_24912,N_24905);
or UO_1458 (O_1458,N_24912,N_24862);
nor UO_1459 (O_1459,N_24985,N_24834);
or UO_1460 (O_1460,N_24975,N_24979);
or UO_1461 (O_1461,N_24802,N_24974);
nor UO_1462 (O_1462,N_24924,N_24961);
or UO_1463 (O_1463,N_24814,N_24851);
or UO_1464 (O_1464,N_24847,N_24815);
nand UO_1465 (O_1465,N_24955,N_24993);
xor UO_1466 (O_1466,N_24972,N_24976);
and UO_1467 (O_1467,N_24954,N_24802);
nand UO_1468 (O_1468,N_24969,N_24876);
xnor UO_1469 (O_1469,N_24894,N_24963);
or UO_1470 (O_1470,N_24871,N_24887);
nor UO_1471 (O_1471,N_24945,N_24882);
nor UO_1472 (O_1472,N_24954,N_24916);
or UO_1473 (O_1473,N_24864,N_24845);
xor UO_1474 (O_1474,N_24998,N_24910);
xnor UO_1475 (O_1475,N_24904,N_24941);
or UO_1476 (O_1476,N_24816,N_24992);
xnor UO_1477 (O_1477,N_24953,N_24889);
nor UO_1478 (O_1478,N_24935,N_24889);
and UO_1479 (O_1479,N_24961,N_24889);
xor UO_1480 (O_1480,N_24830,N_24997);
nor UO_1481 (O_1481,N_24975,N_24970);
and UO_1482 (O_1482,N_24882,N_24837);
xnor UO_1483 (O_1483,N_24923,N_24989);
and UO_1484 (O_1484,N_24883,N_24885);
nand UO_1485 (O_1485,N_24816,N_24846);
and UO_1486 (O_1486,N_24958,N_24870);
and UO_1487 (O_1487,N_24821,N_24802);
xnor UO_1488 (O_1488,N_24869,N_24958);
or UO_1489 (O_1489,N_24986,N_24902);
and UO_1490 (O_1490,N_24966,N_24807);
xor UO_1491 (O_1491,N_24857,N_24953);
and UO_1492 (O_1492,N_24918,N_24810);
and UO_1493 (O_1493,N_24933,N_24993);
nor UO_1494 (O_1494,N_24867,N_24840);
nor UO_1495 (O_1495,N_24847,N_24800);
nand UO_1496 (O_1496,N_24982,N_24988);
and UO_1497 (O_1497,N_24894,N_24976);
nor UO_1498 (O_1498,N_24921,N_24864);
or UO_1499 (O_1499,N_24955,N_24879);
or UO_1500 (O_1500,N_24893,N_24996);
or UO_1501 (O_1501,N_24904,N_24912);
nor UO_1502 (O_1502,N_24880,N_24845);
nand UO_1503 (O_1503,N_24859,N_24967);
nor UO_1504 (O_1504,N_24888,N_24898);
nand UO_1505 (O_1505,N_24859,N_24838);
and UO_1506 (O_1506,N_24919,N_24866);
xor UO_1507 (O_1507,N_24898,N_24946);
nand UO_1508 (O_1508,N_24942,N_24910);
and UO_1509 (O_1509,N_24980,N_24955);
and UO_1510 (O_1510,N_24940,N_24824);
nor UO_1511 (O_1511,N_24986,N_24829);
nand UO_1512 (O_1512,N_24914,N_24821);
or UO_1513 (O_1513,N_24882,N_24993);
nor UO_1514 (O_1514,N_24856,N_24819);
nor UO_1515 (O_1515,N_24862,N_24928);
nand UO_1516 (O_1516,N_24982,N_24816);
nand UO_1517 (O_1517,N_24906,N_24821);
nand UO_1518 (O_1518,N_24844,N_24805);
nand UO_1519 (O_1519,N_24946,N_24826);
or UO_1520 (O_1520,N_24978,N_24907);
or UO_1521 (O_1521,N_24909,N_24949);
nor UO_1522 (O_1522,N_24972,N_24826);
nor UO_1523 (O_1523,N_24908,N_24816);
and UO_1524 (O_1524,N_24859,N_24944);
nor UO_1525 (O_1525,N_24926,N_24922);
and UO_1526 (O_1526,N_24996,N_24955);
xnor UO_1527 (O_1527,N_24846,N_24897);
nand UO_1528 (O_1528,N_24853,N_24940);
xnor UO_1529 (O_1529,N_24936,N_24900);
and UO_1530 (O_1530,N_24929,N_24968);
or UO_1531 (O_1531,N_24847,N_24967);
or UO_1532 (O_1532,N_24927,N_24912);
and UO_1533 (O_1533,N_24846,N_24819);
xnor UO_1534 (O_1534,N_24863,N_24803);
xnor UO_1535 (O_1535,N_24937,N_24838);
or UO_1536 (O_1536,N_24823,N_24826);
and UO_1537 (O_1537,N_24829,N_24816);
and UO_1538 (O_1538,N_24911,N_24854);
xnor UO_1539 (O_1539,N_24909,N_24974);
xnor UO_1540 (O_1540,N_24895,N_24929);
xnor UO_1541 (O_1541,N_24972,N_24802);
nor UO_1542 (O_1542,N_24995,N_24982);
xor UO_1543 (O_1543,N_24893,N_24926);
nand UO_1544 (O_1544,N_24916,N_24996);
xor UO_1545 (O_1545,N_24965,N_24957);
or UO_1546 (O_1546,N_24936,N_24935);
xnor UO_1547 (O_1547,N_24969,N_24996);
or UO_1548 (O_1548,N_24902,N_24954);
nand UO_1549 (O_1549,N_24829,N_24926);
and UO_1550 (O_1550,N_24938,N_24882);
xnor UO_1551 (O_1551,N_24905,N_24963);
or UO_1552 (O_1552,N_24994,N_24854);
and UO_1553 (O_1553,N_24982,N_24839);
and UO_1554 (O_1554,N_24816,N_24905);
or UO_1555 (O_1555,N_24926,N_24851);
or UO_1556 (O_1556,N_24873,N_24827);
nor UO_1557 (O_1557,N_24955,N_24857);
nor UO_1558 (O_1558,N_24923,N_24973);
xor UO_1559 (O_1559,N_24892,N_24814);
and UO_1560 (O_1560,N_24931,N_24830);
xor UO_1561 (O_1561,N_24830,N_24843);
nand UO_1562 (O_1562,N_24928,N_24906);
xor UO_1563 (O_1563,N_24937,N_24898);
nor UO_1564 (O_1564,N_24986,N_24876);
and UO_1565 (O_1565,N_24933,N_24907);
xnor UO_1566 (O_1566,N_24971,N_24869);
nand UO_1567 (O_1567,N_24895,N_24981);
nor UO_1568 (O_1568,N_24810,N_24834);
and UO_1569 (O_1569,N_24912,N_24842);
or UO_1570 (O_1570,N_24992,N_24841);
nand UO_1571 (O_1571,N_24926,N_24903);
and UO_1572 (O_1572,N_24925,N_24922);
or UO_1573 (O_1573,N_24945,N_24901);
nand UO_1574 (O_1574,N_24838,N_24862);
xnor UO_1575 (O_1575,N_24949,N_24862);
and UO_1576 (O_1576,N_24972,N_24936);
nand UO_1577 (O_1577,N_24963,N_24882);
xor UO_1578 (O_1578,N_24904,N_24848);
and UO_1579 (O_1579,N_24859,N_24976);
or UO_1580 (O_1580,N_24803,N_24813);
or UO_1581 (O_1581,N_24869,N_24920);
or UO_1582 (O_1582,N_24978,N_24855);
and UO_1583 (O_1583,N_24990,N_24913);
xnor UO_1584 (O_1584,N_24834,N_24848);
and UO_1585 (O_1585,N_24889,N_24968);
or UO_1586 (O_1586,N_24900,N_24810);
and UO_1587 (O_1587,N_24929,N_24988);
and UO_1588 (O_1588,N_24939,N_24853);
xor UO_1589 (O_1589,N_24889,N_24801);
or UO_1590 (O_1590,N_24990,N_24915);
nor UO_1591 (O_1591,N_24857,N_24848);
nor UO_1592 (O_1592,N_24939,N_24828);
nand UO_1593 (O_1593,N_24879,N_24941);
and UO_1594 (O_1594,N_24804,N_24829);
and UO_1595 (O_1595,N_24837,N_24864);
and UO_1596 (O_1596,N_24996,N_24942);
and UO_1597 (O_1597,N_24812,N_24959);
nand UO_1598 (O_1598,N_24962,N_24941);
and UO_1599 (O_1599,N_24941,N_24947);
and UO_1600 (O_1600,N_24928,N_24821);
nand UO_1601 (O_1601,N_24869,N_24977);
xor UO_1602 (O_1602,N_24837,N_24883);
and UO_1603 (O_1603,N_24934,N_24902);
and UO_1604 (O_1604,N_24824,N_24882);
or UO_1605 (O_1605,N_24808,N_24942);
nor UO_1606 (O_1606,N_24803,N_24978);
nor UO_1607 (O_1607,N_24863,N_24903);
xor UO_1608 (O_1608,N_24917,N_24906);
nor UO_1609 (O_1609,N_24966,N_24905);
or UO_1610 (O_1610,N_24971,N_24974);
xnor UO_1611 (O_1611,N_24842,N_24860);
nor UO_1612 (O_1612,N_24914,N_24882);
nor UO_1613 (O_1613,N_24929,N_24928);
and UO_1614 (O_1614,N_24993,N_24949);
and UO_1615 (O_1615,N_24937,N_24918);
or UO_1616 (O_1616,N_24960,N_24982);
nor UO_1617 (O_1617,N_24978,N_24973);
or UO_1618 (O_1618,N_24888,N_24938);
or UO_1619 (O_1619,N_24890,N_24908);
or UO_1620 (O_1620,N_24828,N_24901);
nand UO_1621 (O_1621,N_24841,N_24883);
or UO_1622 (O_1622,N_24954,N_24966);
xor UO_1623 (O_1623,N_24987,N_24807);
and UO_1624 (O_1624,N_24861,N_24963);
and UO_1625 (O_1625,N_24894,N_24880);
xnor UO_1626 (O_1626,N_24903,N_24831);
or UO_1627 (O_1627,N_24974,N_24953);
xor UO_1628 (O_1628,N_24814,N_24832);
or UO_1629 (O_1629,N_24872,N_24914);
and UO_1630 (O_1630,N_24986,N_24950);
nor UO_1631 (O_1631,N_24805,N_24972);
and UO_1632 (O_1632,N_24902,N_24938);
or UO_1633 (O_1633,N_24934,N_24890);
nand UO_1634 (O_1634,N_24850,N_24917);
nor UO_1635 (O_1635,N_24921,N_24900);
xnor UO_1636 (O_1636,N_24907,N_24912);
or UO_1637 (O_1637,N_24925,N_24940);
xor UO_1638 (O_1638,N_24920,N_24811);
or UO_1639 (O_1639,N_24839,N_24802);
xor UO_1640 (O_1640,N_24911,N_24977);
xnor UO_1641 (O_1641,N_24931,N_24932);
or UO_1642 (O_1642,N_24984,N_24974);
nor UO_1643 (O_1643,N_24840,N_24823);
and UO_1644 (O_1644,N_24906,N_24810);
and UO_1645 (O_1645,N_24855,N_24840);
or UO_1646 (O_1646,N_24880,N_24964);
xor UO_1647 (O_1647,N_24858,N_24888);
and UO_1648 (O_1648,N_24984,N_24901);
and UO_1649 (O_1649,N_24870,N_24837);
and UO_1650 (O_1650,N_24873,N_24940);
and UO_1651 (O_1651,N_24872,N_24844);
xnor UO_1652 (O_1652,N_24839,N_24824);
xor UO_1653 (O_1653,N_24843,N_24927);
nand UO_1654 (O_1654,N_24875,N_24909);
nand UO_1655 (O_1655,N_24917,N_24841);
nand UO_1656 (O_1656,N_24832,N_24997);
nor UO_1657 (O_1657,N_24982,N_24851);
and UO_1658 (O_1658,N_24960,N_24905);
xor UO_1659 (O_1659,N_24862,N_24929);
or UO_1660 (O_1660,N_24976,N_24815);
and UO_1661 (O_1661,N_24923,N_24843);
nand UO_1662 (O_1662,N_24894,N_24814);
nor UO_1663 (O_1663,N_24890,N_24904);
nand UO_1664 (O_1664,N_24882,N_24856);
xor UO_1665 (O_1665,N_24866,N_24975);
or UO_1666 (O_1666,N_24898,N_24985);
xnor UO_1667 (O_1667,N_24939,N_24954);
nor UO_1668 (O_1668,N_24943,N_24922);
nand UO_1669 (O_1669,N_24822,N_24827);
nor UO_1670 (O_1670,N_24931,N_24874);
nor UO_1671 (O_1671,N_24911,N_24894);
or UO_1672 (O_1672,N_24930,N_24839);
xnor UO_1673 (O_1673,N_24875,N_24934);
and UO_1674 (O_1674,N_24986,N_24926);
and UO_1675 (O_1675,N_24870,N_24979);
or UO_1676 (O_1676,N_24841,N_24993);
or UO_1677 (O_1677,N_24989,N_24985);
or UO_1678 (O_1678,N_24856,N_24985);
or UO_1679 (O_1679,N_24998,N_24981);
or UO_1680 (O_1680,N_24877,N_24892);
nor UO_1681 (O_1681,N_24966,N_24953);
nand UO_1682 (O_1682,N_24983,N_24991);
and UO_1683 (O_1683,N_24847,N_24987);
xor UO_1684 (O_1684,N_24870,N_24996);
or UO_1685 (O_1685,N_24802,N_24828);
xor UO_1686 (O_1686,N_24905,N_24909);
xor UO_1687 (O_1687,N_24981,N_24990);
nand UO_1688 (O_1688,N_24868,N_24978);
nand UO_1689 (O_1689,N_24899,N_24893);
or UO_1690 (O_1690,N_24906,N_24891);
nor UO_1691 (O_1691,N_24835,N_24976);
and UO_1692 (O_1692,N_24828,N_24874);
nand UO_1693 (O_1693,N_24845,N_24813);
or UO_1694 (O_1694,N_24988,N_24959);
or UO_1695 (O_1695,N_24848,N_24938);
and UO_1696 (O_1696,N_24883,N_24896);
and UO_1697 (O_1697,N_24930,N_24826);
or UO_1698 (O_1698,N_24832,N_24875);
xnor UO_1699 (O_1699,N_24995,N_24954);
and UO_1700 (O_1700,N_24919,N_24984);
xor UO_1701 (O_1701,N_24930,N_24965);
and UO_1702 (O_1702,N_24896,N_24892);
and UO_1703 (O_1703,N_24857,N_24962);
nor UO_1704 (O_1704,N_24954,N_24963);
nor UO_1705 (O_1705,N_24827,N_24843);
nor UO_1706 (O_1706,N_24846,N_24824);
and UO_1707 (O_1707,N_24907,N_24923);
nor UO_1708 (O_1708,N_24850,N_24847);
or UO_1709 (O_1709,N_24830,N_24894);
xnor UO_1710 (O_1710,N_24807,N_24958);
xor UO_1711 (O_1711,N_24913,N_24955);
or UO_1712 (O_1712,N_24982,N_24932);
nor UO_1713 (O_1713,N_24850,N_24925);
xor UO_1714 (O_1714,N_24857,N_24870);
nand UO_1715 (O_1715,N_24858,N_24873);
nand UO_1716 (O_1716,N_24890,N_24925);
or UO_1717 (O_1717,N_24942,N_24891);
or UO_1718 (O_1718,N_24958,N_24959);
nand UO_1719 (O_1719,N_24896,N_24931);
nand UO_1720 (O_1720,N_24810,N_24821);
and UO_1721 (O_1721,N_24935,N_24838);
and UO_1722 (O_1722,N_24829,N_24967);
or UO_1723 (O_1723,N_24957,N_24801);
xor UO_1724 (O_1724,N_24909,N_24946);
nor UO_1725 (O_1725,N_24800,N_24902);
and UO_1726 (O_1726,N_24907,N_24858);
xnor UO_1727 (O_1727,N_24850,N_24995);
and UO_1728 (O_1728,N_24819,N_24972);
nor UO_1729 (O_1729,N_24981,N_24965);
nor UO_1730 (O_1730,N_24858,N_24921);
xnor UO_1731 (O_1731,N_24823,N_24853);
xnor UO_1732 (O_1732,N_24847,N_24812);
or UO_1733 (O_1733,N_24801,N_24952);
or UO_1734 (O_1734,N_24820,N_24980);
and UO_1735 (O_1735,N_24969,N_24982);
nor UO_1736 (O_1736,N_24993,N_24831);
or UO_1737 (O_1737,N_24915,N_24843);
or UO_1738 (O_1738,N_24837,N_24875);
or UO_1739 (O_1739,N_24878,N_24831);
nor UO_1740 (O_1740,N_24853,N_24857);
and UO_1741 (O_1741,N_24920,N_24907);
and UO_1742 (O_1742,N_24939,N_24873);
nor UO_1743 (O_1743,N_24966,N_24982);
xor UO_1744 (O_1744,N_24893,N_24816);
nand UO_1745 (O_1745,N_24863,N_24867);
nand UO_1746 (O_1746,N_24888,N_24893);
xnor UO_1747 (O_1747,N_24884,N_24894);
xor UO_1748 (O_1748,N_24836,N_24838);
nand UO_1749 (O_1749,N_24933,N_24869);
xor UO_1750 (O_1750,N_24981,N_24822);
xnor UO_1751 (O_1751,N_24921,N_24927);
and UO_1752 (O_1752,N_24979,N_24912);
xor UO_1753 (O_1753,N_24908,N_24991);
xor UO_1754 (O_1754,N_24835,N_24951);
nand UO_1755 (O_1755,N_24968,N_24912);
nand UO_1756 (O_1756,N_24864,N_24919);
nand UO_1757 (O_1757,N_24953,N_24928);
xor UO_1758 (O_1758,N_24878,N_24835);
or UO_1759 (O_1759,N_24874,N_24949);
nor UO_1760 (O_1760,N_24845,N_24950);
nor UO_1761 (O_1761,N_24884,N_24958);
nor UO_1762 (O_1762,N_24857,N_24944);
xnor UO_1763 (O_1763,N_24974,N_24923);
nor UO_1764 (O_1764,N_24932,N_24926);
nor UO_1765 (O_1765,N_24965,N_24851);
or UO_1766 (O_1766,N_24856,N_24952);
and UO_1767 (O_1767,N_24872,N_24909);
nor UO_1768 (O_1768,N_24924,N_24849);
nor UO_1769 (O_1769,N_24923,N_24878);
and UO_1770 (O_1770,N_24995,N_24803);
and UO_1771 (O_1771,N_24951,N_24963);
nand UO_1772 (O_1772,N_24905,N_24914);
xor UO_1773 (O_1773,N_24856,N_24974);
nor UO_1774 (O_1774,N_24975,N_24859);
nor UO_1775 (O_1775,N_24991,N_24889);
or UO_1776 (O_1776,N_24958,N_24844);
nand UO_1777 (O_1777,N_24984,N_24829);
and UO_1778 (O_1778,N_24883,N_24893);
nand UO_1779 (O_1779,N_24974,N_24844);
nand UO_1780 (O_1780,N_24927,N_24872);
nand UO_1781 (O_1781,N_24931,N_24934);
or UO_1782 (O_1782,N_24916,N_24822);
and UO_1783 (O_1783,N_24902,N_24952);
nor UO_1784 (O_1784,N_24936,N_24980);
nand UO_1785 (O_1785,N_24914,N_24932);
or UO_1786 (O_1786,N_24836,N_24903);
nor UO_1787 (O_1787,N_24928,N_24960);
xnor UO_1788 (O_1788,N_24938,N_24821);
xor UO_1789 (O_1789,N_24839,N_24854);
xor UO_1790 (O_1790,N_24865,N_24894);
and UO_1791 (O_1791,N_24885,N_24982);
xor UO_1792 (O_1792,N_24829,N_24942);
and UO_1793 (O_1793,N_24909,N_24932);
nand UO_1794 (O_1794,N_24883,N_24967);
nor UO_1795 (O_1795,N_24956,N_24848);
nor UO_1796 (O_1796,N_24928,N_24852);
nand UO_1797 (O_1797,N_24838,N_24844);
and UO_1798 (O_1798,N_24833,N_24987);
or UO_1799 (O_1799,N_24920,N_24888);
and UO_1800 (O_1800,N_24859,N_24864);
xor UO_1801 (O_1801,N_24983,N_24814);
xnor UO_1802 (O_1802,N_24975,N_24942);
nand UO_1803 (O_1803,N_24939,N_24925);
nor UO_1804 (O_1804,N_24863,N_24810);
nor UO_1805 (O_1805,N_24895,N_24911);
and UO_1806 (O_1806,N_24913,N_24958);
nand UO_1807 (O_1807,N_24992,N_24877);
and UO_1808 (O_1808,N_24942,N_24805);
and UO_1809 (O_1809,N_24804,N_24971);
nor UO_1810 (O_1810,N_24935,N_24932);
or UO_1811 (O_1811,N_24861,N_24935);
and UO_1812 (O_1812,N_24967,N_24895);
nand UO_1813 (O_1813,N_24833,N_24810);
xor UO_1814 (O_1814,N_24926,N_24860);
nor UO_1815 (O_1815,N_24901,N_24917);
nand UO_1816 (O_1816,N_24948,N_24964);
or UO_1817 (O_1817,N_24876,N_24830);
or UO_1818 (O_1818,N_24922,N_24944);
and UO_1819 (O_1819,N_24927,N_24871);
or UO_1820 (O_1820,N_24929,N_24907);
nor UO_1821 (O_1821,N_24896,N_24967);
xnor UO_1822 (O_1822,N_24919,N_24942);
and UO_1823 (O_1823,N_24870,N_24884);
nor UO_1824 (O_1824,N_24944,N_24976);
and UO_1825 (O_1825,N_24979,N_24904);
and UO_1826 (O_1826,N_24828,N_24934);
nor UO_1827 (O_1827,N_24938,N_24854);
and UO_1828 (O_1828,N_24826,N_24982);
xor UO_1829 (O_1829,N_24972,N_24969);
nand UO_1830 (O_1830,N_24807,N_24886);
xnor UO_1831 (O_1831,N_24916,N_24933);
and UO_1832 (O_1832,N_24928,N_24836);
or UO_1833 (O_1833,N_24849,N_24960);
xnor UO_1834 (O_1834,N_24829,N_24826);
or UO_1835 (O_1835,N_24852,N_24872);
xor UO_1836 (O_1836,N_24829,N_24920);
or UO_1837 (O_1837,N_24989,N_24806);
and UO_1838 (O_1838,N_24823,N_24930);
nand UO_1839 (O_1839,N_24972,N_24988);
xor UO_1840 (O_1840,N_24865,N_24982);
and UO_1841 (O_1841,N_24902,N_24823);
nor UO_1842 (O_1842,N_24882,N_24828);
nor UO_1843 (O_1843,N_24984,N_24899);
or UO_1844 (O_1844,N_24870,N_24967);
xor UO_1845 (O_1845,N_24810,N_24985);
nor UO_1846 (O_1846,N_24900,N_24870);
nand UO_1847 (O_1847,N_24977,N_24975);
nor UO_1848 (O_1848,N_24940,N_24875);
nand UO_1849 (O_1849,N_24821,N_24812);
xor UO_1850 (O_1850,N_24997,N_24893);
nor UO_1851 (O_1851,N_24993,N_24948);
xnor UO_1852 (O_1852,N_24849,N_24912);
nor UO_1853 (O_1853,N_24920,N_24970);
or UO_1854 (O_1854,N_24819,N_24826);
and UO_1855 (O_1855,N_24920,N_24813);
nand UO_1856 (O_1856,N_24900,N_24867);
xor UO_1857 (O_1857,N_24908,N_24811);
xnor UO_1858 (O_1858,N_24809,N_24993);
xor UO_1859 (O_1859,N_24971,N_24856);
xor UO_1860 (O_1860,N_24902,N_24955);
nand UO_1861 (O_1861,N_24898,N_24995);
or UO_1862 (O_1862,N_24952,N_24803);
nor UO_1863 (O_1863,N_24990,N_24923);
and UO_1864 (O_1864,N_24868,N_24965);
xnor UO_1865 (O_1865,N_24932,N_24801);
nand UO_1866 (O_1866,N_24912,N_24911);
nand UO_1867 (O_1867,N_24837,N_24908);
and UO_1868 (O_1868,N_24822,N_24989);
or UO_1869 (O_1869,N_24857,N_24824);
nand UO_1870 (O_1870,N_24836,N_24839);
nand UO_1871 (O_1871,N_24981,N_24941);
nor UO_1872 (O_1872,N_24831,N_24810);
xor UO_1873 (O_1873,N_24995,N_24994);
nor UO_1874 (O_1874,N_24998,N_24845);
xor UO_1875 (O_1875,N_24955,N_24806);
and UO_1876 (O_1876,N_24942,N_24981);
nand UO_1877 (O_1877,N_24898,N_24803);
nor UO_1878 (O_1878,N_24911,N_24914);
or UO_1879 (O_1879,N_24909,N_24987);
nor UO_1880 (O_1880,N_24904,N_24971);
and UO_1881 (O_1881,N_24928,N_24801);
and UO_1882 (O_1882,N_24927,N_24962);
nand UO_1883 (O_1883,N_24993,N_24905);
nor UO_1884 (O_1884,N_24805,N_24912);
xor UO_1885 (O_1885,N_24803,N_24894);
nor UO_1886 (O_1886,N_24907,N_24991);
and UO_1887 (O_1887,N_24818,N_24814);
or UO_1888 (O_1888,N_24904,N_24872);
nor UO_1889 (O_1889,N_24842,N_24852);
and UO_1890 (O_1890,N_24959,N_24826);
nand UO_1891 (O_1891,N_24812,N_24879);
or UO_1892 (O_1892,N_24865,N_24834);
or UO_1893 (O_1893,N_24919,N_24812);
or UO_1894 (O_1894,N_24962,N_24866);
and UO_1895 (O_1895,N_24975,N_24889);
xnor UO_1896 (O_1896,N_24866,N_24821);
and UO_1897 (O_1897,N_24982,N_24829);
xor UO_1898 (O_1898,N_24808,N_24952);
nand UO_1899 (O_1899,N_24811,N_24828);
nor UO_1900 (O_1900,N_24859,N_24951);
nor UO_1901 (O_1901,N_24870,N_24841);
nand UO_1902 (O_1902,N_24982,N_24849);
nand UO_1903 (O_1903,N_24905,N_24945);
or UO_1904 (O_1904,N_24934,N_24858);
and UO_1905 (O_1905,N_24841,N_24852);
nor UO_1906 (O_1906,N_24887,N_24872);
and UO_1907 (O_1907,N_24927,N_24820);
or UO_1908 (O_1908,N_24987,N_24980);
nor UO_1909 (O_1909,N_24914,N_24970);
and UO_1910 (O_1910,N_24815,N_24965);
nor UO_1911 (O_1911,N_24869,N_24915);
xnor UO_1912 (O_1912,N_24819,N_24832);
nand UO_1913 (O_1913,N_24808,N_24907);
nand UO_1914 (O_1914,N_24899,N_24913);
and UO_1915 (O_1915,N_24993,N_24927);
nor UO_1916 (O_1916,N_24822,N_24825);
nand UO_1917 (O_1917,N_24827,N_24832);
xor UO_1918 (O_1918,N_24957,N_24969);
nor UO_1919 (O_1919,N_24950,N_24835);
xor UO_1920 (O_1920,N_24917,N_24993);
and UO_1921 (O_1921,N_24841,N_24846);
nand UO_1922 (O_1922,N_24991,N_24845);
or UO_1923 (O_1923,N_24915,N_24954);
and UO_1924 (O_1924,N_24809,N_24883);
xor UO_1925 (O_1925,N_24907,N_24898);
nand UO_1926 (O_1926,N_24808,N_24920);
xor UO_1927 (O_1927,N_24998,N_24809);
xnor UO_1928 (O_1928,N_24842,N_24876);
and UO_1929 (O_1929,N_24805,N_24935);
and UO_1930 (O_1930,N_24856,N_24824);
and UO_1931 (O_1931,N_24900,N_24892);
xor UO_1932 (O_1932,N_24841,N_24911);
or UO_1933 (O_1933,N_24869,N_24936);
nor UO_1934 (O_1934,N_24918,N_24805);
nand UO_1935 (O_1935,N_24937,N_24834);
or UO_1936 (O_1936,N_24802,N_24929);
xor UO_1937 (O_1937,N_24955,N_24967);
nor UO_1938 (O_1938,N_24812,N_24908);
nor UO_1939 (O_1939,N_24878,N_24889);
nand UO_1940 (O_1940,N_24921,N_24901);
xor UO_1941 (O_1941,N_24852,N_24912);
nor UO_1942 (O_1942,N_24904,N_24845);
xnor UO_1943 (O_1943,N_24917,N_24903);
nor UO_1944 (O_1944,N_24964,N_24974);
nor UO_1945 (O_1945,N_24920,N_24908);
or UO_1946 (O_1946,N_24896,N_24984);
nand UO_1947 (O_1947,N_24893,N_24998);
nand UO_1948 (O_1948,N_24966,N_24802);
or UO_1949 (O_1949,N_24998,N_24833);
nor UO_1950 (O_1950,N_24862,N_24806);
nand UO_1951 (O_1951,N_24930,N_24828);
or UO_1952 (O_1952,N_24956,N_24918);
and UO_1953 (O_1953,N_24866,N_24989);
nand UO_1954 (O_1954,N_24862,N_24819);
and UO_1955 (O_1955,N_24865,N_24885);
and UO_1956 (O_1956,N_24821,N_24978);
xnor UO_1957 (O_1957,N_24877,N_24881);
nand UO_1958 (O_1958,N_24914,N_24857);
and UO_1959 (O_1959,N_24885,N_24802);
nand UO_1960 (O_1960,N_24991,N_24951);
and UO_1961 (O_1961,N_24965,N_24946);
nor UO_1962 (O_1962,N_24989,N_24800);
xor UO_1963 (O_1963,N_24865,N_24965);
and UO_1964 (O_1964,N_24879,N_24895);
nor UO_1965 (O_1965,N_24934,N_24976);
or UO_1966 (O_1966,N_24816,N_24986);
xor UO_1967 (O_1967,N_24893,N_24978);
nor UO_1968 (O_1968,N_24815,N_24895);
xnor UO_1969 (O_1969,N_24802,N_24932);
nor UO_1970 (O_1970,N_24844,N_24869);
or UO_1971 (O_1971,N_24939,N_24936);
xor UO_1972 (O_1972,N_24848,N_24908);
and UO_1973 (O_1973,N_24845,N_24980);
or UO_1974 (O_1974,N_24921,N_24861);
xor UO_1975 (O_1975,N_24923,N_24985);
and UO_1976 (O_1976,N_24863,N_24977);
nand UO_1977 (O_1977,N_24947,N_24916);
and UO_1978 (O_1978,N_24811,N_24802);
nor UO_1979 (O_1979,N_24831,N_24859);
nand UO_1980 (O_1980,N_24874,N_24893);
nor UO_1981 (O_1981,N_24822,N_24875);
or UO_1982 (O_1982,N_24869,N_24959);
xnor UO_1983 (O_1983,N_24852,N_24814);
and UO_1984 (O_1984,N_24943,N_24997);
xnor UO_1985 (O_1985,N_24806,N_24881);
nor UO_1986 (O_1986,N_24891,N_24997);
xor UO_1987 (O_1987,N_24885,N_24976);
xor UO_1988 (O_1988,N_24831,N_24882);
xnor UO_1989 (O_1989,N_24880,N_24942);
or UO_1990 (O_1990,N_24998,N_24805);
or UO_1991 (O_1991,N_24896,N_24989);
nand UO_1992 (O_1992,N_24842,N_24922);
or UO_1993 (O_1993,N_24959,N_24982);
and UO_1994 (O_1994,N_24874,N_24903);
nand UO_1995 (O_1995,N_24813,N_24980);
or UO_1996 (O_1996,N_24895,N_24812);
xor UO_1997 (O_1997,N_24988,N_24917);
xnor UO_1998 (O_1998,N_24982,N_24974);
and UO_1999 (O_1999,N_24931,N_24899);
nor UO_2000 (O_2000,N_24934,N_24900);
nand UO_2001 (O_2001,N_24806,N_24947);
or UO_2002 (O_2002,N_24871,N_24949);
and UO_2003 (O_2003,N_24832,N_24854);
xor UO_2004 (O_2004,N_24907,N_24880);
or UO_2005 (O_2005,N_24961,N_24957);
xor UO_2006 (O_2006,N_24933,N_24935);
or UO_2007 (O_2007,N_24938,N_24981);
nand UO_2008 (O_2008,N_24994,N_24849);
or UO_2009 (O_2009,N_24993,N_24869);
nand UO_2010 (O_2010,N_24802,N_24898);
nor UO_2011 (O_2011,N_24935,N_24860);
nor UO_2012 (O_2012,N_24809,N_24927);
or UO_2013 (O_2013,N_24996,N_24904);
nand UO_2014 (O_2014,N_24918,N_24970);
nor UO_2015 (O_2015,N_24970,N_24926);
nand UO_2016 (O_2016,N_24870,N_24899);
nand UO_2017 (O_2017,N_24979,N_24895);
or UO_2018 (O_2018,N_24829,N_24860);
nand UO_2019 (O_2019,N_24843,N_24907);
nor UO_2020 (O_2020,N_24953,N_24930);
nor UO_2021 (O_2021,N_24883,N_24915);
nor UO_2022 (O_2022,N_24988,N_24823);
nand UO_2023 (O_2023,N_24804,N_24947);
xor UO_2024 (O_2024,N_24807,N_24872);
nand UO_2025 (O_2025,N_24822,N_24983);
xnor UO_2026 (O_2026,N_24921,N_24842);
or UO_2027 (O_2027,N_24992,N_24931);
and UO_2028 (O_2028,N_24826,N_24847);
xnor UO_2029 (O_2029,N_24834,N_24806);
nand UO_2030 (O_2030,N_24856,N_24842);
nand UO_2031 (O_2031,N_24973,N_24943);
xnor UO_2032 (O_2032,N_24845,N_24890);
xnor UO_2033 (O_2033,N_24981,N_24957);
xor UO_2034 (O_2034,N_24871,N_24824);
or UO_2035 (O_2035,N_24897,N_24968);
or UO_2036 (O_2036,N_24809,N_24804);
nand UO_2037 (O_2037,N_24907,N_24805);
or UO_2038 (O_2038,N_24914,N_24823);
and UO_2039 (O_2039,N_24860,N_24921);
and UO_2040 (O_2040,N_24821,N_24801);
xor UO_2041 (O_2041,N_24852,N_24922);
nand UO_2042 (O_2042,N_24944,N_24847);
nor UO_2043 (O_2043,N_24962,N_24993);
xnor UO_2044 (O_2044,N_24967,N_24842);
nand UO_2045 (O_2045,N_24970,N_24909);
nor UO_2046 (O_2046,N_24897,N_24956);
xnor UO_2047 (O_2047,N_24981,N_24857);
and UO_2048 (O_2048,N_24809,N_24897);
and UO_2049 (O_2049,N_24915,N_24908);
nor UO_2050 (O_2050,N_24905,N_24959);
nand UO_2051 (O_2051,N_24994,N_24875);
and UO_2052 (O_2052,N_24985,N_24984);
xor UO_2053 (O_2053,N_24821,N_24813);
nand UO_2054 (O_2054,N_24957,N_24822);
or UO_2055 (O_2055,N_24912,N_24803);
nand UO_2056 (O_2056,N_24881,N_24822);
nand UO_2057 (O_2057,N_24821,N_24814);
nor UO_2058 (O_2058,N_24978,N_24990);
or UO_2059 (O_2059,N_24862,N_24956);
and UO_2060 (O_2060,N_24855,N_24860);
xnor UO_2061 (O_2061,N_24823,N_24820);
nor UO_2062 (O_2062,N_24894,N_24970);
xnor UO_2063 (O_2063,N_24841,N_24949);
and UO_2064 (O_2064,N_24836,N_24963);
nand UO_2065 (O_2065,N_24864,N_24866);
and UO_2066 (O_2066,N_24842,N_24880);
xnor UO_2067 (O_2067,N_24850,N_24947);
and UO_2068 (O_2068,N_24802,N_24814);
and UO_2069 (O_2069,N_24921,N_24953);
or UO_2070 (O_2070,N_24876,N_24924);
nor UO_2071 (O_2071,N_24991,N_24862);
nand UO_2072 (O_2072,N_24982,N_24904);
and UO_2073 (O_2073,N_24937,N_24883);
nand UO_2074 (O_2074,N_24843,N_24983);
nand UO_2075 (O_2075,N_24985,N_24815);
nor UO_2076 (O_2076,N_24866,N_24932);
xor UO_2077 (O_2077,N_24893,N_24921);
or UO_2078 (O_2078,N_24860,N_24979);
or UO_2079 (O_2079,N_24948,N_24879);
nand UO_2080 (O_2080,N_24873,N_24904);
and UO_2081 (O_2081,N_24868,N_24972);
and UO_2082 (O_2082,N_24891,N_24995);
nor UO_2083 (O_2083,N_24910,N_24939);
or UO_2084 (O_2084,N_24828,N_24980);
nor UO_2085 (O_2085,N_24938,N_24857);
and UO_2086 (O_2086,N_24958,N_24813);
or UO_2087 (O_2087,N_24928,N_24991);
xnor UO_2088 (O_2088,N_24950,N_24935);
or UO_2089 (O_2089,N_24910,N_24917);
and UO_2090 (O_2090,N_24872,N_24977);
xor UO_2091 (O_2091,N_24853,N_24916);
nor UO_2092 (O_2092,N_24816,N_24918);
nand UO_2093 (O_2093,N_24888,N_24865);
and UO_2094 (O_2094,N_24968,N_24873);
nor UO_2095 (O_2095,N_24811,N_24999);
xnor UO_2096 (O_2096,N_24940,N_24946);
or UO_2097 (O_2097,N_24880,N_24803);
and UO_2098 (O_2098,N_24986,N_24813);
nor UO_2099 (O_2099,N_24905,N_24964);
xnor UO_2100 (O_2100,N_24957,N_24800);
xnor UO_2101 (O_2101,N_24882,N_24912);
xnor UO_2102 (O_2102,N_24900,N_24841);
xnor UO_2103 (O_2103,N_24942,N_24941);
nand UO_2104 (O_2104,N_24808,N_24992);
nor UO_2105 (O_2105,N_24846,N_24902);
xnor UO_2106 (O_2106,N_24915,N_24886);
nor UO_2107 (O_2107,N_24966,N_24885);
nand UO_2108 (O_2108,N_24897,N_24977);
xor UO_2109 (O_2109,N_24804,N_24924);
nor UO_2110 (O_2110,N_24803,N_24906);
and UO_2111 (O_2111,N_24979,N_24991);
nand UO_2112 (O_2112,N_24845,N_24900);
or UO_2113 (O_2113,N_24937,N_24854);
nand UO_2114 (O_2114,N_24811,N_24870);
and UO_2115 (O_2115,N_24820,N_24932);
xor UO_2116 (O_2116,N_24938,N_24830);
xor UO_2117 (O_2117,N_24956,N_24966);
and UO_2118 (O_2118,N_24951,N_24911);
xnor UO_2119 (O_2119,N_24991,N_24870);
or UO_2120 (O_2120,N_24955,N_24919);
or UO_2121 (O_2121,N_24947,N_24970);
nand UO_2122 (O_2122,N_24885,N_24884);
or UO_2123 (O_2123,N_24869,N_24951);
and UO_2124 (O_2124,N_24824,N_24837);
nand UO_2125 (O_2125,N_24863,N_24812);
nand UO_2126 (O_2126,N_24915,N_24857);
nand UO_2127 (O_2127,N_24983,N_24802);
nor UO_2128 (O_2128,N_24851,N_24930);
nand UO_2129 (O_2129,N_24979,N_24928);
and UO_2130 (O_2130,N_24930,N_24923);
xnor UO_2131 (O_2131,N_24983,N_24896);
nand UO_2132 (O_2132,N_24821,N_24878);
or UO_2133 (O_2133,N_24829,N_24849);
nor UO_2134 (O_2134,N_24873,N_24977);
nand UO_2135 (O_2135,N_24974,N_24865);
xor UO_2136 (O_2136,N_24958,N_24952);
and UO_2137 (O_2137,N_24994,N_24928);
nor UO_2138 (O_2138,N_24947,N_24982);
and UO_2139 (O_2139,N_24816,N_24899);
and UO_2140 (O_2140,N_24927,N_24815);
xor UO_2141 (O_2141,N_24923,N_24810);
and UO_2142 (O_2142,N_24842,N_24819);
xor UO_2143 (O_2143,N_24869,N_24966);
nand UO_2144 (O_2144,N_24891,N_24864);
nand UO_2145 (O_2145,N_24809,N_24888);
xnor UO_2146 (O_2146,N_24943,N_24979);
nand UO_2147 (O_2147,N_24943,N_24952);
or UO_2148 (O_2148,N_24927,N_24943);
xor UO_2149 (O_2149,N_24960,N_24927);
nand UO_2150 (O_2150,N_24936,N_24977);
or UO_2151 (O_2151,N_24962,N_24934);
xor UO_2152 (O_2152,N_24925,N_24854);
xor UO_2153 (O_2153,N_24908,N_24826);
xor UO_2154 (O_2154,N_24930,N_24958);
or UO_2155 (O_2155,N_24817,N_24872);
nor UO_2156 (O_2156,N_24905,N_24904);
nand UO_2157 (O_2157,N_24843,N_24914);
and UO_2158 (O_2158,N_24959,N_24861);
xor UO_2159 (O_2159,N_24885,N_24900);
nand UO_2160 (O_2160,N_24987,N_24816);
nand UO_2161 (O_2161,N_24814,N_24879);
xnor UO_2162 (O_2162,N_24809,N_24832);
nor UO_2163 (O_2163,N_24812,N_24889);
nand UO_2164 (O_2164,N_24808,N_24897);
xor UO_2165 (O_2165,N_24858,N_24816);
xor UO_2166 (O_2166,N_24992,N_24940);
and UO_2167 (O_2167,N_24802,N_24900);
or UO_2168 (O_2168,N_24938,N_24937);
nand UO_2169 (O_2169,N_24915,N_24999);
and UO_2170 (O_2170,N_24858,N_24987);
or UO_2171 (O_2171,N_24889,N_24966);
or UO_2172 (O_2172,N_24810,N_24916);
xnor UO_2173 (O_2173,N_24911,N_24856);
or UO_2174 (O_2174,N_24878,N_24929);
xor UO_2175 (O_2175,N_24989,N_24860);
xnor UO_2176 (O_2176,N_24832,N_24934);
or UO_2177 (O_2177,N_24882,N_24964);
or UO_2178 (O_2178,N_24951,N_24879);
xnor UO_2179 (O_2179,N_24978,N_24832);
xor UO_2180 (O_2180,N_24920,N_24817);
nor UO_2181 (O_2181,N_24988,N_24904);
nor UO_2182 (O_2182,N_24920,N_24864);
and UO_2183 (O_2183,N_24998,N_24966);
and UO_2184 (O_2184,N_24822,N_24913);
and UO_2185 (O_2185,N_24928,N_24941);
and UO_2186 (O_2186,N_24979,N_24966);
nor UO_2187 (O_2187,N_24979,N_24869);
and UO_2188 (O_2188,N_24996,N_24932);
nand UO_2189 (O_2189,N_24990,N_24940);
or UO_2190 (O_2190,N_24963,N_24832);
nand UO_2191 (O_2191,N_24889,N_24960);
nor UO_2192 (O_2192,N_24811,N_24967);
and UO_2193 (O_2193,N_24934,N_24865);
nand UO_2194 (O_2194,N_24853,N_24800);
nand UO_2195 (O_2195,N_24896,N_24894);
nand UO_2196 (O_2196,N_24917,N_24892);
nand UO_2197 (O_2197,N_24866,N_24944);
and UO_2198 (O_2198,N_24928,N_24874);
and UO_2199 (O_2199,N_24899,N_24865);
nor UO_2200 (O_2200,N_24869,N_24910);
xnor UO_2201 (O_2201,N_24847,N_24912);
and UO_2202 (O_2202,N_24961,N_24980);
nand UO_2203 (O_2203,N_24936,N_24966);
nor UO_2204 (O_2204,N_24977,N_24971);
and UO_2205 (O_2205,N_24900,N_24973);
and UO_2206 (O_2206,N_24834,N_24827);
nor UO_2207 (O_2207,N_24910,N_24827);
nand UO_2208 (O_2208,N_24986,N_24842);
nand UO_2209 (O_2209,N_24838,N_24884);
nor UO_2210 (O_2210,N_24869,N_24935);
xor UO_2211 (O_2211,N_24954,N_24938);
xor UO_2212 (O_2212,N_24981,N_24936);
and UO_2213 (O_2213,N_24807,N_24910);
and UO_2214 (O_2214,N_24939,N_24908);
or UO_2215 (O_2215,N_24862,N_24918);
nor UO_2216 (O_2216,N_24959,N_24964);
or UO_2217 (O_2217,N_24863,N_24949);
nor UO_2218 (O_2218,N_24987,N_24925);
nor UO_2219 (O_2219,N_24868,N_24896);
and UO_2220 (O_2220,N_24971,N_24991);
xnor UO_2221 (O_2221,N_24823,N_24922);
and UO_2222 (O_2222,N_24932,N_24981);
xor UO_2223 (O_2223,N_24926,N_24878);
nor UO_2224 (O_2224,N_24894,N_24834);
and UO_2225 (O_2225,N_24837,N_24929);
or UO_2226 (O_2226,N_24953,N_24852);
and UO_2227 (O_2227,N_24880,N_24862);
or UO_2228 (O_2228,N_24820,N_24832);
nand UO_2229 (O_2229,N_24950,N_24919);
xor UO_2230 (O_2230,N_24868,N_24939);
nand UO_2231 (O_2231,N_24848,N_24907);
nor UO_2232 (O_2232,N_24987,N_24961);
and UO_2233 (O_2233,N_24961,N_24939);
xor UO_2234 (O_2234,N_24933,N_24948);
nor UO_2235 (O_2235,N_24951,N_24801);
xor UO_2236 (O_2236,N_24952,N_24881);
nand UO_2237 (O_2237,N_24990,N_24806);
nor UO_2238 (O_2238,N_24904,N_24976);
or UO_2239 (O_2239,N_24856,N_24906);
xor UO_2240 (O_2240,N_24960,N_24978);
and UO_2241 (O_2241,N_24902,N_24895);
or UO_2242 (O_2242,N_24875,N_24936);
and UO_2243 (O_2243,N_24879,N_24976);
and UO_2244 (O_2244,N_24875,N_24968);
or UO_2245 (O_2245,N_24827,N_24811);
nor UO_2246 (O_2246,N_24880,N_24835);
xor UO_2247 (O_2247,N_24831,N_24805);
xor UO_2248 (O_2248,N_24874,N_24981);
nand UO_2249 (O_2249,N_24979,N_24931);
xnor UO_2250 (O_2250,N_24924,N_24822);
and UO_2251 (O_2251,N_24943,N_24901);
nor UO_2252 (O_2252,N_24827,N_24957);
and UO_2253 (O_2253,N_24886,N_24936);
and UO_2254 (O_2254,N_24846,N_24951);
nor UO_2255 (O_2255,N_24942,N_24878);
and UO_2256 (O_2256,N_24997,N_24864);
and UO_2257 (O_2257,N_24977,N_24996);
or UO_2258 (O_2258,N_24913,N_24868);
xnor UO_2259 (O_2259,N_24804,N_24889);
xnor UO_2260 (O_2260,N_24804,N_24923);
nor UO_2261 (O_2261,N_24815,N_24848);
or UO_2262 (O_2262,N_24953,N_24924);
xnor UO_2263 (O_2263,N_24888,N_24895);
xor UO_2264 (O_2264,N_24843,N_24832);
or UO_2265 (O_2265,N_24893,N_24993);
nor UO_2266 (O_2266,N_24944,N_24931);
and UO_2267 (O_2267,N_24993,N_24894);
nand UO_2268 (O_2268,N_24827,N_24998);
nor UO_2269 (O_2269,N_24888,N_24883);
nor UO_2270 (O_2270,N_24844,N_24839);
nand UO_2271 (O_2271,N_24994,N_24809);
xnor UO_2272 (O_2272,N_24961,N_24849);
nand UO_2273 (O_2273,N_24896,N_24853);
xor UO_2274 (O_2274,N_24882,N_24835);
nand UO_2275 (O_2275,N_24890,N_24910);
xnor UO_2276 (O_2276,N_24911,N_24936);
nor UO_2277 (O_2277,N_24935,N_24891);
nor UO_2278 (O_2278,N_24911,N_24996);
nor UO_2279 (O_2279,N_24939,N_24826);
and UO_2280 (O_2280,N_24949,N_24887);
xnor UO_2281 (O_2281,N_24993,N_24930);
or UO_2282 (O_2282,N_24962,N_24888);
nor UO_2283 (O_2283,N_24975,N_24856);
or UO_2284 (O_2284,N_24870,N_24827);
xor UO_2285 (O_2285,N_24811,N_24928);
and UO_2286 (O_2286,N_24925,N_24826);
or UO_2287 (O_2287,N_24962,N_24994);
or UO_2288 (O_2288,N_24839,N_24999);
or UO_2289 (O_2289,N_24861,N_24885);
or UO_2290 (O_2290,N_24938,N_24823);
nand UO_2291 (O_2291,N_24966,N_24835);
nor UO_2292 (O_2292,N_24883,N_24856);
xnor UO_2293 (O_2293,N_24919,N_24898);
nor UO_2294 (O_2294,N_24901,N_24987);
nand UO_2295 (O_2295,N_24847,N_24958);
and UO_2296 (O_2296,N_24954,N_24898);
or UO_2297 (O_2297,N_24937,N_24879);
nor UO_2298 (O_2298,N_24862,N_24812);
or UO_2299 (O_2299,N_24904,N_24824);
or UO_2300 (O_2300,N_24987,N_24966);
and UO_2301 (O_2301,N_24935,N_24911);
xnor UO_2302 (O_2302,N_24879,N_24807);
and UO_2303 (O_2303,N_24948,N_24860);
or UO_2304 (O_2304,N_24914,N_24937);
xor UO_2305 (O_2305,N_24913,N_24887);
xnor UO_2306 (O_2306,N_24815,N_24997);
or UO_2307 (O_2307,N_24816,N_24994);
or UO_2308 (O_2308,N_24950,N_24838);
or UO_2309 (O_2309,N_24812,N_24976);
xnor UO_2310 (O_2310,N_24903,N_24934);
xor UO_2311 (O_2311,N_24938,N_24970);
nor UO_2312 (O_2312,N_24919,N_24972);
xor UO_2313 (O_2313,N_24986,N_24929);
and UO_2314 (O_2314,N_24895,N_24996);
nor UO_2315 (O_2315,N_24834,N_24820);
nor UO_2316 (O_2316,N_24999,N_24933);
xnor UO_2317 (O_2317,N_24840,N_24903);
and UO_2318 (O_2318,N_24851,N_24945);
and UO_2319 (O_2319,N_24998,N_24879);
xor UO_2320 (O_2320,N_24946,N_24841);
nand UO_2321 (O_2321,N_24919,N_24816);
nor UO_2322 (O_2322,N_24910,N_24886);
xor UO_2323 (O_2323,N_24830,N_24866);
nor UO_2324 (O_2324,N_24910,N_24933);
xor UO_2325 (O_2325,N_24865,N_24915);
nand UO_2326 (O_2326,N_24839,N_24804);
xnor UO_2327 (O_2327,N_24928,N_24951);
or UO_2328 (O_2328,N_24946,N_24959);
nand UO_2329 (O_2329,N_24969,N_24854);
nor UO_2330 (O_2330,N_24894,N_24889);
or UO_2331 (O_2331,N_24997,N_24984);
and UO_2332 (O_2332,N_24917,N_24895);
xnor UO_2333 (O_2333,N_24807,N_24904);
or UO_2334 (O_2334,N_24978,N_24853);
nor UO_2335 (O_2335,N_24881,N_24890);
nand UO_2336 (O_2336,N_24810,N_24950);
xnor UO_2337 (O_2337,N_24978,N_24963);
and UO_2338 (O_2338,N_24973,N_24826);
xor UO_2339 (O_2339,N_24914,N_24935);
nand UO_2340 (O_2340,N_24805,N_24802);
nand UO_2341 (O_2341,N_24818,N_24918);
and UO_2342 (O_2342,N_24979,N_24998);
xnor UO_2343 (O_2343,N_24939,N_24941);
and UO_2344 (O_2344,N_24895,N_24953);
and UO_2345 (O_2345,N_24921,N_24885);
nand UO_2346 (O_2346,N_24949,N_24803);
nor UO_2347 (O_2347,N_24802,N_24838);
or UO_2348 (O_2348,N_24806,N_24958);
nand UO_2349 (O_2349,N_24987,N_24910);
or UO_2350 (O_2350,N_24813,N_24942);
and UO_2351 (O_2351,N_24924,N_24932);
or UO_2352 (O_2352,N_24916,N_24932);
nand UO_2353 (O_2353,N_24975,N_24953);
nand UO_2354 (O_2354,N_24856,N_24838);
nand UO_2355 (O_2355,N_24944,N_24897);
and UO_2356 (O_2356,N_24995,N_24919);
nand UO_2357 (O_2357,N_24816,N_24842);
nor UO_2358 (O_2358,N_24988,N_24895);
nand UO_2359 (O_2359,N_24905,N_24898);
xnor UO_2360 (O_2360,N_24857,N_24894);
xnor UO_2361 (O_2361,N_24971,N_24901);
or UO_2362 (O_2362,N_24895,N_24869);
nand UO_2363 (O_2363,N_24896,N_24929);
nor UO_2364 (O_2364,N_24832,N_24992);
and UO_2365 (O_2365,N_24858,N_24983);
nand UO_2366 (O_2366,N_24962,N_24995);
nor UO_2367 (O_2367,N_24891,N_24982);
nand UO_2368 (O_2368,N_24916,N_24931);
xnor UO_2369 (O_2369,N_24924,N_24841);
and UO_2370 (O_2370,N_24846,N_24971);
nand UO_2371 (O_2371,N_24871,N_24800);
or UO_2372 (O_2372,N_24892,N_24997);
nand UO_2373 (O_2373,N_24800,N_24988);
xor UO_2374 (O_2374,N_24817,N_24976);
nand UO_2375 (O_2375,N_24929,N_24844);
or UO_2376 (O_2376,N_24987,N_24823);
nand UO_2377 (O_2377,N_24831,N_24842);
and UO_2378 (O_2378,N_24821,N_24807);
or UO_2379 (O_2379,N_24923,N_24939);
nor UO_2380 (O_2380,N_24882,N_24995);
or UO_2381 (O_2381,N_24864,N_24954);
or UO_2382 (O_2382,N_24919,N_24882);
nand UO_2383 (O_2383,N_24973,N_24825);
or UO_2384 (O_2384,N_24954,N_24991);
xnor UO_2385 (O_2385,N_24804,N_24886);
nor UO_2386 (O_2386,N_24932,N_24912);
xnor UO_2387 (O_2387,N_24988,N_24803);
or UO_2388 (O_2388,N_24916,N_24891);
nand UO_2389 (O_2389,N_24832,N_24817);
nand UO_2390 (O_2390,N_24822,N_24809);
xnor UO_2391 (O_2391,N_24800,N_24834);
nand UO_2392 (O_2392,N_24959,N_24820);
nand UO_2393 (O_2393,N_24876,N_24883);
xor UO_2394 (O_2394,N_24899,N_24942);
nand UO_2395 (O_2395,N_24944,N_24921);
or UO_2396 (O_2396,N_24866,N_24935);
and UO_2397 (O_2397,N_24979,N_24896);
nand UO_2398 (O_2398,N_24989,N_24933);
xor UO_2399 (O_2399,N_24953,N_24842);
and UO_2400 (O_2400,N_24996,N_24868);
and UO_2401 (O_2401,N_24932,N_24825);
nand UO_2402 (O_2402,N_24984,N_24875);
and UO_2403 (O_2403,N_24956,N_24994);
nor UO_2404 (O_2404,N_24928,N_24882);
or UO_2405 (O_2405,N_24888,N_24856);
nor UO_2406 (O_2406,N_24813,N_24870);
nor UO_2407 (O_2407,N_24830,N_24919);
or UO_2408 (O_2408,N_24841,N_24866);
xnor UO_2409 (O_2409,N_24940,N_24857);
and UO_2410 (O_2410,N_24910,N_24854);
nand UO_2411 (O_2411,N_24942,N_24892);
nand UO_2412 (O_2412,N_24841,N_24805);
nand UO_2413 (O_2413,N_24887,N_24961);
xor UO_2414 (O_2414,N_24859,N_24999);
and UO_2415 (O_2415,N_24851,N_24903);
or UO_2416 (O_2416,N_24947,N_24835);
or UO_2417 (O_2417,N_24991,N_24923);
and UO_2418 (O_2418,N_24880,N_24860);
and UO_2419 (O_2419,N_24837,N_24813);
or UO_2420 (O_2420,N_24873,N_24916);
nand UO_2421 (O_2421,N_24810,N_24983);
nand UO_2422 (O_2422,N_24959,N_24859);
xnor UO_2423 (O_2423,N_24801,N_24808);
nand UO_2424 (O_2424,N_24811,N_24959);
and UO_2425 (O_2425,N_24980,N_24865);
xor UO_2426 (O_2426,N_24916,N_24974);
nand UO_2427 (O_2427,N_24899,N_24932);
or UO_2428 (O_2428,N_24905,N_24987);
or UO_2429 (O_2429,N_24935,N_24905);
nand UO_2430 (O_2430,N_24831,N_24823);
xnor UO_2431 (O_2431,N_24878,N_24951);
nand UO_2432 (O_2432,N_24811,N_24924);
and UO_2433 (O_2433,N_24928,N_24999);
or UO_2434 (O_2434,N_24838,N_24826);
nand UO_2435 (O_2435,N_24800,N_24849);
xnor UO_2436 (O_2436,N_24958,N_24867);
xor UO_2437 (O_2437,N_24815,N_24891);
xor UO_2438 (O_2438,N_24808,N_24926);
and UO_2439 (O_2439,N_24996,N_24849);
and UO_2440 (O_2440,N_24827,N_24902);
or UO_2441 (O_2441,N_24978,N_24890);
nand UO_2442 (O_2442,N_24900,N_24926);
nand UO_2443 (O_2443,N_24821,N_24850);
and UO_2444 (O_2444,N_24810,N_24978);
xnor UO_2445 (O_2445,N_24820,N_24833);
nor UO_2446 (O_2446,N_24937,N_24842);
xor UO_2447 (O_2447,N_24913,N_24903);
or UO_2448 (O_2448,N_24961,N_24847);
xor UO_2449 (O_2449,N_24958,N_24863);
and UO_2450 (O_2450,N_24940,N_24928);
and UO_2451 (O_2451,N_24807,N_24969);
nand UO_2452 (O_2452,N_24995,N_24886);
nand UO_2453 (O_2453,N_24874,N_24915);
xor UO_2454 (O_2454,N_24993,N_24885);
nand UO_2455 (O_2455,N_24962,N_24990);
or UO_2456 (O_2456,N_24840,N_24916);
and UO_2457 (O_2457,N_24871,N_24936);
nor UO_2458 (O_2458,N_24819,N_24891);
and UO_2459 (O_2459,N_24958,N_24932);
nor UO_2460 (O_2460,N_24985,N_24906);
nand UO_2461 (O_2461,N_24971,N_24998);
nor UO_2462 (O_2462,N_24885,N_24971);
or UO_2463 (O_2463,N_24923,N_24832);
or UO_2464 (O_2464,N_24941,N_24858);
xor UO_2465 (O_2465,N_24815,N_24940);
and UO_2466 (O_2466,N_24870,N_24927);
nand UO_2467 (O_2467,N_24985,N_24945);
nand UO_2468 (O_2468,N_24974,N_24849);
nand UO_2469 (O_2469,N_24970,N_24810);
nand UO_2470 (O_2470,N_24935,N_24853);
nand UO_2471 (O_2471,N_24820,N_24854);
nor UO_2472 (O_2472,N_24912,N_24944);
or UO_2473 (O_2473,N_24961,N_24833);
or UO_2474 (O_2474,N_24972,N_24857);
nor UO_2475 (O_2475,N_24805,N_24860);
xor UO_2476 (O_2476,N_24936,N_24962);
nand UO_2477 (O_2477,N_24906,N_24999);
nor UO_2478 (O_2478,N_24965,N_24881);
nor UO_2479 (O_2479,N_24958,N_24842);
xnor UO_2480 (O_2480,N_24958,N_24946);
xnor UO_2481 (O_2481,N_24995,N_24862);
and UO_2482 (O_2482,N_24973,N_24939);
nor UO_2483 (O_2483,N_24836,N_24948);
and UO_2484 (O_2484,N_24867,N_24812);
nor UO_2485 (O_2485,N_24882,N_24984);
nor UO_2486 (O_2486,N_24872,N_24985);
xnor UO_2487 (O_2487,N_24846,N_24911);
or UO_2488 (O_2488,N_24828,N_24885);
nor UO_2489 (O_2489,N_24931,N_24917);
nor UO_2490 (O_2490,N_24935,N_24882);
or UO_2491 (O_2491,N_24809,N_24893);
and UO_2492 (O_2492,N_24834,N_24863);
and UO_2493 (O_2493,N_24942,N_24825);
or UO_2494 (O_2494,N_24991,N_24836);
nor UO_2495 (O_2495,N_24991,N_24936);
and UO_2496 (O_2496,N_24932,N_24811);
nand UO_2497 (O_2497,N_24956,N_24867);
or UO_2498 (O_2498,N_24882,N_24840);
and UO_2499 (O_2499,N_24810,N_24959);
or UO_2500 (O_2500,N_24995,N_24915);
xor UO_2501 (O_2501,N_24964,N_24918);
or UO_2502 (O_2502,N_24875,N_24929);
nand UO_2503 (O_2503,N_24900,N_24838);
xnor UO_2504 (O_2504,N_24887,N_24931);
nand UO_2505 (O_2505,N_24834,N_24841);
nor UO_2506 (O_2506,N_24986,N_24962);
or UO_2507 (O_2507,N_24891,N_24860);
nand UO_2508 (O_2508,N_24947,N_24805);
nor UO_2509 (O_2509,N_24986,N_24932);
xor UO_2510 (O_2510,N_24888,N_24928);
nand UO_2511 (O_2511,N_24861,N_24930);
and UO_2512 (O_2512,N_24987,N_24874);
nor UO_2513 (O_2513,N_24881,N_24920);
nand UO_2514 (O_2514,N_24836,N_24809);
or UO_2515 (O_2515,N_24942,N_24914);
and UO_2516 (O_2516,N_24831,N_24969);
xor UO_2517 (O_2517,N_24997,N_24854);
and UO_2518 (O_2518,N_24933,N_24879);
and UO_2519 (O_2519,N_24927,N_24868);
and UO_2520 (O_2520,N_24923,N_24945);
or UO_2521 (O_2521,N_24989,N_24939);
nand UO_2522 (O_2522,N_24922,N_24889);
nor UO_2523 (O_2523,N_24969,N_24877);
and UO_2524 (O_2524,N_24992,N_24896);
nand UO_2525 (O_2525,N_24814,N_24824);
nand UO_2526 (O_2526,N_24952,N_24843);
nand UO_2527 (O_2527,N_24895,N_24843);
nand UO_2528 (O_2528,N_24852,N_24838);
and UO_2529 (O_2529,N_24849,N_24962);
and UO_2530 (O_2530,N_24923,N_24875);
xor UO_2531 (O_2531,N_24809,N_24863);
nor UO_2532 (O_2532,N_24853,N_24862);
nor UO_2533 (O_2533,N_24958,N_24995);
and UO_2534 (O_2534,N_24954,N_24856);
and UO_2535 (O_2535,N_24872,N_24888);
or UO_2536 (O_2536,N_24911,N_24822);
or UO_2537 (O_2537,N_24965,N_24960);
nand UO_2538 (O_2538,N_24930,N_24901);
xor UO_2539 (O_2539,N_24915,N_24807);
xnor UO_2540 (O_2540,N_24964,N_24901);
or UO_2541 (O_2541,N_24947,N_24834);
and UO_2542 (O_2542,N_24883,N_24814);
nor UO_2543 (O_2543,N_24838,N_24807);
nand UO_2544 (O_2544,N_24875,N_24864);
nor UO_2545 (O_2545,N_24867,N_24981);
or UO_2546 (O_2546,N_24890,N_24906);
nand UO_2547 (O_2547,N_24958,N_24827);
nor UO_2548 (O_2548,N_24911,N_24871);
or UO_2549 (O_2549,N_24831,N_24964);
nand UO_2550 (O_2550,N_24990,N_24830);
nand UO_2551 (O_2551,N_24971,N_24949);
nand UO_2552 (O_2552,N_24898,N_24883);
or UO_2553 (O_2553,N_24826,N_24806);
and UO_2554 (O_2554,N_24802,N_24807);
xor UO_2555 (O_2555,N_24953,N_24940);
or UO_2556 (O_2556,N_24945,N_24995);
nor UO_2557 (O_2557,N_24819,N_24983);
and UO_2558 (O_2558,N_24914,N_24979);
xor UO_2559 (O_2559,N_24942,N_24963);
and UO_2560 (O_2560,N_24872,N_24863);
nand UO_2561 (O_2561,N_24831,N_24888);
or UO_2562 (O_2562,N_24871,N_24977);
and UO_2563 (O_2563,N_24903,N_24919);
xor UO_2564 (O_2564,N_24983,N_24940);
nor UO_2565 (O_2565,N_24997,N_24985);
nand UO_2566 (O_2566,N_24821,N_24915);
or UO_2567 (O_2567,N_24930,N_24959);
or UO_2568 (O_2568,N_24824,N_24953);
or UO_2569 (O_2569,N_24932,N_24867);
and UO_2570 (O_2570,N_24874,N_24932);
or UO_2571 (O_2571,N_24961,N_24809);
nand UO_2572 (O_2572,N_24997,N_24926);
xnor UO_2573 (O_2573,N_24855,N_24868);
nand UO_2574 (O_2574,N_24922,N_24948);
nand UO_2575 (O_2575,N_24933,N_24973);
nand UO_2576 (O_2576,N_24830,N_24806);
or UO_2577 (O_2577,N_24860,N_24848);
and UO_2578 (O_2578,N_24878,N_24871);
or UO_2579 (O_2579,N_24801,N_24878);
nand UO_2580 (O_2580,N_24886,N_24978);
and UO_2581 (O_2581,N_24819,N_24971);
nand UO_2582 (O_2582,N_24833,N_24938);
or UO_2583 (O_2583,N_24848,N_24920);
nor UO_2584 (O_2584,N_24938,N_24864);
or UO_2585 (O_2585,N_24900,N_24975);
nor UO_2586 (O_2586,N_24825,N_24820);
and UO_2587 (O_2587,N_24878,N_24898);
and UO_2588 (O_2588,N_24964,N_24915);
or UO_2589 (O_2589,N_24823,N_24970);
nor UO_2590 (O_2590,N_24833,N_24850);
and UO_2591 (O_2591,N_24890,N_24858);
and UO_2592 (O_2592,N_24901,N_24865);
nand UO_2593 (O_2593,N_24853,N_24913);
nand UO_2594 (O_2594,N_24966,N_24902);
xor UO_2595 (O_2595,N_24881,N_24830);
and UO_2596 (O_2596,N_24825,N_24805);
nand UO_2597 (O_2597,N_24855,N_24998);
or UO_2598 (O_2598,N_24978,N_24971);
nand UO_2599 (O_2599,N_24834,N_24819);
nand UO_2600 (O_2600,N_24831,N_24931);
or UO_2601 (O_2601,N_24859,N_24955);
nand UO_2602 (O_2602,N_24827,N_24933);
nor UO_2603 (O_2603,N_24853,N_24914);
or UO_2604 (O_2604,N_24887,N_24903);
and UO_2605 (O_2605,N_24912,N_24964);
nand UO_2606 (O_2606,N_24918,N_24842);
nand UO_2607 (O_2607,N_24999,N_24882);
or UO_2608 (O_2608,N_24945,N_24906);
or UO_2609 (O_2609,N_24851,N_24835);
and UO_2610 (O_2610,N_24999,N_24940);
nor UO_2611 (O_2611,N_24867,N_24988);
nand UO_2612 (O_2612,N_24886,N_24930);
xor UO_2613 (O_2613,N_24849,N_24971);
nand UO_2614 (O_2614,N_24960,N_24846);
xor UO_2615 (O_2615,N_24885,N_24896);
xnor UO_2616 (O_2616,N_24806,N_24880);
or UO_2617 (O_2617,N_24936,N_24888);
nand UO_2618 (O_2618,N_24895,N_24897);
nor UO_2619 (O_2619,N_24995,N_24829);
and UO_2620 (O_2620,N_24963,N_24926);
or UO_2621 (O_2621,N_24849,N_24917);
and UO_2622 (O_2622,N_24805,N_24811);
nand UO_2623 (O_2623,N_24989,N_24865);
nor UO_2624 (O_2624,N_24880,N_24951);
nand UO_2625 (O_2625,N_24935,N_24826);
or UO_2626 (O_2626,N_24828,N_24960);
xnor UO_2627 (O_2627,N_24980,N_24918);
and UO_2628 (O_2628,N_24892,N_24859);
xor UO_2629 (O_2629,N_24877,N_24852);
and UO_2630 (O_2630,N_24868,N_24853);
nor UO_2631 (O_2631,N_24825,N_24923);
or UO_2632 (O_2632,N_24852,N_24811);
nor UO_2633 (O_2633,N_24879,N_24834);
and UO_2634 (O_2634,N_24820,N_24936);
nand UO_2635 (O_2635,N_24990,N_24952);
nand UO_2636 (O_2636,N_24936,N_24826);
nor UO_2637 (O_2637,N_24807,N_24978);
xor UO_2638 (O_2638,N_24840,N_24827);
and UO_2639 (O_2639,N_24936,N_24845);
xnor UO_2640 (O_2640,N_24840,N_24919);
or UO_2641 (O_2641,N_24819,N_24962);
xor UO_2642 (O_2642,N_24887,N_24874);
nand UO_2643 (O_2643,N_24998,N_24950);
or UO_2644 (O_2644,N_24996,N_24972);
nor UO_2645 (O_2645,N_24887,N_24936);
nor UO_2646 (O_2646,N_24939,N_24885);
nand UO_2647 (O_2647,N_24802,N_24813);
nor UO_2648 (O_2648,N_24964,N_24872);
xor UO_2649 (O_2649,N_24915,N_24892);
nand UO_2650 (O_2650,N_24974,N_24830);
nor UO_2651 (O_2651,N_24991,N_24833);
nor UO_2652 (O_2652,N_24995,N_24956);
and UO_2653 (O_2653,N_24973,N_24817);
and UO_2654 (O_2654,N_24963,N_24858);
nor UO_2655 (O_2655,N_24883,N_24994);
nand UO_2656 (O_2656,N_24813,N_24857);
nand UO_2657 (O_2657,N_24916,N_24946);
nand UO_2658 (O_2658,N_24891,N_24940);
or UO_2659 (O_2659,N_24897,N_24858);
or UO_2660 (O_2660,N_24958,N_24857);
nand UO_2661 (O_2661,N_24813,N_24855);
or UO_2662 (O_2662,N_24877,N_24900);
nand UO_2663 (O_2663,N_24965,N_24826);
xnor UO_2664 (O_2664,N_24807,N_24826);
or UO_2665 (O_2665,N_24823,N_24906);
nand UO_2666 (O_2666,N_24809,N_24820);
and UO_2667 (O_2667,N_24985,N_24816);
nor UO_2668 (O_2668,N_24843,N_24833);
xor UO_2669 (O_2669,N_24857,N_24964);
nor UO_2670 (O_2670,N_24881,N_24853);
or UO_2671 (O_2671,N_24897,N_24936);
nand UO_2672 (O_2672,N_24915,N_24842);
nand UO_2673 (O_2673,N_24906,N_24956);
nor UO_2674 (O_2674,N_24931,N_24924);
nand UO_2675 (O_2675,N_24982,N_24901);
and UO_2676 (O_2676,N_24890,N_24899);
nand UO_2677 (O_2677,N_24929,N_24889);
xnor UO_2678 (O_2678,N_24845,N_24816);
and UO_2679 (O_2679,N_24956,N_24915);
or UO_2680 (O_2680,N_24847,N_24876);
xnor UO_2681 (O_2681,N_24932,N_24920);
or UO_2682 (O_2682,N_24816,N_24958);
nand UO_2683 (O_2683,N_24926,N_24905);
or UO_2684 (O_2684,N_24867,N_24860);
nand UO_2685 (O_2685,N_24947,N_24922);
nand UO_2686 (O_2686,N_24949,N_24927);
nor UO_2687 (O_2687,N_24897,N_24883);
and UO_2688 (O_2688,N_24930,N_24999);
xor UO_2689 (O_2689,N_24988,N_24971);
or UO_2690 (O_2690,N_24942,N_24986);
or UO_2691 (O_2691,N_24990,N_24948);
or UO_2692 (O_2692,N_24937,N_24886);
xor UO_2693 (O_2693,N_24926,N_24850);
xnor UO_2694 (O_2694,N_24961,N_24951);
or UO_2695 (O_2695,N_24805,N_24867);
nor UO_2696 (O_2696,N_24827,N_24949);
or UO_2697 (O_2697,N_24848,N_24819);
and UO_2698 (O_2698,N_24975,N_24808);
or UO_2699 (O_2699,N_24991,N_24996);
nand UO_2700 (O_2700,N_24808,N_24875);
nand UO_2701 (O_2701,N_24842,N_24885);
nand UO_2702 (O_2702,N_24884,N_24997);
xnor UO_2703 (O_2703,N_24940,N_24951);
nor UO_2704 (O_2704,N_24902,N_24904);
nand UO_2705 (O_2705,N_24875,N_24997);
xor UO_2706 (O_2706,N_24921,N_24943);
and UO_2707 (O_2707,N_24971,N_24987);
or UO_2708 (O_2708,N_24943,N_24850);
and UO_2709 (O_2709,N_24947,N_24811);
nor UO_2710 (O_2710,N_24926,N_24973);
xor UO_2711 (O_2711,N_24997,N_24825);
xor UO_2712 (O_2712,N_24973,N_24875);
and UO_2713 (O_2713,N_24835,N_24876);
xor UO_2714 (O_2714,N_24930,N_24868);
or UO_2715 (O_2715,N_24965,N_24966);
nand UO_2716 (O_2716,N_24833,N_24839);
xnor UO_2717 (O_2717,N_24897,N_24803);
nor UO_2718 (O_2718,N_24853,N_24806);
xor UO_2719 (O_2719,N_24948,N_24846);
and UO_2720 (O_2720,N_24910,N_24820);
xnor UO_2721 (O_2721,N_24897,N_24865);
nor UO_2722 (O_2722,N_24822,N_24900);
or UO_2723 (O_2723,N_24904,N_24960);
xnor UO_2724 (O_2724,N_24847,N_24970);
nor UO_2725 (O_2725,N_24852,N_24850);
and UO_2726 (O_2726,N_24896,N_24837);
xnor UO_2727 (O_2727,N_24837,N_24968);
nand UO_2728 (O_2728,N_24972,N_24852);
nand UO_2729 (O_2729,N_24846,N_24966);
xor UO_2730 (O_2730,N_24896,N_24850);
and UO_2731 (O_2731,N_24946,N_24811);
nor UO_2732 (O_2732,N_24925,N_24920);
nor UO_2733 (O_2733,N_24926,N_24902);
nand UO_2734 (O_2734,N_24912,N_24909);
nor UO_2735 (O_2735,N_24982,N_24831);
or UO_2736 (O_2736,N_24882,N_24909);
nor UO_2737 (O_2737,N_24979,N_24862);
xnor UO_2738 (O_2738,N_24818,N_24841);
nand UO_2739 (O_2739,N_24800,N_24939);
and UO_2740 (O_2740,N_24853,N_24879);
nand UO_2741 (O_2741,N_24896,N_24900);
xnor UO_2742 (O_2742,N_24859,N_24836);
or UO_2743 (O_2743,N_24956,N_24911);
xnor UO_2744 (O_2744,N_24803,N_24935);
and UO_2745 (O_2745,N_24925,N_24889);
or UO_2746 (O_2746,N_24936,N_24964);
nor UO_2747 (O_2747,N_24849,N_24986);
xnor UO_2748 (O_2748,N_24948,N_24935);
or UO_2749 (O_2749,N_24982,N_24953);
or UO_2750 (O_2750,N_24875,N_24890);
xnor UO_2751 (O_2751,N_24836,N_24830);
or UO_2752 (O_2752,N_24865,N_24814);
xor UO_2753 (O_2753,N_24979,N_24871);
or UO_2754 (O_2754,N_24931,N_24821);
and UO_2755 (O_2755,N_24922,N_24841);
and UO_2756 (O_2756,N_24858,N_24966);
nor UO_2757 (O_2757,N_24921,N_24886);
xor UO_2758 (O_2758,N_24875,N_24814);
and UO_2759 (O_2759,N_24918,N_24961);
or UO_2760 (O_2760,N_24908,N_24804);
or UO_2761 (O_2761,N_24871,N_24891);
nand UO_2762 (O_2762,N_24919,N_24886);
xnor UO_2763 (O_2763,N_24940,N_24886);
and UO_2764 (O_2764,N_24858,N_24914);
and UO_2765 (O_2765,N_24832,N_24845);
nand UO_2766 (O_2766,N_24981,N_24887);
or UO_2767 (O_2767,N_24806,N_24949);
xor UO_2768 (O_2768,N_24835,N_24889);
or UO_2769 (O_2769,N_24841,N_24901);
or UO_2770 (O_2770,N_24918,N_24846);
or UO_2771 (O_2771,N_24838,N_24957);
or UO_2772 (O_2772,N_24800,N_24872);
xnor UO_2773 (O_2773,N_24851,N_24866);
and UO_2774 (O_2774,N_24912,N_24930);
or UO_2775 (O_2775,N_24930,N_24969);
nand UO_2776 (O_2776,N_24979,N_24949);
or UO_2777 (O_2777,N_24808,N_24827);
xnor UO_2778 (O_2778,N_24832,N_24958);
and UO_2779 (O_2779,N_24996,N_24923);
xor UO_2780 (O_2780,N_24952,N_24940);
nor UO_2781 (O_2781,N_24812,N_24999);
or UO_2782 (O_2782,N_24869,N_24881);
nand UO_2783 (O_2783,N_24873,N_24958);
or UO_2784 (O_2784,N_24979,N_24875);
xor UO_2785 (O_2785,N_24917,N_24916);
nand UO_2786 (O_2786,N_24907,N_24842);
xnor UO_2787 (O_2787,N_24929,N_24852);
xor UO_2788 (O_2788,N_24987,N_24947);
or UO_2789 (O_2789,N_24843,N_24970);
or UO_2790 (O_2790,N_24977,N_24950);
nor UO_2791 (O_2791,N_24859,N_24914);
xnor UO_2792 (O_2792,N_24906,N_24935);
nor UO_2793 (O_2793,N_24842,N_24853);
nor UO_2794 (O_2794,N_24832,N_24961);
nand UO_2795 (O_2795,N_24888,N_24950);
xor UO_2796 (O_2796,N_24835,N_24981);
and UO_2797 (O_2797,N_24817,N_24818);
xor UO_2798 (O_2798,N_24916,N_24987);
xor UO_2799 (O_2799,N_24997,N_24999);
or UO_2800 (O_2800,N_24851,N_24914);
nand UO_2801 (O_2801,N_24983,N_24828);
xor UO_2802 (O_2802,N_24968,N_24823);
xor UO_2803 (O_2803,N_24875,N_24938);
and UO_2804 (O_2804,N_24983,N_24911);
or UO_2805 (O_2805,N_24921,N_24883);
and UO_2806 (O_2806,N_24885,N_24954);
nand UO_2807 (O_2807,N_24922,N_24883);
nand UO_2808 (O_2808,N_24958,N_24866);
xnor UO_2809 (O_2809,N_24823,N_24916);
nand UO_2810 (O_2810,N_24955,N_24805);
xnor UO_2811 (O_2811,N_24849,N_24932);
nand UO_2812 (O_2812,N_24905,N_24947);
and UO_2813 (O_2813,N_24825,N_24852);
xnor UO_2814 (O_2814,N_24892,N_24861);
xor UO_2815 (O_2815,N_24966,N_24926);
nor UO_2816 (O_2816,N_24860,N_24817);
and UO_2817 (O_2817,N_24929,N_24914);
and UO_2818 (O_2818,N_24929,N_24863);
or UO_2819 (O_2819,N_24909,N_24814);
nor UO_2820 (O_2820,N_24867,N_24918);
xnor UO_2821 (O_2821,N_24992,N_24902);
nand UO_2822 (O_2822,N_24843,N_24950);
xor UO_2823 (O_2823,N_24883,N_24971);
nand UO_2824 (O_2824,N_24942,N_24966);
xor UO_2825 (O_2825,N_24983,N_24938);
nor UO_2826 (O_2826,N_24996,N_24949);
or UO_2827 (O_2827,N_24975,N_24976);
and UO_2828 (O_2828,N_24814,N_24963);
xor UO_2829 (O_2829,N_24898,N_24964);
nand UO_2830 (O_2830,N_24916,N_24817);
xor UO_2831 (O_2831,N_24874,N_24921);
xor UO_2832 (O_2832,N_24855,N_24983);
nand UO_2833 (O_2833,N_24891,N_24886);
nand UO_2834 (O_2834,N_24844,N_24878);
nand UO_2835 (O_2835,N_24889,N_24955);
and UO_2836 (O_2836,N_24983,N_24968);
xnor UO_2837 (O_2837,N_24922,N_24825);
nand UO_2838 (O_2838,N_24945,N_24863);
and UO_2839 (O_2839,N_24904,N_24991);
nor UO_2840 (O_2840,N_24993,N_24825);
nor UO_2841 (O_2841,N_24967,N_24909);
or UO_2842 (O_2842,N_24928,N_24867);
nor UO_2843 (O_2843,N_24981,N_24912);
xor UO_2844 (O_2844,N_24991,N_24846);
xnor UO_2845 (O_2845,N_24834,N_24808);
xor UO_2846 (O_2846,N_24859,N_24996);
or UO_2847 (O_2847,N_24841,N_24842);
or UO_2848 (O_2848,N_24809,N_24828);
xnor UO_2849 (O_2849,N_24921,N_24965);
or UO_2850 (O_2850,N_24918,N_24986);
nand UO_2851 (O_2851,N_24918,N_24957);
nand UO_2852 (O_2852,N_24979,N_24967);
or UO_2853 (O_2853,N_24939,N_24878);
nor UO_2854 (O_2854,N_24965,N_24812);
nor UO_2855 (O_2855,N_24958,N_24804);
or UO_2856 (O_2856,N_24885,N_24868);
and UO_2857 (O_2857,N_24807,N_24897);
nand UO_2858 (O_2858,N_24846,N_24958);
nand UO_2859 (O_2859,N_24808,N_24913);
xor UO_2860 (O_2860,N_24929,N_24942);
nand UO_2861 (O_2861,N_24856,N_24993);
nand UO_2862 (O_2862,N_24836,N_24852);
or UO_2863 (O_2863,N_24957,N_24953);
nor UO_2864 (O_2864,N_24965,N_24923);
or UO_2865 (O_2865,N_24925,N_24928);
nand UO_2866 (O_2866,N_24941,N_24973);
xnor UO_2867 (O_2867,N_24951,N_24934);
or UO_2868 (O_2868,N_24944,N_24949);
or UO_2869 (O_2869,N_24877,N_24927);
nand UO_2870 (O_2870,N_24904,N_24997);
or UO_2871 (O_2871,N_24809,N_24864);
nand UO_2872 (O_2872,N_24996,N_24889);
or UO_2873 (O_2873,N_24869,N_24939);
and UO_2874 (O_2874,N_24938,N_24885);
xnor UO_2875 (O_2875,N_24833,N_24982);
or UO_2876 (O_2876,N_24809,N_24980);
nor UO_2877 (O_2877,N_24933,N_24974);
nand UO_2878 (O_2878,N_24940,N_24806);
nor UO_2879 (O_2879,N_24981,N_24896);
xnor UO_2880 (O_2880,N_24819,N_24894);
nand UO_2881 (O_2881,N_24972,N_24913);
or UO_2882 (O_2882,N_24918,N_24833);
nand UO_2883 (O_2883,N_24867,N_24846);
and UO_2884 (O_2884,N_24942,N_24928);
nor UO_2885 (O_2885,N_24876,N_24970);
or UO_2886 (O_2886,N_24809,N_24981);
nand UO_2887 (O_2887,N_24866,N_24856);
xor UO_2888 (O_2888,N_24982,N_24943);
nor UO_2889 (O_2889,N_24904,N_24876);
nand UO_2890 (O_2890,N_24993,N_24806);
xnor UO_2891 (O_2891,N_24852,N_24999);
nand UO_2892 (O_2892,N_24955,N_24814);
nor UO_2893 (O_2893,N_24893,N_24914);
or UO_2894 (O_2894,N_24836,N_24915);
and UO_2895 (O_2895,N_24801,N_24906);
or UO_2896 (O_2896,N_24932,N_24941);
or UO_2897 (O_2897,N_24941,N_24890);
or UO_2898 (O_2898,N_24817,N_24951);
or UO_2899 (O_2899,N_24807,N_24836);
nor UO_2900 (O_2900,N_24994,N_24977);
and UO_2901 (O_2901,N_24909,N_24969);
and UO_2902 (O_2902,N_24867,N_24905);
nor UO_2903 (O_2903,N_24995,N_24997);
xor UO_2904 (O_2904,N_24968,N_24826);
or UO_2905 (O_2905,N_24941,N_24884);
nor UO_2906 (O_2906,N_24962,N_24944);
or UO_2907 (O_2907,N_24985,N_24873);
or UO_2908 (O_2908,N_24860,N_24875);
or UO_2909 (O_2909,N_24816,N_24879);
nand UO_2910 (O_2910,N_24829,N_24915);
nand UO_2911 (O_2911,N_24905,N_24802);
or UO_2912 (O_2912,N_24875,N_24897);
xnor UO_2913 (O_2913,N_24919,N_24946);
or UO_2914 (O_2914,N_24985,N_24937);
xor UO_2915 (O_2915,N_24853,N_24920);
and UO_2916 (O_2916,N_24916,N_24888);
xnor UO_2917 (O_2917,N_24887,N_24940);
or UO_2918 (O_2918,N_24859,N_24846);
nor UO_2919 (O_2919,N_24957,N_24817);
and UO_2920 (O_2920,N_24933,N_24880);
or UO_2921 (O_2921,N_24880,N_24962);
nor UO_2922 (O_2922,N_24878,N_24925);
nor UO_2923 (O_2923,N_24909,N_24849);
and UO_2924 (O_2924,N_24991,N_24803);
and UO_2925 (O_2925,N_24875,N_24886);
and UO_2926 (O_2926,N_24892,N_24927);
nor UO_2927 (O_2927,N_24817,N_24850);
and UO_2928 (O_2928,N_24834,N_24895);
xnor UO_2929 (O_2929,N_24882,N_24881);
and UO_2930 (O_2930,N_24983,N_24873);
xor UO_2931 (O_2931,N_24825,N_24853);
nor UO_2932 (O_2932,N_24955,N_24851);
xor UO_2933 (O_2933,N_24935,N_24840);
nor UO_2934 (O_2934,N_24819,N_24902);
nand UO_2935 (O_2935,N_24923,N_24976);
or UO_2936 (O_2936,N_24833,N_24912);
nand UO_2937 (O_2937,N_24874,N_24845);
nand UO_2938 (O_2938,N_24869,N_24873);
nor UO_2939 (O_2939,N_24885,N_24910);
or UO_2940 (O_2940,N_24812,N_24884);
xnor UO_2941 (O_2941,N_24944,N_24970);
nor UO_2942 (O_2942,N_24934,N_24921);
nand UO_2943 (O_2943,N_24857,N_24859);
or UO_2944 (O_2944,N_24932,N_24939);
nor UO_2945 (O_2945,N_24816,N_24903);
xnor UO_2946 (O_2946,N_24831,N_24832);
xor UO_2947 (O_2947,N_24818,N_24974);
and UO_2948 (O_2948,N_24882,N_24822);
nor UO_2949 (O_2949,N_24960,N_24839);
xor UO_2950 (O_2950,N_24932,N_24879);
xor UO_2951 (O_2951,N_24957,N_24889);
xor UO_2952 (O_2952,N_24994,N_24801);
nand UO_2953 (O_2953,N_24972,N_24899);
xnor UO_2954 (O_2954,N_24902,N_24969);
nor UO_2955 (O_2955,N_24835,N_24841);
or UO_2956 (O_2956,N_24890,N_24840);
or UO_2957 (O_2957,N_24914,N_24837);
nor UO_2958 (O_2958,N_24941,N_24847);
or UO_2959 (O_2959,N_24933,N_24878);
xor UO_2960 (O_2960,N_24979,N_24906);
and UO_2961 (O_2961,N_24820,N_24997);
nor UO_2962 (O_2962,N_24881,N_24990);
and UO_2963 (O_2963,N_24917,N_24963);
nand UO_2964 (O_2964,N_24949,N_24919);
nand UO_2965 (O_2965,N_24938,N_24846);
nor UO_2966 (O_2966,N_24931,N_24888);
nand UO_2967 (O_2967,N_24983,N_24827);
nand UO_2968 (O_2968,N_24885,N_24959);
and UO_2969 (O_2969,N_24836,N_24923);
nor UO_2970 (O_2970,N_24981,N_24841);
xnor UO_2971 (O_2971,N_24966,N_24941);
nand UO_2972 (O_2972,N_24910,N_24806);
and UO_2973 (O_2973,N_24954,N_24984);
xor UO_2974 (O_2974,N_24808,N_24895);
and UO_2975 (O_2975,N_24948,N_24994);
and UO_2976 (O_2976,N_24921,N_24898);
xor UO_2977 (O_2977,N_24865,N_24847);
nor UO_2978 (O_2978,N_24862,N_24902);
and UO_2979 (O_2979,N_24953,N_24911);
nor UO_2980 (O_2980,N_24995,N_24989);
or UO_2981 (O_2981,N_24975,N_24941);
xor UO_2982 (O_2982,N_24995,N_24885);
nor UO_2983 (O_2983,N_24827,N_24931);
nor UO_2984 (O_2984,N_24984,N_24872);
and UO_2985 (O_2985,N_24905,N_24842);
nand UO_2986 (O_2986,N_24894,N_24986);
xor UO_2987 (O_2987,N_24879,N_24830);
or UO_2988 (O_2988,N_24939,N_24808);
nand UO_2989 (O_2989,N_24842,N_24872);
xor UO_2990 (O_2990,N_24991,N_24814);
or UO_2991 (O_2991,N_24831,N_24998);
nor UO_2992 (O_2992,N_24941,N_24907);
nor UO_2993 (O_2993,N_24942,N_24890);
nand UO_2994 (O_2994,N_24829,N_24820);
or UO_2995 (O_2995,N_24967,N_24820);
or UO_2996 (O_2996,N_24994,N_24968);
or UO_2997 (O_2997,N_24863,N_24980);
xnor UO_2998 (O_2998,N_24936,N_24873);
xnor UO_2999 (O_2999,N_24864,N_24822);
endmodule