module basic_2500_25000_3000_125_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
xor U0 (N_0,In_1805,In_1286);
or U1 (N_1,In_2454,In_1703);
and U2 (N_2,In_1298,In_1190);
or U3 (N_3,In_1831,In_1880);
xor U4 (N_4,In_678,In_801);
and U5 (N_5,In_1213,In_1311);
nor U6 (N_6,In_799,In_1982);
xor U7 (N_7,In_2175,In_1818);
nor U8 (N_8,In_1525,In_478);
xnor U9 (N_9,In_462,In_1524);
nor U10 (N_10,In_1841,In_2464);
xnor U11 (N_11,In_2111,In_2030);
nor U12 (N_12,In_50,In_1523);
and U13 (N_13,In_1346,In_1074);
xnor U14 (N_14,In_1835,In_1948);
nor U15 (N_15,In_444,In_1887);
and U16 (N_16,In_683,In_1317);
and U17 (N_17,In_2140,In_403);
or U18 (N_18,In_429,In_1145);
nand U19 (N_19,In_103,In_2047);
nand U20 (N_20,In_398,In_452);
xor U21 (N_21,In_624,In_447);
or U22 (N_22,In_1438,In_1641);
and U23 (N_23,In_2142,In_976);
or U24 (N_24,In_2444,In_823);
nor U25 (N_25,In_198,In_148);
and U26 (N_26,In_658,In_641);
or U27 (N_27,In_1811,In_2399);
and U28 (N_28,In_1586,In_1284);
or U29 (N_29,In_36,In_391);
xnor U30 (N_30,In_1119,In_1856);
and U31 (N_31,In_1776,In_1384);
xnor U32 (N_32,In_703,In_773);
xor U33 (N_33,In_1543,In_622);
or U34 (N_34,In_1508,In_519);
xor U35 (N_35,In_2099,In_1810);
xnor U36 (N_36,In_1371,In_964);
nand U37 (N_37,In_433,In_1464);
xnor U38 (N_38,In_105,In_2096);
or U39 (N_39,In_535,In_1072);
nand U40 (N_40,In_1808,In_77);
nor U41 (N_41,In_2103,In_1191);
and U42 (N_42,In_66,In_432);
or U43 (N_43,In_1514,In_1949);
or U44 (N_44,In_2133,In_1839);
xor U45 (N_45,In_757,In_1106);
nor U46 (N_46,In_2062,In_1062);
nand U47 (N_47,In_257,In_680);
xnor U48 (N_48,In_1239,In_640);
and U49 (N_49,In_1915,In_459);
nor U50 (N_50,In_2429,In_158);
or U51 (N_51,In_1069,In_142);
xnor U52 (N_52,In_239,In_407);
nand U53 (N_53,In_379,In_2234);
or U54 (N_54,In_2194,In_1279);
or U55 (N_55,In_189,In_673);
xnor U56 (N_56,In_975,In_492);
nor U57 (N_57,In_1201,In_359);
nor U58 (N_58,In_1959,In_581);
nor U59 (N_59,In_1352,In_589);
or U60 (N_60,In_613,In_1614);
xnor U61 (N_61,In_1969,In_2008);
xnor U62 (N_62,In_372,In_90);
and U63 (N_63,In_438,In_1096);
or U64 (N_64,In_2421,In_39);
and U65 (N_65,In_895,In_2180);
nand U66 (N_66,In_917,In_1903);
nor U67 (N_67,In_950,In_1061);
nor U68 (N_68,In_902,In_605);
and U69 (N_69,In_1075,In_143);
xnor U70 (N_70,In_2431,In_109);
nor U71 (N_71,In_604,In_1488);
xor U72 (N_72,In_2017,In_2045);
nor U73 (N_73,In_1789,In_872);
and U74 (N_74,In_106,In_223);
xor U75 (N_75,In_301,In_999);
xnor U76 (N_76,In_1954,In_75);
nor U77 (N_77,In_911,In_25);
nand U78 (N_78,In_1761,In_237);
nor U79 (N_79,In_534,In_2182);
or U80 (N_80,In_590,In_650);
xnor U81 (N_81,In_1169,In_2317);
and U82 (N_82,In_855,In_939);
xor U83 (N_83,In_967,In_200);
nand U84 (N_84,In_1046,In_1058);
or U85 (N_85,In_783,In_1288);
nor U86 (N_86,In_974,In_1866);
nand U87 (N_87,In_120,In_254);
xnor U88 (N_88,In_1531,In_491);
and U89 (N_89,In_2488,In_207);
nand U90 (N_90,In_1055,In_1477);
nor U91 (N_91,In_108,In_34);
nand U92 (N_92,In_2442,In_1573);
nor U93 (N_93,In_928,In_921);
and U94 (N_94,In_953,In_990);
nand U95 (N_95,In_378,In_1217);
xor U96 (N_96,In_1581,In_1180);
and U97 (N_97,In_1219,In_1952);
xor U98 (N_98,In_162,In_2400);
nand U99 (N_99,In_1094,In_24);
nand U100 (N_100,In_1901,In_1362);
nand U101 (N_101,In_865,In_399);
xor U102 (N_102,In_1893,In_843);
xor U103 (N_103,In_1676,In_2087);
and U104 (N_104,In_2296,In_11);
nand U105 (N_105,In_933,In_2134);
nand U106 (N_106,In_451,In_83);
or U107 (N_107,In_2119,In_1842);
and U108 (N_108,In_194,In_576);
nor U109 (N_109,In_1374,In_297);
or U110 (N_110,In_819,In_185);
or U111 (N_111,In_664,In_1391);
and U112 (N_112,In_1146,In_636);
xnor U113 (N_113,In_1649,In_814);
and U114 (N_114,In_742,In_1924);
and U115 (N_115,In_1370,In_1481);
nand U116 (N_116,In_1174,In_635);
or U117 (N_117,In_436,In_2010);
nor U118 (N_118,In_2039,In_2208);
nor U119 (N_119,In_1824,In_419);
and U120 (N_120,In_116,In_2348);
or U121 (N_121,In_1913,In_1056);
xnor U122 (N_122,In_1702,In_569);
or U123 (N_123,In_335,In_1256);
nor U124 (N_124,In_212,In_1771);
nor U125 (N_125,In_1474,In_2462);
nand U126 (N_126,In_1020,In_1136);
or U127 (N_127,In_147,In_875);
or U128 (N_128,In_434,In_2128);
and U129 (N_129,In_2229,In_2426);
xor U130 (N_130,In_1829,In_1621);
or U131 (N_131,In_1153,In_2334);
nand U132 (N_132,In_1002,In_948);
or U133 (N_133,In_82,In_1411);
nand U134 (N_134,In_1602,In_2218);
and U135 (N_135,In_934,In_2281);
xnor U136 (N_136,In_1998,In_1116);
nor U137 (N_137,In_494,In_495);
nand U138 (N_138,In_838,In_2388);
nor U139 (N_139,In_1783,In_765);
xnor U140 (N_140,In_1232,In_520);
nand U141 (N_141,In_353,In_2210);
xnor U142 (N_142,In_1128,In_9);
nand U143 (N_143,In_114,In_1744);
or U144 (N_144,In_2040,In_1348);
and U145 (N_145,In_1950,In_259);
nor U146 (N_146,In_1125,In_1502);
or U147 (N_147,In_123,In_30);
xor U148 (N_148,In_1325,In_2490);
or U149 (N_149,In_1738,In_724);
nand U150 (N_150,In_722,In_1571);
nor U151 (N_151,In_1353,In_43);
xor U152 (N_152,In_1026,In_552);
nand U153 (N_153,In_1022,In_1506);
and U154 (N_154,In_1579,In_2223);
nor U155 (N_155,In_1343,In_2434);
and U156 (N_156,In_1678,In_562);
nor U157 (N_157,In_863,In_653);
nor U158 (N_158,In_1861,In_1);
and U159 (N_159,In_2084,In_1890);
and U160 (N_160,In_749,In_1513);
nor U161 (N_161,In_585,In_654);
nand U162 (N_162,In_2065,In_2201);
xnor U163 (N_163,In_1588,In_1512);
xor U164 (N_164,In_1942,In_1447);
nand U165 (N_165,In_2171,In_2420);
nand U166 (N_166,In_652,In_1705);
nor U167 (N_167,In_2287,In_1469);
and U168 (N_168,In_1051,In_1764);
nor U169 (N_169,In_1553,In_1150);
and U170 (N_170,In_949,In_2012);
or U171 (N_171,In_1028,In_392);
xnor U172 (N_172,In_1511,In_515);
nor U173 (N_173,In_512,In_2109);
xnor U174 (N_174,In_1987,In_352);
or U175 (N_175,In_1659,In_1635);
xnor U176 (N_176,In_1986,In_637);
xnor U177 (N_177,In_1908,In_2004);
nor U178 (N_178,In_346,In_2006);
and U179 (N_179,In_445,In_764);
nand U180 (N_180,In_2225,In_1114);
and U181 (N_181,In_1991,In_2410);
or U182 (N_182,In_2067,In_1547);
nor U183 (N_183,In_2104,In_1312);
nor U184 (N_184,In_446,In_815);
nor U185 (N_185,In_19,In_2107);
xnor U186 (N_186,In_2167,In_1953);
or U187 (N_187,In_1170,In_1463);
and U188 (N_188,In_1580,In_1912);
or U189 (N_189,In_140,In_2112);
or U190 (N_190,In_1570,In_2493);
nand U191 (N_191,In_2397,In_2301);
nand U192 (N_192,In_228,In_420);
and U193 (N_193,In_2494,In_2492);
and U194 (N_194,In_1455,In_1091);
nand U195 (N_195,In_238,In_2372);
and U196 (N_196,In_1409,In_1630);
nor U197 (N_197,In_1535,In_1309);
nor U198 (N_198,In_2110,In_1643);
or U199 (N_199,In_1875,In_49);
nor U200 (N_200,In_784,In_2054);
or U201 (N_201,In_1426,In_218);
or U202 (N_202,In_572,In_2079);
nor U203 (N_203,In_1961,N_197);
nor U204 (N_204,In_631,In_2115);
nor U205 (N_205,In_1567,In_970);
or U206 (N_206,In_1124,In_1461);
nand U207 (N_207,In_1395,In_1478);
nand U208 (N_208,In_1857,In_1656);
xor U209 (N_209,In_2286,In_1210);
nor U210 (N_210,In_2451,In_1040);
nand U211 (N_211,In_425,In_1574);
or U212 (N_212,In_595,In_827);
nor U213 (N_213,In_1785,In_596);
and U214 (N_214,In_1404,In_205);
nor U215 (N_215,In_348,In_2059);
xnor U216 (N_216,N_98,In_2335);
or U217 (N_217,In_2252,In_1425);
or U218 (N_218,In_575,In_1714);
or U219 (N_219,In_2144,N_191);
or U220 (N_220,In_376,N_139);
and U221 (N_221,In_2181,In_1819);
nor U222 (N_222,In_1501,In_1840);
xor U223 (N_223,In_265,In_339);
nor U224 (N_224,In_122,In_2455);
nor U225 (N_225,In_1604,N_80);
xor U226 (N_226,In_1359,In_1483);
xor U227 (N_227,In_2015,In_1238);
nand U228 (N_228,In_560,In_161);
nor U229 (N_229,In_2389,In_1721);
xnor U230 (N_230,In_693,In_1454);
or U231 (N_231,N_101,In_1710);
or U232 (N_232,In_18,In_1847);
and U233 (N_233,In_1175,In_145);
or U234 (N_234,In_1328,In_417);
nor U235 (N_235,In_2190,N_30);
and U236 (N_236,N_67,In_1648);
nand U237 (N_237,In_2364,In_1204);
nand U238 (N_238,In_144,In_2319);
nor U239 (N_239,In_1448,In_2336);
or U240 (N_240,In_2374,In_195);
xor U241 (N_241,In_750,In_7);
or U242 (N_242,In_221,In_2253);
nor U243 (N_243,In_573,In_510);
xor U244 (N_244,In_1383,In_1110);
nand U245 (N_245,In_532,In_775);
or U246 (N_246,In_689,In_1797);
or U247 (N_247,In_362,In_541);
or U248 (N_248,In_609,N_153);
xnor U249 (N_249,N_62,In_695);
nor U250 (N_250,In_2153,In_649);
and U251 (N_251,In_518,In_474);
xor U252 (N_252,In_2418,In_1679);
or U253 (N_253,In_1979,In_1009);
xnor U254 (N_254,In_507,In_1895);
xor U255 (N_255,In_1014,In_1830);
nor U256 (N_256,In_763,In_1498);
xnor U257 (N_257,In_356,In_2056);
and U258 (N_258,In_2356,In_1539);
or U259 (N_259,In_243,In_1769);
nand U260 (N_260,In_1715,N_192);
nor U261 (N_261,In_367,In_1759);
nand U262 (N_262,In_1613,In_2269);
or U263 (N_263,In_2100,In_845);
and U264 (N_264,In_1792,In_793);
nand U265 (N_265,In_1126,In_1342);
nor U266 (N_266,In_1372,In_2354);
xor U267 (N_267,In_965,In_1419);
and U268 (N_268,In_606,In_1526);
nor U269 (N_269,In_1670,In_2118);
and U270 (N_270,N_178,In_2246);
nand U271 (N_271,In_453,In_1225);
nor U272 (N_272,In_1534,In_176);
xnor U273 (N_273,In_1216,In_973);
and U274 (N_274,In_995,In_2178);
xnor U275 (N_275,In_1121,In_1964);
nand U276 (N_276,In_1149,In_737);
or U277 (N_277,In_1820,In_304);
or U278 (N_278,In_488,In_769);
nand U279 (N_279,In_1140,In_73);
nor U280 (N_280,In_38,In_861);
or U281 (N_281,In_1510,In_1701);
nand U282 (N_282,In_208,In_1322);
nand U283 (N_283,In_17,In_2166);
nor U284 (N_284,In_306,In_1938);
xor U285 (N_285,In_1177,In_2394);
xnor U286 (N_286,In_2129,N_149);
and U287 (N_287,In_2452,In_862);
or U288 (N_288,In_1931,In_1159);
and U289 (N_289,In_61,N_89);
xnor U290 (N_290,In_1537,In_661);
and U291 (N_291,In_214,In_219);
nand U292 (N_292,In_2385,In_944);
and U293 (N_293,In_651,N_83);
nor U294 (N_294,In_582,In_1379);
nand U295 (N_295,In_1450,In_2072);
or U296 (N_296,N_78,In_1885);
nand U297 (N_297,In_324,In_821);
xnor U298 (N_298,N_106,In_1947);
nor U299 (N_299,In_1054,In_1444);
nor U300 (N_300,In_733,In_564);
and U301 (N_301,In_2474,In_1031);
xor U302 (N_302,In_72,In_1584);
and U303 (N_303,In_901,In_70);
nor U304 (N_304,In_1092,In_1664);
or U305 (N_305,In_2361,In_1565);
nor U306 (N_306,In_426,In_1476);
xnor U307 (N_307,In_2390,In_956);
or U308 (N_308,N_20,In_1929);
xnor U309 (N_309,In_2273,N_45);
or U310 (N_310,In_130,In_2468);
nor U311 (N_311,In_1289,In_945);
xnor U312 (N_312,In_1723,In_260);
nand U313 (N_313,In_1407,In_1237);
nand U314 (N_314,In_991,In_1415);
or U315 (N_315,In_818,In_963);
nor U316 (N_316,In_2159,In_2185);
or U317 (N_317,In_1479,In_1197);
nand U318 (N_318,In_333,In_128);
nor U319 (N_319,N_168,In_2176);
nand U320 (N_320,In_2288,N_154);
xor U321 (N_321,N_88,In_547);
and U322 (N_322,In_1057,In_1249);
nor U323 (N_323,In_1324,In_707);
nand U324 (N_324,In_1902,In_892);
and U325 (N_325,In_1754,In_487);
and U326 (N_326,In_1631,N_97);
or U327 (N_327,In_1264,In_1970);
or U328 (N_328,In_209,In_1142);
or U329 (N_329,In_758,In_1202);
and U330 (N_330,In_943,In_2057);
nand U331 (N_331,In_1465,In_1432);
or U332 (N_332,In_727,In_1434);
nand U333 (N_333,In_688,In_559);
nand U334 (N_334,In_1120,In_2359);
nor U335 (N_335,N_199,In_593);
nor U336 (N_336,In_316,N_100);
nor U337 (N_337,In_565,N_61);
nor U338 (N_338,In_5,In_2033);
and U339 (N_339,In_2487,In_2041);
and U340 (N_340,In_2211,In_135);
xor U341 (N_341,In_2127,In_1049);
nor U342 (N_342,In_46,In_2352);
nand U343 (N_343,In_511,In_1962);
and U344 (N_344,In_52,In_1578);
and U345 (N_345,In_1876,In_1240);
or U346 (N_346,In_2204,In_164);
xor U347 (N_347,In_48,In_505);
and U348 (N_348,In_2274,In_279);
or U349 (N_349,In_1722,In_831);
nor U350 (N_350,In_1320,In_263);
and U351 (N_351,In_1285,In_897);
xnor U352 (N_352,In_681,In_2060);
or U353 (N_353,In_1662,N_4);
nand U354 (N_354,In_1082,In_74);
xnor U355 (N_355,In_1171,In_2165);
nand U356 (N_356,In_197,In_694);
nor U357 (N_357,In_1794,In_454);
xnor U358 (N_358,In_1341,In_1380);
nor U359 (N_359,In_28,In_2415);
or U360 (N_360,N_105,In_1816);
nand U361 (N_361,In_1994,In_1538);
xor U362 (N_362,In_1853,In_2480);
nor U363 (N_363,In_2262,In_1480);
xor U364 (N_364,In_1747,In_1354);
nand U365 (N_365,In_327,In_516);
and U366 (N_366,In_235,In_1826);
nand U367 (N_367,In_2071,In_668);
and U368 (N_368,In_1178,In_1780);
nor U369 (N_369,In_1520,In_1209);
or U370 (N_370,In_1349,In_2380);
nand U371 (N_371,In_1109,In_699);
xor U372 (N_372,In_2247,In_2440);
and U373 (N_373,In_538,In_2236);
nand U374 (N_374,In_413,In_2089);
nand U375 (N_375,In_2308,In_684);
and U376 (N_376,In_231,In_1946);
xnor U377 (N_377,In_163,In_633);
or U378 (N_378,In_1129,In_601);
nand U379 (N_379,In_2376,In_1412);
or U380 (N_380,In_1263,In_2463);
xnor U381 (N_381,N_161,In_986);
or U382 (N_382,In_57,In_1823);
nand U383 (N_383,In_2164,In_92);
nor U384 (N_384,In_171,In_95);
or U385 (N_385,In_1500,In_726);
and U386 (N_386,N_5,In_1303);
nand U387 (N_387,N_174,In_925);
or U388 (N_388,N_91,In_253);
or U389 (N_389,In_1073,In_930);
or U390 (N_390,In_2321,In_1030);
and U391 (N_391,In_2126,In_2342);
nor U392 (N_392,In_800,In_2407);
nand U393 (N_393,In_614,In_473);
nand U394 (N_394,In_1420,In_1442);
nor U395 (N_395,In_828,N_55);
nor U396 (N_396,In_931,In_834);
and U397 (N_397,In_80,N_32);
nor U398 (N_398,In_1926,In_251);
nor U399 (N_399,In_331,In_2358);
and U400 (N_400,In_1386,In_1609);
xnor U401 (N_401,In_1541,In_281);
and U402 (N_402,N_96,In_1398);
xor U403 (N_403,In_645,In_1837);
and U404 (N_404,In_824,In_1713);
nor U405 (N_405,N_59,N_217);
nand U406 (N_406,In_1261,In_1984);
or U407 (N_407,In_803,N_163);
or U408 (N_408,In_1977,N_111);
xnor U409 (N_409,In_272,In_1027);
nor U410 (N_410,N_276,N_297);
and U411 (N_411,In_1605,N_294);
nor U412 (N_412,In_2401,In_186);
or U413 (N_413,In_2331,In_312);
and U414 (N_414,In_1687,In_1768);
xnor U415 (N_415,In_2228,In_155);
and U416 (N_416,In_712,In_530);
xnor U417 (N_417,In_2235,In_1000);
and U418 (N_418,In_245,In_522);
xnor U419 (N_419,In_1692,In_2163);
nand U420 (N_420,In_1332,In_1458);
and U421 (N_421,In_829,In_2315);
nand U422 (N_422,In_206,In_2282);
nor U423 (N_423,In_172,In_1033);
and U424 (N_424,In_1559,In_2428);
nand U425 (N_425,In_1417,In_211);
xnor U426 (N_426,In_1854,In_2101);
nor U427 (N_427,In_400,N_359);
nand U428 (N_428,In_924,In_880);
xor U429 (N_429,In_1019,In_390);
or U430 (N_430,In_1653,In_2299);
and U431 (N_431,In_2123,In_625);
nand U432 (N_432,In_2349,In_470);
or U433 (N_433,In_1295,N_390);
or U434 (N_434,In_851,N_315);
nor U435 (N_435,In_1208,In_785);
nor U436 (N_436,In_2082,N_104);
or U437 (N_437,In_1900,N_179);
or U438 (N_438,In_1011,N_397);
and U439 (N_439,N_295,N_44);
xor U440 (N_440,In_2151,In_127);
nor U441 (N_441,N_303,In_1084);
nor U442 (N_442,In_1672,In_1657);
or U443 (N_443,In_1048,In_777);
or U444 (N_444,In_1452,In_2195);
and U445 (N_445,In_2466,N_74);
xnor U446 (N_446,N_300,In_1728);
and U447 (N_447,In_2156,In_296);
or U448 (N_448,In_169,In_743);
and U449 (N_449,In_1727,In_812);
or U450 (N_450,In_957,In_1135);
xnor U451 (N_451,In_1522,In_1891);
xor U452 (N_452,In_2485,N_129);
nand U453 (N_453,In_1967,In_947);
and U454 (N_454,In_2275,In_1366);
and U455 (N_455,In_1421,In_1944);
xor U456 (N_456,In_940,In_183);
and U457 (N_457,In_586,In_1509);
nor U458 (N_458,In_2261,In_718);
and U459 (N_459,In_837,In_1302);
and U460 (N_460,N_47,In_2097);
and U461 (N_461,In_2192,In_2362);
and U462 (N_462,In_1930,In_1973);
nor U463 (N_463,In_2121,In_450);
nand U464 (N_464,In_227,In_2360);
or U465 (N_465,In_1922,In_258);
or U466 (N_466,In_354,In_93);
nand U467 (N_467,In_1896,In_1003);
and U468 (N_468,In_410,N_220);
xor U469 (N_469,In_1244,In_1992);
and U470 (N_470,In_1925,N_254);
xor U471 (N_471,N_257,In_698);
or U472 (N_472,In_809,In_2387);
and U473 (N_473,In_485,In_754);
nor U474 (N_474,In_1377,N_248);
nand U475 (N_475,In_242,In_2449);
xor U476 (N_476,In_958,In_959);
and U477 (N_477,In_461,N_326);
xor U478 (N_478,N_85,In_1607);
or U479 (N_479,N_348,In_2432);
nand U480 (N_480,In_993,In_2081);
xnor U481 (N_481,In_232,In_177);
or U482 (N_482,In_2471,In_962);
xnor U483 (N_483,In_580,In_1551);
and U484 (N_484,In_1381,In_10);
xnor U485 (N_485,In_141,In_1603);
and U486 (N_486,N_127,In_364);
nor U487 (N_487,In_2481,In_388);
or U488 (N_488,In_846,In_2341);
xnor U489 (N_489,In_882,In_1636);
xnor U490 (N_490,In_1935,N_235);
xnor U491 (N_491,In_705,N_259);
or U492 (N_492,In_1867,N_350);
and U493 (N_493,In_2307,In_289);
and U494 (N_494,In_2091,In_676);
xor U495 (N_495,N_293,In_692);
nand U496 (N_496,In_667,In_154);
and U497 (N_497,N_394,In_1195);
and U498 (N_498,In_2222,In_910);
xor U499 (N_499,In_1963,In_891);
nor U500 (N_500,In_1214,N_15);
and U501 (N_501,In_303,In_1267);
or U502 (N_502,In_2384,In_380);
nand U503 (N_503,In_496,In_546);
and U504 (N_504,In_1305,In_1774);
and U505 (N_505,In_178,In_1212);
nand U506 (N_506,In_960,N_169);
nand U507 (N_507,In_224,In_1331);
xor U508 (N_508,In_2458,In_1223);
and U509 (N_509,N_165,N_382);
or U510 (N_510,In_545,In_1194);
and U511 (N_511,In_802,N_281);
xor U512 (N_512,In_842,In_1314);
nand U513 (N_513,In_1360,In_2186);
xor U514 (N_514,In_2037,In_1215);
nor U515 (N_515,In_2227,N_214);
and U516 (N_516,N_279,In_696);
xor U517 (N_517,N_312,In_840);
nor U518 (N_518,N_274,In_1257);
xnor U519 (N_519,In_96,In_1700);
or U520 (N_520,In_1181,In_329);
nand U521 (N_521,In_1008,In_961);
xor U522 (N_522,In_1358,In_0);
or U523 (N_523,In_266,In_2244);
and U524 (N_524,In_187,N_113);
nor U525 (N_525,In_283,In_1750);
or U526 (N_526,In_797,In_1394);
xor U527 (N_527,In_414,In_317);
nor U528 (N_528,In_268,In_22);
or U529 (N_529,In_2138,In_2338);
nand U530 (N_530,In_753,In_406);
xnor U531 (N_531,In_905,In_1532);
xor U532 (N_532,In_250,In_2219);
nand U533 (N_533,In_1006,In_340);
nand U534 (N_534,In_2489,In_1410);
nor U535 (N_535,N_112,In_3);
nor U536 (N_536,N_6,N_2);
nand U537 (N_537,In_662,In_1844);
nor U538 (N_538,In_1587,In_885);
nor U539 (N_539,In_203,N_366);
nor U540 (N_540,In_2024,In_1832);
and U541 (N_541,In_996,In_1628);
or U542 (N_542,In_2251,In_1528);
or U543 (N_543,In_719,In_556);
nand U544 (N_544,In_1554,In_1042);
nor U545 (N_545,In_1801,In_1319);
xor U546 (N_546,In_2447,In_2027);
nand U547 (N_547,In_1872,In_1400);
nor U548 (N_548,In_500,In_150);
nor U549 (N_549,N_159,In_1800);
or U550 (N_550,In_156,N_56);
nor U551 (N_551,In_2411,In_1441);
xnor U552 (N_552,N_72,In_248);
nor U553 (N_553,In_1230,In_1858);
or U554 (N_554,In_1064,In_2239);
nand U555 (N_555,In_2050,In_2333);
nor U556 (N_556,In_1749,In_1067);
xor U557 (N_557,In_1650,In_56);
and U558 (N_558,In_2196,In_1242);
nor U559 (N_559,In_735,In_1200);
or U560 (N_560,In_2238,In_1918);
nor U561 (N_561,In_76,In_167);
or U562 (N_562,In_2476,N_336);
or U563 (N_563,In_833,In_1937);
nand U564 (N_564,N_160,N_204);
and U565 (N_565,In_107,In_126);
and U566 (N_566,N_189,In_2009);
and U567 (N_567,In_1467,In_2300);
nor U568 (N_568,In_794,In_2114);
or U569 (N_569,In_1158,In_2266);
nor U570 (N_570,In_1996,N_12);
nor U571 (N_571,In_2169,In_1164);
and U572 (N_572,In_2002,In_841);
nor U573 (N_573,In_639,In_1684);
nand U574 (N_574,In_1742,In_21);
xnor U575 (N_575,In_2409,In_351);
nor U576 (N_576,N_263,N_65);
or U577 (N_577,In_100,In_1806);
nor U578 (N_578,In_1486,N_216);
or U579 (N_579,In_71,In_110);
nand U580 (N_580,In_1694,N_256);
and U581 (N_581,In_412,In_466);
nor U582 (N_582,In_971,In_1066);
nor U583 (N_583,In_2245,In_832);
and U584 (N_584,In_1160,In_1645);
xnor U585 (N_585,In_2486,In_1873);
nor U586 (N_586,In_739,In_1590);
xor U587 (N_587,In_2168,In_1849);
xnor U588 (N_588,N_115,In_760);
and U589 (N_589,In_2309,In_1758);
and U590 (N_590,N_398,In_1141);
xnor U591 (N_591,In_2403,In_2365);
or U592 (N_592,In_1596,In_2283);
xor U593 (N_593,In_1732,In_1730);
xor U594 (N_594,In_2026,In_2353);
nand U595 (N_595,In_2343,In_2231);
xnor U596 (N_596,In_2305,In_2131);
xor U597 (N_597,In_920,In_202);
or U598 (N_598,In_184,In_1327);
xnor U599 (N_599,In_1919,In_1920);
nor U600 (N_600,In_2272,In_1699);
nand U601 (N_601,In_1775,In_2416);
and U602 (N_602,In_482,In_987);
and U603 (N_603,In_1910,In_1888);
and U604 (N_604,In_2073,In_1886);
nor U605 (N_605,In_830,In_1668);
and U606 (N_606,N_108,In_136);
or U607 (N_607,N_182,In_2044);
nor U608 (N_608,N_565,In_225);
xor U609 (N_609,In_1139,N_242);
and U610 (N_610,N_476,In_682);
nand U611 (N_611,In_1235,In_1485);
or U612 (N_612,N_207,N_7);
and U613 (N_613,In_526,In_2417);
nand U614 (N_614,In_2293,N_132);
or U615 (N_615,In_498,N_213);
or U616 (N_616,N_226,N_241);
and U617 (N_617,In_782,In_778);
xnor U618 (N_618,In_2070,In_117);
nand U619 (N_619,In_913,In_1321);
nor U620 (N_620,In_1870,In_932);
or U621 (N_621,In_2200,In_428);
or U622 (N_622,In_1134,In_1205);
xnor U623 (N_623,In_2061,In_2439);
and U624 (N_624,In_2183,N_578);
xnor U625 (N_625,N_320,N_227);
or U626 (N_626,In_1179,In_1548);
nor U627 (N_627,In_2386,In_1446);
nand U628 (N_628,In_1737,In_293);
or U629 (N_629,N_511,N_252);
or U630 (N_630,In_1023,N_285);
and U631 (N_631,In_1610,In_431);
nand U632 (N_632,In_394,N_441);
nand U633 (N_633,In_2497,In_1229);
or U634 (N_634,In_740,In_1770);
nand U635 (N_635,In_1640,N_531);
nor U636 (N_636,In_1490,N_313);
xnor U637 (N_637,In_342,In_1294);
or U638 (N_638,N_555,In_2313);
nand U639 (N_639,In_44,N_8);
nor U640 (N_640,In_2198,N_210);
nor U641 (N_641,In_847,In_1851);
nand U642 (N_642,In_1709,In_2295);
or U643 (N_643,In_536,In_1995);
nor U644 (N_644,In_430,In_1731);
nand U645 (N_645,In_539,In_1651);
nand U646 (N_646,In_1098,N_166);
nand U647 (N_647,In_1459,In_2145);
nor U648 (N_648,In_2035,In_2080);
and U649 (N_649,In_1560,N_423);
or U650 (N_650,In_139,In_1864);
nor U651 (N_651,N_304,N_465);
or U652 (N_652,In_1845,In_2294);
nor U653 (N_653,In_173,N_595);
nor U654 (N_654,In_1113,In_630);
or U655 (N_655,In_249,N_575);
xor U656 (N_656,N_583,In_157);
nor U657 (N_657,In_168,N_19);
or U658 (N_658,In_1392,In_900);
and U659 (N_659,In_2068,In_1071);
xor U660 (N_660,In_524,In_2157);
and U661 (N_661,In_1976,In_1720);
nand U662 (N_662,N_121,In_627);
nand U663 (N_663,In_687,In_881);
nand U664 (N_664,In_373,N_334);
nor U665 (N_665,N_272,In_440);
nand U666 (N_666,N_401,N_228);
nand U667 (N_667,In_165,N_515);
or U668 (N_668,In_313,N_434);
nand U669 (N_669,In_2135,In_566);
nor U670 (N_670,In_2143,N_299);
and U671 (N_671,In_383,In_1743);
or U672 (N_672,In_1663,In_1494);
nor U673 (N_673,N_208,In_55);
nor U674 (N_674,N_292,In_1907);
xor U675 (N_675,N_338,N_411);
nand U676 (N_676,In_1796,In_2098);
nand U677 (N_677,In_252,In_1233);
or U678 (N_678,N_448,In_2377);
or U679 (N_679,N_314,In_1304);
nand U680 (N_680,In_1639,In_69);
and U681 (N_681,N_215,In_382);
and U682 (N_682,In_1669,In_192);
and U683 (N_683,In_437,In_679);
and U684 (N_684,In_421,In_1492);
nor U685 (N_685,N_145,In_273);
xnor U686 (N_686,In_1250,In_1367);
and U687 (N_687,In_153,N_466);
and U688 (N_688,In_1884,N_184);
or U689 (N_689,In_2048,N_521);
xor U690 (N_690,In_610,In_2435);
xnor U691 (N_691,N_49,N_54);
and U692 (N_692,In_1187,In_1583);
xor U693 (N_693,In_1255,In_751);
and U694 (N_694,In_657,N_580);
or U695 (N_695,In_1878,In_1271);
and U696 (N_696,In_501,N_358);
and U697 (N_697,In_477,N_233);
xor U698 (N_698,N_1,N_477);
nand U699 (N_699,In_463,In_1496);
nand U700 (N_700,N_288,In_2132);
and U701 (N_701,In_1234,N_193);
nor U702 (N_702,In_795,In_375);
and U703 (N_703,In_1222,In_2477);
and U704 (N_704,N_267,In_2124);
or U705 (N_705,In_1365,In_836);
and U706 (N_706,N_291,In_1070);
xor U707 (N_707,N_34,In_1183);
nand U708 (N_708,In_588,In_1788);
and U709 (N_709,In_587,N_138);
nand U710 (N_710,In_508,In_86);
and U711 (N_711,N_135,In_2173);
nor U712 (N_712,N_391,In_2460);
nand U713 (N_713,In_2046,In_1282);
nand U714 (N_714,In_1017,In_2214);
xnor U715 (N_715,In_2482,In_2001);
nand U716 (N_716,In_1231,In_2478);
nand U717 (N_717,N_414,In_529);
nor U718 (N_718,In_1777,In_1290);
nor U719 (N_719,In_1456,N_144);
or U720 (N_720,In_1751,In_448);
xor U721 (N_721,In_1276,N_33);
nor U722 (N_722,In_857,In_734);
nor U723 (N_723,In_2470,In_1617);
nand U724 (N_724,In_874,In_2155);
nand U725 (N_725,In_2158,In_1147);
nor U726 (N_726,In_1218,In_449);
or U727 (N_727,N_86,N_481);
xnor U728 (N_728,In_792,In_318);
xnor U729 (N_729,In_2265,In_648);
xor U730 (N_730,In_1882,In_2496);
xor U731 (N_731,In_1445,In_15);
or U732 (N_732,In_1624,In_2453);
or U733 (N_733,In_2226,In_2220);
and U734 (N_734,N_539,In_166);
nand U735 (N_735,In_2312,In_321);
xor U736 (N_736,N_231,In_65);
nand U737 (N_737,In_386,In_1162);
or U738 (N_738,In_1495,In_513);
nand U739 (N_739,N_377,In_563);
nand U740 (N_740,In_721,In_1193);
nand U741 (N_741,In_2414,In_608);
nand U742 (N_742,In_951,In_292);
nor U743 (N_743,N_581,In_2193);
nand U744 (N_744,In_643,In_350);
nor U745 (N_745,In_1345,N_373);
nand U746 (N_746,In_744,N_553);
and U747 (N_747,In_1313,N_495);
and U748 (N_748,In_14,In_915);
or U749 (N_749,In_2303,N_124);
xor U750 (N_750,N_318,N_187);
nor U751 (N_751,In_1173,In_1784);
nor U752 (N_752,In_497,In_1600);
nor U753 (N_753,N_428,In_2086);
and U754 (N_754,In_1683,In_2013);
or U755 (N_755,In_2034,N_130);
xnor U756 (N_756,In_468,In_1300);
and U757 (N_757,In_929,In_1156);
xor U758 (N_758,In_1546,In_642);
xnor U759 (N_759,In_1561,In_33);
nor U760 (N_760,In_1622,In_229);
nand U761 (N_761,N_90,In_54);
nor U762 (N_762,N_363,N_64);
xnor U763 (N_763,In_1152,N_277);
or U764 (N_764,In_1382,In_551);
or U765 (N_765,In_1063,N_381);
nand U766 (N_766,N_346,In_2221);
and U767 (N_767,In_1041,N_410);
nand U768 (N_768,In_1729,In_1674);
nor U769 (N_769,N_369,N_508);
or U770 (N_770,In_1736,In_1766);
nor U771 (N_771,N_492,In_2154);
or U772 (N_772,N_497,In_1988);
and U773 (N_773,In_1632,In_503);
xnor U774 (N_774,In_2069,In_2499);
or U775 (N_775,In_1453,In_1385);
or U776 (N_776,In_759,N_408);
nand U777 (N_777,In_981,In_287);
or U778 (N_778,In_2215,In_1616);
and U779 (N_779,In_1122,In_720);
nor U780 (N_780,In_1266,In_2405);
nor U781 (N_781,In_984,In_1130);
and U782 (N_782,N_430,In_1827);
or U783 (N_783,In_1734,In_756);
nor U784 (N_784,In_1983,N_335);
and U785 (N_785,N_562,N_475);
nor U786 (N_786,In_1236,In_2278);
nor U787 (N_787,In_1422,N_589);
or U788 (N_788,In_2191,In_1457);
or U789 (N_789,In_338,N_446);
nand U790 (N_790,In_1576,In_1081);
nor U791 (N_791,In_2150,In_2311);
nand U792 (N_792,In_2328,N_286);
nand U793 (N_793,In_424,N_478);
nand U794 (N_794,N_546,In_2177);
nor U795 (N_795,N_404,N_339);
and U796 (N_796,In_1413,N_224);
and U797 (N_797,N_230,N_523);
and U798 (N_798,N_137,In_1874);
or U799 (N_799,In_1491,In_115);
xnor U800 (N_800,In_1843,N_379);
and U801 (N_801,N_711,In_298);
nor U802 (N_802,N_316,N_650);
nor U803 (N_803,N_548,In_817);
and U804 (N_804,N_729,N_616);
nand U805 (N_805,N_400,N_399);
or U806 (N_806,In_1090,In_592);
nand U807 (N_807,N_632,N_721);
and U808 (N_808,In_671,N_460);
or U809 (N_809,In_686,In_1269);
nand U810 (N_810,In_942,In_2324);
nand U811 (N_811,In_2381,N_413);
xor U812 (N_812,In_310,N_775);
nor U813 (N_813,In_361,In_2199);
nand U814 (N_814,In_1036,In_1773);
xnor U815 (N_815,In_323,N_795);
xnor U816 (N_816,N_31,In_670);
or U817 (N_817,N_150,In_853);
or U818 (N_818,In_1206,In_1403);
xnor U819 (N_819,In_89,In_2028);
nand U820 (N_820,N_790,N_668);
or U821 (N_821,In_2213,In_2368);
nand U822 (N_822,In_1623,In_1591);
xnor U823 (N_823,In_1323,N_143);
nand U824 (N_824,In_1032,N_58);
nand U825 (N_825,In_1698,N_456);
nand U826 (N_826,In_804,In_2162);
and U827 (N_827,In_1226,In_299);
and U828 (N_828,In_484,In_2350);
and U829 (N_829,N_225,In_860);
or U830 (N_830,In_322,In_883);
nand U831 (N_831,In_2423,In_389);
xnor U832 (N_832,In_1595,N_71);
and U833 (N_833,In_906,In_387);
or U834 (N_834,In_1658,In_160);
nor U835 (N_835,In_1836,N_13);
nor U836 (N_836,In_591,In_1397);
nor U837 (N_837,In_2472,In_1039);
xnor U838 (N_838,In_1940,N_374);
and U839 (N_839,N_579,In_1575);
xor U840 (N_840,In_806,In_2241);
nor U841 (N_841,In_1005,In_711);
nand U842 (N_842,N_436,In_1137);
or U843 (N_843,N_35,In_1497);
and U844 (N_844,N_70,In_1462);
nor U845 (N_845,In_1790,In_997);
nor U846 (N_846,N_550,N_648);
and U847 (N_847,In_2443,In_1254);
or U848 (N_848,In_1253,N_21);
nand U849 (N_849,In_660,N_158);
or U850 (N_850,In_728,In_2259);
or U851 (N_851,In_343,In_1566);
xor U852 (N_852,In_1932,In_1990);
xor U853 (N_853,In_1246,In_531);
nor U854 (N_854,N_509,N_461);
or U855 (N_855,N_99,In_1956);
and U856 (N_856,In_1038,In_521);
nand U857 (N_857,In_1093,In_40);
or U858 (N_858,In_146,In_1102);
nand U859 (N_859,In_255,N_619);
or U860 (N_860,In_1748,In_1361);
or U861 (N_861,In_458,N_43);
or U862 (N_862,In_1350,N_38);
xor U863 (N_863,In_807,In_1634);
or U864 (N_864,In_561,In_2457);
nand U865 (N_865,N_46,In_1065);
xnor U866 (N_866,In_210,In_441);
or U867 (N_867,In_1521,In_472);
xor U868 (N_868,In_1338,N_333);
nor U869 (N_869,N_666,In_1335);
or U870 (N_870,N_688,N_710);
and U871 (N_871,In_300,N_596);
nor U872 (N_872,In_67,N_439);
nor U873 (N_873,N_747,N_637);
nand U874 (N_874,N_560,N_375);
nor U875 (N_875,N_141,N_652);
or U876 (N_876,In_385,N_758);
xnor U877 (N_877,N_499,In_2085);
xor U878 (N_878,N_679,N_754);
and U879 (N_879,N_368,In_1726);
nand U880 (N_880,In_884,In_97);
nand U881 (N_881,N_689,In_663);
and U882 (N_882,In_2436,In_923);
nor U883 (N_883,N_357,N_457);
nand U884 (N_884,In_2029,N_664);
and U885 (N_885,N_114,In_848);
xnor U886 (N_886,In_1879,In_365);
xnor U887 (N_887,In_1778,In_79);
xor U888 (N_888,In_26,In_1248);
xnor U889 (N_889,N_622,In_1503);
and U890 (N_890,N_574,In_730);
and U891 (N_891,In_334,In_1405);
xnor U892 (N_892,In_852,N_667);
or U893 (N_893,In_1283,In_936);
or U894 (N_894,N_755,In_1330);
nand U895 (N_895,N_693,In_2240);
xnor U896 (N_896,In_1273,N_380);
or U897 (N_897,In_755,In_1906);
nor U898 (N_898,In_2433,In_2023);
or U899 (N_899,N_612,In_1291);
nor U900 (N_900,In_825,N_424);
xnor U901 (N_901,N_792,In_181);
or U902 (N_902,N_324,In_977);
or U903 (N_903,N_392,In_1101);
or U904 (N_904,In_45,N_512);
nand U905 (N_905,In_1939,In_319);
xor U906 (N_906,In_2290,In_859);
xor U907 (N_907,In_1618,In_1516);
xnor U908 (N_908,In_899,In_35);
and U909 (N_909,In_1838,In_282);
or U910 (N_910,In_1133,In_509);
or U911 (N_911,In_1557,In_182);
xnor U912 (N_912,In_2318,In_766);
nor U913 (N_913,In_347,In_1435);
and U914 (N_914,N_432,In_1277);
nand U915 (N_915,N_682,N_331);
or U916 (N_916,In_13,In_1544);
nor U917 (N_917,N_633,N_791);
and U918 (N_918,N_566,N_654);
and U919 (N_919,N_606,In_1035);
nor U920 (N_920,In_826,In_20);
and U921 (N_921,In_1746,In_1782);
or U922 (N_922,In_2120,N_534);
nand U923 (N_923,In_2445,In_616);
nand U924 (N_924,N_42,In_599);
and U925 (N_925,In_2088,In_2000);
nand U926 (N_926,N_704,N_734);
or U927 (N_927,In_1654,N_493);
and U928 (N_928,N_745,In_2329);
xor U929 (N_929,In_723,In_1489);
or U930 (N_930,N_490,In_761);
nor U931 (N_931,In_656,In_1104);
nor U932 (N_932,In_201,In_1647);
nand U933 (N_933,In_435,In_659);
or U934 (N_934,In_1828,In_2264);
nor U935 (N_935,N_341,N_780);
and U936 (N_936,In_1015,In_1540);
nor U937 (N_937,In_1708,In_31);
or U938 (N_938,In_918,In_2031);
or U939 (N_939,In_1821,In_1652);
xor U940 (N_940,In_2136,In_1833);
nor U941 (N_941,N_395,In_276);
nor U942 (N_942,N_325,N_356);
nand U943 (N_943,N_222,In_1860);
xor U944 (N_944,In_514,N_715);
and U945 (N_945,N_94,In_669);
nand U946 (N_946,In_355,In_1804);
nand U947 (N_947,In_1184,In_1911);
and U948 (N_948,N_544,In_2051);
xor U949 (N_949,N_670,In_985);
xor U950 (N_950,In_717,In_1719);
nor U951 (N_951,In_701,N_376);
xor U952 (N_952,In_1518,N_706);
xnor U953 (N_953,In_2393,N_699);
nor U954 (N_954,In_619,In_1985);
nor U955 (N_955,In_2036,In_1118);
xor U956 (N_956,N_195,In_1060);
nor U957 (N_957,In_2011,In_1245);
nand U958 (N_958,N_530,In_1993);
and U959 (N_959,In_603,N_445);
and U960 (N_960,N_568,N_156);
and U961 (N_961,In_908,In_644);
xnor U962 (N_962,N_587,N_351);
xnor U963 (N_963,In_256,In_2233);
or U964 (N_964,N_205,In_1917);
and U965 (N_965,In_1127,In_1364);
nand U966 (N_966,N_79,In_1877);
nand U967 (N_967,N_776,In_879);
nand U968 (N_968,N_784,In_955);
or U969 (N_969,In_715,In_1786);
and U970 (N_970,N_396,In_2032);
and U971 (N_971,In_1301,In_938);
and U972 (N_972,In_553,N_799);
nand U973 (N_973,In_1968,In_1198);
nand U974 (N_974,N_655,In_275);
and U975 (N_975,In_170,In_1642);
or U976 (N_976,In_2160,In_2424);
xor U977 (N_977,In_1241,In_204);
nand U978 (N_978,N_122,N_151);
nor U979 (N_979,In_2203,N_723);
xor U980 (N_980,In_288,N_720);
nor U981 (N_981,N_147,In_330);
and U982 (N_982,In_2212,N_232);
and U983 (N_983,In_2042,N_540);
nand U984 (N_984,N_438,N_642);
or U985 (N_985,In_638,In_234);
nand U986 (N_986,In_2019,In_280);
nand U987 (N_987,N_777,In_2320);
or U988 (N_988,N_384,In_1018);
nand U989 (N_989,In_2479,In_1340);
and U990 (N_990,In_1572,In_193);
xnor U991 (N_991,N_234,In_402);
nor U992 (N_992,In_1268,In_1545);
nand U993 (N_993,In_1689,In_1752);
nand U994 (N_994,In_623,N_455);
and U995 (N_995,In_1424,In_1989);
nand U996 (N_996,In_2419,N_532);
nand U997 (N_997,In_1199,In_457);
nand U998 (N_998,In_1529,In_1834);
and U999 (N_999,N_332,N_177);
nand U1000 (N_1000,In_1308,N_525);
or U1001 (N_1001,In_1262,In_134);
and U1002 (N_1002,In_1451,In_159);
or U1003 (N_1003,In_262,In_1176);
and U1004 (N_1004,In_1688,In_381);
nor U1005 (N_1005,N_95,In_1278);
nor U1006 (N_1006,N_601,N_317);
nand U1007 (N_1007,In_811,In_1336);
and U1008 (N_1008,N_522,In_1471);
nand U1009 (N_1009,N_81,In_2076);
and U1010 (N_1010,N_269,In_2327);
nand U1011 (N_1011,In_655,In_1185);
nand U1012 (N_1012,N_916,In_2279);
xor U1013 (N_1013,N_772,In_1577);
xor U1014 (N_1014,In_2148,N_278);
xnor U1015 (N_1015,In_1166,N_571);
xor U1016 (N_1016,In_2179,N_963);
and U1017 (N_1017,N_327,In_597);
xnor U1018 (N_1018,N_593,N_815);
xor U1019 (N_1019,N_761,In_729);
or U1020 (N_1020,In_493,In_1085);
nand U1021 (N_1021,N_789,N_942);
and U1022 (N_1022,In_2406,In_2473);
nand U1023 (N_1023,In_1123,In_2412);
xor U1024 (N_1024,N_898,N_63);
nor U1025 (N_1025,N_724,N_561);
and U1026 (N_1026,N_806,N_503);
and U1027 (N_1027,In_979,In_455);
and U1028 (N_1028,N_524,N_516);
and U1029 (N_1029,In_1997,In_927);
nand U1030 (N_1030,In_1725,In_1718);
nand U1031 (N_1031,N_841,In_1889);
nand U1032 (N_1032,In_672,In_2106);
and U1033 (N_1033,In_904,N_282);
nand U1034 (N_1034,In_584,N_118);
or U1035 (N_1035,N_202,N_698);
and U1036 (N_1036,N_588,N_737);
nor U1037 (N_1037,In_1484,N_886);
or U1038 (N_1038,In_1306,N_984);
or U1039 (N_1039,In_2189,In_1131);
xnor U1040 (N_1040,In_702,N_211);
or U1041 (N_1041,N_196,N_301);
nor U1042 (N_1042,In_1807,In_980);
nor U1043 (N_1043,In_486,N_905);
and U1044 (N_1044,In_1852,In_1757);
or U1045 (N_1045,N_321,N_653);
and U1046 (N_1046,N_473,N_569);
and U1047 (N_1047,In_876,N_422);
xor U1048 (N_1048,N_329,In_2117);
nor U1049 (N_1049,In_762,In_506);
or U1050 (N_1050,N_635,In_1080);
nand U1051 (N_1051,In_558,N_762);
nand U1052 (N_1052,In_41,N_923);
xor U1053 (N_1053,N_922,In_1552);
nor U1054 (N_1054,In_2357,In_1661);
and U1055 (N_1055,In_1975,N_617);
nor U1056 (N_1056,In_1224,N_28);
or U1057 (N_1057,In_978,N_440);
nand U1058 (N_1058,In_620,In_2188);
xnor U1059 (N_1059,In_1318,In_748);
nand U1060 (N_1060,N_676,In_1431);
nand U1061 (N_1061,N_692,In_725);
xor U1062 (N_1062,In_2332,N_846);
xnor U1063 (N_1063,N_330,N_774);
nand U1064 (N_1064,N_549,In_216);
xor U1065 (N_1065,In_968,N_519);
nand U1066 (N_1066,N_802,N_874);
xor U1067 (N_1067,N_554,In_1515);
nand U1068 (N_1068,In_1904,In_2216);
nor U1069 (N_1069,N_444,N_973);
xor U1070 (N_1070,In_1629,N_866);
or U1071 (N_1071,N_406,N_935);
nand U1072 (N_1072,N_188,N_502);
nand U1073 (N_1073,In_632,In_1077);
or U1074 (N_1074,In_230,N_171);
xnor U1075 (N_1075,N_709,In_1339);
and U1076 (N_1076,N_305,In_1793);
nor U1077 (N_1077,In_1487,N_703);
nor U1078 (N_1078,In_363,N_117);
and U1079 (N_1079,N_822,In_1375);
nor U1080 (N_1080,In_710,In_416);
or U1081 (N_1081,In_215,N_491);
nor U1082 (N_1082,In_1690,N_966);
nand U1083 (N_1083,In_527,N_757);
nand U1084 (N_1084,In_896,In_2408);
and U1085 (N_1085,N_983,In_666);
xor U1086 (N_1086,N_887,N_832);
nor U1087 (N_1087,In_1763,In_914);
or U1088 (N_1088,In_1972,In_1601);
xor U1089 (N_1089,In_174,N_718);
and U1090 (N_1090,In_697,In_2025);
and U1091 (N_1091,In_2459,N_322);
nor U1092 (N_1092,N_513,N_547);
nand U1093 (N_1093,In_125,In_810);
or U1094 (N_1094,N_982,In_337);
xor U1095 (N_1095,In_1869,In_1707);
xor U1096 (N_1096,N_237,In_1865);
or U1097 (N_1097,In_137,In_1592);
xor U1098 (N_1098,N_268,In_2351);
or U1099 (N_1099,In_2323,N_639);
or U1100 (N_1100,N_337,In_2149);
or U1101 (N_1101,In_1099,N_749);
or U1102 (N_1102,In_2018,N_895);
xor U1103 (N_1103,In_567,N_603);
nand U1104 (N_1104,N_186,N_892);
or U1105 (N_1105,In_1619,In_1389);
and U1106 (N_1106,N_68,In_894);
nand U1107 (N_1107,In_844,N_783);
xor U1108 (N_1108,In_798,In_328);
nand U1109 (N_1109,N_148,In_1756);
and U1110 (N_1110,N_765,In_118);
and U1111 (N_1111,N_782,In_732);
nor U1112 (N_1112,In_2271,In_1280);
nor U1113 (N_1113,In_533,In_1103);
or U1114 (N_1114,N_930,In_1625);
or U1115 (N_1115,N_599,In_708);
nor U1116 (N_1116,N_636,In_396);
nor U1117 (N_1117,N_510,In_886);
nor U1118 (N_1118,In_2347,In_469);
nor U1119 (N_1119,In_2020,In_1221);
nor U1120 (N_1120,N_464,In_1376);
nand U1121 (N_1121,In_2243,N_681);
nand U1122 (N_1122,In_2105,In_1021);
xnor U1123 (N_1123,In_2469,N_591);
xnor U1124 (N_1124,N_538,In_1871);
nand U1125 (N_1125,N_393,N_728);
nand U1126 (N_1126,In_418,In_1107);
xor U1127 (N_1127,N_798,In_612);
xor U1128 (N_1128,In_916,N_740);
xor U1129 (N_1129,In_1088,In_2043);
nand U1130 (N_1130,In_890,N_958);
xnor U1131 (N_1131,N_201,In_2297);
xor U1132 (N_1132,In_113,N_14);
nor U1133 (N_1133,N_157,N_997);
and U1134 (N_1134,N_949,In_647);
or U1135 (N_1135,In_2064,In_543);
xor U1136 (N_1136,In_1402,N_500);
or U1137 (N_1137,N_823,In_2250);
and U1138 (N_1138,N_742,In_1251);
nand U1139 (N_1139,N_882,N_103);
nand U1140 (N_1140,N_736,In_87);
nand U1141 (N_1141,N_496,N_306);
nor U1142 (N_1142,In_1167,In_119);
or U1143 (N_1143,In_839,In_358);
xnor U1144 (N_1144,In_47,In_1633);
or U1145 (N_1145,In_1711,N_602);
nand U1146 (N_1146,N_727,N_656);
xnor U1147 (N_1147,N_976,N_767);
and U1148 (N_1148,N_378,N_200);
nor U1149 (N_1149,In_277,In_774);
xnor U1150 (N_1150,N_385,In_1037);
nor U1151 (N_1151,In_1585,In_731);
and U1152 (N_1152,In_1505,N_442);
nor U1153 (N_1153,In_2276,In_1059);
xor U1154 (N_1154,N_649,In_467);
nand U1155 (N_1155,N_751,In_2016);
xnor U1156 (N_1156,In_1165,N_469);
or U1157 (N_1157,N_311,In_2078);
nand U1158 (N_1158,In_138,N_435);
and U1159 (N_1159,In_267,N_701);
xnor U1160 (N_1160,In_983,In_101);
nor U1161 (N_1161,N_684,N_92);
nor U1162 (N_1162,In_2425,N_828);
xor U1163 (N_1163,In_747,N_861);
nand U1164 (N_1164,N_821,In_1499);
and U1165 (N_1165,N_941,In_2392);
and U1166 (N_1166,N_628,N_672);
nor U1167 (N_1167,In_37,N_273);
and U1168 (N_1168,In_779,In_907);
or U1169 (N_1169,N_825,In_709);
xor U1170 (N_1170,N_167,N_170);
xor U1171 (N_1171,N_934,In_690);
xor U1172 (N_1172,N_454,N_770);
or U1173 (N_1173,In_1957,In_2456);
or U1174 (N_1174,In_1597,N_506);
xnor U1175 (N_1175,N_944,In_345);
or U1176 (N_1176,N_911,In_2249);
and U1177 (N_1177,N_750,N_533);
and U1178 (N_1178,N_708,In_213);
or U1179 (N_1179,In_1739,N_936);
or U1180 (N_1180,In_1753,N_675);
nand U1181 (N_1181,N_134,N_819);
nor U1182 (N_1182,In_926,In_2289);
xnor U1183 (N_1183,In_1569,N_858);
or U1184 (N_1184,N_173,N_125);
xor U1185 (N_1185,N_529,In_2113);
nand U1186 (N_1186,In_1357,In_1010);
and U1187 (N_1187,N_155,N_618);
or U1188 (N_1188,N_778,In_401);
xnor U1189 (N_1189,N_808,In_1390);
nand U1190 (N_1190,In_738,In_1855);
xnor U1191 (N_1191,In_68,N_779);
nor U1192 (N_1192,In_2270,In_1293);
or U1193 (N_1193,In_471,In_395);
and U1194 (N_1194,In_1862,In_415);
and U1195 (N_1195,N_426,In_1921);
nand U1196 (N_1196,In_1013,N_697);
xnor U1197 (N_1197,In_1296,In_2263);
nand U1198 (N_1198,N_884,N_484);
and U1199 (N_1199,N_812,In_1016);
nor U1200 (N_1200,N_471,N_76);
nor U1201 (N_1201,N_1105,N_405);
nand U1202 (N_1202,In_1086,In_393);
nor U1203 (N_1203,In_1555,N_1183);
nand U1204 (N_1204,N_283,In_577);
nand U1205 (N_1205,In_714,N_258);
or U1206 (N_1206,N_1046,In_1803);
xor U1207 (N_1207,N_1051,N_623);
nand U1208 (N_1208,In_2052,N_287);
nor U1209 (N_1209,In_2430,N_559);
nor U1210 (N_1210,In_1666,In_835);
and U1211 (N_1211,In_1418,In_822);
and U1212 (N_1212,In_2172,In_1646);
nand U1213 (N_1213,N_1072,N_243);
xor U1214 (N_1214,N_556,In_1220);
nand U1215 (N_1215,In_2292,N_453);
nand U1216 (N_1216,N_1197,In_315);
or U1217 (N_1217,N_631,In_816);
nor U1218 (N_1218,In_1868,N_1098);
xor U1219 (N_1219,N_1016,N_1047);
nand U1220 (N_1220,N_867,In_1504);
nand U1221 (N_1221,In_2391,N_726);
and U1222 (N_1222,N_1157,In_1076);
and U1223 (N_1223,In_704,In_2083);
xnor U1224 (N_1224,N_609,In_1517);
nor U1225 (N_1225,In_2355,In_1568);
nor U1226 (N_1226,In_1620,N_1026);
xor U1227 (N_1227,In_621,N_180);
or U1228 (N_1228,N_1123,N_860);
xnor U1229 (N_1229,N_939,N_1160);
or U1230 (N_1230,N_908,In_523);
and U1231 (N_1231,N_1086,N_1064);
xnor U1232 (N_1232,In_32,In_1760);
nor U1233 (N_1233,In_464,In_1691);
nand U1234 (N_1234,In_1111,N_1002);
and U1235 (N_1235,N_700,N_1093);
nand U1236 (N_1236,N_903,N_1114);
nand U1237 (N_1237,In_946,N_927);
xor U1238 (N_1238,N_959,In_326);
xor U1239 (N_1239,In_411,N_768);
nor U1240 (N_1240,In_1564,N_24);
and U1241 (N_1241,N_896,N_600);
nor U1242 (N_1242,N_77,In_790);
nor U1243 (N_1243,N_264,In_954);
nand U1244 (N_1244,In_675,N_1023);
nand U1245 (N_1245,N_1126,N_1190);
and U1246 (N_1246,N_1144,In_1024);
xor U1247 (N_1247,N_289,In_291);
nand U1248 (N_1248,In_371,In_2413);
and U1249 (N_1249,In_1905,N_27);
nor U1250 (N_1250,In_261,N_489);
xor U1251 (N_1251,In_871,In_2267);
nor U1252 (N_1252,N_1166,In_867);
nor U1253 (N_1253,N_1048,In_1034);
nand U1254 (N_1254,In_1706,In_4);
nand U1255 (N_1255,In_2038,N_868);
nor U1256 (N_1256,N_1067,N_1041);
nand U1257 (N_1257,N_1020,In_370);
nor U1258 (N_1258,N_48,In_483);
nand U1259 (N_1259,N_479,N_1176);
xnor U1260 (N_1260,In_1281,In_2375);
xnor U1261 (N_1261,In_864,N_1085);
and U1262 (N_1262,In_2310,In_941);
or U1263 (N_1263,In_295,In_2402);
nand U1264 (N_1264,In_222,N_1088);
xnor U1265 (N_1265,In_369,N_412);
nand U1266 (N_1266,N_1124,In_53);
nor U1267 (N_1267,N_181,In_1265);
or U1268 (N_1268,N_753,In_1172);
nor U1269 (N_1269,In_1530,N_176);
or U1270 (N_1270,N_66,N_1029);
or U1271 (N_1271,N_764,In_2346);
nand U1272 (N_1272,N_123,N_629);
or U1273 (N_1273,In_1637,N_342);
nor U1274 (N_1274,In_1196,N_1054);
or U1275 (N_1275,In_1791,In_2367);
nor U1276 (N_1276,In_736,In_2139);
xor U1277 (N_1277,In_607,In_152);
nor U1278 (N_1278,In_2277,N_843);
or U1279 (N_1279,In_2461,N_75);
xnor U1280 (N_1280,N_164,N_296);
xnor U1281 (N_1281,In_1767,In_1533);
or U1282 (N_1282,In_1717,In_2398);
and U1283 (N_1283,N_890,In_1025);
nand U1284 (N_1284,In_1363,In_796);
and U1285 (N_1285,N_918,In_2005);
nand U1286 (N_1286,In_1598,N_255);
nor U1287 (N_1287,N_1036,N_610);
and U1288 (N_1288,N_732,N_683);
nand U1289 (N_1289,N_344,N_611);
and U1290 (N_1290,In_1682,N_567);
or U1291 (N_1291,N_480,In_549);
nor U1292 (N_1292,In_909,N_891);
nand U1293 (N_1293,N_979,N_1080);
or U1294 (N_1294,In_594,N_1019);
nor U1295 (N_1295,N_630,In_1047);
and U1296 (N_1296,N_323,N_1040);
xnor U1297 (N_1297,In_1772,In_752);
nand U1298 (N_1298,In_58,In_745);
nor U1299 (N_1299,N_759,N_1152);
and U1300 (N_1300,In_2339,N_909);
nand U1301 (N_1301,N_133,In_1999);
or U1302 (N_1302,N_852,In_2232);
nand U1303 (N_1303,In_1536,In_2302);
and U1304 (N_1304,N_131,N_838);
and U1305 (N_1305,In_1693,In_2325);
nand U1306 (N_1306,N_467,In_1337);
nand U1307 (N_1307,N_1027,N_1159);
xor U1308 (N_1308,N_931,N_1011);
nand U1309 (N_1309,N_1116,In_1437);
nand U1310 (N_1310,N_535,In_1401);
nand U1311 (N_1311,N_309,N_947);
or U1312 (N_1312,N_907,N_298);
and U1313 (N_1313,In_2491,N_870);
and U1314 (N_1314,In_1850,In_1741);
nand U1315 (N_1315,In_311,In_1326);
xor U1316 (N_1316,N_807,N_69);
and U1317 (N_1317,In_2146,In_691);
xnor U1318 (N_1318,N_594,In_969);
and U1319 (N_1319,N_910,In_1971);
xnor U1320 (N_1320,In_16,N_960);
or U1321 (N_1321,N_872,N_505);
and U1322 (N_1322,N_834,N_518);
nand U1323 (N_1323,N_447,In_247);
or U1324 (N_1324,N_1194,N_26);
and U1325 (N_1325,N_848,In_674);
nand U1326 (N_1326,In_1112,In_226);
xnor U1327 (N_1327,In_2248,In_270);
and U1328 (N_1328,In_919,N_433);
nand U1329 (N_1329,In_713,In_1189);
nor U1330 (N_1330,In_59,N_128);
or U1331 (N_1331,In_1960,In_1333);
nand U1332 (N_1332,In_1936,In_1316);
and U1333 (N_1333,In_787,In_1740);
nand U1334 (N_1334,N_796,In_2230);
or U1335 (N_1335,N_863,N_831);
and U1336 (N_1336,In_2340,In_1809);
xnor U1337 (N_1337,N_739,N_659);
or U1338 (N_1338,In_246,In_1433);
nand U1339 (N_1339,N_586,N_657);
xnor U1340 (N_1340,In_1148,In_27);
nand U1341 (N_1341,N_51,N_290);
and U1342 (N_1342,N_40,N_744);
xnor U1343 (N_1343,In_2448,N_712);
nand U1344 (N_1344,In_2366,N_386);
xor U1345 (N_1345,In_1144,N_1014);
xnor U1346 (N_1346,In_2498,N_563);
xnor U1347 (N_1347,N_970,N_921);
or U1348 (N_1348,N_894,In_29);
or U1349 (N_1349,N_730,In_1660);
or U1350 (N_1350,In_1965,In_2063);
nand U1351 (N_1351,In_583,N_1084);
or U1352 (N_1352,N_1112,N_590);
xor U1353 (N_1353,N_827,N_140);
or U1354 (N_1354,In_517,N_948);
or U1355 (N_1355,In_1151,In_2363);
and U1356 (N_1356,N_573,N_873);
and U1357 (N_1357,In_1941,N_1005);
and U1358 (N_1358,In_903,N_975);
nand U1359 (N_1359,N_968,In_868);
and U1360 (N_1360,N_185,N_1001);
xnor U1361 (N_1361,N_1115,N_1131);
nand U1362 (N_1362,In_618,N_388);
xnor U1363 (N_1363,N_901,N_713);
nand U1364 (N_1364,N_809,N_1148);
and U1365 (N_1365,N_107,N_1175);
or U1366 (N_1366,In_84,N_1099);
and U1367 (N_1367,N_236,N_897);
nor U1368 (N_1368,In_1427,N_1170);
xnor U1369 (N_1369,N_722,In_405);
nand U1370 (N_1370,In_1894,In_502);
and U1371 (N_1371,N_1171,N_926);
nand U1372 (N_1372,N_1151,In_1428);
nand U1373 (N_1373,In_294,In_384);
nor U1374 (N_1374,N_360,N_1089);
or U1375 (N_1375,In_1100,N_245);
nor U1376 (N_1376,In_1399,In_1562);
nor U1377 (N_1377,N_1119,N_714);
xor U1378 (N_1378,N_943,N_793);
and U1379 (N_1379,In_2209,N_1132);
xor U1380 (N_1380,In_1097,In_1429);
and U1381 (N_1381,In_1299,N_429);
nor U1382 (N_1382,N_864,In_1615);
or U1383 (N_1383,N_472,N_1169);
and U1384 (N_1384,In_937,In_1599);
xor U1385 (N_1385,In_1822,N_1033);
and U1386 (N_1386,N_1172,In_1787);
xnor U1387 (N_1387,N_1179,In_1329);
or U1388 (N_1388,N_452,N_551);
nor U1389 (N_1389,In_554,N_262);
nand U1390 (N_1390,N_1021,N_1096);
nand U1391 (N_1391,N_1195,N_933);
nand U1392 (N_1392,N_371,In_2224);
nand U1393 (N_1393,N_349,In_2256);
nand U1394 (N_1394,N_845,In_1155);
and U1395 (N_1395,In_2130,N_365);
or U1396 (N_1396,In_2147,N_1150);
and U1397 (N_1397,N_1017,N_1030);
or U1398 (N_1398,In_1550,N_354);
nor U1399 (N_1399,In_1934,N_416);
nor U1400 (N_1400,In_741,In_1154);
or U1401 (N_1401,N_1293,In_1443);
xnor U1402 (N_1402,N_1079,N_1184);
and U1403 (N_1403,In_1274,In_2258);
or U1404 (N_1404,N_1062,N_265);
nor U1405 (N_1405,N_913,In_873);
and U1406 (N_1406,In_475,N_1333);
nor U1407 (N_1407,N_1285,N_250);
or U1408 (N_1408,N_353,N_1104);
nand U1409 (N_1409,N_1140,In_1943);
nand U1410 (N_1410,In_2446,In_994);
nand U1411 (N_1411,N_787,N_1204);
xor U1412 (N_1412,N_674,N_1037);
xor U1413 (N_1413,N_881,N_1068);
xor U1414 (N_1414,In_2075,N_1289);
xnor U1415 (N_1415,N_427,In_2484);
nand U1416 (N_1416,In_1812,N_1317);
or U1417 (N_1417,N_1224,N_1209);
nor U1418 (N_1418,In_241,N_1181);
or U1419 (N_1419,In_781,N_1125);
or U1420 (N_1420,N_1288,N_1127);
and U1421 (N_1421,In_611,N_995);
nand U1422 (N_1422,N_1241,N_431);
xnor U1423 (N_1423,N_18,N_1376);
or U1424 (N_1424,In_542,N_1060);
nor U1425 (N_1425,In_2116,In_2450);
or U1426 (N_1426,In_1814,N_1003);
or U1427 (N_1427,N_889,N_1368);
nand U1428 (N_1428,In_377,N_1164);
nand U1429 (N_1429,N_564,In_1083);
xnor U1430 (N_1430,In_1466,N_572);
or U1431 (N_1431,In_1802,N_370);
or U1432 (N_1432,N_1167,N_800);
or U1433 (N_1433,In_1745,In_2137);
xor U1434 (N_1434,N_1297,N_1373);
nor U1435 (N_1435,N_501,In_2022);
nand U1436 (N_1436,N_1270,N_1185);
and U1437 (N_1437,N_116,N_645);
nand U1438 (N_1438,In_236,N_627);
or U1439 (N_1439,N_974,In_2161);
nand U1440 (N_1440,N_1387,N_937);
nor U1441 (N_1441,In_1044,In_2467);
or U1442 (N_1442,In_2092,N_665);
or U1443 (N_1443,N_977,In_1899);
and U1444 (N_1444,N_950,N_486);
nand U1445 (N_1445,N_1042,N_920);
and U1446 (N_1446,N_940,In_578);
or U1447 (N_1447,N_1313,N_813);
nor U1448 (N_1448,N_16,N_760);
nor U1449 (N_1449,N_854,N_1326);
nor U1450 (N_1450,N_998,N_229);
nand U1451 (N_1451,In_767,N_218);
xnor U1452 (N_1452,In_2306,In_922);
xnor U1453 (N_1453,In_1423,N_1363);
xor U1454 (N_1454,N_1292,N_437);
xnor U1455 (N_1455,N_22,In_336);
xnor U1456 (N_1456,N_856,N_1208);
nor U1457 (N_1457,In_646,In_2141);
nand U1458 (N_1458,N_1281,In_856);
and U1459 (N_1459,In_121,N_625);
or U1460 (N_1460,In_2049,N_914);
nor U1461 (N_1461,N_1073,N_1143);
nand U1462 (N_1462,N_626,N_1393);
xor U1463 (N_1463,In_188,In_423);
or U1464 (N_1464,N_526,N_1316);
nand U1465 (N_1465,In_357,N_1111);
and U1466 (N_1466,N_1121,N_592);
nand U1467 (N_1467,N_1233,N_1158);
xnor U1468 (N_1468,N_1396,In_1052);
nand U1469 (N_1469,N_364,N_1044);
or U1470 (N_1470,In_1779,In_133);
nor U1471 (N_1471,N_1028,In_1927);
xor U1472 (N_1472,N_1246,In_1798);
xnor U1473 (N_1473,N_956,In_2014);
nand U1474 (N_1474,N_980,In_2066);
nand U1475 (N_1475,N_1237,In_537);
and U1476 (N_1476,N_842,N_904);
and U1477 (N_1477,N_1381,N_136);
xor U1478 (N_1478,N_837,In_344);
and U1479 (N_1479,N_1065,N_1269);
nor U1480 (N_1480,In_2268,N_993);
nand U1481 (N_1481,N_1378,In_1089);
nor U1482 (N_1482,In_1612,In_1627);
xnor U1483 (N_1483,N_1307,N_1335);
or U1484 (N_1484,N_82,In_966);
xnor U1485 (N_1485,N_641,N_1232);
or U1486 (N_1486,In_898,In_131);
xor U1487 (N_1487,N_1198,In_1287);
nand U1488 (N_1488,In_286,In_23);
xor U1489 (N_1489,In_1493,N_60);
xnor U1490 (N_1490,N_836,In_1408);
or U1491 (N_1491,In_481,In_1117);
and U1492 (N_1492,In_877,N_990);
and U1493 (N_1493,N_1009,In_1243);
nand U1494 (N_1494,In_2404,In_1686);
xnor U1495 (N_1495,N_788,In_332);
nor U1496 (N_1496,In_1315,In_579);
or U1497 (N_1497,In_716,N_1302);
or U1498 (N_1498,In_2202,In_1712);
and U1499 (N_1499,N_1133,In_2197);
xor U1500 (N_1500,N_971,In_2441);
and U1501 (N_1501,N_1355,N_661);
and U1502 (N_1502,N_855,In_888);
or U1503 (N_1503,N_1103,N_1216);
or U1504 (N_1504,In_1473,In_2174);
nor U1505 (N_1505,In_768,In_1898);
nand U1506 (N_1506,In_1883,In_366);
and U1507 (N_1507,N_110,N_1049);
or U1508 (N_1508,N_621,N_1082);
nand U1509 (N_1509,N_1228,In_1227);
and U1510 (N_1510,N_829,In_1735);
and U1511 (N_1511,N_945,In_2465);
or U1512 (N_1512,In_269,In_1697);
nand U1513 (N_1513,N_1364,N_1279);
xor U1514 (N_1514,N_1092,N_1202);
or U1515 (N_1515,N_246,In_2373);
xnor U1516 (N_1516,In_112,N_1076);
xnor U1517 (N_1517,N_219,N_1155);
or U1518 (N_1518,N_1253,N_1238);
nor U1519 (N_1519,In_1846,N_1214);
nor U1520 (N_1520,N_251,N_1015);
xnor U1521 (N_1521,N_485,N_542);
nand U1522 (N_1522,N_1383,N_1258);
nor U1523 (N_1523,In_1733,In_1482);
nand U1524 (N_1524,N_1018,N_1296);
xor U1525 (N_1525,In_1007,N_1318);
nor U1526 (N_1526,N_1039,N_1180);
nor U1527 (N_1527,N_183,N_543);
or U1528 (N_1528,In_1716,In_1916);
or U1529 (N_1529,N_658,In_1472);
nand U1530 (N_1530,In_99,N_175);
nor U1531 (N_1531,In_2369,N_957);
nand U1532 (N_1532,N_1245,N_952);
nand U1533 (N_1533,N_805,N_1182);
or U1534 (N_1534,N_25,In_102);
nor U1535 (N_1535,N_1366,N_1388);
or U1536 (N_1536,N_310,In_480);
xor U1537 (N_1537,N_646,N_162);
nor U1538 (N_1538,N_1141,N_585);
nand U1539 (N_1539,N_981,N_1163);
xor U1540 (N_1540,In_1563,N_797);
nand U1541 (N_1541,N_87,N_1319);
xor U1542 (N_1542,In_1355,N_1379);
nor U1543 (N_1543,In_2255,N_1192);
xor U1544 (N_1544,N_41,N_558);
nor U1545 (N_1545,N_1249,N_1053);
nand U1546 (N_1546,In_935,In_1347);
nand U1547 (N_1547,N_1095,In_60);
nor U1548 (N_1548,In_244,N_1399);
or U1549 (N_1549,In_2187,In_820);
and U1550 (N_1550,N_463,N_402);
and U1551 (N_1551,In_1665,N_1322);
nor U1552 (N_1552,In_63,In_1252);
xor U1553 (N_1553,N_1341,In_1671);
or U1554 (N_1554,N_541,N_705);
and U1555 (N_1555,N_620,In_1186);
xor U1556 (N_1556,N_203,N_361);
nand U1557 (N_1557,In_1393,N_1235);
or U1558 (N_1558,N_769,N_1294);
or U1559 (N_1559,N_190,In_1440);
xnor U1560 (N_1560,In_190,N_340);
or U1561 (N_1561,In_504,N_1007);
nand U1562 (N_1562,In_1863,N_443);
xor U1563 (N_1563,In_2371,In_1368);
or U1564 (N_1564,N_1142,In_1680);
or U1565 (N_1565,N_816,N_260);
or U1566 (N_1566,N_238,N_1043);
nor U1567 (N_1567,N_389,N_1251);
or U1568 (N_1568,N_875,N_417);
nor U1569 (N_1569,N_835,N_1255);
xnor U1570 (N_1570,In_179,In_889);
nand U1571 (N_1571,N_483,In_1087);
and U1572 (N_1572,In_422,N_1200);
xor U1573 (N_1573,In_571,In_878);
or U1574 (N_1574,In_489,N_1102);
or U1575 (N_1575,In_866,In_1001);
and U1576 (N_1576,N_1225,N_1331);
xor U1577 (N_1577,N_517,In_1053);
nor U1578 (N_1578,In_404,In_2095);
or U1579 (N_1579,N_247,N_119);
nand U1580 (N_1580,In_789,N_604);
nand U1581 (N_1581,N_1050,In_2003);
nand U1582 (N_1582,In_557,N_1134);
xnor U1583 (N_1583,N_1203,N_1059);
or U1584 (N_1584,N_731,In_8);
and U1585 (N_1585,N_1045,In_617);
and U1586 (N_1586,In_2298,In_1272);
nor U1587 (N_1587,In_2383,N_372);
and U1588 (N_1588,In_998,In_2285);
nor U1589 (N_1589,N_961,N_1300);
or U1590 (N_1590,N_1078,N_415);
nand U1591 (N_1591,In_220,In_308);
xnor U1592 (N_1592,N_1365,In_149);
nand U1593 (N_1593,N_719,N_1052);
and U1594 (N_1594,N_1263,N_810);
nor U1595 (N_1595,N_1117,N_1022);
nor U1596 (N_1596,In_1344,In_151);
nor U1597 (N_1597,N_1315,N_1122);
nor U1598 (N_1598,In_1594,In_746);
nand U1599 (N_1599,In_771,N_853);
nor U1600 (N_1600,N_1513,N_1257);
nand U1601 (N_1601,N_1519,N_1162);
or U1602 (N_1602,N_660,N_1361);
or U1603 (N_1603,N_1284,N_253);
nand U1604 (N_1604,N_1451,N_84);
and U1605 (N_1605,N_915,N_1427);
or U1606 (N_1606,In_1439,N_1286);
xnor U1607 (N_1607,In_442,N_1342);
and U1608 (N_1608,In_869,In_1589);
nor U1609 (N_1609,N_1345,In_374);
or U1610 (N_1610,In_285,In_12);
or U1611 (N_1611,N_1529,In_2152);
or U1612 (N_1612,In_2291,N_1524);
nand U1613 (N_1613,In_1527,In_1951);
nand U1614 (N_1614,In_1582,In_1681);
and U1615 (N_1615,In_952,In_525);
nand U1616 (N_1616,In_1825,N_1530);
nand U1617 (N_1617,N_1201,N_451);
and U1618 (N_1618,N_1538,In_1542);
nor U1619 (N_1619,N_1504,N_1324);
or U1620 (N_1620,N_1437,In_1115);
or U1621 (N_1621,In_2053,N_1499);
or U1622 (N_1622,In_788,N_1586);
and U1623 (N_1623,In_2284,N_1455);
nor U1624 (N_1624,N_1502,In_677);
nand U1625 (N_1625,In_602,N_1024);
nand U1626 (N_1626,N_878,N_1572);
xnor U1627 (N_1627,N_1304,N_1438);
xor U1628 (N_1628,N_39,In_132);
xor U1629 (N_1629,N_694,N_1496);
and U1630 (N_1630,In_982,N_1215);
xor U1631 (N_1631,N_1434,N_1392);
nor U1632 (N_1632,In_2184,N_1398);
and U1633 (N_1633,N_1421,N_1574);
or U1634 (N_1634,N_735,N_1485);
nand U1635 (N_1635,N_1484,In_1406);
nor U1636 (N_1636,N_647,N_746);
nand U1637 (N_1637,In_2345,In_1755);
nor U1638 (N_1638,N_1474,N_240);
xor U1639 (N_1639,N_1526,N_1479);
nor U1640 (N_1640,N_752,N_1311);
and U1641 (N_1641,In_2379,N_343);
nand U1642 (N_1642,N_1219,N_17);
nor U1643 (N_1643,N_1509,N_1303);
xor U1644 (N_1644,N_900,In_1270);
xor U1645 (N_1645,N_52,N_680);
nand U1646 (N_1646,In_2122,N_275);
xor U1647 (N_1647,In_104,In_2170);
nor U1648 (N_1648,N_36,In_626);
and U1649 (N_1649,In_628,N_1008);
nor U1650 (N_1650,In_1974,N_458);
xnor U1651 (N_1651,In_2055,In_2427);
and U1652 (N_1652,N_1448,In_544);
xnor U1653 (N_1653,N_1578,N_449);
xnor U1654 (N_1654,N_1356,In_191);
or U1655 (N_1655,N_407,In_1799);
xnor U1656 (N_1656,N_1561,N_1535);
and U1657 (N_1657,In_443,In_1685);
or U1658 (N_1658,N_1384,N_3);
nor U1659 (N_1659,N_1153,N_102);
nor U1660 (N_1660,N_1120,N_1012);
xor U1661 (N_1661,In_780,N_1268);
nor U1662 (N_1662,N_1357,N_1222);
xor U1663 (N_1663,In_1914,N_1013);
nor U1664 (N_1664,N_419,N_1436);
nor U1665 (N_1665,N_1557,N_978);
and U1666 (N_1666,N_1488,In_2206);
nand U1667 (N_1667,N_1400,N_50);
and U1668 (N_1668,N_172,N_1391);
nand U1669 (N_1669,N_514,N_1465);
or U1670 (N_1670,N_1066,N_1478);
nand U1671 (N_1671,In_772,N_801);
nand U1672 (N_1672,N_1339,N_917);
xor U1673 (N_1673,N_1410,N_1518);
nor U1674 (N_1674,N_528,N_142);
xnor U1675 (N_1675,N_1505,N_474);
nand U1676 (N_1676,N_1495,N_1147);
xor U1677 (N_1677,In_2094,N_1308);
or U1678 (N_1678,N_643,N_1463);
nand U1679 (N_1679,In_91,N_1594);
or U1680 (N_1680,In_2090,In_124);
nand U1681 (N_1681,N_1309,N_902);
nor U1682 (N_1682,N_1058,N_1422);
and U1683 (N_1683,N_1113,In_2217);
and U1684 (N_1684,N_1406,In_1004);
nand U1685 (N_1685,N_1470,In_465);
nand U1686 (N_1686,N_1034,N_1108);
nor U1687 (N_1687,In_1762,N_953);
or U1688 (N_1688,N_1441,In_2382);
and U1689 (N_1689,In_1704,N_1403);
or U1690 (N_1690,N_498,N_1234);
nand U1691 (N_1691,N_880,In_1460);
xor U1692 (N_1692,In_427,In_1933);
or U1693 (N_1693,N_1385,N_527);
nand U1694 (N_1694,In_1430,N_1446);
nor U1695 (N_1695,In_1881,N_23);
nor U1696 (N_1696,In_700,In_1079);
or U1697 (N_1697,In_1655,In_360);
nor U1698 (N_1698,N_1454,N_1358);
and U1699 (N_1699,N_152,N_1559);
and U1700 (N_1700,In_1980,In_175);
or U1701 (N_1701,N_1178,N_888);
and U1702 (N_1702,In_2058,N_1588);
or U1703 (N_1703,N_545,In_1724);
xor U1704 (N_1704,N_126,N_1522);
nand U1705 (N_1705,In_1945,N_1231);
xnor U1706 (N_1706,N_1282,In_1387);
nand U1707 (N_1707,N_1374,N_1032);
nor U1708 (N_1708,N_1212,N_1503);
nor U1709 (N_1709,N_1584,N_1106);
nand U1710 (N_1710,In_912,In_490);
or U1711 (N_1711,N_1469,N_929);
or U1712 (N_1712,In_786,In_1955);
nand U1713 (N_1713,N_876,N_1031);
nor U1714 (N_1714,In_2254,N_1248);
xor U1715 (N_1715,N_638,N_738);
nand U1716 (N_1716,N_1382,N_1301);
or U1717 (N_1717,N_1390,N_1273);
or U1718 (N_1718,N_1407,N_1587);
xnor U1719 (N_1719,In_320,In_1556);
nand U1720 (N_1720,N_1532,N_1264);
nand U1721 (N_1721,In_1470,In_615);
xnor U1722 (N_1722,N_1456,N_1329);
and U1723 (N_1723,N_1408,N_883);
and U1724 (N_1724,N_1320,N_1107);
and U1725 (N_1725,N_1490,In_1859);
or U1726 (N_1726,N_239,N_1372);
xnor U1727 (N_1727,N_1186,N_817);
xnor U1728 (N_1728,N_785,N_367);
nor U1729 (N_1729,In_233,N_644);
or U1730 (N_1730,N_954,N_209);
xnor U1731 (N_1731,N_1542,In_397);
or U1732 (N_1732,N_1555,N_1254);
nand U1733 (N_1733,In_2378,In_1188);
or U1734 (N_1734,In_284,N_1261);
and U1735 (N_1735,In_1765,N_1305);
or U1736 (N_1736,N_1128,In_1923);
and U1737 (N_1737,N_893,N_1556);
or U1738 (N_1738,N_985,In_1369);
and U1739 (N_1739,In_199,N_1492);
and U1740 (N_1740,N_1283,N_1189);
or U1741 (N_1741,In_81,N_308);
and U1742 (N_1742,N_743,N_1590);
xnor U1743 (N_1743,In_791,N_271);
and U1744 (N_1744,N_1343,In_1981);
xnor U1745 (N_1745,N_1508,N_1428);
and U1746 (N_1746,In_2344,N_1210);
nor U1747 (N_1747,N_1517,N_1598);
or U1748 (N_1748,In_665,N_1161);
xnor U1749 (N_1749,N_1006,N_1321);
and U1750 (N_1750,N_1154,N_1135);
xnor U1751 (N_1751,N_830,In_1163);
and U1752 (N_1752,N_1325,N_756);
or U1753 (N_1753,N_1347,N_818);
and U1754 (N_1754,N_1330,N_608);
xor U1755 (N_1755,N_1063,In_989);
nand U1756 (N_1756,N_1511,N_570);
nand U1757 (N_1757,N_1352,In_1157);
or U1758 (N_1758,In_854,N_671);
xnor U1759 (N_1759,N_1536,In_1207);
xor U1760 (N_1760,N_1431,N_1118);
and U1761 (N_1761,N_1416,In_409);
or U1762 (N_1762,In_1045,In_1356);
xor U1763 (N_1763,In_1449,N_1291);
xor U1764 (N_1764,N_1554,N_1548);
nand U1765 (N_1765,N_1443,In_1558);
nor U1766 (N_1766,In_1897,In_992);
xor U1767 (N_1767,N_1340,N_1493);
or U1768 (N_1768,In_1781,N_1250);
xor U1769 (N_1769,N_1071,In_271);
and U1770 (N_1770,In_1848,N_1459);
nand U1771 (N_1771,N_1570,N_1259);
nand U1772 (N_1772,N_1444,In_568);
and U1773 (N_1773,In_887,N_57);
nand U1774 (N_1774,N_919,In_850);
xor U1775 (N_1775,N_1440,In_1334);
or U1776 (N_1776,N_1544,N_972);
xor U1777 (N_1777,N_1458,In_307);
and U1778 (N_1778,In_1396,N_1074);
xnor U1779 (N_1779,N_1165,In_1307);
nand U1780 (N_1780,In_51,N_1461);
or U1781 (N_1781,In_1310,In_540);
nand U1782 (N_1782,In_1043,In_1644);
nor U1783 (N_1783,N_733,N_244);
or U1784 (N_1784,In_88,N_932);
nand U1785 (N_1785,N_1247,In_1258);
nand U1786 (N_1786,N_859,N_1240);
xnor U1787 (N_1787,N_1295,In_1203);
xnor U1788 (N_1788,In_2207,N_1447);
nor U1789 (N_1789,In_305,N_1395);
nand U1790 (N_1790,N_409,In_2337);
xor U1791 (N_1791,N_1205,N_663);
nand U1792 (N_1792,N_1109,N_1299);
nand U1793 (N_1793,N_1573,N_1010);
nor U1794 (N_1794,N_1547,N_987);
xor U1795 (N_1795,N_1221,N_1487);
nor U1796 (N_1796,In_368,In_555);
and U1797 (N_1797,In_2395,N_1267);
nor U1798 (N_1798,In_2102,N_1596);
xnor U1799 (N_1799,In_476,N_851);
and U1800 (N_1800,N_1777,N_302);
nand U1801 (N_1801,N_1707,In_1966);
and U1802 (N_1802,N_1213,N_1697);
and U1803 (N_1803,N_1429,In_1475);
nand U1804 (N_1804,N_582,N_1742);
xor U1805 (N_1805,In_2074,N_470);
nor U1806 (N_1806,N_1749,In_240);
nand U1807 (N_1807,N_1498,N_1420);
nand U1808 (N_1808,N_1660,N_1786);
xnor U1809 (N_1809,N_1661,In_1677);
and U1810 (N_1810,N_1276,N_1218);
xnor U1811 (N_1811,N_1386,In_460);
xnor U1812 (N_1812,N_1227,N_319);
nand U1813 (N_1813,In_302,N_1056);
nand U1814 (N_1814,N_1701,N_1759);
or U1815 (N_1815,N_1553,N_1655);
or U1816 (N_1816,N_1683,N_1433);
nor U1817 (N_1817,N_1671,N_1632);
and U1818 (N_1818,N_1754,In_1416);
nor U1819 (N_1819,N_879,N_850);
nor U1820 (N_1820,N_1610,In_2125);
xor U1821 (N_1821,N_1424,N_1613);
nand U1822 (N_1822,N_1537,N_1314);
nand U1823 (N_1823,N_1298,N_520);
or U1824 (N_1824,N_1362,In_1161);
nand U1825 (N_1825,N_1637,N_1647);
nand U1826 (N_1826,In_2205,N_1277);
xor U1827 (N_1827,N_1776,N_1617);
nand U1828 (N_1828,N_194,In_706);
and U1829 (N_1829,In_893,N_1793);
nand U1830 (N_1830,N_1649,In_1105);
nor U1831 (N_1831,N_1512,N_1719);
nor U1832 (N_1832,In_1351,N_1272);
xnor U1833 (N_1833,N_1353,In_1813);
or U1834 (N_1834,In_972,N_1145);
xor U1835 (N_1835,In_1593,N_1728);
nand U1836 (N_1836,N_1401,N_986);
xnor U1837 (N_1837,N_989,N_362);
nor U1838 (N_1838,N_781,N_462);
xnor U1839 (N_1839,N_1580,N_1405);
or U1840 (N_1840,N_1507,N_1612);
or U1841 (N_1841,N_1732,N_1706);
xor U1842 (N_1842,N_1752,N_1738);
and U1843 (N_1843,N_552,N_1566);
nor U1844 (N_1844,N_347,In_2077);
or U1845 (N_1845,N_1745,N_678);
xor U1846 (N_1846,N_1717,N_1643);
xor U1847 (N_1847,In_2304,N_1653);
and U1848 (N_1848,N_1534,N_1327);
nor U1849 (N_1849,In_1673,N_824);
nand U1850 (N_1850,N_1782,N_1389);
nand U1851 (N_1851,N_1780,N_1644);
nor U1852 (N_1852,In_2260,In_574);
nand U1853 (N_1853,N_1336,N_1725);
nand U1854 (N_1854,N_1727,N_1097);
and U1855 (N_1855,In_1795,N_717);
nand U1856 (N_1856,N_1792,N_1271);
nor U1857 (N_1857,N_1500,N_345);
xor U1858 (N_1858,N_1789,N_584);
nand U1859 (N_1859,N_964,N_1367);
and U1860 (N_1860,In_1414,N_1607);
nor U1861 (N_1861,N_73,N_1730);
xnor U1862 (N_1862,In_180,N_839);
and U1863 (N_1863,N_1623,N_696);
xor U1864 (N_1864,N_1100,N_1191);
nand U1865 (N_1865,N_1476,N_1412);
xnor U1866 (N_1866,In_598,N_669);
nand U1867 (N_1867,N_1081,N_1672);
nor U1868 (N_1868,In_2322,In_2422);
nor U1869 (N_1869,N_1256,N_1592);
nand U1870 (N_1870,N_1418,N_1312);
xnor U1871 (N_1871,In_988,N_662);
and U1872 (N_1872,N_1691,N_1760);
and U1873 (N_1873,In_196,N_1615);
or U1874 (N_1874,N_1252,N_1230);
xnor U1875 (N_1875,N_1638,N_576);
nand U1876 (N_1876,N_1266,N_1582);
nand U1877 (N_1877,N_10,N_1664);
nand U1878 (N_1878,N_1287,N_1666);
nor U1879 (N_1879,In_1675,N_1724);
xnor U1880 (N_1880,N_1662,N_1236);
or U1881 (N_1881,In_42,N_1371);
nor U1882 (N_1882,N_1101,In_2495);
and U1883 (N_1883,N_1415,In_1132);
nand U1884 (N_1884,N_946,N_1543);
and U1885 (N_1885,N_1673,N_1430);
nand U1886 (N_1886,N_1229,N_1494);
nand U1887 (N_1887,In_439,N_221);
nor U1888 (N_1888,N_1467,N_1757);
nor U1889 (N_1889,N_261,N_1568);
or U1890 (N_1890,N_1619,In_1626);
xnor U1891 (N_1891,N_1571,N_607);
xnor U1892 (N_1892,N_1435,N_1796);
nor U1893 (N_1893,In_1815,In_1373);
and U1894 (N_1894,In_2330,N_1713);
or U1895 (N_1895,N_741,N_1631);
or U1896 (N_1896,N_1539,N_1771);
xor U1897 (N_1897,N_1658,In_1638);
nand U1898 (N_1898,In_1549,N_1714);
nor U1899 (N_1899,N_1639,N_965);
or U1900 (N_1900,N_1654,N_1591);
xnor U1901 (N_1901,N_1627,N_1462);
and U1902 (N_1902,In_770,N_1274);
or U1903 (N_1903,N_1693,N_1149);
and U1904 (N_1904,N_1648,N_1703);
nor U1905 (N_1905,N_1773,In_2021);
and U1906 (N_1906,N_1334,In_1068);
or U1907 (N_1907,N_1700,N_766);
or U1908 (N_1908,N_1774,In_1958);
nand U1909 (N_1909,N_1663,N_849);
nand U1910 (N_1910,N_1531,N_1000);
or U1911 (N_1911,In_813,N_1567);
nand U1912 (N_1912,In_805,N_690);
and U1913 (N_1913,N_1576,N_1477);
nor U1914 (N_1914,N_1442,N_280);
and U1915 (N_1915,In_2483,N_1729);
or U1916 (N_1916,In_1696,N_1709);
and U1917 (N_1917,N_1748,N_1091);
or U1918 (N_1918,N_1645,N_1758);
and U1919 (N_1919,N_1533,N_598);
nand U1920 (N_1920,N_955,N_1747);
nand U1921 (N_1921,In_2437,N_1377);
nor U1922 (N_1922,N_1694,In_1168);
xnor U1923 (N_1923,N_1207,N_1370);
nor U1924 (N_1924,N_1763,N_1715);
nand U1925 (N_1925,N_1278,N_771);
and U1926 (N_1926,N_418,N_597);
nor U1927 (N_1927,N_1682,N_487);
and U1928 (N_1928,N_1737,In_1050);
or U1929 (N_1929,In_550,N_624);
nor U1930 (N_1930,N_1621,N_1482);
nand U1931 (N_1931,N_212,N_1736);
and U1932 (N_1932,N_383,N_1608);
or U1933 (N_1933,N_1640,N_847);
nor U1934 (N_1934,N_1332,N_1794);
or U1935 (N_1935,N_468,In_1667);
and U1936 (N_1936,N_37,N_938);
or U1937 (N_1937,N_865,N_1740);
nor U1938 (N_1938,N_906,N_1702);
nor U1939 (N_1939,In_1928,N_1489);
nor U1940 (N_1940,N_1635,In_776);
and U1941 (N_1941,N_862,In_456);
nor U1942 (N_1942,N_1223,N_1690);
nand U1943 (N_1943,N_1411,N_1349);
and U1944 (N_1944,N_1328,N_1211);
and U1945 (N_1945,In_217,N_1226);
or U1946 (N_1946,In_325,In_2242);
or U1947 (N_1947,N_1545,N_1723);
nor U1948 (N_1948,In_2326,N_1244);
or U1949 (N_1949,N_686,N_1597);
xor U1950 (N_1950,N_1798,N_1310);
and U1951 (N_1951,N_109,N_1668);
or U1952 (N_1952,In_1519,N_1687);
or U1953 (N_1953,N_1761,N_1744);
xnor U1954 (N_1954,N_840,In_1211);
and U1955 (N_1955,N_1243,N_651);
nand U1956 (N_1956,N_1090,N_1670);
nor U1957 (N_1957,N_1025,N_1600);
or U1958 (N_1958,N_1359,In_1143);
and U1959 (N_1959,N_928,N_1473);
nand U1960 (N_1960,N_748,N_1472);
nor U1961 (N_1961,N_1739,In_849);
nor U1962 (N_1962,N_605,In_408);
or U1963 (N_1963,In_98,N_1785);
xnor U1964 (N_1964,N_352,N_1712);
and U1965 (N_1965,N_1603,In_274);
nand U1966 (N_1966,N_1188,N_557);
and U1967 (N_1967,N_1480,In_629);
nand U1968 (N_1968,In_1292,N_1523);
xnor U1969 (N_1969,N_1346,In_2475);
or U1970 (N_1970,In_278,N_249);
or U1971 (N_1971,N_1550,N_1563);
nor U1972 (N_1972,N_877,N_1775);
nand U1973 (N_1973,N_1795,N_1756);
and U1974 (N_1974,N_1720,N_999);
or U1975 (N_1975,N_1070,N_1577);
and U1976 (N_1976,In_1507,N_991);
nor U1977 (N_1977,In_1695,N_1575);
nand U1978 (N_1978,N_615,N_459);
nor U1979 (N_1979,N_1769,N_685);
or U1980 (N_1980,N_1684,N_504);
nand U1981 (N_1981,N_763,N_844);
or U1982 (N_1982,N_1419,N_53);
nand U1983 (N_1983,N_1779,N_1772);
or U1984 (N_1984,N_1280,N_1710);
xor U1985 (N_1985,N_1698,N_1540);
xnor U1986 (N_1986,N_1616,In_1260);
and U1987 (N_1987,N_1650,In_2438);
and U1988 (N_1988,N_899,In_479);
nor U1989 (N_1989,N_1784,N_988);
xor U1990 (N_1990,In_290,N_1510);
xor U1991 (N_1991,N_1369,In_1078);
nand U1992 (N_1992,N_924,N_1035);
xor U1993 (N_1993,N_1491,N_1681);
nor U1994 (N_1994,In_858,N_1716);
and U1995 (N_1995,N_1569,N_1551);
nand U1996 (N_1996,N_1514,In_548);
or U1997 (N_1997,N_1692,N_1602);
xor U1998 (N_1998,N_1679,N_1338);
and U1999 (N_1999,N_1156,N_1726);
nand U2000 (N_2000,N_871,N_1583);
nand U2001 (N_2001,N_1380,N_1828);
and U2002 (N_2002,N_1903,N_1940);
nand U2003 (N_2003,N_1686,N_1999);
and U2004 (N_2004,N_1452,N_1680);
or U2005 (N_2005,In_111,N_1860);
nor U2006 (N_2006,N_857,N_1483);
or U2007 (N_2007,N_1075,N_1193);
nor U2008 (N_2008,N_1604,N_1846);
nand U2009 (N_2009,N_328,N_1956);
nor U2010 (N_2010,N_1705,N_1871);
or U2011 (N_2011,N_1558,In_2396);
or U2012 (N_2012,N_1667,N_1004);
xor U2013 (N_2013,N_1527,N_270);
xnor U2014 (N_2014,N_1933,N_1625);
xor U2015 (N_2015,In_1275,N_1875);
nor U2016 (N_2016,N_1677,N_1624);
xnor U2017 (N_2017,N_1965,N_1764);
and U2018 (N_2018,N_1768,N_1886);
xnor U2019 (N_2019,N_1976,N_1375);
xnor U2020 (N_2020,N_1822,N_1946);
nor U2021 (N_2021,N_1925,N_1967);
nor U2022 (N_2022,N_403,N_1909);
and U2023 (N_2023,In_2007,N_1960);
or U2024 (N_2024,N_1136,In_1468);
xnor U2025 (N_2025,N_146,N_1939);
and U2026 (N_2026,In_2280,N_1077);
nand U2027 (N_2027,N_1481,N_1404);
xor U2028 (N_2028,N_1674,N_450);
nand U2029 (N_2029,N_1174,N_1815);
xnor U2030 (N_2030,N_1541,N_1926);
xor U2031 (N_2031,N_1242,N_687);
and U2032 (N_2032,N_1920,N_1652);
nand U2033 (N_2033,N_1515,N_1595);
or U2034 (N_2034,N_1818,N_1528);
nor U2035 (N_2035,N_1453,N_1426);
nor U2036 (N_2036,N_1872,N_1741);
and U2037 (N_2037,N_1892,N_1975);
nor U2038 (N_2038,N_634,N_1913);
nand U2039 (N_2039,N_1110,In_808);
xnor U2040 (N_2040,N_1853,N_1980);
or U2041 (N_2041,N_1402,N_1599);
nand U2042 (N_2042,N_1893,N_1589);
nor U2043 (N_2043,In_64,In_634);
nor U2044 (N_2044,N_803,N_1560);
xor U2045 (N_2045,N_885,In_1182);
or U2046 (N_2046,N_1460,N_1953);
nand U2047 (N_2047,N_1620,N_1685);
xor U2048 (N_2048,N_1998,N_1626);
nand U2049 (N_2049,N_1839,In_85);
and U2050 (N_2050,N_1622,N_1506);
or U2051 (N_2051,N_1445,N_1425);
nor U2052 (N_2052,N_421,N_1989);
nor U2053 (N_2053,N_1858,N_1177);
and U2054 (N_2054,N_1781,N_1832);
xnor U2055 (N_2055,N_1290,N_1838);
and U2056 (N_2056,N_223,N_1579);
xnor U2057 (N_2057,N_1833,N_1981);
or U2058 (N_2058,N_1819,N_1486);
nand U2059 (N_2059,N_1963,N_1521);
xor U2060 (N_2060,N_707,In_1108);
and U2061 (N_2061,N_1830,N_1843);
nand U2062 (N_2062,N_640,N_1921);
nand U2063 (N_2063,N_1932,In_499);
or U2064 (N_2064,N_1413,N_811);
and U2065 (N_2065,N_1951,N_1651);
and U2066 (N_2066,N_1605,N_1897);
and U2067 (N_2067,N_1911,N_613);
nor U2068 (N_2068,N_1905,In_94);
nand U2069 (N_2069,N_1766,N_1961);
or U2070 (N_2070,N_1944,N_1783);
xnor U2071 (N_2071,N_1414,N_1936);
and U2072 (N_2072,N_702,N_307);
xor U2073 (N_2073,N_1857,N_1907);
or U2074 (N_2074,N_1889,N_1825);
and U2075 (N_2075,N_1601,N_1912);
or U2076 (N_2076,N_1906,N_1806);
nor U2077 (N_2077,N_1770,N_1952);
nand U2078 (N_2078,N_1850,N_1394);
nor U2079 (N_2079,In_341,N_1988);
and U2080 (N_2080,N_1146,N_1884);
xnor U2081 (N_2081,N_1870,N_773);
or U2082 (N_2082,N_695,N_1895);
or U2083 (N_2083,N_1704,N_1869);
nand U2084 (N_2084,N_1417,In_2314);
xor U2085 (N_2085,In_1095,In_1297);
or U2086 (N_2086,N_1862,N_1265);
xnor U2087 (N_2087,N_1471,N_1721);
nand U2088 (N_2088,N_1904,N_537);
nand U2089 (N_2089,N_1957,In_2316);
or U2090 (N_2090,N_1820,N_1938);
nand U2091 (N_2091,N_1929,N_1409);
xnor U2092 (N_2092,N_1955,N_1807);
or U2093 (N_2093,N_1829,N_1811);
or U2094 (N_2094,N_1220,N_1919);
nand U2095 (N_2095,N_1835,N_1924);
nand U2096 (N_2096,N_967,N_1676);
and U2097 (N_2097,N_1734,N_1791);
and U2098 (N_2098,N_1803,N_1038);
xor U2099 (N_2099,N_1805,N_1630);
or U2100 (N_2100,In_1378,N_1778);
nand U2101 (N_2101,N_1982,N_1606);
nor U2102 (N_2102,N_1562,In_314);
xor U2103 (N_2103,N_1996,N_1995);
or U2104 (N_2104,N_1788,N_1217);
or U2105 (N_2105,N_969,N_1851);
and U2106 (N_2106,In_1388,N_1611);
nand U2107 (N_2107,N_1129,N_1997);
xor U2108 (N_2108,N_1934,N_387);
xnor U2109 (N_2109,In_1228,N_1877);
xnor U2110 (N_2110,N_1199,N_1549);
nor U2111 (N_2111,N_1977,N_1450);
nor U2112 (N_2112,N_1765,N_1564);
nor U2113 (N_2113,N_1468,N_1935);
and U2114 (N_2114,N_1863,N_1735);
nor U2115 (N_2115,N_1239,N_1708);
xor U2116 (N_2116,N_1618,N_1882);
and U2117 (N_2117,N_1915,N_1950);
and U2118 (N_2118,N_1733,N_1432);
xnor U2119 (N_2119,N_482,N_826);
xor U2120 (N_2120,N_1970,N_1196);
xnor U2121 (N_2121,N_1449,N_1609);
xnor U2122 (N_2122,N_1057,N_1350);
or U2123 (N_2123,N_1898,N_1646);
xnor U2124 (N_2124,In_309,N_488);
nand U2125 (N_2125,N_814,N_1525);
and U2126 (N_2126,N_1834,N_1464);
and U2127 (N_2127,N_1873,In_1259);
or U2128 (N_2128,N_1847,N_1337);
and U2129 (N_2129,N_1900,In_2);
nand U2130 (N_2130,N_725,N_1816);
or U2131 (N_2131,N_1069,N_1750);
xnor U2132 (N_2132,N_1348,N_1917);
nor U2133 (N_2133,In_349,N_1767);
xor U2134 (N_2134,N_1812,N_1187);
xor U2135 (N_2135,N_1351,In_1029);
nand U2136 (N_2136,N_1642,N_9);
and U2137 (N_2137,N_1993,N_925);
xnor U2138 (N_2138,N_1840,N_1991);
or U2139 (N_2139,In_1817,N_1878);
and U2140 (N_2140,N_1922,N_1813);
xor U2141 (N_2141,N_951,N_1804);
or U2142 (N_2142,N_266,N_996);
or U2143 (N_2143,N_1699,N_1948);
nor U2144 (N_2144,N_1821,N_1746);
xor U2145 (N_2145,N_1881,N_1641);
nor U2146 (N_2146,N_1094,N_1801);
xnor U2147 (N_2147,N_1718,In_685);
nand U2148 (N_2148,N_1883,N_1137);
nor U2149 (N_2149,N_1958,N_1665);
xnor U2150 (N_2150,N_1856,N_1753);
or U2151 (N_2151,N_1947,N_869);
nor U2152 (N_2152,N_1962,N_994);
xnor U2153 (N_2153,In_6,N_1636);
or U2154 (N_2154,N_1930,N_1397);
nand U2155 (N_2155,In_1892,N_1979);
nand U2156 (N_2156,N_1987,In_600);
and U2157 (N_2157,N_1823,N_1323);
nor U2158 (N_2158,N_1306,In_78);
or U2159 (N_2159,N_1876,N_1262);
xnor U2160 (N_2160,N_1865,In_2237);
xor U2161 (N_2161,N_507,N_1520);
and U2162 (N_2162,N_1565,N_1852);
nor U2163 (N_2163,N_673,N_677);
nand U2164 (N_2164,N_1972,N_1844);
and U2165 (N_2165,N_1802,N_786);
or U2166 (N_2166,N_536,N_1475);
nand U2167 (N_2167,In_1608,N_912);
and U2168 (N_2168,N_11,N_1984);
nor U2169 (N_2169,N_198,N_1899);
and U2170 (N_2170,N_1867,N_206);
and U2171 (N_2171,N_1581,N_1516);
nor U2172 (N_2172,N_1901,N_1659);
xor U2173 (N_2173,N_614,N_1790);
nand U2174 (N_2174,N_1799,N_1836);
nand U2175 (N_2175,In_2108,N_1914);
nor U2176 (N_2176,N_1678,In_528);
nor U2177 (N_2177,N_1614,N_1810);
and U2178 (N_2178,In_570,N_1675);
nand U2179 (N_2179,N_820,N_1593);
xor U2180 (N_2180,N_1887,In_264);
xnor U2181 (N_2181,N_1743,N_1827);
nor U2182 (N_2182,N_1800,N_1890);
and U2183 (N_2183,N_1923,In_1611);
xor U2184 (N_2184,N_962,N_1848);
nor U2185 (N_2185,N_1842,N_1260);
nand U2186 (N_2186,N_1695,N_1689);
or U2187 (N_2187,N_1845,N_1354);
and U2188 (N_2188,N_1894,N_1910);
or U2189 (N_2189,N_1864,N_1173);
xnor U2190 (N_2190,In_2370,N_1994);
nand U2191 (N_2191,N_794,N_1139);
nor U2192 (N_2192,N_1130,N_1855);
xor U2193 (N_2193,N_1969,N_1497);
or U2194 (N_2194,N_1722,N_1751);
nor U2195 (N_2195,N_1206,N_1902);
or U2196 (N_2196,In_62,N_1891);
nor U2197 (N_2197,N_1837,N_1949);
nor U2198 (N_2198,N_1943,N_1360);
xnor U2199 (N_2199,N_577,N_1629);
or U2200 (N_2200,N_2184,N_2029);
nand U2201 (N_2201,N_2156,N_2150);
nand U2202 (N_2202,N_2147,N_2151);
nand U2203 (N_2203,N_1992,N_2049);
nor U2204 (N_2204,N_2187,N_2102);
and U2205 (N_2205,N_2176,N_2007);
xnor U2206 (N_2206,N_1931,N_2189);
and U2207 (N_2207,N_2063,N_2155);
nand U2208 (N_2208,N_355,N_2173);
or U2209 (N_2209,N_2044,N_2071);
nand U2210 (N_2210,N_1083,In_1012);
or U2211 (N_2211,N_2137,N_2115);
and U2212 (N_2212,N_2038,N_2074);
or U2213 (N_2213,N_1918,N_2105);
and U2214 (N_2214,N_2011,N_2170);
and U2215 (N_2215,N_2103,N_2160);
or U2216 (N_2216,N_1896,N_1964);
nor U2217 (N_2217,N_1439,N_2000);
or U2218 (N_2218,N_2032,N_2037);
nor U2219 (N_2219,N_1657,N_1669);
and U2220 (N_2220,N_2081,N_1809);
or U2221 (N_2221,N_1826,N_2001);
nand U2222 (N_2222,N_2169,N_2121);
nand U2223 (N_2223,N_2174,In_1247);
and U2224 (N_2224,N_2122,N_1978);
xor U2225 (N_2225,N_2139,N_2027);
nand U2226 (N_2226,N_2062,N_1055);
nand U2227 (N_2227,N_2118,N_2153);
and U2228 (N_2228,N_2191,N_2060);
nor U2229 (N_2229,N_2181,N_2177);
or U2230 (N_2230,N_804,N_2164);
nor U2231 (N_2231,N_2073,N_2019);
and U2232 (N_2232,N_1466,N_1971);
or U2233 (N_2233,N_1168,N_2086);
and U2234 (N_2234,N_833,N_2182);
nand U2235 (N_2235,N_1990,N_2085);
or U2236 (N_2236,N_2058,N_2119);
nor U2237 (N_2237,N_1868,N_2024);
xnor U2238 (N_2238,N_2140,N_2092);
and U2239 (N_2239,N_2047,N_1731);
and U2240 (N_2240,N_2075,N_2087);
and U2241 (N_2241,N_1762,N_1849);
and U2242 (N_2242,N_425,N_2022);
nor U2243 (N_2243,N_1854,In_1909);
and U2244 (N_2244,N_1888,N_494);
nand U2245 (N_2245,N_2065,N_2077);
or U2246 (N_2246,N_1959,N_2057);
xor U2247 (N_2247,N_2059,N_2040);
nand U2248 (N_2248,N_1928,N_1808);
xnor U2249 (N_2249,N_2141,N_2123);
or U2250 (N_2250,N_2113,N_1880);
nor U2251 (N_2251,N_2104,N_1908);
xnor U2252 (N_2252,N_1344,N_1879);
nor U2253 (N_2253,N_2048,N_2129);
and U2254 (N_2254,In_1138,N_2117);
and U2255 (N_2255,N_2034,N_2179);
xnor U2256 (N_2256,N_2114,N_2194);
and U2257 (N_2257,N_2076,N_2012);
xor U2258 (N_2258,N_1973,N_120);
nand U2259 (N_2259,N_1501,N_2046);
or U2260 (N_2260,N_2185,N_2133);
nand U2261 (N_2261,N_2023,N_2069);
nor U2262 (N_2262,In_1606,N_2192);
nand U2263 (N_2263,In_1192,N_2042);
nand U2264 (N_2264,N_2134,N_1711);
xnor U2265 (N_2265,N_2198,N_2107);
and U2266 (N_2266,N_2175,N_2003);
nor U2267 (N_2267,N_2013,N_2018);
nor U2268 (N_2268,N_1945,N_2142);
nor U2269 (N_2269,N_2143,N_2148);
nor U2270 (N_2270,N_2017,N_2010);
nor U2271 (N_2271,N_2083,N_1423);
xor U2272 (N_2272,N_2052,N_2193);
nand U2273 (N_2273,N_1942,N_2157);
or U2274 (N_2274,N_1941,N_2196);
nor U2275 (N_2275,N_2149,N_2068);
and U2276 (N_2276,N_2180,N_2172);
nor U2277 (N_2277,N_2014,N_2199);
nand U2278 (N_2278,N_2090,N_1831);
and U2279 (N_2279,N_1552,N_2144);
or U2280 (N_2280,N_2162,N_2171);
xor U2281 (N_2281,N_284,N_2099);
xor U2282 (N_2282,N_1696,N_2043);
nand U2283 (N_2283,N_691,N_2135);
and U2284 (N_2284,N_2120,N_1859);
and U2285 (N_2285,N_2030,N_2015);
or U2286 (N_2286,N_2056,N_2124);
or U2287 (N_2287,N_2067,N_2091);
nor U2288 (N_2288,N_2009,N_1861);
nor U2289 (N_2289,N_2021,N_2039);
nand U2290 (N_2290,N_1138,N_1817);
or U2291 (N_2291,N_1937,N_2097);
and U2292 (N_2292,N_2112,N_2095);
nand U2293 (N_2293,N_2008,N_1633);
or U2294 (N_2294,N_2002,N_1885);
xor U2295 (N_2295,N_2020,N_1966);
nor U2296 (N_2296,N_2109,N_1628);
nand U2297 (N_2297,N_2078,N_1983);
nor U2298 (N_2298,N_2146,N_2152);
and U2299 (N_2299,N_93,N_1866);
nor U2300 (N_2300,In_870,In_2093);
nand U2301 (N_2301,In_2257,N_1968);
nand U2302 (N_2302,N_2035,N_1787);
and U2303 (N_2303,N_1457,N_2004);
xor U2304 (N_2304,N_2158,N_2033);
or U2305 (N_2305,N_1634,N_716);
or U2306 (N_2306,N_1824,N_2054);
and U2307 (N_2307,N_1755,N_1585);
xor U2308 (N_2308,N_2111,N_2082);
xnor U2309 (N_2309,N_2110,N_2166);
nand U2310 (N_2310,N_2006,N_2050);
nor U2311 (N_2311,N_1986,N_1814);
nand U2312 (N_2312,N_2190,N_2167);
and U2313 (N_2313,N_2064,N_1974);
and U2314 (N_2314,N_2168,N_2061);
and U2315 (N_2315,N_1688,N_420);
and U2316 (N_2316,N_2036,N_2125);
and U2317 (N_2317,N_2098,N_2093);
nand U2318 (N_2318,N_2138,N_1985);
or U2319 (N_2319,N_2197,N_2094);
xor U2320 (N_2320,N_2188,N_2072);
nor U2321 (N_2321,In_1436,N_2088);
nor U2322 (N_2322,N_2128,N_2096);
and U2323 (N_2323,N_1841,N_2186);
nor U2324 (N_2324,N_1927,N_1916);
and U2325 (N_2325,N_2136,N_1275);
nand U2326 (N_2326,N_1546,N_2159);
nor U2327 (N_2327,N_2165,N_2116);
and U2328 (N_2328,N_2100,N_2079);
nand U2329 (N_2329,N_2055,N_2005);
or U2330 (N_2330,N_2145,N_1954);
xnor U2331 (N_2331,N_2132,N_2026);
and U2332 (N_2332,N_2028,N_2127);
or U2333 (N_2333,N_2106,N_2016);
nand U2334 (N_2334,N_2051,N_1087);
xor U2335 (N_2335,N_29,N_2126);
xor U2336 (N_2336,N_2084,In_129);
xor U2337 (N_2337,N_2154,In_1978);
nor U2338 (N_2338,N_2163,N_0);
nor U2339 (N_2339,N_2183,N_2108);
xnor U2340 (N_2340,N_2101,N_2070);
and U2341 (N_2341,N_2161,N_1656);
xnor U2342 (N_2342,N_2053,N_2066);
nor U2343 (N_2343,N_2080,N_1797);
xor U2344 (N_2344,N_992,N_1061);
nor U2345 (N_2345,N_2195,N_2178);
and U2346 (N_2346,N_2031,N_2131);
nand U2347 (N_2347,N_2130,N_2089);
xnor U2348 (N_2348,N_2025,N_1874);
nor U2349 (N_2349,N_2045,N_2041);
nor U2350 (N_2350,N_2023,N_1696);
xor U2351 (N_2351,N_716,N_2010);
and U2352 (N_2352,N_1879,N_2177);
nor U2353 (N_2353,N_1983,N_2011);
xnor U2354 (N_2354,N_1423,N_2054);
nor U2355 (N_2355,N_2162,N_2003);
and U2356 (N_2356,N_2019,N_2022);
xnor U2357 (N_2357,N_2007,N_2179);
nand U2358 (N_2358,N_2155,N_2030);
and U2359 (N_2359,N_2187,N_2043);
nand U2360 (N_2360,N_2100,N_2037);
nand U2361 (N_2361,N_2184,N_2138);
xor U2362 (N_2362,N_2014,N_2139);
xnor U2363 (N_2363,N_804,N_2094);
or U2364 (N_2364,N_2083,N_2199);
and U2365 (N_2365,N_2143,N_2188);
nor U2366 (N_2366,N_2190,N_2184);
and U2367 (N_2367,N_2140,N_2136);
and U2368 (N_2368,N_2132,N_1888);
nand U2369 (N_2369,N_2111,N_2015);
and U2370 (N_2370,N_2054,N_2135);
nand U2371 (N_2371,N_1945,N_2069);
nand U2372 (N_2372,N_2136,N_1656);
xor U2373 (N_2373,N_2021,N_2043);
nand U2374 (N_2374,N_804,N_2123);
and U2375 (N_2375,N_1824,N_1731);
and U2376 (N_2376,N_2192,N_1896);
or U2377 (N_2377,N_2173,N_1854);
nor U2378 (N_2378,N_2172,N_2079);
xnor U2379 (N_2379,N_2009,N_2199);
and U2380 (N_2380,N_2054,N_2092);
and U2381 (N_2381,N_1731,N_2005);
or U2382 (N_2382,N_1888,N_2144);
xnor U2383 (N_2383,N_2136,N_2127);
nand U2384 (N_2384,N_2168,N_2115);
and U2385 (N_2385,N_2157,N_1809);
or U2386 (N_2386,N_2118,N_2003);
and U2387 (N_2387,N_2115,N_2095);
or U2388 (N_2388,N_691,N_2126);
and U2389 (N_2389,N_2032,N_2123);
nor U2390 (N_2390,N_1908,N_2105);
nand U2391 (N_2391,N_2117,N_2105);
nor U2392 (N_2392,N_2059,N_2052);
nand U2393 (N_2393,N_1501,N_2182);
nand U2394 (N_2394,N_355,N_1826);
and U2395 (N_2395,N_2177,N_2087);
xnor U2396 (N_2396,N_2088,N_2098);
xor U2397 (N_2397,N_2125,N_284);
nand U2398 (N_2398,N_2096,N_2168);
nor U2399 (N_2399,N_1824,N_2017);
nand U2400 (N_2400,N_2305,N_2355);
or U2401 (N_2401,N_2360,N_2388);
and U2402 (N_2402,N_2343,N_2251);
nand U2403 (N_2403,N_2242,N_2308);
and U2404 (N_2404,N_2259,N_2203);
nor U2405 (N_2405,N_2255,N_2312);
or U2406 (N_2406,N_2279,N_2366);
or U2407 (N_2407,N_2336,N_2219);
or U2408 (N_2408,N_2359,N_2322);
or U2409 (N_2409,N_2392,N_2281);
nor U2410 (N_2410,N_2361,N_2250);
nor U2411 (N_2411,N_2221,N_2233);
xnor U2412 (N_2412,N_2228,N_2260);
nor U2413 (N_2413,N_2254,N_2362);
or U2414 (N_2414,N_2277,N_2289);
nor U2415 (N_2415,N_2396,N_2363);
or U2416 (N_2416,N_2399,N_2364);
nand U2417 (N_2417,N_2280,N_2339);
xnor U2418 (N_2418,N_2344,N_2301);
or U2419 (N_2419,N_2303,N_2218);
or U2420 (N_2420,N_2356,N_2377);
xnor U2421 (N_2421,N_2236,N_2341);
xnor U2422 (N_2422,N_2306,N_2394);
or U2423 (N_2423,N_2370,N_2235);
nor U2424 (N_2424,N_2201,N_2249);
or U2425 (N_2425,N_2342,N_2263);
nand U2426 (N_2426,N_2224,N_2398);
and U2427 (N_2427,N_2348,N_2294);
and U2428 (N_2428,N_2223,N_2207);
nor U2429 (N_2429,N_2220,N_2213);
xnor U2430 (N_2430,N_2371,N_2243);
nor U2431 (N_2431,N_2258,N_2252);
or U2432 (N_2432,N_2321,N_2372);
xor U2433 (N_2433,N_2317,N_2212);
nand U2434 (N_2434,N_2315,N_2205);
and U2435 (N_2435,N_2332,N_2202);
xor U2436 (N_2436,N_2314,N_2264);
and U2437 (N_2437,N_2239,N_2271);
xnor U2438 (N_2438,N_2318,N_2253);
nor U2439 (N_2439,N_2267,N_2387);
and U2440 (N_2440,N_2351,N_2240);
or U2441 (N_2441,N_2381,N_2204);
nand U2442 (N_2442,N_2266,N_2230);
or U2443 (N_2443,N_2310,N_2272);
or U2444 (N_2444,N_2304,N_2347);
and U2445 (N_2445,N_2323,N_2302);
nand U2446 (N_2446,N_2273,N_2328);
nor U2447 (N_2447,N_2345,N_2295);
or U2448 (N_2448,N_2285,N_2278);
or U2449 (N_2449,N_2313,N_2270);
and U2450 (N_2450,N_2275,N_2241);
nand U2451 (N_2451,N_2214,N_2375);
nor U2452 (N_2452,N_2385,N_2261);
xor U2453 (N_2453,N_2324,N_2293);
or U2454 (N_2454,N_2291,N_2299);
nand U2455 (N_2455,N_2300,N_2282);
and U2456 (N_2456,N_2311,N_2217);
nor U2457 (N_2457,N_2382,N_2244);
xnor U2458 (N_2458,N_2206,N_2290);
and U2459 (N_2459,N_2379,N_2376);
or U2460 (N_2460,N_2330,N_2286);
nor U2461 (N_2461,N_2354,N_2390);
or U2462 (N_2462,N_2262,N_2333);
nor U2463 (N_2463,N_2393,N_2391);
and U2464 (N_2464,N_2209,N_2357);
and U2465 (N_2465,N_2231,N_2319);
nor U2466 (N_2466,N_2352,N_2232);
and U2467 (N_2467,N_2208,N_2326);
and U2468 (N_2468,N_2349,N_2340);
or U2469 (N_2469,N_2383,N_2316);
xnor U2470 (N_2470,N_2229,N_2397);
xnor U2471 (N_2471,N_2380,N_2374);
or U2472 (N_2472,N_2327,N_2337);
nor U2473 (N_2473,N_2325,N_2269);
nor U2474 (N_2474,N_2265,N_2225);
or U2475 (N_2475,N_2395,N_2338);
nand U2476 (N_2476,N_2222,N_2353);
and U2477 (N_2477,N_2248,N_2296);
nand U2478 (N_2478,N_2226,N_2274);
xor U2479 (N_2479,N_2256,N_2384);
nand U2480 (N_2480,N_2329,N_2386);
and U2481 (N_2481,N_2215,N_2238);
xnor U2482 (N_2482,N_2210,N_2350);
or U2483 (N_2483,N_2245,N_2257);
xnor U2484 (N_2484,N_2346,N_2292);
nand U2485 (N_2485,N_2246,N_2227);
nand U2486 (N_2486,N_2358,N_2283);
and U2487 (N_2487,N_2378,N_2268);
nor U2488 (N_2488,N_2334,N_2320);
nor U2489 (N_2489,N_2276,N_2309);
or U2490 (N_2490,N_2211,N_2216);
nand U2491 (N_2491,N_2247,N_2234);
or U2492 (N_2492,N_2287,N_2373);
nor U2493 (N_2493,N_2367,N_2331);
or U2494 (N_2494,N_2368,N_2365);
nand U2495 (N_2495,N_2237,N_2200);
nor U2496 (N_2496,N_2389,N_2369);
xnor U2497 (N_2497,N_2297,N_2284);
or U2498 (N_2498,N_2307,N_2288);
and U2499 (N_2499,N_2335,N_2298);
nand U2500 (N_2500,N_2272,N_2387);
and U2501 (N_2501,N_2250,N_2252);
nor U2502 (N_2502,N_2298,N_2220);
nor U2503 (N_2503,N_2328,N_2224);
nand U2504 (N_2504,N_2347,N_2261);
and U2505 (N_2505,N_2297,N_2280);
xor U2506 (N_2506,N_2338,N_2377);
or U2507 (N_2507,N_2227,N_2376);
and U2508 (N_2508,N_2347,N_2328);
nor U2509 (N_2509,N_2332,N_2255);
or U2510 (N_2510,N_2375,N_2282);
and U2511 (N_2511,N_2390,N_2300);
nand U2512 (N_2512,N_2306,N_2357);
and U2513 (N_2513,N_2302,N_2282);
or U2514 (N_2514,N_2258,N_2347);
nand U2515 (N_2515,N_2219,N_2296);
nor U2516 (N_2516,N_2311,N_2375);
or U2517 (N_2517,N_2323,N_2347);
nor U2518 (N_2518,N_2390,N_2218);
nand U2519 (N_2519,N_2211,N_2326);
nor U2520 (N_2520,N_2314,N_2239);
xor U2521 (N_2521,N_2235,N_2305);
or U2522 (N_2522,N_2362,N_2218);
nand U2523 (N_2523,N_2230,N_2275);
nand U2524 (N_2524,N_2378,N_2223);
or U2525 (N_2525,N_2241,N_2298);
and U2526 (N_2526,N_2266,N_2274);
or U2527 (N_2527,N_2361,N_2305);
nand U2528 (N_2528,N_2367,N_2385);
or U2529 (N_2529,N_2377,N_2394);
or U2530 (N_2530,N_2343,N_2302);
xnor U2531 (N_2531,N_2362,N_2235);
and U2532 (N_2532,N_2328,N_2352);
or U2533 (N_2533,N_2307,N_2398);
nor U2534 (N_2534,N_2244,N_2300);
nor U2535 (N_2535,N_2384,N_2398);
or U2536 (N_2536,N_2269,N_2340);
nor U2537 (N_2537,N_2205,N_2386);
and U2538 (N_2538,N_2398,N_2238);
nor U2539 (N_2539,N_2347,N_2203);
nor U2540 (N_2540,N_2372,N_2207);
and U2541 (N_2541,N_2213,N_2261);
nor U2542 (N_2542,N_2321,N_2225);
and U2543 (N_2543,N_2379,N_2340);
nor U2544 (N_2544,N_2232,N_2363);
and U2545 (N_2545,N_2202,N_2318);
nor U2546 (N_2546,N_2343,N_2348);
and U2547 (N_2547,N_2312,N_2388);
nor U2548 (N_2548,N_2301,N_2355);
nand U2549 (N_2549,N_2252,N_2212);
or U2550 (N_2550,N_2206,N_2296);
or U2551 (N_2551,N_2213,N_2379);
and U2552 (N_2552,N_2387,N_2307);
and U2553 (N_2553,N_2358,N_2256);
xor U2554 (N_2554,N_2340,N_2280);
nor U2555 (N_2555,N_2206,N_2268);
and U2556 (N_2556,N_2397,N_2357);
xnor U2557 (N_2557,N_2235,N_2272);
xnor U2558 (N_2558,N_2330,N_2361);
nand U2559 (N_2559,N_2361,N_2265);
or U2560 (N_2560,N_2399,N_2248);
xor U2561 (N_2561,N_2299,N_2345);
nand U2562 (N_2562,N_2280,N_2286);
or U2563 (N_2563,N_2366,N_2275);
and U2564 (N_2564,N_2277,N_2212);
and U2565 (N_2565,N_2303,N_2244);
or U2566 (N_2566,N_2220,N_2295);
nor U2567 (N_2567,N_2211,N_2287);
nand U2568 (N_2568,N_2318,N_2234);
nand U2569 (N_2569,N_2326,N_2265);
nor U2570 (N_2570,N_2383,N_2366);
nor U2571 (N_2571,N_2303,N_2217);
nand U2572 (N_2572,N_2229,N_2303);
nor U2573 (N_2573,N_2359,N_2396);
and U2574 (N_2574,N_2261,N_2315);
xnor U2575 (N_2575,N_2266,N_2299);
xnor U2576 (N_2576,N_2389,N_2365);
xnor U2577 (N_2577,N_2315,N_2227);
xor U2578 (N_2578,N_2248,N_2220);
or U2579 (N_2579,N_2232,N_2358);
nand U2580 (N_2580,N_2345,N_2390);
nor U2581 (N_2581,N_2301,N_2292);
or U2582 (N_2582,N_2302,N_2303);
and U2583 (N_2583,N_2334,N_2315);
nor U2584 (N_2584,N_2247,N_2212);
and U2585 (N_2585,N_2339,N_2232);
nand U2586 (N_2586,N_2395,N_2224);
nand U2587 (N_2587,N_2332,N_2334);
nor U2588 (N_2588,N_2270,N_2277);
nand U2589 (N_2589,N_2256,N_2351);
nand U2590 (N_2590,N_2315,N_2383);
or U2591 (N_2591,N_2327,N_2349);
nor U2592 (N_2592,N_2235,N_2203);
and U2593 (N_2593,N_2378,N_2217);
and U2594 (N_2594,N_2359,N_2306);
or U2595 (N_2595,N_2383,N_2389);
and U2596 (N_2596,N_2393,N_2280);
xor U2597 (N_2597,N_2341,N_2233);
nand U2598 (N_2598,N_2218,N_2313);
and U2599 (N_2599,N_2357,N_2310);
or U2600 (N_2600,N_2595,N_2521);
and U2601 (N_2601,N_2453,N_2518);
and U2602 (N_2602,N_2420,N_2427);
and U2603 (N_2603,N_2436,N_2487);
or U2604 (N_2604,N_2559,N_2474);
nor U2605 (N_2605,N_2426,N_2432);
xor U2606 (N_2606,N_2570,N_2440);
nand U2607 (N_2607,N_2523,N_2552);
xor U2608 (N_2608,N_2499,N_2478);
or U2609 (N_2609,N_2409,N_2539);
nor U2610 (N_2610,N_2462,N_2491);
nor U2611 (N_2611,N_2567,N_2533);
and U2612 (N_2612,N_2415,N_2592);
nand U2613 (N_2613,N_2553,N_2482);
nor U2614 (N_2614,N_2502,N_2524);
nor U2615 (N_2615,N_2546,N_2484);
or U2616 (N_2616,N_2438,N_2483);
nand U2617 (N_2617,N_2517,N_2446);
nor U2618 (N_2618,N_2434,N_2461);
nor U2619 (N_2619,N_2503,N_2562);
xnor U2620 (N_2620,N_2443,N_2405);
nor U2621 (N_2621,N_2451,N_2560);
nor U2622 (N_2622,N_2515,N_2413);
xor U2623 (N_2623,N_2442,N_2454);
and U2624 (N_2624,N_2508,N_2568);
nand U2625 (N_2625,N_2460,N_2536);
or U2626 (N_2626,N_2537,N_2526);
and U2627 (N_2627,N_2444,N_2489);
nand U2628 (N_2628,N_2516,N_2572);
nor U2629 (N_2629,N_2410,N_2469);
nor U2630 (N_2630,N_2419,N_2540);
or U2631 (N_2631,N_2557,N_2598);
or U2632 (N_2632,N_2425,N_2479);
nor U2633 (N_2633,N_2582,N_2578);
or U2634 (N_2634,N_2428,N_2447);
xnor U2635 (N_2635,N_2556,N_2541);
or U2636 (N_2636,N_2543,N_2450);
xor U2637 (N_2637,N_2531,N_2538);
nor U2638 (N_2638,N_2457,N_2441);
and U2639 (N_2639,N_2558,N_2509);
and U2640 (N_2640,N_2527,N_2514);
or U2641 (N_2641,N_2576,N_2510);
and U2642 (N_2642,N_2455,N_2548);
nand U2643 (N_2643,N_2593,N_2501);
nand U2644 (N_2644,N_2472,N_2412);
nand U2645 (N_2645,N_2403,N_2530);
xnor U2646 (N_2646,N_2549,N_2481);
nor U2647 (N_2647,N_2414,N_2470);
nand U2648 (N_2648,N_2555,N_2411);
nor U2649 (N_2649,N_2416,N_2590);
nand U2650 (N_2650,N_2587,N_2554);
and U2651 (N_2651,N_2421,N_2506);
and U2652 (N_2652,N_2542,N_2563);
nand U2653 (N_2653,N_2594,N_2597);
nand U2654 (N_2654,N_2429,N_2465);
nor U2655 (N_2655,N_2439,N_2473);
and U2656 (N_2656,N_2423,N_2494);
nor U2657 (N_2657,N_2433,N_2456);
or U2658 (N_2658,N_2529,N_2458);
nor U2659 (N_2659,N_2519,N_2532);
or U2660 (N_2660,N_2586,N_2512);
and U2661 (N_2661,N_2596,N_2485);
nor U2662 (N_2662,N_2545,N_2430);
nand U2663 (N_2663,N_2476,N_2422);
nand U2664 (N_2664,N_2401,N_2564);
nand U2665 (N_2665,N_2589,N_2488);
xnor U2666 (N_2666,N_2581,N_2561);
xnor U2667 (N_2667,N_2466,N_2575);
nand U2668 (N_2668,N_2467,N_2477);
or U2669 (N_2669,N_2551,N_2402);
or U2670 (N_2670,N_2580,N_2573);
and U2671 (N_2671,N_2585,N_2475);
xnor U2672 (N_2672,N_2497,N_2407);
nor U2673 (N_2673,N_2535,N_2550);
or U2674 (N_2674,N_2464,N_2449);
nand U2675 (N_2675,N_2500,N_2471);
nand U2676 (N_2676,N_2404,N_2431);
and U2677 (N_2677,N_2507,N_2498);
and U2678 (N_2678,N_2584,N_2408);
nor U2679 (N_2679,N_2406,N_2493);
nand U2680 (N_2680,N_2591,N_2486);
and U2681 (N_2681,N_2463,N_2599);
nor U2682 (N_2682,N_2424,N_2492);
nor U2683 (N_2683,N_2490,N_2566);
or U2684 (N_2684,N_2496,N_2480);
nand U2685 (N_2685,N_2520,N_2435);
nand U2686 (N_2686,N_2534,N_2565);
or U2687 (N_2687,N_2448,N_2525);
xnor U2688 (N_2688,N_2571,N_2522);
nor U2689 (N_2689,N_2437,N_2579);
xor U2690 (N_2690,N_2588,N_2544);
and U2691 (N_2691,N_2528,N_2505);
and U2692 (N_2692,N_2400,N_2574);
nand U2693 (N_2693,N_2468,N_2495);
nor U2694 (N_2694,N_2547,N_2417);
nor U2695 (N_2695,N_2569,N_2459);
nor U2696 (N_2696,N_2583,N_2445);
xor U2697 (N_2697,N_2513,N_2418);
nand U2698 (N_2698,N_2452,N_2504);
and U2699 (N_2699,N_2577,N_2511);
or U2700 (N_2700,N_2548,N_2572);
nor U2701 (N_2701,N_2599,N_2545);
xor U2702 (N_2702,N_2549,N_2577);
xor U2703 (N_2703,N_2581,N_2590);
or U2704 (N_2704,N_2561,N_2536);
or U2705 (N_2705,N_2550,N_2487);
and U2706 (N_2706,N_2590,N_2579);
and U2707 (N_2707,N_2481,N_2516);
xnor U2708 (N_2708,N_2469,N_2549);
and U2709 (N_2709,N_2489,N_2466);
and U2710 (N_2710,N_2512,N_2574);
xnor U2711 (N_2711,N_2445,N_2575);
nor U2712 (N_2712,N_2554,N_2490);
nor U2713 (N_2713,N_2576,N_2497);
nand U2714 (N_2714,N_2484,N_2443);
nor U2715 (N_2715,N_2508,N_2587);
xnor U2716 (N_2716,N_2427,N_2434);
and U2717 (N_2717,N_2451,N_2524);
nand U2718 (N_2718,N_2567,N_2505);
xnor U2719 (N_2719,N_2477,N_2433);
nand U2720 (N_2720,N_2447,N_2486);
nor U2721 (N_2721,N_2513,N_2498);
xor U2722 (N_2722,N_2553,N_2579);
xor U2723 (N_2723,N_2462,N_2469);
xnor U2724 (N_2724,N_2589,N_2593);
and U2725 (N_2725,N_2456,N_2539);
and U2726 (N_2726,N_2434,N_2493);
nand U2727 (N_2727,N_2480,N_2486);
or U2728 (N_2728,N_2474,N_2449);
xor U2729 (N_2729,N_2408,N_2455);
nor U2730 (N_2730,N_2589,N_2547);
nor U2731 (N_2731,N_2451,N_2542);
nor U2732 (N_2732,N_2463,N_2462);
or U2733 (N_2733,N_2481,N_2511);
xor U2734 (N_2734,N_2595,N_2409);
nor U2735 (N_2735,N_2474,N_2410);
and U2736 (N_2736,N_2403,N_2534);
nor U2737 (N_2737,N_2501,N_2460);
and U2738 (N_2738,N_2477,N_2453);
nor U2739 (N_2739,N_2429,N_2561);
xor U2740 (N_2740,N_2425,N_2514);
xor U2741 (N_2741,N_2534,N_2483);
nor U2742 (N_2742,N_2460,N_2431);
and U2743 (N_2743,N_2472,N_2455);
nand U2744 (N_2744,N_2582,N_2432);
and U2745 (N_2745,N_2478,N_2434);
xnor U2746 (N_2746,N_2418,N_2443);
and U2747 (N_2747,N_2539,N_2537);
or U2748 (N_2748,N_2468,N_2471);
xor U2749 (N_2749,N_2470,N_2538);
and U2750 (N_2750,N_2402,N_2488);
or U2751 (N_2751,N_2596,N_2409);
or U2752 (N_2752,N_2440,N_2451);
nand U2753 (N_2753,N_2573,N_2514);
and U2754 (N_2754,N_2484,N_2403);
and U2755 (N_2755,N_2447,N_2457);
xnor U2756 (N_2756,N_2414,N_2599);
or U2757 (N_2757,N_2562,N_2548);
nand U2758 (N_2758,N_2420,N_2429);
nor U2759 (N_2759,N_2485,N_2521);
xnor U2760 (N_2760,N_2494,N_2407);
or U2761 (N_2761,N_2463,N_2532);
nor U2762 (N_2762,N_2581,N_2567);
xor U2763 (N_2763,N_2541,N_2510);
xor U2764 (N_2764,N_2508,N_2576);
or U2765 (N_2765,N_2589,N_2438);
or U2766 (N_2766,N_2472,N_2440);
nor U2767 (N_2767,N_2572,N_2555);
nand U2768 (N_2768,N_2496,N_2454);
or U2769 (N_2769,N_2412,N_2466);
or U2770 (N_2770,N_2475,N_2403);
xnor U2771 (N_2771,N_2564,N_2412);
nor U2772 (N_2772,N_2530,N_2535);
and U2773 (N_2773,N_2568,N_2495);
nand U2774 (N_2774,N_2435,N_2480);
or U2775 (N_2775,N_2489,N_2463);
xnor U2776 (N_2776,N_2430,N_2444);
and U2777 (N_2777,N_2428,N_2525);
nor U2778 (N_2778,N_2414,N_2512);
xnor U2779 (N_2779,N_2483,N_2527);
xor U2780 (N_2780,N_2478,N_2439);
nand U2781 (N_2781,N_2452,N_2583);
nand U2782 (N_2782,N_2487,N_2594);
xor U2783 (N_2783,N_2574,N_2485);
nand U2784 (N_2784,N_2425,N_2511);
xnor U2785 (N_2785,N_2579,N_2460);
or U2786 (N_2786,N_2479,N_2478);
and U2787 (N_2787,N_2577,N_2515);
nand U2788 (N_2788,N_2558,N_2568);
nor U2789 (N_2789,N_2492,N_2527);
and U2790 (N_2790,N_2484,N_2547);
nor U2791 (N_2791,N_2513,N_2465);
and U2792 (N_2792,N_2536,N_2594);
nand U2793 (N_2793,N_2421,N_2571);
and U2794 (N_2794,N_2401,N_2463);
xor U2795 (N_2795,N_2485,N_2559);
or U2796 (N_2796,N_2575,N_2589);
xor U2797 (N_2797,N_2401,N_2444);
or U2798 (N_2798,N_2496,N_2477);
nand U2799 (N_2799,N_2452,N_2581);
xnor U2800 (N_2800,N_2741,N_2790);
and U2801 (N_2801,N_2622,N_2670);
or U2802 (N_2802,N_2648,N_2700);
nor U2803 (N_2803,N_2632,N_2638);
nand U2804 (N_2804,N_2631,N_2663);
or U2805 (N_2805,N_2653,N_2644);
or U2806 (N_2806,N_2623,N_2633);
and U2807 (N_2807,N_2765,N_2776);
or U2808 (N_2808,N_2699,N_2789);
xor U2809 (N_2809,N_2715,N_2779);
and U2810 (N_2810,N_2636,N_2620);
xor U2811 (N_2811,N_2796,N_2701);
nor U2812 (N_2812,N_2756,N_2630);
xnor U2813 (N_2813,N_2769,N_2680);
nor U2814 (N_2814,N_2608,N_2637);
or U2815 (N_2815,N_2786,N_2723);
nand U2816 (N_2816,N_2752,N_2654);
nor U2817 (N_2817,N_2649,N_2783);
and U2818 (N_2818,N_2628,N_2621);
nor U2819 (N_2819,N_2661,N_2727);
nand U2820 (N_2820,N_2774,N_2736);
nand U2821 (N_2821,N_2662,N_2791);
nand U2822 (N_2822,N_2696,N_2728);
and U2823 (N_2823,N_2753,N_2611);
nand U2824 (N_2824,N_2754,N_2751);
or U2825 (N_2825,N_2665,N_2619);
xnor U2826 (N_2826,N_2777,N_2685);
nand U2827 (N_2827,N_2759,N_2625);
nand U2828 (N_2828,N_2764,N_2758);
and U2829 (N_2829,N_2677,N_2612);
xor U2830 (N_2830,N_2771,N_2650);
and U2831 (N_2831,N_2775,N_2749);
nand U2832 (N_2832,N_2626,N_2799);
xor U2833 (N_2833,N_2613,N_2610);
and U2834 (N_2834,N_2675,N_2747);
and U2835 (N_2835,N_2710,N_2683);
nand U2836 (N_2836,N_2725,N_2798);
or U2837 (N_2837,N_2716,N_2643);
and U2838 (N_2838,N_2651,N_2645);
xor U2839 (N_2839,N_2690,N_2718);
or U2840 (N_2840,N_2618,N_2748);
nand U2841 (N_2841,N_2688,N_2770);
xor U2842 (N_2842,N_2714,N_2713);
or U2843 (N_2843,N_2604,N_2672);
nand U2844 (N_2844,N_2787,N_2763);
nor U2845 (N_2845,N_2682,N_2689);
and U2846 (N_2846,N_2657,N_2659);
nand U2847 (N_2847,N_2743,N_2703);
and U2848 (N_2848,N_2660,N_2724);
xor U2849 (N_2849,N_2746,N_2635);
xor U2850 (N_2850,N_2684,N_2772);
xor U2851 (N_2851,N_2629,N_2679);
or U2852 (N_2852,N_2707,N_2755);
or U2853 (N_2853,N_2721,N_2600);
nand U2854 (N_2854,N_2793,N_2706);
xnor U2855 (N_2855,N_2607,N_2784);
nand U2856 (N_2856,N_2687,N_2639);
or U2857 (N_2857,N_2615,N_2726);
xor U2858 (N_2858,N_2691,N_2674);
nand U2859 (N_2859,N_2795,N_2719);
xor U2860 (N_2860,N_2780,N_2722);
xor U2861 (N_2861,N_2602,N_2609);
and U2862 (N_2862,N_2603,N_2734);
or U2863 (N_2863,N_2750,N_2617);
or U2864 (N_2864,N_2761,N_2708);
nor U2865 (N_2865,N_2788,N_2616);
and U2866 (N_2866,N_2642,N_2739);
nor U2867 (N_2867,N_2656,N_2712);
or U2868 (N_2868,N_2720,N_2605);
and U2869 (N_2869,N_2705,N_2695);
nor U2870 (N_2870,N_2792,N_2737);
nor U2871 (N_2871,N_2673,N_2697);
xor U2872 (N_2872,N_2767,N_2666);
and U2873 (N_2873,N_2732,N_2797);
or U2874 (N_2874,N_2669,N_2729);
xor U2875 (N_2875,N_2778,N_2676);
or U2876 (N_2876,N_2733,N_2702);
or U2877 (N_2877,N_2773,N_2785);
and U2878 (N_2878,N_2717,N_2641);
nor U2879 (N_2879,N_2693,N_2782);
or U2880 (N_2880,N_2614,N_2757);
and U2881 (N_2881,N_2735,N_2731);
nand U2882 (N_2882,N_2768,N_2667);
and U2883 (N_2883,N_2601,N_2738);
nand U2884 (N_2884,N_2742,N_2709);
nand U2885 (N_2885,N_2681,N_2794);
or U2886 (N_2886,N_2655,N_2781);
or U2887 (N_2887,N_2762,N_2686);
and U2888 (N_2888,N_2698,N_2652);
nand U2889 (N_2889,N_2704,N_2627);
xnor U2890 (N_2890,N_2634,N_2606);
nor U2891 (N_2891,N_2694,N_2678);
nor U2892 (N_2892,N_2745,N_2646);
xnor U2893 (N_2893,N_2664,N_2640);
and U2894 (N_2894,N_2740,N_2624);
or U2895 (N_2895,N_2766,N_2692);
xnor U2896 (N_2896,N_2711,N_2647);
or U2897 (N_2897,N_2671,N_2730);
nand U2898 (N_2898,N_2744,N_2668);
xnor U2899 (N_2899,N_2658,N_2760);
nor U2900 (N_2900,N_2646,N_2694);
xnor U2901 (N_2901,N_2604,N_2733);
nor U2902 (N_2902,N_2622,N_2633);
and U2903 (N_2903,N_2633,N_2763);
and U2904 (N_2904,N_2660,N_2644);
xnor U2905 (N_2905,N_2603,N_2750);
nand U2906 (N_2906,N_2754,N_2676);
nor U2907 (N_2907,N_2647,N_2673);
and U2908 (N_2908,N_2723,N_2764);
nand U2909 (N_2909,N_2703,N_2675);
nand U2910 (N_2910,N_2751,N_2606);
and U2911 (N_2911,N_2768,N_2728);
nand U2912 (N_2912,N_2778,N_2632);
nor U2913 (N_2913,N_2615,N_2735);
or U2914 (N_2914,N_2690,N_2720);
nand U2915 (N_2915,N_2719,N_2631);
xor U2916 (N_2916,N_2675,N_2643);
and U2917 (N_2917,N_2688,N_2746);
and U2918 (N_2918,N_2716,N_2730);
or U2919 (N_2919,N_2727,N_2678);
or U2920 (N_2920,N_2766,N_2627);
nand U2921 (N_2921,N_2654,N_2642);
nand U2922 (N_2922,N_2785,N_2629);
and U2923 (N_2923,N_2646,N_2728);
nand U2924 (N_2924,N_2639,N_2702);
nand U2925 (N_2925,N_2657,N_2623);
nor U2926 (N_2926,N_2692,N_2711);
and U2927 (N_2927,N_2601,N_2718);
nor U2928 (N_2928,N_2765,N_2667);
xnor U2929 (N_2929,N_2639,N_2707);
or U2930 (N_2930,N_2687,N_2737);
xor U2931 (N_2931,N_2639,N_2718);
nor U2932 (N_2932,N_2764,N_2785);
nor U2933 (N_2933,N_2699,N_2610);
xnor U2934 (N_2934,N_2722,N_2697);
nor U2935 (N_2935,N_2697,N_2601);
xor U2936 (N_2936,N_2705,N_2684);
nand U2937 (N_2937,N_2758,N_2737);
and U2938 (N_2938,N_2761,N_2643);
nor U2939 (N_2939,N_2786,N_2705);
nor U2940 (N_2940,N_2707,N_2715);
nor U2941 (N_2941,N_2665,N_2714);
or U2942 (N_2942,N_2776,N_2626);
nand U2943 (N_2943,N_2750,N_2609);
or U2944 (N_2944,N_2615,N_2678);
and U2945 (N_2945,N_2668,N_2708);
nand U2946 (N_2946,N_2600,N_2779);
or U2947 (N_2947,N_2719,N_2793);
xnor U2948 (N_2948,N_2635,N_2662);
xor U2949 (N_2949,N_2628,N_2603);
and U2950 (N_2950,N_2716,N_2606);
or U2951 (N_2951,N_2611,N_2635);
or U2952 (N_2952,N_2759,N_2607);
and U2953 (N_2953,N_2674,N_2618);
or U2954 (N_2954,N_2762,N_2630);
or U2955 (N_2955,N_2708,N_2758);
or U2956 (N_2956,N_2732,N_2607);
nor U2957 (N_2957,N_2617,N_2630);
nand U2958 (N_2958,N_2746,N_2710);
nand U2959 (N_2959,N_2793,N_2742);
or U2960 (N_2960,N_2662,N_2673);
and U2961 (N_2961,N_2631,N_2723);
nand U2962 (N_2962,N_2723,N_2777);
nor U2963 (N_2963,N_2708,N_2607);
nand U2964 (N_2964,N_2773,N_2713);
nor U2965 (N_2965,N_2764,N_2690);
nor U2966 (N_2966,N_2663,N_2625);
nand U2967 (N_2967,N_2761,N_2676);
nand U2968 (N_2968,N_2623,N_2762);
nand U2969 (N_2969,N_2771,N_2697);
xor U2970 (N_2970,N_2631,N_2693);
and U2971 (N_2971,N_2740,N_2717);
or U2972 (N_2972,N_2681,N_2672);
xor U2973 (N_2973,N_2663,N_2715);
or U2974 (N_2974,N_2613,N_2713);
nand U2975 (N_2975,N_2614,N_2760);
and U2976 (N_2976,N_2783,N_2678);
and U2977 (N_2977,N_2718,N_2659);
or U2978 (N_2978,N_2708,N_2706);
and U2979 (N_2979,N_2684,N_2680);
nor U2980 (N_2980,N_2620,N_2704);
nand U2981 (N_2981,N_2749,N_2766);
nor U2982 (N_2982,N_2702,N_2738);
and U2983 (N_2983,N_2767,N_2677);
or U2984 (N_2984,N_2658,N_2765);
and U2985 (N_2985,N_2630,N_2707);
xnor U2986 (N_2986,N_2620,N_2710);
nor U2987 (N_2987,N_2725,N_2626);
or U2988 (N_2988,N_2665,N_2701);
nor U2989 (N_2989,N_2638,N_2601);
nor U2990 (N_2990,N_2674,N_2729);
or U2991 (N_2991,N_2739,N_2732);
and U2992 (N_2992,N_2781,N_2715);
nor U2993 (N_2993,N_2634,N_2702);
xnor U2994 (N_2994,N_2736,N_2622);
or U2995 (N_2995,N_2790,N_2695);
nand U2996 (N_2996,N_2639,N_2714);
nor U2997 (N_2997,N_2612,N_2694);
nand U2998 (N_2998,N_2693,N_2753);
nor U2999 (N_2999,N_2746,N_2772);
xor U3000 (N_3000,N_2893,N_2975);
or U3001 (N_3001,N_2926,N_2974);
or U3002 (N_3002,N_2971,N_2873);
nand U3003 (N_3003,N_2827,N_2900);
and U3004 (N_3004,N_2833,N_2991);
and U3005 (N_3005,N_2892,N_2826);
or U3006 (N_3006,N_2931,N_2929);
and U3007 (N_3007,N_2885,N_2865);
or U3008 (N_3008,N_2895,N_2949);
nor U3009 (N_3009,N_2845,N_2838);
or U3010 (N_3010,N_2839,N_2836);
xor U3011 (N_3011,N_2829,N_2902);
and U3012 (N_3012,N_2808,N_2846);
nor U3013 (N_3013,N_2901,N_2913);
nand U3014 (N_3014,N_2921,N_2855);
xnor U3015 (N_3015,N_2994,N_2987);
nand U3016 (N_3016,N_2939,N_2946);
and U3017 (N_3017,N_2867,N_2807);
nand U3018 (N_3018,N_2822,N_2915);
nand U3019 (N_3019,N_2878,N_2819);
or U3020 (N_3020,N_2925,N_2831);
nand U3021 (N_3021,N_2993,N_2961);
or U3022 (N_3022,N_2945,N_2872);
nor U3023 (N_3023,N_2898,N_2928);
or U3024 (N_3024,N_2924,N_2851);
nor U3025 (N_3025,N_2979,N_2957);
nor U3026 (N_3026,N_2909,N_2992);
or U3027 (N_3027,N_2857,N_2950);
and U3028 (N_3028,N_2881,N_2815);
nor U3029 (N_3029,N_2968,N_2882);
nor U3030 (N_3030,N_2932,N_2821);
xnor U3031 (N_3031,N_2964,N_2800);
xnor U3032 (N_3032,N_2868,N_2955);
nand U3033 (N_3033,N_2880,N_2983);
or U3034 (N_3034,N_2914,N_2848);
or U3035 (N_3035,N_2875,N_2804);
nand U3036 (N_3036,N_2956,N_2859);
nor U3037 (N_3037,N_2918,N_2896);
nor U3038 (N_3038,N_2816,N_2934);
or U3039 (N_3039,N_2911,N_2830);
nor U3040 (N_3040,N_2995,N_2876);
nor U3041 (N_3041,N_2986,N_2920);
and U3042 (N_3042,N_2990,N_2814);
or U3043 (N_3043,N_2935,N_2801);
or U3044 (N_3044,N_2907,N_2905);
xor U3045 (N_3045,N_2812,N_2840);
nand U3046 (N_3046,N_2863,N_2809);
nand U3047 (N_3047,N_2847,N_2982);
and U3048 (N_3048,N_2954,N_2817);
and U3049 (N_3049,N_2943,N_2823);
nor U3050 (N_3050,N_2874,N_2985);
or U3051 (N_3051,N_2835,N_2960);
nor U3052 (N_3052,N_2866,N_2852);
and U3053 (N_3053,N_2832,N_2988);
and U3054 (N_3054,N_2977,N_2912);
nand U3055 (N_3055,N_2941,N_2999);
and U3056 (N_3056,N_2879,N_2825);
nor U3057 (N_3057,N_2891,N_2903);
nor U3058 (N_3058,N_2978,N_2937);
or U3059 (N_3059,N_2916,N_2818);
xnor U3060 (N_3060,N_2938,N_2853);
or U3061 (N_3061,N_2856,N_2810);
and U3062 (N_3062,N_2894,N_2989);
and U3063 (N_3063,N_2862,N_2890);
nand U3064 (N_3064,N_2972,N_2843);
nor U3065 (N_3065,N_2861,N_2919);
nand U3066 (N_3066,N_2869,N_2927);
and U3067 (N_3067,N_2886,N_2922);
and U3068 (N_3068,N_2969,N_2813);
nand U3069 (N_3069,N_2811,N_2981);
and U3070 (N_3070,N_2837,N_2802);
and U3071 (N_3071,N_2998,N_2834);
or U3072 (N_3072,N_2959,N_2951);
xor U3073 (N_3073,N_2963,N_2970);
nand U3074 (N_3074,N_2850,N_2897);
or U3075 (N_3075,N_2858,N_2883);
nor U3076 (N_3076,N_2820,N_2967);
xor U3077 (N_3077,N_2980,N_2854);
nand U3078 (N_3078,N_2803,N_2887);
xor U3079 (N_3079,N_2888,N_2864);
and U3080 (N_3080,N_2976,N_2884);
and U3081 (N_3081,N_2849,N_2910);
nor U3082 (N_3082,N_2944,N_2997);
nor U3083 (N_3083,N_2973,N_2966);
xnor U3084 (N_3084,N_2940,N_2923);
nand U3085 (N_3085,N_2953,N_2952);
or U3086 (N_3086,N_2933,N_2870);
or U3087 (N_3087,N_2860,N_2842);
and U3088 (N_3088,N_2844,N_2828);
or U3089 (N_3089,N_2906,N_2899);
or U3090 (N_3090,N_2877,N_2947);
nor U3091 (N_3091,N_2908,N_2936);
xor U3092 (N_3092,N_2996,N_2824);
xnor U3093 (N_3093,N_2917,N_2871);
nand U3094 (N_3094,N_2984,N_2889);
and U3095 (N_3095,N_2958,N_2942);
xor U3096 (N_3096,N_2962,N_2904);
xnor U3097 (N_3097,N_2841,N_2930);
or U3098 (N_3098,N_2805,N_2806);
or U3099 (N_3099,N_2965,N_2948);
nand U3100 (N_3100,N_2841,N_2817);
and U3101 (N_3101,N_2877,N_2982);
and U3102 (N_3102,N_2854,N_2958);
and U3103 (N_3103,N_2930,N_2807);
and U3104 (N_3104,N_2933,N_2816);
nand U3105 (N_3105,N_2828,N_2992);
and U3106 (N_3106,N_2841,N_2871);
nand U3107 (N_3107,N_2894,N_2945);
and U3108 (N_3108,N_2885,N_2804);
nor U3109 (N_3109,N_2981,N_2886);
nand U3110 (N_3110,N_2958,N_2851);
nand U3111 (N_3111,N_2859,N_2851);
and U3112 (N_3112,N_2839,N_2826);
nor U3113 (N_3113,N_2855,N_2960);
xnor U3114 (N_3114,N_2943,N_2837);
xnor U3115 (N_3115,N_2928,N_2872);
and U3116 (N_3116,N_2943,N_2817);
xor U3117 (N_3117,N_2874,N_2889);
nor U3118 (N_3118,N_2976,N_2929);
nand U3119 (N_3119,N_2927,N_2923);
and U3120 (N_3120,N_2900,N_2971);
nor U3121 (N_3121,N_2926,N_2936);
xor U3122 (N_3122,N_2996,N_2951);
nand U3123 (N_3123,N_2913,N_2912);
xor U3124 (N_3124,N_2901,N_2886);
and U3125 (N_3125,N_2863,N_2956);
nand U3126 (N_3126,N_2916,N_2893);
and U3127 (N_3127,N_2904,N_2988);
nor U3128 (N_3128,N_2860,N_2978);
xnor U3129 (N_3129,N_2906,N_2866);
nor U3130 (N_3130,N_2920,N_2963);
nand U3131 (N_3131,N_2905,N_2829);
or U3132 (N_3132,N_2847,N_2891);
and U3133 (N_3133,N_2860,N_2920);
xnor U3134 (N_3134,N_2815,N_2849);
and U3135 (N_3135,N_2986,N_2851);
and U3136 (N_3136,N_2893,N_2819);
and U3137 (N_3137,N_2947,N_2852);
and U3138 (N_3138,N_2815,N_2915);
nand U3139 (N_3139,N_2860,N_2912);
xor U3140 (N_3140,N_2846,N_2891);
nor U3141 (N_3141,N_2895,N_2963);
or U3142 (N_3142,N_2918,N_2891);
nor U3143 (N_3143,N_2990,N_2887);
xnor U3144 (N_3144,N_2900,N_2864);
or U3145 (N_3145,N_2865,N_2973);
nor U3146 (N_3146,N_2931,N_2901);
nand U3147 (N_3147,N_2802,N_2942);
xnor U3148 (N_3148,N_2858,N_2851);
xnor U3149 (N_3149,N_2915,N_2895);
xor U3150 (N_3150,N_2969,N_2911);
and U3151 (N_3151,N_2911,N_2937);
nor U3152 (N_3152,N_2824,N_2861);
xnor U3153 (N_3153,N_2957,N_2840);
xnor U3154 (N_3154,N_2886,N_2960);
nand U3155 (N_3155,N_2873,N_2862);
xnor U3156 (N_3156,N_2825,N_2922);
or U3157 (N_3157,N_2903,N_2938);
or U3158 (N_3158,N_2984,N_2885);
xnor U3159 (N_3159,N_2970,N_2805);
xor U3160 (N_3160,N_2880,N_2914);
nand U3161 (N_3161,N_2865,N_2956);
and U3162 (N_3162,N_2866,N_2987);
nor U3163 (N_3163,N_2983,N_2819);
nor U3164 (N_3164,N_2944,N_2898);
nand U3165 (N_3165,N_2935,N_2833);
and U3166 (N_3166,N_2934,N_2948);
nand U3167 (N_3167,N_2887,N_2849);
and U3168 (N_3168,N_2999,N_2887);
xor U3169 (N_3169,N_2979,N_2939);
nand U3170 (N_3170,N_2858,N_2885);
xor U3171 (N_3171,N_2980,N_2897);
nor U3172 (N_3172,N_2887,N_2926);
nor U3173 (N_3173,N_2927,N_2863);
or U3174 (N_3174,N_2873,N_2851);
nand U3175 (N_3175,N_2839,N_2875);
and U3176 (N_3176,N_2864,N_2822);
and U3177 (N_3177,N_2957,N_2927);
xor U3178 (N_3178,N_2885,N_2893);
xor U3179 (N_3179,N_2911,N_2824);
and U3180 (N_3180,N_2896,N_2814);
xor U3181 (N_3181,N_2834,N_2822);
and U3182 (N_3182,N_2970,N_2860);
nand U3183 (N_3183,N_2935,N_2989);
nand U3184 (N_3184,N_2871,N_2890);
or U3185 (N_3185,N_2877,N_2975);
nand U3186 (N_3186,N_2898,N_2998);
nor U3187 (N_3187,N_2934,N_2898);
nor U3188 (N_3188,N_2841,N_2823);
nand U3189 (N_3189,N_2991,N_2990);
xor U3190 (N_3190,N_2958,N_2909);
xor U3191 (N_3191,N_2823,N_2994);
or U3192 (N_3192,N_2968,N_2921);
nor U3193 (N_3193,N_2831,N_2938);
and U3194 (N_3194,N_2929,N_2843);
nor U3195 (N_3195,N_2802,N_2801);
nand U3196 (N_3196,N_2888,N_2840);
and U3197 (N_3197,N_2948,N_2827);
or U3198 (N_3198,N_2947,N_2828);
nor U3199 (N_3199,N_2804,N_2890);
xnor U3200 (N_3200,N_3152,N_3138);
nand U3201 (N_3201,N_3162,N_3098);
nor U3202 (N_3202,N_3159,N_3108);
xnor U3203 (N_3203,N_3051,N_3131);
and U3204 (N_3204,N_3189,N_3004);
nor U3205 (N_3205,N_3082,N_3022);
nand U3206 (N_3206,N_3062,N_3199);
or U3207 (N_3207,N_3115,N_3101);
xnor U3208 (N_3208,N_3096,N_3192);
and U3209 (N_3209,N_3070,N_3044);
and U3210 (N_3210,N_3064,N_3078);
xor U3211 (N_3211,N_3126,N_3030);
xnor U3212 (N_3212,N_3128,N_3157);
or U3213 (N_3213,N_3144,N_3017);
and U3214 (N_3214,N_3155,N_3151);
nand U3215 (N_3215,N_3085,N_3196);
nor U3216 (N_3216,N_3120,N_3088);
nor U3217 (N_3217,N_3198,N_3186);
and U3218 (N_3218,N_3054,N_3055);
and U3219 (N_3219,N_3160,N_3073);
nand U3220 (N_3220,N_3146,N_3080);
nand U3221 (N_3221,N_3041,N_3086);
xor U3222 (N_3222,N_3066,N_3117);
or U3223 (N_3223,N_3188,N_3009);
or U3224 (N_3224,N_3110,N_3191);
or U3225 (N_3225,N_3037,N_3149);
nor U3226 (N_3226,N_3053,N_3076);
or U3227 (N_3227,N_3165,N_3141);
or U3228 (N_3228,N_3031,N_3087);
nand U3229 (N_3229,N_3173,N_3020);
nor U3230 (N_3230,N_3172,N_3068);
or U3231 (N_3231,N_3019,N_3118);
or U3232 (N_3232,N_3002,N_3097);
or U3233 (N_3233,N_3021,N_3140);
nand U3234 (N_3234,N_3023,N_3099);
nor U3235 (N_3235,N_3018,N_3190);
xor U3236 (N_3236,N_3167,N_3125);
nand U3237 (N_3237,N_3181,N_3038);
or U3238 (N_3238,N_3012,N_3061);
nand U3239 (N_3239,N_3119,N_3195);
or U3240 (N_3240,N_3164,N_3049);
xnor U3241 (N_3241,N_3001,N_3133);
and U3242 (N_3242,N_3089,N_3102);
or U3243 (N_3243,N_3067,N_3175);
nor U3244 (N_3244,N_3079,N_3077);
xnor U3245 (N_3245,N_3043,N_3123);
or U3246 (N_3246,N_3168,N_3193);
nand U3247 (N_3247,N_3011,N_3134);
nand U3248 (N_3248,N_3033,N_3107);
and U3249 (N_3249,N_3035,N_3136);
nor U3250 (N_3250,N_3187,N_3130);
and U3251 (N_3251,N_3100,N_3007);
xor U3252 (N_3252,N_3046,N_3059);
xnor U3253 (N_3253,N_3015,N_3025);
nor U3254 (N_3254,N_3135,N_3180);
and U3255 (N_3255,N_3006,N_3153);
xnor U3256 (N_3256,N_3045,N_3042);
nand U3257 (N_3257,N_3161,N_3026);
nand U3258 (N_3258,N_3048,N_3127);
nor U3259 (N_3259,N_3150,N_3013);
nor U3260 (N_3260,N_3032,N_3095);
and U3261 (N_3261,N_3036,N_3103);
nor U3262 (N_3262,N_3094,N_3072);
nand U3263 (N_3263,N_3116,N_3163);
xor U3264 (N_3264,N_3091,N_3005);
nand U3265 (N_3265,N_3174,N_3142);
or U3266 (N_3266,N_3111,N_3063);
nand U3267 (N_3267,N_3084,N_3197);
nor U3268 (N_3268,N_3178,N_3122);
nand U3269 (N_3269,N_3093,N_3171);
nor U3270 (N_3270,N_3081,N_3158);
and U3271 (N_3271,N_3039,N_3003);
or U3272 (N_3272,N_3132,N_3124);
nand U3273 (N_3273,N_3145,N_3027);
xor U3274 (N_3274,N_3182,N_3139);
xnor U3275 (N_3275,N_3069,N_3154);
or U3276 (N_3276,N_3166,N_3074);
xnor U3277 (N_3277,N_3092,N_3137);
or U3278 (N_3278,N_3113,N_3156);
and U3279 (N_3279,N_3000,N_3040);
nand U3280 (N_3280,N_3010,N_3028);
nor U3281 (N_3281,N_3143,N_3075);
and U3282 (N_3282,N_3029,N_3176);
nand U3283 (N_3283,N_3052,N_3034);
xnor U3284 (N_3284,N_3185,N_3016);
or U3285 (N_3285,N_3184,N_3083);
xor U3286 (N_3286,N_3183,N_3058);
nor U3287 (N_3287,N_3106,N_3014);
or U3288 (N_3288,N_3104,N_3169);
or U3289 (N_3289,N_3109,N_3047);
or U3290 (N_3290,N_3177,N_3024);
xnor U3291 (N_3291,N_3057,N_3121);
or U3292 (N_3292,N_3060,N_3148);
nor U3293 (N_3293,N_3065,N_3090);
and U3294 (N_3294,N_3170,N_3129);
nand U3295 (N_3295,N_3147,N_3105);
and U3296 (N_3296,N_3008,N_3050);
nor U3297 (N_3297,N_3056,N_3114);
nand U3298 (N_3298,N_3179,N_3194);
nor U3299 (N_3299,N_3071,N_3112);
and U3300 (N_3300,N_3171,N_3058);
or U3301 (N_3301,N_3191,N_3134);
xor U3302 (N_3302,N_3147,N_3099);
nand U3303 (N_3303,N_3172,N_3023);
and U3304 (N_3304,N_3083,N_3029);
nor U3305 (N_3305,N_3094,N_3000);
nand U3306 (N_3306,N_3057,N_3027);
nand U3307 (N_3307,N_3055,N_3003);
xor U3308 (N_3308,N_3101,N_3184);
xor U3309 (N_3309,N_3105,N_3135);
xor U3310 (N_3310,N_3182,N_3097);
nor U3311 (N_3311,N_3051,N_3094);
nor U3312 (N_3312,N_3103,N_3123);
nor U3313 (N_3313,N_3089,N_3112);
nand U3314 (N_3314,N_3025,N_3104);
xnor U3315 (N_3315,N_3198,N_3022);
and U3316 (N_3316,N_3182,N_3087);
nand U3317 (N_3317,N_3060,N_3180);
and U3318 (N_3318,N_3006,N_3035);
or U3319 (N_3319,N_3079,N_3140);
xor U3320 (N_3320,N_3125,N_3153);
or U3321 (N_3321,N_3186,N_3106);
nor U3322 (N_3322,N_3011,N_3106);
nand U3323 (N_3323,N_3022,N_3020);
nor U3324 (N_3324,N_3031,N_3164);
nor U3325 (N_3325,N_3158,N_3116);
nor U3326 (N_3326,N_3170,N_3039);
xor U3327 (N_3327,N_3180,N_3148);
xor U3328 (N_3328,N_3121,N_3028);
xor U3329 (N_3329,N_3083,N_3127);
nand U3330 (N_3330,N_3193,N_3197);
xor U3331 (N_3331,N_3049,N_3099);
and U3332 (N_3332,N_3141,N_3090);
nor U3333 (N_3333,N_3019,N_3125);
xor U3334 (N_3334,N_3184,N_3060);
xor U3335 (N_3335,N_3178,N_3197);
nor U3336 (N_3336,N_3014,N_3175);
or U3337 (N_3337,N_3003,N_3071);
or U3338 (N_3338,N_3123,N_3186);
and U3339 (N_3339,N_3063,N_3156);
nor U3340 (N_3340,N_3076,N_3075);
and U3341 (N_3341,N_3157,N_3180);
xor U3342 (N_3342,N_3185,N_3097);
nor U3343 (N_3343,N_3047,N_3121);
nand U3344 (N_3344,N_3123,N_3018);
nor U3345 (N_3345,N_3177,N_3011);
and U3346 (N_3346,N_3010,N_3160);
nand U3347 (N_3347,N_3012,N_3068);
nand U3348 (N_3348,N_3189,N_3061);
or U3349 (N_3349,N_3071,N_3189);
nor U3350 (N_3350,N_3130,N_3163);
and U3351 (N_3351,N_3086,N_3046);
or U3352 (N_3352,N_3197,N_3065);
or U3353 (N_3353,N_3017,N_3081);
or U3354 (N_3354,N_3020,N_3064);
xor U3355 (N_3355,N_3036,N_3045);
nand U3356 (N_3356,N_3099,N_3051);
and U3357 (N_3357,N_3166,N_3137);
nor U3358 (N_3358,N_3159,N_3014);
xor U3359 (N_3359,N_3158,N_3015);
and U3360 (N_3360,N_3035,N_3071);
xnor U3361 (N_3361,N_3042,N_3085);
or U3362 (N_3362,N_3151,N_3103);
or U3363 (N_3363,N_3066,N_3120);
nor U3364 (N_3364,N_3022,N_3059);
and U3365 (N_3365,N_3069,N_3175);
or U3366 (N_3366,N_3099,N_3015);
nor U3367 (N_3367,N_3120,N_3191);
and U3368 (N_3368,N_3066,N_3060);
nor U3369 (N_3369,N_3117,N_3055);
nand U3370 (N_3370,N_3000,N_3093);
nand U3371 (N_3371,N_3038,N_3175);
or U3372 (N_3372,N_3053,N_3035);
or U3373 (N_3373,N_3196,N_3118);
and U3374 (N_3374,N_3075,N_3102);
and U3375 (N_3375,N_3144,N_3117);
nand U3376 (N_3376,N_3017,N_3127);
nor U3377 (N_3377,N_3058,N_3128);
nor U3378 (N_3378,N_3039,N_3032);
nand U3379 (N_3379,N_3099,N_3093);
xnor U3380 (N_3380,N_3159,N_3186);
or U3381 (N_3381,N_3025,N_3199);
xnor U3382 (N_3382,N_3111,N_3062);
and U3383 (N_3383,N_3122,N_3171);
and U3384 (N_3384,N_3013,N_3008);
nand U3385 (N_3385,N_3170,N_3010);
and U3386 (N_3386,N_3116,N_3127);
xnor U3387 (N_3387,N_3030,N_3059);
nor U3388 (N_3388,N_3018,N_3172);
or U3389 (N_3389,N_3052,N_3022);
nand U3390 (N_3390,N_3118,N_3110);
nand U3391 (N_3391,N_3046,N_3138);
and U3392 (N_3392,N_3055,N_3145);
nand U3393 (N_3393,N_3119,N_3156);
nand U3394 (N_3394,N_3056,N_3071);
nor U3395 (N_3395,N_3175,N_3070);
or U3396 (N_3396,N_3183,N_3175);
xnor U3397 (N_3397,N_3103,N_3061);
nor U3398 (N_3398,N_3099,N_3066);
or U3399 (N_3399,N_3055,N_3183);
or U3400 (N_3400,N_3296,N_3236);
nand U3401 (N_3401,N_3216,N_3309);
nand U3402 (N_3402,N_3294,N_3240);
nand U3403 (N_3403,N_3267,N_3223);
and U3404 (N_3404,N_3200,N_3331);
and U3405 (N_3405,N_3318,N_3237);
xnor U3406 (N_3406,N_3242,N_3396);
nor U3407 (N_3407,N_3367,N_3293);
xnor U3408 (N_3408,N_3299,N_3230);
or U3409 (N_3409,N_3364,N_3370);
and U3410 (N_3410,N_3284,N_3297);
xor U3411 (N_3411,N_3311,N_3202);
nand U3412 (N_3412,N_3306,N_3265);
or U3413 (N_3413,N_3390,N_3330);
xnor U3414 (N_3414,N_3234,N_3208);
nand U3415 (N_3415,N_3385,N_3273);
or U3416 (N_3416,N_3361,N_3372);
and U3417 (N_3417,N_3206,N_3269);
nor U3418 (N_3418,N_3247,N_3352);
nand U3419 (N_3419,N_3212,N_3277);
nand U3420 (N_3420,N_3347,N_3376);
and U3421 (N_3421,N_3368,N_3349);
nand U3422 (N_3422,N_3259,N_3374);
nor U3423 (N_3423,N_3335,N_3345);
xor U3424 (N_3424,N_3399,N_3346);
nor U3425 (N_3425,N_3220,N_3365);
and U3426 (N_3426,N_3351,N_3298);
and U3427 (N_3427,N_3302,N_3384);
and U3428 (N_3428,N_3389,N_3283);
nand U3429 (N_3429,N_3257,N_3360);
or U3430 (N_3430,N_3334,N_3362);
and U3431 (N_3431,N_3343,N_3313);
nor U3432 (N_3432,N_3300,N_3373);
xor U3433 (N_3433,N_3369,N_3337);
nand U3434 (N_3434,N_3244,N_3336);
nand U3435 (N_3435,N_3214,N_3217);
nor U3436 (N_3436,N_3357,N_3204);
or U3437 (N_3437,N_3316,N_3276);
nand U3438 (N_3438,N_3226,N_3323);
xnor U3439 (N_3439,N_3201,N_3387);
and U3440 (N_3440,N_3232,N_3210);
nand U3441 (N_3441,N_3315,N_3308);
and U3442 (N_3442,N_3388,N_3326);
nand U3443 (N_3443,N_3270,N_3227);
xor U3444 (N_3444,N_3224,N_3295);
and U3445 (N_3445,N_3281,N_3286);
nor U3446 (N_3446,N_3325,N_3246);
nand U3447 (N_3447,N_3391,N_3222);
nand U3448 (N_3448,N_3339,N_3386);
nand U3449 (N_3449,N_3287,N_3307);
or U3450 (N_3450,N_3203,N_3310);
or U3451 (N_3451,N_3383,N_3393);
or U3452 (N_3452,N_3243,N_3312);
or U3453 (N_3453,N_3380,N_3348);
xnor U3454 (N_3454,N_3285,N_3272);
xnor U3455 (N_3455,N_3342,N_3278);
nor U3456 (N_3456,N_3356,N_3241);
xor U3457 (N_3457,N_3274,N_3324);
nand U3458 (N_3458,N_3350,N_3397);
and U3459 (N_3459,N_3275,N_3303);
and U3460 (N_3460,N_3262,N_3394);
nand U3461 (N_3461,N_3250,N_3215);
nand U3462 (N_3462,N_3205,N_3377);
nand U3463 (N_3463,N_3255,N_3305);
or U3464 (N_3464,N_3353,N_3245);
xnor U3465 (N_3465,N_3379,N_3225);
xor U3466 (N_3466,N_3378,N_3258);
or U3467 (N_3467,N_3218,N_3366);
or U3468 (N_3468,N_3340,N_3291);
nand U3469 (N_3469,N_3261,N_3332);
and U3470 (N_3470,N_3253,N_3280);
nor U3471 (N_3471,N_3292,N_3327);
or U3472 (N_3472,N_3333,N_3231);
nand U3473 (N_3473,N_3375,N_3322);
xor U3474 (N_3474,N_3358,N_3359);
nor U3475 (N_3475,N_3282,N_3252);
or U3476 (N_3476,N_3354,N_3314);
xor U3477 (N_3477,N_3338,N_3256);
nor U3478 (N_3478,N_3251,N_3392);
nand U3479 (N_3479,N_3211,N_3395);
xnor U3480 (N_3480,N_3355,N_3329);
or U3481 (N_3481,N_3233,N_3371);
and U3482 (N_3482,N_3239,N_3279);
nor U3483 (N_3483,N_3320,N_3317);
and U3484 (N_3484,N_3228,N_3304);
or U3485 (N_3485,N_3249,N_3207);
nand U3486 (N_3486,N_3381,N_3264);
nor U3487 (N_3487,N_3271,N_3229);
xor U3488 (N_3488,N_3248,N_3219);
nor U3489 (N_3489,N_3235,N_3268);
nor U3490 (N_3490,N_3289,N_3209);
nor U3491 (N_3491,N_3254,N_3363);
nor U3492 (N_3492,N_3328,N_3238);
nand U3493 (N_3493,N_3382,N_3301);
or U3494 (N_3494,N_3260,N_3321);
xnor U3495 (N_3495,N_3221,N_3398);
or U3496 (N_3496,N_3290,N_3288);
or U3497 (N_3497,N_3263,N_3266);
nor U3498 (N_3498,N_3344,N_3213);
xnor U3499 (N_3499,N_3341,N_3319);
or U3500 (N_3500,N_3309,N_3232);
xnor U3501 (N_3501,N_3234,N_3211);
nor U3502 (N_3502,N_3391,N_3206);
or U3503 (N_3503,N_3243,N_3297);
and U3504 (N_3504,N_3283,N_3307);
xnor U3505 (N_3505,N_3366,N_3309);
xnor U3506 (N_3506,N_3209,N_3332);
nor U3507 (N_3507,N_3213,N_3363);
nand U3508 (N_3508,N_3291,N_3218);
nor U3509 (N_3509,N_3327,N_3363);
xor U3510 (N_3510,N_3256,N_3213);
nor U3511 (N_3511,N_3350,N_3382);
nand U3512 (N_3512,N_3269,N_3372);
nand U3513 (N_3513,N_3210,N_3346);
xnor U3514 (N_3514,N_3310,N_3341);
and U3515 (N_3515,N_3207,N_3215);
xnor U3516 (N_3516,N_3302,N_3340);
xnor U3517 (N_3517,N_3396,N_3252);
and U3518 (N_3518,N_3398,N_3291);
or U3519 (N_3519,N_3350,N_3333);
nor U3520 (N_3520,N_3225,N_3321);
nor U3521 (N_3521,N_3361,N_3390);
and U3522 (N_3522,N_3246,N_3322);
xnor U3523 (N_3523,N_3277,N_3230);
and U3524 (N_3524,N_3280,N_3316);
or U3525 (N_3525,N_3344,N_3374);
or U3526 (N_3526,N_3380,N_3314);
nand U3527 (N_3527,N_3304,N_3363);
and U3528 (N_3528,N_3296,N_3331);
nand U3529 (N_3529,N_3294,N_3356);
xor U3530 (N_3530,N_3292,N_3363);
nand U3531 (N_3531,N_3332,N_3235);
or U3532 (N_3532,N_3212,N_3247);
nor U3533 (N_3533,N_3241,N_3254);
nand U3534 (N_3534,N_3334,N_3229);
nor U3535 (N_3535,N_3215,N_3255);
and U3536 (N_3536,N_3230,N_3312);
xnor U3537 (N_3537,N_3266,N_3368);
nor U3538 (N_3538,N_3387,N_3210);
nor U3539 (N_3539,N_3319,N_3249);
nand U3540 (N_3540,N_3247,N_3263);
xor U3541 (N_3541,N_3205,N_3298);
nor U3542 (N_3542,N_3371,N_3224);
nor U3543 (N_3543,N_3347,N_3340);
or U3544 (N_3544,N_3217,N_3212);
and U3545 (N_3545,N_3221,N_3324);
and U3546 (N_3546,N_3342,N_3373);
nand U3547 (N_3547,N_3227,N_3279);
nor U3548 (N_3548,N_3228,N_3235);
or U3549 (N_3549,N_3349,N_3364);
nor U3550 (N_3550,N_3213,N_3371);
or U3551 (N_3551,N_3385,N_3218);
xor U3552 (N_3552,N_3222,N_3311);
xor U3553 (N_3553,N_3386,N_3243);
nor U3554 (N_3554,N_3366,N_3227);
xor U3555 (N_3555,N_3326,N_3364);
xnor U3556 (N_3556,N_3377,N_3215);
nor U3557 (N_3557,N_3250,N_3239);
or U3558 (N_3558,N_3210,N_3297);
xnor U3559 (N_3559,N_3300,N_3243);
and U3560 (N_3560,N_3396,N_3333);
nor U3561 (N_3561,N_3218,N_3259);
nand U3562 (N_3562,N_3243,N_3320);
or U3563 (N_3563,N_3350,N_3219);
xnor U3564 (N_3564,N_3277,N_3250);
nand U3565 (N_3565,N_3374,N_3387);
or U3566 (N_3566,N_3318,N_3329);
xnor U3567 (N_3567,N_3218,N_3354);
or U3568 (N_3568,N_3206,N_3361);
nor U3569 (N_3569,N_3308,N_3275);
xnor U3570 (N_3570,N_3304,N_3233);
and U3571 (N_3571,N_3205,N_3246);
xor U3572 (N_3572,N_3267,N_3381);
and U3573 (N_3573,N_3332,N_3284);
nor U3574 (N_3574,N_3370,N_3262);
or U3575 (N_3575,N_3362,N_3368);
or U3576 (N_3576,N_3396,N_3278);
and U3577 (N_3577,N_3201,N_3211);
nand U3578 (N_3578,N_3214,N_3389);
xor U3579 (N_3579,N_3358,N_3242);
nand U3580 (N_3580,N_3274,N_3320);
nor U3581 (N_3581,N_3329,N_3310);
nor U3582 (N_3582,N_3261,N_3223);
xnor U3583 (N_3583,N_3266,N_3379);
nor U3584 (N_3584,N_3289,N_3296);
nor U3585 (N_3585,N_3278,N_3229);
nand U3586 (N_3586,N_3362,N_3373);
and U3587 (N_3587,N_3227,N_3363);
xor U3588 (N_3588,N_3326,N_3303);
nand U3589 (N_3589,N_3335,N_3210);
xnor U3590 (N_3590,N_3215,N_3204);
nor U3591 (N_3591,N_3300,N_3325);
xnor U3592 (N_3592,N_3352,N_3396);
nand U3593 (N_3593,N_3231,N_3395);
xor U3594 (N_3594,N_3317,N_3283);
or U3595 (N_3595,N_3243,N_3232);
or U3596 (N_3596,N_3333,N_3220);
nand U3597 (N_3597,N_3310,N_3212);
or U3598 (N_3598,N_3338,N_3339);
xnor U3599 (N_3599,N_3311,N_3245);
nand U3600 (N_3600,N_3434,N_3494);
xor U3601 (N_3601,N_3573,N_3410);
nand U3602 (N_3602,N_3577,N_3499);
xnor U3603 (N_3603,N_3433,N_3580);
or U3604 (N_3604,N_3563,N_3482);
or U3605 (N_3605,N_3404,N_3422);
and U3606 (N_3606,N_3441,N_3464);
nor U3607 (N_3607,N_3564,N_3590);
xor U3608 (N_3608,N_3436,N_3487);
or U3609 (N_3609,N_3475,N_3593);
nor U3610 (N_3610,N_3540,N_3570);
nand U3611 (N_3611,N_3530,N_3560);
nand U3612 (N_3612,N_3510,N_3412);
or U3613 (N_3613,N_3443,N_3448);
and U3614 (N_3614,N_3445,N_3595);
xor U3615 (N_3615,N_3428,N_3546);
and U3616 (N_3616,N_3496,N_3416);
or U3617 (N_3617,N_3501,N_3488);
nand U3618 (N_3618,N_3551,N_3437);
xor U3619 (N_3619,N_3431,N_3402);
and U3620 (N_3620,N_3552,N_3489);
xnor U3621 (N_3621,N_3584,N_3537);
or U3622 (N_3622,N_3506,N_3513);
and U3623 (N_3623,N_3451,N_3414);
or U3624 (N_3624,N_3524,N_3481);
or U3625 (N_3625,N_3541,N_3518);
xor U3626 (N_3626,N_3531,N_3574);
and U3627 (N_3627,N_3472,N_3596);
xnor U3628 (N_3628,N_3405,N_3559);
nor U3629 (N_3629,N_3533,N_3585);
or U3630 (N_3630,N_3539,N_3588);
xnor U3631 (N_3631,N_3519,N_3523);
nand U3632 (N_3632,N_3421,N_3424);
nand U3633 (N_3633,N_3480,N_3446);
xor U3634 (N_3634,N_3592,N_3490);
nor U3635 (N_3635,N_3581,N_3558);
or U3636 (N_3636,N_3430,N_3575);
or U3637 (N_3637,N_3548,N_3538);
xnor U3638 (N_3638,N_3442,N_3527);
nand U3639 (N_3639,N_3586,N_3543);
and U3640 (N_3640,N_3400,N_3429);
and U3641 (N_3641,N_3555,N_3497);
or U3642 (N_3642,N_3417,N_3526);
nor U3643 (N_3643,N_3589,N_3521);
or U3644 (N_3644,N_3520,N_3484);
and U3645 (N_3645,N_3572,N_3425);
and U3646 (N_3646,N_3544,N_3498);
nand U3647 (N_3647,N_3591,N_3495);
nor U3648 (N_3648,N_3471,N_3435);
and U3649 (N_3649,N_3568,N_3542);
or U3650 (N_3650,N_3511,N_3594);
or U3651 (N_3651,N_3411,N_3587);
nor U3652 (N_3652,N_3504,N_3505);
or U3653 (N_3653,N_3427,N_3535);
or U3654 (N_3654,N_3478,N_3469);
nor U3655 (N_3655,N_3420,N_3432);
or U3656 (N_3656,N_3565,N_3569);
nand U3657 (N_3657,N_3479,N_3525);
nand U3658 (N_3658,N_3502,N_3576);
nand U3659 (N_3659,N_3514,N_3458);
nor U3660 (N_3660,N_3406,N_3407);
nor U3661 (N_3661,N_3452,N_3419);
xnor U3662 (N_3662,N_3566,N_3578);
xor U3663 (N_3663,N_3466,N_3455);
or U3664 (N_3664,N_3461,N_3439);
xor U3665 (N_3665,N_3440,N_3508);
xor U3666 (N_3666,N_3485,N_3457);
xor U3667 (N_3667,N_3460,N_3477);
nor U3668 (N_3668,N_3597,N_3545);
or U3669 (N_3669,N_3459,N_3486);
nor U3670 (N_3670,N_3557,N_3515);
nand U3671 (N_3671,N_3522,N_3553);
nor U3672 (N_3672,N_3467,N_3536);
and U3673 (N_3673,N_3491,N_3426);
xor U3674 (N_3674,N_3423,N_3456);
nand U3675 (N_3675,N_3474,N_3550);
or U3676 (N_3676,N_3401,N_3476);
or U3677 (N_3677,N_3403,N_3447);
xnor U3678 (N_3678,N_3562,N_3468);
nand U3679 (N_3679,N_3507,N_3579);
xor U3680 (N_3680,N_3509,N_3465);
nand U3681 (N_3681,N_3438,N_3444);
nand U3682 (N_3682,N_3549,N_3554);
nand U3683 (N_3683,N_3529,N_3598);
or U3684 (N_3684,N_3450,N_3492);
nor U3685 (N_3685,N_3453,N_3582);
nand U3686 (N_3686,N_3415,N_3463);
or U3687 (N_3687,N_3483,N_3547);
nor U3688 (N_3688,N_3470,N_3462);
and U3689 (N_3689,N_3512,N_3449);
nand U3690 (N_3690,N_3517,N_3503);
and U3691 (N_3691,N_3413,N_3454);
nor U3692 (N_3692,N_3418,N_3528);
or U3693 (N_3693,N_3500,N_3532);
nand U3694 (N_3694,N_3556,N_3473);
nor U3695 (N_3695,N_3583,N_3409);
xnor U3696 (N_3696,N_3571,N_3599);
and U3697 (N_3697,N_3408,N_3561);
nor U3698 (N_3698,N_3567,N_3493);
and U3699 (N_3699,N_3534,N_3516);
or U3700 (N_3700,N_3484,N_3553);
nand U3701 (N_3701,N_3552,N_3597);
and U3702 (N_3702,N_3523,N_3429);
nand U3703 (N_3703,N_3573,N_3499);
and U3704 (N_3704,N_3456,N_3431);
xor U3705 (N_3705,N_3453,N_3569);
xor U3706 (N_3706,N_3545,N_3566);
nand U3707 (N_3707,N_3417,N_3464);
nand U3708 (N_3708,N_3437,N_3582);
nor U3709 (N_3709,N_3435,N_3417);
or U3710 (N_3710,N_3520,N_3406);
and U3711 (N_3711,N_3573,N_3524);
and U3712 (N_3712,N_3493,N_3423);
or U3713 (N_3713,N_3408,N_3462);
and U3714 (N_3714,N_3441,N_3446);
nor U3715 (N_3715,N_3467,N_3583);
or U3716 (N_3716,N_3565,N_3482);
nand U3717 (N_3717,N_3462,N_3414);
nor U3718 (N_3718,N_3556,N_3432);
xor U3719 (N_3719,N_3448,N_3408);
and U3720 (N_3720,N_3543,N_3557);
xor U3721 (N_3721,N_3591,N_3560);
nor U3722 (N_3722,N_3573,N_3566);
and U3723 (N_3723,N_3531,N_3427);
nor U3724 (N_3724,N_3527,N_3410);
or U3725 (N_3725,N_3544,N_3475);
xnor U3726 (N_3726,N_3430,N_3508);
or U3727 (N_3727,N_3493,N_3418);
nor U3728 (N_3728,N_3495,N_3469);
and U3729 (N_3729,N_3484,N_3574);
nand U3730 (N_3730,N_3486,N_3520);
nor U3731 (N_3731,N_3570,N_3498);
xor U3732 (N_3732,N_3540,N_3453);
nand U3733 (N_3733,N_3579,N_3517);
xor U3734 (N_3734,N_3593,N_3471);
xnor U3735 (N_3735,N_3526,N_3423);
nor U3736 (N_3736,N_3540,N_3475);
nor U3737 (N_3737,N_3571,N_3452);
nor U3738 (N_3738,N_3403,N_3444);
nor U3739 (N_3739,N_3449,N_3438);
and U3740 (N_3740,N_3485,N_3490);
and U3741 (N_3741,N_3418,N_3476);
nand U3742 (N_3742,N_3433,N_3522);
nor U3743 (N_3743,N_3516,N_3486);
and U3744 (N_3744,N_3483,N_3556);
nor U3745 (N_3745,N_3568,N_3554);
or U3746 (N_3746,N_3506,N_3534);
or U3747 (N_3747,N_3462,N_3574);
or U3748 (N_3748,N_3575,N_3516);
and U3749 (N_3749,N_3527,N_3454);
nand U3750 (N_3750,N_3574,N_3416);
and U3751 (N_3751,N_3513,N_3467);
or U3752 (N_3752,N_3520,N_3462);
and U3753 (N_3753,N_3400,N_3408);
nand U3754 (N_3754,N_3579,N_3505);
or U3755 (N_3755,N_3542,N_3406);
and U3756 (N_3756,N_3480,N_3442);
or U3757 (N_3757,N_3480,N_3526);
or U3758 (N_3758,N_3509,N_3503);
nor U3759 (N_3759,N_3486,N_3437);
xnor U3760 (N_3760,N_3428,N_3498);
or U3761 (N_3761,N_3444,N_3491);
and U3762 (N_3762,N_3412,N_3432);
nand U3763 (N_3763,N_3569,N_3530);
nand U3764 (N_3764,N_3437,N_3589);
xnor U3765 (N_3765,N_3477,N_3423);
or U3766 (N_3766,N_3598,N_3567);
and U3767 (N_3767,N_3535,N_3501);
and U3768 (N_3768,N_3505,N_3593);
nor U3769 (N_3769,N_3450,N_3547);
or U3770 (N_3770,N_3490,N_3452);
nor U3771 (N_3771,N_3541,N_3505);
nand U3772 (N_3772,N_3574,N_3450);
and U3773 (N_3773,N_3426,N_3488);
xor U3774 (N_3774,N_3403,N_3402);
and U3775 (N_3775,N_3529,N_3517);
or U3776 (N_3776,N_3511,N_3414);
and U3777 (N_3777,N_3477,N_3512);
xor U3778 (N_3778,N_3576,N_3574);
and U3779 (N_3779,N_3521,N_3418);
or U3780 (N_3780,N_3514,N_3505);
nor U3781 (N_3781,N_3420,N_3582);
or U3782 (N_3782,N_3543,N_3570);
nand U3783 (N_3783,N_3524,N_3501);
nor U3784 (N_3784,N_3492,N_3585);
xor U3785 (N_3785,N_3593,N_3520);
or U3786 (N_3786,N_3459,N_3411);
xnor U3787 (N_3787,N_3421,N_3478);
and U3788 (N_3788,N_3585,N_3576);
nor U3789 (N_3789,N_3432,N_3460);
nor U3790 (N_3790,N_3499,N_3463);
nor U3791 (N_3791,N_3491,N_3480);
nor U3792 (N_3792,N_3434,N_3547);
nor U3793 (N_3793,N_3464,N_3418);
nor U3794 (N_3794,N_3548,N_3523);
xnor U3795 (N_3795,N_3575,N_3442);
or U3796 (N_3796,N_3557,N_3416);
nand U3797 (N_3797,N_3424,N_3552);
or U3798 (N_3798,N_3434,N_3590);
and U3799 (N_3799,N_3489,N_3554);
nor U3800 (N_3800,N_3665,N_3651);
or U3801 (N_3801,N_3750,N_3771);
or U3802 (N_3802,N_3721,N_3763);
and U3803 (N_3803,N_3624,N_3641);
nand U3804 (N_3804,N_3616,N_3751);
or U3805 (N_3805,N_3769,N_3717);
nand U3806 (N_3806,N_3785,N_3738);
and U3807 (N_3807,N_3735,N_3797);
or U3808 (N_3808,N_3658,N_3676);
and U3809 (N_3809,N_3646,N_3737);
or U3810 (N_3810,N_3696,N_3654);
and U3811 (N_3811,N_3795,N_3663);
nor U3812 (N_3812,N_3683,N_3749);
xnor U3813 (N_3813,N_3793,N_3601);
xnor U3814 (N_3814,N_3698,N_3690);
or U3815 (N_3815,N_3762,N_3739);
xnor U3816 (N_3816,N_3635,N_3652);
or U3817 (N_3817,N_3620,N_3758);
xnor U3818 (N_3818,N_3639,N_3653);
and U3819 (N_3819,N_3714,N_3732);
or U3820 (N_3820,N_3674,N_3767);
or U3821 (N_3821,N_3669,N_3764);
xnor U3822 (N_3822,N_3789,N_3796);
nand U3823 (N_3823,N_3702,N_3727);
and U3824 (N_3824,N_3685,N_3680);
nand U3825 (N_3825,N_3678,N_3642);
xnor U3826 (N_3826,N_3661,N_3686);
xnor U3827 (N_3827,N_3756,N_3621);
xnor U3828 (N_3828,N_3792,N_3660);
or U3829 (N_3829,N_3656,N_3668);
or U3830 (N_3830,N_3780,N_3723);
or U3831 (N_3831,N_3693,N_3672);
nor U3832 (N_3832,N_3775,N_3779);
and U3833 (N_3833,N_3606,N_3611);
or U3834 (N_3834,N_3741,N_3703);
and U3835 (N_3835,N_3742,N_3794);
nand U3836 (N_3836,N_3720,N_3689);
and U3837 (N_3837,N_3608,N_3743);
nand U3838 (N_3838,N_3664,N_3655);
nand U3839 (N_3839,N_3744,N_3766);
nand U3840 (N_3840,N_3691,N_3711);
xor U3841 (N_3841,N_3715,N_3784);
xor U3842 (N_3842,N_3768,N_3716);
or U3843 (N_3843,N_3776,N_3773);
nor U3844 (N_3844,N_3778,N_3709);
nand U3845 (N_3845,N_3697,N_3623);
and U3846 (N_3846,N_3707,N_3631);
or U3847 (N_3847,N_3729,N_3677);
xor U3848 (N_3848,N_3682,N_3791);
xnor U3849 (N_3849,N_3734,N_3605);
and U3850 (N_3850,N_3619,N_3788);
xor U3851 (N_3851,N_3650,N_3618);
nor U3852 (N_3852,N_3670,N_3798);
and U3853 (N_3853,N_3722,N_3745);
xor U3854 (N_3854,N_3603,N_3740);
nand U3855 (N_3855,N_3644,N_3713);
nor U3856 (N_3856,N_3673,N_3671);
nor U3857 (N_3857,N_3787,N_3799);
xnor U3858 (N_3858,N_3600,N_3705);
nor U3859 (N_3859,N_3694,N_3736);
or U3860 (N_3860,N_3681,N_3752);
nand U3861 (N_3861,N_3636,N_3687);
or U3862 (N_3862,N_3638,N_3725);
nand U3863 (N_3863,N_3633,N_3626);
nor U3864 (N_3864,N_3710,N_3700);
nor U3865 (N_3865,N_3790,N_3781);
and U3866 (N_3866,N_3634,N_3637);
nand U3867 (N_3867,N_3753,N_3774);
or U3868 (N_3868,N_3667,N_3726);
xor U3869 (N_3869,N_3602,N_3783);
nand U3870 (N_3870,N_3706,N_3640);
nor U3871 (N_3871,N_3628,N_3712);
or U3872 (N_3872,N_3632,N_3719);
nand U3873 (N_3873,N_3748,N_3610);
nor U3874 (N_3874,N_3645,N_3657);
nand U3875 (N_3875,N_3666,N_3679);
and U3876 (N_3876,N_3731,N_3695);
xor U3877 (N_3877,N_3688,N_3614);
nand U3878 (N_3878,N_3708,N_3625);
nor U3879 (N_3879,N_3733,N_3772);
xor U3880 (N_3880,N_3786,N_3704);
or U3881 (N_3881,N_3615,N_3629);
and U3882 (N_3882,N_3609,N_3684);
and U3883 (N_3883,N_3648,N_3612);
nand U3884 (N_3884,N_3757,N_3659);
nand U3885 (N_3885,N_3627,N_3761);
or U3886 (N_3886,N_3613,N_3730);
xor U3887 (N_3887,N_3777,N_3782);
xor U3888 (N_3888,N_3692,N_3647);
nor U3889 (N_3889,N_3662,N_3643);
and U3890 (N_3890,N_3724,N_3622);
xor U3891 (N_3891,N_3765,N_3699);
or U3892 (N_3892,N_3630,N_3728);
or U3893 (N_3893,N_3755,N_3649);
nand U3894 (N_3894,N_3617,N_3746);
nand U3895 (N_3895,N_3701,N_3754);
nand U3896 (N_3896,N_3607,N_3718);
nand U3897 (N_3897,N_3747,N_3760);
or U3898 (N_3898,N_3770,N_3759);
xnor U3899 (N_3899,N_3604,N_3675);
or U3900 (N_3900,N_3647,N_3663);
xnor U3901 (N_3901,N_3797,N_3646);
and U3902 (N_3902,N_3622,N_3773);
nand U3903 (N_3903,N_3691,N_3608);
nand U3904 (N_3904,N_3753,N_3776);
nand U3905 (N_3905,N_3715,N_3749);
xor U3906 (N_3906,N_3675,N_3784);
or U3907 (N_3907,N_3770,N_3620);
xor U3908 (N_3908,N_3634,N_3620);
nand U3909 (N_3909,N_3693,N_3684);
nor U3910 (N_3910,N_3693,N_3654);
and U3911 (N_3911,N_3771,N_3638);
nor U3912 (N_3912,N_3715,N_3772);
or U3913 (N_3913,N_3630,N_3724);
nand U3914 (N_3914,N_3691,N_3754);
or U3915 (N_3915,N_3727,N_3722);
xnor U3916 (N_3916,N_3672,N_3753);
nor U3917 (N_3917,N_3642,N_3768);
nand U3918 (N_3918,N_3715,N_3798);
nand U3919 (N_3919,N_3740,N_3772);
nand U3920 (N_3920,N_3612,N_3643);
nand U3921 (N_3921,N_3628,N_3661);
nand U3922 (N_3922,N_3670,N_3751);
and U3923 (N_3923,N_3669,N_3781);
nand U3924 (N_3924,N_3725,N_3796);
xor U3925 (N_3925,N_3755,N_3660);
xor U3926 (N_3926,N_3716,N_3772);
or U3927 (N_3927,N_3644,N_3693);
or U3928 (N_3928,N_3641,N_3672);
xnor U3929 (N_3929,N_3781,N_3663);
and U3930 (N_3930,N_3770,N_3677);
and U3931 (N_3931,N_3783,N_3738);
and U3932 (N_3932,N_3605,N_3675);
and U3933 (N_3933,N_3672,N_3613);
xor U3934 (N_3934,N_3713,N_3646);
and U3935 (N_3935,N_3660,N_3628);
xnor U3936 (N_3936,N_3641,N_3770);
or U3937 (N_3937,N_3721,N_3792);
and U3938 (N_3938,N_3742,N_3639);
xor U3939 (N_3939,N_3665,N_3617);
or U3940 (N_3940,N_3792,N_3640);
xor U3941 (N_3941,N_3719,N_3601);
nand U3942 (N_3942,N_3769,N_3629);
and U3943 (N_3943,N_3634,N_3677);
nand U3944 (N_3944,N_3661,N_3609);
xor U3945 (N_3945,N_3620,N_3649);
and U3946 (N_3946,N_3623,N_3681);
nand U3947 (N_3947,N_3660,N_3790);
or U3948 (N_3948,N_3776,N_3635);
or U3949 (N_3949,N_3642,N_3721);
and U3950 (N_3950,N_3704,N_3766);
xnor U3951 (N_3951,N_3646,N_3694);
xor U3952 (N_3952,N_3669,N_3727);
or U3953 (N_3953,N_3603,N_3689);
or U3954 (N_3954,N_3626,N_3782);
nand U3955 (N_3955,N_3762,N_3766);
or U3956 (N_3956,N_3738,N_3672);
nand U3957 (N_3957,N_3774,N_3766);
and U3958 (N_3958,N_3694,N_3649);
xnor U3959 (N_3959,N_3794,N_3685);
and U3960 (N_3960,N_3755,N_3736);
xor U3961 (N_3961,N_3694,N_3659);
nand U3962 (N_3962,N_3663,N_3639);
nand U3963 (N_3963,N_3748,N_3756);
or U3964 (N_3964,N_3630,N_3611);
xnor U3965 (N_3965,N_3793,N_3669);
xor U3966 (N_3966,N_3705,N_3752);
or U3967 (N_3967,N_3783,N_3767);
nor U3968 (N_3968,N_3793,N_3639);
nor U3969 (N_3969,N_3795,N_3643);
nand U3970 (N_3970,N_3723,N_3607);
and U3971 (N_3971,N_3664,N_3630);
nor U3972 (N_3972,N_3643,N_3679);
nor U3973 (N_3973,N_3660,N_3607);
or U3974 (N_3974,N_3650,N_3745);
xor U3975 (N_3975,N_3625,N_3633);
nand U3976 (N_3976,N_3755,N_3776);
nor U3977 (N_3977,N_3798,N_3643);
xnor U3978 (N_3978,N_3624,N_3781);
nand U3979 (N_3979,N_3630,N_3613);
xor U3980 (N_3980,N_3711,N_3750);
nor U3981 (N_3981,N_3655,N_3616);
or U3982 (N_3982,N_3733,N_3693);
or U3983 (N_3983,N_3661,N_3703);
or U3984 (N_3984,N_3610,N_3631);
xnor U3985 (N_3985,N_3790,N_3761);
or U3986 (N_3986,N_3713,N_3679);
and U3987 (N_3987,N_3633,N_3756);
and U3988 (N_3988,N_3620,N_3752);
nor U3989 (N_3989,N_3680,N_3776);
or U3990 (N_3990,N_3775,N_3723);
nor U3991 (N_3991,N_3661,N_3689);
xor U3992 (N_3992,N_3648,N_3611);
and U3993 (N_3993,N_3796,N_3747);
nand U3994 (N_3994,N_3788,N_3610);
xnor U3995 (N_3995,N_3733,N_3703);
nand U3996 (N_3996,N_3734,N_3686);
and U3997 (N_3997,N_3747,N_3622);
or U3998 (N_3998,N_3762,N_3652);
xnor U3999 (N_3999,N_3790,N_3626);
nor U4000 (N_4000,N_3843,N_3882);
nor U4001 (N_4001,N_3866,N_3839);
nand U4002 (N_4002,N_3811,N_3926);
nor U4003 (N_4003,N_3928,N_3841);
xnor U4004 (N_4004,N_3842,N_3845);
and U4005 (N_4005,N_3984,N_3911);
xor U4006 (N_4006,N_3986,N_3831);
or U4007 (N_4007,N_3904,N_3947);
and U4008 (N_4008,N_3899,N_3962);
xnor U4009 (N_4009,N_3992,N_3980);
nor U4010 (N_4010,N_3914,N_3906);
xnor U4011 (N_4011,N_3963,N_3876);
nor U4012 (N_4012,N_3924,N_3971);
nand U4013 (N_4013,N_3837,N_3864);
and U4014 (N_4014,N_3959,N_3951);
and U4015 (N_4015,N_3927,N_3868);
and U4016 (N_4016,N_3826,N_3820);
and U4017 (N_4017,N_3885,N_3872);
nand U4018 (N_4018,N_3808,N_3832);
and U4019 (N_4019,N_3920,N_3828);
or U4020 (N_4020,N_3853,N_3895);
nand U4021 (N_4021,N_3821,N_3819);
nor U4022 (N_4022,N_3897,N_3929);
nand U4023 (N_4023,N_3827,N_3877);
nand U4024 (N_4024,N_3881,N_3810);
nor U4025 (N_4025,N_3848,N_3887);
and U4026 (N_4026,N_3941,N_3874);
nand U4027 (N_4027,N_3950,N_3917);
or U4028 (N_4028,N_3939,N_3835);
nand U4029 (N_4029,N_3990,N_3993);
xnor U4030 (N_4030,N_3847,N_3910);
and U4031 (N_4031,N_3970,N_3954);
and U4032 (N_4032,N_3890,N_3800);
or U4033 (N_4033,N_3932,N_3921);
or U4034 (N_4034,N_3915,N_3907);
nand U4035 (N_4035,N_3936,N_3849);
nor U4036 (N_4036,N_3940,N_3858);
nand U4037 (N_4037,N_3974,N_3884);
and U4038 (N_4038,N_3838,N_3972);
xor U4039 (N_4039,N_3802,N_3893);
nor U4040 (N_4040,N_3998,N_3809);
xnor U4041 (N_4041,N_3969,N_3931);
nor U4042 (N_4042,N_3806,N_3807);
nand U4043 (N_4043,N_3916,N_3844);
nor U4044 (N_4044,N_3854,N_3836);
and U4045 (N_4045,N_3812,N_3825);
or U4046 (N_4046,N_3840,N_3818);
nor U4047 (N_4047,N_3933,N_3894);
nand U4048 (N_4048,N_3883,N_3803);
nor U4049 (N_4049,N_3829,N_3948);
xnor U4050 (N_4050,N_3973,N_3822);
nor U4051 (N_4051,N_3923,N_3982);
or U4052 (N_4052,N_3801,N_3979);
xor U4053 (N_4053,N_3909,N_3988);
or U4054 (N_4054,N_3913,N_3863);
and U4055 (N_4055,N_3865,N_3912);
or U4056 (N_4056,N_3851,N_3997);
nand U4057 (N_4057,N_3871,N_3815);
nor U4058 (N_4058,N_3945,N_3952);
or U4059 (N_4059,N_3955,N_3857);
and U4060 (N_4060,N_3855,N_3975);
and U4061 (N_4061,N_3892,N_3976);
or U4062 (N_4062,N_3824,N_3956);
nor U4063 (N_4063,N_3953,N_3942);
and U4064 (N_4064,N_3891,N_3859);
and U4065 (N_4065,N_3861,N_3987);
nor U4066 (N_4066,N_3850,N_3995);
or U4067 (N_4067,N_3900,N_3934);
nor U4068 (N_4068,N_3817,N_3878);
xnor U4069 (N_4069,N_3994,N_3977);
xor U4070 (N_4070,N_3846,N_3814);
and U4071 (N_4071,N_3949,N_3922);
nand U4072 (N_4072,N_3961,N_3898);
nand U4073 (N_4073,N_3985,N_3925);
and U4074 (N_4074,N_3879,N_3880);
and U4075 (N_4075,N_3908,N_3935);
nand U4076 (N_4076,N_3957,N_3938);
xnor U4077 (N_4077,N_3862,N_3834);
or U4078 (N_4078,N_3902,N_3918);
nor U4079 (N_4079,N_3965,N_3968);
nor U4080 (N_4080,N_3989,N_3816);
xnor U4081 (N_4081,N_3852,N_3813);
or U4082 (N_4082,N_3856,N_3991);
or U4083 (N_4083,N_3943,N_3805);
nand U4084 (N_4084,N_3919,N_3804);
or U4085 (N_4085,N_3960,N_3981);
nor U4086 (N_4086,N_3946,N_3888);
xnor U4087 (N_4087,N_3873,N_3983);
and U4088 (N_4088,N_3930,N_3966);
and U4089 (N_4089,N_3958,N_3967);
or U4090 (N_4090,N_3944,N_3833);
and U4091 (N_4091,N_3867,N_3870);
xnor U4092 (N_4092,N_3889,N_3937);
and U4093 (N_4093,N_3999,N_3964);
or U4094 (N_4094,N_3905,N_3823);
nor U4095 (N_4095,N_3886,N_3860);
nand U4096 (N_4096,N_3903,N_3996);
or U4097 (N_4097,N_3869,N_3978);
nand U4098 (N_4098,N_3896,N_3901);
or U4099 (N_4099,N_3830,N_3875);
nor U4100 (N_4100,N_3861,N_3828);
or U4101 (N_4101,N_3951,N_3974);
nand U4102 (N_4102,N_3891,N_3896);
and U4103 (N_4103,N_3885,N_3829);
nand U4104 (N_4104,N_3903,N_3824);
nor U4105 (N_4105,N_3814,N_3839);
and U4106 (N_4106,N_3996,N_3808);
nand U4107 (N_4107,N_3984,N_3912);
nand U4108 (N_4108,N_3968,N_3813);
or U4109 (N_4109,N_3916,N_3854);
or U4110 (N_4110,N_3962,N_3888);
nand U4111 (N_4111,N_3888,N_3935);
xor U4112 (N_4112,N_3995,N_3808);
xor U4113 (N_4113,N_3878,N_3919);
or U4114 (N_4114,N_3921,N_3834);
or U4115 (N_4115,N_3908,N_3804);
and U4116 (N_4116,N_3969,N_3983);
or U4117 (N_4117,N_3950,N_3844);
and U4118 (N_4118,N_3917,N_3814);
nor U4119 (N_4119,N_3846,N_3861);
or U4120 (N_4120,N_3943,N_3831);
nor U4121 (N_4121,N_3814,N_3982);
or U4122 (N_4122,N_3804,N_3810);
nor U4123 (N_4123,N_3960,N_3881);
nand U4124 (N_4124,N_3816,N_3937);
or U4125 (N_4125,N_3806,N_3937);
xor U4126 (N_4126,N_3925,N_3898);
or U4127 (N_4127,N_3950,N_3998);
and U4128 (N_4128,N_3944,N_3904);
and U4129 (N_4129,N_3897,N_3834);
nor U4130 (N_4130,N_3830,N_3855);
nand U4131 (N_4131,N_3930,N_3988);
or U4132 (N_4132,N_3992,N_3904);
and U4133 (N_4133,N_3990,N_3919);
or U4134 (N_4134,N_3883,N_3818);
nor U4135 (N_4135,N_3912,N_3928);
or U4136 (N_4136,N_3934,N_3939);
nor U4137 (N_4137,N_3859,N_3801);
nand U4138 (N_4138,N_3928,N_3842);
nand U4139 (N_4139,N_3833,N_3846);
nor U4140 (N_4140,N_3907,N_3985);
and U4141 (N_4141,N_3821,N_3933);
xnor U4142 (N_4142,N_3888,N_3814);
and U4143 (N_4143,N_3934,N_3800);
or U4144 (N_4144,N_3938,N_3839);
and U4145 (N_4145,N_3833,N_3815);
nor U4146 (N_4146,N_3930,N_3816);
or U4147 (N_4147,N_3832,N_3800);
and U4148 (N_4148,N_3964,N_3866);
and U4149 (N_4149,N_3983,N_3945);
nand U4150 (N_4150,N_3931,N_3971);
nor U4151 (N_4151,N_3863,N_3921);
nand U4152 (N_4152,N_3867,N_3970);
xor U4153 (N_4153,N_3868,N_3978);
or U4154 (N_4154,N_3929,N_3981);
or U4155 (N_4155,N_3895,N_3995);
and U4156 (N_4156,N_3826,N_3866);
nand U4157 (N_4157,N_3878,N_3883);
or U4158 (N_4158,N_3873,N_3824);
nor U4159 (N_4159,N_3927,N_3941);
nor U4160 (N_4160,N_3981,N_3940);
or U4161 (N_4161,N_3809,N_3824);
nand U4162 (N_4162,N_3997,N_3979);
nand U4163 (N_4163,N_3828,N_3919);
and U4164 (N_4164,N_3952,N_3877);
nand U4165 (N_4165,N_3845,N_3875);
xnor U4166 (N_4166,N_3975,N_3962);
and U4167 (N_4167,N_3972,N_3921);
or U4168 (N_4168,N_3973,N_3988);
and U4169 (N_4169,N_3973,N_3904);
or U4170 (N_4170,N_3893,N_3811);
xnor U4171 (N_4171,N_3825,N_3826);
nor U4172 (N_4172,N_3896,N_3867);
and U4173 (N_4173,N_3979,N_3904);
xor U4174 (N_4174,N_3866,N_3852);
xor U4175 (N_4175,N_3991,N_3889);
nor U4176 (N_4176,N_3917,N_3894);
nand U4177 (N_4177,N_3915,N_3964);
and U4178 (N_4178,N_3968,N_3850);
nand U4179 (N_4179,N_3859,N_3836);
nor U4180 (N_4180,N_3801,N_3808);
xor U4181 (N_4181,N_3824,N_3864);
and U4182 (N_4182,N_3976,N_3937);
xnor U4183 (N_4183,N_3866,N_3965);
or U4184 (N_4184,N_3975,N_3856);
nor U4185 (N_4185,N_3859,N_3855);
xnor U4186 (N_4186,N_3985,N_3992);
xor U4187 (N_4187,N_3925,N_3927);
nor U4188 (N_4188,N_3800,N_3925);
nor U4189 (N_4189,N_3931,N_3936);
nand U4190 (N_4190,N_3911,N_3874);
or U4191 (N_4191,N_3933,N_3955);
xor U4192 (N_4192,N_3998,N_3870);
nand U4193 (N_4193,N_3892,N_3838);
xor U4194 (N_4194,N_3951,N_3808);
and U4195 (N_4195,N_3985,N_3845);
nand U4196 (N_4196,N_3862,N_3803);
nand U4197 (N_4197,N_3826,N_3930);
nor U4198 (N_4198,N_3892,N_3971);
xor U4199 (N_4199,N_3943,N_3811);
and U4200 (N_4200,N_4181,N_4016);
xor U4201 (N_4201,N_4076,N_4073);
nor U4202 (N_4202,N_4055,N_4144);
nand U4203 (N_4203,N_4135,N_4088);
or U4204 (N_4204,N_4023,N_4183);
nor U4205 (N_4205,N_4000,N_4081);
or U4206 (N_4206,N_4011,N_4138);
xor U4207 (N_4207,N_4130,N_4166);
xnor U4208 (N_4208,N_4025,N_4077);
nor U4209 (N_4209,N_4137,N_4096);
nor U4210 (N_4210,N_4048,N_4087);
nor U4211 (N_4211,N_4017,N_4172);
xor U4212 (N_4212,N_4101,N_4156);
nor U4213 (N_4213,N_4067,N_4019);
nand U4214 (N_4214,N_4071,N_4116);
xnor U4215 (N_4215,N_4054,N_4127);
xnor U4216 (N_4216,N_4038,N_4113);
xor U4217 (N_4217,N_4089,N_4056);
or U4218 (N_4218,N_4028,N_4098);
or U4219 (N_4219,N_4005,N_4074);
nor U4220 (N_4220,N_4112,N_4122);
xor U4221 (N_4221,N_4008,N_4029);
and U4222 (N_4222,N_4150,N_4182);
xor U4223 (N_4223,N_4118,N_4104);
or U4224 (N_4224,N_4111,N_4084);
and U4225 (N_4225,N_4036,N_4190);
nand U4226 (N_4226,N_4102,N_4179);
or U4227 (N_4227,N_4194,N_4106);
xor U4228 (N_4228,N_4198,N_4175);
or U4229 (N_4229,N_4153,N_4132);
nand U4230 (N_4230,N_4032,N_4047);
nand U4231 (N_4231,N_4070,N_4050);
or U4232 (N_4232,N_4053,N_4066);
or U4233 (N_4233,N_4045,N_4063);
or U4234 (N_4234,N_4131,N_4035);
and U4235 (N_4235,N_4020,N_4100);
nor U4236 (N_4236,N_4110,N_4191);
or U4237 (N_4237,N_4124,N_4155);
and U4238 (N_4238,N_4037,N_4001);
xnor U4239 (N_4239,N_4146,N_4061);
and U4240 (N_4240,N_4064,N_4007);
and U4241 (N_4241,N_4014,N_4117);
xnor U4242 (N_4242,N_4143,N_4006);
nor U4243 (N_4243,N_4126,N_4092);
xnor U4244 (N_4244,N_4044,N_4069);
nand U4245 (N_4245,N_4107,N_4180);
xnor U4246 (N_4246,N_4168,N_4164);
nor U4247 (N_4247,N_4105,N_4159);
nor U4248 (N_4248,N_4018,N_4128);
nor U4249 (N_4249,N_4068,N_4094);
xnor U4250 (N_4250,N_4060,N_4040);
and U4251 (N_4251,N_4157,N_4171);
xor U4252 (N_4252,N_4141,N_4115);
nand U4253 (N_4253,N_4174,N_4186);
and U4254 (N_4254,N_4031,N_4108);
nor U4255 (N_4255,N_4123,N_4004);
nor U4256 (N_4256,N_4009,N_4042);
or U4257 (N_4257,N_4078,N_4161);
nor U4258 (N_4258,N_4039,N_4046);
or U4259 (N_4259,N_4072,N_4187);
or U4260 (N_4260,N_4043,N_4059);
and U4261 (N_4261,N_4151,N_4149);
xnor U4262 (N_4262,N_4010,N_4079);
nor U4263 (N_4263,N_4169,N_4121);
nand U4264 (N_4264,N_4003,N_4120);
xnor U4265 (N_4265,N_4027,N_4030);
or U4266 (N_4266,N_4086,N_4196);
nand U4267 (N_4267,N_4133,N_4154);
nand U4268 (N_4268,N_4125,N_4002);
and U4269 (N_4269,N_4170,N_4022);
xor U4270 (N_4270,N_4049,N_4142);
nand U4271 (N_4271,N_4114,N_4099);
and U4272 (N_4272,N_4093,N_4197);
and U4273 (N_4273,N_4041,N_4195);
nor U4274 (N_4274,N_4015,N_4162);
or U4275 (N_4275,N_4177,N_4024);
nand U4276 (N_4276,N_4134,N_4058);
and U4277 (N_4277,N_4012,N_4192);
or U4278 (N_4278,N_4145,N_4026);
and U4279 (N_4279,N_4158,N_4057);
nor U4280 (N_4280,N_4152,N_4021);
xnor U4281 (N_4281,N_4095,N_4140);
nand U4282 (N_4282,N_4052,N_4051);
and U4283 (N_4283,N_4083,N_4062);
or U4284 (N_4284,N_4184,N_4080);
or U4285 (N_4285,N_4167,N_4189);
or U4286 (N_4286,N_4082,N_4091);
xor U4287 (N_4287,N_4033,N_4163);
and U4288 (N_4288,N_4147,N_4199);
and U4289 (N_4289,N_4136,N_4129);
nand U4290 (N_4290,N_4075,N_4148);
or U4291 (N_4291,N_4065,N_4013);
xor U4292 (N_4292,N_4165,N_4097);
nor U4293 (N_4293,N_4193,N_4085);
nand U4294 (N_4294,N_4139,N_4119);
or U4295 (N_4295,N_4103,N_4173);
or U4296 (N_4296,N_4178,N_4109);
and U4297 (N_4297,N_4188,N_4160);
or U4298 (N_4298,N_4090,N_4185);
or U4299 (N_4299,N_4034,N_4176);
xnor U4300 (N_4300,N_4085,N_4152);
nor U4301 (N_4301,N_4062,N_4045);
nand U4302 (N_4302,N_4186,N_4191);
nor U4303 (N_4303,N_4073,N_4176);
and U4304 (N_4304,N_4070,N_4043);
nor U4305 (N_4305,N_4109,N_4099);
and U4306 (N_4306,N_4018,N_4155);
nor U4307 (N_4307,N_4040,N_4113);
nand U4308 (N_4308,N_4159,N_4195);
nand U4309 (N_4309,N_4174,N_4142);
xor U4310 (N_4310,N_4049,N_4077);
nand U4311 (N_4311,N_4018,N_4161);
and U4312 (N_4312,N_4126,N_4107);
nor U4313 (N_4313,N_4086,N_4149);
xor U4314 (N_4314,N_4062,N_4058);
nand U4315 (N_4315,N_4175,N_4153);
nor U4316 (N_4316,N_4164,N_4062);
or U4317 (N_4317,N_4184,N_4109);
nor U4318 (N_4318,N_4066,N_4187);
and U4319 (N_4319,N_4094,N_4035);
and U4320 (N_4320,N_4060,N_4017);
xnor U4321 (N_4321,N_4038,N_4055);
or U4322 (N_4322,N_4095,N_4102);
or U4323 (N_4323,N_4059,N_4183);
nor U4324 (N_4324,N_4071,N_4166);
or U4325 (N_4325,N_4038,N_4137);
nor U4326 (N_4326,N_4140,N_4037);
xor U4327 (N_4327,N_4148,N_4000);
nand U4328 (N_4328,N_4015,N_4000);
and U4329 (N_4329,N_4027,N_4153);
xnor U4330 (N_4330,N_4025,N_4016);
or U4331 (N_4331,N_4025,N_4068);
nand U4332 (N_4332,N_4108,N_4181);
xnor U4333 (N_4333,N_4054,N_4106);
and U4334 (N_4334,N_4054,N_4158);
nand U4335 (N_4335,N_4143,N_4092);
and U4336 (N_4336,N_4109,N_4176);
xnor U4337 (N_4337,N_4001,N_4052);
xor U4338 (N_4338,N_4167,N_4099);
or U4339 (N_4339,N_4114,N_4116);
and U4340 (N_4340,N_4093,N_4031);
and U4341 (N_4341,N_4141,N_4090);
or U4342 (N_4342,N_4176,N_4030);
nor U4343 (N_4343,N_4159,N_4139);
nor U4344 (N_4344,N_4086,N_4000);
or U4345 (N_4345,N_4026,N_4116);
or U4346 (N_4346,N_4168,N_4004);
nand U4347 (N_4347,N_4014,N_4087);
xnor U4348 (N_4348,N_4101,N_4060);
nand U4349 (N_4349,N_4193,N_4144);
or U4350 (N_4350,N_4108,N_4073);
and U4351 (N_4351,N_4076,N_4181);
xor U4352 (N_4352,N_4192,N_4073);
nor U4353 (N_4353,N_4055,N_4002);
and U4354 (N_4354,N_4148,N_4185);
and U4355 (N_4355,N_4164,N_4153);
nand U4356 (N_4356,N_4176,N_4011);
nand U4357 (N_4357,N_4112,N_4171);
xor U4358 (N_4358,N_4091,N_4041);
nor U4359 (N_4359,N_4096,N_4134);
and U4360 (N_4360,N_4014,N_4133);
or U4361 (N_4361,N_4109,N_4037);
nor U4362 (N_4362,N_4107,N_4127);
nor U4363 (N_4363,N_4114,N_4028);
and U4364 (N_4364,N_4126,N_4157);
nor U4365 (N_4365,N_4050,N_4090);
nor U4366 (N_4366,N_4150,N_4076);
nand U4367 (N_4367,N_4067,N_4160);
or U4368 (N_4368,N_4116,N_4146);
nor U4369 (N_4369,N_4116,N_4143);
xnor U4370 (N_4370,N_4154,N_4193);
nand U4371 (N_4371,N_4023,N_4196);
xnor U4372 (N_4372,N_4185,N_4140);
nand U4373 (N_4373,N_4095,N_4081);
xnor U4374 (N_4374,N_4157,N_4035);
xor U4375 (N_4375,N_4150,N_4067);
or U4376 (N_4376,N_4077,N_4017);
nand U4377 (N_4377,N_4021,N_4029);
nor U4378 (N_4378,N_4013,N_4026);
or U4379 (N_4379,N_4018,N_4045);
xor U4380 (N_4380,N_4087,N_4065);
xnor U4381 (N_4381,N_4065,N_4049);
or U4382 (N_4382,N_4031,N_4174);
or U4383 (N_4383,N_4120,N_4088);
nor U4384 (N_4384,N_4193,N_4062);
nand U4385 (N_4385,N_4182,N_4059);
and U4386 (N_4386,N_4108,N_4141);
nand U4387 (N_4387,N_4081,N_4045);
and U4388 (N_4388,N_4194,N_4040);
or U4389 (N_4389,N_4175,N_4174);
nor U4390 (N_4390,N_4147,N_4143);
or U4391 (N_4391,N_4099,N_4165);
and U4392 (N_4392,N_4015,N_4139);
nor U4393 (N_4393,N_4170,N_4106);
xnor U4394 (N_4394,N_4038,N_4194);
and U4395 (N_4395,N_4085,N_4045);
nor U4396 (N_4396,N_4189,N_4061);
nand U4397 (N_4397,N_4086,N_4148);
and U4398 (N_4398,N_4110,N_4092);
nor U4399 (N_4399,N_4120,N_4018);
xor U4400 (N_4400,N_4246,N_4267);
nor U4401 (N_4401,N_4222,N_4233);
xor U4402 (N_4402,N_4227,N_4206);
and U4403 (N_4403,N_4303,N_4279);
nor U4404 (N_4404,N_4358,N_4200);
nor U4405 (N_4405,N_4263,N_4272);
nor U4406 (N_4406,N_4215,N_4384);
nand U4407 (N_4407,N_4205,N_4350);
nor U4408 (N_4408,N_4321,N_4307);
xor U4409 (N_4409,N_4361,N_4310);
or U4410 (N_4410,N_4323,N_4380);
nand U4411 (N_4411,N_4290,N_4301);
and U4412 (N_4412,N_4232,N_4309);
or U4413 (N_4413,N_4241,N_4395);
xnor U4414 (N_4414,N_4218,N_4292);
nor U4415 (N_4415,N_4208,N_4293);
nor U4416 (N_4416,N_4304,N_4203);
and U4417 (N_4417,N_4357,N_4393);
xor U4418 (N_4418,N_4397,N_4236);
xor U4419 (N_4419,N_4362,N_4229);
xor U4420 (N_4420,N_4398,N_4312);
and U4421 (N_4421,N_4258,N_4287);
nor U4422 (N_4422,N_4237,N_4231);
nand U4423 (N_4423,N_4319,N_4225);
or U4424 (N_4424,N_4392,N_4250);
nor U4425 (N_4425,N_4217,N_4212);
or U4426 (N_4426,N_4219,N_4318);
xnor U4427 (N_4427,N_4360,N_4344);
nor U4428 (N_4428,N_4269,N_4281);
nor U4429 (N_4429,N_4276,N_4235);
and U4430 (N_4430,N_4371,N_4343);
or U4431 (N_4431,N_4342,N_4253);
and U4432 (N_4432,N_4265,N_4373);
and U4433 (N_4433,N_4228,N_4314);
nor U4434 (N_4434,N_4221,N_4389);
nand U4435 (N_4435,N_4369,N_4341);
xor U4436 (N_4436,N_4282,N_4224);
nand U4437 (N_4437,N_4214,N_4266);
nor U4438 (N_4438,N_4268,N_4377);
nor U4439 (N_4439,N_4340,N_4247);
and U4440 (N_4440,N_4299,N_4347);
nand U4441 (N_4441,N_4336,N_4252);
nand U4442 (N_4442,N_4313,N_4326);
or U4443 (N_4443,N_4370,N_4349);
or U4444 (N_4444,N_4353,N_4201);
and U4445 (N_4445,N_4328,N_4375);
and U4446 (N_4446,N_4382,N_4285);
nor U4447 (N_4447,N_4283,N_4274);
xor U4448 (N_4448,N_4262,N_4345);
or U4449 (N_4449,N_4348,N_4331);
nand U4450 (N_4450,N_4234,N_4351);
xnor U4451 (N_4451,N_4352,N_4248);
nor U4452 (N_4452,N_4338,N_4325);
and U4453 (N_4453,N_4363,N_4335);
or U4454 (N_4454,N_4239,N_4278);
nor U4455 (N_4455,N_4381,N_4238);
nor U4456 (N_4456,N_4305,N_4365);
and U4457 (N_4457,N_4264,N_4273);
nand U4458 (N_4458,N_4211,N_4220);
nand U4459 (N_4459,N_4324,N_4315);
nand U4460 (N_4460,N_4296,N_4245);
nand U4461 (N_4461,N_4280,N_4391);
or U4462 (N_4462,N_4223,N_4275);
nor U4463 (N_4463,N_4254,N_4387);
nand U4464 (N_4464,N_4368,N_4256);
or U4465 (N_4465,N_4306,N_4284);
xor U4466 (N_4466,N_4202,N_4322);
and U4467 (N_4467,N_4346,N_4337);
or U4468 (N_4468,N_4288,N_4367);
nand U4469 (N_4469,N_4251,N_4354);
xnor U4470 (N_4470,N_4244,N_4210);
and U4471 (N_4471,N_4317,N_4230);
or U4472 (N_4472,N_4249,N_4355);
or U4473 (N_4473,N_4374,N_4207);
xnor U4474 (N_4474,N_4300,N_4383);
and U4475 (N_4475,N_4386,N_4240);
nor U4476 (N_4476,N_4286,N_4366);
xnor U4477 (N_4477,N_4294,N_4379);
xor U4478 (N_4478,N_4308,N_4334);
nand U4479 (N_4479,N_4255,N_4356);
nand U4480 (N_4480,N_4242,N_4297);
nand U4481 (N_4481,N_4243,N_4332);
or U4482 (N_4482,N_4390,N_4364);
and U4483 (N_4483,N_4376,N_4320);
or U4484 (N_4484,N_4260,N_4333);
nor U4485 (N_4485,N_4257,N_4311);
xnor U4486 (N_4486,N_4372,N_4359);
or U4487 (N_4487,N_4271,N_4291);
and U4488 (N_4488,N_4399,N_4204);
xor U4489 (N_4489,N_4226,N_4378);
and U4490 (N_4490,N_4316,N_4209);
nor U4491 (N_4491,N_4327,N_4394);
or U4492 (N_4492,N_4385,N_4213);
nand U4493 (N_4493,N_4330,N_4277);
nor U4494 (N_4494,N_4329,N_4388);
nand U4495 (N_4495,N_4396,N_4259);
xnor U4496 (N_4496,N_4339,N_4302);
nand U4497 (N_4497,N_4216,N_4270);
xor U4498 (N_4498,N_4261,N_4289);
and U4499 (N_4499,N_4298,N_4295);
or U4500 (N_4500,N_4370,N_4236);
xor U4501 (N_4501,N_4216,N_4376);
xor U4502 (N_4502,N_4207,N_4216);
nand U4503 (N_4503,N_4304,N_4221);
and U4504 (N_4504,N_4283,N_4213);
nand U4505 (N_4505,N_4363,N_4208);
nor U4506 (N_4506,N_4346,N_4355);
and U4507 (N_4507,N_4273,N_4231);
or U4508 (N_4508,N_4234,N_4286);
nand U4509 (N_4509,N_4222,N_4253);
xnor U4510 (N_4510,N_4361,N_4266);
and U4511 (N_4511,N_4386,N_4376);
or U4512 (N_4512,N_4363,N_4352);
nand U4513 (N_4513,N_4357,N_4362);
and U4514 (N_4514,N_4337,N_4278);
nand U4515 (N_4515,N_4274,N_4387);
xor U4516 (N_4516,N_4357,N_4257);
or U4517 (N_4517,N_4393,N_4352);
nor U4518 (N_4518,N_4314,N_4325);
xor U4519 (N_4519,N_4206,N_4326);
nand U4520 (N_4520,N_4246,N_4373);
or U4521 (N_4521,N_4273,N_4238);
nor U4522 (N_4522,N_4267,N_4321);
nand U4523 (N_4523,N_4317,N_4353);
nor U4524 (N_4524,N_4249,N_4238);
or U4525 (N_4525,N_4287,N_4206);
nand U4526 (N_4526,N_4398,N_4212);
nand U4527 (N_4527,N_4363,N_4399);
or U4528 (N_4528,N_4220,N_4230);
nor U4529 (N_4529,N_4358,N_4311);
nor U4530 (N_4530,N_4248,N_4263);
and U4531 (N_4531,N_4309,N_4337);
or U4532 (N_4532,N_4267,N_4207);
nor U4533 (N_4533,N_4305,N_4388);
or U4534 (N_4534,N_4354,N_4390);
nor U4535 (N_4535,N_4210,N_4381);
and U4536 (N_4536,N_4294,N_4328);
nor U4537 (N_4537,N_4319,N_4238);
and U4538 (N_4538,N_4214,N_4344);
xnor U4539 (N_4539,N_4221,N_4384);
and U4540 (N_4540,N_4392,N_4223);
nor U4541 (N_4541,N_4251,N_4395);
nand U4542 (N_4542,N_4308,N_4271);
xor U4543 (N_4543,N_4242,N_4286);
and U4544 (N_4544,N_4393,N_4362);
nand U4545 (N_4545,N_4245,N_4336);
and U4546 (N_4546,N_4357,N_4269);
or U4547 (N_4547,N_4218,N_4380);
xor U4548 (N_4548,N_4266,N_4257);
nand U4549 (N_4549,N_4297,N_4352);
nand U4550 (N_4550,N_4210,N_4354);
nand U4551 (N_4551,N_4337,N_4355);
nor U4552 (N_4552,N_4372,N_4239);
xnor U4553 (N_4553,N_4211,N_4319);
xnor U4554 (N_4554,N_4270,N_4289);
nor U4555 (N_4555,N_4204,N_4345);
nor U4556 (N_4556,N_4314,N_4290);
or U4557 (N_4557,N_4365,N_4309);
and U4558 (N_4558,N_4279,N_4220);
xor U4559 (N_4559,N_4245,N_4223);
xnor U4560 (N_4560,N_4337,N_4273);
nand U4561 (N_4561,N_4269,N_4237);
or U4562 (N_4562,N_4234,N_4209);
nor U4563 (N_4563,N_4368,N_4255);
xnor U4564 (N_4564,N_4249,N_4344);
and U4565 (N_4565,N_4361,N_4223);
xnor U4566 (N_4566,N_4370,N_4212);
or U4567 (N_4567,N_4207,N_4290);
and U4568 (N_4568,N_4204,N_4254);
xor U4569 (N_4569,N_4214,N_4391);
or U4570 (N_4570,N_4331,N_4295);
or U4571 (N_4571,N_4348,N_4387);
nand U4572 (N_4572,N_4256,N_4316);
or U4573 (N_4573,N_4294,N_4201);
and U4574 (N_4574,N_4256,N_4340);
nor U4575 (N_4575,N_4222,N_4380);
xor U4576 (N_4576,N_4354,N_4201);
nand U4577 (N_4577,N_4263,N_4285);
and U4578 (N_4578,N_4205,N_4259);
or U4579 (N_4579,N_4233,N_4279);
and U4580 (N_4580,N_4226,N_4389);
and U4581 (N_4581,N_4387,N_4201);
xor U4582 (N_4582,N_4311,N_4250);
or U4583 (N_4583,N_4346,N_4307);
xor U4584 (N_4584,N_4346,N_4387);
nor U4585 (N_4585,N_4251,N_4228);
nand U4586 (N_4586,N_4373,N_4370);
nand U4587 (N_4587,N_4383,N_4282);
nor U4588 (N_4588,N_4312,N_4319);
xor U4589 (N_4589,N_4384,N_4278);
and U4590 (N_4590,N_4240,N_4230);
nor U4591 (N_4591,N_4323,N_4369);
xor U4592 (N_4592,N_4368,N_4238);
nand U4593 (N_4593,N_4218,N_4215);
or U4594 (N_4594,N_4302,N_4378);
xnor U4595 (N_4595,N_4323,N_4359);
nand U4596 (N_4596,N_4202,N_4220);
or U4597 (N_4597,N_4246,N_4399);
nor U4598 (N_4598,N_4379,N_4381);
or U4599 (N_4599,N_4306,N_4222);
xor U4600 (N_4600,N_4575,N_4559);
nor U4601 (N_4601,N_4495,N_4568);
xnor U4602 (N_4602,N_4524,N_4457);
nand U4603 (N_4603,N_4408,N_4541);
or U4604 (N_4604,N_4522,N_4525);
or U4605 (N_4605,N_4445,N_4427);
or U4606 (N_4606,N_4499,N_4484);
or U4607 (N_4607,N_4456,N_4583);
or U4608 (N_4608,N_4501,N_4515);
xor U4609 (N_4609,N_4438,N_4562);
or U4610 (N_4610,N_4506,N_4556);
nor U4611 (N_4611,N_4472,N_4433);
or U4612 (N_4612,N_4406,N_4443);
xnor U4613 (N_4613,N_4404,N_4550);
or U4614 (N_4614,N_4436,N_4584);
xnor U4615 (N_4615,N_4448,N_4444);
xor U4616 (N_4616,N_4597,N_4591);
xnor U4617 (N_4617,N_4598,N_4538);
or U4618 (N_4618,N_4567,N_4463);
nor U4619 (N_4619,N_4578,N_4498);
nand U4620 (N_4620,N_4486,N_4534);
or U4621 (N_4621,N_4485,N_4529);
or U4622 (N_4622,N_4442,N_4503);
and U4623 (N_4623,N_4405,N_4439);
nor U4624 (N_4624,N_4470,N_4455);
and U4625 (N_4625,N_4544,N_4533);
xor U4626 (N_4626,N_4458,N_4451);
nor U4627 (N_4627,N_4482,N_4402);
or U4628 (N_4628,N_4518,N_4423);
nand U4629 (N_4629,N_4514,N_4537);
or U4630 (N_4630,N_4409,N_4579);
nor U4631 (N_4631,N_4466,N_4573);
nand U4632 (N_4632,N_4415,N_4547);
and U4633 (N_4633,N_4587,N_4527);
xor U4634 (N_4634,N_4450,N_4526);
nor U4635 (N_4635,N_4545,N_4507);
nor U4636 (N_4636,N_4400,N_4516);
and U4637 (N_4637,N_4464,N_4413);
and U4638 (N_4638,N_4581,N_4407);
nor U4639 (N_4639,N_4582,N_4539);
and U4640 (N_4640,N_4435,N_4555);
nor U4641 (N_4641,N_4403,N_4596);
nand U4642 (N_4642,N_4558,N_4494);
and U4643 (N_4643,N_4546,N_4447);
nand U4644 (N_4644,N_4434,N_4508);
or U4645 (N_4645,N_4401,N_4563);
or U4646 (N_4646,N_4549,N_4461);
nor U4647 (N_4647,N_4577,N_4580);
and U4648 (N_4648,N_4521,N_4512);
and U4649 (N_4649,N_4557,N_4569);
nor U4650 (N_4650,N_4417,N_4560);
and U4651 (N_4651,N_4505,N_4449);
and U4652 (N_4652,N_4475,N_4571);
nor U4653 (N_4653,N_4459,N_4412);
or U4654 (N_4654,N_4523,N_4590);
xor U4655 (N_4655,N_4471,N_4532);
or U4656 (N_4656,N_4429,N_4502);
or U4657 (N_4657,N_4465,N_4418);
or U4658 (N_4658,N_4410,N_4430);
xor U4659 (N_4659,N_4425,N_4421);
nor U4660 (N_4660,N_4460,N_4510);
or U4661 (N_4661,N_4595,N_4586);
nand U4662 (N_4662,N_4420,N_4432);
nand U4663 (N_4663,N_4599,N_4479);
xnor U4664 (N_4664,N_4511,N_4452);
and U4665 (N_4665,N_4565,N_4572);
and U4666 (N_4666,N_4488,N_4419);
and U4667 (N_4667,N_4492,N_4491);
xnor U4668 (N_4668,N_4530,N_4422);
and U4669 (N_4669,N_4589,N_4481);
or U4670 (N_4670,N_4594,N_4536);
nor U4671 (N_4671,N_4519,N_4493);
nor U4672 (N_4672,N_4548,N_4564);
or U4673 (N_4673,N_4416,N_4478);
xor U4674 (N_4674,N_4496,N_4552);
nor U4675 (N_4675,N_4428,N_4480);
nor U4676 (N_4676,N_4476,N_4504);
xor U4677 (N_4677,N_4468,N_4477);
nand U4678 (N_4678,N_4540,N_4411);
nand U4679 (N_4679,N_4553,N_4474);
or U4680 (N_4680,N_4440,N_4469);
and U4681 (N_4681,N_4513,N_4520);
nand U4682 (N_4682,N_4489,N_4500);
xor U4683 (N_4683,N_4588,N_4431);
xnor U4684 (N_4684,N_4509,N_4592);
and U4685 (N_4685,N_4437,N_4531);
or U4686 (N_4686,N_4453,N_4551);
or U4687 (N_4687,N_4554,N_4446);
xnor U4688 (N_4688,N_4542,N_4497);
or U4689 (N_4689,N_4483,N_4576);
or U4690 (N_4690,N_4517,N_4570);
nand U4691 (N_4691,N_4467,N_4593);
nand U4692 (N_4692,N_4441,N_4528);
xor U4693 (N_4693,N_4426,N_4585);
nor U4694 (N_4694,N_4490,N_4487);
and U4695 (N_4695,N_4543,N_4454);
and U4696 (N_4696,N_4414,N_4424);
nand U4697 (N_4697,N_4535,N_4462);
xnor U4698 (N_4698,N_4566,N_4574);
nor U4699 (N_4699,N_4473,N_4561);
nor U4700 (N_4700,N_4464,N_4496);
and U4701 (N_4701,N_4550,N_4484);
nand U4702 (N_4702,N_4407,N_4548);
nor U4703 (N_4703,N_4483,N_4509);
or U4704 (N_4704,N_4563,N_4586);
nand U4705 (N_4705,N_4461,N_4454);
xor U4706 (N_4706,N_4424,N_4493);
and U4707 (N_4707,N_4559,N_4414);
or U4708 (N_4708,N_4596,N_4567);
and U4709 (N_4709,N_4588,N_4593);
xor U4710 (N_4710,N_4455,N_4541);
or U4711 (N_4711,N_4567,N_4545);
or U4712 (N_4712,N_4487,N_4557);
and U4713 (N_4713,N_4456,N_4497);
xor U4714 (N_4714,N_4561,N_4440);
xor U4715 (N_4715,N_4578,N_4565);
xnor U4716 (N_4716,N_4587,N_4515);
or U4717 (N_4717,N_4420,N_4576);
xnor U4718 (N_4718,N_4465,N_4491);
nor U4719 (N_4719,N_4471,N_4524);
or U4720 (N_4720,N_4471,N_4400);
or U4721 (N_4721,N_4404,N_4483);
or U4722 (N_4722,N_4536,N_4502);
or U4723 (N_4723,N_4430,N_4573);
xnor U4724 (N_4724,N_4477,N_4540);
xor U4725 (N_4725,N_4540,N_4512);
nor U4726 (N_4726,N_4421,N_4579);
nand U4727 (N_4727,N_4503,N_4435);
xnor U4728 (N_4728,N_4452,N_4411);
or U4729 (N_4729,N_4490,N_4499);
or U4730 (N_4730,N_4464,N_4429);
nand U4731 (N_4731,N_4428,N_4409);
and U4732 (N_4732,N_4564,N_4471);
nor U4733 (N_4733,N_4451,N_4400);
or U4734 (N_4734,N_4587,N_4468);
and U4735 (N_4735,N_4455,N_4565);
nor U4736 (N_4736,N_4490,N_4521);
nor U4737 (N_4737,N_4531,N_4421);
xor U4738 (N_4738,N_4537,N_4532);
nor U4739 (N_4739,N_4542,N_4537);
and U4740 (N_4740,N_4571,N_4527);
nor U4741 (N_4741,N_4585,N_4512);
nor U4742 (N_4742,N_4487,N_4581);
and U4743 (N_4743,N_4497,N_4458);
xor U4744 (N_4744,N_4583,N_4498);
nand U4745 (N_4745,N_4474,N_4539);
and U4746 (N_4746,N_4567,N_4441);
xnor U4747 (N_4747,N_4457,N_4552);
or U4748 (N_4748,N_4549,N_4494);
and U4749 (N_4749,N_4516,N_4595);
xnor U4750 (N_4750,N_4590,N_4596);
and U4751 (N_4751,N_4594,N_4531);
nand U4752 (N_4752,N_4445,N_4406);
or U4753 (N_4753,N_4453,N_4415);
nor U4754 (N_4754,N_4548,N_4491);
and U4755 (N_4755,N_4497,N_4479);
and U4756 (N_4756,N_4572,N_4467);
or U4757 (N_4757,N_4501,N_4442);
xor U4758 (N_4758,N_4519,N_4549);
and U4759 (N_4759,N_4432,N_4555);
or U4760 (N_4760,N_4497,N_4423);
nand U4761 (N_4761,N_4545,N_4543);
and U4762 (N_4762,N_4470,N_4567);
or U4763 (N_4763,N_4487,N_4578);
or U4764 (N_4764,N_4547,N_4584);
nor U4765 (N_4765,N_4436,N_4435);
xor U4766 (N_4766,N_4591,N_4558);
or U4767 (N_4767,N_4473,N_4497);
and U4768 (N_4768,N_4549,N_4596);
and U4769 (N_4769,N_4471,N_4583);
xor U4770 (N_4770,N_4552,N_4544);
and U4771 (N_4771,N_4575,N_4524);
nor U4772 (N_4772,N_4539,N_4440);
xor U4773 (N_4773,N_4588,N_4568);
nand U4774 (N_4774,N_4551,N_4483);
or U4775 (N_4775,N_4533,N_4585);
nand U4776 (N_4776,N_4563,N_4567);
nor U4777 (N_4777,N_4445,N_4557);
nand U4778 (N_4778,N_4555,N_4455);
or U4779 (N_4779,N_4546,N_4590);
or U4780 (N_4780,N_4576,N_4584);
nand U4781 (N_4781,N_4408,N_4539);
xnor U4782 (N_4782,N_4440,N_4589);
nand U4783 (N_4783,N_4558,N_4453);
and U4784 (N_4784,N_4466,N_4433);
and U4785 (N_4785,N_4558,N_4405);
and U4786 (N_4786,N_4407,N_4566);
nor U4787 (N_4787,N_4409,N_4576);
xnor U4788 (N_4788,N_4520,N_4524);
xnor U4789 (N_4789,N_4520,N_4410);
nand U4790 (N_4790,N_4400,N_4522);
nor U4791 (N_4791,N_4401,N_4580);
nand U4792 (N_4792,N_4415,N_4504);
nand U4793 (N_4793,N_4570,N_4466);
or U4794 (N_4794,N_4546,N_4553);
nor U4795 (N_4795,N_4535,N_4466);
and U4796 (N_4796,N_4476,N_4593);
and U4797 (N_4797,N_4476,N_4459);
nand U4798 (N_4798,N_4403,N_4467);
and U4799 (N_4799,N_4429,N_4555);
nor U4800 (N_4800,N_4753,N_4759);
nor U4801 (N_4801,N_4655,N_4679);
xor U4802 (N_4802,N_4796,N_4692);
nor U4803 (N_4803,N_4720,N_4686);
nor U4804 (N_4804,N_4780,N_4631);
xor U4805 (N_4805,N_4701,N_4747);
xnor U4806 (N_4806,N_4710,N_4785);
or U4807 (N_4807,N_4738,N_4647);
and U4808 (N_4808,N_4777,N_4616);
nand U4809 (N_4809,N_4676,N_4607);
nor U4810 (N_4810,N_4706,N_4769);
xnor U4811 (N_4811,N_4755,N_4629);
or U4812 (N_4812,N_4766,N_4661);
xor U4813 (N_4813,N_4762,N_4649);
nor U4814 (N_4814,N_4671,N_4693);
and U4815 (N_4815,N_4688,N_4602);
and U4816 (N_4816,N_4640,N_4719);
xnor U4817 (N_4817,N_4788,N_4713);
xnor U4818 (N_4818,N_4746,N_4767);
and U4819 (N_4819,N_4639,N_4757);
nand U4820 (N_4820,N_4638,N_4623);
or U4821 (N_4821,N_4636,N_4748);
and U4822 (N_4822,N_4600,N_4716);
xor U4823 (N_4823,N_4681,N_4617);
nor U4824 (N_4824,N_4737,N_4756);
xnor U4825 (N_4825,N_4630,N_4749);
nor U4826 (N_4826,N_4615,N_4684);
and U4827 (N_4827,N_4683,N_4610);
nand U4828 (N_4828,N_4694,N_4625);
or U4829 (N_4829,N_4699,N_4744);
nand U4830 (N_4830,N_4611,N_4745);
xor U4831 (N_4831,N_4674,N_4687);
and U4832 (N_4832,N_4726,N_4722);
xnor U4833 (N_4833,N_4714,N_4680);
nor U4834 (N_4834,N_4735,N_4650);
xnor U4835 (N_4835,N_4739,N_4705);
and U4836 (N_4836,N_4606,N_4794);
xor U4837 (N_4837,N_4624,N_4670);
nand U4838 (N_4838,N_4758,N_4613);
and U4839 (N_4839,N_4682,N_4729);
and U4840 (N_4840,N_4743,N_4768);
and U4841 (N_4841,N_4677,N_4678);
and U4842 (N_4842,N_4724,N_4775);
nand U4843 (N_4843,N_4626,N_4695);
nand U4844 (N_4844,N_4628,N_4787);
or U4845 (N_4845,N_4637,N_4761);
or U4846 (N_4846,N_4730,N_4651);
and U4847 (N_4847,N_4782,N_4657);
nand U4848 (N_4848,N_4792,N_4660);
or U4849 (N_4849,N_4642,N_4634);
nor U4850 (N_4850,N_4632,N_4712);
or U4851 (N_4851,N_4786,N_4641);
nor U4852 (N_4852,N_4609,N_4605);
or U4853 (N_4853,N_4668,N_4622);
nand U4854 (N_4854,N_4643,N_4633);
xnor U4855 (N_4855,N_4608,N_4619);
or U4856 (N_4856,N_4635,N_4601);
nand U4857 (N_4857,N_4750,N_4709);
nor U4858 (N_4858,N_4618,N_4763);
nand U4859 (N_4859,N_4715,N_4793);
nor U4860 (N_4860,N_4778,N_4790);
xor U4861 (N_4861,N_4659,N_4789);
nand U4862 (N_4862,N_4603,N_4673);
nand U4863 (N_4863,N_4653,N_4760);
or U4864 (N_4864,N_4667,N_4742);
nor U4865 (N_4865,N_4690,N_4654);
and U4866 (N_4866,N_4741,N_4644);
xor U4867 (N_4867,N_4791,N_4799);
xnor U4868 (N_4868,N_4685,N_4752);
xor U4869 (N_4869,N_4736,N_4703);
or U4870 (N_4870,N_4740,N_4721);
and U4871 (N_4871,N_4765,N_4689);
xnor U4872 (N_4872,N_4697,N_4732);
xnor U4873 (N_4873,N_4773,N_4734);
nand U4874 (N_4874,N_4604,N_4731);
or U4875 (N_4875,N_4648,N_4621);
or U4876 (N_4876,N_4784,N_4774);
xnor U4877 (N_4877,N_4658,N_4620);
nand U4878 (N_4878,N_4797,N_4718);
and U4879 (N_4879,N_4675,N_4795);
and U4880 (N_4880,N_4771,N_4754);
and U4881 (N_4881,N_4711,N_4770);
nor U4882 (N_4882,N_4727,N_4776);
and U4883 (N_4883,N_4725,N_4696);
nor U4884 (N_4884,N_4783,N_4672);
xnor U4885 (N_4885,N_4691,N_4707);
and U4886 (N_4886,N_4627,N_4698);
nor U4887 (N_4887,N_4779,N_4700);
and U4888 (N_4888,N_4798,N_4733);
or U4889 (N_4889,N_4662,N_4764);
xnor U4890 (N_4890,N_4663,N_4702);
xnor U4891 (N_4891,N_4717,N_4645);
or U4892 (N_4892,N_4652,N_4704);
and U4893 (N_4893,N_4612,N_4751);
xor U4894 (N_4894,N_4646,N_4669);
nand U4895 (N_4895,N_4708,N_4664);
or U4896 (N_4896,N_4723,N_4614);
xor U4897 (N_4897,N_4666,N_4656);
nor U4898 (N_4898,N_4772,N_4665);
or U4899 (N_4899,N_4728,N_4781);
or U4900 (N_4900,N_4798,N_4636);
nand U4901 (N_4901,N_4788,N_4628);
nand U4902 (N_4902,N_4721,N_4760);
or U4903 (N_4903,N_4624,N_4771);
or U4904 (N_4904,N_4798,N_4625);
or U4905 (N_4905,N_4615,N_4643);
xnor U4906 (N_4906,N_4712,N_4780);
and U4907 (N_4907,N_4753,N_4660);
nand U4908 (N_4908,N_4779,N_4747);
and U4909 (N_4909,N_4797,N_4756);
xnor U4910 (N_4910,N_4742,N_4618);
nor U4911 (N_4911,N_4719,N_4795);
or U4912 (N_4912,N_4746,N_4620);
nand U4913 (N_4913,N_4653,N_4797);
xor U4914 (N_4914,N_4799,N_4727);
nand U4915 (N_4915,N_4727,N_4710);
or U4916 (N_4916,N_4651,N_4765);
xor U4917 (N_4917,N_4652,N_4769);
nand U4918 (N_4918,N_4618,N_4631);
nor U4919 (N_4919,N_4794,N_4659);
xor U4920 (N_4920,N_4606,N_4692);
or U4921 (N_4921,N_4661,N_4613);
and U4922 (N_4922,N_4701,N_4639);
or U4923 (N_4923,N_4628,N_4731);
xnor U4924 (N_4924,N_4792,N_4699);
xnor U4925 (N_4925,N_4750,N_4731);
xor U4926 (N_4926,N_4677,N_4698);
nor U4927 (N_4927,N_4656,N_4667);
nand U4928 (N_4928,N_4761,N_4732);
nand U4929 (N_4929,N_4669,N_4752);
or U4930 (N_4930,N_4762,N_4659);
or U4931 (N_4931,N_4610,N_4732);
and U4932 (N_4932,N_4767,N_4757);
or U4933 (N_4933,N_4732,N_4793);
nor U4934 (N_4934,N_4794,N_4770);
nand U4935 (N_4935,N_4695,N_4733);
xor U4936 (N_4936,N_4627,N_4648);
xor U4937 (N_4937,N_4640,N_4708);
and U4938 (N_4938,N_4732,N_4615);
nand U4939 (N_4939,N_4660,N_4688);
nor U4940 (N_4940,N_4722,N_4785);
or U4941 (N_4941,N_4702,N_4631);
nand U4942 (N_4942,N_4603,N_4634);
xor U4943 (N_4943,N_4734,N_4657);
xor U4944 (N_4944,N_4715,N_4757);
nand U4945 (N_4945,N_4737,N_4622);
and U4946 (N_4946,N_4788,N_4682);
nor U4947 (N_4947,N_4636,N_4677);
nor U4948 (N_4948,N_4691,N_4696);
nand U4949 (N_4949,N_4730,N_4793);
nand U4950 (N_4950,N_4672,N_4650);
nor U4951 (N_4951,N_4646,N_4618);
or U4952 (N_4952,N_4725,N_4730);
and U4953 (N_4953,N_4679,N_4740);
nor U4954 (N_4954,N_4662,N_4700);
and U4955 (N_4955,N_4719,N_4617);
nand U4956 (N_4956,N_4765,N_4720);
nand U4957 (N_4957,N_4648,N_4732);
and U4958 (N_4958,N_4698,N_4720);
nor U4959 (N_4959,N_4691,N_4760);
or U4960 (N_4960,N_4737,N_4620);
nor U4961 (N_4961,N_4792,N_4647);
nor U4962 (N_4962,N_4757,N_4700);
nand U4963 (N_4963,N_4678,N_4666);
nand U4964 (N_4964,N_4683,N_4667);
or U4965 (N_4965,N_4675,N_4770);
nor U4966 (N_4966,N_4781,N_4664);
xor U4967 (N_4967,N_4664,N_4711);
xor U4968 (N_4968,N_4766,N_4645);
and U4969 (N_4969,N_4715,N_4627);
xnor U4970 (N_4970,N_4654,N_4635);
nor U4971 (N_4971,N_4635,N_4770);
nor U4972 (N_4972,N_4712,N_4677);
and U4973 (N_4973,N_4697,N_4739);
nor U4974 (N_4974,N_4706,N_4717);
nand U4975 (N_4975,N_4772,N_4639);
nand U4976 (N_4976,N_4701,N_4771);
nand U4977 (N_4977,N_4680,N_4654);
nand U4978 (N_4978,N_4763,N_4775);
nand U4979 (N_4979,N_4773,N_4710);
xor U4980 (N_4980,N_4795,N_4615);
and U4981 (N_4981,N_4607,N_4604);
nor U4982 (N_4982,N_4730,N_4616);
or U4983 (N_4983,N_4681,N_4786);
nand U4984 (N_4984,N_4725,N_4609);
nor U4985 (N_4985,N_4647,N_4613);
xnor U4986 (N_4986,N_4654,N_4774);
and U4987 (N_4987,N_4644,N_4685);
and U4988 (N_4988,N_4763,N_4746);
and U4989 (N_4989,N_4609,N_4769);
or U4990 (N_4990,N_4777,N_4754);
and U4991 (N_4991,N_4645,N_4744);
nor U4992 (N_4992,N_4716,N_4781);
nand U4993 (N_4993,N_4798,N_4631);
or U4994 (N_4994,N_4735,N_4785);
nor U4995 (N_4995,N_4793,N_4789);
xor U4996 (N_4996,N_4757,N_4710);
nor U4997 (N_4997,N_4665,N_4750);
or U4998 (N_4998,N_4778,N_4628);
or U4999 (N_4999,N_4628,N_4762);
and U5000 (N_5000,N_4943,N_4822);
nor U5001 (N_5001,N_4934,N_4996);
xnor U5002 (N_5002,N_4995,N_4868);
or U5003 (N_5003,N_4832,N_4931);
nand U5004 (N_5004,N_4951,N_4813);
nand U5005 (N_5005,N_4829,N_4876);
nor U5006 (N_5006,N_4836,N_4979);
or U5007 (N_5007,N_4874,N_4940);
and U5008 (N_5008,N_4916,N_4816);
nand U5009 (N_5009,N_4877,N_4898);
nand U5010 (N_5010,N_4911,N_4809);
or U5011 (N_5011,N_4972,N_4899);
xor U5012 (N_5012,N_4805,N_4867);
xnor U5013 (N_5013,N_4992,N_4850);
xnor U5014 (N_5014,N_4925,N_4861);
and U5015 (N_5015,N_4833,N_4930);
or U5016 (N_5016,N_4962,N_4878);
or U5017 (N_5017,N_4844,N_4970);
or U5018 (N_5018,N_4839,N_4815);
and U5019 (N_5019,N_4825,N_4827);
xor U5020 (N_5020,N_4862,N_4982);
xnor U5021 (N_5021,N_4986,N_4887);
xor U5022 (N_5022,N_4977,N_4855);
xnor U5023 (N_5023,N_4811,N_4854);
and U5024 (N_5024,N_4849,N_4923);
xor U5025 (N_5025,N_4856,N_4921);
xor U5026 (N_5026,N_4935,N_4913);
nor U5027 (N_5027,N_4924,N_4857);
nand U5028 (N_5028,N_4946,N_4869);
and U5029 (N_5029,N_4910,N_4864);
or U5030 (N_5030,N_4853,N_4893);
nor U5031 (N_5031,N_4941,N_4994);
nand U5032 (N_5032,N_4831,N_4875);
nor U5033 (N_5033,N_4843,N_4882);
xor U5034 (N_5034,N_4858,N_4880);
or U5035 (N_5035,N_4942,N_4947);
nor U5036 (N_5036,N_4802,N_4957);
or U5037 (N_5037,N_4803,N_4965);
nor U5038 (N_5038,N_4976,N_4903);
nor U5039 (N_5039,N_4914,N_4800);
or U5040 (N_5040,N_4840,N_4929);
xor U5041 (N_5041,N_4901,N_4985);
or U5042 (N_5042,N_4902,N_4904);
or U5043 (N_5043,N_4889,N_4872);
xor U5044 (N_5044,N_4975,N_4871);
nor U5045 (N_5045,N_4961,N_4888);
and U5046 (N_5046,N_4884,N_4828);
nand U5047 (N_5047,N_4971,N_4955);
and U5048 (N_5048,N_4989,N_4915);
xor U5049 (N_5049,N_4860,N_4895);
or U5050 (N_5050,N_4906,N_4987);
nor U5051 (N_5051,N_4936,N_4973);
nand U5052 (N_5052,N_4966,N_4993);
and U5053 (N_5053,N_4919,N_4846);
nor U5054 (N_5054,N_4883,N_4808);
or U5055 (N_5055,N_4963,N_4819);
nor U5056 (N_5056,N_4845,N_4807);
xnor U5057 (N_5057,N_4907,N_4909);
nand U5058 (N_5058,N_4848,N_4926);
or U5059 (N_5059,N_4897,N_4852);
nor U5060 (N_5060,N_4870,N_4806);
or U5061 (N_5061,N_4933,N_4959);
and U5062 (N_5062,N_4842,N_4964);
or U5063 (N_5063,N_4981,N_4801);
xor U5064 (N_5064,N_4841,N_4824);
nor U5065 (N_5065,N_4866,N_4810);
xor U5066 (N_5066,N_4863,N_4918);
nor U5067 (N_5067,N_4873,N_4818);
nor U5068 (N_5068,N_4920,N_4837);
or U5069 (N_5069,N_4859,N_4894);
nor U5070 (N_5070,N_4958,N_4980);
and U5071 (N_5071,N_4838,N_4988);
or U5072 (N_5072,N_4984,N_4983);
nand U5073 (N_5073,N_4890,N_4812);
xor U5074 (N_5074,N_4851,N_4820);
nor U5075 (N_5075,N_4952,N_4881);
xor U5076 (N_5076,N_4967,N_4932);
or U5077 (N_5077,N_4990,N_4922);
or U5078 (N_5078,N_4956,N_4847);
and U5079 (N_5079,N_4891,N_4991);
nand U5080 (N_5080,N_4835,N_4998);
or U5081 (N_5081,N_4969,N_4939);
nand U5082 (N_5082,N_4826,N_4950);
and U5083 (N_5083,N_4821,N_4949);
xor U5084 (N_5084,N_4948,N_4978);
or U5085 (N_5085,N_4908,N_4945);
or U5086 (N_5086,N_4927,N_4896);
xnor U5087 (N_5087,N_4917,N_4886);
and U5088 (N_5088,N_4960,N_4944);
nand U5089 (N_5089,N_4823,N_4834);
nand U5090 (N_5090,N_4968,N_4954);
and U5091 (N_5091,N_4928,N_4830);
nand U5092 (N_5092,N_4937,N_4905);
or U5093 (N_5093,N_4892,N_4814);
or U5094 (N_5094,N_4804,N_4974);
or U5095 (N_5095,N_4865,N_4817);
nor U5096 (N_5096,N_4938,N_4900);
and U5097 (N_5097,N_4885,N_4953);
and U5098 (N_5098,N_4997,N_4912);
xor U5099 (N_5099,N_4999,N_4879);
nor U5100 (N_5100,N_4812,N_4813);
nor U5101 (N_5101,N_4846,N_4957);
nand U5102 (N_5102,N_4964,N_4863);
xnor U5103 (N_5103,N_4920,N_4864);
nor U5104 (N_5104,N_4960,N_4829);
xnor U5105 (N_5105,N_4927,N_4816);
nand U5106 (N_5106,N_4815,N_4887);
nor U5107 (N_5107,N_4945,N_4941);
xnor U5108 (N_5108,N_4928,N_4991);
xor U5109 (N_5109,N_4826,N_4866);
nor U5110 (N_5110,N_4965,N_4837);
xor U5111 (N_5111,N_4962,N_4849);
xor U5112 (N_5112,N_4907,N_4861);
xnor U5113 (N_5113,N_4958,N_4846);
and U5114 (N_5114,N_4914,N_4845);
or U5115 (N_5115,N_4896,N_4955);
xnor U5116 (N_5116,N_4904,N_4892);
or U5117 (N_5117,N_4837,N_4853);
nor U5118 (N_5118,N_4871,N_4951);
nand U5119 (N_5119,N_4821,N_4905);
xor U5120 (N_5120,N_4927,N_4939);
or U5121 (N_5121,N_4838,N_4952);
nand U5122 (N_5122,N_4958,N_4876);
and U5123 (N_5123,N_4906,N_4845);
nor U5124 (N_5124,N_4893,N_4832);
or U5125 (N_5125,N_4863,N_4938);
xnor U5126 (N_5126,N_4981,N_4909);
nand U5127 (N_5127,N_4995,N_4964);
and U5128 (N_5128,N_4950,N_4981);
xnor U5129 (N_5129,N_4965,N_4978);
nand U5130 (N_5130,N_4894,N_4993);
nand U5131 (N_5131,N_4859,N_4858);
nor U5132 (N_5132,N_4968,N_4852);
xnor U5133 (N_5133,N_4834,N_4897);
nor U5134 (N_5134,N_4926,N_4961);
nor U5135 (N_5135,N_4997,N_4999);
xnor U5136 (N_5136,N_4983,N_4830);
xnor U5137 (N_5137,N_4889,N_4845);
or U5138 (N_5138,N_4845,N_4881);
and U5139 (N_5139,N_4805,N_4988);
nor U5140 (N_5140,N_4876,N_4971);
nand U5141 (N_5141,N_4809,N_4937);
xnor U5142 (N_5142,N_4910,N_4871);
or U5143 (N_5143,N_4998,N_4806);
or U5144 (N_5144,N_4856,N_4922);
nand U5145 (N_5145,N_4867,N_4987);
and U5146 (N_5146,N_4925,N_4922);
nor U5147 (N_5147,N_4906,N_4994);
nor U5148 (N_5148,N_4892,N_4943);
and U5149 (N_5149,N_4821,N_4868);
or U5150 (N_5150,N_4820,N_4941);
xor U5151 (N_5151,N_4812,N_4950);
nand U5152 (N_5152,N_4914,N_4876);
or U5153 (N_5153,N_4940,N_4953);
or U5154 (N_5154,N_4938,N_4953);
nand U5155 (N_5155,N_4967,N_4976);
xnor U5156 (N_5156,N_4800,N_4995);
nor U5157 (N_5157,N_4961,N_4927);
nand U5158 (N_5158,N_4826,N_4952);
nor U5159 (N_5159,N_4902,N_4907);
nor U5160 (N_5160,N_4968,N_4904);
xor U5161 (N_5161,N_4936,N_4958);
or U5162 (N_5162,N_4801,N_4895);
nand U5163 (N_5163,N_4906,N_4803);
and U5164 (N_5164,N_4961,N_4817);
and U5165 (N_5165,N_4895,N_4936);
and U5166 (N_5166,N_4885,N_4952);
and U5167 (N_5167,N_4846,N_4820);
and U5168 (N_5168,N_4973,N_4852);
or U5169 (N_5169,N_4945,N_4825);
or U5170 (N_5170,N_4887,N_4945);
xnor U5171 (N_5171,N_4957,N_4903);
nand U5172 (N_5172,N_4906,N_4957);
or U5173 (N_5173,N_4855,N_4861);
nor U5174 (N_5174,N_4950,N_4922);
nor U5175 (N_5175,N_4829,N_4935);
xnor U5176 (N_5176,N_4966,N_4883);
nor U5177 (N_5177,N_4954,N_4882);
and U5178 (N_5178,N_4919,N_4970);
nor U5179 (N_5179,N_4841,N_4819);
xnor U5180 (N_5180,N_4906,N_4842);
or U5181 (N_5181,N_4847,N_4977);
xor U5182 (N_5182,N_4850,N_4817);
nand U5183 (N_5183,N_4931,N_4857);
nand U5184 (N_5184,N_4958,N_4922);
nor U5185 (N_5185,N_4832,N_4916);
or U5186 (N_5186,N_4801,N_4955);
xor U5187 (N_5187,N_4962,N_4841);
xnor U5188 (N_5188,N_4968,N_4919);
nand U5189 (N_5189,N_4867,N_4869);
and U5190 (N_5190,N_4998,N_4876);
and U5191 (N_5191,N_4846,N_4801);
and U5192 (N_5192,N_4906,N_4826);
or U5193 (N_5193,N_4957,N_4853);
nand U5194 (N_5194,N_4923,N_4833);
nor U5195 (N_5195,N_4984,N_4929);
nor U5196 (N_5196,N_4855,N_4901);
nor U5197 (N_5197,N_4936,N_4851);
and U5198 (N_5198,N_4833,N_4862);
nor U5199 (N_5199,N_4953,N_4979);
or U5200 (N_5200,N_5010,N_5142);
or U5201 (N_5201,N_5018,N_5144);
nand U5202 (N_5202,N_5091,N_5140);
nand U5203 (N_5203,N_5190,N_5128);
xor U5204 (N_5204,N_5112,N_5113);
xor U5205 (N_5205,N_5141,N_5179);
nor U5206 (N_5206,N_5007,N_5106);
and U5207 (N_5207,N_5092,N_5115);
xnor U5208 (N_5208,N_5148,N_5089);
nor U5209 (N_5209,N_5118,N_5064);
and U5210 (N_5210,N_5097,N_5029);
xnor U5211 (N_5211,N_5172,N_5197);
xor U5212 (N_5212,N_5182,N_5013);
nor U5213 (N_5213,N_5024,N_5124);
nor U5214 (N_5214,N_5175,N_5105);
and U5215 (N_5215,N_5099,N_5093);
or U5216 (N_5216,N_5102,N_5178);
and U5217 (N_5217,N_5021,N_5187);
nor U5218 (N_5218,N_5169,N_5137);
nor U5219 (N_5219,N_5146,N_5065);
xor U5220 (N_5220,N_5167,N_5181);
nand U5221 (N_5221,N_5051,N_5038);
and U5222 (N_5222,N_5012,N_5121);
or U5223 (N_5223,N_5080,N_5019);
nand U5224 (N_5224,N_5067,N_5173);
nand U5225 (N_5225,N_5189,N_5101);
nor U5226 (N_5226,N_5071,N_5129);
xor U5227 (N_5227,N_5006,N_5163);
xnor U5228 (N_5228,N_5005,N_5035);
xnor U5229 (N_5229,N_5122,N_5055);
nor U5230 (N_5230,N_5104,N_5094);
and U5231 (N_5231,N_5161,N_5083);
or U5232 (N_5232,N_5044,N_5098);
and U5233 (N_5233,N_5086,N_5192);
nand U5234 (N_5234,N_5139,N_5174);
xnor U5235 (N_5235,N_5068,N_5108);
and U5236 (N_5236,N_5009,N_5049);
nand U5237 (N_5237,N_5156,N_5147);
nor U5238 (N_5238,N_5033,N_5057);
nand U5239 (N_5239,N_5069,N_5061);
nor U5240 (N_5240,N_5082,N_5131);
or U5241 (N_5241,N_5053,N_5070);
and U5242 (N_5242,N_5001,N_5056);
xor U5243 (N_5243,N_5031,N_5088);
and U5244 (N_5244,N_5123,N_5133);
xnor U5245 (N_5245,N_5110,N_5165);
nor U5246 (N_5246,N_5109,N_5151);
and U5247 (N_5247,N_5039,N_5183);
nor U5248 (N_5248,N_5134,N_5062);
nor U5249 (N_5249,N_5160,N_5117);
nand U5250 (N_5250,N_5095,N_5125);
nand U5251 (N_5251,N_5199,N_5048);
nor U5252 (N_5252,N_5132,N_5041);
nand U5253 (N_5253,N_5008,N_5025);
xor U5254 (N_5254,N_5042,N_5162);
nand U5255 (N_5255,N_5020,N_5046);
and U5256 (N_5256,N_5050,N_5157);
or U5257 (N_5257,N_5194,N_5154);
xor U5258 (N_5258,N_5196,N_5130);
xnor U5259 (N_5259,N_5164,N_5054);
nand U5260 (N_5260,N_5177,N_5026);
xnor U5261 (N_5261,N_5153,N_5058);
xnor U5262 (N_5262,N_5000,N_5060);
xnor U5263 (N_5263,N_5032,N_5120);
nor U5264 (N_5264,N_5081,N_5073);
or U5265 (N_5265,N_5036,N_5176);
or U5266 (N_5266,N_5184,N_5072);
nor U5267 (N_5267,N_5103,N_5087);
xor U5268 (N_5268,N_5168,N_5047);
nand U5269 (N_5269,N_5111,N_5074);
nor U5270 (N_5270,N_5066,N_5180);
nor U5271 (N_5271,N_5107,N_5002);
or U5272 (N_5272,N_5059,N_5185);
nand U5273 (N_5273,N_5126,N_5004);
or U5274 (N_5274,N_5127,N_5014);
and U5275 (N_5275,N_5052,N_5150);
xor U5276 (N_5276,N_5037,N_5076);
nor U5277 (N_5277,N_5034,N_5043);
nand U5278 (N_5278,N_5016,N_5186);
or U5279 (N_5279,N_5030,N_5096);
or U5280 (N_5280,N_5166,N_5155);
and U5281 (N_5281,N_5170,N_5045);
and U5282 (N_5282,N_5193,N_5022);
nor U5283 (N_5283,N_5138,N_5100);
nor U5284 (N_5284,N_5090,N_5063);
and U5285 (N_5285,N_5171,N_5017);
and U5286 (N_5286,N_5078,N_5023);
xnor U5287 (N_5287,N_5011,N_5040);
nor U5288 (N_5288,N_5015,N_5135);
and U5289 (N_5289,N_5158,N_5145);
nand U5290 (N_5290,N_5003,N_5075);
or U5291 (N_5291,N_5116,N_5079);
or U5292 (N_5292,N_5188,N_5085);
nor U5293 (N_5293,N_5195,N_5077);
xnor U5294 (N_5294,N_5028,N_5119);
and U5295 (N_5295,N_5191,N_5084);
nor U5296 (N_5296,N_5198,N_5159);
nor U5297 (N_5297,N_5152,N_5114);
nor U5298 (N_5298,N_5136,N_5143);
and U5299 (N_5299,N_5027,N_5149);
nand U5300 (N_5300,N_5051,N_5117);
xor U5301 (N_5301,N_5094,N_5031);
nand U5302 (N_5302,N_5092,N_5151);
nor U5303 (N_5303,N_5074,N_5110);
xor U5304 (N_5304,N_5164,N_5110);
nand U5305 (N_5305,N_5163,N_5003);
and U5306 (N_5306,N_5177,N_5057);
or U5307 (N_5307,N_5131,N_5186);
nor U5308 (N_5308,N_5195,N_5173);
xor U5309 (N_5309,N_5135,N_5125);
nand U5310 (N_5310,N_5187,N_5041);
nand U5311 (N_5311,N_5091,N_5073);
nand U5312 (N_5312,N_5139,N_5062);
nor U5313 (N_5313,N_5196,N_5072);
or U5314 (N_5314,N_5184,N_5062);
or U5315 (N_5315,N_5179,N_5008);
nand U5316 (N_5316,N_5009,N_5014);
nand U5317 (N_5317,N_5088,N_5087);
and U5318 (N_5318,N_5017,N_5034);
nor U5319 (N_5319,N_5160,N_5068);
nand U5320 (N_5320,N_5015,N_5121);
nor U5321 (N_5321,N_5169,N_5155);
or U5322 (N_5322,N_5173,N_5170);
or U5323 (N_5323,N_5042,N_5010);
and U5324 (N_5324,N_5104,N_5024);
xnor U5325 (N_5325,N_5008,N_5046);
nand U5326 (N_5326,N_5054,N_5096);
and U5327 (N_5327,N_5174,N_5079);
or U5328 (N_5328,N_5146,N_5190);
xnor U5329 (N_5329,N_5048,N_5083);
xnor U5330 (N_5330,N_5085,N_5179);
xor U5331 (N_5331,N_5011,N_5110);
xor U5332 (N_5332,N_5170,N_5050);
or U5333 (N_5333,N_5101,N_5103);
xnor U5334 (N_5334,N_5011,N_5084);
xor U5335 (N_5335,N_5023,N_5178);
nor U5336 (N_5336,N_5194,N_5075);
and U5337 (N_5337,N_5184,N_5188);
nand U5338 (N_5338,N_5111,N_5016);
and U5339 (N_5339,N_5075,N_5150);
nor U5340 (N_5340,N_5161,N_5042);
nand U5341 (N_5341,N_5047,N_5085);
xor U5342 (N_5342,N_5066,N_5129);
xnor U5343 (N_5343,N_5075,N_5170);
and U5344 (N_5344,N_5121,N_5066);
and U5345 (N_5345,N_5058,N_5039);
nand U5346 (N_5346,N_5199,N_5113);
or U5347 (N_5347,N_5096,N_5184);
xor U5348 (N_5348,N_5036,N_5174);
nand U5349 (N_5349,N_5045,N_5149);
or U5350 (N_5350,N_5184,N_5111);
and U5351 (N_5351,N_5072,N_5063);
and U5352 (N_5352,N_5195,N_5178);
xor U5353 (N_5353,N_5150,N_5092);
and U5354 (N_5354,N_5014,N_5115);
xor U5355 (N_5355,N_5154,N_5185);
xnor U5356 (N_5356,N_5042,N_5071);
nor U5357 (N_5357,N_5064,N_5165);
and U5358 (N_5358,N_5191,N_5165);
xnor U5359 (N_5359,N_5060,N_5002);
and U5360 (N_5360,N_5059,N_5138);
nand U5361 (N_5361,N_5158,N_5199);
nor U5362 (N_5362,N_5048,N_5086);
xor U5363 (N_5363,N_5145,N_5147);
nor U5364 (N_5364,N_5107,N_5037);
xnor U5365 (N_5365,N_5009,N_5182);
nand U5366 (N_5366,N_5034,N_5127);
nor U5367 (N_5367,N_5070,N_5045);
and U5368 (N_5368,N_5027,N_5029);
and U5369 (N_5369,N_5001,N_5008);
nand U5370 (N_5370,N_5034,N_5021);
and U5371 (N_5371,N_5036,N_5043);
nor U5372 (N_5372,N_5128,N_5142);
and U5373 (N_5373,N_5127,N_5053);
and U5374 (N_5374,N_5162,N_5182);
and U5375 (N_5375,N_5016,N_5067);
or U5376 (N_5376,N_5191,N_5092);
xor U5377 (N_5377,N_5060,N_5193);
and U5378 (N_5378,N_5012,N_5139);
xnor U5379 (N_5379,N_5085,N_5061);
nor U5380 (N_5380,N_5131,N_5051);
and U5381 (N_5381,N_5118,N_5001);
or U5382 (N_5382,N_5075,N_5017);
or U5383 (N_5383,N_5141,N_5099);
nor U5384 (N_5384,N_5008,N_5185);
xor U5385 (N_5385,N_5007,N_5197);
xor U5386 (N_5386,N_5000,N_5148);
and U5387 (N_5387,N_5183,N_5143);
nor U5388 (N_5388,N_5043,N_5111);
and U5389 (N_5389,N_5129,N_5046);
nand U5390 (N_5390,N_5182,N_5163);
xor U5391 (N_5391,N_5131,N_5038);
nand U5392 (N_5392,N_5077,N_5198);
and U5393 (N_5393,N_5119,N_5120);
and U5394 (N_5394,N_5039,N_5052);
and U5395 (N_5395,N_5126,N_5185);
xnor U5396 (N_5396,N_5196,N_5127);
or U5397 (N_5397,N_5118,N_5125);
or U5398 (N_5398,N_5092,N_5042);
or U5399 (N_5399,N_5022,N_5038);
or U5400 (N_5400,N_5387,N_5346);
nor U5401 (N_5401,N_5386,N_5293);
and U5402 (N_5402,N_5361,N_5333);
xor U5403 (N_5403,N_5235,N_5266);
nand U5404 (N_5404,N_5323,N_5339);
xnor U5405 (N_5405,N_5231,N_5268);
or U5406 (N_5406,N_5320,N_5294);
nand U5407 (N_5407,N_5221,N_5274);
nand U5408 (N_5408,N_5390,N_5314);
nor U5409 (N_5409,N_5232,N_5362);
xor U5410 (N_5410,N_5297,N_5327);
nor U5411 (N_5411,N_5313,N_5223);
nand U5412 (N_5412,N_5256,N_5355);
nand U5413 (N_5413,N_5210,N_5248);
nor U5414 (N_5414,N_5379,N_5318);
and U5415 (N_5415,N_5385,N_5282);
nor U5416 (N_5416,N_5272,N_5321);
xnor U5417 (N_5417,N_5396,N_5352);
or U5418 (N_5418,N_5254,N_5369);
nand U5419 (N_5419,N_5269,N_5204);
xnor U5420 (N_5420,N_5239,N_5317);
nor U5421 (N_5421,N_5226,N_5324);
or U5422 (N_5422,N_5307,N_5374);
nand U5423 (N_5423,N_5329,N_5257);
nor U5424 (N_5424,N_5335,N_5344);
or U5425 (N_5425,N_5222,N_5359);
nor U5426 (N_5426,N_5356,N_5299);
xnor U5427 (N_5427,N_5399,N_5300);
nor U5428 (N_5428,N_5393,N_5380);
nand U5429 (N_5429,N_5206,N_5229);
or U5430 (N_5430,N_5275,N_5236);
nand U5431 (N_5431,N_5276,N_5265);
nor U5432 (N_5432,N_5306,N_5325);
xnor U5433 (N_5433,N_5338,N_5261);
and U5434 (N_5434,N_5383,N_5241);
and U5435 (N_5435,N_5371,N_5331);
xnor U5436 (N_5436,N_5259,N_5215);
xor U5437 (N_5437,N_5243,N_5285);
or U5438 (N_5438,N_5292,N_5308);
nand U5439 (N_5439,N_5301,N_5351);
or U5440 (N_5440,N_5394,N_5234);
or U5441 (N_5441,N_5290,N_5367);
and U5442 (N_5442,N_5279,N_5287);
xor U5443 (N_5443,N_5332,N_5214);
nor U5444 (N_5444,N_5341,N_5263);
nor U5445 (N_5445,N_5357,N_5304);
or U5446 (N_5446,N_5373,N_5382);
nor U5447 (N_5447,N_5247,N_5368);
nand U5448 (N_5448,N_5208,N_5310);
and U5449 (N_5449,N_5364,N_5337);
and U5450 (N_5450,N_5334,N_5233);
or U5451 (N_5451,N_5312,N_5316);
nor U5452 (N_5452,N_5278,N_5209);
and U5453 (N_5453,N_5391,N_5353);
nor U5454 (N_5454,N_5205,N_5258);
or U5455 (N_5455,N_5225,N_5381);
xor U5456 (N_5456,N_5377,N_5271);
xnor U5457 (N_5457,N_5395,N_5200);
or U5458 (N_5458,N_5349,N_5280);
and U5459 (N_5459,N_5207,N_5330);
nand U5460 (N_5460,N_5343,N_5216);
xor U5461 (N_5461,N_5217,N_5267);
and U5462 (N_5462,N_5245,N_5251);
xnor U5463 (N_5463,N_5260,N_5360);
xnor U5464 (N_5464,N_5246,N_5283);
or U5465 (N_5465,N_5220,N_5237);
nor U5466 (N_5466,N_5296,N_5201);
and U5467 (N_5467,N_5262,N_5319);
xnor U5468 (N_5468,N_5302,N_5281);
nand U5469 (N_5469,N_5366,N_5218);
and U5470 (N_5470,N_5326,N_5284);
nor U5471 (N_5471,N_5219,N_5378);
nor U5472 (N_5472,N_5291,N_5264);
and U5473 (N_5473,N_5244,N_5342);
nor U5474 (N_5474,N_5336,N_5348);
nor U5475 (N_5475,N_5384,N_5370);
and U5476 (N_5476,N_5289,N_5340);
or U5477 (N_5477,N_5311,N_5286);
nor U5478 (N_5478,N_5270,N_5238);
and U5479 (N_5479,N_5212,N_5224);
nand U5480 (N_5480,N_5303,N_5288);
and U5481 (N_5481,N_5358,N_5392);
and U5482 (N_5482,N_5249,N_5230);
xnor U5483 (N_5483,N_5255,N_5240);
nor U5484 (N_5484,N_5354,N_5345);
or U5485 (N_5485,N_5277,N_5253);
and U5486 (N_5486,N_5376,N_5322);
nand U5487 (N_5487,N_5372,N_5315);
xnor U5488 (N_5488,N_5389,N_5365);
or U5489 (N_5489,N_5228,N_5388);
xor U5490 (N_5490,N_5213,N_5250);
nor U5491 (N_5491,N_5252,N_5350);
and U5492 (N_5492,N_5328,N_5273);
and U5493 (N_5493,N_5347,N_5309);
nand U5494 (N_5494,N_5398,N_5305);
or U5495 (N_5495,N_5203,N_5227);
and U5496 (N_5496,N_5202,N_5397);
nor U5497 (N_5497,N_5363,N_5298);
xnor U5498 (N_5498,N_5295,N_5375);
or U5499 (N_5499,N_5242,N_5211);
nand U5500 (N_5500,N_5244,N_5399);
or U5501 (N_5501,N_5352,N_5320);
or U5502 (N_5502,N_5211,N_5200);
nor U5503 (N_5503,N_5214,N_5253);
or U5504 (N_5504,N_5376,N_5226);
nor U5505 (N_5505,N_5376,N_5268);
nor U5506 (N_5506,N_5343,N_5321);
xnor U5507 (N_5507,N_5329,N_5302);
or U5508 (N_5508,N_5215,N_5256);
nor U5509 (N_5509,N_5205,N_5213);
nor U5510 (N_5510,N_5293,N_5266);
and U5511 (N_5511,N_5275,N_5324);
and U5512 (N_5512,N_5242,N_5245);
nand U5513 (N_5513,N_5308,N_5374);
or U5514 (N_5514,N_5337,N_5363);
nor U5515 (N_5515,N_5278,N_5280);
or U5516 (N_5516,N_5312,N_5384);
xnor U5517 (N_5517,N_5296,N_5214);
xnor U5518 (N_5518,N_5382,N_5311);
and U5519 (N_5519,N_5236,N_5360);
or U5520 (N_5520,N_5316,N_5398);
and U5521 (N_5521,N_5285,N_5386);
or U5522 (N_5522,N_5249,N_5321);
xor U5523 (N_5523,N_5208,N_5348);
nor U5524 (N_5524,N_5311,N_5314);
nand U5525 (N_5525,N_5298,N_5323);
xnor U5526 (N_5526,N_5272,N_5259);
nand U5527 (N_5527,N_5388,N_5263);
xor U5528 (N_5528,N_5300,N_5362);
nand U5529 (N_5529,N_5246,N_5399);
or U5530 (N_5530,N_5282,N_5213);
and U5531 (N_5531,N_5278,N_5255);
nand U5532 (N_5532,N_5329,N_5300);
or U5533 (N_5533,N_5367,N_5349);
nor U5534 (N_5534,N_5372,N_5387);
and U5535 (N_5535,N_5339,N_5325);
nor U5536 (N_5536,N_5336,N_5390);
nor U5537 (N_5537,N_5298,N_5209);
nor U5538 (N_5538,N_5258,N_5249);
nor U5539 (N_5539,N_5346,N_5312);
nor U5540 (N_5540,N_5328,N_5351);
nor U5541 (N_5541,N_5215,N_5224);
xor U5542 (N_5542,N_5210,N_5316);
and U5543 (N_5543,N_5332,N_5370);
nand U5544 (N_5544,N_5347,N_5224);
xnor U5545 (N_5545,N_5370,N_5388);
and U5546 (N_5546,N_5235,N_5335);
xnor U5547 (N_5547,N_5368,N_5208);
and U5548 (N_5548,N_5235,N_5222);
or U5549 (N_5549,N_5278,N_5367);
xor U5550 (N_5550,N_5271,N_5362);
and U5551 (N_5551,N_5311,N_5250);
nor U5552 (N_5552,N_5221,N_5244);
and U5553 (N_5553,N_5203,N_5302);
nor U5554 (N_5554,N_5236,N_5240);
nand U5555 (N_5555,N_5329,N_5247);
xor U5556 (N_5556,N_5261,N_5207);
xor U5557 (N_5557,N_5247,N_5305);
xor U5558 (N_5558,N_5314,N_5329);
nor U5559 (N_5559,N_5250,N_5298);
nand U5560 (N_5560,N_5263,N_5354);
nor U5561 (N_5561,N_5272,N_5313);
nor U5562 (N_5562,N_5295,N_5256);
xnor U5563 (N_5563,N_5326,N_5350);
nand U5564 (N_5564,N_5284,N_5390);
xor U5565 (N_5565,N_5231,N_5377);
xnor U5566 (N_5566,N_5246,N_5335);
or U5567 (N_5567,N_5342,N_5285);
and U5568 (N_5568,N_5247,N_5323);
or U5569 (N_5569,N_5285,N_5282);
and U5570 (N_5570,N_5312,N_5365);
or U5571 (N_5571,N_5206,N_5325);
nand U5572 (N_5572,N_5340,N_5307);
and U5573 (N_5573,N_5225,N_5388);
nand U5574 (N_5574,N_5369,N_5374);
and U5575 (N_5575,N_5365,N_5275);
and U5576 (N_5576,N_5236,N_5314);
or U5577 (N_5577,N_5257,N_5366);
nand U5578 (N_5578,N_5264,N_5334);
nor U5579 (N_5579,N_5391,N_5280);
nand U5580 (N_5580,N_5370,N_5241);
nor U5581 (N_5581,N_5266,N_5268);
and U5582 (N_5582,N_5239,N_5396);
or U5583 (N_5583,N_5208,N_5241);
nand U5584 (N_5584,N_5334,N_5288);
xnor U5585 (N_5585,N_5368,N_5225);
or U5586 (N_5586,N_5204,N_5387);
nand U5587 (N_5587,N_5315,N_5344);
or U5588 (N_5588,N_5239,N_5283);
and U5589 (N_5589,N_5350,N_5386);
nor U5590 (N_5590,N_5333,N_5222);
or U5591 (N_5591,N_5314,N_5347);
and U5592 (N_5592,N_5264,N_5352);
and U5593 (N_5593,N_5257,N_5327);
nor U5594 (N_5594,N_5202,N_5365);
nand U5595 (N_5595,N_5343,N_5335);
nand U5596 (N_5596,N_5271,N_5369);
or U5597 (N_5597,N_5253,N_5373);
and U5598 (N_5598,N_5355,N_5352);
and U5599 (N_5599,N_5394,N_5329);
nor U5600 (N_5600,N_5510,N_5585);
or U5601 (N_5601,N_5455,N_5506);
nand U5602 (N_5602,N_5565,N_5581);
nor U5603 (N_5603,N_5476,N_5519);
and U5604 (N_5604,N_5497,N_5401);
and U5605 (N_5605,N_5486,N_5549);
xnor U5606 (N_5606,N_5422,N_5590);
xor U5607 (N_5607,N_5515,N_5427);
xor U5608 (N_5608,N_5461,N_5413);
xor U5609 (N_5609,N_5457,N_5584);
xnor U5610 (N_5610,N_5553,N_5542);
nor U5611 (N_5611,N_5552,N_5580);
nor U5612 (N_5612,N_5573,N_5406);
xnor U5613 (N_5613,N_5592,N_5494);
nand U5614 (N_5614,N_5582,N_5561);
nor U5615 (N_5615,N_5591,N_5458);
xor U5616 (N_5616,N_5444,N_5471);
xor U5617 (N_5617,N_5564,N_5452);
or U5618 (N_5618,N_5490,N_5547);
xor U5619 (N_5619,N_5492,N_5480);
xor U5620 (N_5620,N_5501,N_5470);
xor U5621 (N_5621,N_5570,N_5556);
xor U5622 (N_5622,N_5467,N_5560);
or U5623 (N_5623,N_5508,N_5432);
nand U5624 (N_5624,N_5466,N_5438);
nand U5625 (N_5625,N_5571,N_5424);
xnor U5626 (N_5626,N_5563,N_5450);
nor U5627 (N_5627,N_5441,N_5495);
nor U5628 (N_5628,N_5541,N_5437);
or U5629 (N_5629,N_5434,N_5447);
and U5630 (N_5630,N_5483,N_5578);
and U5631 (N_5631,N_5421,N_5576);
nor U5632 (N_5632,N_5416,N_5456);
or U5633 (N_5633,N_5535,N_5558);
or U5634 (N_5634,N_5446,N_5451);
and U5635 (N_5635,N_5513,N_5420);
nand U5636 (N_5636,N_5496,N_5543);
and U5637 (N_5637,N_5472,N_5539);
nand U5638 (N_5638,N_5431,N_5551);
nor U5639 (N_5639,N_5555,N_5598);
and U5640 (N_5640,N_5454,N_5465);
nand U5641 (N_5641,N_5599,N_5531);
nand U5642 (N_5642,N_5514,N_5517);
nand U5643 (N_5643,N_5597,N_5586);
xnor U5644 (N_5644,N_5493,N_5522);
nand U5645 (N_5645,N_5562,N_5426);
nor U5646 (N_5646,N_5469,N_5527);
nand U5647 (N_5647,N_5512,N_5453);
nor U5648 (N_5648,N_5546,N_5418);
nand U5649 (N_5649,N_5588,N_5503);
or U5650 (N_5650,N_5429,N_5489);
nor U5651 (N_5651,N_5462,N_5499);
xor U5652 (N_5652,N_5537,N_5567);
or U5653 (N_5653,N_5464,N_5538);
nand U5654 (N_5654,N_5579,N_5521);
or U5655 (N_5655,N_5593,N_5554);
xnor U5656 (N_5656,N_5491,N_5435);
nor U5657 (N_5657,N_5526,N_5474);
nand U5658 (N_5658,N_5442,N_5568);
or U5659 (N_5659,N_5475,N_5516);
and U5660 (N_5660,N_5544,N_5414);
or U5661 (N_5661,N_5403,N_5595);
xor U5662 (N_5662,N_5507,N_5448);
and U5663 (N_5663,N_5540,N_5463);
or U5664 (N_5664,N_5478,N_5589);
or U5665 (N_5665,N_5459,N_5407);
and U5666 (N_5666,N_5566,N_5504);
nand U5667 (N_5667,N_5410,N_5485);
nor U5668 (N_5668,N_5550,N_5428);
nor U5669 (N_5669,N_5415,N_5572);
and U5670 (N_5670,N_5408,N_5409);
and U5671 (N_5671,N_5502,N_5587);
nor U5672 (N_5672,N_5439,N_5524);
nor U5673 (N_5673,N_5473,N_5430);
and U5674 (N_5674,N_5532,N_5411);
and U5675 (N_5675,N_5569,N_5436);
nor U5676 (N_5676,N_5534,N_5575);
nand U5677 (N_5677,N_5520,N_5594);
and U5678 (N_5678,N_5484,N_5533);
and U5679 (N_5679,N_5412,N_5583);
xnor U5680 (N_5680,N_5518,N_5530);
xor U5681 (N_5681,N_5445,N_5525);
nand U5682 (N_5682,N_5487,N_5557);
nand U5683 (N_5683,N_5400,N_5419);
nand U5684 (N_5684,N_5402,N_5498);
xor U5685 (N_5685,N_5404,N_5468);
and U5686 (N_5686,N_5511,N_5500);
nor U5687 (N_5687,N_5536,N_5577);
and U5688 (N_5688,N_5482,N_5529);
xor U5689 (N_5689,N_5481,N_5449);
or U5690 (N_5690,N_5574,N_5423);
or U5691 (N_5691,N_5488,N_5440);
and U5692 (N_5692,N_5528,N_5405);
nor U5693 (N_5693,N_5460,N_5443);
and U5694 (N_5694,N_5505,N_5559);
and U5695 (N_5695,N_5596,N_5417);
and U5696 (N_5696,N_5477,N_5548);
nor U5697 (N_5697,N_5523,N_5479);
nor U5698 (N_5698,N_5545,N_5433);
nand U5699 (N_5699,N_5509,N_5425);
nor U5700 (N_5700,N_5595,N_5576);
xnor U5701 (N_5701,N_5555,N_5429);
xnor U5702 (N_5702,N_5551,N_5449);
nand U5703 (N_5703,N_5469,N_5575);
or U5704 (N_5704,N_5480,N_5488);
or U5705 (N_5705,N_5446,N_5503);
nor U5706 (N_5706,N_5456,N_5512);
xnor U5707 (N_5707,N_5454,N_5500);
nor U5708 (N_5708,N_5560,N_5542);
and U5709 (N_5709,N_5522,N_5558);
and U5710 (N_5710,N_5540,N_5556);
nor U5711 (N_5711,N_5413,N_5570);
and U5712 (N_5712,N_5442,N_5542);
and U5713 (N_5713,N_5475,N_5451);
or U5714 (N_5714,N_5494,N_5515);
nand U5715 (N_5715,N_5406,N_5432);
or U5716 (N_5716,N_5547,N_5536);
xnor U5717 (N_5717,N_5476,N_5483);
xor U5718 (N_5718,N_5502,N_5437);
xor U5719 (N_5719,N_5463,N_5558);
nand U5720 (N_5720,N_5409,N_5470);
and U5721 (N_5721,N_5458,N_5408);
nor U5722 (N_5722,N_5441,N_5595);
or U5723 (N_5723,N_5412,N_5401);
xnor U5724 (N_5724,N_5492,N_5459);
nor U5725 (N_5725,N_5554,N_5497);
nand U5726 (N_5726,N_5536,N_5506);
or U5727 (N_5727,N_5475,N_5587);
and U5728 (N_5728,N_5565,N_5470);
nor U5729 (N_5729,N_5464,N_5535);
xor U5730 (N_5730,N_5486,N_5552);
nor U5731 (N_5731,N_5536,N_5546);
or U5732 (N_5732,N_5441,N_5527);
nor U5733 (N_5733,N_5538,N_5472);
nand U5734 (N_5734,N_5525,N_5562);
nand U5735 (N_5735,N_5444,N_5483);
nand U5736 (N_5736,N_5448,N_5585);
nand U5737 (N_5737,N_5415,N_5559);
nor U5738 (N_5738,N_5515,N_5509);
nor U5739 (N_5739,N_5499,N_5524);
nand U5740 (N_5740,N_5563,N_5522);
or U5741 (N_5741,N_5528,N_5532);
or U5742 (N_5742,N_5595,N_5408);
nor U5743 (N_5743,N_5429,N_5535);
and U5744 (N_5744,N_5566,N_5478);
or U5745 (N_5745,N_5545,N_5407);
and U5746 (N_5746,N_5545,N_5478);
and U5747 (N_5747,N_5532,N_5515);
nor U5748 (N_5748,N_5592,N_5476);
nand U5749 (N_5749,N_5448,N_5411);
or U5750 (N_5750,N_5479,N_5439);
or U5751 (N_5751,N_5541,N_5570);
or U5752 (N_5752,N_5457,N_5435);
nand U5753 (N_5753,N_5459,N_5544);
xnor U5754 (N_5754,N_5555,N_5579);
nand U5755 (N_5755,N_5533,N_5416);
and U5756 (N_5756,N_5568,N_5472);
xor U5757 (N_5757,N_5571,N_5545);
nor U5758 (N_5758,N_5598,N_5496);
nor U5759 (N_5759,N_5542,N_5535);
xnor U5760 (N_5760,N_5556,N_5436);
nand U5761 (N_5761,N_5507,N_5519);
or U5762 (N_5762,N_5544,N_5489);
xnor U5763 (N_5763,N_5582,N_5576);
xnor U5764 (N_5764,N_5533,N_5594);
and U5765 (N_5765,N_5536,N_5464);
xor U5766 (N_5766,N_5597,N_5400);
nand U5767 (N_5767,N_5433,N_5570);
and U5768 (N_5768,N_5476,N_5536);
nand U5769 (N_5769,N_5516,N_5500);
xor U5770 (N_5770,N_5525,N_5571);
and U5771 (N_5771,N_5548,N_5493);
or U5772 (N_5772,N_5522,N_5530);
nand U5773 (N_5773,N_5531,N_5585);
nand U5774 (N_5774,N_5554,N_5553);
nand U5775 (N_5775,N_5456,N_5443);
nand U5776 (N_5776,N_5551,N_5435);
nor U5777 (N_5777,N_5534,N_5452);
nand U5778 (N_5778,N_5562,N_5457);
nand U5779 (N_5779,N_5535,N_5564);
or U5780 (N_5780,N_5504,N_5547);
nor U5781 (N_5781,N_5578,N_5530);
and U5782 (N_5782,N_5412,N_5540);
nor U5783 (N_5783,N_5580,N_5506);
or U5784 (N_5784,N_5593,N_5420);
nor U5785 (N_5785,N_5444,N_5558);
and U5786 (N_5786,N_5456,N_5445);
or U5787 (N_5787,N_5516,N_5418);
or U5788 (N_5788,N_5556,N_5586);
nor U5789 (N_5789,N_5478,N_5435);
or U5790 (N_5790,N_5432,N_5425);
nor U5791 (N_5791,N_5434,N_5458);
or U5792 (N_5792,N_5596,N_5402);
and U5793 (N_5793,N_5419,N_5406);
xnor U5794 (N_5794,N_5488,N_5452);
and U5795 (N_5795,N_5469,N_5520);
xor U5796 (N_5796,N_5561,N_5420);
nor U5797 (N_5797,N_5572,N_5505);
nor U5798 (N_5798,N_5516,N_5434);
xor U5799 (N_5799,N_5572,N_5419);
and U5800 (N_5800,N_5787,N_5767);
and U5801 (N_5801,N_5789,N_5611);
nand U5802 (N_5802,N_5655,N_5690);
and U5803 (N_5803,N_5790,N_5642);
nor U5804 (N_5804,N_5673,N_5719);
nor U5805 (N_5805,N_5601,N_5630);
and U5806 (N_5806,N_5720,N_5739);
nand U5807 (N_5807,N_5618,N_5710);
and U5808 (N_5808,N_5638,N_5620);
nor U5809 (N_5809,N_5625,N_5712);
or U5810 (N_5810,N_5704,N_5725);
nor U5811 (N_5811,N_5634,N_5771);
or U5812 (N_5812,N_5628,N_5758);
and U5813 (N_5813,N_5766,N_5764);
nor U5814 (N_5814,N_5784,N_5751);
xnor U5815 (N_5815,N_5732,N_5614);
nand U5816 (N_5816,N_5721,N_5747);
or U5817 (N_5817,N_5686,N_5716);
xor U5818 (N_5818,N_5746,N_5694);
and U5819 (N_5819,N_5759,N_5603);
xnor U5820 (N_5820,N_5661,N_5665);
or U5821 (N_5821,N_5714,N_5692);
nand U5822 (N_5822,N_5757,N_5762);
or U5823 (N_5823,N_5668,N_5777);
xnor U5824 (N_5824,N_5627,N_5731);
nor U5825 (N_5825,N_5676,N_5616);
xnor U5826 (N_5826,N_5602,N_5624);
nand U5827 (N_5827,N_5608,N_5640);
and U5828 (N_5828,N_5717,N_5795);
xnor U5829 (N_5829,N_5708,N_5650);
nand U5830 (N_5830,N_5735,N_5631);
xnor U5831 (N_5831,N_5643,N_5670);
nor U5832 (N_5832,N_5781,N_5775);
nand U5833 (N_5833,N_5701,N_5666);
xor U5834 (N_5834,N_5609,N_5632);
nand U5835 (N_5835,N_5730,N_5768);
or U5836 (N_5836,N_5709,N_5700);
xnor U5837 (N_5837,N_5723,N_5754);
nand U5838 (N_5838,N_5707,N_5644);
and U5839 (N_5839,N_5679,N_5606);
nor U5840 (N_5840,N_5617,N_5728);
nor U5841 (N_5841,N_5729,N_5744);
or U5842 (N_5842,N_5683,N_5761);
nor U5843 (N_5843,N_5669,N_5755);
and U5844 (N_5844,N_5741,N_5626);
and U5845 (N_5845,N_5696,N_5615);
and U5846 (N_5846,N_5785,N_5654);
nand U5847 (N_5847,N_5782,N_5693);
or U5848 (N_5848,N_5748,N_5659);
and U5849 (N_5849,N_5718,N_5623);
or U5850 (N_5850,N_5796,N_5791);
xor U5851 (N_5851,N_5786,N_5662);
nor U5852 (N_5852,N_5778,N_5793);
nand U5853 (N_5853,N_5736,N_5687);
nor U5854 (N_5854,N_5733,N_5647);
or U5855 (N_5855,N_5613,N_5672);
nand U5856 (N_5856,N_5619,N_5702);
xor U5857 (N_5857,N_5753,N_5715);
xor U5858 (N_5858,N_5776,N_5722);
or U5859 (N_5859,N_5695,N_5724);
or U5860 (N_5860,N_5671,N_5674);
nor U5861 (N_5861,N_5621,N_5685);
and U5862 (N_5862,N_5773,N_5635);
nand U5863 (N_5863,N_5691,N_5794);
or U5864 (N_5864,N_5798,N_5664);
xor U5865 (N_5865,N_5779,N_5646);
and U5866 (N_5866,N_5726,N_5633);
nand U5867 (N_5867,N_5760,N_5607);
nor U5868 (N_5868,N_5698,N_5610);
nand U5869 (N_5869,N_5689,N_5697);
nand U5870 (N_5870,N_5629,N_5713);
or U5871 (N_5871,N_5651,N_5639);
nand U5872 (N_5872,N_5663,N_5788);
or U5873 (N_5873,N_5641,N_5682);
nand U5874 (N_5874,N_5749,N_5648);
and U5875 (N_5875,N_5675,N_5737);
xnor U5876 (N_5876,N_5765,N_5783);
nor U5877 (N_5877,N_5622,N_5770);
nand U5878 (N_5878,N_5750,N_5792);
nor U5879 (N_5879,N_5660,N_5769);
or U5880 (N_5880,N_5743,N_5774);
nor U5881 (N_5881,N_5645,N_5780);
xor U5882 (N_5882,N_5742,N_5797);
nand U5883 (N_5883,N_5734,N_5703);
xor U5884 (N_5884,N_5667,N_5699);
nand U5885 (N_5885,N_5637,N_5605);
xor U5886 (N_5886,N_5727,N_5740);
nand U5887 (N_5887,N_5711,N_5636);
or U5888 (N_5888,N_5678,N_5752);
or U5889 (N_5889,N_5772,N_5688);
nor U5890 (N_5890,N_5658,N_5677);
or U5891 (N_5891,N_5705,N_5612);
and U5892 (N_5892,N_5656,N_5604);
and U5893 (N_5893,N_5684,N_5657);
nand U5894 (N_5894,N_5680,N_5763);
or U5895 (N_5895,N_5745,N_5652);
nor U5896 (N_5896,N_5681,N_5649);
xor U5897 (N_5897,N_5756,N_5738);
nor U5898 (N_5898,N_5706,N_5653);
and U5899 (N_5899,N_5600,N_5799);
xnor U5900 (N_5900,N_5778,N_5733);
and U5901 (N_5901,N_5753,N_5680);
xor U5902 (N_5902,N_5776,N_5680);
or U5903 (N_5903,N_5739,N_5674);
or U5904 (N_5904,N_5633,N_5605);
xnor U5905 (N_5905,N_5634,N_5669);
and U5906 (N_5906,N_5747,N_5781);
nor U5907 (N_5907,N_5760,N_5653);
xor U5908 (N_5908,N_5769,N_5655);
nand U5909 (N_5909,N_5748,N_5762);
nor U5910 (N_5910,N_5786,N_5644);
and U5911 (N_5911,N_5779,N_5774);
xnor U5912 (N_5912,N_5609,N_5784);
or U5913 (N_5913,N_5793,N_5792);
or U5914 (N_5914,N_5734,N_5773);
or U5915 (N_5915,N_5700,N_5664);
nand U5916 (N_5916,N_5690,N_5684);
nor U5917 (N_5917,N_5685,N_5780);
or U5918 (N_5918,N_5796,N_5636);
nor U5919 (N_5919,N_5784,N_5741);
or U5920 (N_5920,N_5643,N_5796);
nand U5921 (N_5921,N_5760,N_5658);
nor U5922 (N_5922,N_5732,N_5686);
nor U5923 (N_5923,N_5624,N_5751);
nor U5924 (N_5924,N_5767,N_5626);
nor U5925 (N_5925,N_5793,N_5711);
or U5926 (N_5926,N_5793,N_5676);
nor U5927 (N_5927,N_5650,N_5748);
xor U5928 (N_5928,N_5726,N_5713);
or U5929 (N_5929,N_5709,N_5679);
and U5930 (N_5930,N_5697,N_5705);
nand U5931 (N_5931,N_5761,N_5707);
nor U5932 (N_5932,N_5752,N_5670);
and U5933 (N_5933,N_5759,N_5614);
or U5934 (N_5934,N_5633,N_5690);
nand U5935 (N_5935,N_5652,N_5784);
nor U5936 (N_5936,N_5694,N_5728);
and U5937 (N_5937,N_5674,N_5784);
nand U5938 (N_5938,N_5721,N_5639);
nor U5939 (N_5939,N_5691,N_5710);
or U5940 (N_5940,N_5730,N_5726);
xor U5941 (N_5941,N_5625,N_5724);
nand U5942 (N_5942,N_5785,N_5636);
nor U5943 (N_5943,N_5748,N_5760);
or U5944 (N_5944,N_5745,N_5624);
and U5945 (N_5945,N_5713,N_5641);
or U5946 (N_5946,N_5755,N_5775);
xor U5947 (N_5947,N_5741,N_5606);
xor U5948 (N_5948,N_5637,N_5721);
nand U5949 (N_5949,N_5681,N_5608);
and U5950 (N_5950,N_5798,N_5614);
xnor U5951 (N_5951,N_5619,N_5792);
nor U5952 (N_5952,N_5608,N_5782);
xnor U5953 (N_5953,N_5780,N_5667);
or U5954 (N_5954,N_5625,N_5740);
and U5955 (N_5955,N_5778,N_5606);
nand U5956 (N_5956,N_5668,N_5769);
or U5957 (N_5957,N_5713,N_5650);
or U5958 (N_5958,N_5731,N_5637);
xnor U5959 (N_5959,N_5741,N_5780);
nand U5960 (N_5960,N_5791,N_5600);
or U5961 (N_5961,N_5786,N_5624);
nor U5962 (N_5962,N_5743,N_5660);
xor U5963 (N_5963,N_5780,N_5606);
and U5964 (N_5964,N_5740,N_5711);
nor U5965 (N_5965,N_5788,N_5626);
nand U5966 (N_5966,N_5766,N_5623);
xor U5967 (N_5967,N_5767,N_5738);
xnor U5968 (N_5968,N_5689,N_5746);
and U5969 (N_5969,N_5665,N_5691);
and U5970 (N_5970,N_5702,N_5668);
nand U5971 (N_5971,N_5704,N_5669);
nor U5972 (N_5972,N_5768,N_5660);
and U5973 (N_5973,N_5733,N_5624);
and U5974 (N_5974,N_5677,N_5760);
nand U5975 (N_5975,N_5605,N_5727);
nor U5976 (N_5976,N_5734,N_5742);
nand U5977 (N_5977,N_5626,N_5613);
or U5978 (N_5978,N_5634,N_5653);
nand U5979 (N_5979,N_5637,N_5714);
nor U5980 (N_5980,N_5727,N_5777);
or U5981 (N_5981,N_5726,N_5651);
or U5982 (N_5982,N_5790,N_5666);
xnor U5983 (N_5983,N_5665,N_5749);
nand U5984 (N_5984,N_5634,N_5788);
nor U5985 (N_5985,N_5673,N_5683);
nand U5986 (N_5986,N_5785,N_5688);
or U5987 (N_5987,N_5724,N_5634);
nor U5988 (N_5988,N_5749,N_5669);
and U5989 (N_5989,N_5606,N_5768);
xor U5990 (N_5990,N_5691,N_5614);
and U5991 (N_5991,N_5721,N_5719);
xor U5992 (N_5992,N_5756,N_5750);
and U5993 (N_5993,N_5688,N_5685);
and U5994 (N_5994,N_5637,N_5707);
nand U5995 (N_5995,N_5790,N_5791);
or U5996 (N_5996,N_5733,N_5611);
and U5997 (N_5997,N_5637,N_5751);
and U5998 (N_5998,N_5612,N_5660);
nor U5999 (N_5999,N_5697,N_5753);
nand U6000 (N_6000,N_5985,N_5806);
and U6001 (N_6001,N_5822,N_5872);
nor U6002 (N_6002,N_5960,N_5810);
nand U6003 (N_6003,N_5841,N_5910);
or U6004 (N_6004,N_5832,N_5988);
and U6005 (N_6005,N_5840,N_5905);
nor U6006 (N_6006,N_5979,N_5989);
nor U6007 (N_6007,N_5878,N_5833);
nor U6008 (N_6008,N_5811,N_5802);
nand U6009 (N_6009,N_5939,N_5819);
xor U6010 (N_6010,N_5996,N_5858);
xor U6011 (N_6011,N_5909,N_5801);
or U6012 (N_6012,N_5900,N_5886);
and U6013 (N_6013,N_5937,N_5958);
or U6014 (N_6014,N_5834,N_5890);
nand U6015 (N_6015,N_5889,N_5980);
nand U6016 (N_6016,N_5997,N_5827);
nor U6017 (N_6017,N_5826,N_5955);
xor U6018 (N_6018,N_5998,N_5856);
xnor U6019 (N_6019,N_5943,N_5902);
or U6020 (N_6020,N_5863,N_5982);
nand U6021 (N_6021,N_5987,N_5920);
nor U6022 (N_6022,N_5865,N_5869);
and U6023 (N_6023,N_5864,N_5807);
nand U6024 (N_6024,N_5966,N_5950);
and U6025 (N_6025,N_5884,N_5971);
nor U6026 (N_6026,N_5928,N_5887);
nand U6027 (N_6027,N_5927,N_5843);
nor U6028 (N_6028,N_5867,N_5944);
and U6029 (N_6029,N_5963,N_5837);
nand U6030 (N_6030,N_5951,N_5967);
xor U6031 (N_6031,N_5929,N_5804);
nand U6032 (N_6032,N_5809,N_5895);
and U6033 (N_6033,N_5915,N_5981);
and U6034 (N_6034,N_5829,N_5824);
nand U6035 (N_6035,N_5906,N_5954);
and U6036 (N_6036,N_5870,N_5994);
xnor U6037 (N_6037,N_5965,N_5962);
xnor U6038 (N_6038,N_5879,N_5800);
and U6039 (N_6039,N_5855,N_5970);
nor U6040 (N_6040,N_5846,N_5968);
nor U6041 (N_6041,N_5978,N_5896);
xnor U6042 (N_6042,N_5934,N_5861);
or U6043 (N_6043,N_5931,N_5916);
nand U6044 (N_6044,N_5859,N_5977);
nand U6045 (N_6045,N_5918,N_5913);
xnor U6046 (N_6046,N_5991,N_5976);
and U6047 (N_6047,N_5821,N_5930);
nor U6048 (N_6048,N_5877,N_5825);
nor U6049 (N_6049,N_5972,N_5904);
or U6050 (N_6050,N_5844,N_5953);
nand U6051 (N_6051,N_5875,N_5866);
and U6052 (N_6052,N_5961,N_5942);
nand U6053 (N_6053,N_5888,N_5848);
or U6054 (N_6054,N_5813,N_5914);
nor U6055 (N_6055,N_5986,N_5815);
nand U6056 (N_6056,N_5897,N_5993);
and U6057 (N_6057,N_5990,N_5876);
xnor U6058 (N_6058,N_5803,N_5999);
and U6059 (N_6059,N_5830,N_5892);
or U6060 (N_6060,N_5932,N_5828);
and U6061 (N_6061,N_5992,N_5912);
or U6062 (N_6062,N_5818,N_5964);
nor U6063 (N_6063,N_5836,N_5947);
nand U6064 (N_6064,N_5823,N_5862);
or U6065 (N_6065,N_5868,N_5940);
or U6066 (N_6066,N_5917,N_5849);
or U6067 (N_6067,N_5949,N_5894);
and U6068 (N_6068,N_5926,N_5903);
and U6069 (N_6069,N_5919,N_5983);
and U6070 (N_6070,N_5995,N_5885);
nor U6071 (N_6071,N_5839,N_5957);
and U6072 (N_6072,N_5881,N_5974);
nand U6073 (N_6073,N_5899,N_5969);
nand U6074 (N_6074,N_5907,N_5923);
nand U6075 (N_6075,N_5984,N_5874);
xnor U6076 (N_6076,N_5883,N_5973);
xor U6077 (N_6077,N_5945,N_5805);
nor U6078 (N_6078,N_5852,N_5901);
or U6079 (N_6079,N_5835,N_5921);
xor U6080 (N_6080,N_5882,N_5952);
nand U6081 (N_6081,N_5814,N_5941);
nor U6082 (N_6082,N_5851,N_5935);
and U6083 (N_6083,N_5959,N_5831);
and U6084 (N_6084,N_5857,N_5975);
xor U6085 (N_6085,N_5956,N_5880);
or U6086 (N_6086,N_5871,N_5842);
nand U6087 (N_6087,N_5850,N_5938);
or U6088 (N_6088,N_5816,N_5820);
and U6089 (N_6089,N_5845,N_5936);
xor U6090 (N_6090,N_5853,N_5898);
nor U6091 (N_6091,N_5817,N_5812);
xnor U6092 (N_6092,N_5946,N_5924);
and U6093 (N_6093,N_5933,N_5854);
xor U6094 (N_6094,N_5838,N_5922);
and U6095 (N_6095,N_5908,N_5808);
nor U6096 (N_6096,N_5873,N_5948);
or U6097 (N_6097,N_5847,N_5911);
nor U6098 (N_6098,N_5925,N_5893);
or U6099 (N_6099,N_5860,N_5891);
and U6100 (N_6100,N_5808,N_5960);
xnor U6101 (N_6101,N_5988,N_5871);
nor U6102 (N_6102,N_5914,N_5904);
and U6103 (N_6103,N_5865,N_5951);
nand U6104 (N_6104,N_5817,N_5844);
nor U6105 (N_6105,N_5964,N_5887);
and U6106 (N_6106,N_5817,N_5944);
or U6107 (N_6107,N_5927,N_5806);
nor U6108 (N_6108,N_5833,N_5972);
nor U6109 (N_6109,N_5891,N_5988);
and U6110 (N_6110,N_5937,N_5878);
xnor U6111 (N_6111,N_5921,N_5881);
nand U6112 (N_6112,N_5923,N_5949);
nand U6113 (N_6113,N_5885,N_5976);
nand U6114 (N_6114,N_5944,N_5866);
xnor U6115 (N_6115,N_5858,N_5980);
xnor U6116 (N_6116,N_5940,N_5924);
or U6117 (N_6117,N_5841,N_5800);
nor U6118 (N_6118,N_5859,N_5902);
and U6119 (N_6119,N_5961,N_5900);
nand U6120 (N_6120,N_5981,N_5900);
or U6121 (N_6121,N_5807,N_5806);
or U6122 (N_6122,N_5922,N_5983);
nor U6123 (N_6123,N_5864,N_5800);
or U6124 (N_6124,N_5921,N_5966);
nand U6125 (N_6125,N_5975,N_5900);
and U6126 (N_6126,N_5963,N_5815);
nand U6127 (N_6127,N_5907,N_5896);
xor U6128 (N_6128,N_5864,N_5985);
nand U6129 (N_6129,N_5923,N_5821);
and U6130 (N_6130,N_5890,N_5934);
nor U6131 (N_6131,N_5916,N_5844);
and U6132 (N_6132,N_5929,N_5945);
nand U6133 (N_6133,N_5950,N_5866);
nor U6134 (N_6134,N_5923,N_5846);
and U6135 (N_6135,N_5865,N_5837);
xnor U6136 (N_6136,N_5919,N_5953);
or U6137 (N_6137,N_5996,N_5944);
and U6138 (N_6138,N_5908,N_5919);
and U6139 (N_6139,N_5962,N_5899);
xnor U6140 (N_6140,N_5852,N_5820);
nor U6141 (N_6141,N_5980,N_5801);
xor U6142 (N_6142,N_5899,N_5919);
or U6143 (N_6143,N_5984,N_5986);
and U6144 (N_6144,N_5887,N_5813);
and U6145 (N_6145,N_5961,N_5824);
and U6146 (N_6146,N_5967,N_5860);
nand U6147 (N_6147,N_5969,N_5979);
or U6148 (N_6148,N_5803,N_5986);
nand U6149 (N_6149,N_5959,N_5812);
nor U6150 (N_6150,N_5813,N_5840);
nor U6151 (N_6151,N_5846,N_5961);
and U6152 (N_6152,N_5873,N_5946);
nor U6153 (N_6153,N_5868,N_5983);
nand U6154 (N_6154,N_5948,N_5950);
xnor U6155 (N_6155,N_5920,N_5877);
and U6156 (N_6156,N_5931,N_5869);
and U6157 (N_6157,N_5814,N_5959);
and U6158 (N_6158,N_5959,N_5975);
and U6159 (N_6159,N_5903,N_5824);
xor U6160 (N_6160,N_5979,N_5982);
nand U6161 (N_6161,N_5831,N_5802);
and U6162 (N_6162,N_5869,N_5937);
nor U6163 (N_6163,N_5871,N_5890);
nand U6164 (N_6164,N_5914,N_5841);
and U6165 (N_6165,N_5905,N_5903);
nand U6166 (N_6166,N_5966,N_5895);
or U6167 (N_6167,N_5800,N_5973);
or U6168 (N_6168,N_5940,N_5965);
nor U6169 (N_6169,N_5830,N_5876);
xnor U6170 (N_6170,N_5858,N_5956);
xor U6171 (N_6171,N_5871,N_5990);
or U6172 (N_6172,N_5897,N_5964);
and U6173 (N_6173,N_5946,N_5891);
xnor U6174 (N_6174,N_5877,N_5974);
and U6175 (N_6175,N_5918,N_5809);
and U6176 (N_6176,N_5880,N_5928);
xor U6177 (N_6177,N_5815,N_5891);
nor U6178 (N_6178,N_5946,N_5837);
or U6179 (N_6179,N_5831,N_5855);
nand U6180 (N_6180,N_5991,N_5923);
xnor U6181 (N_6181,N_5817,N_5985);
nand U6182 (N_6182,N_5930,N_5815);
xor U6183 (N_6183,N_5864,N_5845);
and U6184 (N_6184,N_5900,N_5927);
nor U6185 (N_6185,N_5962,N_5979);
or U6186 (N_6186,N_5886,N_5840);
xnor U6187 (N_6187,N_5855,N_5901);
xnor U6188 (N_6188,N_5858,N_5907);
or U6189 (N_6189,N_5949,N_5950);
or U6190 (N_6190,N_5965,N_5996);
xor U6191 (N_6191,N_5809,N_5907);
and U6192 (N_6192,N_5820,N_5930);
xnor U6193 (N_6193,N_5929,N_5992);
and U6194 (N_6194,N_5848,N_5931);
or U6195 (N_6195,N_5872,N_5803);
or U6196 (N_6196,N_5869,N_5911);
or U6197 (N_6197,N_5818,N_5929);
nand U6198 (N_6198,N_5853,N_5822);
or U6199 (N_6199,N_5942,N_5992);
nor U6200 (N_6200,N_6106,N_6195);
xnor U6201 (N_6201,N_6126,N_6002);
nor U6202 (N_6202,N_6061,N_6148);
or U6203 (N_6203,N_6004,N_6167);
or U6204 (N_6204,N_6144,N_6054);
and U6205 (N_6205,N_6181,N_6138);
xor U6206 (N_6206,N_6058,N_6119);
nor U6207 (N_6207,N_6162,N_6090);
nor U6208 (N_6208,N_6068,N_6073);
and U6209 (N_6209,N_6011,N_6030);
or U6210 (N_6210,N_6176,N_6182);
nor U6211 (N_6211,N_6093,N_6036);
or U6212 (N_6212,N_6001,N_6077);
and U6213 (N_6213,N_6033,N_6016);
nor U6214 (N_6214,N_6067,N_6059);
nor U6215 (N_6215,N_6187,N_6082);
or U6216 (N_6216,N_6051,N_6183);
nand U6217 (N_6217,N_6198,N_6112);
and U6218 (N_6218,N_6168,N_6013);
xnor U6219 (N_6219,N_6034,N_6153);
nand U6220 (N_6220,N_6110,N_6186);
and U6221 (N_6221,N_6133,N_6015);
xor U6222 (N_6222,N_6164,N_6008);
nand U6223 (N_6223,N_6185,N_6180);
or U6224 (N_6224,N_6146,N_6111);
nand U6225 (N_6225,N_6159,N_6129);
nor U6226 (N_6226,N_6085,N_6042);
and U6227 (N_6227,N_6199,N_6097);
xor U6228 (N_6228,N_6005,N_6116);
or U6229 (N_6229,N_6139,N_6171);
nor U6230 (N_6230,N_6197,N_6184);
or U6231 (N_6231,N_6044,N_6160);
nor U6232 (N_6232,N_6052,N_6057);
or U6233 (N_6233,N_6079,N_6134);
and U6234 (N_6234,N_6192,N_6143);
and U6235 (N_6235,N_6029,N_6190);
nand U6236 (N_6236,N_6047,N_6131);
xor U6237 (N_6237,N_6173,N_6071);
or U6238 (N_6238,N_6132,N_6156);
nand U6239 (N_6239,N_6101,N_6046);
nand U6240 (N_6240,N_6124,N_6194);
and U6241 (N_6241,N_6012,N_6019);
and U6242 (N_6242,N_6069,N_6127);
or U6243 (N_6243,N_6095,N_6084);
nor U6244 (N_6244,N_6125,N_6086);
and U6245 (N_6245,N_6010,N_6123);
and U6246 (N_6246,N_6122,N_6083);
nor U6247 (N_6247,N_6063,N_6107);
nor U6248 (N_6248,N_6128,N_6074);
xor U6249 (N_6249,N_6028,N_6163);
nand U6250 (N_6250,N_6141,N_6024);
and U6251 (N_6251,N_6196,N_6165);
and U6252 (N_6252,N_6121,N_6150);
and U6253 (N_6253,N_6103,N_6161);
nand U6254 (N_6254,N_6092,N_6145);
and U6255 (N_6255,N_6076,N_6050);
or U6256 (N_6256,N_6026,N_6154);
nor U6257 (N_6257,N_6039,N_6035);
or U6258 (N_6258,N_6175,N_6066);
or U6259 (N_6259,N_6078,N_6009);
or U6260 (N_6260,N_6096,N_6191);
nor U6261 (N_6261,N_6064,N_6006);
and U6262 (N_6262,N_6149,N_6018);
or U6263 (N_6263,N_6170,N_6100);
nand U6264 (N_6264,N_6102,N_6089);
nand U6265 (N_6265,N_6023,N_6022);
and U6266 (N_6266,N_6081,N_6087);
nand U6267 (N_6267,N_6178,N_6048);
and U6268 (N_6268,N_6135,N_6055);
and U6269 (N_6269,N_6045,N_6113);
and U6270 (N_6270,N_6040,N_6105);
nor U6271 (N_6271,N_6037,N_6003);
or U6272 (N_6272,N_6031,N_6130);
and U6273 (N_6273,N_6179,N_6080);
nand U6274 (N_6274,N_6169,N_6152);
xor U6275 (N_6275,N_6025,N_6109);
and U6276 (N_6276,N_6104,N_6060);
nand U6277 (N_6277,N_6065,N_6193);
or U6278 (N_6278,N_6114,N_6117);
nor U6279 (N_6279,N_6157,N_6099);
nor U6280 (N_6280,N_6108,N_6174);
and U6281 (N_6281,N_6038,N_6142);
and U6282 (N_6282,N_6155,N_6043);
nand U6283 (N_6283,N_6041,N_6118);
and U6284 (N_6284,N_6136,N_6062);
nand U6285 (N_6285,N_6088,N_6007);
xnor U6286 (N_6286,N_6115,N_6032);
nor U6287 (N_6287,N_6166,N_6091);
xnor U6288 (N_6288,N_6188,N_6056);
nor U6289 (N_6289,N_6000,N_6094);
or U6290 (N_6290,N_6151,N_6140);
nand U6291 (N_6291,N_6137,N_6020);
and U6292 (N_6292,N_6027,N_6172);
nor U6293 (N_6293,N_6189,N_6014);
xnor U6294 (N_6294,N_6070,N_6072);
or U6295 (N_6295,N_6075,N_6098);
nor U6296 (N_6296,N_6120,N_6053);
or U6297 (N_6297,N_6177,N_6158);
nand U6298 (N_6298,N_6049,N_6017);
xnor U6299 (N_6299,N_6147,N_6021);
and U6300 (N_6300,N_6011,N_6039);
or U6301 (N_6301,N_6104,N_6174);
xor U6302 (N_6302,N_6040,N_6098);
nand U6303 (N_6303,N_6121,N_6034);
or U6304 (N_6304,N_6133,N_6058);
nor U6305 (N_6305,N_6138,N_6029);
xnor U6306 (N_6306,N_6052,N_6123);
xnor U6307 (N_6307,N_6073,N_6040);
nor U6308 (N_6308,N_6058,N_6015);
xnor U6309 (N_6309,N_6059,N_6015);
or U6310 (N_6310,N_6187,N_6049);
nand U6311 (N_6311,N_6110,N_6023);
nor U6312 (N_6312,N_6145,N_6064);
nand U6313 (N_6313,N_6039,N_6128);
and U6314 (N_6314,N_6040,N_6171);
xor U6315 (N_6315,N_6143,N_6151);
or U6316 (N_6316,N_6057,N_6174);
and U6317 (N_6317,N_6169,N_6114);
nand U6318 (N_6318,N_6194,N_6030);
xnor U6319 (N_6319,N_6045,N_6050);
xor U6320 (N_6320,N_6145,N_6044);
xnor U6321 (N_6321,N_6166,N_6090);
and U6322 (N_6322,N_6037,N_6039);
or U6323 (N_6323,N_6080,N_6154);
nand U6324 (N_6324,N_6049,N_6051);
and U6325 (N_6325,N_6032,N_6170);
xnor U6326 (N_6326,N_6112,N_6156);
nor U6327 (N_6327,N_6160,N_6117);
nand U6328 (N_6328,N_6154,N_6185);
nor U6329 (N_6329,N_6046,N_6100);
and U6330 (N_6330,N_6197,N_6004);
and U6331 (N_6331,N_6078,N_6178);
and U6332 (N_6332,N_6141,N_6198);
xor U6333 (N_6333,N_6056,N_6131);
and U6334 (N_6334,N_6143,N_6059);
or U6335 (N_6335,N_6129,N_6028);
xnor U6336 (N_6336,N_6182,N_6130);
xor U6337 (N_6337,N_6075,N_6157);
nand U6338 (N_6338,N_6179,N_6118);
nand U6339 (N_6339,N_6142,N_6198);
nor U6340 (N_6340,N_6109,N_6118);
xor U6341 (N_6341,N_6083,N_6159);
nand U6342 (N_6342,N_6125,N_6062);
or U6343 (N_6343,N_6092,N_6167);
xor U6344 (N_6344,N_6019,N_6047);
and U6345 (N_6345,N_6177,N_6148);
xor U6346 (N_6346,N_6073,N_6149);
and U6347 (N_6347,N_6041,N_6069);
xnor U6348 (N_6348,N_6180,N_6171);
nand U6349 (N_6349,N_6112,N_6147);
and U6350 (N_6350,N_6143,N_6052);
nor U6351 (N_6351,N_6190,N_6140);
nand U6352 (N_6352,N_6032,N_6177);
xnor U6353 (N_6353,N_6185,N_6140);
nor U6354 (N_6354,N_6184,N_6018);
xor U6355 (N_6355,N_6012,N_6171);
and U6356 (N_6356,N_6165,N_6029);
nor U6357 (N_6357,N_6095,N_6075);
and U6358 (N_6358,N_6014,N_6086);
nand U6359 (N_6359,N_6194,N_6185);
or U6360 (N_6360,N_6041,N_6086);
nand U6361 (N_6361,N_6130,N_6099);
nor U6362 (N_6362,N_6047,N_6030);
or U6363 (N_6363,N_6155,N_6105);
or U6364 (N_6364,N_6117,N_6170);
and U6365 (N_6365,N_6009,N_6046);
and U6366 (N_6366,N_6195,N_6183);
and U6367 (N_6367,N_6111,N_6128);
nand U6368 (N_6368,N_6046,N_6130);
xnor U6369 (N_6369,N_6130,N_6114);
and U6370 (N_6370,N_6110,N_6046);
or U6371 (N_6371,N_6024,N_6065);
xor U6372 (N_6372,N_6011,N_6111);
xor U6373 (N_6373,N_6050,N_6135);
nor U6374 (N_6374,N_6019,N_6169);
nand U6375 (N_6375,N_6167,N_6081);
nor U6376 (N_6376,N_6177,N_6144);
nor U6377 (N_6377,N_6132,N_6074);
xnor U6378 (N_6378,N_6026,N_6131);
and U6379 (N_6379,N_6156,N_6037);
nand U6380 (N_6380,N_6095,N_6117);
nor U6381 (N_6381,N_6133,N_6054);
nand U6382 (N_6382,N_6005,N_6166);
nand U6383 (N_6383,N_6135,N_6020);
and U6384 (N_6384,N_6019,N_6189);
xor U6385 (N_6385,N_6033,N_6093);
or U6386 (N_6386,N_6105,N_6148);
and U6387 (N_6387,N_6146,N_6145);
or U6388 (N_6388,N_6087,N_6172);
nand U6389 (N_6389,N_6198,N_6143);
nand U6390 (N_6390,N_6126,N_6194);
nor U6391 (N_6391,N_6043,N_6135);
nor U6392 (N_6392,N_6090,N_6035);
and U6393 (N_6393,N_6039,N_6090);
xnor U6394 (N_6394,N_6008,N_6059);
xor U6395 (N_6395,N_6137,N_6033);
nand U6396 (N_6396,N_6117,N_6076);
xor U6397 (N_6397,N_6189,N_6178);
nor U6398 (N_6398,N_6070,N_6105);
nor U6399 (N_6399,N_6195,N_6189);
nor U6400 (N_6400,N_6200,N_6343);
nor U6401 (N_6401,N_6204,N_6206);
nand U6402 (N_6402,N_6370,N_6309);
xnor U6403 (N_6403,N_6313,N_6383);
xnor U6404 (N_6404,N_6306,N_6212);
and U6405 (N_6405,N_6201,N_6341);
xnor U6406 (N_6406,N_6220,N_6258);
nand U6407 (N_6407,N_6355,N_6296);
nor U6408 (N_6408,N_6224,N_6262);
or U6409 (N_6409,N_6269,N_6295);
or U6410 (N_6410,N_6395,N_6356);
nand U6411 (N_6411,N_6273,N_6392);
xnor U6412 (N_6412,N_6297,N_6257);
nor U6413 (N_6413,N_6222,N_6242);
nor U6414 (N_6414,N_6332,N_6333);
or U6415 (N_6415,N_6217,N_6229);
or U6416 (N_6416,N_6219,N_6346);
nand U6417 (N_6417,N_6259,N_6256);
nor U6418 (N_6418,N_6216,N_6228);
nor U6419 (N_6419,N_6300,N_6202);
nand U6420 (N_6420,N_6391,N_6213);
or U6421 (N_6421,N_6267,N_6307);
and U6422 (N_6422,N_6397,N_6365);
nand U6423 (N_6423,N_6246,N_6353);
nand U6424 (N_6424,N_6270,N_6374);
nand U6425 (N_6425,N_6369,N_6239);
nor U6426 (N_6426,N_6208,N_6381);
nand U6427 (N_6427,N_6382,N_6394);
xor U6428 (N_6428,N_6248,N_6203);
and U6429 (N_6429,N_6334,N_6275);
xnor U6430 (N_6430,N_6310,N_6235);
nor U6431 (N_6431,N_6327,N_6266);
nor U6432 (N_6432,N_6260,N_6360);
nor U6433 (N_6433,N_6389,N_6373);
nor U6434 (N_6434,N_6247,N_6322);
or U6435 (N_6435,N_6312,N_6286);
nand U6436 (N_6436,N_6387,N_6323);
and U6437 (N_6437,N_6276,N_6291);
xnor U6438 (N_6438,N_6338,N_6398);
nor U6439 (N_6439,N_6264,N_6372);
nor U6440 (N_6440,N_6284,N_6348);
and U6441 (N_6441,N_6265,N_6301);
and U6442 (N_6442,N_6311,N_6384);
nand U6443 (N_6443,N_6298,N_6320);
nand U6444 (N_6444,N_6350,N_6345);
and U6445 (N_6445,N_6376,N_6349);
xor U6446 (N_6446,N_6240,N_6321);
nand U6447 (N_6447,N_6351,N_6319);
or U6448 (N_6448,N_6302,N_6223);
nand U6449 (N_6449,N_6249,N_6299);
and U6450 (N_6450,N_6364,N_6231);
nor U6451 (N_6451,N_6336,N_6377);
nand U6452 (N_6452,N_6214,N_6324);
nor U6453 (N_6453,N_6316,N_6263);
and U6454 (N_6454,N_6268,N_6358);
nor U6455 (N_6455,N_6388,N_6207);
nand U6456 (N_6456,N_6238,N_6362);
xnor U6457 (N_6457,N_6236,N_6271);
xor U6458 (N_6458,N_6304,N_6234);
and U6459 (N_6459,N_6386,N_6352);
xor U6460 (N_6460,N_6283,N_6314);
nor U6461 (N_6461,N_6308,N_6274);
xnor U6462 (N_6462,N_6385,N_6337);
xor U6463 (N_6463,N_6303,N_6261);
xor U6464 (N_6464,N_6252,N_6230);
or U6465 (N_6465,N_6347,N_6232);
xor U6466 (N_6466,N_6244,N_6254);
or U6467 (N_6467,N_6330,N_6318);
nor U6468 (N_6468,N_6344,N_6294);
and U6469 (N_6469,N_6277,N_6378);
or U6470 (N_6470,N_6237,N_6335);
or U6471 (N_6471,N_6329,N_6226);
nand U6472 (N_6472,N_6280,N_6278);
xor U6473 (N_6473,N_6251,N_6342);
nand U6474 (N_6474,N_6250,N_6288);
and U6475 (N_6475,N_6287,N_6315);
nor U6476 (N_6476,N_6326,N_6357);
or U6477 (N_6477,N_6361,N_6281);
and U6478 (N_6478,N_6210,N_6241);
xnor U6479 (N_6479,N_6255,N_6218);
and U6480 (N_6480,N_6399,N_6340);
and U6481 (N_6481,N_6367,N_6221);
or U6482 (N_6482,N_6375,N_6317);
and U6483 (N_6483,N_6205,N_6290);
xor U6484 (N_6484,N_6289,N_6396);
xor U6485 (N_6485,N_6243,N_6380);
nand U6486 (N_6486,N_6339,N_6359);
or U6487 (N_6487,N_6211,N_6209);
nand U6488 (N_6488,N_6282,N_6390);
nor U6489 (N_6489,N_6371,N_6279);
and U6490 (N_6490,N_6368,N_6393);
nand U6491 (N_6491,N_6305,N_6253);
and U6492 (N_6492,N_6215,N_6331);
nand U6493 (N_6493,N_6233,N_6379);
xor U6494 (N_6494,N_6293,N_6325);
xor U6495 (N_6495,N_6227,N_6328);
and U6496 (N_6496,N_6285,N_6366);
xor U6497 (N_6497,N_6354,N_6363);
xor U6498 (N_6498,N_6272,N_6292);
nand U6499 (N_6499,N_6245,N_6225);
and U6500 (N_6500,N_6255,N_6254);
nand U6501 (N_6501,N_6257,N_6255);
nand U6502 (N_6502,N_6307,N_6251);
and U6503 (N_6503,N_6397,N_6392);
and U6504 (N_6504,N_6287,N_6320);
nand U6505 (N_6505,N_6393,N_6222);
or U6506 (N_6506,N_6301,N_6378);
or U6507 (N_6507,N_6232,N_6378);
xor U6508 (N_6508,N_6329,N_6386);
xnor U6509 (N_6509,N_6391,N_6291);
nand U6510 (N_6510,N_6207,N_6206);
xor U6511 (N_6511,N_6271,N_6223);
or U6512 (N_6512,N_6319,N_6286);
xnor U6513 (N_6513,N_6291,N_6301);
nand U6514 (N_6514,N_6237,N_6322);
and U6515 (N_6515,N_6298,N_6228);
nand U6516 (N_6516,N_6234,N_6348);
xnor U6517 (N_6517,N_6331,N_6241);
nand U6518 (N_6518,N_6383,N_6229);
or U6519 (N_6519,N_6262,N_6202);
xnor U6520 (N_6520,N_6242,N_6254);
nor U6521 (N_6521,N_6239,N_6206);
xor U6522 (N_6522,N_6347,N_6391);
nor U6523 (N_6523,N_6232,N_6390);
nor U6524 (N_6524,N_6222,N_6215);
and U6525 (N_6525,N_6236,N_6357);
xor U6526 (N_6526,N_6223,N_6290);
xor U6527 (N_6527,N_6219,N_6304);
nor U6528 (N_6528,N_6300,N_6219);
xor U6529 (N_6529,N_6226,N_6283);
xor U6530 (N_6530,N_6288,N_6364);
xnor U6531 (N_6531,N_6290,N_6382);
nor U6532 (N_6532,N_6328,N_6301);
and U6533 (N_6533,N_6272,N_6273);
xnor U6534 (N_6534,N_6274,N_6261);
nor U6535 (N_6535,N_6326,N_6277);
xnor U6536 (N_6536,N_6264,N_6325);
xor U6537 (N_6537,N_6266,N_6397);
nor U6538 (N_6538,N_6313,N_6361);
xnor U6539 (N_6539,N_6204,N_6263);
nor U6540 (N_6540,N_6309,N_6252);
nor U6541 (N_6541,N_6280,N_6228);
or U6542 (N_6542,N_6278,N_6392);
nand U6543 (N_6543,N_6329,N_6348);
and U6544 (N_6544,N_6261,N_6310);
xor U6545 (N_6545,N_6334,N_6225);
nand U6546 (N_6546,N_6268,N_6372);
nand U6547 (N_6547,N_6386,N_6381);
or U6548 (N_6548,N_6248,N_6320);
nand U6549 (N_6549,N_6278,N_6219);
xnor U6550 (N_6550,N_6284,N_6233);
nor U6551 (N_6551,N_6252,N_6384);
or U6552 (N_6552,N_6386,N_6294);
and U6553 (N_6553,N_6350,N_6333);
nand U6554 (N_6554,N_6336,N_6304);
or U6555 (N_6555,N_6201,N_6346);
nor U6556 (N_6556,N_6255,N_6223);
or U6557 (N_6557,N_6298,N_6366);
nand U6558 (N_6558,N_6386,N_6373);
nand U6559 (N_6559,N_6384,N_6332);
nand U6560 (N_6560,N_6329,N_6260);
nor U6561 (N_6561,N_6301,N_6228);
or U6562 (N_6562,N_6378,N_6289);
nand U6563 (N_6563,N_6386,N_6364);
or U6564 (N_6564,N_6376,N_6324);
nor U6565 (N_6565,N_6292,N_6274);
nand U6566 (N_6566,N_6296,N_6348);
nor U6567 (N_6567,N_6337,N_6225);
nor U6568 (N_6568,N_6336,N_6378);
nor U6569 (N_6569,N_6338,N_6320);
nor U6570 (N_6570,N_6386,N_6334);
or U6571 (N_6571,N_6231,N_6242);
and U6572 (N_6572,N_6247,N_6229);
or U6573 (N_6573,N_6369,N_6317);
and U6574 (N_6574,N_6260,N_6269);
and U6575 (N_6575,N_6286,N_6214);
and U6576 (N_6576,N_6312,N_6225);
xnor U6577 (N_6577,N_6314,N_6218);
or U6578 (N_6578,N_6383,N_6306);
or U6579 (N_6579,N_6325,N_6335);
and U6580 (N_6580,N_6361,N_6375);
or U6581 (N_6581,N_6248,N_6237);
xor U6582 (N_6582,N_6240,N_6340);
and U6583 (N_6583,N_6311,N_6271);
xnor U6584 (N_6584,N_6273,N_6231);
or U6585 (N_6585,N_6395,N_6375);
xnor U6586 (N_6586,N_6359,N_6256);
xnor U6587 (N_6587,N_6390,N_6249);
and U6588 (N_6588,N_6388,N_6317);
or U6589 (N_6589,N_6319,N_6313);
nand U6590 (N_6590,N_6281,N_6345);
nand U6591 (N_6591,N_6217,N_6243);
and U6592 (N_6592,N_6321,N_6348);
xor U6593 (N_6593,N_6314,N_6336);
or U6594 (N_6594,N_6318,N_6201);
nor U6595 (N_6595,N_6327,N_6252);
xnor U6596 (N_6596,N_6240,N_6261);
xor U6597 (N_6597,N_6285,N_6375);
or U6598 (N_6598,N_6213,N_6257);
nor U6599 (N_6599,N_6215,N_6254);
and U6600 (N_6600,N_6518,N_6428);
nor U6601 (N_6601,N_6484,N_6437);
nand U6602 (N_6602,N_6406,N_6441);
nand U6603 (N_6603,N_6550,N_6508);
xor U6604 (N_6604,N_6528,N_6551);
and U6605 (N_6605,N_6473,N_6521);
nand U6606 (N_6606,N_6458,N_6403);
and U6607 (N_6607,N_6448,N_6542);
nor U6608 (N_6608,N_6444,N_6439);
nand U6609 (N_6609,N_6497,N_6523);
and U6610 (N_6610,N_6558,N_6430);
nand U6611 (N_6611,N_6513,N_6574);
xor U6612 (N_6612,N_6567,N_6548);
nand U6613 (N_6613,N_6522,N_6418);
nor U6614 (N_6614,N_6557,N_6517);
nor U6615 (N_6615,N_6553,N_6405);
nor U6616 (N_6616,N_6472,N_6449);
nor U6617 (N_6617,N_6464,N_6564);
and U6618 (N_6618,N_6594,N_6586);
and U6619 (N_6619,N_6488,N_6531);
nand U6620 (N_6620,N_6493,N_6581);
or U6621 (N_6621,N_6547,N_6544);
nand U6622 (N_6622,N_6585,N_6505);
xnor U6623 (N_6623,N_6571,N_6489);
or U6624 (N_6624,N_6525,N_6582);
nand U6625 (N_6625,N_6541,N_6552);
xor U6626 (N_6626,N_6471,N_6487);
and U6627 (N_6627,N_6535,N_6573);
nand U6628 (N_6628,N_6409,N_6465);
xor U6629 (N_6629,N_6411,N_6483);
or U6630 (N_6630,N_6402,N_6407);
or U6631 (N_6631,N_6534,N_6556);
xnor U6632 (N_6632,N_6529,N_6445);
nand U6633 (N_6633,N_6422,N_6593);
nor U6634 (N_6634,N_6532,N_6587);
nand U6635 (N_6635,N_6579,N_6434);
and U6636 (N_6636,N_6500,N_6492);
nand U6637 (N_6637,N_6530,N_6427);
xnor U6638 (N_6638,N_6527,N_6577);
nand U6639 (N_6639,N_6435,N_6485);
xor U6640 (N_6640,N_6597,N_6503);
nor U6641 (N_6641,N_6561,N_6506);
or U6642 (N_6642,N_6459,N_6545);
xnor U6643 (N_6643,N_6533,N_6447);
nand U6644 (N_6644,N_6537,N_6572);
nor U6645 (N_6645,N_6570,N_6560);
nand U6646 (N_6646,N_6524,N_6494);
or U6647 (N_6647,N_6401,N_6455);
nand U6648 (N_6648,N_6470,N_6596);
or U6649 (N_6649,N_6477,N_6511);
and U6650 (N_6650,N_6568,N_6495);
nand U6651 (N_6651,N_6463,N_6539);
or U6652 (N_6652,N_6466,N_6566);
nor U6653 (N_6653,N_6519,N_6433);
xor U6654 (N_6654,N_6423,N_6520);
or U6655 (N_6655,N_6436,N_6595);
and U6656 (N_6656,N_6486,N_6549);
nor U6657 (N_6657,N_6468,N_6509);
nor U6658 (N_6658,N_6569,N_6588);
nand U6659 (N_6659,N_6443,N_6496);
nand U6660 (N_6660,N_6408,N_6512);
nand U6661 (N_6661,N_6414,N_6559);
xor U6662 (N_6662,N_6478,N_6424);
nand U6663 (N_6663,N_6481,N_6526);
or U6664 (N_6664,N_6546,N_6590);
nand U6665 (N_6665,N_6457,N_6565);
nand U6666 (N_6666,N_6454,N_6499);
or U6667 (N_6667,N_6514,N_6446);
or U6668 (N_6668,N_6507,N_6419);
nand U6669 (N_6669,N_6538,N_6589);
xor U6670 (N_6670,N_6461,N_6562);
and U6671 (N_6671,N_6504,N_6501);
nor U6672 (N_6672,N_6450,N_6469);
nor U6673 (N_6673,N_6479,N_6460);
nor U6674 (N_6674,N_6467,N_6462);
nand U6675 (N_6675,N_6554,N_6515);
and U6676 (N_6676,N_6498,N_6599);
and U6677 (N_6677,N_6555,N_6475);
and U6678 (N_6678,N_6510,N_6591);
nand U6679 (N_6679,N_6563,N_6491);
nor U6680 (N_6680,N_6442,N_6420);
nand U6681 (N_6681,N_6429,N_6516);
and U6682 (N_6682,N_6400,N_6416);
nor U6683 (N_6683,N_6412,N_6598);
and U6684 (N_6684,N_6410,N_6425);
or U6685 (N_6685,N_6440,N_6474);
nor U6686 (N_6686,N_6583,N_6580);
and U6687 (N_6687,N_6432,N_6536);
nor U6688 (N_6688,N_6421,N_6426);
or U6689 (N_6689,N_6456,N_6431);
and U6690 (N_6690,N_6417,N_6592);
and U6691 (N_6691,N_6490,N_6576);
nand U6692 (N_6692,N_6413,N_6404);
nand U6693 (N_6693,N_6540,N_6415);
nor U6694 (N_6694,N_6502,N_6451);
or U6695 (N_6695,N_6578,N_6482);
or U6696 (N_6696,N_6575,N_6438);
nor U6697 (N_6697,N_6453,N_6476);
or U6698 (N_6698,N_6480,N_6543);
xnor U6699 (N_6699,N_6584,N_6452);
or U6700 (N_6700,N_6585,N_6574);
nand U6701 (N_6701,N_6596,N_6525);
nand U6702 (N_6702,N_6409,N_6549);
or U6703 (N_6703,N_6445,N_6565);
or U6704 (N_6704,N_6595,N_6565);
nor U6705 (N_6705,N_6559,N_6565);
or U6706 (N_6706,N_6446,N_6535);
xor U6707 (N_6707,N_6592,N_6577);
or U6708 (N_6708,N_6535,N_6441);
xnor U6709 (N_6709,N_6554,N_6499);
nor U6710 (N_6710,N_6448,N_6400);
and U6711 (N_6711,N_6504,N_6537);
xor U6712 (N_6712,N_6543,N_6586);
xnor U6713 (N_6713,N_6521,N_6412);
nor U6714 (N_6714,N_6530,N_6518);
or U6715 (N_6715,N_6550,N_6581);
or U6716 (N_6716,N_6551,N_6410);
or U6717 (N_6717,N_6426,N_6471);
xor U6718 (N_6718,N_6513,N_6484);
and U6719 (N_6719,N_6540,N_6407);
and U6720 (N_6720,N_6409,N_6470);
nand U6721 (N_6721,N_6454,N_6537);
and U6722 (N_6722,N_6489,N_6536);
nand U6723 (N_6723,N_6458,N_6533);
nand U6724 (N_6724,N_6423,N_6474);
nor U6725 (N_6725,N_6507,N_6554);
and U6726 (N_6726,N_6450,N_6594);
nand U6727 (N_6727,N_6593,N_6580);
nor U6728 (N_6728,N_6455,N_6535);
nand U6729 (N_6729,N_6455,N_6544);
or U6730 (N_6730,N_6583,N_6570);
and U6731 (N_6731,N_6433,N_6573);
and U6732 (N_6732,N_6465,N_6536);
and U6733 (N_6733,N_6501,N_6523);
and U6734 (N_6734,N_6406,N_6516);
xnor U6735 (N_6735,N_6592,N_6483);
nand U6736 (N_6736,N_6435,N_6518);
nand U6737 (N_6737,N_6431,N_6599);
nand U6738 (N_6738,N_6472,N_6467);
nand U6739 (N_6739,N_6591,N_6541);
nor U6740 (N_6740,N_6551,N_6477);
or U6741 (N_6741,N_6485,N_6546);
xor U6742 (N_6742,N_6561,N_6453);
and U6743 (N_6743,N_6504,N_6580);
and U6744 (N_6744,N_6489,N_6447);
xnor U6745 (N_6745,N_6541,N_6558);
and U6746 (N_6746,N_6427,N_6567);
nand U6747 (N_6747,N_6520,N_6450);
nand U6748 (N_6748,N_6473,N_6496);
nand U6749 (N_6749,N_6467,N_6524);
nor U6750 (N_6750,N_6467,N_6530);
nand U6751 (N_6751,N_6560,N_6464);
and U6752 (N_6752,N_6458,N_6468);
and U6753 (N_6753,N_6551,N_6476);
and U6754 (N_6754,N_6439,N_6557);
xor U6755 (N_6755,N_6422,N_6464);
or U6756 (N_6756,N_6581,N_6566);
nand U6757 (N_6757,N_6442,N_6426);
nor U6758 (N_6758,N_6444,N_6598);
and U6759 (N_6759,N_6559,N_6576);
or U6760 (N_6760,N_6565,N_6426);
nor U6761 (N_6761,N_6543,N_6513);
or U6762 (N_6762,N_6540,N_6521);
nand U6763 (N_6763,N_6493,N_6522);
xnor U6764 (N_6764,N_6522,N_6412);
nand U6765 (N_6765,N_6543,N_6519);
and U6766 (N_6766,N_6501,N_6545);
or U6767 (N_6767,N_6452,N_6462);
nor U6768 (N_6768,N_6533,N_6593);
or U6769 (N_6769,N_6507,N_6514);
nand U6770 (N_6770,N_6405,N_6429);
or U6771 (N_6771,N_6414,N_6549);
and U6772 (N_6772,N_6526,N_6509);
and U6773 (N_6773,N_6561,N_6582);
or U6774 (N_6774,N_6592,N_6409);
or U6775 (N_6775,N_6463,N_6504);
nand U6776 (N_6776,N_6493,N_6482);
nor U6777 (N_6777,N_6462,N_6456);
nor U6778 (N_6778,N_6590,N_6565);
xnor U6779 (N_6779,N_6580,N_6476);
or U6780 (N_6780,N_6581,N_6565);
or U6781 (N_6781,N_6545,N_6511);
or U6782 (N_6782,N_6415,N_6501);
nand U6783 (N_6783,N_6418,N_6404);
xor U6784 (N_6784,N_6479,N_6524);
xnor U6785 (N_6785,N_6458,N_6400);
and U6786 (N_6786,N_6576,N_6413);
or U6787 (N_6787,N_6552,N_6538);
nor U6788 (N_6788,N_6556,N_6457);
nand U6789 (N_6789,N_6460,N_6476);
nand U6790 (N_6790,N_6493,N_6412);
and U6791 (N_6791,N_6508,N_6411);
nor U6792 (N_6792,N_6599,N_6482);
nor U6793 (N_6793,N_6455,N_6478);
nor U6794 (N_6794,N_6416,N_6538);
nor U6795 (N_6795,N_6518,N_6474);
xor U6796 (N_6796,N_6470,N_6549);
or U6797 (N_6797,N_6520,N_6566);
nor U6798 (N_6798,N_6460,N_6450);
nand U6799 (N_6799,N_6561,N_6480);
or U6800 (N_6800,N_6661,N_6608);
or U6801 (N_6801,N_6733,N_6627);
nand U6802 (N_6802,N_6667,N_6754);
and U6803 (N_6803,N_6629,N_6664);
xnor U6804 (N_6804,N_6726,N_6637);
xor U6805 (N_6805,N_6751,N_6618);
or U6806 (N_6806,N_6706,N_6695);
xnor U6807 (N_6807,N_6756,N_6764);
xor U6808 (N_6808,N_6709,N_6747);
nor U6809 (N_6809,N_6769,N_6630);
xor U6810 (N_6810,N_6788,N_6621);
and U6811 (N_6811,N_6723,N_6654);
and U6812 (N_6812,N_6720,N_6659);
nand U6813 (N_6813,N_6744,N_6643);
xor U6814 (N_6814,N_6644,N_6717);
xnor U6815 (N_6815,N_6741,N_6796);
and U6816 (N_6816,N_6632,N_6722);
xnor U6817 (N_6817,N_6727,N_6694);
xor U6818 (N_6818,N_6680,N_6714);
and U6819 (N_6819,N_6609,N_6776);
or U6820 (N_6820,N_6772,N_6739);
or U6821 (N_6821,N_6790,N_6711);
nand U6822 (N_6822,N_6732,N_6781);
nand U6823 (N_6823,N_6639,N_6755);
nand U6824 (N_6824,N_6686,N_6691);
and U6825 (N_6825,N_6628,N_6604);
xor U6826 (N_6826,N_6652,N_6645);
and U6827 (N_6827,N_6683,N_6716);
nand U6828 (N_6828,N_6619,N_6689);
nor U6829 (N_6829,N_6729,N_6673);
nor U6830 (N_6830,N_6681,N_6672);
nand U6831 (N_6831,N_6740,N_6657);
and U6832 (N_6832,N_6668,N_6771);
nand U6833 (N_6833,N_6633,N_6752);
or U6834 (N_6834,N_6622,N_6669);
xor U6835 (N_6835,N_6782,N_6725);
xnor U6836 (N_6836,N_6762,N_6665);
or U6837 (N_6837,N_6712,N_6617);
nor U6838 (N_6838,N_6784,N_6750);
or U6839 (N_6839,N_6738,N_6647);
xor U6840 (N_6840,N_6786,N_6724);
or U6841 (N_6841,N_6783,N_6703);
nor U6842 (N_6842,N_6611,N_6760);
xor U6843 (N_6843,N_6603,N_6615);
or U6844 (N_6844,N_6670,N_6682);
nand U6845 (N_6845,N_6698,N_6770);
nor U6846 (N_6846,N_6613,N_6692);
and U6847 (N_6847,N_6768,N_6651);
or U6848 (N_6848,N_6702,N_6605);
or U6849 (N_6849,N_6758,N_6777);
or U6850 (N_6850,N_6749,N_6761);
nand U6851 (N_6851,N_6773,N_6614);
or U6852 (N_6852,N_6640,N_6623);
nand U6853 (N_6853,N_6631,N_6798);
or U6854 (N_6854,N_6648,N_6636);
nand U6855 (N_6855,N_6693,N_6678);
and U6856 (N_6856,N_6721,N_6779);
and U6857 (N_6857,N_6757,N_6701);
nand U6858 (N_6858,N_6778,N_6635);
nor U6859 (N_6859,N_6699,N_6616);
xnor U6860 (N_6860,N_6728,N_6697);
nor U6861 (N_6861,N_6660,N_6625);
nor U6862 (N_6862,N_6679,N_6685);
or U6863 (N_6863,N_6704,N_6797);
nor U6864 (N_6864,N_6663,N_6675);
or U6865 (N_6865,N_6734,N_6687);
nor U6866 (N_6866,N_6748,N_6737);
xor U6867 (N_6867,N_6787,N_6650);
xnor U6868 (N_6868,N_6656,N_6601);
and U6869 (N_6869,N_6666,N_6602);
and U6870 (N_6870,N_6634,N_6763);
or U6871 (N_6871,N_6759,N_6774);
and U6872 (N_6872,N_6638,N_6684);
nand U6873 (N_6873,N_6794,N_6612);
nand U6874 (N_6874,N_6658,N_6662);
xnor U6875 (N_6875,N_6655,N_6710);
nor U6876 (N_6876,N_6765,N_6606);
or U6877 (N_6877,N_6696,N_6610);
nor U6878 (N_6878,N_6646,N_6767);
xnor U6879 (N_6879,N_6653,N_6642);
xor U6880 (N_6880,N_6745,N_6719);
nand U6881 (N_6881,N_6793,N_6792);
nand U6882 (N_6882,N_6735,N_6641);
nor U6883 (N_6883,N_6700,N_6775);
or U6884 (N_6884,N_6708,N_6743);
nand U6885 (N_6885,N_6713,N_6746);
nand U6886 (N_6886,N_6707,N_6799);
nor U6887 (N_6887,N_6715,N_6736);
xnor U6888 (N_6888,N_6766,N_6674);
and U6889 (N_6889,N_6785,N_6742);
nor U6890 (N_6890,N_6753,N_6600);
xnor U6891 (N_6891,N_6791,N_6730);
xor U6892 (N_6892,N_6649,N_6690);
nor U6893 (N_6893,N_6620,N_6718);
or U6894 (N_6894,N_6624,N_6607);
or U6895 (N_6895,N_6677,N_6795);
or U6896 (N_6896,N_6676,N_6731);
xor U6897 (N_6897,N_6789,N_6626);
or U6898 (N_6898,N_6705,N_6780);
or U6899 (N_6899,N_6671,N_6688);
nor U6900 (N_6900,N_6780,N_6676);
nor U6901 (N_6901,N_6609,N_6703);
xor U6902 (N_6902,N_6601,N_6630);
nand U6903 (N_6903,N_6734,N_6633);
or U6904 (N_6904,N_6716,N_6709);
nor U6905 (N_6905,N_6796,N_6633);
or U6906 (N_6906,N_6659,N_6676);
xnor U6907 (N_6907,N_6613,N_6767);
nor U6908 (N_6908,N_6634,N_6626);
or U6909 (N_6909,N_6779,N_6745);
or U6910 (N_6910,N_6733,N_6614);
or U6911 (N_6911,N_6721,N_6658);
nor U6912 (N_6912,N_6624,N_6771);
xnor U6913 (N_6913,N_6607,N_6687);
or U6914 (N_6914,N_6703,N_6660);
nand U6915 (N_6915,N_6622,N_6739);
nand U6916 (N_6916,N_6731,N_6775);
xor U6917 (N_6917,N_6654,N_6771);
nor U6918 (N_6918,N_6769,N_6787);
nand U6919 (N_6919,N_6642,N_6624);
nor U6920 (N_6920,N_6669,N_6603);
or U6921 (N_6921,N_6703,N_6687);
nor U6922 (N_6922,N_6627,N_6791);
nand U6923 (N_6923,N_6664,N_6610);
nand U6924 (N_6924,N_6613,N_6779);
nand U6925 (N_6925,N_6680,N_6782);
or U6926 (N_6926,N_6704,N_6765);
nand U6927 (N_6927,N_6646,N_6748);
and U6928 (N_6928,N_6651,N_6621);
nand U6929 (N_6929,N_6740,N_6698);
and U6930 (N_6930,N_6686,N_6722);
nor U6931 (N_6931,N_6762,N_6715);
nand U6932 (N_6932,N_6728,N_6679);
nor U6933 (N_6933,N_6669,N_6765);
xor U6934 (N_6934,N_6779,N_6723);
nand U6935 (N_6935,N_6732,N_6607);
or U6936 (N_6936,N_6619,N_6654);
nor U6937 (N_6937,N_6782,N_6674);
and U6938 (N_6938,N_6742,N_6799);
nand U6939 (N_6939,N_6674,N_6761);
or U6940 (N_6940,N_6643,N_6666);
nor U6941 (N_6941,N_6662,N_6756);
nand U6942 (N_6942,N_6616,N_6656);
nor U6943 (N_6943,N_6632,N_6749);
or U6944 (N_6944,N_6656,N_6681);
nor U6945 (N_6945,N_6795,N_6608);
or U6946 (N_6946,N_6623,N_6689);
and U6947 (N_6947,N_6629,N_6619);
nand U6948 (N_6948,N_6731,N_6689);
xnor U6949 (N_6949,N_6675,N_6741);
and U6950 (N_6950,N_6707,N_6623);
nand U6951 (N_6951,N_6620,N_6794);
or U6952 (N_6952,N_6627,N_6765);
nor U6953 (N_6953,N_6709,N_6641);
nor U6954 (N_6954,N_6746,N_6640);
nor U6955 (N_6955,N_6671,N_6663);
nor U6956 (N_6956,N_6636,N_6791);
xnor U6957 (N_6957,N_6628,N_6639);
nand U6958 (N_6958,N_6706,N_6623);
or U6959 (N_6959,N_6675,N_6769);
nor U6960 (N_6960,N_6665,N_6658);
nor U6961 (N_6961,N_6632,N_6713);
nor U6962 (N_6962,N_6691,N_6649);
nor U6963 (N_6963,N_6632,N_6696);
nor U6964 (N_6964,N_6696,N_6789);
nand U6965 (N_6965,N_6774,N_6739);
nor U6966 (N_6966,N_6778,N_6648);
xor U6967 (N_6967,N_6799,N_6698);
or U6968 (N_6968,N_6788,N_6716);
xor U6969 (N_6969,N_6769,N_6637);
and U6970 (N_6970,N_6643,N_6701);
nand U6971 (N_6971,N_6730,N_6778);
xor U6972 (N_6972,N_6740,N_6601);
nor U6973 (N_6973,N_6717,N_6679);
and U6974 (N_6974,N_6757,N_6687);
or U6975 (N_6975,N_6781,N_6766);
nor U6976 (N_6976,N_6662,N_6717);
and U6977 (N_6977,N_6663,N_6763);
and U6978 (N_6978,N_6625,N_6631);
nand U6979 (N_6979,N_6686,N_6676);
xnor U6980 (N_6980,N_6618,N_6609);
and U6981 (N_6981,N_6603,N_6679);
nor U6982 (N_6982,N_6602,N_6744);
nand U6983 (N_6983,N_6630,N_6600);
or U6984 (N_6984,N_6772,N_6730);
and U6985 (N_6985,N_6643,N_6640);
nand U6986 (N_6986,N_6601,N_6673);
and U6987 (N_6987,N_6662,N_6798);
nor U6988 (N_6988,N_6766,N_6786);
xor U6989 (N_6989,N_6669,N_6790);
nor U6990 (N_6990,N_6620,N_6784);
nor U6991 (N_6991,N_6693,N_6683);
and U6992 (N_6992,N_6746,N_6728);
or U6993 (N_6993,N_6663,N_6783);
xor U6994 (N_6994,N_6763,N_6617);
nand U6995 (N_6995,N_6678,N_6698);
nand U6996 (N_6996,N_6648,N_6661);
xnor U6997 (N_6997,N_6734,N_6721);
xor U6998 (N_6998,N_6651,N_6657);
nand U6999 (N_6999,N_6635,N_6723);
nor U7000 (N_7000,N_6944,N_6843);
nor U7001 (N_7001,N_6979,N_6858);
nand U7002 (N_7002,N_6970,N_6855);
nor U7003 (N_7003,N_6811,N_6960);
nand U7004 (N_7004,N_6930,N_6985);
nand U7005 (N_7005,N_6896,N_6829);
and U7006 (N_7006,N_6969,N_6941);
and U7007 (N_7007,N_6998,N_6994);
nand U7008 (N_7008,N_6816,N_6916);
xnor U7009 (N_7009,N_6844,N_6889);
and U7010 (N_7010,N_6923,N_6906);
xnor U7011 (N_7011,N_6937,N_6929);
and U7012 (N_7012,N_6847,N_6903);
nand U7013 (N_7013,N_6886,N_6950);
nor U7014 (N_7014,N_6962,N_6856);
nand U7015 (N_7015,N_6940,N_6810);
nor U7016 (N_7016,N_6824,N_6907);
nor U7017 (N_7017,N_6832,N_6933);
xnor U7018 (N_7018,N_6943,N_6982);
nor U7019 (N_7019,N_6804,N_6992);
nand U7020 (N_7020,N_6917,N_6865);
nand U7021 (N_7021,N_6851,N_6838);
and U7022 (N_7022,N_6961,N_6915);
nand U7023 (N_7023,N_6890,N_6904);
and U7024 (N_7024,N_6808,N_6883);
xnor U7025 (N_7025,N_6813,N_6828);
and U7026 (N_7026,N_6955,N_6871);
and U7027 (N_7027,N_6836,N_6814);
and U7028 (N_7028,N_6866,N_6964);
and U7029 (N_7029,N_6873,N_6956);
xnor U7030 (N_7030,N_6949,N_6803);
and U7031 (N_7031,N_6875,N_6819);
and U7032 (N_7032,N_6862,N_6909);
nor U7033 (N_7033,N_6809,N_6919);
nor U7034 (N_7034,N_6882,N_6936);
nand U7035 (N_7035,N_6966,N_6869);
nand U7036 (N_7036,N_6820,N_6864);
and U7037 (N_7037,N_6894,N_6993);
xor U7038 (N_7038,N_6876,N_6918);
nand U7039 (N_7039,N_6931,N_6818);
and U7040 (N_7040,N_6958,N_6850);
nor U7041 (N_7041,N_6854,N_6957);
nand U7042 (N_7042,N_6984,N_6912);
or U7043 (N_7043,N_6861,N_6800);
and U7044 (N_7044,N_6852,N_6908);
nand U7045 (N_7045,N_6983,N_6849);
nor U7046 (N_7046,N_6973,N_6892);
nor U7047 (N_7047,N_6833,N_6996);
and U7048 (N_7048,N_6939,N_6948);
nand U7049 (N_7049,N_6951,N_6897);
nand U7050 (N_7050,N_6924,N_6953);
xnor U7051 (N_7051,N_6870,N_6934);
xor U7052 (N_7052,N_6834,N_6860);
nor U7053 (N_7053,N_6830,N_6842);
xor U7054 (N_7054,N_6997,N_6999);
and U7055 (N_7055,N_6990,N_6853);
nor U7056 (N_7056,N_6839,N_6891);
and U7057 (N_7057,N_6900,N_6878);
and U7058 (N_7058,N_6801,N_6802);
nor U7059 (N_7059,N_6926,N_6857);
or U7060 (N_7060,N_6938,N_6974);
nor U7061 (N_7061,N_6986,N_6825);
or U7062 (N_7062,N_6863,N_6885);
and U7063 (N_7063,N_6905,N_6911);
and U7064 (N_7064,N_6965,N_6823);
xor U7065 (N_7065,N_6927,N_6988);
nor U7066 (N_7066,N_6822,N_6935);
xor U7067 (N_7067,N_6976,N_6846);
and U7068 (N_7068,N_6946,N_6848);
and U7069 (N_7069,N_6928,N_6963);
xnor U7070 (N_7070,N_6901,N_6835);
nor U7071 (N_7071,N_6920,N_6805);
xor U7072 (N_7072,N_6975,N_6872);
and U7073 (N_7073,N_6815,N_6902);
or U7074 (N_7074,N_6977,N_6837);
nor U7075 (N_7075,N_6831,N_6995);
nor U7076 (N_7076,N_6913,N_6867);
nor U7077 (N_7077,N_6991,N_6812);
xnor U7078 (N_7078,N_6981,N_6972);
and U7079 (N_7079,N_6922,N_6840);
xnor U7080 (N_7080,N_6968,N_6910);
nor U7081 (N_7081,N_6859,N_6880);
xor U7082 (N_7082,N_6899,N_6868);
or U7083 (N_7083,N_6874,N_6879);
nand U7084 (N_7084,N_6989,N_6893);
xor U7085 (N_7085,N_6932,N_6942);
or U7086 (N_7086,N_6807,N_6959);
nand U7087 (N_7087,N_6952,N_6877);
nand U7088 (N_7088,N_6881,N_6978);
and U7089 (N_7089,N_6826,N_6827);
and U7090 (N_7090,N_6884,N_6925);
xnor U7091 (N_7091,N_6817,N_6841);
nor U7092 (N_7092,N_6887,N_6967);
xnor U7093 (N_7093,N_6914,N_6954);
nor U7094 (N_7094,N_6947,N_6895);
and U7095 (N_7095,N_6971,N_6806);
xnor U7096 (N_7096,N_6888,N_6921);
nand U7097 (N_7097,N_6980,N_6821);
or U7098 (N_7098,N_6945,N_6987);
or U7099 (N_7099,N_6845,N_6898);
nor U7100 (N_7100,N_6902,N_6993);
nand U7101 (N_7101,N_6938,N_6932);
xor U7102 (N_7102,N_6818,N_6949);
nand U7103 (N_7103,N_6835,N_6895);
or U7104 (N_7104,N_6898,N_6813);
nor U7105 (N_7105,N_6945,N_6921);
nand U7106 (N_7106,N_6872,N_6890);
and U7107 (N_7107,N_6842,N_6948);
or U7108 (N_7108,N_6813,N_6971);
nand U7109 (N_7109,N_6872,N_6999);
nand U7110 (N_7110,N_6901,N_6949);
and U7111 (N_7111,N_6861,N_6884);
nand U7112 (N_7112,N_6974,N_6898);
nor U7113 (N_7113,N_6851,N_6806);
xnor U7114 (N_7114,N_6943,N_6814);
nor U7115 (N_7115,N_6972,N_6886);
and U7116 (N_7116,N_6836,N_6847);
xnor U7117 (N_7117,N_6896,N_6960);
nor U7118 (N_7118,N_6875,N_6858);
nand U7119 (N_7119,N_6843,N_6802);
nand U7120 (N_7120,N_6906,N_6874);
nor U7121 (N_7121,N_6872,N_6957);
nand U7122 (N_7122,N_6961,N_6987);
and U7123 (N_7123,N_6867,N_6920);
xor U7124 (N_7124,N_6849,N_6897);
and U7125 (N_7125,N_6863,N_6948);
nor U7126 (N_7126,N_6822,N_6942);
and U7127 (N_7127,N_6982,N_6891);
xor U7128 (N_7128,N_6917,N_6896);
nor U7129 (N_7129,N_6816,N_6882);
nand U7130 (N_7130,N_6909,N_6951);
and U7131 (N_7131,N_6828,N_6891);
nor U7132 (N_7132,N_6836,N_6971);
nand U7133 (N_7133,N_6817,N_6843);
nor U7134 (N_7134,N_6990,N_6960);
nor U7135 (N_7135,N_6931,N_6848);
nand U7136 (N_7136,N_6944,N_6875);
xor U7137 (N_7137,N_6845,N_6865);
nand U7138 (N_7138,N_6910,N_6975);
nor U7139 (N_7139,N_6884,N_6952);
nand U7140 (N_7140,N_6909,N_6807);
and U7141 (N_7141,N_6958,N_6978);
nand U7142 (N_7142,N_6903,N_6826);
nor U7143 (N_7143,N_6912,N_6909);
nand U7144 (N_7144,N_6885,N_6814);
or U7145 (N_7145,N_6953,N_6844);
or U7146 (N_7146,N_6885,N_6963);
or U7147 (N_7147,N_6879,N_6978);
or U7148 (N_7148,N_6988,N_6864);
and U7149 (N_7149,N_6895,N_6898);
nor U7150 (N_7150,N_6839,N_6947);
nor U7151 (N_7151,N_6992,N_6944);
nand U7152 (N_7152,N_6996,N_6811);
nor U7153 (N_7153,N_6987,N_6957);
or U7154 (N_7154,N_6940,N_6843);
and U7155 (N_7155,N_6853,N_6916);
nor U7156 (N_7156,N_6947,N_6890);
nor U7157 (N_7157,N_6830,N_6800);
xnor U7158 (N_7158,N_6823,N_6970);
xor U7159 (N_7159,N_6976,N_6877);
or U7160 (N_7160,N_6995,N_6869);
nor U7161 (N_7161,N_6887,N_6976);
and U7162 (N_7162,N_6866,N_6897);
and U7163 (N_7163,N_6824,N_6848);
or U7164 (N_7164,N_6930,N_6929);
nor U7165 (N_7165,N_6937,N_6868);
nand U7166 (N_7166,N_6902,N_6831);
nor U7167 (N_7167,N_6868,N_6863);
nand U7168 (N_7168,N_6840,N_6857);
or U7169 (N_7169,N_6881,N_6914);
nand U7170 (N_7170,N_6970,N_6990);
and U7171 (N_7171,N_6926,N_6874);
and U7172 (N_7172,N_6897,N_6996);
nand U7173 (N_7173,N_6999,N_6965);
nand U7174 (N_7174,N_6954,N_6863);
and U7175 (N_7175,N_6825,N_6872);
and U7176 (N_7176,N_6806,N_6814);
nor U7177 (N_7177,N_6969,N_6904);
and U7178 (N_7178,N_6861,N_6925);
nor U7179 (N_7179,N_6817,N_6876);
and U7180 (N_7180,N_6899,N_6800);
nor U7181 (N_7181,N_6830,N_6990);
nand U7182 (N_7182,N_6837,N_6934);
nand U7183 (N_7183,N_6853,N_6924);
and U7184 (N_7184,N_6932,N_6909);
nand U7185 (N_7185,N_6918,N_6987);
or U7186 (N_7186,N_6883,N_6868);
and U7187 (N_7187,N_6997,N_6846);
nand U7188 (N_7188,N_6951,N_6858);
and U7189 (N_7189,N_6840,N_6942);
or U7190 (N_7190,N_6802,N_6836);
and U7191 (N_7191,N_6917,N_6991);
or U7192 (N_7192,N_6950,N_6919);
and U7193 (N_7193,N_6981,N_6955);
and U7194 (N_7194,N_6964,N_6862);
nand U7195 (N_7195,N_6981,N_6851);
xor U7196 (N_7196,N_6857,N_6927);
and U7197 (N_7197,N_6937,N_6874);
xor U7198 (N_7198,N_6851,N_6997);
and U7199 (N_7199,N_6943,N_6835);
xor U7200 (N_7200,N_7135,N_7074);
or U7201 (N_7201,N_7073,N_7032);
or U7202 (N_7202,N_7152,N_7124);
and U7203 (N_7203,N_7104,N_7047);
nor U7204 (N_7204,N_7025,N_7099);
xor U7205 (N_7205,N_7151,N_7182);
nor U7206 (N_7206,N_7024,N_7183);
nand U7207 (N_7207,N_7156,N_7103);
nor U7208 (N_7208,N_7089,N_7023);
nor U7209 (N_7209,N_7030,N_7133);
or U7210 (N_7210,N_7038,N_7014);
xor U7211 (N_7211,N_7018,N_7148);
xnor U7212 (N_7212,N_7168,N_7070);
and U7213 (N_7213,N_7029,N_7011);
or U7214 (N_7214,N_7009,N_7082);
nand U7215 (N_7215,N_7096,N_7052);
and U7216 (N_7216,N_7002,N_7054);
or U7217 (N_7217,N_7128,N_7092);
xnor U7218 (N_7218,N_7109,N_7123);
or U7219 (N_7219,N_7193,N_7006);
or U7220 (N_7220,N_7060,N_7196);
nand U7221 (N_7221,N_7134,N_7066);
nand U7222 (N_7222,N_7131,N_7067);
and U7223 (N_7223,N_7107,N_7088);
nand U7224 (N_7224,N_7010,N_7149);
nor U7225 (N_7225,N_7061,N_7116);
nor U7226 (N_7226,N_7186,N_7097);
nor U7227 (N_7227,N_7034,N_7114);
nand U7228 (N_7228,N_7187,N_7055);
xor U7229 (N_7229,N_7068,N_7164);
xnor U7230 (N_7230,N_7085,N_7162);
or U7231 (N_7231,N_7001,N_7053);
and U7232 (N_7232,N_7105,N_7167);
and U7233 (N_7233,N_7174,N_7078);
nor U7234 (N_7234,N_7062,N_7185);
xnor U7235 (N_7235,N_7170,N_7136);
and U7236 (N_7236,N_7019,N_7065);
nor U7237 (N_7237,N_7050,N_7081);
and U7238 (N_7238,N_7080,N_7181);
or U7239 (N_7239,N_7090,N_7084);
and U7240 (N_7240,N_7057,N_7137);
or U7241 (N_7241,N_7138,N_7076);
and U7242 (N_7242,N_7157,N_7100);
and U7243 (N_7243,N_7013,N_7049);
or U7244 (N_7244,N_7111,N_7069);
or U7245 (N_7245,N_7031,N_7027);
or U7246 (N_7246,N_7077,N_7017);
xnor U7247 (N_7247,N_7033,N_7176);
xor U7248 (N_7248,N_7035,N_7072);
and U7249 (N_7249,N_7037,N_7016);
and U7250 (N_7250,N_7122,N_7173);
or U7251 (N_7251,N_7042,N_7110);
nor U7252 (N_7252,N_7003,N_7153);
and U7253 (N_7253,N_7108,N_7101);
xnor U7254 (N_7254,N_7058,N_7087);
nor U7255 (N_7255,N_7071,N_7094);
nor U7256 (N_7256,N_7188,N_7147);
xor U7257 (N_7257,N_7091,N_7194);
nor U7258 (N_7258,N_7045,N_7121);
and U7259 (N_7259,N_7172,N_7175);
nor U7260 (N_7260,N_7159,N_7169);
or U7261 (N_7261,N_7140,N_7117);
nor U7262 (N_7262,N_7075,N_7192);
or U7263 (N_7263,N_7020,N_7040);
xnor U7264 (N_7264,N_7189,N_7007);
nor U7265 (N_7265,N_7043,N_7132);
xor U7266 (N_7266,N_7093,N_7015);
xnor U7267 (N_7267,N_7141,N_7056);
nand U7268 (N_7268,N_7142,N_7028);
nor U7269 (N_7269,N_7163,N_7041);
and U7270 (N_7270,N_7048,N_7130);
and U7271 (N_7271,N_7051,N_7064);
nor U7272 (N_7272,N_7198,N_7171);
nor U7273 (N_7273,N_7086,N_7026);
or U7274 (N_7274,N_7197,N_7102);
or U7275 (N_7275,N_7021,N_7144);
nand U7276 (N_7276,N_7146,N_7005);
and U7277 (N_7277,N_7046,N_7036);
and U7278 (N_7278,N_7044,N_7098);
nand U7279 (N_7279,N_7059,N_7079);
nand U7280 (N_7280,N_7139,N_7115);
nand U7281 (N_7281,N_7083,N_7166);
and U7282 (N_7282,N_7063,N_7195);
nor U7283 (N_7283,N_7154,N_7126);
nor U7284 (N_7284,N_7145,N_7119);
nor U7285 (N_7285,N_7004,N_7129);
nand U7286 (N_7286,N_7118,N_7095);
and U7287 (N_7287,N_7039,N_7177);
or U7288 (N_7288,N_7012,N_7022);
xnor U7289 (N_7289,N_7106,N_7000);
and U7290 (N_7290,N_7184,N_7158);
nand U7291 (N_7291,N_7127,N_7120);
nor U7292 (N_7292,N_7150,N_7180);
or U7293 (N_7293,N_7155,N_7191);
nand U7294 (N_7294,N_7125,N_7199);
nand U7295 (N_7295,N_7113,N_7008);
nor U7296 (N_7296,N_7112,N_7165);
xnor U7297 (N_7297,N_7161,N_7143);
nand U7298 (N_7298,N_7190,N_7178);
xnor U7299 (N_7299,N_7160,N_7179);
and U7300 (N_7300,N_7175,N_7059);
xnor U7301 (N_7301,N_7067,N_7070);
or U7302 (N_7302,N_7037,N_7106);
or U7303 (N_7303,N_7114,N_7177);
xnor U7304 (N_7304,N_7158,N_7020);
nor U7305 (N_7305,N_7087,N_7121);
or U7306 (N_7306,N_7064,N_7122);
nand U7307 (N_7307,N_7080,N_7100);
xor U7308 (N_7308,N_7024,N_7009);
and U7309 (N_7309,N_7092,N_7165);
nand U7310 (N_7310,N_7182,N_7053);
or U7311 (N_7311,N_7066,N_7065);
nor U7312 (N_7312,N_7111,N_7120);
nand U7313 (N_7313,N_7147,N_7137);
xor U7314 (N_7314,N_7014,N_7065);
nor U7315 (N_7315,N_7101,N_7045);
and U7316 (N_7316,N_7024,N_7102);
nor U7317 (N_7317,N_7165,N_7091);
xnor U7318 (N_7318,N_7042,N_7195);
or U7319 (N_7319,N_7164,N_7085);
or U7320 (N_7320,N_7047,N_7186);
xor U7321 (N_7321,N_7180,N_7132);
xor U7322 (N_7322,N_7137,N_7020);
nand U7323 (N_7323,N_7150,N_7101);
or U7324 (N_7324,N_7185,N_7136);
xor U7325 (N_7325,N_7103,N_7066);
and U7326 (N_7326,N_7164,N_7095);
and U7327 (N_7327,N_7058,N_7091);
and U7328 (N_7328,N_7005,N_7007);
nor U7329 (N_7329,N_7103,N_7150);
xor U7330 (N_7330,N_7109,N_7096);
xnor U7331 (N_7331,N_7123,N_7077);
nand U7332 (N_7332,N_7106,N_7048);
and U7333 (N_7333,N_7007,N_7081);
nand U7334 (N_7334,N_7189,N_7008);
xnor U7335 (N_7335,N_7111,N_7139);
xor U7336 (N_7336,N_7182,N_7146);
xor U7337 (N_7337,N_7088,N_7069);
xor U7338 (N_7338,N_7083,N_7061);
and U7339 (N_7339,N_7103,N_7170);
and U7340 (N_7340,N_7067,N_7119);
nor U7341 (N_7341,N_7139,N_7037);
nor U7342 (N_7342,N_7012,N_7133);
nor U7343 (N_7343,N_7060,N_7057);
xnor U7344 (N_7344,N_7081,N_7047);
xor U7345 (N_7345,N_7064,N_7159);
nor U7346 (N_7346,N_7185,N_7039);
nand U7347 (N_7347,N_7197,N_7170);
nand U7348 (N_7348,N_7062,N_7159);
or U7349 (N_7349,N_7171,N_7133);
nand U7350 (N_7350,N_7015,N_7162);
or U7351 (N_7351,N_7093,N_7170);
xor U7352 (N_7352,N_7146,N_7095);
nand U7353 (N_7353,N_7035,N_7065);
nor U7354 (N_7354,N_7189,N_7126);
and U7355 (N_7355,N_7130,N_7014);
xnor U7356 (N_7356,N_7095,N_7153);
or U7357 (N_7357,N_7172,N_7113);
and U7358 (N_7358,N_7157,N_7046);
nand U7359 (N_7359,N_7104,N_7141);
and U7360 (N_7360,N_7098,N_7126);
xor U7361 (N_7361,N_7104,N_7149);
nor U7362 (N_7362,N_7119,N_7054);
nor U7363 (N_7363,N_7119,N_7125);
xor U7364 (N_7364,N_7173,N_7176);
nor U7365 (N_7365,N_7079,N_7176);
or U7366 (N_7366,N_7030,N_7080);
or U7367 (N_7367,N_7056,N_7083);
xnor U7368 (N_7368,N_7196,N_7125);
nand U7369 (N_7369,N_7001,N_7032);
and U7370 (N_7370,N_7117,N_7118);
or U7371 (N_7371,N_7170,N_7148);
nor U7372 (N_7372,N_7040,N_7019);
nor U7373 (N_7373,N_7055,N_7075);
nor U7374 (N_7374,N_7147,N_7013);
xnor U7375 (N_7375,N_7158,N_7035);
nand U7376 (N_7376,N_7039,N_7053);
nor U7377 (N_7377,N_7072,N_7173);
nor U7378 (N_7378,N_7033,N_7137);
nor U7379 (N_7379,N_7177,N_7144);
nand U7380 (N_7380,N_7139,N_7152);
or U7381 (N_7381,N_7125,N_7034);
xor U7382 (N_7382,N_7005,N_7045);
xor U7383 (N_7383,N_7086,N_7153);
nand U7384 (N_7384,N_7010,N_7033);
and U7385 (N_7385,N_7095,N_7189);
or U7386 (N_7386,N_7101,N_7151);
and U7387 (N_7387,N_7046,N_7165);
and U7388 (N_7388,N_7014,N_7028);
nand U7389 (N_7389,N_7103,N_7076);
nand U7390 (N_7390,N_7005,N_7163);
xor U7391 (N_7391,N_7005,N_7001);
or U7392 (N_7392,N_7047,N_7100);
nand U7393 (N_7393,N_7156,N_7147);
nand U7394 (N_7394,N_7048,N_7175);
nand U7395 (N_7395,N_7197,N_7049);
nor U7396 (N_7396,N_7096,N_7139);
and U7397 (N_7397,N_7040,N_7083);
and U7398 (N_7398,N_7104,N_7014);
nand U7399 (N_7399,N_7066,N_7048);
and U7400 (N_7400,N_7221,N_7235);
nand U7401 (N_7401,N_7383,N_7294);
and U7402 (N_7402,N_7303,N_7355);
and U7403 (N_7403,N_7397,N_7232);
xnor U7404 (N_7404,N_7217,N_7359);
and U7405 (N_7405,N_7352,N_7348);
nor U7406 (N_7406,N_7277,N_7317);
xor U7407 (N_7407,N_7305,N_7373);
nand U7408 (N_7408,N_7205,N_7256);
xor U7409 (N_7409,N_7349,N_7295);
or U7410 (N_7410,N_7372,N_7275);
or U7411 (N_7411,N_7318,N_7357);
or U7412 (N_7412,N_7356,N_7395);
nand U7413 (N_7413,N_7308,N_7274);
nand U7414 (N_7414,N_7262,N_7310);
xnor U7415 (N_7415,N_7398,N_7371);
or U7416 (N_7416,N_7381,N_7346);
xor U7417 (N_7417,N_7269,N_7396);
nand U7418 (N_7418,N_7242,N_7370);
and U7419 (N_7419,N_7273,N_7286);
nand U7420 (N_7420,N_7204,N_7234);
and U7421 (N_7421,N_7288,N_7211);
or U7422 (N_7422,N_7306,N_7216);
nand U7423 (N_7423,N_7347,N_7284);
nand U7424 (N_7424,N_7362,N_7343);
xnor U7425 (N_7425,N_7309,N_7297);
nor U7426 (N_7426,N_7272,N_7394);
or U7427 (N_7427,N_7330,N_7248);
xnor U7428 (N_7428,N_7313,N_7307);
nand U7429 (N_7429,N_7293,N_7287);
nor U7430 (N_7430,N_7257,N_7241);
nand U7431 (N_7431,N_7292,N_7304);
and U7432 (N_7432,N_7333,N_7227);
nor U7433 (N_7433,N_7378,N_7276);
nand U7434 (N_7434,N_7223,N_7249);
nand U7435 (N_7435,N_7326,N_7264);
nor U7436 (N_7436,N_7393,N_7354);
nand U7437 (N_7437,N_7368,N_7200);
and U7438 (N_7438,N_7229,N_7341);
xnor U7439 (N_7439,N_7238,N_7351);
xnor U7440 (N_7440,N_7376,N_7328);
xor U7441 (N_7441,N_7283,N_7331);
and U7442 (N_7442,N_7375,N_7296);
or U7443 (N_7443,N_7327,N_7209);
or U7444 (N_7444,N_7360,N_7246);
and U7445 (N_7445,N_7300,N_7301);
and U7446 (N_7446,N_7334,N_7207);
xor U7447 (N_7447,N_7374,N_7320);
and U7448 (N_7448,N_7335,N_7332);
xor U7449 (N_7449,N_7243,N_7261);
xor U7450 (N_7450,N_7312,N_7202);
nand U7451 (N_7451,N_7392,N_7298);
and U7452 (N_7452,N_7319,N_7278);
or U7453 (N_7453,N_7263,N_7377);
and U7454 (N_7454,N_7338,N_7218);
nor U7455 (N_7455,N_7206,N_7281);
and U7456 (N_7456,N_7363,N_7389);
nand U7457 (N_7457,N_7228,N_7361);
nor U7458 (N_7458,N_7390,N_7266);
nor U7459 (N_7459,N_7350,N_7254);
or U7460 (N_7460,N_7358,N_7267);
nand U7461 (N_7461,N_7280,N_7255);
nand U7462 (N_7462,N_7231,N_7384);
nor U7463 (N_7463,N_7322,N_7399);
nand U7464 (N_7464,N_7299,N_7220);
or U7465 (N_7465,N_7265,N_7302);
xor U7466 (N_7466,N_7289,N_7282);
nor U7467 (N_7467,N_7285,N_7208);
xor U7468 (N_7468,N_7279,N_7260);
or U7469 (N_7469,N_7244,N_7239);
xnor U7470 (N_7470,N_7215,N_7224);
nand U7471 (N_7471,N_7268,N_7240);
nor U7472 (N_7472,N_7236,N_7291);
nand U7473 (N_7473,N_7323,N_7271);
xor U7474 (N_7474,N_7344,N_7290);
nor U7475 (N_7475,N_7380,N_7201);
xnor U7476 (N_7476,N_7245,N_7367);
nand U7477 (N_7477,N_7382,N_7219);
nor U7478 (N_7478,N_7315,N_7250);
nand U7479 (N_7479,N_7270,N_7364);
nor U7480 (N_7480,N_7339,N_7316);
and U7481 (N_7481,N_7337,N_7222);
nand U7482 (N_7482,N_7252,N_7247);
or U7483 (N_7483,N_7251,N_7336);
or U7484 (N_7484,N_7225,N_7226);
or U7485 (N_7485,N_7237,N_7366);
and U7486 (N_7486,N_7387,N_7388);
nor U7487 (N_7487,N_7324,N_7353);
and U7488 (N_7488,N_7379,N_7391);
and U7489 (N_7489,N_7314,N_7325);
nor U7490 (N_7490,N_7214,N_7210);
xnor U7491 (N_7491,N_7345,N_7365);
or U7492 (N_7492,N_7258,N_7385);
xnor U7493 (N_7493,N_7340,N_7212);
nand U7494 (N_7494,N_7329,N_7369);
nor U7495 (N_7495,N_7203,N_7386);
nand U7496 (N_7496,N_7321,N_7311);
xor U7497 (N_7497,N_7342,N_7213);
xor U7498 (N_7498,N_7253,N_7230);
nor U7499 (N_7499,N_7233,N_7259);
nand U7500 (N_7500,N_7387,N_7275);
and U7501 (N_7501,N_7390,N_7220);
or U7502 (N_7502,N_7377,N_7311);
or U7503 (N_7503,N_7372,N_7340);
nor U7504 (N_7504,N_7338,N_7287);
nor U7505 (N_7505,N_7347,N_7346);
or U7506 (N_7506,N_7270,N_7331);
xnor U7507 (N_7507,N_7223,N_7254);
and U7508 (N_7508,N_7318,N_7208);
nor U7509 (N_7509,N_7298,N_7256);
or U7510 (N_7510,N_7379,N_7208);
nand U7511 (N_7511,N_7297,N_7247);
nor U7512 (N_7512,N_7366,N_7316);
or U7513 (N_7513,N_7377,N_7391);
or U7514 (N_7514,N_7343,N_7303);
nand U7515 (N_7515,N_7375,N_7261);
nor U7516 (N_7516,N_7246,N_7261);
and U7517 (N_7517,N_7241,N_7288);
xnor U7518 (N_7518,N_7332,N_7222);
xnor U7519 (N_7519,N_7377,N_7362);
nand U7520 (N_7520,N_7324,N_7317);
nand U7521 (N_7521,N_7205,N_7239);
and U7522 (N_7522,N_7368,N_7335);
xor U7523 (N_7523,N_7248,N_7280);
and U7524 (N_7524,N_7214,N_7249);
xnor U7525 (N_7525,N_7303,N_7329);
nand U7526 (N_7526,N_7276,N_7256);
or U7527 (N_7527,N_7259,N_7271);
nor U7528 (N_7528,N_7311,N_7364);
nand U7529 (N_7529,N_7345,N_7232);
nand U7530 (N_7530,N_7315,N_7345);
nand U7531 (N_7531,N_7313,N_7373);
and U7532 (N_7532,N_7248,N_7325);
xnor U7533 (N_7533,N_7275,N_7360);
and U7534 (N_7534,N_7303,N_7398);
nand U7535 (N_7535,N_7370,N_7339);
or U7536 (N_7536,N_7353,N_7289);
or U7537 (N_7537,N_7385,N_7214);
and U7538 (N_7538,N_7276,N_7236);
nor U7539 (N_7539,N_7392,N_7387);
nand U7540 (N_7540,N_7349,N_7300);
and U7541 (N_7541,N_7304,N_7243);
nor U7542 (N_7542,N_7286,N_7224);
xor U7543 (N_7543,N_7278,N_7357);
xnor U7544 (N_7544,N_7299,N_7296);
nand U7545 (N_7545,N_7291,N_7213);
and U7546 (N_7546,N_7215,N_7333);
xor U7547 (N_7547,N_7273,N_7330);
nand U7548 (N_7548,N_7293,N_7220);
xnor U7549 (N_7549,N_7201,N_7291);
nor U7550 (N_7550,N_7352,N_7223);
xnor U7551 (N_7551,N_7264,N_7353);
and U7552 (N_7552,N_7322,N_7200);
nor U7553 (N_7553,N_7378,N_7212);
nor U7554 (N_7554,N_7250,N_7221);
and U7555 (N_7555,N_7268,N_7211);
xor U7556 (N_7556,N_7357,N_7343);
nor U7557 (N_7557,N_7278,N_7314);
nor U7558 (N_7558,N_7279,N_7234);
and U7559 (N_7559,N_7231,N_7367);
and U7560 (N_7560,N_7220,N_7356);
or U7561 (N_7561,N_7217,N_7372);
xnor U7562 (N_7562,N_7393,N_7209);
nand U7563 (N_7563,N_7283,N_7394);
xnor U7564 (N_7564,N_7203,N_7245);
or U7565 (N_7565,N_7375,N_7226);
xor U7566 (N_7566,N_7335,N_7205);
and U7567 (N_7567,N_7233,N_7246);
xor U7568 (N_7568,N_7214,N_7200);
or U7569 (N_7569,N_7297,N_7277);
nand U7570 (N_7570,N_7349,N_7253);
nand U7571 (N_7571,N_7384,N_7292);
nor U7572 (N_7572,N_7250,N_7283);
nand U7573 (N_7573,N_7209,N_7304);
or U7574 (N_7574,N_7263,N_7367);
and U7575 (N_7575,N_7325,N_7378);
or U7576 (N_7576,N_7269,N_7354);
and U7577 (N_7577,N_7367,N_7323);
and U7578 (N_7578,N_7200,N_7356);
or U7579 (N_7579,N_7366,N_7240);
or U7580 (N_7580,N_7367,N_7307);
and U7581 (N_7581,N_7377,N_7249);
and U7582 (N_7582,N_7304,N_7342);
xor U7583 (N_7583,N_7272,N_7254);
nand U7584 (N_7584,N_7389,N_7335);
xnor U7585 (N_7585,N_7395,N_7324);
and U7586 (N_7586,N_7362,N_7221);
and U7587 (N_7587,N_7216,N_7282);
or U7588 (N_7588,N_7204,N_7351);
or U7589 (N_7589,N_7331,N_7290);
nand U7590 (N_7590,N_7245,N_7332);
or U7591 (N_7591,N_7291,N_7396);
or U7592 (N_7592,N_7206,N_7353);
xor U7593 (N_7593,N_7248,N_7372);
xor U7594 (N_7594,N_7245,N_7339);
and U7595 (N_7595,N_7322,N_7211);
and U7596 (N_7596,N_7249,N_7317);
xnor U7597 (N_7597,N_7213,N_7318);
nand U7598 (N_7598,N_7367,N_7246);
nor U7599 (N_7599,N_7307,N_7249);
xnor U7600 (N_7600,N_7432,N_7496);
nand U7601 (N_7601,N_7504,N_7499);
nor U7602 (N_7602,N_7588,N_7541);
xnor U7603 (N_7603,N_7539,N_7484);
nand U7604 (N_7604,N_7520,N_7551);
or U7605 (N_7605,N_7509,N_7597);
xor U7606 (N_7606,N_7571,N_7569);
or U7607 (N_7607,N_7452,N_7595);
xnor U7608 (N_7608,N_7489,N_7456);
xnor U7609 (N_7609,N_7559,N_7493);
or U7610 (N_7610,N_7421,N_7556);
nand U7611 (N_7611,N_7529,N_7408);
xor U7612 (N_7612,N_7563,N_7587);
and U7613 (N_7613,N_7464,N_7513);
xor U7614 (N_7614,N_7526,N_7430);
or U7615 (N_7615,N_7424,N_7583);
and U7616 (N_7616,N_7417,N_7445);
nor U7617 (N_7617,N_7514,N_7572);
or U7618 (N_7618,N_7593,N_7468);
and U7619 (N_7619,N_7470,N_7429);
nor U7620 (N_7620,N_7506,N_7462);
and U7621 (N_7621,N_7522,N_7411);
nor U7622 (N_7622,N_7546,N_7535);
xnor U7623 (N_7623,N_7442,N_7431);
or U7624 (N_7624,N_7540,N_7533);
or U7625 (N_7625,N_7441,N_7550);
xnor U7626 (N_7626,N_7423,N_7498);
nor U7627 (N_7627,N_7422,N_7425);
nand U7628 (N_7628,N_7419,N_7573);
nor U7629 (N_7629,N_7538,N_7492);
or U7630 (N_7630,N_7549,N_7501);
nor U7631 (N_7631,N_7505,N_7534);
or U7632 (N_7632,N_7508,N_7525);
nor U7633 (N_7633,N_7443,N_7400);
or U7634 (N_7634,N_7524,N_7457);
nand U7635 (N_7635,N_7482,N_7448);
and U7636 (N_7636,N_7580,N_7471);
or U7637 (N_7637,N_7519,N_7568);
nand U7638 (N_7638,N_7469,N_7491);
or U7639 (N_7639,N_7455,N_7490);
nand U7640 (N_7640,N_7502,N_7545);
nand U7641 (N_7641,N_7548,N_7420);
and U7642 (N_7642,N_7585,N_7570);
or U7643 (N_7643,N_7599,N_7437);
nor U7644 (N_7644,N_7507,N_7454);
nor U7645 (N_7645,N_7497,N_7561);
xor U7646 (N_7646,N_7584,N_7465);
or U7647 (N_7647,N_7521,N_7510);
nand U7648 (N_7648,N_7512,N_7594);
nand U7649 (N_7649,N_7434,N_7516);
or U7650 (N_7650,N_7591,N_7449);
or U7651 (N_7651,N_7460,N_7574);
xnor U7652 (N_7652,N_7447,N_7418);
xnor U7653 (N_7653,N_7494,N_7495);
xnor U7654 (N_7654,N_7586,N_7481);
nand U7655 (N_7655,N_7415,N_7477);
and U7656 (N_7656,N_7433,N_7459);
nor U7657 (N_7657,N_7589,N_7557);
xnor U7658 (N_7658,N_7410,N_7527);
nand U7659 (N_7659,N_7552,N_7426);
xor U7660 (N_7660,N_7518,N_7560);
or U7661 (N_7661,N_7414,N_7537);
and U7662 (N_7662,N_7466,N_7436);
xnor U7663 (N_7663,N_7467,N_7547);
and U7664 (N_7664,N_7439,N_7473);
xor U7665 (N_7665,N_7566,N_7528);
and U7666 (N_7666,N_7554,N_7590);
xor U7667 (N_7667,N_7413,N_7485);
xnor U7668 (N_7668,N_7567,N_7401);
and U7669 (N_7669,N_7412,N_7487);
nor U7670 (N_7670,N_7444,N_7479);
or U7671 (N_7671,N_7403,N_7446);
nor U7672 (N_7672,N_7438,N_7451);
or U7673 (N_7673,N_7543,N_7577);
xor U7674 (N_7674,N_7517,N_7483);
nor U7675 (N_7675,N_7582,N_7402);
xnor U7676 (N_7676,N_7486,N_7503);
or U7677 (N_7677,N_7564,N_7428);
and U7678 (N_7678,N_7435,N_7592);
nor U7679 (N_7679,N_7536,N_7450);
nor U7680 (N_7680,N_7515,N_7596);
xor U7681 (N_7681,N_7579,N_7531);
nor U7682 (N_7682,N_7461,N_7475);
xor U7683 (N_7683,N_7530,N_7578);
nor U7684 (N_7684,N_7565,N_7480);
xor U7685 (N_7685,N_7488,N_7405);
and U7686 (N_7686,N_7532,N_7463);
or U7687 (N_7687,N_7558,N_7511);
nor U7688 (N_7688,N_7500,N_7404);
or U7689 (N_7689,N_7553,N_7542);
xnor U7690 (N_7690,N_7555,N_7409);
xor U7691 (N_7691,N_7416,N_7523);
and U7692 (N_7692,N_7544,N_7562);
and U7693 (N_7693,N_7458,N_7581);
xor U7694 (N_7694,N_7427,N_7440);
and U7695 (N_7695,N_7476,N_7575);
and U7696 (N_7696,N_7453,N_7407);
nand U7697 (N_7697,N_7598,N_7474);
nor U7698 (N_7698,N_7478,N_7576);
nand U7699 (N_7699,N_7406,N_7472);
and U7700 (N_7700,N_7446,N_7489);
nand U7701 (N_7701,N_7569,N_7576);
and U7702 (N_7702,N_7525,N_7521);
xnor U7703 (N_7703,N_7559,N_7567);
and U7704 (N_7704,N_7487,N_7491);
nand U7705 (N_7705,N_7474,N_7488);
or U7706 (N_7706,N_7568,N_7433);
xor U7707 (N_7707,N_7435,N_7474);
or U7708 (N_7708,N_7511,N_7451);
or U7709 (N_7709,N_7512,N_7437);
nand U7710 (N_7710,N_7426,N_7575);
xor U7711 (N_7711,N_7540,N_7400);
xnor U7712 (N_7712,N_7461,N_7413);
nand U7713 (N_7713,N_7488,N_7548);
xor U7714 (N_7714,N_7495,N_7530);
or U7715 (N_7715,N_7510,N_7523);
or U7716 (N_7716,N_7459,N_7536);
or U7717 (N_7717,N_7443,N_7484);
xor U7718 (N_7718,N_7553,N_7567);
nor U7719 (N_7719,N_7403,N_7420);
nand U7720 (N_7720,N_7456,N_7588);
and U7721 (N_7721,N_7500,N_7561);
xnor U7722 (N_7722,N_7429,N_7478);
nor U7723 (N_7723,N_7466,N_7523);
nor U7724 (N_7724,N_7592,N_7579);
nand U7725 (N_7725,N_7598,N_7402);
xor U7726 (N_7726,N_7515,N_7542);
nor U7727 (N_7727,N_7462,N_7508);
nor U7728 (N_7728,N_7423,N_7543);
xnor U7729 (N_7729,N_7540,N_7403);
nor U7730 (N_7730,N_7470,N_7549);
and U7731 (N_7731,N_7535,N_7490);
xor U7732 (N_7732,N_7516,N_7530);
and U7733 (N_7733,N_7559,N_7507);
nor U7734 (N_7734,N_7522,N_7405);
nor U7735 (N_7735,N_7492,N_7406);
or U7736 (N_7736,N_7467,N_7561);
nand U7737 (N_7737,N_7576,N_7587);
nand U7738 (N_7738,N_7551,N_7569);
xnor U7739 (N_7739,N_7437,N_7483);
xor U7740 (N_7740,N_7444,N_7554);
and U7741 (N_7741,N_7535,N_7552);
xor U7742 (N_7742,N_7499,N_7469);
nor U7743 (N_7743,N_7554,N_7526);
or U7744 (N_7744,N_7523,N_7595);
and U7745 (N_7745,N_7469,N_7517);
nor U7746 (N_7746,N_7406,N_7518);
nand U7747 (N_7747,N_7580,N_7538);
or U7748 (N_7748,N_7569,N_7493);
xnor U7749 (N_7749,N_7529,N_7487);
or U7750 (N_7750,N_7450,N_7427);
or U7751 (N_7751,N_7507,N_7442);
xor U7752 (N_7752,N_7412,N_7443);
xnor U7753 (N_7753,N_7443,N_7545);
xor U7754 (N_7754,N_7492,N_7467);
or U7755 (N_7755,N_7559,N_7479);
xnor U7756 (N_7756,N_7423,N_7474);
nand U7757 (N_7757,N_7472,N_7403);
nand U7758 (N_7758,N_7577,N_7593);
xor U7759 (N_7759,N_7543,N_7572);
nor U7760 (N_7760,N_7590,N_7557);
nor U7761 (N_7761,N_7518,N_7548);
or U7762 (N_7762,N_7454,N_7550);
xnor U7763 (N_7763,N_7592,N_7469);
or U7764 (N_7764,N_7580,N_7478);
nor U7765 (N_7765,N_7538,N_7577);
xnor U7766 (N_7766,N_7532,N_7510);
nor U7767 (N_7767,N_7437,N_7404);
xor U7768 (N_7768,N_7477,N_7454);
nand U7769 (N_7769,N_7560,N_7509);
and U7770 (N_7770,N_7496,N_7486);
or U7771 (N_7771,N_7589,N_7418);
nor U7772 (N_7772,N_7535,N_7520);
nor U7773 (N_7773,N_7417,N_7588);
or U7774 (N_7774,N_7467,N_7504);
xnor U7775 (N_7775,N_7509,N_7491);
nor U7776 (N_7776,N_7526,N_7543);
nand U7777 (N_7777,N_7451,N_7483);
or U7778 (N_7778,N_7423,N_7590);
and U7779 (N_7779,N_7569,N_7505);
nand U7780 (N_7780,N_7503,N_7408);
and U7781 (N_7781,N_7422,N_7473);
xor U7782 (N_7782,N_7468,N_7565);
or U7783 (N_7783,N_7413,N_7513);
nor U7784 (N_7784,N_7412,N_7561);
nor U7785 (N_7785,N_7496,N_7421);
or U7786 (N_7786,N_7483,N_7495);
xnor U7787 (N_7787,N_7524,N_7423);
xor U7788 (N_7788,N_7508,N_7532);
and U7789 (N_7789,N_7447,N_7505);
xnor U7790 (N_7790,N_7417,N_7414);
xor U7791 (N_7791,N_7490,N_7443);
and U7792 (N_7792,N_7483,N_7477);
nor U7793 (N_7793,N_7404,N_7487);
nor U7794 (N_7794,N_7575,N_7464);
nand U7795 (N_7795,N_7455,N_7492);
and U7796 (N_7796,N_7548,N_7494);
and U7797 (N_7797,N_7523,N_7501);
xnor U7798 (N_7798,N_7409,N_7468);
and U7799 (N_7799,N_7425,N_7458);
nor U7800 (N_7800,N_7670,N_7600);
or U7801 (N_7801,N_7698,N_7758);
nor U7802 (N_7802,N_7784,N_7781);
xnor U7803 (N_7803,N_7696,N_7796);
nor U7804 (N_7804,N_7793,N_7773);
and U7805 (N_7805,N_7635,N_7638);
and U7806 (N_7806,N_7734,N_7690);
xor U7807 (N_7807,N_7684,N_7617);
or U7808 (N_7808,N_7632,N_7641);
and U7809 (N_7809,N_7707,N_7752);
xor U7810 (N_7810,N_7790,N_7779);
and U7811 (N_7811,N_7627,N_7605);
nand U7812 (N_7812,N_7644,N_7611);
or U7813 (N_7813,N_7675,N_7765);
or U7814 (N_7814,N_7626,N_7689);
nor U7815 (N_7815,N_7722,N_7649);
and U7816 (N_7816,N_7747,N_7667);
xnor U7817 (N_7817,N_7629,N_7685);
and U7818 (N_7818,N_7705,N_7770);
nand U7819 (N_7819,N_7709,N_7662);
and U7820 (N_7820,N_7769,N_7609);
or U7821 (N_7821,N_7672,N_7652);
and U7822 (N_7822,N_7625,N_7688);
xor U7823 (N_7823,N_7787,N_7761);
or U7824 (N_7824,N_7785,N_7701);
or U7825 (N_7825,N_7634,N_7703);
or U7826 (N_7826,N_7633,N_7771);
nor U7827 (N_7827,N_7648,N_7735);
or U7828 (N_7828,N_7711,N_7687);
nand U7829 (N_7829,N_7668,N_7748);
nor U7830 (N_7830,N_7733,N_7608);
or U7831 (N_7831,N_7620,N_7673);
and U7832 (N_7832,N_7653,N_7724);
or U7833 (N_7833,N_7789,N_7622);
nand U7834 (N_7834,N_7727,N_7739);
xnor U7835 (N_7835,N_7694,N_7794);
xnor U7836 (N_7836,N_7767,N_7618);
xnor U7837 (N_7837,N_7657,N_7725);
nor U7838 (N_7838,N_7777,N_7732);
or U7839 (N_7839,N_7660,N_7683);
nor U7840 (N_7840,N_7716,N_7655);
or U7841 (N_7841,N_7762,N_7750);
nand U7842 (N_7842,N_7702,N_7776);
nand U7843 (N_7843,N_7754,N_7603);
nand U7844 (N_7844,N_7792,N_7745);
nor U7845 (N_7845,N_7678,N_7602);
or U7846 (N_7846,N_7676,N_7743);
and U7847 (N_7847,N_7778,N_7719);
nor U7848 (N_7848,N_7640,N_7788);
or U7849 (N_7849,N_7606,N_7646);
or U7850 (N_7850,N_7636,N_7738);
and U7851 (N_7851,N_7797,N_7729);
xor U7852 (N_7852,N_7666,N_7749);
nand U7853 (N_7853,N_7669,N_7686);
or U7854 (N_7854,N_7766,N_7615);
nor U7855 (N_7855,N_7621,N_7737);
nor U7856 (N_7856,N_7730,N_7714);
and U7857 (N_7857,N_7616,N_7717);
nand U7858 (N_7858,N_7751,N_7718);
and U7859 (N_7859,N_7713,N_7623);
nand U7860 (N_7860,N_7708,N_7742);
nand U7861 (N_7861,N_7680,N_7613);
xnor U7862 (N_7862,N_7682,N_7741);
nand U7863 (N_7863,N_7775,N_7723);
nor U7864 (N_7864,N_7783,N_7628);
or U7865 (N_7865,N_7647,N_7643);
nand U7866 (N_7866,N_7757,N_7755);
or U7867 (N_7867,N_7658,N_7674);
and U7868 (N_7868,N_7607,N_7665);
xnor U7869 (N_7869,N_7610,N_7721);
xnor U7870 (N_7870,N_7726,N_7782);
and U7871 (N_7871,N_7661,N_7759);
nor U7872 (N_7872,N_7645,N_7706);
or U7873 (N_7873,N_7699,N_7756);
nor U7874 (N_7874,N_7798,N_7677);
xnor U7875 (N_7875,N_7692,N_7601);
nand U7876 (N_7876,N_7671,N_7760);
xnor U7877 (N_7877,N_7799,N_7651);
nor U7878 (N_7878,N_7619,N_7780);
xnor U7879 (N_7879,N_7630,N_7720);
and U7880 (N_7880,N_7728,N_7614);
nor U7881 (N_7881,N_7740,N_7681);
xor U7882 (N_7882,N_7763,N_7786);
nor U7883 (N_7883,N_7791,N_7637);
and U7884 (N_7884,N_7679,N_7774);
or U7885 (N_7885,N_7704,N_7631);
and U7886 (N_7886,N_7659,N_7715);
nor U7887 (N_7887,N_7712,N_7656);
nand U7888 (N_7888,N_7693,N_7795);
xnor U7889 (N_7889,N_7664,N_7710);
or U7890 (N_7890,N_7663,N_7642);
nor U7891 (N_7891,N_7731,N_7744);
or U7892 (N_7892,N_7654,N_7746);
nand U7893 (N_7893,N_7639,N_7697);
nor U7894 (N_7894,N_7772,N_7700);
and U7895 (N_7895,N_7753,N_7624);
nor U7896 (N_7896,N_7764,N_7612);
and U7897 (N_7897,N_7691,N_7695);
nor U7898 (N_7898,N_7650,N_7768);
xnor U7899 (N_7899,N_7736,N_7604);
or U7900 (N_7900,N_7748,N_7652);
nand U7901 (N_7901,N_7630,N_7743);
and U7902 (N_7902,N_7782,N_7707);
xnor U7903 (N_7903,N_7712,N_7757);
or U7904 (N_7904,N_7714,N_7614);
or U7905 (N_7905,N_7750,N_7773);
nor U7906 (N_7906,N_7723,N_7650);
xor U7907 (N_7907,N_7744,N_7724);
nor U7908 (N_7908,N_7724,N_7730);
and U7909 (N_7909,N_7734,N_7669);
nor U7910 (N_7910,N_7771,N_7610);
nand U7911 (N_7911,N_7638,N_7636);
or U7912 (N_7912,N_7667,N_7602);
and U7913 (N_7913,N_7731,N_7728);
and U7914 (N_7914,N_7618,N_7775);
nand U7915 (N_7915,N_7604,N_7648);
nor U7916 (N_7916,N_7670,N_7662);
or U7917 (N_7917,N_7645,N_7757);
or U7918 (N_7918,N_7652,N_7701);
and U7919 (N_7919,N_7733,N_7780);
xnor U7920 (N_7920,N_7678,N_7677);
xnor U7921 (N_7921,N_7696,N_7664);
nor U7922 (N_7922,N_7718,N_7710);
or U7923 (N_7923,N_7679,N_7786);
nand U7924 (N_7924,N_7759,N_7726);
xor U7925 (N_7925,N_7609,N_7652);
and U7926 (N_7926,N_7645,N_7686);
nand U7927 (N_7927,N_7752,N_7781);
and U7928 (N_7928,N_7622,N_7763);
nor U7929 (N_7929,N_7650,N_7678);
nand U7930 (N_7930,N_7635,N_7758);
nor U7931 (N_7931,N_7785,N_7657);
and U7932 (N_7932,N_7727,N_7704);
nor U7933 (N_7933,N_7724,N_7742);
nand U7934 (N_7934,N_7655,N_7772);
nor U7935 (N_7935,N_7647,N_7661);
xor U7936 (N_7936,N_7761,N_7665);
nor U7937 (N_7937,N_7674,N_7651);
nor U7938 (N_7938,N_7764,N_7791);
nor U7939 (N_7939,N_7714,N_7652);
nor U7940 (N_7940,N_7673,N_7635);
xor U7941 (N_7941,N_7776,N_7679);
xnor U7942 (N_7942,N_7710,N_7769);
nand U7943 (N_7943,N_7700,N_7645);
xor U7944 (N_7944,N_7735,N_7633);
xnor U7945 (N_7945,N_7727,N_7606);
nand U7946 (N_7946,N_7685,N_7650);
nand U7947 (N_7947,N_7636,N_7715);
xor U7948 (N_7948,N_7747,N_7746);
nor U7949 (N_7949,N_7776,N_7735);
nor U7950 (N_7950,N_7740,N_7743);
nand U7951 (N_7951,N_7684,N_7716);
xor U7952 (N_7952,N_7646,N_7726);
nand U7953 (N_7953,N_7666,N_7637);
nor U7954 (N_7954,N_7795,N_7729);
or U7955 (N_7955,N_7741,N_7773);
nor U7956 (N_7956,N_7648,N_7736);
nor U7957 (N_7957,N_7610,N_7664);
nand U7958 (N_7958,N_7688,N_7780);
nand U7959 (N_7959,N_7794,N_7772);
or U7960 (N_7960,N_7782,N_7614);
nand U7961 (N_7961,N_7680,N_7717);
nand U7962 (N_7962,N_7752,N_7632);
nor U7963 (N_7963,N_7725,N_7749);
nor U7964 (N_7964,N_7613,N_7715);
nand U7965 (N_7965,N_7738,N_7681);
and U7966 (N_7966,N_7721,N_7685);
nor U7967 (N_7967,N_7785,N_7781);
and U7968 (N_7968,N_7765,N_7707);
xor U7969 (N_7969,N_7763,N_7628);
and U7970 (N_7970,N_7676,N_7686);
and U7971 (N_7971,N_7679,N_7754);
nand U7972 (N_7972,N_7688,N_7719);
nand U7973 (N_7973,N_7719,N_7756);
nand U7974 (N_7974,N_7788,N_7744);
xor U7975 (N_7975,N_7701,N_7628);
nand U7976 (N_7976,N_7616,N_7688);
and U7977 (N_7977,N_7730,N_7773);
or U7978 (N_7978,N_7776,N_7653);
nand U7979 (N_7979,N_7656,N_7745);
nand U7980 (N_7980,N_7653,N_7684);
xnor U7981 (N_7981,N_7799,N_7797);
and U7982 (N_7982,N_7631,N_7772);
nand U7983 (N_7983,N_7784,N_7762);
or U7984 (N_7984,N_7793,N_7700);
xor U7985 (N_7985,N_7664,N_7604);
and U7986 (N_7986,N_7751,N_7764);
xnor U7987 (N_7987,N_7788,N_7677);
nor U7988 (N_7988,N_7696,N_7605);
xnor U7989 (N_7989,N_7613,N_7706);
or U7990 (N_7990,N_7663,N_7788);
nor U7991 (N_7991,N_7612,N_7603);
nand U7992 (N_7992,N_7767,N_7729);
nand U7993 (N_7993,N_7623,N_7790);
nor U7994 (N_7994,N_7772,N_7691);
nor U7995 (N_7995,N_7698,N_7680);
nand U7996 (N_7996,N_7673,N_7657);
xor U7997 (N_7997,N_7762,N_7748);
xnor U7998 (N_7998,N_7706,N_7786);
or U7999 (N_7999,N_7736,N_7666);
or U8000 (N_8000,N_7990,N_7866);
nor U8001 (N_8001,N_7842,N_7983);
xor U8002 (N_8002,N_7836,N_7854);
and U8003 (N_8003,N_7903,N_7997);
and U8004 (N_8004,N_7880,N_7814);
nor U8005 (N_8005,N_7909,N_7907);
and U8006 (N_8006,N_7930,N_7887);
xor U8007 (N_8007,N_7897,N_7989);
nor U8008 (N_8008,N_7871,N_7980);
nor U8009 (N_8009,N_7899,N_7927);
and U8010 (N_8010,N_7925,N_7968);
xnor U8011 (N_8011,N_7803,N_7827);
xor U8012 (N_8012,N_7815,N_7920);
xnor U8013 (N_8013,N_7935,N_7851);
nand U8014 (N_8014,N_7853,N_7807);
or U8015 (N_8015,N_7912,N_7900);
or U8016 (N_8016,N_7921,N_7963);
xnor U8017 (N_8017,N_7894,N_7808);
or U8018 (N_8018,N_7870,N_7933);
nand U8019 (N_8019,N_7860,N_7949);
nor U8020 (N_8020,N_7821,N_7872);
nand U8021 (N_8021,N_7800,N_7916);
or U8022 (N_8022,N_7878,N_7959);
nor U8023 (N_8023,N_7883,N_7896);
nand U8024 (N_8024,N_7868,N_7859);
xnor U8025 (N_8025,N_7943,N_7919);
nor U8026 (N_8026,N_7984,N_7809);
and U8027 (N_8027,N_7946,N_7975);
and U8028 (N_8028,N_7951,N_7802);
xnor U8029 (N_8029,N_7857,N_7955);
or U8030 (N_8030,N_7826,N_7822);
xor U8031 (N_8031,N_7960,N_7956);
nand U8032 (N_8032,N_7941,N_7844);
nand U8033 (N_8033,N_7901,N_7986);
nor U8034 (N_8034,N_7938,N_7879);
nand U8035 (N_8035,N_7995,N_7806);
and U8036 (N_8036,N_7936,N_7974);
nand U8037 (N_8037,N_7873,N_7819);
xnor U8038 (N_8038,N_7876,N_7944);
xnor U8039 (N_8039,N_7817,N_7856);
xor U8040 (N_8040,N_7987,N_7863);
xor U8041 (N_8041,N_7978,N_7877);
or U8042 (N_8042,N_7805,N_7843);
nand U8043 (N_8043,N_7926,N_7874);
xor U8044 (N_8044,N_7906,N_7966);
and U8045 (N_8045,N_7824,N_7939);
nor U8046 (N_8046,N_7838,N_7950);
and U8047 (N_8047,N_7964,N_7917);
or U8048 (N_8048,N_7829,N_7841);
nand U8049 (N_8049,N_7910,N_7839);
or U8050 (N_8050,N_7820,N_7845);
or U8051 (N_8051,N_7840,N_7848);
xnor U8052 (N_8052,N_7849,N_7888);
or U8053 (N_8053,N_7985,N_7816);
nand U8054 (N_8054,N_7923,N_7837);
nand U8055 (N_8055,N_7818,N_7847);
nor U8056 (N_8056,N_7971,N_7831);
nand U8057 (N_8057,N_7981,N_7922);
nor U8058 (N_8058,N_7858,N_7988);
nand U8059 (N_8059,N_7893,N_7890);
and U8060 (N_8060,N_7813,N_7965);
nand U8061 (N_8061,N_7828,N_7957);
nor U8062 (N_8062,N_7993,N_7958);
nand U8063 (N_8063,N_7929,N_7905);
or U8064 (N_8064,N_7823,N_7867);
and U8065 (N_8065,N_7865,N_7942);
and U8066 (N_8066,N_7810,N_7996);
or U8067 (N_8067,N_7846,N_7931);
nand U8068 (N_8068,N_7886,N_7928);
xor U8069 (N_8069,N_7885,N_7947);
nand U8070 (N_8070,N_7972,N_7913);
xnor U8071 (N_8071,N_7908,N_7861);
xnor U8072 (N_8072,N_7804,N_7855);
nand U8073 (N_8073,N_7898,N_7869);
and U8074 (N_8074,N_7895,N_7862);
and U8075 (N_8075,N_7875,N_7991);
nor U8076 (N_8076,N_7832,N_7911);
nand U8077 (N_8077,N_7934,N_7999);
nand U8078 (N_8078,N_7992,N_7850);
or U8079 (N_8079,N_7882,N_7970);
nor U8080 (N_8080,N_7924,N_7953);
and U8081 (N_8081,N_7998,N_7967);
xor U8082 (N_8082,N_7940,N_7945);
and U8083 (N_8083,N_7852,N_7948);
nor U8084 (N_8084,N_7973,N_7918);
nor U8085 (N_8085,N_7915,N_7889);
xnor U8086 (N_8086,N_7932,N_7891);
or U8087 (N_8087,N_7977,N_7801);
nand U8088 (N_8088,N_7834,N_7962);
and U8089 (N_8089,N_7835,N_7954);
and U8090 (N_8090,N_7937,N_7830);
nand U8091 (N_8091,N_7969,N_7952);
nor U8092 (N_8092,N_7904,N_7812);
or U8093 (N_8093,N_7994,N_7982);
or U8094 (N_8094,N_7892,N_7811);
and U8095 (N_8095,N_7881,N_7825);
xor U8096 (N_8096,N_7902,N_7833);
nand U8097 (N_8097,N_7864,N_7961);
and U8098 (N_8098,N_7979,N_7976);
nor U8099 (N_8099,N_7914,N_7884);
nand U8100 (N_8100,N_7989,N_7894);
and U8101 (N_8101,N_7855,N_7991);
nor U8102 (N_8102,N_7933,N_7982);
xnor U8103 (N_8103,N_7829,N_7819);
xor U8104 (N_8104,N_7904,N_7991);
and U8105 (N_8105,N_7898,N_7879);
nor U8106 (N_8106,N_7839,N_7929);
and U8107 (N_8107,N_7849,N_7944);
nor U8108 (N_8108,N_7846,N_7935);
and U8109 (N_8109,N_7887,N_7859);
xnor U8110 (N_8110,N_7997,N_7963);
nor U8111 (N_8111,N_7906,N_7848);
nor U8112 (N_8112,N_7808,N_7812);
nor U8113 (N_8113,N_7910,N_7865);
and U8114 (N_8114,N_7993,N_7808);
or U8115 (N_8115,N_7936,N_7922);
nor U8116 (N_8116,N_7937,N_7940);
and U8117 (N_8117,N_7862,N_7807);
xor U8118 (N_8118,N_7829,N_7854);
and U8119 (N_8119,N_7843,N_7811);
and U8120 (N_8120,N_7860,N_7832);
and U8121 (N_8121,N_7943,N_7847);
xor U8122 (N_8122,N_7905,N_7955);
and U8123 (N_8123,N_7846,N_7940);
nand U8124 (N_8124,N_7870,N_7974);
nand U8125 (N_8125,N_7861,N_7895);
nand U8126 (N_8126,N_7990,N_7900);
nor U8127 (N_8127,N_7824,N_7960);
nand U8128 (N_8128,N_7900,N_7949);
nor U8129 (N_8129,N_7930,N_7812);
nor U8130 (N_8130,N_7838,N_7929);
nor U8131 (N_8131,N_7916,N_7860);
xnor U8132 (N_8132,N_7886,N_7840);
xor U8133 (N_8133,N_7962,N_7938);
nand U8134 (N_8134,N_7903,N_7868);
nand U8135 (N_8135,N_7943,N_7897);
xnor U8136 (N_8136,N_7868,N_7930);
nor U8137 (N_8137,N_7976,N_7918);
nand U8138 (N_8138,N_7914,N_7962);
or U8139 (N_8139,N_7990,N_7813);
or U8140 (N_8140,N_7803,N_7992);
nor U8141 (N_8141,N_7856,N_7833);
xnor U8142 (N_8142,N_7910,N_7987);
and U8143 (N_8143,N_7997,N_7821);
xnor U8144 (N_8144,N_7828,N_7849);
nor U8145 (N_8145,N_7913,N_7958);
nor U8146 (N_8146,N_7941,N_7952);
or U8147 (N_8147,N_7964,N_7867);
xor U8148 (N_8148,N_7989,N_7979);
or U8149 (N_8149,N_7939,N_7806);
nand U8150 (N_8150,N_7839,N_7987);
nand U8151 (N_8151,N_7935,N_7830);
nand U8152 (N_8152,N_7952,N_7990);
and U8153 (N_8153,N_7960,N_7937);
xnor U8154 (N_8154,N_7820,N_7976);
and U8155 (N_8155,N_7874,N_7921);
or U8156 (N_8156,N_7865,N_7871);
nor U8157 (N_8157,N_7911,N_7803);
and U8158 (N_8158,N_7914,N_7851);
xnor U8159 (N_8159,N_7887,N_7839);
and U8160 (N_8160,N_7867,N_7932);
xor U8161 (N_8161,N_7984,N_7805);
nor U8162 (N_8162,N_7932,N_7879);
or U8163 (N_8163,N_7890,N_7899);
nand U8164 (N_8164,N_7904,N_7871);
and U8165 (N_8165,N_7978,N_7913);
nor U8166 (N_8166,N_7952,N_7870);
and U8167 (N_8167,N_7990,N_7829);
and U8168 (N_8168,N_7960,N_7931);
and U8169 (N_8169,N_7896,N_7920);
or U8170 (N_8170,N_7845,N_7949);
or U8171 (N_8171,N_7969,N_7922);
nand U8172 (N_8172,N_7975,N_7951);
xor U8173 (N_8173,N_7871,N_7959);
and U8174 (N_8174,N_7890,N_7905);
and U8175 (N_8175,N_7859,N_7831);
and U8176 (N_8176,N_7962,N_7835);
nor U8177 (N_8177,N_7852,N_7879);
nor U8178 (N_8178,N_7951,N_7906);
and U8179 (N_8179,N_7810,N_7938);
or U8180 (N_8180,N_7856,N_7881);
xor U8181 (N_8181,N_7997,N_7934);
nand U8182 (N_8182,N_7985,N_7972);
nand U8183 (N_8183,N_7891,N_7881);
nor U8184 (N_8184,N_7900,N_7807);
or U8185 (N_8185,N_7921,N_7808);
or U8186 (N_8186,N_7960,N_7996);
and U8187 (N_8187,N_7897,N_7828);
nor U8188 (N_8188,N_7807,N_7941);
nand U8189 (N_8189,N_7937,N_7870);
or U8190 (N_8190,N_7951,N_7851);
xnor U8191 (N_8191,N_7932,N_7875);
nor U8192 (N_8192,N_7883,N_7922);
nand U8193 (N_8193,N_7893,N_7995);
nor U8194 (N_8194,N_7945,N_7924);
nor U8195 (N_8195,N_7944,N_7992);
and U8196 (N_8196,N_7859,N_7923);
or U8197 (N_8197,N_7916,N_7977);
xor U8198 (N_8198,N_7926,N_7803);
xnor U8199 (N_8199,N_7849,N_7979);
or U8200 (N_8200,N_8114,N_8052);
nor U8201 (N_8201,N_8037,N_8175);
xnor U8202 (N_8202,N_8156,N_8002);
xnor U8203 (N_8203,N_8011,N_8196);
nor U8204 (N_8204,N_8091,N_8053);
xor U8205 (N_8205,N_8050,N_8061);
or U8206 (N_8206,N_8044,N_8104);
or U8207 (N_8207,N_8157,N_8000);
nand U8208 (N_8208,N_8151,N_8186);
nor U8209 (N_8209,N_8164,N_8135);
nor U8210 (N_8210,N_8194,N_8064);
and U8211 (N_8211,N_8159,N_8008);
and U8212 (N_8212,N_8132,N_8129);
nor U8213 (N_8213,N_8118,N_8025);
or U8214 (N_8214,N_8088,N_8145);
nand U8215 (N_8215,N_8069,N_8169);
xor U8216 (N_8216,N_8067,N_8084);
or U8217 (N_8217,N_8060,N_8009);
nand U8218 (N_8218,N_8144,N_8099);
and U8219 (N_8219,N_8184,N_8040);
nand U8220 (N_8220,N_8036,N_8139);
nor U8221 (N_8221,N_8134,N_8119);
nor U8222 (N_8222,N_8172,N_8005);
nor U8223 (N_8223,N_8142,N_8120);
nand U8224 (N_8224,N_8078,N_8199);
or U8225 (N_8225,N_8116,N_8162);
xnor U8226 (N_8226,N_8133,N_8087);
nand U8227 (N_8227,N_8038,N_8013);
nand U8228 (N_8228,N_8131,N_8115);
nor U8229 (N_8229,N_8148,N_8046);
or U8230 (N_8230,N_8062,N_8123);
xnor U8231 (N_8231,N_8063,N_8168);
nor U8232 (N_8232,N_8143,N_8049);
or U8233 (N_8233,N_8066,N_8072);
nor U8234 (N_8234,N_8020,N_8090);
or U8235 (N_8235,N_8146,N_8039);
and U8236 (N_8236,N_8147,N_8018);
or U8237 (N_8237,N_8071,N_8101);
xnor U8238 (N_8238,N_8163,N_8195);
and U8239 (N_8239,N_8180,N_8103);
xnor U8240 (N_8240,N_8010,N_8034);
or U8241 (N_8241,N_8054,N_8045);
and U8242 (N_8242,N_8117,N_8198);
xnor U8243 (N_8243,N_8181,N_8153);
and U8244 (N_8244,N_8140,N_8155);
nor U8245 (N_8245,N_8122,N_8188);
or U8246 (N_8246,N_8176,N_8001);
or U8247 (N_8247,N_8055,N_8125);
xor U8248 (N_8248,N_8003,N_8007);
nand U8249 (N_8249,N_8185,N_8160);
and U8250 (N_8250,N_8017,N_8097);
xor U8251 (N_8251,N_8189,N_8056);
xnor U8252 (N_8252,N_8109,N_8089);
xnor U8253 (N_8253,N_8086,N_8124);
xor U8254 (N_8254,N_8048,N_8150);
xor U8255 (N_8255,N_8057,N_8179);
nor U8256 (N_8256,N_8076,N_8149);
xor U8257 (N_8257,N_8178,N_8107);
or U8258 (N_8258,N_8065,N_8126);
or U8259 (N_8259,N_8127,N_8158);
xor U8260 (N_8260,N_8190,N_8141);
or U8261 (N_8261,N_8079,N_8080);
xnor U8262 (N_8262,N_8170,N_8033);
nand U8263 (N_8263,N_8043,N_8058);
nor U8264 (N_8264,N_8183,N_8171);
nor U8265 (N_8265,N_8022,N_8081);
nand U8266 (N_8266,N_8083,N_8095);
xor U8267 (N_8267,N_8192,N_8024);
nand U8268 (N_8268,N_8173,N_8014);
nand U8269 (N_8269,N_8138,N_8073);
or U8270 (N_8270,N_8004,N_8051);
and U8271 (N_8271,N_8047,N_8074);
nor U8272 (N_8272,N_8077,N_8102);
xnor U8273 (N_8273,N_8012,N_8113);
xor U8274 (N_8274,N_8137,N_8085);
nor U8275 (N_8275,N_8177,N_8030);
nand U8276 (N_8276,N_8059,N_8015);
nand U8277 (N_8277,N_8174,N_8021);
nand U8278 (N_8278,N_8075,N_8092);
and U8279 (N_8279,N_8098,N_8197);
or U8280 (N_8280,N_8032,N_8093);
xor U8281 (N_8281,N_8019,N_8110);
and U8282 (N_8282,N_8121,N_8035);
xnor U8283 (N_8283,N_8128,N_8130);
or U8284 (N_8284,N_8136,N_8031);
xor U8285 (N_8285,N_8027,N_8152);
and U8286 (N_8286,N_8154,N_8006);
and U8287 (N_8287,N_8068,N_8112);
xor U8288 (N_8288,N_8029,N_8165);
and U8289 (N_8289,N_8191,N_8193);
xnor U8290 (N_8290,N_8182,N_8100);
and U8291 (N_8291,N_8042,N_8028);
nor U8292 (N_8292,N_8106,N_8041);
or U8293 (N_8293,N_8070,N_8096);
nor U8294 (N_8294,N_8108,N_8105);
and U8295 (N_8295,N_8167,N_8016);
or U8296 (N_8296,N_8161,N_8111);
xor U8297 (N_8297,N_8023,N_8187);
or U8298 (N_8298,N_8082,N_8094);
nand U8299 (N_8299,N_8026,N_8166);
nor U8300 (N_8300,N_8114,N_8127);
and U8301 (N_8301,N_8101,N_8103);
or U8302 (N_8302,N_8020,N_8131);
or U8303 (N_8303,N_8085,N_8022);
xnor U8304 (N_8304,N_8015,N_8179);
or U8305 (N_8305,N_8177,N_8183);
nand U8306 (N_8306,N_8056,N_8047);
or U8307 (N_8307,N_8017,N_8023);
or U8308 (N_8308,N_8008,N_8078);
or U8309 (N_8309,N_8152,N_8173);
or U8310 (N_8310,N_8083,N_8157);
and U8311 (N_8311,N_8122,N_8059);
nor U8312 (N_8312,N_8187,N_8002);
or U8313 (N_8313,N_8094,N_8104);
nor U8314 (N_8314,N_8146,N_8144);
nor U8315 (N_8315,N_8185,N_8129);
and U8316 (N_8316,N_8037,N_8192);
xor U8317 (N_8317,N_8054,N_8196);
nor U8318 (N_8318,N_8051,N_8197);
nor U8319 (N_8319,N_8012,N_8184);
nor U8320 (N_8320,N_8129,N_8164);
xnor U8321 (N_8321,N_8097,N_8198);
or U8322 (N_8322,N_8158,N_8095);
xor U8323 (N_8323,N_8017,N_8138);
nand U8324 (N_8324,N_8165,N_8116);
nor U8325 (N_8325,N_8129,N_8045);
and U8326 (N_8326,N_8166,N_8169);
or U8327 (N_8327,N_8080,N_8159);
xnor U8328 (N_8328,N_8176,N_8156);
xnor U8329 (N_8329,N_8023,N_8068);
xnor U8330 (N_8330,N_8082,N_8178);
xnor U8331 (N_8331,N_8042,N_8199);
nand U8332 (N_8332,N_8077,N_8054);
and U8333 (N_8333,N_8138,N_8015);
and U8334 (N_8334,N_8142,N_8140);
nand U8335 (N_8335,N_8156,N_8102);
xor U8336 (N_8336,N_8176,N_8190);
nand U8337 (N_8337,N_8136,N_8078);
xor U8338 (N_8338,N_8190,N_8057);
nand U8339 (N_8339,N_8099,N_8102);
xnor U8340 (N_8340,N_8139,N_8021);
nor U8341 (N_8341,N_8104,N_8010);
and U8342 (N_8342,N_8174,N_8009);
and U8343 (N_8343,N_8176,N_8076);
and U8344 (N_8344,N_8030,N_8025);
nor U8345 (N_8345,N_8013,N_8095);
nor U8346 (N_8346,N_8017,N_8074);
nand U8347 (N_8347,N_8078,N_8037);
nor U8348 (N_8348,N_8160,N_8046);
nand U8349 (N_8349,N_8155,N_8104);
nand U8350 (N_8350,N_8187,N_8005);
nand U8351 (N_8351,N_8151,N_8104);
nor U8352 (N_8352,N_8034,N_8043);
nand U8353 (N_8353,N_8060,N_8045);
xor U8354 (N_8354,N_8111,N_8072);
and U8355 (N_8355,N_8012,N_8001);
nor U8356 (N_8356,N_8048,N_8056);
xnor U8357 (N_8357,N_8147,N_8055);
and U8358 (N_8358,N_8043,N_8188);
xnor U8359 (N_8359,N_8192,N_8187);
xnor U8360 (N_8360,N_8060,N_8007);
or U8361 (N_8361,N_8197,N_8007);
nor U8362 (N_8362,N_8158,N_8103);
nand U8363 (N_8363,N_8187,N_8176);
or U8364 (N_8364,N_8132,N_8133);
xor U8365 (N_8365,N_8077,N_8160);
nor U8366 (N_8366,N_8086,N_8067);
nor U8367 (N_8367,N_8002,N_8136);
nand U8368 (N_8368,N_8052,N_8021);
xor U8369 (N_8369,N_8073,N_8035);
nand U8370 (N_8370,N_8008,N_8031);
or U8371 (N_8371,N_8197,N_8086);
nor U8372 (N_8372,N_8087,N_8100);
nor U8373 (N_8373,N_8005,N_8122);
and U8374 (N_8374,N_8111,N_8074);
and U8375 (N_8375,N_8000,N_8190);
or U8376 (N_8376,N_8133,N_8131);
nor U8377 (N_8377,N_8104,N_8084);
or U8378 (N_8378,N_8147,N_8006);
xor U8379 (N_8379,N_8128,N_8015);
nand U8380 (N_8380,N_8024,N_8106);
and U8381 (N_8381,N_8114,N_8065);
nand U8382 (N_8382,N_8194,N_8193);
nor U8383 (N_8383,N_8081,N_8192);
xnor U8384 (N_8384,N_8084,N_8106);
nor U8385 (N_8385,N_8066,N_8165);
nor U8386 (N_8386,N_8097,N_8152);
xor U8387 (N_8387,N_8024,N_8023);
and U8388 (N_8388,N_8148,N_8158);
or U8389 (N_8389,N_8193,N_8105);
xnor U8390 (N_8390,N_8077,N_8185);
nand U8391 (N_8391,N_8075,N_8045);
and U8392 (N_8392,N_8121,N_8094);
or U8393 (N_8393,N_8114,N_8137);
xor U8394 (N_8394,N_8049,N_8039);
xor U8395 (N_8395,N_8154,N_8059);
or U8396 (N_8396,N_8030,N_8150);
nor U8397 (N_8397,N_8011,N_8143);
nor U8398 (N_8398,N_8182,N_8139);
or U8399 (N_8399,N_8022,N_8062);
nand U8400 (N_8400,N_8264,N_8345);
nor U8401 (N_8401,N_8392,N_8250);
nor U8402 (N_8402,N_8332,N_8339);
nand U8403 (N_8403,N_8260,N_8299);
nand U8404 (N_8404,N_8362,N_8388);
xnor U8405 (N_8405,N_8301,N_8204);
nor U8406 (N_8406,N_8237,N_8317);
xnor U8407 (N_8407,N_8391,N_8273);
nor U8408 (N_8408,N_8266,N_8303);
and U8409 (N_8409,N_8398,N_8351);
xnor U8410 (N_8410,N_8342,N_8312);
nand U8411 (N_8411,N_8349,N_8220);
xor U8412 (N_8412,N_8360,N_8319);
xor U8413 (N_8413,N_8336,N_8385);
or U8414 (N_8414,N_8308,N_8348);
xor U8415 (N_8415,N_8207,N_8363);
xnor U8416 (N_8416,N_8283,N_8328);
xor U8417 (N_8417,N_8245,N_8272);
or U8418 (N_8418,N_8321,N_8395);
and U8419 (N_8419,N_8233,N_8213);
nand U8420 (N_8420,N_8252,N_8274);
nor U8421 (N_8421,N_8277,N_8282);
xnor U8422 (N_8422,N_8209,N_8218);
nand U8423 (N_8423,N_8353,N_8370);
or U8424 (N_8424,N_8227,N_8307);
nor U8425 (N_8425,N_8287,N_8323);
nand U8426 (N_8426,N_8367,N_8206);
nor U8427 (N_8427,N_8275,N_8344);
xnor U8428 (N_8428,N_8366,N_8211);
and U8429 (N_8429,N_8201,N_8270);
xor U8430 (N_8430,N_8341,N_8311);
and U8431 (N_8431,N_8340,N_8390);
nor U8432 (N_8432,N_8239,N_8280);
xor U8433 (N_8433,N_8259,N_8249);
nor U8434 (N_8434,N_8399,N_8210);
nor U8435 (N_8435,N_8276,N_8315);
or U8436 (N_8436,N_8373,N_8305);
or U8437 (N_8437,N_8347,N_8352);
and U8438 (N_8438,N_8372,N_8318);
or U8439 (N_8439,N_8313,N_8236);
nand U8440 (N_8440,N_8295,N_8286);
nor U8441 (N_8441,N_8267,N_8258);
nor U8442 (N_8442,N_8214,N_8224);
nor U8443 (N_8443,N_8288,N_8394);
and U8444 (N_8444,N_8350,N_8205);
nor U8445 (N_8445,N_8256,N_8316);
or U8446 (N_8446,N_8310,N_8242);
or U8447 (N_8447,N_8383,N_8369);
nor U8448 (N_8448,N_8247,N_8330);
nand U8449 (N_8449,N_8225,N_8263);
nand U8450 (N_8450,N_8231,N_8281);
and U8451 (N_8451,N_8298,N_8331);
xnor U8452 (N_8452,N_8386,N_8255);
or U8453 (N_8453,N_8229,N_8377);
and U8454 (N_8454,N_8324,N_8300);
nand U8455 (N_8455,N_8269,N_8235);
or U8456 (N_8456,N_8384,N_8257);
nand U8457 (N_8457,N_8254,N_8382);
nor U8458 (N_8458,N_8243,N_8346);
or U8459 (N_8459,N_8238,N_8361);
or U8460 (N_8460,N_8304,N_8234);
or U8461 (N_8461,N_8291,N_8320);
xnor U8462 (N_8462,N_8396,N_8327);
and U8463 (N_8463,N_8221,N_8248);
nor U8464 (N_8464,N_8240,N_8358);
xnor U8465 (N_8465,N_8359,N_8379);
nand U8466 (N_8466,N_8329,N_8357);
or U8467 (N_8467,N_8226,N_8334);
and U8468 (N_8468,N_8293,N_8222);
or U8469 (N_8469,N_8326,N_8387);
xnor U8470 (N_8470,N_8380,N_8355);
nor U8471 (N_8471,N_8228,N_8376);
nand U8472 (N_8472,N_8217,N_8306);
or U8473 (N_8473,N_8325,N_8381);
nand U8474 (N_8474,N_8261,N_8268);
xnor U8475 (N_8475,N_8314,N_8297);
nand U8476 (N_8476,N_8200,N_8230);
nor U8477 (N_8477,N_8309,N_8393);
or U8478 (N_8478,N_8338,N_8368);
xnor U8479 (N_8479,N_8364,N_8262);
and U8480 (N_8480,N_8223,N_8253);
nor U8481 (N_8481,N_8333,N_8292);
xor U8482 (N_8482,N_8271,N_8212);
xnor U8483 (N_8483,N_8215,N_8251);
nor U8484 (N_8484,N_8374,N_8335);
nand U8485 (N_8485,N_8208,N_8289);
nor U8486 (N_8486,N_8265,N_8343);
nand U8487 (N_8487,N_8375,N_8216);
nor U8488 (N_8488,N_8290,N_8244);
nor U8489 (N_8489,N_8219,N_8397);
or U8490 (N_8490,N_8356,N_8284);
xor U8491 (N_8491,N_8322,N_8202);
nand U8492 (N_8492,N_8294,N_8285);
or U8493 (N_8493,N_8378,N_8241);
or U8494 (N_8494,N_8389,N_8278);
nor U8495 (N_8495,N_8203,N_8371);
nand U8496 (N_8496,N_8302,N_8296);
or U8497 (N_8497,N_8365,N_8279);
xnor U8498 (N_8498,N_8246,N_8354);
nand U8499 (N_8499,N_8337,N_8232);
nand U8500 (N_8500,N_8328,N_8315);
xnor U8501 (N_8501,N_8297,N_8352);
xor U8502 (N_8502,N_8250,N_8328);
nor U8503 (N_8503,N_8251,N_8212);
nand U8504 (N_8504,N_8375,N_8236);
nand U8505 (N_8505,N_8282,N_8341);
nand U8506 (N_8506,N_8326,N_8213);
and U8507 (N_8507,N_8250,N_8398);
xor U8508 (N_8508,N_8251,N_8384);
or U8509 (N_8509,N_8351,N_8306);
or U8510 (N_8510,N_8377,N_8305);
and U8511 (N_8511,N_8372,N_8216);
nor U8512 (N_8512,N_8279,N_8235);
nand U8513 (N_8513,N_8317,N_8273);
xor U8514 (N_8514,N_8282,N_8252);
nand U8515 (N_8515,N_8258,N_8200);
or U8516 (N_8516,N_8395,N_8349);
nand U8517 (N_8517,N_8269,N_8264);
or U8518 (N_8518,N_8222,N_8381);
xor U8519 (N_8519,N_8367,N_8374);
xor U8520 (N_8520,N_8284,N_8281);
xor U8521 (N_8521,N_8236,N_8365);
xor U8522 (N_8522,N_8228,N_8254);
nor U8523 (N_8523,N_8336,N_8375);
or U8524 (N_8524,N_8272,N_8354);
nor U8525 (N_8525,N_8384,N_8367);
and U8526 (N_8526,N_8294,N_8251);
nor U8527 (N_8527,N_8357,N_8380);
and U8528 (N_8528,N_8208,N_8281);
nand U8529 (N_8529,N_8225,N_8371);
xnor U8530 (N_8530,N_8260,N_8311);
nor U8531 (N_8531,N_8249,N_8281);
nand U8532 (N_8532,N_8255,N_8394);
nor U8533 (N_8533,N_8236,N_8322);
nand U8534 (N_8534,N_8358,N_8317);
nor U8535 (N_8535,N_8380,N_8320);
xor U8536 (N_8536,N_8223,N_8364);
nor U8537 (N_8537,N_8363,N_8231);
xnor U8538 (N_8538,N_8293,N_8389);
and U8539 (N_8539,N_8295,N_8330);
or U8540 (N_8540,N_8328,N_8270);
xor U8541 (N_8541,N_8374,N_8260);
or U8542 (N_8542,N_8354,N_8286);
or U8543 (N_8543,N_8364,N_8374);
xnor U8544 (N_8544,N_8281,N_8259);
or U8545 (N_8545,N_8227,N_8373);
or U8546 (N_8546,N_8368,N_8229);
xor U8547 (N_8547,N_8209,N_8360);
nor U8548 (N_8548,N_8211,N_8380);
xor U8549 (N_8549,N_8361,N_8200);
or U8550 (N_8550,N_8263,N_8365);
or U8551 (N_8551,N_8306,N_8246);
nand U8552 (N_8552,N_8353,N_8395);
xnor U8553 (N_8553,N_8395,N_8355);
nand U8554 (N_8554,N_8361,N_8268);
xnor U8555 (N_8555,N_8310,N_8334);
and U8556 (N_8556,N_8311,N_8357);
or U8557 (N_8557,N_8368,N_8340);
nand U8558 (N_8558,N_8278,N_8284);
or U8559 (N_8559,N_8364,N_8203);
xnor U8560 (N_8560,N_8209,N_8368);
or U8561 (N_8561,N_8377,N_8335);
and U8562 (N_8562,N_8263,N_8254);
xor U8563 (N_8563,N_8236,N_8210);
and U8564 (N_8564,N_8237,N_8299);
nand U8565 (N_8565,N_8258,N_8352);
xnor U8566 (N_8566,N_8245,N_8264);
nor U8567 (N_8567,N_8295,N_8288);
nand U8568 (N_8568,N_8395,N_8292);
or U8569 (N_8569,N_8314,N_8313);
nor U8570 (N_8570,N_8259,N_8223);
and U8571 (N_8571,N_8232,N_8395);
or U8572 (N_8572,N_8238,N_8225);
or U8573 (N_8573,N_8298,N_8313);
or U8574 (N_8574,N_8293,N_8363);
nor U8575 (N_8575,N_8211,N_8229);
or U8576 (N_8576,N_8219,N_8375);
nor U8577 (N_8577,N_8360,N_8362);
and U8578 (N_8578,N_8347,N_8230);
nor U8579 (N_8579,N_8347,N_8315);
nor U8580 (N_8580,N_8375,N_8231);
nor U8581 (N_8581,N_8339,N_8373);
nor U8582 (N_8582,N_8294,N_8290);
and U8583 (N_8583,N_8221,N_8321);
xnor U8584 (N_8584,N_8226,N_8219);
nand U8585 (N_8585,N_8378,N_8248);
xnor U8586 (N_8586,N_8398,N_8392);
nor U8587 (N_8587,N_8366,N_8320);
xor U8588 (N_8588,N_8326,N_8281);
nand U8589 (N_8589,N_8263,N_8235);
and U8590 (N_8590,N_8349,N_8251);
or U8591 (N_8591,N_8386,N_8279);
nor U8592 (N_8592,N_8309,N_8298);
nand U8593 (N_8593,N_8265,N_8232);
and U8594 (N_8594,N_8343,N_8358);
or U8595 (N_8595,N_8203,N_8227);
or U8596 (N_8596,N_8268,N_8202);
nor U8597 (N_8597,N_8281,N_8211);
nand U8598 (N_8598,N_8366,N_8231);
xnor U8599 (N_8599,N_8369,N_8351);
nand U8600 (N_8600,N_8519,N_8524);
or U8601 (N_8601,N_8483,N_8549);
or U8602 (N_8602,N_8468,N_8571);
nand U8603 (N_8603,N_8494,N_8504);
and U8604 (N_8604,N_8499,N_8560);
and U8605 (N_8605,N_8540,N_8591);
xor U8606 (N_8606,N_8430,N_8428);
or U8607 (N_8607,N_8570,N_8528);
and U8608 (N_8608,N_8522,N_8464);
xor U8609 (N_8609,N_8520,N_8594);
xor U8610 (N_8610,N_8424,N_8467);
nand U8611 (N_8611,N_8492,N_8409);
xor U8612 (N_8612,N_8505,N_8568);
or U8613 (N_8613,N_8586,N_8403);
xnor U8614 (N_8614,N_8421,N_8407);
xor U8615 (N_8615,N_8523,N_8542);
and U8616 (N_8616,N_8443,N_8441);
or U8617 (N_8617,N_8497,N_8412);
xnor U8618 (N_8618,N_8429,N_8511);
nand U8619 (N_8619,N_8416,N_8580);
and U8620 (N_8620,N_8425,N_8454);
nor U8621 (N_8621,N_8547,N_8525);
nor U8622 (N_8622,N_8556,N_8593);
nand U8623 (N_8623,N_8419,N_8455);
xnor U8624 (N_8624,N_8402,N_8436);
nor U8625 (N_8625,N_8590,N_8431);
and U8626 (N_8626,N_8582,N_8588);
and U8627 (N_8627,N_8587,N_8501);
nand U8628 (N_8628,N_8413,N_8411);
nand U8629 (N_8629,N_8485,N_8521);
or U8630 (N_8630,N_8566,N_8446);
nor U8631 (N_8631,N_8539,N_8529);
nand U8632 (N_8632,N_8562,N_8526);
and U8633 (N_8633,N_8400,N_8434);
nor U8634 (N_8634,N_8487,N_8432);
and U8635 (N_8635,N_8466,N_8415);
or U8636 (N_8636,N_8496,N_8548);
xnor U8637 (N_8637,N_8410,N_8583);
xnor U8638 (N_8638,N_8546,N_8442);
nand U8639 (N_8639,N_8445,N_8489);
or U8640 (N_8640,N_8417,N_8453);
nor U8641 (N_8641,N_8532,N_8543);
nand U8642 (N_8642,N_8498,N_8545);
and U8643 (N_8643,N_8473,N_8535);
xor U8644 (N_8644,N_8476,N_8598);
xnor U8645 (N_8645,N_8506,N_8584);
nor U8646 (N_8646,N_8507,N_8479);
and U8647 (N_8647,N_8564,N_8533);
or U8648 (N_8648,N_8437,N_8401);
xnor U8649 (N_8649,N_8555,N_8508);
or U8650 (N_8650,N_8527,N_8449);
nand U8651 (N_8651,N_8444,N_8552);
nor U8652 (N_8652,N_8551,N_8544);
and U8653 (N_8653,N_8484,N_8558);
xnor U8654 (N_8654,N_8510,N_8460);
xor U8655 (N_8655,N_8472,N_8541);
nor U8656 (N_8656,N_8530,N_8537);
or U8657 (N_8657,N_8477,N_8567);
or U8658 (N_8658,N_8516,N_8486);
or U8659 (N_8659,N_8518,N_8592);
or U8660 (N_8660,N_8481,N_8482);
and U8661 (N_8661,N_8517,N_8463);
nand U8662 (N_8662,N_8578,N_8475);
nor U8663 (N_8663,N_8509,N_8561);
xnor U8664 (N_8664,N_8420,N_8534);
or U8665 (N_8665,N_8465,N_8565);
nand U8666 (N_8666,N_8559,N_8576);
nor U8667 (N_8667,N_8435,N_8480);
and U8668 (N_8668,N_8438,N_8563);
nand U8669 (N_8669,N_8423,N_8513);
nand U8670 (N_8670,N_8433,N_8554);
xnor U8671 (N_8671,N_8448,N_8488);
xor U8672 (N_8672,N_8447,N_8422);
xnor U8673 (N_8673,N_8462,N_8469);
xnor U8674 (N_8674,N_8531,N_8585);
and U8675 (N_8675,N_8406,N_8404);
nor U8676 (N_8676,N_8495,N_8490);
xor U8677 (N_8677,N_8572,N_8502);
xor U8678 (N_8678,N_8599,N_8575);
nor U8679 (N_8679,N_8408,N_8457);
nor U8680 (N_8680,N_8451,N_8470);
nor U8681 (N_8681,N_8474,N_8515);
nand U8682 (N_8682,N_8456,N_8500);
and U8683 (N_8683,N_8589,N_8557);
or U8684 (N_8684,N_8596,N_8569);
xor U8685 (N_8685,N_8478,N_8512);
or U8686 (N_8686,N_8418,N_8450);
or U8687 (N_8687,N_8581,N_8426);
or U8688 (N_8688,N_8459,N_8553);
nand U8689 (N_8689,N_8439,N_8493);
nand U8690 (N_8690,N_8597,N_8579);
and U8691 (N_8691,N_8514,N_8471);
nor U8692 (N_8692,N_8405,N_8414);
nor U8693 (N_8693,N_8458,N_8503);
or U8694 (N_8694,N_8538,N_8427);
nand U8695 (N_8695,N_8440,N_8461);
nor U8696 (N_8696,N_8491,N_8595);
nor U8697 (N_8697,N_8577,N_8550);
xnor U8698 (N_8698,N_8536,N_8452);
and U8699 (N_8699,N_8573,N_8574);
and U8700 (N_8700,N_8583,N_8403);
xnor U8701 (N_8701,N_8544,N_8541);
and U8702 (N_8702,N_8446,N_8402);
nor U8703 (N_8703,N_8421,N_8427);
and U8704 (N_8704,N_8572,N_8598);
and U8705 (N_8705,N_8405,N_8540);
or U8706 (N_8706,N_8500,N_8578);
nand U8707 (N_8707,N_8534,N_8431);
nand U8708 (N_8708,N_8448,N_8402);
nand U8709 (N_8709,N_8480,N_8559);
nor U8710 (N_8710,N_8439,N_8538);
and U8711 (N_8711,N_8566,N_8557);
nor U8712 (N_8712,N_8470,N_8410);
nor U8713 (N_8713,N_8510,N_8585);
xnor U8714 (N_8714,N_8549,N_8429);
nor U8715 (N_8715,N_8516,N_8583);
nor U8716 (N_8716,N_8595,N_8525);
or U8717 (N_8717,N_8462,N_8438);
or U8718 (N_8718,N_8414,N_8586);
and U8719 (N_8719,N_8451,N_8580);
xor U8720 (N_8720,N_8573,N_8503);
xnor U8721 (N_8721,N_8503,N_8530);
nand U8722 (N_8722,N_8534,N_8519);
and U8723 (N_8723,N_8477,N_8585);
nor U8724 (N_8724,N_8452,N_8598);
nand U8725 (N_8725,N_8475,N_8500);
nor U8726 (N_8726,N_8505,N_8430);
xnor U8727 (N_8727,N_8592,N_8419);
xor U8728 (N_8728,N_8579,N_8441);
or U8729 (N_8729,N_8514,N_8421);
xor U8730 (N_8730,N_8446,N_8410);
and U8731 (N_8731,N_8532,N_8585);
and U8732 (N_8732,N_8476,N_8552);
nand U8733 (N_8733,N_8492,N_8547);
and U8734 (N_8734,N_8525,N_8496);
nor U8735 (N_8735,N_8422,N_8592);
or U8736 (N_8736,N_8533,N_8596);
xor U8737 (N_8737,N_8416,N_8523);
or U8738 (N_8738,N_8460,N_8419);
or U8739 (N_8739,N_8492,N_8497);
nand U8740 (N_8740,N_8506,N_8427);
xor U8741 (N_8741,N_8466,N_8474);
xor U8742 (N_8742,N_8429,N_8536);
xor U8743 (N_8743,N_8550,N_8494);
xnor U8744 (N_8744,N_8586,N_8439);
or U8745 (N_8745,N_8417,N_8400);
nor U8746 (N_8746,N_8433,N_8453);
or U8747 (N_8747,N_8472,N_8418);
xnor U8748 (N_8748,N_8431,N_8511);
or U8749 (N_8749,N_8513,N_8405);
nand U8750 (N_8750,N_8498,N_8598);
nand U8751 (N_8751,N_8548,N_8453);
nor U8752 (N_8752,N_8416,N_8404);
or U8753 (N_8753,N_8534,N_8524);
nor U8754 (N_8754,N_8551,N_8433);
xor U8755 (N_8755,N_8448,N_8537);
xor U8756 (N_8756,N_8476,N_8479);
xor U8757 (N_8757,N_8580,N_8515);
xor U8758 (N_8758,N_8572,N_8499);
nand U8759 (N_8759,N_8455,N_8408);
and U8760 (N_8760,N_8470,N_8480);
nor U8761 (N_8761,N_8506,N_8572);
xnor U8762 (N_8762,N_8430,N_8477);
xor U8763 (N_8763,N_8415,N_8566);
nor U8764 (N_8764,N_8477,N_8450);
or U8765 (N_8765,N_8566,N_8560);
nand U8766 (N_8766,N_8567,N_8513);
nor U8767 (N_8767,N_8461,N_8557);
or U8768 (N_8768,N_8576,N_8473);
nor U8769 (N_8769,N_8499,N_8426);
nand U8770 (N_8770,N_8408,N_8434);
nor U8771 (N_8771,N_8469,N_8588);
nor U8772 (N_8772,N_8435,N_8575);
xnor U8773 (N_8773,N_8519,N_8400);
nor U8774 (N_8774,N_8520,N_8513);
nor U8775 (N_8775,N_8433,N_8512);
xor U8776 (N_8776,N_8466,N_8514);
nand U8777 (N_8777,N_8500,N_8478);
or U8778 (N_8778,N_8555,N_8416);
and U8779 (N_8779,N_8580,N_8550);
nand U8780 (N_8780,N_8436,N_8505);
xnor U8781 (N_8781,N_8402,N_8542);
xnor U8782 (N_8782,N_8451,N_8490);
and U8783 (N_8783,N_8481,N_8517);
and U8784 (N_8784,N_8454,N_8509);
and U8785 (N_8785,N_8567,N_8558);
or U8786 (N_8786,N_8473,N_8560);
or U8787 (N_8787,N_8492,N_8472);
and U8788 (N_8788,N_8509,N_8428);
xor U8789 (N_8789,N_8475,N_8566);
xor U8790 (N_8790,N_8429,N_8542);
nor U8791 (N_8791,N_8550,N_8488);
or U8792 (N_8792,N_8446,N_8587);
nand U8793 (N_8793,N_8502,N_8508);
xor U8794 (N_8794,N_8410,N_8554);
xor U8795 (N_8795,N_8411,N_8581);
nor U8796 (N_8796,N_8476,N_8443);
and U8797 (N_8797,N_8513,N_8495);
nor U8798 (N_8798,N_8410,N_8494);
or U8799 (N_8799,N_8466,N_8465);
and U8800 (N_8800,N_8679,N_8738);
nand U8801 (N_8801,N_8767,N_8658);
nor U8802 (N_8802,N_8702,N_8778);
and U8803 (N_8803,N_8615,N_8717);
or U8804 (N_8804,N_8781,N_8613);
or U8805 (N_8805,N_8796,N_8725);
or U8806 (N_8806,N_8712,N_8713);
and U8807 (N_8807,N_8697,N_8633);
nor U8808 (N_8808,N_8783,N_8771);
or U8809 (N_8809,N_8625,N_8718);
nor U8810 (N_8810,N_8657,N_8762);
and U8811 (N_8811,N_8793,N_8775);
nand U8812 (N_8812,N_8648,N_8608);
or U8813 (N_8813,N_8678,N_8690);
nor U8814 (N_8814,N_8790,N_8716);
xor U8815 (N_8815,N_8766,N_8644);
or U8816 (N_8816,N_8704,N_8681);
nand U8817 (N_8817,N_8668,N_8662);
and U8818 (N_8818,N_8784,N_8720);
xnor U8819 (N_8819,N_8683,N_8753);
and U8820 (N_8820,N_8671,N_8741);
nand U8821 (N_8821,N_8721,N_8643);
or U8822 (N_8822,N_8743,N_8711);
or U8823 (N_8823,N_8669,N_8707);
and U8824 (N_8824,N_8664,N_8730);
xor U8825 (N_8825,N_8611,N_8618);
xor U8826 (N_8826,N_8777,N_8659);
and U8827 (N_8827,N_8774,N_8645);
nor U8828 (N_8828,N_8715,N_8769);
nor U8829 (N_8829,N_8626,N_8792);
nor U8830 (N_8830,N_8699,N_8619);
nand U8831 (N_8831,N_8772,N_8752);
and U8832 (N_8832,N_8627,N_8734);
and U8833 (N_8833,N_8764,N_8677);
and U8834 (N_8834,N_8749,N_8731);
and U8835 (N_8835,N_8761,N_8785);
or U8836 (N_8836,N_8634,N_8651);
nand U8837 (N_8837,N_8791,N_8685);
nor U8838 (N_8838,N_8632,N_8603);
xnor U8839 (N_8839,N_8672,N_8691);
nand U8840 (N_8840,N_8750,N_8795);
nor U8841 (N_8841,N_8710,N_8757);
and U8842 (N_8842,N_8705,N_8649);
xor U8843 (N_8843,N_8675,N_8676);
nand U8844 (N_8844,N_8745,N_8622);
xor U8845 (N_8845,N_8620,N_8663);
nand U8846 (N_8846,N_8700,N_8751);
nor U8847 (N_8847,N_8639,N_8709);
xor U8848 (N_8848,N_8740,N_8661);
xor U8849 (N_8849,N_8742,N_8698);
or U8850 (N_8850,N_8798,N_8797);
nor U8851 (N_8851,N_8760,N_8727);
nand U8852 (N_8852,N_8708,N_8744);
xor U8853 (N_8853,N_8674,N_8794);
nand U8854 (N_8854,N_8736,N_8748);
xor U8855 (N_8855,N_8688,N_8600);
nand U8856 (N_8856,N_8637,N_8650);
or U8857 (N_8857,N_8682,N_8696);
nor U8858 (N_8858,N_8636,N_8621);
nand U8859 (N_8859,N_8780,N_8601);
xor U8860 (N_8860,N_8602,N_8779);
nand U8861 (N_8861,N_8733,N_8693);
nand U8862 (N_8862,N_8703,N_8723);
nor U8863 (N_8863,N_8695,N_8799);
nor U8864 (N_8864,N_8630,N_8729);
nor U8865 (N_8865,N_8694,N_8635);
and U8866 (N_8866,N_8692,N_8673);
nor U8867 (N_8867,N_8786,N_8670);
and U8868 (N_8868,N_8624,N_8789);
xor U8869 (N_8869,N_8655,N_8647);
xnor U8870 (N_8870,N_8638,N_8641);
and U8871 (N_8871,N_8628,N_8763);
and U8872 (N_8872,N_8656,N_8640);
nand U8873 (N_8873,N_8646,N_8684);
xnor U8874 (N_8874,N_8680,N_8667);
nand U8875 (N_8875,N_8714,N_8623);
or U8876 (N_8876,N_8701,N_8758);
nor U8877 (N_8877,N_8768,N_8689);
xor U8878 (N_8878,N_8614,N_8739);
nor U8879 (N_8879,N_8687,N_8732);
or U8880 (N_8880,N_8631,N_8756);
xor U8881 (N_8881,N_8719,N_8787);
and U8882 (N_8882,N_8610,N_8724);
and U8883 (N_8883,N_8735,N_8617);
and U8884 (N_8884,N_8686,N_8607);
nor U8885 (N_8885,N_8629,N_8747);
nand U8886 (N_8886,N_8782,N_8665);
nor U8887 (N_8887,N_8605,N_8737);
or U8888 (N_8888,N_8754,N_8706);
and U8889 (N_8889,N_8612,N_8606);
and U8890 (N_8890,N_8773,N_8746);
nor U8891 (N_8891,N_8616,N_8642);
or U8892 (N_8892,N_8666,N_8770);
nor U8893 (N_8893,N_8788,N_8604);
nand U8894 (N_8894,N_8755,N_8765);
and U8895 (N_8895,N_8726,N_8722);
nor U8896 (N_8896,N_8728,N_8654);
or U8897 (N_8897,N_8759,N_8776);
or U8898 (N_8898,N_8652,N_8653);
or U8899 (N_8899,N_8609,N_8660);
xor U8900 (N_8900,N_8675,N_8621);
xnor U8901 (N_8901,N_8633,N_8672);
nand U8902 (N_8902,N_8798,N_8709);
nand U8903 (N_8903,N_8616,N_8714);
or U8904 (N_8904,N_8688,N_8797);
and U8905 (N_8905,N_8678,N_8741);
nand U8906 (N_8906,N_8798,N_8707);
xor U8907 (N_8907,N_8777,N_8766);
nand U8908 (N_8908,N_8671,N_8779);
and U8909 (N_8909,N_8709,N_8615);
and U8910 (N_8910,N_8794,N_8627);
and U8911 (N_8911,N_8781,N_8722);
xor U8912 (N_8912,N_8771,N_8784);
xor U8913 (N_8913,N_8703,N_8697);
nand U8914 (N_8914,N_8747,N_8727);
or U8915 (N_8915,N_8740,N_8624);
nor U8916 (N_8916,N_8766,N_8681);
and U8917 (N_8917,N_8787,N_8709);
xnor U8918 (N_8918,N_8748,N_8796);
and U8919 (N_8919,N_8691,N_8776);
nor U8920 (N_8920,N_8694,N_8685);
nor U8921 (N_8921,N_8631,N_8724);
or U8922 (N_8922,N_8795,N_8654);
nand U8923 (N_8923,N_8661,N_8776);
nor U8924 (N_8924,N_8734,N_8715);
nand U8925 (N_8925,N_8656,N_8729);
xor U8926 (N_8926,N_8702,N_8729);
and U8927 (N_8927,N_8777,N_8748);
xnor U8928 (N_8928,N_8777,N_8634);
and U8929 (N_8929,N_8725,N_8682);
nand U8930 (N_8930,N_8785,N_8618);
nand U8931 (N_8931,N_8666,N_8613);
xnor U8932 (N_8932,N_8762,N_8607);
and U8933 (N_8933,N_8755,N_8778);
or U8934 (N_8934,N_8776,N_8733);
and U8935 (N_8935,N_8751,N_8719);
nand U8936 (N_8936,N_8782,N_8613);
or U8937 (N_8937,N_8746,N_8732);
or U8938 (N_8938,N_8617,N_8637);
or U8939 (N_8939,N_8626,N_8793);
nor U8940 (N_8940,N_8652,N_8723);
and U8941 (N_8941,N_8782,N_8651);
and U8942 (N_8942,N_8729,N_8638);
nand U8943 (N_8943,N_8614,N_8664);
nor U8944 (N_8944,N_8780,N_8649);
nor U8945 (N_8945,N_8627,N_8795);
xor U8946 (N_8946,N_8787,N_8658);
xor U8947 (N_8947,N_8794,N_8619);
nor U8948 (N_8948,N_8601,N_8776);
and U8949 (N_8949,N_8638,N_8689);
and U8950 (N_8950,N_8670,N_8766);
xor U8951 (N_8951,N_8650,N_8724);
and U8952 (N_8952,N_8645,N_8605);
nand U8953 (N_8953,N_8600,N_8678);
xnor U8954 (N_8954,N_8737,N_8630);
or U8955 (N_8955,N_8762,N_8610);
nor U8956 (N_8956,N_8695,N_8653);
nor U8957 (N_8957,N_8777,N_8626);
nor U8958 (N_8958,N_8724,N_8640);
xor U8959 (N_8959,N_8763,N_8685);
nor U8960 (N_8960,N_8610,N_8740);
or U8961 (N_8961,N_8609,N_8634);
xnor U8962 (N_8962,N_8745,N_8741);
nand U8963 (N_8963,N_8679,N_8642);
xor U8964 (N_8964,N_8750,N_8773);
and U8965 (N_8965,N_8628,N_8685);
xor U8966 (N_8966,N_8646,N_8633);
nor U8967 (N_8967,N_8750,N_8693);
nand U8968 (N_8968,N_8607,N_8766);
and U8969 (N_8969,N_8685,N_8661);
nor U8970 (N_8970,N_8610,N_8680);
or U8971 (N_8971,N_8783,N_8637);
nor U8972 (N_8972,N_8656,N_8769);
or U8973 (N_8973,N_8755,N_8742);
nor U8974 (N_8974,N_8690,N_8763);
or U8975 (N_8975,N_8788,N_8618);
nor U8976 (N_8976,N_8795,N_8609);
and U8977 (N_8977,N_8756,N_8731);
nand U8978 (N_8978,N_8714,N_8691);
or U8979 (N_8979,N_8677,N_8623);
nor U8980 (N_8980,N_8767,N_8780);
xor U8981 (N_8981,N_8737,N_8751);
xor U8982 (N_8982,N_8648,N_8759);
xor U8983 (N_8983,N_8640,N_8784);
nor U8984 (N_8984,N_8690,N_8655);
nor U8985 (N_8985,N_8620,N_8667);
and U8986 (N_8986,N_8668,N_8739);
nand U8987 (N_8987,N_8796,N_8706);
xnor U8988 (N_8988,N_8670,N_8687);
or U8989 (N_8989,N_8628,N_8723);
and U8990 (N_8990,N_8676,N_8608);
or U8991 (N_8991,N_8650,N_8707);
or U8992 (N_8992,N_8789,N_8601);
nand U8993 (N_8993,N_8625,N_8686);
or U8994 (N_8994,N_8757,N_8796);
or U8995 (N_8995,N_8627,N_8745);
nor U8996 (N_8996,N_8775,N_8742);
xnor U8997 (N_8997,N_8768,N_8747);
nor U8998 (N_8998,N_8645,N_8708);
nand U8999 (N_8999,N_8639,N_8797);
nor U9000 (N_9000,N_8897,N_8976);
nor U9001 (N_9001,N_8834,N_8998);
or U9002 (N_9002,N_8810,N_8974);
and U9003 (N_9003,N_8882,N_8957);
or U9004 (N_9004,N_8970,N_8826);
nor U9005 (N_9005,N_8914,N_8903);
or U9006 (N_9006,N_8991,N_8954);
xnor U9007 (N_9007,N_8868,N_8931);
and U9008 (N_9008,N_8862,N_8953);
or U9009 (N_9009,N_8888,N_8873);
and U9010 (N_9010,N_8987,N_8945);
xnor U9011 (N_9011,N_8892,N_8857);
or U9012 (N_9012,N_8825,N_8912);
and U9013 (N_9013,N_8889,N_8930);
xnor U9014 (N_9014,N_8967,N_8969);
and U9015 (N_9015,N_8869,N_8994);
and U9016 (N_9016,N_8828,N_8922);
nor U9017 (N_9017,N_8803,N_8858);
xor U9018 (N_9018,N_8900,N_8846);
nor U9019 (N_9019,N_8937,N_8962);
nor U9020 (N_9020,N_8805,N_8812);
xnor U9021 (N_9021,N_8843,N_8879);
xor U9022 (N_9022,N_8815,N_8850);
or U9023 (N_9023,N_8997,N_8839);
xnor U9024 (N_9024,N_8916,N_8919);
xnor U9025 (N_9025,N_8877,N_8844);
nand U9026 (N_9026,N_8866,N_8872);
xnor U9027 (N_9027,N_8951,N_8980);
or U9028 (N_9028,N_8935,N_8949);
nor U9029 (N_9029,N_8856,N_8863);
or U9030 (N_9030,N_8943,N_8800);
or U9031 (N_9031,N_8847,N_8999);
nand U9032 (N_9032,N_8848,N_8822);
nor U9033 (N_9033,N_8896,N_8865);
or U9034 (N_9034,N_8852,N_8979);
nor U9035 (N_9035,N_8905,N_8838);
and U9036 (N_9036,N_8944,N_8878);
and U9037 (N_9037,N_8824,N_8929);
xor U9038 (N_9038,N_8817,N_8819);
nand U9039 (N_9039,N_8818,N_8915);
nor U9040 (N_9040,N_8885,N_8958);
or U9041 (N_9041,N_8933,N_8904);
nand U9042 (N_9042,N_8936,N_8978);
nor U9043 (N_9043,N_8995,N_8870);
nor U9044 (N_9044,N_8895,N_8876);
xnor U9045 (N_9045,N_8984,N_8926);
xnor U9046 (N_9046,N_8910,N_8963);
nand U9047 (N_9047,N_8938,N_8830);
and U9048 (N_9048,N_8851,N_8906);
nand U9049 (N_9049,N_8845,N_8874);
or U9050 (N_9050,N_8940,N_8939);
nor U9051 (N_9051,N_8941,N_8855);
xnor U9052 (N_9052,N_8881,N_8948);
nand U9053 (N_9053,N_8801,N_8871);
nor U9054 (N_9054,N_8809,N_8802);
and U9055 (N_9055,N_8861,N_8902);
xnor U9056 (N_9056,N_8966,N_8985);
or U9057 (N_9057,N_8835,N_8911);
or U9058 (N_9058,N_8956,N_8917);
nand U9059 (N_9059,N_8981,N_8833);
nand U9060 (N_9060,N_8836,N_8859);
nor U9061 (N_9061,N_8921,N_8955);
and U9062 (N_9062,N_8925,N_8989);
or U9063 (N_9063,N_8832,N_8831);
nor U9064 (N_9064,N_8960,N_8913);
or U9065 (N_9065,N_8886,N_8808);
nand U9066 (N_9066,N_8840,N_8952);
or U9067 (N_9067,N_8827,N_8927);
nor U9068 (N_9068,N_8829,N_8883);
and U9069 (N_9069,N_8982,N_8806);
or U9070 (N_9070,N_8977,N_8814);
nor U9071 (N_9071,N_8901,N_8990);
nor U9072 (N_9072,N_8934,N_8988);
xnor U9073 (N_9073,N_8853,N_8946);
and U9074 (N_9074,N_8964,N_8993);
or U9075 (N_9075,N_8924,N_8908);
nor U9076 (N_9076,N_8959,N_8983);
nand U9077 (N_9077,N_8986,N_8899);
and U9078 (N_9078,N_8961,N_8884);
or U9079 (N_9079,N_8894,N_8820);
nand U9080 (N_9080,N_8880,N_8816);
nor U9081 (N_9081,N_8932,N_8975);
nor U9082 (N_9082,N_8972,N_8968);
or U9083 (N_9083,N_8860,N_8807);
nor U9084 (N_9084,N_8849,N_8875);
nor U9085 (N_9085,N_8837,N_8923);
xor U9086 (N_9086,N_8907,N_8854);
nand U9087 (N_9087,N_8804,N_8973);
nand U9088 (N_9088,N_8928,N_8909);
or U9089 (N_9089,N_8965,N_8992);
or U9090 (N_9090,N_8887,N_8890);
xor U9091 (N_9091,N_8813,N_8920);
nand U9092 (N_9092,N_8971,N_8918);
or U9093 (N_9093,N_8891,N_8950);
nand U9094 (N_9094,N_8821,N_8947);
or U9095 (N_9095,N_8942,N_8842);
nor U9096 (N_9096,N_8898,N_8841);
or U9097 (N_9097,N_8823,N_8893);
nand U9098 (N_9098,N_8811,N_8996);
and U9099 (N_9099,N_8864,N_8867);
nand U9100 (N_9100,N_8861,N_8977);
nand U9101 (N_9101,N_8860,N_8923);
nand U9102 (N_9102,N_8863,N_8899);
or U9103 (N_9103,N_8944,N_8975);
and U9104 (N_9104,N_8897,N_8862);
nand U9105 (N_9105,N_8955,N_8992);
and U9106 (N_9106,N_8931,N_8967);
nand U9107 (N_9107,N_8822,N_8906);
and U9108 (N_9108,N_8917,N_8830);
nor U9109 (N_9109,N_8851,N_8924);
xnor U9110 (N_9110,N_8993,N_8900);
nand U9111 (N_9111,N_8830,N_8800);
xor U9112 (N_9112,N_8829,N_8854);
nor U9113 (N_9113,N_8967,N_8830);
or U9114 (N_9114,N_8975,N_8955);
nand U9115 (N_9115,N_8991,N_8802);
xor U9116 (N_9116,N_8917,N_8850);
nor U9117 (N_9117,N_8827,N_8979);
or U9118 (N_9118,N_8966,N_8886);
nor U9119 (N_9119,N_8915,N_8926);
nand U9120 (N_9120,N_8939,N_8925);
nor U9121 (N_9121,N_8949,N_8926);
and U9122 (N_9122,N_8995,N_8977);
nand U9123 (N_9123,N_8896,N_8957);
and U9124 (N_9124,N_8930,N_8941);
nor U9125 (N_9125,N_8929,N_8830);
nor U9126 (N_9126,N_8940,N_8914);
xnor U9127 (N_9127,N_8821,N_8939);
and U9128 (N_9128,N_8852,N_8940);
nand U9129 (N_9129,N_8982,N_8916);
and U9130 (N_9130,N_8941,N_8813);
nor U9131 (N_9131,N_8922,N_8892);
and U9132 (N_9132,N_8841,N_8880);
xnor U9133 (N_9133,N_8926,N_8822);
and U9134 (N_9134,N_8869,N_8983);
xor U9135 (N_9135,N_8890,N_8862);
xnor U9136 (N_9136,N_8887,N_8884);
nand U9137 (N_9137,N_8988,N_8956);
nand U9138 (N_9138,N_8896,N_8813);
or U9139 (N_9139,N_8965,N_8936);
nand U9140 (N_9140,N_8965,N_8924);
nor U9141 (N_9141,N_8937,N_8810);
nand U9142 (N_9142,N_8878,N_8904);
nand U9143 (N_9143,N_8845,N_8823);
nor U9144 (N_9144,N_8869,N_8809);
and U9145 (N_9145,N_8952,N_8816);
or U9146 (N_9146,N_8866,N_8897);
xnor U9147 (N_9147,N_8972,N_8917);
and U9148 (N_9148,N_8897,N_8838);
xor U9149 (N_9149,N_8805,N_8962);
xor U9150 (N_9150,N_8862,N_8879);
nand U9151 (N_9151,N_8997,N_8859);
nand U9152 (N_9152,N_8896,N_8818);
and U9153 (N_9153,N_8808,N_8971);
and U9154 (N_9154,N_8881,N_8951);
nand U9155 (N_9155,N_8976,N_8962);
nand U9156 (N_9156,N_8847,N_8928);
and U9157 (N_9157,N_8835,N_8848);
and U9158 (N_9158,N_8814,N_8855);
or U9159 (N_9159,N_8866,N_8903);
xor U9160 (N_9160,N_8989,N_8866);
xor U9161 (N_9161,N_8919,N_8943);
or U9162 (N_9162,N_8903,N_8917);
xor U9163 (N_9163,N_8981,N_8992);
xor U9164 (N_9164,N_8837,N_8914);
nor U9165 (N_9165,N_8895,N_8849);
or U9166 (N_9166,N_8975,N_8852);
and U9167 (N_9167,N_8801,N_8944);
and U9168 (N_9168,N_8910,N_8947);
xor U9169 (N_9169,N_8833,N_8940);
xor U9170 (N_9170,N_8861,N_8837);
or U9171 (N_9171,N_8884,N_8882);
nand U9172 (N_9172,N_8818,N_8835);
or U9173 (N_9173,N_8978,N_8847);
nand U9174 (N_9174,N_8989,N_8896);
or U9175 (N_9175,N_8809,N_8901);
xor U9176 (N_9176,N_8802,N_8861);
or U9177 (N_9177,N_8972,N_8966);
or U9178 (N_9178,N_8819,N_8996);
nand U9179 (N_9179,N_8977,N_8999);
xor U9180 (N_9180,N_8906,N_8882);
nor U9181 (N_9181,N_8822,N_8823);
and U9182 (N_9182,N_8888,N_8992);
nor U9183 (N_9183,N_8810,N_8995);
xnor U9184 (N_9184,N_8845,N_8918);
or U9185 (N_9185,N_8911,N_8941);
and U9186 (N_9186,N_8883,N_8952);
nand U9187 (N_9187,N_8891,N_8952);
or U9188 (N_9188,N_8858,N_8994);
and U9189 (N_9189,N_8892,N_8935);
xnor U9190 (N_9190,N_8848,N_8977);
nand U9191 (N_9191,N_8864,N_8850);
and U9192 (N_9192,N_8995,N_8884);
and U9193 (N_9193,N_8927,N_8905);
or U9194 (N_9194,N_8992,N_8985);
nor U9195 (N_9195,N_8875,N_8832);
or U9196 (N_9196,N_8979,N_8967);
nor U9197 (N_9197,N_8881,N_8990);
or U9198 (N_9198,N_8976,N_8830);
or U9199 (N_9199,N_8957,N_8858);
and U9200 (N_9200,N_9183,N_9133);
nand U9201 (N_9201,N_9038,N_9167);
or U9202 (N_9202,N_9077,N_9034);
nor U9203 (N_9203,N_9061,N_9145);
nand U9204 (N_9204,N_9190,N_9069);
or U9205 (N_9205,N_9053,N_9011);
and U9206 (N_9206,N_9114,N_9031);
and U9207 (N_9207,N_9033,N_9189);
or U9208 (N_9208,N_9096,N_9067);
nor U9209 (N_9209,N_9132,N_9087);
nor U9210 (N_9210,N_9057,N_9079);
nand U9211 (N_9211,N_9180,N_9039);
nor U9212 (N_9212,N_9129,N_9122);
xor U9213 (N_9213,N_9004,N_9146);
xnor U9214 (N_9214,N_9107,N_9143);
or U9215 (N_9215,N_9020,N_9176);
or U9216 (N_9216,N_9005,N_9185);
nand U9217 (N_9217,N_9058,N_9121);
or U9218 (N_9218,N_9014,N_9175);
and U9219 (N_9219,N_9120,N_9100);
or U9220 (N_9220,N_9012,N_9163);
or U9221 (N_9221,N_9161,N_9018);
or U9222 (N_9222,N_9010,N_9188);
and U9223 (N_9223,N_9126,N_9098);
nand U9224 (N_9224,N_9088,N_9141);
and U9225 (N_9225,N_9108,N_9128);
nand U9226 (N_9226,N_9134,N_9062);
and U9227 (N_9227,N_9170,N_9097);
and U9228 (N_9228,N_9142,N_9001);
nor U9229 (N_9229,N_9086,N_9023);
nor U9230 (N_9230,N_9042,N_9055);
or U9231 (N_9231,N_9116,N_9144);
nor U9232 (N_9232,N_9191,N_9151);
or U9233 (N_9233,N_9021,N_9184);
or U9234 (N_9234,N_9193,N_9164);
or U9235 (N_9235,N_9169,N_9083);
xnor U9236 (N_9236,N_9019,N_9162);
xnor U9237 (N_9237,N_9150,N_9076);
xor U9238 (N_9238,N_9199,N_9090);
nor U9239 (N_9239,N_9040,N_9194);
xor U9240 (N_9240,N_9159,N_9196);
xnor U9241 (N_9241,N_9147,N_9047);
nor U9242 (N_9242,N_9093,N_9115);
xor U9243 (N_9243,N_9015,N_9008);
nor U9244 (N_9244,N_9095,N_9197);
and U9245 (N_9245,N_9056,N_9138);
xor U9246 (N_9246,N_9006,N_9025);
or U9247 (N_9247,N_9075,N_9137);
xnor U9248 (N_9248,N_9182,N_9152);
and U9249 (N_9249,N_9105,N_9106);
nand U9250 (N_9250,N_9043,N_9174);
or U9251 (N_9251,N_9080,N_9072);
and U9252 (N_9252,N_9037,N_9113);
xnor U9253 (N_9253,N_9073,N_9091);
and U9254 (N_9254,N_9082,N_9064);
or U9255 (N_9255,N_9022,N_9065);
xor U9256 (N_9256,N_9099,N_9111);
xor U9257 (N_9257,N_9028,N_9178);
or U9258 (N_9258,N_9066,N_9109);
and U9259 (N_9259,N_9166,N_9054);
nor U9260 (N_9260,N_9017,N_9172);
or U9261 (N_9261,N_9007,N_9112);
nor U9262 (N_9262,N_9063,N_9177);
nor U9263 (N_9263,N_9101,N_9050);
xor U9264 (N_9264,N_9002,N_9013);
xor U9265 (N_9265,N_9187,N_9181);
xor U9266 (N_9266,N_9110,N_9195);
and U9267 (N_9267,N_9027,N_9059);
nand U9268 (N_9268,N_9044,N_9102);
or U9269 (N_9269,N_9155,N_9060);
xnor U9270 (N_9270,N_9123,N_9168);
nor U9271 (N_9271,N_9000,N_9160);
nand U9272 (N_9272,N_9139,N_9165);
xnor U9273 (N_9273,N_9003,N_9009);
or U9274 (N_9274,N_9078,N_9148);
nand U9275 (N_9275,N_9092,N_9173);
xor U9276 (N_9276,N_9026,N_9046);
nand U9277 (N_9277,N_9081,N_9140);
nand U9278 (N_9278,N_9192,N_9045);
nand U9279 (N_9279,N_9089,N_9156);
or U9280 (N_9280,N_9186,N_9084);
or U9281 (N_9281,N_9131,N_9049);
nor U9282 (N_9282,N_9154,N_9094);
and U9283 (N_9283,N_9029,N_9117);
or U9284 (N_9284,N_9153,N_9158);
nor U9285 (N_9285,N_9085,N_9179);
and U9286 (N_9286,N_9048,N_9135);
or U9287 (N_9287,N_9071,N_9030);
and U9288 (N_9288,N_9035,N_9052);
or U9289 (N_9289,N_9119,N_9074);
and U9290 (N_9290,N_9068,N_9016);
and U9291 (N_9291,N_9149,N_9136);
nand U9292 (N_9292,N_9103,N_9157);
nor U9293 (N_9293,N_9130,N_9041);
and U9294 (N_9294,N_9198,N_9124);
and U9295 (N_9295,N_9127,N_9032);
nor U9296 (N_9296,N_9104,N_9125);
and U9297 (N_9297,N_9118,N_9024);
or U9298 (N_9298,N_9070,N_9051);
or U9299 (N_9299,N_9171,N_9036);
and U9300 (N_9300,N_9103,N_9088);
xnor U9301 (N_9301,N_9068,N_9020);
nor U9302 (N_9302,N_9147,N_9028);
nand U9303 (N_9303,N_9167,N_9069);
or U9304 (N_9304,N_9148,N_9193);
nor U9305 (N_9305,N_9183,N_9074);
nand U9306 (N_9306,N_9018,N_9158);
and U9307 (N_9307,N_9178,N_9015);
nand U9308 (N_9308,N_9187,N_9012);
nand U9309 (N_9309,N_9116,N_9038);
nor U9310 (N_9310,N_9028,N_9185);
xnor U9311 (N_9311,N_9132,N_9181);
nor U9312 (N_9312,N_9115,N_9057);
nand U9313 (N_9313,N_9159,N_9034);
xnor U9314 (N_9314,N_9033,N_9196);
and U9315 (N_9315,N_9099,N_9082);
nor U9316 (N_9316,N_9037,N_9160);
nand U9317 (N_9317,N_9099,N_9003);
nand U9318 (N_9318,N_9159,N_9053);
xnor U9319 (N_9319,N_9127,N_9187);
nor U9320 (N_9320,N_9020,N_9051);
xnor U9321 (N_9321,N_9109,N_9155);
nor U9322 (N_9322,N_9196,N_9122);
or U9323 (N_9323,N_9002,N_9063);
xor U9324 (N_9324,N_9009,N_9175);
or U9325 (N_9325,N_9176,N_9113);
nand U9326 (N_9326,N_9000,N_9050);
or U9327 (N_9327,N_9161,N_9089);
and U9328 (N_9328,N_9021,N_9105);
xor U9329 (N_9329,N_9018,N_9160);
nor U9330 (N_9330,N_9128,N_9157);
xor U9331 (N_9331,N_9029,N_9086);
xnor U9332 (N_9332,N_9025,N_9057);
and U9333 (N_9333,N_9127,N_9106);
and U9334 (N_9334,N_9171,N_9079);
and U9335 (N_9335,N_9057,N_9154);
and U9336 (N_9336,N_9038,N_9181);
nor U9337 (N_9337,N_9048,N_9026);
and U9338 (N_9338,N_9182,N_9094);
nand U9339 (N_9339,N_9114,N_9064);
nand U9340 (N_9340,N_9100,N_9177);
or U9341 (N_9341,N_9058,N_9068);
nand U9342 (N_9342,N_9023,N_9005);
nor U9343 (N_9343,N_9001,N_9178);
nand U9344 (N_9344,N_9021,N_9158);
nor U9345 (N_9345,N_9126,N_9066);
xor U9346 (N_9346,N_9175,N_9134);
nor U9347 (N_9347,N_9144,N_9128);
or U9348 (N_9348,N_9106,N_9160);
and U9349 (N_9349,N_9004,N_9126);
and U9350 (N_9350,N_9085,N_9188);
xor U9351 (N_9351,N_9141,N_9190);
nor U9352 (N_9352,N_9185,N_9104);
or U9353 (N_9353,N_9042,N_9167);
nand U9354 (N_9354,N_9168,N_9013);
or U9355 (N_9355,N_9059,N_9021);
or U9356 (N_9356,N_9122,N_9055);
or U9357 (N_9357,N_9103,N_9108);
or U9358 (N_9358,N_9007,N_9189);
and U9359 (N_9359,N_9110,N_9033);
nand U9360 (N_9360,N_9099,N_9153);
xnor U9361 (N_9361,N_9126,N_9012);
or U9362 (N_9362,N_9148,N_9013);
xor U9363 (N_9363,N_9033,N_9112);
nor U9364 (N_9364,N_9134,N_9131);
nor U9365 (N_9365,N_9142,N_9017);
nand U9366 (N_9366,N_9139,N_9135);
or U9367 (N_9367,N_9199,N_9078);
or U9368 (N_9368,N_9007,N_9124);
nor U9369 (N_9369,N_9154,N_9104);
or U9370 (N_9370,N_9025,N_9083);
nor U9371 (N_9371,N_9028,N_9177);
or U9372 (N_9372,N_9140,N_9079);
or U9373 (N_9373,N_9089,N_9167);
and U9374 (N_9374,N_9038,N_9190);
xnor U9375 (N_9375,N_9108,N_9184);
or U9376 (N_9376,N_9140,N_9136);
xnor U9377 (N_9377,N_9104,N_9084);
and U9378 (N_9378,N_9028,N_9009);
and U9379 (N_9379,N_9149,N_9135);
or U9380 (N_9380,N_9176,N_9160);
and U9381 (N_9381,N_9073,N_9046);
xor U9382 (N_9382,N_9162,N_9033);
nor U9383 (N_9383,N_9153,N_9050);
xor U9384 (N_9384,N_9033,N_9174);
nand U9385 (N_9385,N_9092,N_9165);
xnor U9386 (N_9386,N_9175,N_9094);
and U9387 (N_9387,N_9147,N_9019);
nand U9388 (N_9388,N_9036,N_9022);
nor U9389 (N_9389,N_9135,N_9128);
or U9390 (N_9390,N_9111,N_9042);
nand U9391 (N_9391,N_9042,N_9079);
xnor U9392 (N_9392,N_9046,N_9165);
nand U9393 (N_9393,N_9148,N_9068);
nand U9394 (N_9394,N_9179,N_9076);
nor U9395 (N_9395,N_9144,N_9084);
xor U9396 (N_9396,N_9085,N_9086);
or U9397 (N_9397,N_9171,N_9093);
nor U9398 (N_9398,N_9198,N_9049);
or U9399 (N_9399,N_9196,N_9068);
and U9400 (N_9400,N_9341,N_9245);
and U9401 (N_9401,N_9375,N_9218);
and U9402 (N_9402,N_9275,N_9346);
xnor U9403 (N_9403,N_9387,N_9364);
nand U9404 (N_9404,N_9351,N_9396);
or U9405 (N_9405,N_9269,N_9314);
xnor U9406 (N_9406,N_9271,N_9342);
or U9407 (N_9407,N_9238,N_9259);
or U9408 (N_9408,N_9258,N_9379);
nor U9409 (N_9409,N_9227,N_9250);
nor U9410 (N_9410,N_9260,N_9229);
nand U9411 (N_9411,N_9237,N_9241);
and U9412 (N_9412,N_9323,N_9270);
and U9413 (N_9413,N_9294,N_9251);
nor U9414 (N_9414,N_9284,N_9301);
nand U9415 (N_9415,N_9228,N_9358);
and U9416 (N_9416,N_9272,N_9369);
nor U9417 (N_9417,N_9318,N_9213);
nand U9418 (N_9418,N_9366,N_9279);
nand U9419 (N_9419,N_9378,N_9329);
nor U9420 (N_9420,N_9304,N_9217);
nand U9421 (N_9421,N_9312,N_9222);
nor U9422 (N_9422,N_9298,N_9214);
or U9423 (N_9423,N_9203,N_9281);
or U9424 (N_9424,N_9319,N_9373);
nand U9425 (N_9425,N_9349,N_9209);
nor U9426 (N_9426,N_9255,N_9273);
and U9427 (N_9427,N_9293,N_9321);
xor U9428 (N_9428,N_9360,N_9290);
nor U9429 (N_9429,N_9310,N_9242);
nand U9430 (N_9430,N_9345,N_9359);
nand U9431 (N_9431,N_9362,N_9239);
and U9432 (N_9432,N_9243,N_9338);
or U9433 (N_9433,N_9324,N_9330);
or U9434 (N_9434,N_9320,N_9254);
xor U9435 (N_9435,N_9332,N_9325);
or U9436 (N_9436,N_9328,N_9223);
nor U9437 (N_9437,N_9277,N_9201);
xnor U9438 (N_9438,N_9206,N_9234);
nor U9439 (N_9439,N_9331,N_9386);
nor U9440 (N_9440,N_9215,N_9202);
nand U9441 (N_9441,N_9286,N_9380);
and U9442 (N_9442,N_9232,N_9317);
and U9443 (N_9443,N_9398,N_9305);
or U9444 (N_9444,N_9249,N_9307);
or U9445 (N_9445,N_9252,N_9200);
and U9446 (N_9446,N_9308,N_9268);
and U9447 (N_9447,N_9226,N_9231);
or U9448 (N_9448,N_9287,N_9236);
nand U9449 (N_9449,N_9265,N_9397);
or U9450 (N_9450,N_9207,N_9282);
and U9451 (N_9451,N_9356,N_9235);
or U9452 (N_9452,N_9348,N_9211);
and U9453 (N_9453,N_9306,N_9399);
xnor U9454 (N_9454,N_9302,N_9326);
nor U9455 (N_9455,N_9297,N_9288);
nand U9456 (N_9456,N_9253,N_9322);
nand U9457 (N_9457,N_9343,N_9361);
or U9458 (N_9458,N_9382,N_9266);
or U9459 (N_9459,N_9283,N_9344);
or U9460 (N_9460,N_9205,N_9212);
or U9461 (N_9461,N_9368,N_9274);
or U9462 (N_9462,N_9363,N_9246);
nor U9463 (N_9463,N_9354,N_9225);
xor U9464 (N_9464,N_9390,N_9285);
or U9465 (N_9465,N_9327,N_9370);
nand U9466 (N_9466,N_9292,N_9367);
nor U9467 (N_9467,N_9315,N_9262);
or U9468 (N_9468,N_9371,N_9376);
nand U9469 (N_9469,N_9278,N_9221);
nor U9470 (N_9470,N_9240,N_9256);
or U9471 (N_9471,N_9299,N_9392);
nor U9472 (N_9472,N_9377,N_9357);
nand U9473 (N_9473,N_9220,N_9300);
nor U9474 (N_9474,N_9365,N_9340);
xnor U9475 (N_9475,N_9280,N_9391);
nand U9476 (N_9476,N_9383,N_9267);
xor U9477 (N_9477,N_9289,N_9336);
nor U9478 (N_9478,N_9291,N_9337);
and U9479 (N_9479,N_9219,N_9295);
or U9480 (N_9480,N_9388,N_9385);
nor U9481 (N_9481,N_9374,N_9296);
nand U9482 (N_9482,N_9313,N_9347);
xnor U9483 (N_9483,N_9261,N_9333);
nor U9484 (N_9484,N_9334,N_9233);
nor U9485 (N_9485,N_9224,N_9230);
nand U9486 (N_9486,N_9395,N_9204);
nand U9487 (N_9487,N_9389,N_9208);
xor U9488 (N_9488,N_9216,N_9303);
or U9489 (N_9489,N_9309,N_9352);
nor U9490 (N_9490,N_9394,N_9311);
nor U9491 (N_9491,N_9257,N_9276);
xor U9492 (N_9492,N_9247,N_9339);
or U9493 (N_9493,N_9316,N_9264);
nand U9494 (N_9494,N_9381,N_9248);
xor U9495 (N_9495,N_9384,N_9372);
and U9496 (N_9496,N_9353,N_9355);
nor U9497 (N_9497,N_9263,N_9335);
nand U9498 (N_9498,N_9244,N_9210);
and U9499 (N_9499,N_9350,N_9393);
nor U9500 (N_9500,N_9350,N_9324);
or U9501 (N_9501,N_9209,N_9279);
nor U9502 (N_9502,N_9381,N_9396);
nor U9503 (N_9503,N_9362,N_9250);
or U9504 (N_9504,N_9220,N_9370);
nor U9505 (N_9505,N_9325,N_9204);
and U9506 (N_9506,N_9343,N_9385);
xor U9507 (N_9507,N_9293,N_9217);
nand U9508 (N_9508,N_9271,N_9251);
or U9509 (N_9509,N_9326,N_9203);
nand U9510 (N_9510,N_9343,N_9397);
and U9511 (N_9511,N_9253,N_9205);
xnor U9512 (N_9512,N_9268,N_9339);
or U9513 (N_9513,N_9272,N_9222);
nor U9514 (N_9514,N_9311,N_9218);
or U9515 (N_9515,N_9353,N_9314);
or U9516 (N_9516,N_9220,N_9244);
xnor U9517 (N_9517,N_9351,N_9244);
nor U9518 (N_9518,N_9229,N_9266);
and U9519 (N_9519,N_9267,N_9233);
nor U9520 (N_9520,N_9215,N_9253);
nor U9521 (N_9521,N_9254,N_9274);
nand U9522 (N_9522,N_9227,N_9262);
or U9523 (N_9523,N_9323,N_9252);
nand U9524 (N_9524,N_9381,N_9281);
nand U9525 (N_9525,N_9314,N_9369);
and U9526 (N_9526,N_9251,N_9223);
and U9527 (N_9527,N_9240,N_9212);
nand U9528 (N_9528,N_9398,N_9274);
nand U9529 (N_9529,N_9259,N_9359);
or U9530 (N_9530,N_9384,N_9362);
nand U9531 (N_9531,N_9207,N_9369);
nand U9532 (N_9532,N_9264,N_9350);
or U9533 (N_9533,N_9356,N_9301);
xnor U9534 (N_9534,N_9275,N_9238);
or U9535 (N_9535,N_9203,N_9359);
and U9536 (N_9536,N_9212,N_9358);
or U9537 (N_9537,N_9298,N_9353);
nand U9538 (N_9538,N_9272,N_9311);
or U9539 (N_9539,N_9283,N_9210);
nor U9540 (N_9540,N_9217,N_9207);
and U9541 (N_9541,N_9265,N_9384);
nand U9542 (N_9542,N_9270,N_9262);
and U9543 (N_9543,N_9359,N_9289);
xor U9544 (N_9544,N_9380,N_9307);
and U9545 (N_9545,N_9275,N_9210);
nor U9546 (N_9546,N_9230,N_9233);
nor U9547 (N_9547,N_9259,N_9293);
and U9548 (N_9548,N_9200,N_9381);
xor U9549 (N_9549,N_9238,N_9384);
xnor U9550 (N_9550,N_9224,N_9223);
nand U9551 (N_9551,N_9338,N_9390);
and U9552 (N_9552,N_9261,N_9382);
nand U9553 (N_9553,N_9208,N_9200);
and U9554 (N_9554,N_9371,N_9220);
or U9555 (N_9555,N_9343,N_9260);
nand U9556 (N_9556,N_9278,N_9276);
nor U9557 (N_9557,N_9231,N_9378);
and U9558 (N_9558,N_9217,N_9302);
xor U9559 (N_9559,N_9235,N_9337);
nor U9560 (N_9560,N_9264,N_9391);
nor U9561 (N_9561,N_9359,N_9225);
nor U9562 (N_9562,N_9250,N_9326);
nor U9563 (N_9563,N_9347,N_9342);
nand U9564 (N_9564,N_9291,N_9383);
nor U9565 (N_9565,N_9350,N_9360);
and U9566 (N_9566,N_9212,N_9303);
or U9567 (N_9567,N_9391,N_9380);
xnor U9568 (N_9568,N_9218,N_9208);
nand U9569 (N_9569,N_9236,N_9379);
and U9570 (N_9570,N_9398,N_9209);
nand U9571 (N_9571,N_9236,N_9203);
nor U9572 (N_9572,N_9352,N_9397);
nor U9573 (N_9573,N_9356,N_9300);
xor U9574 (N_9574,N_9344,N_9260);
xor U9575 (N_9575,N_9277,N_9213);
and U9576 (N_9576,N_9214,N_9277);
xnor U9577 (N_9577,N_9249,N_9321);
or U9578 (N_9578,N_9355,N_9269);
and U9579 (N_9579,N_9284,N_9246);
nand U9580 (N_9580,N_9276,N_9350);
nand U9581 (N_9581,N_9348,N_9269);
or U9582 (N_9582,N_9399,N_9326);
xor U9583 (N_9583,N_9377,N_9307);
xor U9584 (N_9584,N_9285,N_9215);
or U9585 (N_9585,N_9345,N_9283);
nor U9586 (N_9586,N_9254,N_9203);
nor U9587 (N_9587,N_9247,N_9382);
xnor U9588 (N_9588,N_9257,N_9390);
and U9589 (N_9589,N_9212,N_9354);
and U9590 (N_9590,N_9371,N_9309);
xor U9591 (N_9591,N_9368,N_9382);
or U9592 (N_9592,N_9291,N_9304);
nand U9593 (N_9593,N_9320,N_9376);
xnor U9594 (N_9594,N_9267,N_9255);
and U9595 (N_9595,N_9253,N_9203);
or U9596 (N_9596,N_9216,N_9262);
nand U9597 (N_9597,N_9354,N_9259);
nor U9598 (N_9598,N_9382,N_9272);
or U9599 (N_9599,N_9237,N_9274);
nor U9600 (N_9600,N_9597,N_9464);
or U9601 (N_9601,N_9401,N_9541);
or U9602 (N_9602,N_9492,N_9524);
nand U9603 (N_9603,N_9544,N_9548);
nand U9604 (N_9604,N_9466,N_9414);
xor U9605 (N_9605,N_9483,N_9552);
and U9606 (N_9606,N_9458,N_9519);
nor U9607 (N_9607,N_9495,N_9506);
and U9608 (N_9608,N_9554,N_9557);
xor U9609 (N_9609,N_9550,N_9522);
xor U9610 (N_9610,N_9555,N_9507);
or U9611 (N_9611,N_9460,N_9482);
nand U9612 (N_9612,N_9537,N_9521);
xnor U9613 (N_9613,N_9543,N_9553);
and U9614 (N_9614,N_9535,N_9516);
or U9615 (N_9615,N_9406,N_9534);
nor U9616 (N_9616,N_9569,N_9585);
and U9617 (N_9617,N_9448,N_9476);
or U9618 (N_9618,N_9591,N_9529);
nand U9619 (N_9619,N_9412,N_9434);
and U9620 (N_9620,N_9579,N_9497);
and U9621 (N_9621,N_9598,N_9411);
xor U9622 (N_9622,N_9580,N_9538);
nor U9623 (N_9623,N_9599,N_9423);
and U9624 (N_9624,N_9461,N_9456);
or U9625 (N_9625,N_9446,N_9515);
nand U9626 (N_9626,N_9508,N_9457);
nand U9627 (N_9627,N_9451,N_9571);
and U9628 (N_9628,N_9408,N_9491);
nor U9629 (N_9629,N_9463,N_9518);
xor U9630 (N_9630,N_9481,N_9422);
and U9631 (N_9631,N_9500,N_9590);
nand U9632 (N_9632,N_9566,N_9442);
nand U9633 (N_9633,N_9578,N_9421);
and U9634 (N_9634,N_9440,N_9587);
and U9635 (N_9635,N_9586,N_9489);
nor U9636 (N_9636,N_9472,N_9542);
and U9637 (N_9637,N_9564,N_9570);
nor U9638 (N_9638,N_9416,N_9575);
and U9639 (N_9639,N_9583,N_9558);
nor U9640 (N_9640,N_9437,N_9525);
and U9641 (N_9641,N_9532,N_9576);
xor U9642 (N_9642,N_9478,N_9431);
or U9643 (N_9643,N_9494,N_9447);
and U9644 (N_9644,N_9547,N_9588);
nor U9645 (N_9645,N_9468,N_9484);
nor U9646 (N_9646,N_9454,N_9498);
and U9647 (N_9647,N_9584,N_9403);
xnor U9648 (N_9648,N_9450,N_9505);
nand U9649 (N_9649,N_9574,N_9487);
nand U9650 (N_9650,N_9510,N_9546);
or U9651 (N_9651,N_9477,N_9509);
nand U9652 (N_9652,N_9444,N_9520);
xor U9653 (N_9653,N_9426,N_9471);
nand U9654 (N_9654,N_9514,N_9473);
or U9655 (N_9655,N_9415,N_9479);
and U9656 (N_9656,N_9418,N_9581);
or U9657 (N_9657,N_9503,N_9582);
nor U9658 (N_9658,N_9474,N_9445);
nor U9659 (N_9659,N_9436,N_9493);
nand U9660 (N_9660,N_9462,N_9568);
xnor U9661 (N_9661,N_9592,N_9435);
nand U9662 (N_9662,N_9486,N_9531);
and U9663 (N_9663,N_9428,N_9488);
nor U9664 (N_9664,N_9572,N_9430);
and U9665 (N_9665,N_9545,N_9556);
nor U9666 (N_9666,N_9549,N_9561);
nand U9667 (N_9667,N_9517,N_9528);
or U9668 (N_9668,N_9470,N_9512);
nor U9669 (N_9669,N_9523,N_9596);
xor U9670 (N_9670,N_9432,N_9499);
nand U9671 (N_9671,N_9490,N_9420);
xnor U9672 (N_9672,N_9441,N_9593);
and U9673 (N_9673,N_9527,N_9409);
nor U9674 (N_9674,N_9413,N_9594);
nand U9675 (N_9675,N_9513,N_9565);
or U9676 (N_9676,N_9443,N_9467);
xor U9677 (N_9677,N_9536,N_9407);
xnor U9678 (N_9678,N_9433,N_9540);
nor U9679 (N_9679,N_9539,N_9496);
or U9680 (N_9680,N_9573,N_9425);
xnor U9681 (N_9681,N_9404,N_9589);
nand U9682 (N_9682,N_9502,N_9427);
xor U9683 (N_9683,N_9504,N_9424);
xor U9684 (N_9684,N_9480,N_9449);
and U9685 (N_9685,N_9551,N_9595);
nand U9686 (N_9686,N_9501,N_9455);
or U9687 (N_9687,N_9563,N_9405);
nor U9688 (N_9688,N_9533,N_9562);
and U9689 (N_9689,N_9465,N_9530);
nand U9690 (N_9690,N_9469,N_9567);
nor U9691 (N_9691,N_9400,N_9452);
nor U9692 (N_9692,N_9439,N_9485);
and U9693 (N_9693,N_9402,N_9511);
nand U9694 (N_9694,N_9560,N_9417);
and U9695 (N_9695,N_9577,N_9559);
nand U9696 (N_9696,N_9438,N_9419);
nand U9697 (N_9697,N_9526,N_9453);
nor U9698 (N_9698,N_9459,N_9429);
xor U9699 (N_9699,N_9475,N_9410);
xor U9700 (N_9700,N_9405,N_9478);
or U9701 (N_9701,N_9581,N_9511);
nand U9702 (N_9702,N_9430,N_9497);
and U9703 (N_9703,N_9521,N_9403);
xnor U9704 (N_9704,N_9411,N_9420);
xor U9705 (N_9705,N_9417,N_9425);
xnor U9706 (N_9706,N_9443,N_9510);
nand U9707 (N_9707,N_9432,N_9410);
nand U9708 (N_9708,N_9555,N_9532);
nor U9709 (N_9709,N_9565,N_9465);
nand U9710 (N_9710,N_9571,N_9406);
nand U9711 (N_9711,N_9563,N_9438);
xnor U9712 (N_9712,N_9430,N_9445);
nor U9713 (N_9713,N_9569,N_9581);
nor U9714 (N_9714,N_9527,N_9505);
and U9715 (N_9715,N_9407,N_9458);
xor U9716 (N_9716,N_9475,N_9583);
and U9717 (N_9717,N_9478,N_9544);
xnor U9718 (N_9718,N_9547,N_9554);
or U9719 (N_9719,N_9541,N_9523);
nand U9720 (N_9720,N_9566,N_9401);
xor U9721 (N_9721,N_9482,N_9461);
xor U9722 (N_9722,N_9536,N_9545);
or U9723 (N_9723,N_9593,N_9419);
or U9724 (N_9724,N_9404,N_9498);
and U9725 (N_9725,N_9454,N_9535);
xnor U9726 (N_9726,N_9459,N_9557);
and U9727 (N_9727,N_9581,N_9500);
xnor U9728 (N_9728,N_9434,N_9508);
xnor U9729 (N_9729,N_9474,N_9446);
nand U9730 (N_9730,N_9407,N_9453);
and U9731 (N_9731,N_9476,N_9591);
nor U9732 (N_9732,N_9415,N_9580);
xor U9733 (N_9733,N_9403,N_9518);
nand U9734 (N_9734,N_9555,N_9448);
and U9735 (N_9735,N_9451,N_9569);
nor U9736 (N_9736,N_9482,N_9530);
or U9737 (N_9737,N_9519,N_9589);
nor U9738 (N_9738,N_9548,N_9453);
and U9739 (N_9739,N_9571,N_9594);
nor U9740 (N_9740,N_9511,N_9449);
nor U9741 (N_9741,N_9544,N_9528);
nand U9742 (N_9742,N_9418,N_9422);
or U9743 (N_9743,N_9483,N_9589);
nor U9744 (N_9744,N_9436,N_9503);
nand U9745 (N_9745,N_9482,N_9579);
or U9746 (N_9746,N_9459,N_9424);
or U9747 (N_9747,N_9587,N_9498);
or U9748 (N_9748,N_9425,N_9476);
or U9749 (N_9749,N_9445,N_9570);
nand U9750 (N_9750,N_9400,N_9537);
or U9751 (N_9751,N_9552,N_9515);
or U9752 (N_9752,N_9425,N_9559);
nor U9753 (N_9753,N_9512,N_9555);
nand U9754 (N_9754,N_9586,N_9520);
nor U9755 (N_9755,N_9526,N_9588);
nor U9756 (N_9756,N_9528,N_9412);
nor U9757 (N_9757,N_9414,N_9576);
or U9758 (N_9758,N_9416,N_9405);
or U9759 (N_9759,N_9578,N_9455);
nor U9760 (N_9760,N_9470,N_9432);
nand U9761 (N_9761,N_9440,N_9502);
nor U9762 (N_9762,N_9425,N_9510);
nor U9763 (N_9763,N_9583,N_9446);
and U9764 (N_9764,N_9497,N_9479);
nand U9765 (N_9765,N_9401,N_9424);
nor U9766 (N_9766,N_9555,N_9585);
and U9767 (N_9767,N_9513,N_9413);
xor U9768 (N_9768,N_9592,N_9570);
nand U9769 (N_9769,N_9420,N_9593);
nor U9770 (N_9770,N_9536,N_9570);
xor U9771 (N_9771,N_9548,N_9577);
or U9772 (N_9772,N_9559,N_9548);
nor U9773 (N_9773,N_9430,N_9411);
or U9774 (N_9774,N_9460,N_9501);
nand U9775 (N_9775,N_9584,N_9483);
and U9776 (N_9776,N_9540,N_9487);
or U9777 (N_9777,N_9401,N_9591);
nand U9778 (N_9778,N_9495,N_9597);
nand U9779 (N_9779,N_9560,N_9588);
nand U9780 (N_9780,N_9546,N_9442);
or U9781 (N_9781,N_9519,N_9526);
nor U9782 (N_9782,N_9475,N_9574);
xor U9783 (N_9783,N_9423,N_9456);
nand U9784 (N_9784,N_9529,N_9531);
or U9785 (N_9785,N_9529,N_9419);
or U9786 (N_9786,N_9544,N_9489);
nor U9787 (N_9787,N_9443,N_9522);
nand U9788 (N_9788,N_9444,N_9585);
nand U9789 (N_9789,N_9560,N_9507);
xnor U9790 (N_9790,N_9493,N_9407);
or U9791 (N_9791,N_9578,N_9580);
and U9792 (N_9792,N_9576,N_9403);
or U9793 (N_9793,N_9544,N_9423);
nor U9794 (N_9794,N_9537,N_9565);
xnor U9795 (N_9795,N_9520,N_9547);
or U9796 (N_9796,N_9510,N_9512);
and U9797 (N_9797,N_9589,N_9512);
and U9798 (N_9798,N_9514,N_9587);
or U9799 (N_9799,N_9495,N_9585);
or U9800 (N_9800,N_9640,N_9657);
and U9801 (N_9801,N_9679,N_9623);
and U9802 (N_9802,N_9691,N_9701);
xnor U9803 (N_9803,N_9608,N_9604);
nand U9804 (N_9804,N_9678,N_9743);
and U9805 (N_9805,N_9719,N_9628);
nor U9806 (N_9806,N_9735,N_9603);
xor U9807 (N_9807,N_9690,N_9726);
xnor U9808 (N_9808,N_9655,N_9765);
nor U9809 (N_9809,N_9667,N_9705);
and U9810 (N_9810,N_9716,N_9758);
xnor U9811 (N_9811,N_9774,N_9730);
and U9812 (N_9812,N_9616,N_9759);
xnor U9813 (N_9813,N_9746,N_9748);
xnor U9814 (N_9814,N_9721,N_9698);
and U9815 (N_9815,N_9702,N_9773);
or U9816 (N_9816,N_9652,N_9600);
or U9817 (N_9817,N_9636,N_9669);
nor U9818 (N_9818,N_9674,N_9683);
nand U9819 (N_9819,N_9728,N_9725);
and U9820 (N_9820,N_9644,N_9639);
xnor U9821 (N_9821,N_9777,N_9724);
and U9822 (N_9822,N_9664,N_9607);
or U9823 (N_9823,N_9794,N_9687);
xnor U9824 (N_9824,N_9780,N_9713);
nand U9825 (N_9825,N_9781,N_9693);
nand U9826 (N_9826,N_9629,N_9731);
nor U9827 (N_9827,N_9785,N_9707);
xnor U9828 (N_9828,N_9680,N_9612);
or U9829 (N_9829,N_9676,N_9789);
nor U9830 (N_9830,N_9602,N_9605);
and U9831 (N_9831,N_9761,N_9709);
xnor U9832 (N_9832,N_9771,N_9723);
or U9833 (N_9833,N_9648,N_9764);
or U9834 (N_9834,N_9606,N_9788);
nand U9835 (N_9835,N_9610,N_9654);
or U9836 (N_9836,N_9710,N_9793);
or U9837 (N_9837,N_9729,N_9766);
nand U9838 (N_9838,N_9708,N_9787);
nand U9839 (N_9839,N_9673,N_9626);
xor U9840 (N_9840,N_9663,N_9712);
nor U9841 (N_9841,N_9656,N_9736);
and U9842 (N_9842,N_9700,N_9763);
nor U9843 (N_9843,N_9670,N_9745);
xor U9844 (N_9844,N_9779,N_9768);
nor U9845 (N_9845,N_9692,N_9711);
or U9846 (N_9846,N_9737,N_9618);
or U9847 (N_9847,N_9643,N_9651);
and U9848 (N_9848,N_9634,N_9672);
or U9849 (N_9849,N_9733,N_9689);
xnor U9850 (N_9850,N_9696,N_9699);
nand U9851 (N_9851,N_9666,N_9649);
and U9852 (N_9852,N_9621,N_9795);
nand U9853 (N_9853,N_9675,N_9792);
nand U9854 (N_9854,N_9770,N_9613);
and U9855 (N_9855,N_9631,N_9688);
nor U9856 (N_9856,N_9681,N_9650);
or U9857 (N_9857,N_9601,N_9630);
xor U9858 (N_9858,N_9677,N_9734);
and U9859 (N_9859,N_9704,N_9622);
xor U9860 (N_9860,N_9614,N_9642);
nor U9861 (N_9861,N_9703,N_9744);
and U9862 (N_9862,N_9750,N_9740);
nor U9863 (N_9863,N_9617,N_9717);
or U9864 (N_9864,N_9760,N_9778);
xnor U9865 (N_9865,N_9671,N_9767);
nand U9866 (N_9866,N_9727,N_9624);
nand U9867 (N_9867,N_9751,N_9762);
nand U9868 (N_9868,N_9796,N_9635);
nor U9869 (N_9869,N_9742,N_9738);
xor U9870 (N_9870,N_9753,N_9658);
or U9871 (N_9871,N_9722,N_9769);
nor U9872 (N_9872,N_9637,N_9633);
and U9873 (N_9873,N_9706,N_9638);
nand U9874 (N_9874,N_9732,N_9632);
and U9875 (N_9875,N_9625,N_9697);
or U9876 (N_9876,N_9627,N_9782);
or U9877 (N_9877,N_9695,N_9754);
xor U9878 (N_9878,N_9645,N_9686);
xnor U9879 (N_9879,N_9609,N_9714);
and U9880 (N_9880,N_9718,N_9755);
nor U9881 (N_9881,N_9661,N_9783);
nor U9882 (N_9882,N_9752,N_9662);
or U9883 (N_9883,N_9720,N_9797);
xor U9884 (N_9884,N_9798,N_9659);
nor U9885 (N_9885,N_9619,N_9747);
nand U9886 (N_9886,N_9653,N_9660);
xnor U9887 (N_9887,N_9799,N_9775);
xor U9888 (N_9888,N_9786,N_9685);
nor U9889 (N_9889,N_9641,N_9668);
and U9890 (N_9890,N_9772,N_9749);
or U9891 (N_9891,N_9620,N_9684);
xnor U9892 (N_9892,N_9694,N_9790);
or U9893 (N_9893,N_9647,N_9665);
or U9894 (N_9894,N_9741,N_9757);
xnor U9895 (N_9895,N_9776,N_9756);
or U9896 (N_9896,N_9682,N_9784);
nand U9897 (N_9897,N_9715,N_9739);
nor U9898 (N_9898,N_9611,N_9791);
and U9899 (N_9899,N_9646,N_9615);
xnor U9900 (N_9900,N_9615,N_9730);
xnor U9901 (N_9901,N_9610,N_9603);
nand U9902 (N_9902,N_9691,N_9779);
nor U9903 (N_9903,N_9628,N_9786);
nor U9904 (N_9904,N_9720,N_9712);
and U9905 (N_9905,N_9737,N_9662);
or U9906 (N_9906,N_9628,N_9751);
or U9907 (N_9907,N_9733,N_9741);
nand U9908 (N_9908,N_9613,N_9750);
xor U9909 (N_9909,N_9767,N_9685);
nor U9910 (N_9910,N_9728,N_9739);
nor U9911 (N_9911,N_9661,N_9769);
nand U9912 (N_9912,N_9704,N_9620);
nand U9913 (N_9913,N_9713,N_9746);
and U9914 (N_9914,N_9763,N_9760);
and U9915 (N_9915,N_9694,N_9704);
or U9916 (N_9916,N_9652,N_9777);
nand U9917 (N_9917,N_9664,N_9703);
and U9918 (N_9918,N_9739,N_9648);
xnor U9919 (N_9919,N_9760,N_9701);
nor U9920 (N_9920,N_9614,N_9693);
nand U9921 (N_9921,N_9778,N_9736);
nor U9922 (N_9922,N_9669,N_9790);
nor U9923 (N_9923,N_9646,N_9683);
nor U9924 (N_9924,N_9672,N_9679);
nor U9925 (N_9925,N_9659,N_9721);
nor U9926 (N_9926,N_9789,N_9608);
xor U9927 (N_9927,N_9613,N_9691);
xnor U9928 (N_9928,N_9696,N_9704);
and U9929 (N_9929,N_9740,N_9667);
or U9930 (N_9930,N_9785,N_9601);
and U9931 (N_9931,N_9790,N_9671);
or U9932 (N_9932,N_9654,N_9705);
nor U9933 (N_9933,N_9623,N_9695);
nor U9934 (N_9934,N_9667,N_9607);
xnor U9935 (N_9935,N_9651,N_9744);
or U9936 (N_9936,N_9709,N_9715);
xnor U9937 (N_9937,N_9647,N_9782);
or U9938 (N_9938,N_9743,N_9642);
nand U9939 (N_9939,N_9692,N_9623);
or U9940 (N_9940,N_9648,N_9797);
nor U9941 (N_9941,N_9608,N_9660);
nor U9942 (N_9942,N_9600,N_9617);
and U9943 (N_9943,N_9684,N_9791);
nor U9944 (N_9944,N_9756,N_9760);
xnor U9945 (N_9945,N_9699,N_9698);
xor U9946 (N_9946,N_9619,N_9620);
nor U9947 (N_9947,N_9637,N_9736);
xnor U9948 (N_9948,N_9640,N_9623);
nor U9949 (N_9949,N_9644,N_9760);
nand U9950 (N_9950,N_9646,N_9798);
or U9951 (N_9951,N_9624,N_9614);
nor U9952 (N_9952,N_9786,N_9627);
or U9953 (N_9953,N_9708,N_9795);
nor U9954 (N_9954,N_9773,N_9701);
and U9955 (N_9955,N_9706,N_9614);
nor U9956 (N_9956,N_9728,N_9752);
and U9957 (N_9957,N_9674,N_9789);
and U9958 (N_9958,N_9674,N_9601);
and U9959 (N_9959,N_9691,N_9644);
or U9960 (N_9960,N_9787,N_9629);
or U9961 (N_9961,N_9643,N_9645);
and U9962 (N_9962,N_9798,N_9720);
or U9963 (N_9963,N_9628,N_9644);
xor U9964 (N_9964,N_9721,N_9715);
and U9965 (N_9965,N_9789,N_9752);
nor U9966 (N_9966,N_9717,N_9671);
and U9967 (N_9967,N_9640,N_9731);
and U9968 (N_9968,N_9734,N_9676);
xor U9969 (N_9969,N_9692,N_9701);
or U9970 (N_9970,N_9714,N_9612);
nor U9971 (N_9971,N_9643,N_9751);
nand U9972 (N_9972,N_9782,N_9700);
or U9973 (N_9973,N_9790,N_9770);
xnor U9974 (N_9974,N_9785,N_9715);
xnor U9975 (N_9975,N_9604,N_9744);
nand U9976 (N_9976,N_9762,N_9634);
nand U9977 (N_9977,N_9730,N_9736);
and U9978 (N_9978,N_9647,N_9646);
or U9979 (N_9979,N_9725,N_9696);
xnor U9980 (N_9980,N_9795,N_9692);
or U9981 (N_9981,N_9610,N_9622);
nand U9982 (N_9982,N_9639,N_9683);
nor U9983 (N_9983,N_9712,N_9691);
xnor U9984 (N_9984,N_9704,N_9638);
nand U9985 (N_9985,N_9782,N_9744);
nor U9986 (N_9986,N_9773,N_9727);
or U9987 (N_9987,N_9639,N_9736);
xor U9988 (N_9988,N_9782,N_9613);
nand U9989 (N_9989,N_9600,N_9692);
nor U9990 (N_9990,N_9655,N_9733);
and U9991 (N_9991,N_9601,N_9656);
nand U9992 (N_9992,N_9645,N_9630);
nor U9993 (N_9993,N_9788,N_9730);
nand U9994 (N_9994,N_9634,N_9643);
nand U9995 (N_9995,N_9779,N_9631);
nand U9996 (N_9996,N_9610,N_9737);
or U9997 (N_9997,N_9694,N_9716);
xor U9998 (N_9998,N_9777,N_9720);
or U9999 (N_9999,N_9691,N_9678);
xor U10000 (N_10000,N_9954,N_9911);
xor U10001 (N_10001,N_9958,N_9840);
nor U10002 (N_10002,N_9968,N_9845);
nand U10003 (N_10003,N_9921,N_9945);
xor U10004 (N_10004,N_9849,N_9878);
and U10005 (N_10005,N_9905,N_9983);
nor U10006 (N_10006,N_9961,N_9836);
and U10007 (N_10007,N_9986,N_9811);
xor U10008 (N_10008,N_9967,N_9852);
and U10009 (N_10009,N_9874,N_9949);
xor U10010 (N_10010,N_9926,N_9941);
nor U10011 (N_10011,N_9864,N_9832);
nand U10012 (N_10012,N_9936,N_9956);
or U10013 (N_10013,N_9960,N_9896);
nor U10014 (N_10014,N_9819,N_9964);
nand U10015 (N_10015,N_9947,N_9839);
nand U10016 (N_10016,N_9856,N_9870);
and U10017 (N_10017,N_9969,N_9813);
nand U10018 (N_10018,N_9898,N_9950);
or U10019 (N_10019,N_9831,N_9837);
xor U10020 (N_10020,N_9952,N_9901);
or U10021 (N_10021,N_9999,N_9988);
nand U10022 (N_10022,N_9903,N_9929);
nand U10023 (N_10023,N_9822,N_9809);
xnor U10024 (N_10024,N_9843,N_9902);
and U10025 (N_10025,N_9972,N_9859);
nand U10026 (N_10026,N_9815,N_9821);
and U10027 (N_10027,N_9881,N_9865);
nor U10028 (N_10028,N_9890,N_9873);
nor U10029 (N_10029,N_9982,N_9869);
nor U10030 (N_10030,N_9900,N_9934);
nand U10031 (N_10031,N_9848,N_9804);
xnor U10032 (N_10032,N_9820,N_9993);
nor U10033 (N_10033,N_9998,N_9933);
nand U10034 (N_10034,N_9876,N_9860);
or U10035 (N_10035,N_9883,N_9892);
and U10036 (N_10036,N_9885,N_9816);
xor U10037 (N_10037,N_9979,N_9850);
or U10038 (N_10038,N_9817,N_9974);
and U10039 (N_10039,N_9909,N_9955);
nand U10040 (N_10040,N_9833,N_9942);
xnor U10041 (N_10041,N_9824,N_9830);
nor U10042 (N_10042,N_9946,N_9910);
and U10043 (N_10043,N_9897,N_9919);
or U10044 (N_10044,N_9932,N_9925);
xnor U10045 (N_10045,N_9963,N_9802);
xor U10046 (N_10046,N_9912,N_9884);
nor U10047 (N_10047,N_9858,N_9818);
nor U10048 (N_10048,N_9827,N_9880);
nand U10049 (N_10049,N_9846,N_9842);
nand U10050 (N_10050,N_9977,N_9978);
and U10051 (N_10051,N_9914,N_9940);
nand U10052 (N_10052,N_9997,N_9957);
and U10053 (N_10053,N_9971,N_9981);
or U10054 (N_10054,N_9801,N_9992);
and U10055 (N_10055,N_9800,N_9995);
or U10056 (N_10056,N_9829,N_9810);
xnor U10057 (N_10057,N_9991,N_9862);
or U10058 (N_10058,N_9923,N_9906);
xnor U10059 (N_10059,N_9990,N_9803);
xor U10060 (N_10060,N_9828,N_9807);
nand U10061 (N_10061,N_9844,N_9826);
and U10062 (N_10062,N_9891,N_9908);
nand U10063 (N_10063,N_9847,N_9976);
and U10064 (N_10064,N_9944,N_9835);
and U10065 (N_10065,N_9989,N_9938);
xor U10066 (N_10066,N_9966,N_9994);
nor U10067 (N_10067,N_9868,N_9975);
nor U10068 (N_10068,N_9922,N_9984);
nand U10069 (N_10069,N_9882,N_9920);
xor U10070 (N_10070,N_9965,N_9853);
xnor U10071 (N_10071,N_9834,N_9943);
xnor U10072 (N_10072,N_9894,N_9893);
xor U10073 (N_10073,N_9875,N_9899);
nor U10074 (N_10074,N_9915,N_9889);
xnor U10075 (N_10075,N_9838,N_9866);
nand U10076 (N_10076,N_9805,N_9857);
nand U10077 (N_10077,N_9867,N_9886);
xor U10078 (N_10078,N_9888,N_9927);
or U10079 (N_10079,N_9987,N_9962);
or U10080 (N_10080,N_9855,N_9973);
nand U10081 (N_10081,N_9935,N_9872);
nand U10082 (N_10082,N_9931,N_9895);
xor U10083 (N_10083,N_9823,N_9996);
and U10084 (N_10084,N_9854,N_9871);
xor U10085 (N_10085,N_9863,N_9861);
and U10086 (N_10086,N_9851,N_9913);
and U10087 (N_10087,N_9937,N_9928);
or U10088 (N_10088,N_9924,N_9904);
or U10089 (N_10089,N_9959,N_9985);
and U10090 (N_10090,N_9877,N_9948);
and U10091 (N_10091,N_9814,N_9812);
and U10092 (N_10092,N_9939,N_9970);
or U10093 (N_10093,N_9951,N_9953);
nor U10094 (N_10094,N_9841,N_9916);
xor U10095 (N_10095,N_9879,N_9887);
nor U10096 (N_10096,N_9930,N_9825);
nor U10097 (N_10097,N_9806,N_9918);
xnor U10098 (N_10098,N_9980,N_9907);
nand U10099 (N_10099,N_9917,N_9808);
or U10100 (N_10100,N_9841,N_9869);
or U10101 (N_10101,N_9877,N_9924);
nand U10102 (N_10102,N_9866,N_9835);
nor U10103 (N_10103,N_9985,N_9848);
nor U10104 (N_10104,N_9980,N_9852);
and U10105 (N_10105,N_9983,N_9908);
or U10106 (N_10106,N_9867,N_9949);
or U10107 (N_10107,N_9808,N_9872);
xnor U10108 (N_10108,N_9973,N_9857);
xor U10109 (N_10109,N_9974,N_9890);
nand U10110 (N_10110,N_9851,N_9837);
xnor U10111 (N_10111,N_9930,N_9946);
nor U10112 (N_10112,N_9926,N_9976);
or U10113 (N_10113,N_9823,N_9887);
nor U10114 (N_10114,N_9805,N_9947);
nor U10115 (N_10115,N_9827,N_9926);
nand U10116 (N_10116,N_9875,N_9921);
and U10117 (N_10117,N_9871,N_9977);
nor U10118 (N_10118,N_9870,N_9992);
nor U10119 (N_10119,N_9800,N_9979);
xor U10120 (N_10120,N_9875,N_9808);
nand U10121 (N_10121,N_9894,N_9829);
or U10122 (N_10122,N_9858,N_9894);
or U10123 (N_10123,N_9872,N_9835);
xor U10124 (N_10124,N_9962,N_9863);
xor U10125 (N_10125,N_9865,N_9912);
xor U10126 (N_10126,N_9817,N_9863);
and U10127 (N_10127,N_9800,N_9842);
nor U10128 (N_10128,N_9880,N_9894);
and U10129 (N_10129,N_9824,N_9823);
nor U10130 (N_10130,N_9997,N_9898);
nor U10131 (N_10131,N_9897,N_9834);
or U10132 (N_10132,N_9829,N_9832);
or U10133 (N_10133,N_9877,N_9854);
nor U10134 (N_10134,N_9946,N_9885);
nor U10135 (N_10135,N_9922,N_9909);
or U10136 (N_10136,N_9908,N_9996);
nand U10137 (N_10137,N_9889,N_9840);
xor U10138 (N_10138,N_9828,N_9900);
or U10139 (N_10139,N_9978,N_9994);
nand U10140 (N_10140,N_9941,N_9822);
xnor U10141 (N_10141,N_9868,N_9976);
and U10142 (N_10142,N_9848,N_9815);
or U10143 (N_10143,N_9884,N_9983);
and U10144 (N_10144,N_9826,N_9966);
xnor U10145 (N_10145,N_9822,N_9827);
and U10146 (N_10146,N_9974,N_9887);
nor U10147 (N_10147,N_9870,N_9827);
xor U10148 (N_10148,N_9814,N_9816);
nand U10149 (N_10149,N_9812,N_9903);
and U10150 (N_10150,N_9885,N_9995);
nor U10151 (N_10151,N_9873,N_9845);
nand U10152 (N_10152,N_9899,N_9814);
and U10153 (N_10153,N_9953,N_9843);
xor U10154 (N_10154,N_9831,N_9990);
and U10155 (N_10155,N_9807,N_9944);
and U10156 (N_10156,N_9889,N_9973);
or U10157 (N_10157,N_9956,N_9900);
and U10158 (N_10158,N_9979,N_9996);
xnor U10159 (N_10159,N_9865,N_9990);
and U10160 (N_10160,N_9959,N_9856);
xor U10161 (N_10161,N_9963,N_9859);
xnor U10162 (N_10162,N_9959,N_9813);
xor U10163 (N_10163,N_9820,N_9911);
or U10164 (N_10164,N_9996,N_9835);
xor U10165 (N_10165,N_9882,N_9899);
xnor U10166 (N_10166,N_9848,N_9991);
xor U10167 (N_10167,N_9852,N_9853);
or U10168 (N_10168,N_9994,N_9951);
nand U10169 (N_10169,N_9962,N_9940);
xnor U10170 (N_10170,N_9922,N_9973);
nand U10171 (N_10171,N_9832,N_9850);
or U10172 (N_10172,N_9909,N_9835);
or U10173 (N_10173,N_9991,N_9910);
or U10174 (N_10174,N_9934,N_9820);
nand U10175 (N_10175,N_9872,N_9893);
and U10176 (N_10176,N_9999,N_9928);
and U10177 (N_10177,N_9984,N_9997);
nand U10178 (N_10178,N_9824,N_9997);
xor U10179 (N_10179,N_9840,N_9861);
nand U10180 (N_10180,N_9956,N_9862);
and U10181 (N_10181,N_9898,N_9923);
nor U10182 (N_10182,N_9835,N_9991);
and U10183 (N_10183,N_9815,N_9914);
nand U10184 (N_10184,N_9990,N_9946);
nand U10185 (N_10185,N_9871,N_9900);
or U10186 (N_10186,N_9804,N_9879);
nor U10187 (N_10187,N_9984,N_9819);
or U10188 (N_10188,N_9846,N_9905);
xnor U10189 (N_10189,N_9803,N_9880);
xor U10190 (N_10190,N_9868,N_9894);
and U10191 (N_10191,N_9829,N_9809);
xnor U10192 (N_10192,N_9834,N_9951);
nand U10193 (N_10193,N_9914,N_9875);
nor U10194 (N_10194,N_9831,N_9857);
or U10195 (N_10195,N_9962,N_9856);
nor U10196 (N_10196,N_9866,N_9937);
and U10197 (N_10197,N_9836,N_9837);
xnor U10198 (N_10198,N_9887,N_9848);
or U10199 (N_10199,N_9896,N_9806);
nand U10200 (N_10200,N_10150,N_10011);
nor U10201 (N_10201,N_10023,N_10051);
or U10202 (N_10202,N_10151,N_10009);
or U10203 (N_10203,N_10123,N_10162);
or U10204 (N_10204,N_10040,N_10153);
or U10205 (N_10205,N_10148,N_10056);
and U10206 (N_10206,N_10144,N_10013);
nor U10207 (N_10207,N_10098,N_10160);
and U10208 (N_10208,N_10124,N_10036);
nand U10209 (N_10209,N_10152,N_10087);
nand U10210 (N_10210,N_10057,N_10169);
nand U10211 (N_10211,N_10074,N_10165);
and U10212 (N_10212,N_10164,N_10018);
xor U10213 (N_10213,N_10022,N_10194);
or U10214 (N_10214,N_10037,N_10048);
xnor U10215 (N_10215,N_10067,N_10174);
or U10216 (N_10216,N_10155,N_10167);
or U10217 (N_10217,N_10100,N_10039);
xor U10218 (N_10218,N_10116,N_10103);
xor U10219 (N_10219,N_10111,N_10091);
nand U10220 (N_10220,N_10170,N_10089);
nor U10221 (N_10221,N_10000,N_10072);
xnor U10222 (N_10222,N_10185,N_10093);
or U10223 (N_10223,N_10120,N_10137);
nand U10224 (N_10224,N_10115,N_10119);
and U10225 (N_10225,N_10135,N_10017);
xor U10226 (N_10226,N_10118,N_10154);
nand U10227 (N_10227,N_10158,N_10113);
nand U10228 (N_10228,N_10092,N_10055);
nor U10229 (N_10229,N_10075,N_10001);
nor U10230 (N_10230,N_10028,N_10142);
xor U10231 (N_10231,N_10102,N_10140);
nand U10232 (N_10232,N_10041,N_10108);
nor U10233 (N_10233,N_10126,N_10043);
or U10234 (N_10234,N_10003,N_10157);
or U10235 (N_10235,N_10012,N_10081);
xnor U10236 (N_10236,N_10183,N_10010);
or U10237 (N_10237,N_10020,N_10026);
nand U10238 (N_10238,N_10143,N_10014);
and U10239 (N_10239,N_10184,N_10095);
and U10240 (N_10240,N_10065,N_10050);
or U10241 (N_10241,N_10085,N_10172);
nor U10242 (N_10242,N_10016,N_10044);
nand U10243 (N_10243,N_10063,N_10180);
nand U10244 (N_10244,N_10117,N_10181);
and U10245 (N_10245,N_10161,N_10145);
xnor U10246 (N_10246,N_10090,N_10045);
xor U10247 (N_10247,N_10035,N_10064);
nand U10248 (N_10248,N_10199,N_10175);
nor U10249 (N_10249,N_10068,N_10008);
xor U10250 (N_10250,N_10192,N_10066);
nand U10251 (N_10251,N_10127,N_10071);
or U10252 (N_10252,N_10019,N_10038);
nand U10253 (N_10253,N_10107,N_10080);
and U10254 (N_10254,N_10134,N_10076);
or U10255 (N_10255,N_10131,N_10125);
or U10256 (N_10256,N_10032,N_10176);
and U10257 (N_10257,N_10191,N_10128);
nor U10258 (N_10258,N_10015,N_10178);
or U10259 (N_10259,N_10189,N_10030);
and U10260 (N_10260,N_10079,N_10069);
and U10261 (N_10261,N_10059,N_10197);
nor U10262 (N_10262,N_10198,N_10195);
and U10263 (N_10263,N_10182,N_10073);
nand U10264 (N_10264,N_10130,N_10086);
nor U10265 (N_10265,N_10058,N_10112);
and U10266 (N_10266,N_10168,N_10042);
nand U10267 (N_10267,N_10196,N_10141);
or U10268 (N_10268,N_10005,N_10149);
nand U10269 (N_10269,N_10159,N_10177);
nor U10270 (N_10270,N_10054,N_10024);
xor U10271 (N_10271,N_10156,N_10088);
nand U10272 (N_10272,N_10046,N_10139);
nor U10273 (N_10273,N_10094,N_10002);
and U10274 (N_10274,N_10060,N_10193);
or U10275 (N_10275,N_10105,N_10007);
and U10276 (N_10276,N_10188,N_10033);
xor U10277 (N_10277,N_10138,N_10077);
and U10278 (N_10278,N_10083,N_10179);
nand U10279 (N_10279,N_10146,N_10096);
and U10280 (N_10280,N_10166,N_10122);
nand U10281 (N_10281,N_10027,N_10047);
nand U10282 (N_10282,N_10099,N_10171);
or U10283 (N_10283,N_10129,N_10006);
nand U10284 (N_10284,N_10121,N_10029);
nand U10285 (N_10285,N_10004,N_10052);
xnor U10286 (N_10286,N_10132,N_10021);
xnor U10287 (N_10287,N_10136,N_10053);
nand U10288 (N_10288,N_10104,N_10163);
and U10289 (N_10289,N_10084,N_10173);
and U10290 (N_10290,N_10187,N_10031);
and U10291 (N_10291,N_10147,N_10025);
nor U10292 (N_10292,N_10061,N_10078);
nand U10293 (N_10293,N_10101,N_10062);
nand U10294 (N_10294,N_10190,N_10110);
or U10295 (N_10295,N_10133,N_10186);
and U10296 (N_10296,N_10109,N_10106);
or U10297 (N_10297,N_10070,N_10034);
xnor U10298 (N_10298,N_10114,N_10082);
nand U10299 (N_10299,N_10049,N_10097);
nand U10300 (N_10300,N_10148,N_10094);
and U10301 (N_10301,N_10084,N_10183);
nor U10302 (N_10302,N_10094,N_10007);
nor U10303 (N_10303,N_10142,N_10151);
xnor U10304 (N_10304,N_10119,N_10110);
nor U10305 (N_10305,N_10130,N_10136);
and U10306 (N_10306,N_10042,N_10072);
or U10307 (N_10307,N_10175,N_10017);
and U10308 (N_10308,N_10183,N_10059);
nand U10309 (N_10309,N_10196,N_10135);
nand U10310 (N_10310,N_10024,N_10139);
xor U10311 (N_10311,N_10100,N_10015);
nand U10312 (N_10312,N_10071,N_10164);
nand U10313 (N_10313,N_10185,N_10169);
or U10314 (N_10314,N_10156,N_10155);
nor U10315 (N_10315,N_10064,N_10106);
or U10316 (N_10316,N_10044,N_10137);
xor U10317 (N_10317,N_10033,N_10193);
nor U10318 (N_10318,N_10086,N_10031);
or U10319 (N_10319,N_10188,N_10110);
and U10320 (N_10320,N_10009,N_10083);
and U10321 (N_10321,N_10193,N_10102);
nor U10322 (N_10322,N_10161,N_10166);
nand U10323 (N_10323,N_10096,N_10132);
nand U10324 (N_10324,N_10198,N_10016);
nor U10325 (N_10325,N_10156,N_10153);
nand U10326 (N_10326,N_10159,N_10196);
nand U10327 (N_10327,N_10083,N_10080);
nand U10328 (N_10328,N_10133,N_10196);
nor U10329 (N_10329,N_10125,N_10048);
nand U10330 (N_10330,N_10110,N_10065);
xor U10331 (N_10331,N_10191,N_10028);
nor U10332 (N_10332,N_10130,N_10013);
and U10333 (N_10333,N_10116,N_10085);
or U10334 (N_10334,N_10018,N_10076);
and U10335 (N_10335,N_10171,N_10081);
xor U10336 (N_10336,N_10193,N_10079);
nand U10337 (N_10337,N_10075,N_10049);
nand U10338 (N_10338,N_10164,N_10056);
xor U10339 (N_10339,N_10138,N_10037);
or U10340 (N_10340,N_10024,N_10000);
nand U10341 (N_10341,N_10099,N_10170);
nor U10342 (N_10342,N_10015,N_10071);
xor U10343 (N_10343,N_10079,N_10162);
nand U10344 (N_10344,N_10127,N_10021);
or U10345 (N_10345,N_10116,N_10000);
or U10346 (N_10346,N_10131,N_10069);
or U10347 (N_10347,N_10087,N_10175);
xnor U10348 (N_10348,N_10058,N_10168);
xor U10349 (N_10349,N_10195,N_10187);
nor U10350 (N_10350,N_10059,N_10055);
nand U10351 (N_10351,N_10138,N_10072);
and U10352 (N_10352,N_10179,N_10060);
nand U10353 (N_10353,N_10187,N_10120);
and U10354 (N_10354,N_10167,N_10050);
xnor U10355 (N_10355,N_10112,N_10120);
nor U10356 (N_10356,N_10046,N_10066);
nor U10357 (N_10357,N_10083,N_10094);
nand U10358 (N_10358,N_10199,N_10039);
or U10359 (N_10359,N_10144,N_10082);
nor U10360 (N_10360,N_10175,N_10144);
or U10361 (N_10361,N_10111,N_10052);
xnor U10362 (N_10362,N_10193,N_10025);
xor U10363 (N_10363,N_10136,N_10158);
nor U10364 (N_10364,N_10194,N_10066);
nand U10365 (N_10365,N_10181,N_10172);
nand U10366 (N_10366,N_10058,N_10030);
nor U10367 (N_10367,N_10063,N_10064);
nor U10368 (N_10368,N_10087,N_10104);
nand U10369 (N_10369,N_10008,N_10167);
xor U10370 (N_10370,N_10059,N_10177);
nand U10371 (N_10371,N_10087,N_10027);
nor U10372 (N_10372,N_10128,N_10015);
nor U10373 (N_10373,N_10117,N_10118);
nor U10374 (N_10374,N_10158,N_10090);
or U10375 (N_10375,N_10087,N_10166);
xnor U10376 (N_10376,N_10170,N_10135);
nor U10377 (N_10377,N_10187,N_10041);
and U10378 (N_10378,N_10097,N_10144);
and U10379 (N_10379,N_10116,N_10119);
xor U10380 (N_10380,N_10085,N_10060);
or U10381 (N_10381,N_10086,N_10005);
xor U10382 (N_10382,N_10090,N_10182);
nand U10383 (N_10383,N_10059,N_10134);
or U10384 (N_10384,N_10016,N_10177);
xor U10385 (N_10385,N_10126,N_10159);
xnor U10386 (N_10386,N_10085,N_10177);
nor U10387 (N_10387,N_10067,N_10176);
or U10388 (N_10388,N_10093,N_10101);
nor U10389 (N_10389,N_10103,N_10060);
xnor U10390 (N_10390,N_10107,N_10028);
nor U10391 (N_10391,N_10169,N_10112);
xor U10392 (N_10392,N_10128,N_10145);
nor U10393 (N_10393,N_10198,N_10111);
and U10394 (N_10394,N_10107,N_10032);
xor U10395 (N_10395,N_10118,N_10151);
and U10396 (N_10396,N_10076,N_10017);
or U10397 (N_10397,N_10137,N_10047);
or U10398 (N_10398,N_10048,N_10035);
nand U10399 (N_10399,N_10031,N_10074);
xnor U10400 (N_10400,N_10387,N_10271);
nor U10401 (N_10401,N_10352,N_10338);
nand U10402 (N_10402,N_10312,N_10249);
and U10403 (N_10403,N_10268,N_10320);
and U10404 (N_10404,N_10398,N_10305);
nor U10405 (N_10405,N_10212,N_10301);
xnor U10406 (N_10406,N_10319,N_10358);
nor U10407 (N_10407,N_10306,N_10228);
xor U10408 (N_10408,N_10347,N_10293);
xnor U10409 (N_10409,N_10351,N_10214);
nand U10410 (N_10410,N_10295,N_10394);
nor U10411 (N_10411,N_10201,N_10231);
and U10412 (N_10412,N_10204,N_10390);
nor U10413 (N_10413,N_10370,N_10247);
xnor U10414 (N_10414,N_10380,N_10286);
or U10415 (N_10415,N_10266,N_10297);
xnor U10416 (N_10416,N_10276,N_10343);
or U10417 (N_10417,N_10315,N_10246);
nor U10418 (N_10418,N_10291,N_10300);
or U10419 (N_10419,N_10244,N_10267);
or U10420 (N_10420,N_10375,N_10367);
or U10421 (N_10421,N_10225,N_10374);
nor U10422 (N_10422,N_10296,N_10383);
nor U10423 (N_10423,N_10357,N_10368);
nor U10424 (N_10424,N_10308,N_10275);
or U10425 (N_10425,N_10200,N_10285);
nand U10426 (N_10426,N_10336,N_10299);
or U10427 (N_10427,N_10226,N_10316);
and U10428 (N_10428,N_10251,N_10393);
xor U10429 (N_10429,N_10223,N_10208);
nand U10430 (N_10430,N_10314,N_10344);
xor U10431 (N_10431,N_10389,N_10211);
nand U10432 (N_10432,N_10378,N_10274);
nand U10433 (N_10433,N_10265,N_10205);
nor U10434 (N_10434,N_10233,N_10288);
nand U10435 (N_10435,N_10245,N_10258);
nor U10436 (N_10436,N_10363,N_10340);
nand U10437 (N_10437,N_10310,N_10294);
xnor U10438 (N_10438,N_10303,N_10302);
nor U10439 (N_10439,N_10345,N_10253);
and U10440 (N_10440,N_10287,N_10384);
or U10441 (N_10441,N_10215,N_10221);
xnor U10442 (N_10442,N_10323,N_10262);
nand U10443 (N_10443,N_10210,N_10330);
and U10444 (N_10444,N_10272,N_10346);
nand U10445 (N_10445,N_10356,N_10348);
xor U10446 (N_10446,N_10385,N_10333);
and U10447 (N_10447,N_10342,N_10373);
xor U10448 (N_10448,N_10311,N_10202);
xor U10449 (N_10449,N_10304,N_10326);
and U10450 (N_10450,N_10354,N_10239);
or U10451 (N_10451,N_10219,N_10361);
and U10452 (N_10452,N_10207,N_10256);
xnor U10453 (N_10453,N_10213,N_10222);
and U10454 (N_10454,N_10282,N_10334);
xnor U10455 (N_10455,N_10335,N_10209);
xor U10456 (N_10456,N_10331,N_10386);
nand U10457 (N_10457,N_10376,N_10349);
and U10458 (N_10458,N_10366,N_10328);
nor U10459 (N_10459,N_10355,N_10360);
and U10460 (N_10460,N_10259,N_10322);
and U10461 (N_10461,N_10261,N_10254);
and U10462 (N_10462,N_10283,N_10317);
and U10463 (N_10463,N_10250,N_10281);
and U10464 (N_10464,N_10290,N_10318);
and U10465 (N_10465,N_10381,N_10224);
and U10466 (N_10466,N_10203,N_10269);
and U10467 (N_10467,N_10371,N_10298);
or U10468 (N_10468,N_10332,N_10257);
nor U10469 (N_10469,N_10327,N_10397);
and U10470 (N_10470,N_10240,N_10284);
nor U10471 (N_10471,N_10237,N_10217);
nor U10472 (N_10472,N_10395,N_10350);
nor U10473 (N_10473,N_10216,N_10292);
and U10474 (N_10474,N_10218,N_10242);
nor U10475 (N_10475,N_10365,N_10382);
nor U10476 (N_10476,N_10372,N_10307);
nand U10477 (N_10477,N_10206,N_10341);
or U10478 (N_10478,N_10377,N_10353);
xnor U10479 (N_10479,N_10362,N_10309);
or U10480 (N_10480,N_10235,N_10324);
nand U10481 (N_10481,N_10229,N_10391);
xnor U10482 (N_10482,N_10238,N_10255);
or U10483 (N_10483,N_10264,N_10329);
or U10484 (N_10484,N_10289,N_10399);
or U10485 (N_10485,N_10359,N_10273);
nand U10486 (N_10486,N_10227,N_10220);
or U10487 (N_10487,N_10278,N_10277);
nand U10488 (N_10488,N_10234,N_10388);
or U10489 (N_10489,N_10396,N_10236);
and U10490 (N_10490,N_10392,N_10325);
nand U10491 (N_10491,N_10260,N_10280);
xnor U10492 (N_10492,N_10263,N_10364);
and U10493 (N_10493,N_10230,N_10243);
nand U10494 (N_10494,N_10241,N_10313);
and U10495 (N_10495,N_10321,N_10339);
or U10496 (N_10496,N_10337,N_10379);
or U10497 (N_10497,N_10232,N_10270);
and U10498 (N_10498,N_10279,N_10252);
xnor U10499 (N_10499,N_10369,N_10248);
and U10500 (N_10500,N_10387,N_10218);
and U10501 (N_10501,N_10382,N_10235);
xnor U10502 (N_10502,N_10340,N_10383);
and U10503 (N_10503,N_10287,N_10266);
or U10504 (N_10504,N_10398,N_10266);
and U10505 (N_10505,N_10258,N_10388);
nand U10506 (N_10506,N_10271,N_10394);
or U10507 (N_10507,N_10221,N_10203);
and U10508 (N_10508,N_10396,N_10344);
nand U10509 (N_10509,N_10251,N_10240);
nand U10510 (N_10510,N_10300,N_10327);
xnor U10511 (N_10511,N_10242,N_10344);
or U10512 (N_10512,N_10330,N_10225);
nand U10513 (N_10513,N_10216,N_10323);
and U10514 (N_10514,N_10324,N_10213);
xor U10515 (N_10515,N_10251,N_10241);
and U10516 (N_10516,N_10388,N_10327);
xor U10517 (N_10517,N_10243,N_10237);
nor U10518 (N_10518,N_10261,N_10303);
nand U10519 (N_10519,N_10247,N_10267);
or U10520 (N_10520,N_10266,N_10250);
and U10521 (N_10521,N_10338,N_10207);
xnor U10522 (N_10522,N_10385,N_10328);
xor U10523 (N_10523,N_10396,N_10276);
nor U10524 (N_10524,N_10250,N_10230);
nor U10525 (N_10525,N_10344,N_10302);
nor U10526 (N_10526,N_10333,N_10232);
or U10527 (N_10527,N_10310,N_10223);
xor U10528 (N_10528,N_10257,N_10341);
or U10529 (N_10529,N_10284,N_10304);
and U10530 (N_10530,N_10250,N_10359);
or U10531 (N_10531,N_10267,N_10256);
and U10532 (N_10532,N_10280,N_10202);
and U10533 (N_10533,N_10394,N_10392);
and U10534 (N_10534,N_10275,N_10364);
xnor U10535 (N_10535,N_10320,N_10226);
and U10536 (N_10536,N_10255,N_10285);
and U10537 (N_10537,N_10230,N_10275);
nand U10538 (N_10538,N_10301,N_10222);
or U10539 (N_10539,N_10357,N_10248);
and U10540 (N_10540,N_10384,N_10364);
xnor U10541 (N_10541,N_10254,N_10255);
nor U10542 (N_10542,N_10337,N_10309);
or U10543 (N_10543,N_10385,N_10341);
xnor U10544 (N_10544,N_10220,N_10337);
or U10545 (N_10545,N_10289,N_10377);
nand U10546 (N_10546,N_10247,N_10237);
and U10547 (N_10547,N_10348,N_10211);
xor U10548 (N_10548,N_10295,N_10317);
xnor U10549 (N_10549,N_10274,N_10264);
xnor U10550 (N_10550,N_10369,N_10230);
nand U10551 (N_10551,N_10260,N_10209);
and U10552 (N_10552,N_10224,N_10217);
or U10553 (N_10553,N_10310,N_10290);
nor U10554 (N_10554,N_10326,N_10275);
nor U10555 (N_10555,N_10218,N_10263);
nand U10556 (N_10556,N_10300,N_10353);
or U10557 (N_10557,N_10248,N_10346);
nand U10558 (N_10558,N_10285,N_10326);
nand U10559 (N_10559,N_10265,N_10206);
xnor U10560 (N_10560,N_10226,N_10313);
or U10561 (N_10561,N_10326,N_10208);
or U10562 (N_10562,N_10391,N_10232);
or U10563 (N_10563,N_10385,N_10332);
or U10564 (N_10564,N_10202,N_10273);
nor U10565 (N_10565,N_10342,N_10270);
and U10566 (N_10566,N_10345,N_10347);
or U10567 (N_10567,N_10258,N_10319);
nor U10568 (N_10568,N_10375,N_10345);
nand U10569 (N_10569,N_10372,N_10275);
nand U10570 (N_10570,N_10255,N_10380);
xor U10571 (N_10571,N_10242,N_10390);
or U10572 (N_10572,N_10393,N_10317);
nand U10573 (N_10573,N_10323,N_10325);
xnor U10574 (N_10574,N_10385,N_10223);
nor U10575 (N_10575,N_10363,N_10341);
or U10576 (N_10576,N_10245,N_10337);
and U10577 (N_10577,N_10351,N_10330);
or U10578 (N_10578,N_10263,N_10319);
xor U10579 (N_10579,N_10275,N_10211);
and U10580 (N_10580,N_10285,N_10305);
or U10581 (N_10581,N_10339,N_10312);
nand U10582 (N_10582,N_10289,N_10221);
or U10583 (N_10583,N_10216,N_10271);
xnor U10584 (N_10584,N_10316,N_10201);
nand U10585 (N_10585,N_10294,N_10215);
nor U10586 (N_10586,N_10352,N_10247);
nor U10587 (N_10587,N_10232,N_10308);
nor U10588 (N_10588,N_10227,N_10216);
or U10589 (N_10589,N_10349,N_10311);
xor U10590 (N_10590,N_10371,N_10382);
nand U10591 (N_10591,N_10224,N_10259);
and U10592 (N_10592,N_10215,N_10289);
xor U10593 (N_10593,N_10350,N_10363);
nand U10594 (N_10594,N_10250,N_10338);
xnor U10595 (N_10595,N_10288,N_10243);
xor U10596 (N_10596,N_10228,N_10383);
xnor U10597 (N_10597,N_10345,N_10331);
or U10598 (N_10598,N_10273,N_10295);
nand U10599 (N_10599,N_10205,N_10392);
nand U10600 (N_10600,N_10510,N_10456);
nand U10601 (N_10601,N_10452,N_10583);
or U10602 (N_10602,N_10439,N_10445);
or U10603 (N_10603,N_10523,N_10418);
nor U10604 (N_10604,N_10547,N_10474);
or U10605 (N_10605,N_10580,N_10434);
nand U10606 (N_10606,N_10514,N_10435);
nand U10607 (N_10607,N_10486,N_10576);
xor U10608 (N_10608,N_10455,N_10424);
nor U10609 (N_10609,N_10417,N_10575);
and U10610 (N_10610,N_10561,N_10488);
and U10611 (N_10611,N_10470,N_10512);
and U10612 (N_10612,N_10536,N_10421);
or U10613 (N_10613,N_10517,N_10578);
or U10614 (N_10614,N_10433,N_10599);
or U10615 (N_10615,N_10581,N_10416);
nor U10616 (N_10616,N_10577,N_10403);
xnor U10617 (N_10617,N_10407,N_10477);
and U10618 (N_10618,N_10595,N_10543);
nor U10619 (N_10619,N_10442,N_10430);
or U10620 (N_10620,N_10461,N_10506);
xor U10621 (N_10621,N_10548,N_10405);
nand U10622 (N_10622,N_10437,N_10485);
xnor U10623 (N_10623,N_10431,N_10492);
nand U10624 (N_10624,N_10473,N_10457);
nand U10625 (N_10625,N_10411,N_10568);
and U10626 (N_10626,N_10436,N_10588);
and U10627 (N_10627,N_10546,N_10410);
xnor U10628 (N_10628,N_10464,N_10467);
and U10629 (N_10629,N_10597,N_10469);
xnor U10630 (N_10630,N_10545,N_10412);
nor U10631 (N_10631,N_10458,N_10446);
xor U10632 (N_10632,N_10402,N_10400);
or U10633 (N_10633,N_10482,N_10489);
and U10634 (N_10634,N_10560,N_10563);
or U10635 (N_10635,N_10462,N_10513);
or U10636 (N_10636,N_10590,N_10524);
and U10637 (N_10637,N_10479,N_10502);
or U10638 (N_10638,N_10549,N_10495);
or U10639 (N_10639,N_10528,N_10592);
nand U10640 (N_10640,N_10539,N_10498);
nand U10641 (N_10641,N_10526,N_10573);
and U10642 (N_10642,N_10422,N_10562);
nor U10643 (N_10643,N_10589,N_10552);
and U10644 (N_10644,N_10420,N_10428);
nand U10645 (N_10645,N_10567,N_10542);
or U10646 (N_10646,N_10448,N_10518);
or U10647 (N_10647,N_10409,N_10509);
nand U10648 (N_10648,N_10504,N_10566);
and U10649 (N_10649,N_10508,N_10465);
and U10650 (N_10650,N_10565,N_10438);
or U10651 (N_10651,N_10443,N_10534);
or U10652 (N_10652,N_10544,N_10564);
nor U10653 (N_10653,N_10587,N_10537);
and U10654 (N_10654,N_10427,N_10538);
nand U10655 (N_10655,N_10463,N_10572);
xor U10656 (N_10656,N_10440,N_10530);
and U10657 (N_10657,N_10529,N_10451);
and U10658 (N_10658,N_10559,N_10532);
or U10659 (N_10659,N_10503,N_10460);
or U10660 (N_10660,N_10419,N_10515);
and U10661 (N_10661,N_10550,N_10525);
xnor U10662 (N_10662,N_10408,N_10475);
or U10663 (N_10663,N_10404,N_10476);
and U10664 (N_10664,N_10401,N_10551);
nand U10665 (N_10665,N_10484,N_10423);
and U10666 (N_10666,N_10406,N_10493);
and U10667 (N_10667,N_10585,N_10535);
and U10668 (N_10668,N_10594,N_10429);
xnor U10669 (N_10669,N_10557,N_10540);
nor U10670 (N_10670,N_10449,N_10533);
nor U10671 (N_10671,N_10491,N_10413);
and U10672 (N_10672,N_10569,N_10432);
or U10673 (N_10673,N_10497,N_10415);
and U10674 (N_10674,N_10505,N_10447);
and U10675 (N_10675,N_10466,N_10553);
or U10676 (N_10676,N_10582,N_10558);
nand U10677 (N_10677,N_10450,N_10579);
xor U10678 (N_10678,N_10441,N_10527);
nand U10679 (N_10679,N_10499,N_10586);
xnor U10680 (N_10680,N_10481,N_10521);
nor U10681 (N_10681,N_10471,N_10500);
nor U10682 (N_10682,N_10472,N_10478);
and U10683 (N_10683,N_10511,N_10570);
or U10684 (N_10684,N_10496,N_10519);
xor U10685 (N_10685,N_10501,N_10531);
xnor U10686 (N_10686,N_10454,N_10494);
and U10687 (N_10687,N_10487,N_10584);
or U10688 (N_10688,N_10591,N_10426);
nor U10689 (N_10689,N_10571,N_10574);
xnor U10690 (N_10690,N_10490,N_10522);
nand U10691 (N_10691,N_10507,N_10596);
nor U10692 (N_10692,N_10459,N_10516);
nor U10693 (N_10693,N_10554,N_10414);
nor U10694 (N_10694,N_10468,N_10480);
nor U10695 (N_10695,N_10520,N_10555);
nand U10696 (N_10696,N_10556,N_10483);
and U10697 (N_10697,N_10593,N_10541);
and U10698 (N_10698,N_10425,N_10453);
or U10699 (N_10699,N_10444,N_10598);
nor U10700 (N_10700,N_10530,N_10453);
or U10701 (N_10701,N_10445,N_10473);
and U10702 (N_10702,N_10496,N_10550);
nand U10703 (N_10703,N_10411,N_10551);
nand U10704 (N_10704,N_10430,N_10492);
nor U10705 (N_10705,N_10537,N_10592);
or U10706 (N_10706,N_10415,N_10444);
xnor U10707 (N_10707,N_10498,N_10495);
nand U10708 (N_10708,N_10552,N_10509);
and U10709 (N_10709,N_10431,N_10521);
xnor U10710 (N_10710,N_10582,N_10432);
xor U10711 (N_10711,N_10407,N_10596);
nand U10712 (N_10712,N_10426,N_10594);
nor U10713 (N_10713,N_10439,N_10576);
xnor U10714 (N_10714,N_10567,N_10447);
or U10715 (N_10715,N_10510,N_10546);
and U10716 (N_10716,N_10554,N_10566);
nor U10717 (N_10717,N_10495,N_10514);
nor U10718 (N_10718,N_10455,N_10447);
nand U10719 (N_10719,N_10590,N_10536);
and U10720 (N_10720,N_10415,N_10572);
nor U10721 (N_10721,N_10551,N_10438);
nor U10722 (N_10722,N_10550,N_10498);
or U10723 (N_10723,N_10587,N_10578);
nor U10724 (N_10724,N_10443,N_10551);
nor U10725 (N_10725,N_10445,N_10475);
nor U10726 (N_10726,N_10418,N_10557);
and U10727 (N_10727,N_10412,N_10431);
xnor U10728 (N_10728,N_10407,N_10594);
nor U10729 (N_10729,N_10445,N_10560);
or U10730 (N_10730,N_10535,N_10566);
or U10731 (N_10731,N_10410,N_10511);
nand U10732 (N_10732,N_10411,N_10489);
and U10733 (N_10733,N_10598,N_10473);
or U10734 (N_10734,N_10529,N_10463);
nand U10735 (N_10735,N_10555,N_10494);
nor U10736 (N_10736,N_10503,N_10542);
nor U10737 (N_10737,N_10543,N_10420);
nor U10738 (N_10738,N_10551,N_10496);
nor U10739 (N_10739,N_10549,N_10472);
nor U10740 (N_10740,N_10438,N_10567);
nor U10741 (N_10741,N_10444,N_10547);
and U10742 (N_10742,N_10576,N_10485);
nor U10743 (N_10743,N_10577,N_10413);
and U10744 (N_10744,N_10509,N_10425);
nor U10745 (N_10745,N_10553,N_10435);
and U10746 (N_10746,N_10420,N_10482);
nand U10747 (N_10747,N_10557,N_10464);
or U10748 (N_10748,N_10571,N_10461);
nor U10749 (N_10749,N_10514,N_10461);
nand U10750 (N_10750,N_10424,N_10589);
xnor U10751 (N_10751,N_10587,N_10417);
nand U10752 (N_10752,N_10413,N_10499);
and U10753 (N_10753,N_10526,N_10578);
xor U10754 (N_10754,N_10505,N_10565);
xor U10755 (N_10755,N_10584,N_10415);
and U10756 (N_10756,N_10405,N_10425);
nand U10757 (N_10757,N_10411,N_10563);
and U10758 (N_10758,N_10418,N_10439);
nand U10759 (N_10759,N_10526,N_10421);
or U10760 (N_10760,N_10545,N_10468);
nor U10761 (N_10761,N_10466,N_10505);
or U10762 (N_10762,N_10455,N_10545);
or U10763 (N_10763,N_10403,N_10484);
or U10764 (N_10764,N_10440,N_10586);
xor U10765 (N_10765,N_10471,N_10416);
xor U10766 (N_10766,N_10555,N_10421);
nor U10767 (N_10767,N_10540,N_10550);
or U10768 (N_10768,N_10427,N_10468);
and U10769 (N_10769,N_10465,N_10422);
or U10770 (N_10770,N_10410,N_10465);
nor U10771 (N_10771,N_10595,N_10575);
nor U10772 (N_10772,N_10430,N_10536);
and U10773 (N_10773,N_10467,N_10413);
nand U10774 (N_10774,N_10418,N_10441);
or U10775 (N_10775,N_10459,N_10541);
nand U10776 (N_10776,N_10533,N_10511);
or U10777 (N_10777,N_10503,N_10525);
nand U10778 (N_10778,N_10531,N_10470);
nor U10779 (N_10779,N_10493,N_10457);
nand U10780 (N_10780,N_10532,N_10502);
xor U10781 (N_10781,N_10542,N_10498);
or U10782 (N_10782,N_10402,N_10442);
nand U10783 (N_10783,N_10543,N_10592);
and U10784 (N_10784,N_10598,N_10405);
nand U10785 (N_10785,N_10412,N_10459);
and U10786 (N_10786,N_10579,N_10484);
or U10787 (N_10787,N_10533,N_10446);
nor U10788 (N_10788,N_10500,N_10451);
nor U10789 (N_10789,N_10481,N_10402);
or U10790 (N_10790,N_10480,N_10599);
nor U10791 (N_10791,N_10467,N_10510);
or U10792 (N_10792,N_10422,N_10489);
nand U10793 (N_10793,N_10440,N_10542);
or U10794 (N_10794,N_10505,N_10542);
nor U10795 (N_10795,N_10541,N_10528);
nor U10796 (N_10796,N_10599,N_10593);
nand U10797 (N_10797,N_10517,N_10428);
nor U10798 (N_10798,N_10428,N_10411);
xor U10799 (N_10799,N_10494,N_10456);
or U10800 (N_10800,N_10704,N_10786);
xor U10801 (N_10801,N_10740,N_10686);
and U10802 (N_10802,N_10620,N_10745);
nor U10803 (N_10803,N_10748,N_10697);
or U10804 (N_10804,N_10691,N_10793);
and U10805 (N_10805,N_10654,N_10653);
xnor U10806 (N_10806,N_10613,N_10669);
xnor U10807 (N_10807,N_10731,N_10795);
and U10808 (N_10808,N_10660,N_10672);
nor U10809 (N_10809,N_10711,N_10758);
or U10810 (N_10810,N_10646,N_10602);
nor U10811 (N_10811,N_10617,N_10724);
xnor U10812 (N_10812,N_10670,N_10750);
and U10813 (N_10813,N_10766,N_10722);
xor U10814 (N_10814,N_10650,N_10744);
nor U10815 (N_10815,N_10727,N_10717);
xnor U10816 (N_10816,N_10623,N_10682);
or U10817 (N_10817,N_10754,N_10796);
and U10818 (N_10818,N_10762,N_10607);
nor U10819 (N_10819,N_10600,N_10657);
or U10820 (N_10820,N_10627,N_10773);
nand U10821 (N_10821,N_10714,N_10785);
nand U10822 (N_10822,N_10619,N_10703);
or U10823 (N_10823,N_10792,N_10688);
nor U10824 (N_10824,N_10708,N_10692);
xor U10825 (N_10825,N_10683,N_10763);
nand U10826 (N_10826,N_10666,N_10713);
and U10827 (N_10827,N_10676,N_10732);
and U10828 (N_10828,N_10733,N_10625);
or U10829 (N_10829,N_10655,N_10614);
nand U10830 (N_10830,N_10626,N_10765);
and U10831 (N_10831,N_10606,N_10684);
or U10832 (N_10832,N_10642,N_10737);
and U10833 (N_10833,N_10680,N_10638);
nand U10834 (N_10834,N_10712,N_10618);
xnor U10835 (N_10835,N_10734,N_10649);
xnor U10836 (N_10836,N_10735,N_10611);
or U10837 (N_10837,N_10757,N_10752);
and U10838 (N_10838,N_10647,N_10636);
xnor U10839 (N_10839,N_10610,N_10756);
nand U10840 (N_10840,N_10782,N_10780);
or U10841 (N_10841,N_10690,N_10742);
nor U10842 (N_10842,N_10759,N_10746);
xor U10843 (N_10843,N_10720,N_10641);
nand U10844 (N_10844,N_10738,N_10685);
xor U10845 (N_10845,N_10687,N_10630);
xnor U10846 (N_10846,N_10609,N_10749);
nor U10847 (N_10847,N_10662,N_10698);
xnor U10848 (N_10848,N_10751,N_10665);
nor U10849 (N_10849,N_10633,N_10729);
and U10850 (N_10850,N_10718,N_10770);
or U10851 (N_10851,N_10689,N_10632);
xor U10852 (N_10852,N_10677,N_10652);
xor U10853 (N_10853,N_10710,N_10634);
or U10854 (N_10854,N_10648,N_10621);
or U10855 (N_10855,N_10747,N_10776);
nand U10856 (N_10856,N_10739,N_10694);
nor U10857 (N_10857,N_10730,N_10679);
and U10858 (N_10858,N_10787,N_10781);
nor U10859 (N_10859,N_10667,N_10701);
and U10860 (N_10860,N_10678,N_10784);
nor U10861 (N_10861,N_10673,N_10719);
and U10862 (N_10862,N_10658,N_10755);
and U10863 (N_10863,N_10772,N_10693);
or U10864 (N_10864,N_10775,N_10774);
or U10865 (N_10865,N_10702,N_10663);
xor U10866 (N_10866,N_10706,N_10699);
nor U10867 (N_10867,N_10664,N_10791);
and U10868 (N_10868,N_10767,N_10707);
and U10869 (N_10869,N_10779,N_10656);
and U10870 (N_10870,N_10651,N_10631);
and U10871 (N_10871,N_10705,N_10790);
or U10872 (N_10872,N_10622,N_10721);
nand U10873 (N_10873,N_10681,N_10696);
or U10874 (N_10874,N_10778,N_10624);
and U10875 (N_10875,N_10764,N_10675);
and U10876 (N_10876,N_10777,N_10797);
or U10877 (N_10877,N_10608,N_10736);
nor U10878 (N_10878,N_10760,N_10643);
xnor U10879 (N_10879,N_10616,N_10640);
and U10880 (N_10880,N_10771,N_10728);
nor U10881 (N_10881,N_10628,N_10798);
xor U10882 (N_10882,N_10661,N_10715);
xor U10883 (N_10883,N_10743,N_10761);
nor U10884 (N_10884,N_10615,N_10635);
nand U10885 (N_10885,N_10799,N_10709);
xor U10886 (N_10886,N_10726,N_10695);
xor U10887 (N_10887,N_10671,N_10629);
and U10888 (N_10888,N_10645,N_10644);
xor U10889 (N_10889,N_10605,N_10604);
and U10890 (N_10890,N_10769,N_10768);
nor U10891 (N_10891,N_10639,N_10637);
nor U10892 (N_10892,N_10783,N_10725);
and U10893 (N_10893,N_10601,N_10723);
and U10894 (N_10894,N_10753,N_10668);
nand U10895 (N_10895,N_10741,N_10788);
nand U10896 (N_10896,N_10700,N_10794);
or U10897 (N_10897,N_10659,N_10789);
xnor U10898 (N_10898,N_10716,N_10674);
nor U10899 (N_10899,N_10603,N_10612);
and U10900 (N_10900,N_10623,N_10768);
and U10901 (N_10901,N_10607,N_10763);
nand U10902 (N_10902,N_10673,N_10605);
nor U10903 (N_10903,N_10723,N_10793);
nand U10904 (N_10904,N_10629,N_10658);
nand U10905 (N_10905,N_10729,N_10769);
or U10906 (N_10906,N_10631,N_10645);
nand U10907 (N_10907,N_10671,N_10638);
nor U10908 (N_10908,N_10701,N_10739);
xor U10909 (N_10909,N_10634,N_10646);
nand U10910 (N_10910,N_10725,N_10784);
or U10911 (N_10911,N_10619,N_10633);
xor U10912 (N_10912,N_10788,N_10697);
xnor U10913 (N_10913,N_10736,N_10777);
and U10914 (N_10914,N_10724,N_10770);
or U10915 (N_10915,N_10785,N_10632);
or U10916 (N_10916,N_10785,N_10742);
xor U10917 (N_10917,N_10654,N_10610);
nor U10918 (N_10918,N_10750,N_10740);
and U10919 (N_10919,N_10707,N_10756);
nand U10920 (N_10920,N_10619,N_10730);
nor U10921 (N_10921,N_10741,N_10770);
or U10922 (N_10922,N_10628,N_10766);
nand U10923 (N_10923,N_10730,N_10759);
xor U10924 (N_10924,N_10760,N_10743);
or U10925 (N_10925,N_10770,N_10799);
and U10926 (N_10926,N_10737,N_10679);
nand U10927 (N_10927,N_10611,N_10682);
nor U10928 (N_10928,N_10736,N_10646);
or U10929 (N_10929,N_10705,N_10627);
nor U10930 (N_10930,N_10652,N_10660);
and U10931 (N_10931,N_10772,N_10609);
nand U10932 (N_10932,N_10679,N_10669);
and U10933 (N_10933,N_10740,N_10769);
nand U10934 (N_10934,N_10724,N_10780);
and U10935 (N_10935,N_10622,N_10785);
nor U10936 (N_10936,N_10617,N_10644);
and U10937 (N_10937,N_10681,N_10607);
nand U10938 (N_10938,N_10696,N_10791);
nor U10939 (N_10939,N_10713,N_10746);
nor U10940 (N_10940,N_10786,N_10797);
or U10941 (N_10941,N_10753,N_10737);
or U10942 (N_10942,N_10757,N_10662);
nand U10943 (N_10943,N_10648,N_10706);
and U10944 (N_10944,N_10673,N_10749);
nor U10945 (N_10945,N_10784,N_10648);
and U10946 (N_10946,N_10793,N_10661);
nor U10947 (N_10947,N_10620,N_10720);
or U10948 (N_10948,N_10674,N_10698);
xnor U10949 (N_10949,N_10664,N_10712);
nand U10950 (N_10950,N_10782,N_10606);
and U10951 (N_10951,N_10733,N_10607);
nand U10952 (N_10952,N_10610,N_10613);
or U10953 (N_10953,N_10726,N_10793);
or U10954 (N_10954,N_10722,N_10645);
and U10955 (N_10955,N_10636,N_10667);
xor U10956 (N_10956,N_10690,N_10696);
nand U10957 (N_10957,N_10719,N_10650);
and U10958 (N_10958,N_10674,N_10682);
or U10959 (N_10959,N_10673,N_10663);
xor U10960 (N_10960,N_10678,N_10751);
and U10961 (N_10961,N_10634,N_10792);
xnor U10962 (N_10962,N_10666,N_10639);
or U10963 (N_10963,N_10690,N_10727);
or U10964 (N_10964,N_10763,N_10773);
nor U10965 (N_10965,N_10714,N_10727);
xnor U10966 (N_10966,N_10668,N_10692);
nor U10967 (N_10967,N_10626,N_10625);
nor U10968 (N_10968,N_10627,N_10728);
or U10969 (N_10969,N_10631,N_10663);
xor U10970 (N_10970,N_10642,N_10739);
and U10971 (N_10971,N_10728,N_10743);
nand U10972 (N_10972,N_10718,N_10603);
nor U10973 (N_10973,N_10646,N_10761);
xor U10974 (N_10974,N_10674,N_10717);
or U10975 (N_10975,N_10675,N_10740);
nor U10976 (N_10976,N_10757,N_10704);
or U10977 (N_10977,N_10654,N_10649);
or U10978 (N_10978,N_10699,N_10778);
nand U10979 (N_10979,N_10683,N_10751);
or U10980 (N_10980,N_10648,N_10679);
xnor U10981 (N_10981,N_10715,N_10683);
xnor U10982 (N_10982,N_10602,N_10783);
nor U10983 (N_10983,N_10603,N_10698);
and U10984 (N_10984,N_10607,N_10672);
nand U10985 (N_10985,N_10761,N_10615);
and U10986 (N_10986,N_10687,N_10747);
or U10987 (N_10987,N_10758,N_10623);
nand U10988 (N_10988,N_10764,N_10752);
nor U10989 (N_10989,N_10701,N_10742);
nor U10990 (N_10990,N_10695,N_10638);
xnor U10991 (N_10991,N_10727,N_10778);
or U10992 (N_10992,N_10712,N_10621);
xor U10993 (N_10993,N_10664,N_10735);
xnor U10994 (N_10994,N_10786,N_10709);
and U10995 (N_10995,N_10657,N_10782);
nor U10996 (N_10996,N_10788,N_10792);
nand U10997 (N_10997,N_10721,N_10753);
nor U10998 (N_10998,N_10748,N_10794);
or U10999 (N_10999,N_10754,N_10688);
or U11000 (N_11000,N_10889,N_10807);
nor U11001 (N_11001,N_10882,N_10865);
or U11002 (N_11002,N_10925,N_10842);
or U11003 (N_11003,N_10816,N_10870);
xor U11004 (N_11004,N_10952,N_10953);
xnor U11005 (N_11005,N_10904,N_10970);
nand U11006 (N_11006,N_10985,N_10828);
or U11007 (N_11007,N_10948,N_10845);
nor U11008 (N_11008,N_10944,N_10976);
nand U11009 (N_11009,N_10871,N_10831);
nor U11010 (N_11010,N_10818,N_10800);
and U11011 (N_11011,N_10884,N_10808);
nand U11012 (N_11012,N_10931,N_10932);
or U11013 (N_11013,N_10911,N_10829);
nand U11014 (N_11014,N_10851,N_10955);
nand U11015 (N_11015,N_10862,N_10959);
or U11016 (N_11016,N_10835,N_10858);
xnor U11017 (N_11017,N_10958,N_10830);
nand U11018 (N_11018,N_10805,N_10941);
or U11019 (N_11019,N_10850,N_10993);
nand U11020 (N_11020,N_10811,N_10900);
nand U11021 (N_11021,N_10975,N_10906);
and U11022 (N_11022,N_10979,N_10936);
and U11023 (N_11023,N_10832,N_10934);
nand U11024 (N_11024,N_10998,N_10815);
nand U11025 (N_11025,N_10864,N_10867);
xor U11026 (N_11026,N_10841,N_10988);
nor U11027 (N_11027,N_10886,N_10892);
nand U11028 (N_11028,N_10847,N_10986);
nor U11029 (N_11029,N_10877,N_10946);
and U11030 (N_11030,N_10846,N_10875);
and U11031 (N_11031,N_10919,N_10987);
or U11032 (N_11032,N_10924,N_10956);
and U11033 (N_11033,N_10945,N_10869);
xor U11034 (N_11034,N_10814,N_10967);
or U11035 (N_11035,N_10881,N_10933);
or U11036 (N_11036,N_10999,N_10969);
and U11037 (N_11037,N_10821,N_10995);
xor U11038 (N_11038,N_10834,N_10839);
xor U11039 (N_11039,N_10950,N_10801);
xor U11040 (N_11040,N_10806,N_10916);
xnor U11041 (N_11041,N_10844,N_10923);
or U11042 (N_11042,N_10960,N_10902);
and U11043 (N_11043,N_10938,N_10973);
or U11044 (N_11044,N_10843,N_10891);
nand U11045 (N_11045,N_10833,N_10957);
nor U11046 (N_11046,N_10826,N_10861);
and U11047 (N_11047,N_10894,N_10927);
xor U11048 (N_11048,N_10812,N_10878);
and U11049 (N_11049,N_10918,N_10823);
nand U11050 (N_11050,N_10863,N_10940);
xor U11051 (N_11051,N_10874,N_10962);
nand U11052 (N_11052,N_10853,N_10819);
nand U11053 (N_11053,N_10939,N_10890);
or U11054 (N_11054,N_10897,N_10898);
and U11055 (N_11055,N_10803,N_10942);
xor U11056 (N_11056,N_10978,N_10926);
nand U11057 (N_11057,N_10947,N_10840);
and U11058 (N_11058,N_10961,N_10930);
or U11059 (N_11059,N_10971,N_10912);
xor U11060 (N_11060,N_10849,N_10943);
nand U11061 (N_11061,N_10836,N_10968);
nor U11062 (N_11062,N_10876,N_10885);
xnor U11063 (N_11063,N_10903,N_10997);
nor U11064 (N_11064,N_10951,N_10905);
nand U11065 (N_11065,N_10852,N_10972);
nand U11066 (N_11066,N_10813,N_10817);
nor U11067 (N_11067,N_10825,N_10901);
and U11068 (N_11068,N_10802,N_10888);
or U11069 (N_11069,N_10983,N_10883);
nor U11070 (N_11070,N_10866,N_10982);
nand U11071 (N_11071,N_10827,N_10954);
and U11072 (N_11072,N_10928,N_10879);
or U11073 (N_11073,N_10915,N_10873);
and U11074 (N_11074,N_10822,N_10872);
nand U11075 (N_11075,N_10963,N_10990);
and U11076 (N_11076,N_10887,N_10989);
xnor U11077 (N_11077,N_10880,N_10856);
nor U11078 (N_11078,N_10820,N_10994);
and U11079 (N_11079,N_10838,N_10977);
nor U11080 (N_11080,N_10935,N_10907);
nor U11081 (N_11081,N_10980,N_10859);
xnor U11082 (N_11082,N_10824,N_10914);
xnor U11083 (N_11083,N_10991,N_10896);
and U11084 (N_11084,N_10984,N_10804);
nor U11085 (N_11085,N_10895,N_10899);
nand U11086 (N_11086,N_10974,N_10855);
nor U11087 (N_11087,N_10893,N_10996);
nor U11088 (N_11088,N_10937,N_10854);
nor U11089 (N_11089,N_10809,N_10992);
xor U11090 (N_11090,N_10913,N_10837);
nor U11091 (N_11091,N_10910,N_10965);
xnor U11092 (N_11092,N_10917,N_10921);
and U11093 (N_11093,N_10868,N_10929);
nor U11094 (N_11094,N_10860,N_10810);
xor U11095 (N_11095,N_10857,N_10922);
nand U11096 (N_11096,N_10920,N_10949);
nor U11097 (N_11097,N_10964,N_10966);
or U11098 (N_11098,N_10909,N_10908);
or U11099 (N_11099,N_10848,N_10981);
nor U11100 (N_11100,N_10860,N_10901);
nor U11101 (N_11101,N_10942,N_10982);
xnor U11102 (N_11102,N_10836,N_10936);
or U11103 (N_11103,N_10848,N_10935);
and U11104 (N_11104,N_10849,N_10999);
nor U11105 (N_11105,N_10986,N_10948);
xnor U11106 (N_11106,N_10984,N_10805);
or U11107 (N_11107,N_10963,N_10848);
and U11108 (N_11108,N_10845,N_10925);
nor U11109 (N_11109,N_10830,N_10810);
xor U11110 (N_11110,N_10962,N_10841);
and U11111 (N_11111,N_10893,N_10990);
nor U11112 (N_11112,N_10931,N_10991);
or U11113 (N_11113,N_10862,N_10883);
nand U11114 (N_11114,N_10936,N_10867);
nor U11115 (N_11115,N_10912,N_10963);
or U11116 (N_11116,N_10834,N_10846);
xor U11117 (N_11117,N_10905,N_10958);
nor U11118 (N_11118,N_10859,N_10981);
nor U11119 (N_11119,N_10942,N_10828);
nand U11120 (N_11120,N_10819,N_10846);
nor U11121 (N_11121,N_10836,N_10882);
xnor U11122 (N_11122,N_10805,N_10886);
or U11123 (N_11123,N_10939,N_10941);
xor U11124 (N_11124,N_10826,N_10966);
or U11125 (N_11125,N_10805,N_10875);
nor U11126 (N_11126,N_10984,N_10976);
nand U11127 (N_11127,N_10828,N_10802);
and U11128 (N_11128,N_10999,N_10841);
and U11129 (N_11129,N_10830,N_10856);
and U11130 (N_11130,N_10823,N_10950);
xor U11131 (N_11131,N_10852,N_10810);
nor U11132 (N_11132,N_10966,N_10840);
nor U11133 (N_11133,N_10836,N_10867);
and U11134 (N_11134,N_10956,N_10821);
or U11135 (N_11135,N_10974,N_10941);
and U11136 (N_11136,N_10852,N_10861);
nand U11137 (N_11137,N_10859,N_10999);
nor U11138 (N_11138,N_10816,N_10980);
nand U11139 (N_11139,N_10961,N_10822);
nand U11140 (N_11140,N_10863,N_10816);
or U11141 (N_11141,N_10949,N_10854);
or U11142 (N_11142,N_10819,N_10925);
nand U11143 (N_11143,N_10819,N_10802);
or U11144 (N_11144,N_10965,N_10914);
nand U11145 (N_11145,N_10907,N_10887);
nand U11146 (N_11146,N_10827,N_10819);
xor U11147 (N_11147,N_10947,N_10849);
and U11148 (N_11148,N_10862,N_10817);
and U11149 (N_11149,N_10907,N_10809);
nor U11150 (N_11150,N_10931,N_10974);
or U11151 (N_11151,N_10806,N_10955);
nor U11152 (N_11152,N_10886,N_10833);
or U11153 (N_11153,N_10852,N_10830);
xnor U11154 (N_11154,N_10964,N_10818);
or U11155 (N_11155,N_10908,N_10914);
xor U11156 (N_11156,N_10979,N_10885);
and U11157 (N_11157,N_10991,N_10933);
or U11158 (N_11158,N_10907,N_10922);
or U11159 (N_11159,N_10870,N_10956);
and U11160 (N_11160,N_10971,N_10853);
or U11161 (N_11161,N_10810,N_10919);
or U11162 (N_11162,N_10885,N_10815);
xnor U11163 (N_11163,N_10927,N_10862);
nor U11164 (N_11164,N_10836,N_10919);
nand U11165 (N_11165,N_10931,N_10838);
or U11166 (N_11166,N_10827,N_10910);
and U11167 (N_11167,N_10895,N_10912);
or U11168 (N_11168,N_10804,N_10899);
nand U11169 (N_11169,N_10824,N_10967);
xor U11170 (N_11170,N_10818,N_10880);
nand U11171 (N_11171,N_10879,N_10826);
and U11172 (N_11172,N_10856,N_10824);
and U11173 (N_11173,N_10961,N_10808);
nor U11174 (N_11174,N_10834,N_10979);
nand U11175 (N_11175,N_10855,N_10927);
nand U11176 (N_11176,N_10904,N_10905);
nand U11177 (N_11177,N_10946,N_10838);
nand U11178 (N_11178,N_10907,N_10855);
and U11179 (N_11179,N_10814,N_10942);
and U11180 (N_11180,N_10889,N_10849);
nand U11181 (N_11181,N_10909,N_10869);
and U11182 (N_11182,N_10869,N_10874);
and U11183 (N_11183,N_10841,N_10860);
nor U11184 (N_11184,N_10881,N_10895);
nor U11185 (N_11185,N_10998,N_10803);
and U11186 (N_11186,N_10888,N_10813);
nand U11187 (N_11187,N_10870,N_10909);
nor U11188 (N_11188,N_10931,N_10826);
nand U11189 (N_11189,N_10903,N_10816);
xnor U11190 (N_11190,N_10983,N_10819);
or U11191 (N_11191,N_10911,N_10809);
nand U11192 (N_11192,N_10903,N_10840);
xor U11193 (N_11193,N_10942,N_10958);
or U11194 (N_11194,N_10892,N_10827);
nor U11195 (N_11195,N_10804,N_10854);
nor U11196 (N_11196,N_10985,N_10906);
or U11197 (N_11197,N_10952,N_10921);
or U11198 (N_11198,N_10982,N_10826);
nor U11199 (N_11199,N_10904,N_10961);
or U11200 (N_11200,N_11129,N_11138);
and U11201 (N_11201,N_11013,N_11080);
nor U11202 (N_11202,N_11065,N_11122);
or U11203 (N_11203,N_11068,N_11160);
nor U11204 (N_11204,N_11182,N_11052);
xnor U11205 (N_11205,N_11055,N_11166);
or U11206 (N_11206,N_11192,N_11021);
or U11207 (N_11207,N_11035,N_11041);
nor U11208 (N_11208,N_11137,N_11007);
nand U11209 (N_11209,N_11092,N_11156);
or U11210 (N_11210,N_11186,N_11164);
and U11211 (N_11211,N_11043,N_11142);
xnor U11212 (N_11212,N_11171,N_11153);
nor U11213 (N_11213,N_11066,N_11109);
nor U11214 (N_11214,N_11016,N_11032);
and U11215 (N_11215,N_11075,N_11012);
nand U11216 (N_11216,N_11159,N_11094);
nor U11217 (N_11217,N_11106,N_11028);
and U11218 (N_11218,N_11090,N_11074);
and U11219 (N_11219,N_11127,N_11133);
xor U11220 (N_11220,N_11185,N_11022);
nand U11221 (N_11221,N_11034,N_11067);
and U11222 (N_11222,N_11108,N_11100);
nor U11223 (N_11223,N_11161,N_11199);
or U11224 (N_11224,N_11151,N_11157);
nor U11225 (N_11225,N_11070,N_11045);
or U11226 (N_11226,N_11145,N_11173);
nand U11227 (N_11227,N_11096,N_11040);
or U11228 (N_11228,N_11063,N_11003);
nor U11229 (N_11229,N_11027,N_11103);
xnor U11230 (N_11230,N_11167,N_11168);
nor U11231 (N_11231,N_11006,N_11169);
nand U11232 (N_11232,N_11078,N_11004);
xnor U11233 (N_11233,N_11158,N_11180);
and U11234 (N_11234,N_11010,N_11190);
and U11235 (N_11235,N_11146,N_11044);
nand U11236 (N_11236,N_11011,N_11001);
nand U11237 (N_11237,N_11076,N_11197);
nand U11238 (N_11238,N_11087,N_11111);
nor U11239 (N_11239,N_11117,N_11069);
and U11240 (N_11240,N_11147,N_11119);
and U11241 (N_11241,N_11097,N_11088);
nand U11242 (N_11242,N_11019,N_11175);
nor U11243 (N_11243,N_11072,N_11120);
and U11244 (N_11244,N_11048,N_11053);
or U11245 (N_11245,N_11023,N_11132);
and U11246 (N_11246,N_11193,N_11149);
nand U11247 (N_11247,N_11046,N_11163);
xnor U11248 (N_11248,N_11126,N_11136);
or U11249 (N_11249,N_11135,N_11150);
or U11250 (N_11250,N_11091,N_11005);
and U11251 (N_11251,N_11110,N_11026);
xor U11252 (N_11252,N_11061,N_11015);
and U11253 (N_11253,N_11077,N_11059);
and U11254 (N_11254,N_11073,N_11071);
xor U11255 (N_11255,N_11189,N_11084);
and U11256 (N_11256,N_11131,N_11064);
and U11257 (N_11257,N_11102,N_11143);
xnor U11258 (N_11258,N_11139,N_11025);
or U11259 (N_11259,N_11017,N_11191);
and U11260 (N_11260,N_11037,N_11085);
or U11261 (N_11261,N_11141,N_11172);
xnor U11262 (N_11262,N_11128,N_11047);
or U11263 (N_11263,N_11009,N_11113);
and U11264 (N_11264,N_11062,N_11123);
nor U11265 (N_11265,N_11174,N_11130);
or U11266 (N_11266,N_11116,N_11148);
nand U11267 (N_11267,N_11039,N_11056);
nand U11268 (N_11268,N_11134,N_11060);
or U11269 (N_11269,N_11124,N_11183);
nand U11270 (N_11270,N_11114,N_11118);
nor U11271 (N_11271,N_11162,N_11042);
nand U11272 (N_11272,N_11029,N_11195);
and U11273 (N_11273,N_11104,N_11030);
or U11274 (N_11274,N_11154,N_11144);
and U11275 (N_11275,N_11165,N_11086);
or U11276 (N_11276,N_11082,N_11051);
and U11277 (N_11277,N_11033,N_11170);
and U11278 (N_11278,N_11036,N_11196);
or U11279 (N_11279,N_11140,N_11014);
and U11280 (N_11280,N_11083,N_11089);
nor U11281 (N_11281,N_11002,N_11152);
or U11282 (N_11282,N_11187,N_11176);
nor U11283 (N_11283,N_11024,N_11018);
or U11284 (N_11284,N_11095,N_11107);
nand U11285 (N_11285,N_11057,N_11038);
and U11286 (N_11286,N_11125,N_11054);
and U11287 (N_11287,N_11079,N_11198);
nand U11288 (N_11288,N_11081,N_11000);
or U11289 (N_11289,N_11008,N_11194);
nand U11290 (N_11290,N_11031,N_11121);
and U11291 (N_11291,N_11101,N_11178);
and U11292 (N_11292,N_11184,N_11058);
nor U11293 (N_11293,N_11098,N_11099);
nand U11294 (N_11294,N_11188,N_11115);
or U11295 (N_11295,N_11112,N_11049);
or U11296 (N_11296,N_11093,N_11181);
and U11297 (N_11297,N_11105,N_11020);
nor U11298 (N_11298,N_11050,N_11177);
nand U11299 (N_11299,N_11179,N_11155);
xnor U11300 (N_11300,N_11052,N_11042);
or U11301 (N_11301,N_11030,N_11130);
nor U11302 (N_11302,N_11160,N_11187);
nand U11303 (N_11303,N_11188,N_11066);
nand U11304 (N_11304,N_11051,N_11004);
nand U11305 (N_11305,N_11060,N_11018);
or U11306 (N_11306,N_11070,N_11091);
or U11307 (N_11307,N_11080,N_11006);
nor U11308 (N_11308,N_11075,N_11097);
xnor U11309 (N_11309,N_11006,N_11017);
or U11310 (N_11310,N_11017,N_11104);
or U11311 (N_11311,N_11096,N_11100);
nor U11312 (N_11312,N_11181,N_11175);
and U11313 (N_11313,N_11199,N_11189);
and U11314 (N_11314,N_11122,N_11088);
nor U11315 (N_11315,N_11050,N_11108);
xnor U11316 (N_11316,N_11143,N_11127);
nand U11317 (N_11317,N_11180,N_11045);
or U11318 (N_11318,N_11169,N_11108);
nand U11319 (N_11319,N_11054,N_11010);
nor U11320 (N_11320,N_11174,N_11032);
xor U11321 (N_11321,N_11083,N_11118);
or U11322 (N_11322,N_11085,N_11067);
and U11323 (N_11323,N_11098,N_11180);
nand U11324 (N_11324,N_11049,N_11069);
and U11325 (N_11325,N_11061,N_11196);
nand U11326 (N_11326,N_11177,N_11151);
or U11327 (N_11327,N_11147,N_11092);
nor U11328 (N_11328,N_11139,N_11056);
or U11329 (N_11329,N_11142,N_11132);
and U11330 (N_11330,N_11127,N_11129);
nand U11331 (N_11331,N_11130,N_11029);
and U11332 (N_11332,N_11015,N_11169);
or U11333 (N_11333,N_11076,N_11018);
xnor U11334 (N_11334,N_11080,N_11180);
xor U11335 (N_11335,N_11004,N_11127);
nand U11336 (N_11336,N_11110,N_11161);
nor U11337 (N_11337,N_11130,N_11028);
nor U11338 (N_11338,N_11003,N_11007);
nor U11339 (N_11339,N_11031,N_11006);
xnor U11340 (N_11340,N_11169,N_11003);
xnor U11341 (N_11341,N_11184,N_11027);
and U11342 (N_11342,N_11066,N_11150);
nand U11343 (N_11343,N_11194,N_11033);
xor U11344 (N_11344,N_11164,N_11182);
nor U11345 (N_11345,N_11095,N_11017);
xnor U11346 (N_11346,N_11191,N_11161);
and U11347 (N_11347,N_11068,N_11126);
nand U11348 (N_11348,N_11089,N_11102);
nand U11349 (N_11349,N_11142,N_11079);
nand U11350 (N_11350,N_11160,N_11171);
nand U11351 (N_11351,N_11058,N_11132);
nor U11352 (N_11352,N_11121,N_11099);
nand U11353 (N_11353,N_11163,N_11189);
nand U11354 (N_11354,N_11119,N_11060);
and U11355 (N_11355,N_11025,N_11076);
or U11356 (N_11356,N_11080,N_11194);
xnor U11357 (N_11357,N_11191,N_11099);
and U11358 (N_11358,N_11113,N_11075);
xor U11359 (N_11359,N_11129,N_11156);
nand U11360 (N_11360,N_11017,N_11183);
nand U11361 (N_11361,N_11137,N_11030);
or U11362 (N_11362,N_11154,N_11132);
nand U11363 (N_11363,N_11108,N_11188);
and U11364 (N_11364,N_11132,N_11060);
nor U11365 (N_11365,N_11191,N_11173);
nand U11366 (N_11366,N_11181,N_11010);
nand U11367 (N_11367,N_11186,N_11080);
nand U11368 (N_11368,N_11054,N_11176);
nor U11369 (N_11369,N_11154,N_11151);
and U11370 (N_11370,N_11003,N_11021);
nand U11371 (N_11371,N_11139,N_11047);
nor U11372 (N_11372,N_11109,N_11019);
nor U11373 (N_11373,N_11002,N_11056);
xor U11374 (N_11374,N_11093,N_11042);
or U11375 (N_11375,N_11194,N_11170);
xor U11376 (N_11376,N_11087,N_11133);
nand U11377 (N_11377,N_11017,N_11175);
or U11378 (N_11378,N_11053,N_11188);
or U11379 (N_11379,N_11170,N_11196);
nor U11380 (N_11380,N_11024,N_11182);
and U11381 (N_11381,N_11055,N_11019);
xnor U11382 (N_11382,N_11018,N_11059);
nand U11383 (N_11383,N_11039,N_11129);
or U11384 (N_11384,N_11074,N_11000);
xor U11385 (N_11385,N_11042,N_11089);
nand U11386 (N_11386,N_11172,N_11136);
nand U11387 (N_11387,N_11087,N_11163);
nor U11388 (N_11388,N_11091,N_11060);
and U11389 (N_11389,N_11089,N_11113);
xnor U11390 (N_11390,N_11155,N_11054);
and U11391 (N_11391,N_11124,N_11144);
nand U11392 (N_11392,N_11038,N_11107);
or U11393 (N_11393,N_11022,N_11042);
or U11394 (N_11394,N_11021,N_11041);
or U11395 (N_11395,N_11070,N_11124);
and U11396 (N_11396,N_11085,N_11191);
and U11397 (N_11397,N_11166,N_11197);
nor U11398 (N_11398,N_11093,N_11163);
nand U11399 (N_11399,N_11129,N_11104);
and U11400 (N_11400,N_11388,N_11340);
xor U11401 (N_11401,N_11364,N_11330);
or U11402 (N_11402,N_11301,N_11251);
or U11403 (N_11403,N_11265,N_11317);
nand U11404 (N_11404,N_11336,N_11331);
nand U11405 (N_11405,N_11332,N_11391);
or U11406 (N_11406,N_11291,N_11360);
nand U11407 (N_11407,N_11215,N_11309);
nand U11408 (N_11408,N_11363,N_11202);
xor U11409 (N_11409,N_11290,N_11289);
and U11410 (N_11410,N_11344,N_11233);
xnor U11411 (N_11411,N_11281,N_11243);
xnor U11412 (N_11412,N_11351,N_11260);
nand U11413 (N_11413,N_11385,N_11314);
or U11414 (N_11414,N_11345,N_11339);
and U11415 (N_11415,N_11218,N_11298);
nand U11416 (N_11416,N_11378,N_11288);
and U11417 (N_11417,N_11230,N_11384);
xnor U11418 (N_11418,N_11312,N_11269);
xnor U11419 (N_11419,N_11252,N_11350);
nor U11420 (N_11420,N_11286,N_11263);
nand U11421 (N_11421,N_11329,N_11337);
or U11422 (N_11422,N_11241,N_11226);
nand U11423 (N_11423,N_11205,N_11315);
xnor U11424 (N_11424,N_11273,N_11280);
nor U11425 (N_11425,N_11200,N_11313);
and U11426 (N_11426,N_11308,N_11392);
nor U11427 (N_11427,N_11250,N_11367);
and U11428 (N_11428,N_11247,N_11348);
and U11429 (N_11429,N_11375,N_11254);
nor U11430 (N_11430,N_11327,N_11246);
nand U11431 (N_11431,N_11212,N_11292);
nor U11432 (N_11432,N_11356,N_11396);
nand U11433 (N_11433,N_11319,N_11262);
and U11434 (N_11434,N_11380,N_11237);
nand U11435 (N_11435,N_11209,N_11379);
and U11436 (N_11436,N_11296,N_11294);
xnor U11437 (N_11437,N_11390,N_11217);
nand U11438 (N_11438,N_11372,N_11220);
or U11439 (N_11439,N_11245,N_11310);
or U11440 (N_11440,N_11321,N_11383);
nand U11441 (N_11441,N_11257,N_11268);
nand U11442 (N_11442,N_11259,N_11213);
xnor U11443 (N_11443,N_11234,N_11341);
or U11444 (N_11444,N_11278,N_11244);
xor U11445 (N_11445,N_11256,N_11300);
or U11446 (N_11446,N_11276,N_11399);
nand U11447 (N_11447,N_11303,N_11343);
or U11448 (N_11448,N_11347,N_11323);
nand U11449 (N_11449,N_11208,N_11362);
nand U11450 (N_11450,N_11302,N_11353);
nor U11451 (N_11451,N_11214,N_11295);
xor U11452 (N_11452,N_11368,N_11222);
nand U11453 (N_11453,N_11357,N_11219);
nand U11454 (N_11454,N_11307,N_11287);
xnor U11455 (N_11455,N_11270,N_11305);
nor U11456 (N_11456,N_11381,N_11395);
nand U11457 (N_11457,N_11334,N_11255);
and U11458 (N_11458,N_11299,N_11297);
or U11459 (N_11459,N_11393,N_11377);
or U11460 (N_11460,N_11322,N_11240);
nor U11461 (N_11461,N_11206,N_11211);
nand U11462 (N_11462,N_11361,N_11324);
xor U11463 (N_11463,N_11369,N_11283);
xor U11464 (N_11464,N_11316,N_11267);
nor U11465 (N_11465,N_11232,N_11201);
nand U11466 (N_11466,N_11387,N_11338);
nor U11467 (N_11467,N_11210,N_11326);
xor U11468 (N_11468,N_11228,N_11376);
and U11469 (N_11469,N_11225,N_11272);
nor U11470 (N_11470,N_11370,N_11318);
nand U11471 (N_11471,N_11227,N_11238);
and U11472 (N_11472,N_11365,N_11374);
nor U11473 (N_11473,N_11271,N_11223);
nand U11474 (N_11474,N_11386,N_11279);
nor U11475 (N_11475,N_11258,N_11358);
xnor U11476 (N_11476,N_11229,N_11320);
xnor U11477 (N_11477,N_11371,N_11274);
nand U11478 (N_11478,N_11311,N_11398);
xnor U11479 (N_11479,N_11285,N_11282);
or U11480 (N_11480,N_11373,N_11355);
nor U11481 (N_11481,N_11382,N_11266);
or U11482 (N_11482,N_11249,N_11207);
nand U11483 (N_11483,N_11352,N_11328);
or U11484 (N_11484,N_11325,N_11275);
nor U11485 (N_11485,N_11204,N_11389);
or U11486 (N_11486,N_11236,N_11224);
xor U11487 (N_11487,N_11349,N_11235);
xnor U11488 (N_11488,N_11253,N_11333);
xor U11489 (N_11489,N_11248,N_11342);
nor U11490 (N_11490,N_11221,N_11277);
xor U11491 (N_11491,N_11304,N_11346);
xor U11492 (N_11492,N_11366,N_11359);
xor U11493 (N_11493,N_11284,N_11394);
nor U11494 (N_11494,N_11216,N_11203);
nand U11495 (N_11495,N_11306,N_11261);
nand U11496 (N_11496,N_11354,N_11335);
xor U11497 (N_11497,N_11397,N_11239);
xor U11498 (N_11498,N_11231,N_11293);
nor U11499 (N_11499,N_11242,N_11264);
and U11500 (N_11500,N_11255,N_11262);
and U11501 (N_11501,N_11352,N_11207);
and U11502 (N_11502,N_11207,N_11363);
nand U11503 (N_11503,N_11286,N_11291);
xor U11504 (N_11504,N_11331,N_11378);
and U11505 (N_11505,N_11293,N_11365);
nand U11506 (N_11506,N_11246,N_11383);
and U11507 (N_11507,N_11236,N_11305);
nand U11508 (N_11508,N_11347,N_11339);
nor U11509 (N_11509,N_11277,N_11251);
or U11510 (N_11510,N_11235,N_11322);
or U11511 (N_11511,N_11254,N_11244);
nor U11512 (N_11512,N_11396,N_11231);
nor U11513 (N_11513,N_11367,N_11257);
and U11514 (N_11514,N_11247,N_11256);
or U11515 (N_11515,N_11263,N_11247);
nor U11516 (N_11516,N_11220,N_11244);
and U11517 (N_11517,N_11289,N_11315);
and U11518 (N_11518,N_11337,N_11309);
and U11519 (N_11519,N_11247,N_11391);
and U11520 (N_11520,N_11396,N_11386);
or U11521 (N_11521,N_11223,N_11348);
nor U11522 (N_11522,N_11378,N_11313);
xor U11523 (N_11523,N_11372,N_11270);
and U11524 (N_11524,N_11286,N_11371);
xor U11525 (N_11525,N_11355,N_11272);
xnor U11526 (N_11526,N_11366,N_11232);
and U11527 (N_11527,N_11354,N_11202);
xnor U11528 (N_11528,N_11258,N_11273);
and U11529 (N_11529,N_11213,N_11273);
and U11530 (N_11530,N_11370,N_11200);
xor U11531 (N_11531,N_11250,N_11318);
xor U11532 (N_11532,N_11274,N_11372);
nor U11533 (N_11533,N_11330,N_11357);
and U11534 (N_11534,N_11335,N_11247);
or U11535 (N_11535,N_11349,N_11353);
nand U11536 (N_11536,N_11356,N_11354);
nor U11537 (N_11537,N_11227,N_11338);
xor U11538 (N_11538,N_11256,N_11279);
nand U11539 (N_11539,N_11359,N_11369);
xor U11540 (N_11540,N_11370,N_11389);
nor U11541 (N_11541,N_11271,N_11292);
xor U11542 (N_11542,N_11321,N_11274);
xor U11543 (N_11543,N_11361,N_11242);
and U11544 (N_11544,N_11363,N_11262);
xnor U11545 (N_11545,N_11332,N_11306);
nor U11546 (N_11546,N_11258,N_11321);
and U11547 (N_11547,N_11237,N_11358);
nor U11548 (N_11548,N_11298,N_11339);
xnor U11549 (N_11549,N_11214,N_11301);
or U11550 (N_11550,N_11244,N_11305);
and U11551 (N_11551,N_11305,N_11357);
and U11552 (N_11552,N_11309,N_11390);
nor U11553 (N_11553,N_11304,N_11313);
and U11554 (N_11554,N_11385,N_11348);
and U11555 (N_11555,N_11310,N_11212);
nor U11556 (N_11556,N_11235,N_11299);
xnor U11557 (N_11557,N_11263,N_11343);
xnor U11558 (N_11558,N_11389,N_11244);
xnor U11559 (N_11559,N_11334,N_11248);
or U11560 (N_11560,N_11348,N_11317);
xor U11561 (N_11561,N_11233,N_11298);
or U11562 (N_11562,N_11371,N_11336);
and U11563 (N_11563,N_11213,N_11228);
nor U11564 (N_11564,N_11376,N_11321);
or U11565 (N_11565,N_11354,N_11309);
xnor U11566 (N_11566,N_11308,N_11363);
nand U11567 (N_11567,N_11235,N_11343);
or U11568 (N_11568,N_11245,N_11225);
nand U11569 (N_11569,N_11240,N_11253);
xor U11570 (N_11570,N_11254,N_11297);
or U11571 (N_11571,N_11223,N_11226);
or U11572 (N_11572,N_11250,N_11209);
xnor U11573 (N_11573,N_11211,N_11333);
or U11574 (N_11574,N_11342,N_11262);
xnor U11575 (N_11575,N_11365,N_11396);
nor U11576 (N_11576,N_11259,N_11343);
nand U11577 (N_11577,N_11288,N_11253);
nor U11578 (N_11578,N_11327,N_11361);
nand U11579 (N_11579,N_11379,N_11363);
and U11580 (N_11580,N_11284,N_11303);
xnor U11581 (N_11581,N_11367,N_11284);
or U11582 (N_11582,N_11246,N_11243);
nor U11583 (N_11583,N_11311,N_11229);
nor U11584 (N_11584,N_11272,N_11374);
and U11585 (N_11585,N_11323,N_11380);
nand U11586 (N_11586,N_11343,N_11365);
or U11587 (N_11587,N_11234,N_11306);
xor U11588 (N_11588,N_11200,N_11301);
xor U11589 (N_11589,N_11263,N_11274);
nand U11590 (N_11590,N_11270,N_11323);
xor U11591 (N_11591,N_11217,N_11319);
nor U11592 (N_11592,N_11214,N_11327);
and U11593 (N_11593,N_11385,N_11349);
and U11594 (N_11594,N_11362,N_11218);
nand U11595 (N_11595,N_11344,N_11290);
xor U11596 (N_11596,N_11251,N_11256);
or U11597 (N_11597,N_11250,N_11374);
and U11598 (N_11598,N_11265,N_11261);
nand U11599 (N_11599,N_11345,N_11304);
nand U11600 (N_11600,N_11577,N_11567);
nor U11601 (N_11601,N_11595,N_11543);
nand U11602 (N_11602,N_11488,N_11433);
and U11603 (N_11603,N_11439,N_11473);
or U11604 (N_11604,N_11479,N_11442);
xor U11605 (N_11605,N_11497,N_11568);
nand U11606 (N_11606,N_11574,N_11520);
nand U11607 (N_11607,N_11485,N_11592);
and U11608 (N_11608,N_11587,N_11448);
or U11609 (N_11609,N_11547,N_11416);
xnor U11610 (N_11610,N_11559,N_11452);
nor U11611 (N_11611,N_11459,N_11414);
xor U11612 (N_11612,N_11591,N_11598);
nor U11613 (N_11613,N_11594,N_11536);
and U11614 (N_11614,N_11447,N_11477);
nor U11615 (N_11615,N_11552,N_11496);
nor U11616 (N_11616,N_11461,N_11548);
and U11617 (N_11617,N_11537,N_11460);
or U11618 (N_11618,N_11554,N_11469);
xnor U11619 (N_11619,N_11407,N_11584);
nor U11620 (N_11620,N_11418,N_11464);
nand U11621 (N_11621,N_11405,N_11470);
nand U11622 (N_11622,N_11476,N_11489);
nand U11623 (N_11623,N_11572,N_11506);
nor U11624 (N_11624,N_11524,N_11504);
or U11625 (N_11625,N_11502,N_11486);
nor U11626 (N_11626,N_11453,N_11589);
xor U11627 (N_11627,N_11435,N_11495);
xnor U11628 (N_11628,N_11417,N_11474);
xor U11629 (N_11629,N_11432,N_11517);
nor U11630 (N_11630,N_11404,N_11492);
nor U11631 (N_11631,N_11560,N_11436);
and U11632 (N_11632,N_11534,N_11446);
or U11633 (N_11633,N_11586,N_11514);
and U11634 (N_11634,N_11593,N_11511);
xor U11635 (N_11635,N_11564,N_11523);
nand U11636 (N_11636,N_11541,N_11546);
and U11637 (N_11637,N_11531,N_11581);
and U11638 (N_11638,N_11599,N_11487);
or U11639 (N_11639,N_11565,N_11458);
or U11640 (N_11640,N_11408,N_11429);
and U11641 (N_11641,N_11467,N_11501);
nand U11642 (N_11642,N_11545,N_11409);
or U11643 (N_11643,N_11573,N_11519);
nor U11644 (N_11644,N_11510,N_11498);
nand U11645 (N_11645,N_11468,N_11596);
xnor U11646 (N_11646,N_11420,N_11438);
xor U11647 (N_11647,N_11553,N_11526);
and U11648 (N_11648,N_11580,N_11529);
nor U11649 (N_11649,N_11450,N_11507);
and U11650 (N_11650,N_11423,N_11579);
or U11651 (N_11651,N_11491,N_11430);
xnor U11652 (N_11652,N_11512,N_11426);
and U11653 (N_11653,N_11434,N_11535);
or U11654 (N_11654,N_11571,N_11411);
xor U11655 (N_11655,N_11466,N_11550);
nor U11656 (N_11656,N_11551,N_11406);
nor U11657 (N_11657,N_11578,N_11410);
nand U11658 (N_11658,N_11522,N_11576);
xnor U11659 (N_11659,N_11431,N_11413);
or U11660 (N_11660,N_11556,N_11437);
nand U11661 (N_11661,N_11482,N_11419);
nand U11662 (N_11662,N_11521,N_11451);
xnor U11663 (N_11663,N_11540,N_11490);
nand U11664 (N_11664,N_11494,N_11445);
and U11665 (N_11665,N_11500,N_11539);
or U11666 (N_11666,N_11528,N_11425);
or U11667 (N_11667,N_11582,N_11527);
or U11668 (N_11668,N_11525,N_11493);
nand U11669 (N_11669,N_11530,N_11538);
nor U11670 (N_11670,N_11428,N_11508);
or U11671 (N_11671,N_11457,N_11475);
nor U11672 (N_11672,N_11585,N_11484);
or U11673 (N_11673,N_11557,N_11505);
xor U11674 (N_11674,N_11561,N_11583);
or U11675 (N_11675,N_11481,N_11562);
nand U11676 (N_11676,N_11516,N_11400);
nor U11677 (N_11677,N_11518,N_11454);
and U11678 (N_11678,N_11421,N_11403);
and U11679 (N_11679,N_11499,N_11412);
xor U11680 (N_11680,N_11455,N_11462);
nand U11681 (N_11681,N_11509,N_11513);
and U11682 (N_11682,N_11597,N_11463);
or U11683 (N_11683,N_11503,N_11544);
nor U11684 (N_11684,N_11515,N_11588);
and U11685 (N_11685,N_11558,N_11533);
nor U11686 (N_11686,N_11449,N_11566);
nor U11687 (N_11687,N_11575,N_11563);
xor U11688 (N_11688,N_11415,N_11440);
xnor U11689 (N_11689,N_11480,N_11401);
nor U11690 (N_11690,N_11532,N_11424);
and U11691 (N_11691,N_11427,N_11443);
and U11692 (N_11692,N_11478,N_11590);
nor U11693 (N_11693,N_11483,N_11472);
and U11694 (N_11694,N_11569,N_11456);
xnor U11695 (N_11695,N_11444,N_11555);
nor U11696 (N_11696,N_11465,N_11402);
or U11697 (N_11697,N_11422,N_11542);
nand U11698 (N_11698,N_11441,N_11549);
and U11699 (N_11699,N_11570,N_11471);
or U11700 (N_11700,N_11594,N_11442);
nor U11701 (N_11701,N_11551,N_11401);
or U11702 (N_11702,N_11414,N_11409);
or U11703 (N_11703,N_11506,N_11524);
nand U11704 (N_11704,N_11447,N_11494);
and U11705 (N_11705,N_11580,N_11594);
and U11706 (N_11706,N_11427,N_11431);
or U11707 (N_11707,N_11572,N_11533);
and U11708 (N_11708,N_11475,N_11484);
and U11709 (N_11709,N_11521,N_11466);
or U11710 (N_11710,N_11482,N_11449);
nor U11711 (N_11711,N_11448,N_11585);
and U11712 (N_11712,N_11580,N_11467);
nand U11713 (N_11713,N_11501,N_11508);
and U11714 (N_11714,N_11475,N_11548);
or U11715 (N_11715,N_11489,N_11584);
nor U11716 (N_11716,N_11547,N_11498);
xnor U11717 (N_11717,N_11437,N_11467);
nor U11718 (N_11718,N_11524,N_11430);
or U11719 (N_11719,N_11592,N_11422);
and U11720 (N_11720,N_11582,N_11571);
nand U11721 (N_11721,N_11576,N_11445);
nor U11722 (N_11722,N_11414,N_11582);
xnor U11723 (N_11723,N_11410,N_11591);
nor U11724 (N_11724,N_11462,N_11540);
and U11725 (N_11725,N_11482,N_11405);
nand U11726 (N_11726,N_11517,N_11527);
or U11727 (N_11727,N_11546,N_11556);
xor U11728 (N_11728,N_11548,N_11504);
nor U11729 (N_11729,N_11466,N_11495);
or U11730 (N_11730,N_11585,N_11413);
nor U11731 (N_11731,N_11424,N_11478);
nor U11732 (N_11732,N_11407,N_11484);
nand U11733 (N_11733,N_11420,N_11550);
or U11734 (N_11734,N_11419,N_11423);
or U11735 (N_11735,N_11443,N_11414);
xnor U11736 (N_11736,N_11531,N_11429);
nand U11737 (N_11737,N_11568,N_11476);
and U11738 (N_11738,N_11598,N_11405);
or U11739 (N_11739,N_11403,N_11565);
xnor U11740 (N_11740,N_11454,N_11540);
and U11741 (N_11741,N_11467,N_11517);
nor U11742 (N_11742,N_11571,N_11572);
nand U11743 (N_11743,N_11552,N_11537);
xor U11744 (N_11744,N_11453,N_11541);
nor U11745 (N_11745,N_11419,N_11593);
nand U11746 (N_11746,N_11533,N_11590);
and U11747 (N_11747,N_11574,N_11539);
and U11748 (N_11748,N_11446,N_11403);
nand U11749 (N_11749,N_11529,N_11425);
xnor U11750 (N_11750,N_11593,N_11592);
nand U11751 (N_11751,N_11561,N_11564);
and U11752 (N_11752,N_11434,N_11415);
nor U11753 (N_11753,N_11506,N_11410);
xor U11754 (N_11754,N_11420,N_11500);
xnor U11755 (N_11755,N_11432,N_11470);
and U11756 (N_11756,N_11515,N_11565);
and U11757 (N_11757,N_11569,N_11508);
xor U11758 (N_11758,N_11511,N_11519);
xor U11759 (N_11759,N_11410,N_11572);
xnor U11760 (N_11760,N_11470,N_11552);
or U11761 (N_11761,N_11412,N_11431);
or U11762 (N_11762,N_11578,N_11418);
or U11763 (N_11763,N_11535,N_11552);
xnor U11764 (N_11764,N_11561,N_11418);
nor U11765 (N_11765,N_11515,N_11594);
nand U11766 (N_11766,N_11536,N_11468);
nor U11767 (N_11767,N_11418,N_11572);
xor U11768 (N_11768,N_11471,N_11439);
xnor U11769 (N_11769,N_11534,N_11458);
and U11770 (N_11770,N_11518,N_11590);
and U11771 (N_11771,N_11437,N_11452);
xnor U11772 (N_11772,N_11497,N_11535);
or U11773 (N_11773,N_11599,N_11458);
and U11774 (N_11774,N_11492,N_11478);
or U11775 (N_11775,N_11526,N_11584);
nand U11776 (N_11776,N_11446,N_11524);
and U11777 (N_11777,N_11456,N_11579);
or U11778 (N_11778,N_11493,N_11481);
and U11779 (N_11779,N_11477,N_11559);
or U11780 (N_11780,N_11433,N_11410);
nand U11781 (N_11781,N_11568,N_11506);
or U11782 (N_11782,N_11596,N_11537);
nor U11783 (N_11783,N_11438,N_11424);
and U11784 (N_11784,N_11439,N_11420);
xor U11785 (N_11785,N_11437,N_11564);
nand U11786 (N_11786,N_11591,N_11438);
nor U11787 (N_11787,N_11428,N_11464);
xor U11788 (N_11788,N_11400,N_11591);
and U11789 (N_11789,N_11507,N_11573);
nor U11790 (N_11790,N_11431,N_11404);
nand U11791 (N_11791,N_11555,N_11523);
and U11792 (N_11792,N_11554,N_11427);
and U11793 (N_11793,N_11431,N_11491);
or U11794 (N_11794,N_11540,N_11486);
and U11795 (N_11795,N_11533,N_11485);
and U11796 (N_11796,N_11570,N_11413);
nor U11797 (N_11797,N_11566,N_11438);
and U11798 (N_11798,N_11535,N_11517);
and U11799 (N_11799,N_11550,N_11598);
or U11800 (N_11800,N_11764,N_11602);
nor U11801 (N_11801,N_11686,N_11648);
xnor U11802 (N_11802,N_11694,N_11754);
nor U11803 (N_11803,N_11612,N_11744);
nor U11804 (N_11804,N_11652,N_11734);
and U11805 (N_11805,N_11723,N_11700);
or U11806 (N_11806,N_11649,N_11758);
nor U11807 (N_11807,N_11607,N_11659);
or U11808 (N_11808,N_11742,N_11685);
xnor U11809 (N_11809,N_11730,N_11769);
nand U11810 (N_11810,N_11663,N_11753);
and U11811 (N_11811,N_11733,N_11710);
nor U11812 (N_11812,N_11795,N_11655);
or U11813 (N_11813,N_11782,N_11774);
nor U11814 (N_11814,N_11608,N_11615);
and U11815 (N_11815,N_11616,N_11731);
nand U11816 (N_11816,N_11631,N_11788);
nor U11817 (N_11817,N_11715,N_11633);
and U11818 (N_11818,N_11772,N_11737);
nand U11819 (N_11819,N_11746,N_11628);
nor U11820 (N_11820,N_11720,N_11722);
nor U11821 (N_11821,N_11667,N_11789);
or U11822 (N_11822,N_11683,N_11630);
nand U11823 (N_11823,N_11711,N_11791);
nand U11824 (N_11824,N_11752,N_11690);
nand U11825 (N_11825,N_11776,N_11678);
and U11826 (N_11826,N_11671,N_11665);
and U11827 (N_11827,N_11757,N_11747);
nand U11828 (N_11828,N_11674,N_11726);
and U11829 (N_11829,N_11799,N_11779);
or U11830 (N_11830,N_11728,N_11692);
xnor U11831 (N_11831,N_11705,N_11793);
nor U11832 (N_11832,N_11617,N_11716);
nand U11833 (N_11833,N_11637,N_11625);
nor U11834 (N_11834,N_11611,N_11677);
nand U11835 (N_11835,N_11698,N_11609);
nor U11836 (N_11836,N_11706,N_11691);
nor U11837 (N_11837,N_11697,N_11725);
nor U11838 (N_11838,N_11606,N_11729);
nor U11839 (N_11839,N_11664,N_11627);
or U11840 (N_11840,N_11778,N_11794);
nand U11841 (N_11841,N_11604,N_11661);
nand U11842 (N_11842,N_11651,N_11657);
or U11843 (N_11843,N_11721,N_11724);
and U11844 (N_11844,N_11750,N_11639);
xnor U11845 (N_11845,N_11626,N_11689);
nor U11846 (N_11846,N_11654,N_11695);
xor U11847 (N_11847,N_11727,N_11660);
and U11848 (N_11848,N_11708,N_11600);
and U11849 (N_11849,N_11636,N_11780);
xnor U11850 (N_11850,N_11714,N_11620);
and U11851 (N_11851,N_11634,N_11771);
nand U11852 (N_11852,N_11669,N_11783);
nor U11853 (N_11853,N_11703,N_11680);
xnor U11854 (N_11854,N_11638,N_11681);
or U11855 (N_11855,N_11653,N_11739);
and U11856 (N_11856,N_11621,N_11672);
nand U11857 (N_11857,N_11662,N_11658);
nand U11858 (N_11858,N_11673,N_11640);
and U11859 (N_11859,N_11601,N_11712);
nand U11860 (N_11860,N_11761,N_11688);
or U11861 (N_11861,N_11767,N_11696);
and U11862 (N_11862,N_11644,N_11777);
nor U11863 (N_11863,N_11699,N_11713);
nand U11864 (N_11864,N_11784,N_11798);
nand U11865 (N_11865,N_11781,N_11738);
nand U11866 (N_11866,N_11701,N_11676);
nand U11867 (N_11867,N_11745,N_11719);
or U11868 (N_11868,N_11785,N_11618);
or U11869 (N_11869,N_11770,N_11623);
nand U11870 (N_11870,N_11787,N_11635);
or U11871 (N_11871,N_11760,N_11763);
nand U11872 (N_11872,N_11736,N_11684);
xor U11873 (N_11873,N_11647,N_11650);
or U11874 (N_11874,N_11702,N_11632);
nand U11875 (N_11875,N_11741,N_11675);
xnor U11876 (N_11876,N_11666,N_11682);
and U11877 (N_11877,N_11624,N_11668);
or U11878 (N_11878,N_11796,N_11619);
xor U11879 (N_11879,N_11718,N_11646);
nand U11880 (N_11880,N_11622,N_11642);
xnor U11881 (N_11881,N_11749,N_11641);
xnor U11882 (N_11882,N_11786,N_11766);
or U11883 (N_11883,N_11740,N_11614);
xnor U11884 (N_11884,N_11709,N_11656);
or U11885 (N_11885,N_11704,N_11748);
nand U11886 (N_11886,N_11768,N_11645);
nor U11887 (N_11887,N_11679,N_11759);
and U11888 (N_11888,N_11687,N_11613);
or U11889 (N_11889,N_11773,N_11756);
or U11890 (N_11890,N_11629,N_11605);
xnor U11891 (N_11891,N_11610,N_11743);
or U11892 (N_11892,N_11790,N_11732);
or U11893 (N_11893,N_11755,N_11775);
nor U11894 (N_11894,N_11797,N_11643);
nor U11895 (N_11895,N_11603,N_11693);
or U11896 (N_11896,N_11670,N_11765);
nor U11897 (N_11897,N_11717,N_11762);
and U11898 (N_11898,N_11735,N_11707);
and U11899 (N_11899,N_11751,N_11792);
and U11900 (N_11900,N_11621,N_11774);
xor U11901 (N_11901,N_11731,N_11640);
or U11902 (N_11902,N_11615,N_11792);
or U11903 (N_11903,N_11633,N_11651);
xor U11904 (N_11904,N_11739,N_11707);
nand U11905 (N_11905,N_11653,N_11630);
and U11906 (N_11906,N_11792,N_11717);
or U11907 (N_11907,N_11700,N_11612);
and U11908 (N_11908,N_11739,N_11663);
xnor U11909 (N_11909,N_11715,N_11773);
nand U11910 (N_11910,N_11618,N_11717);
nand U11911 (N_11911,N_11738,N_11755);
xnor U11912 (N_11912,N_11673,N_11763);
or U11913 (N_11913,N_11691,N_11743);
or U11914 (N_11914,N_11743,N_11785);
and U11915 (N_11915,N_11636,N_11626);
or U11916 (N_11916,N_11620,N_11618);
nand U11917 (N_11917,N_11675,N_11652);
nor U11918 (N_11918,N_11615,N_11767);
nor U11919 (N_11919,N_11704,N_11721);
or U11920 (N_11920,N_11728,N_11619);
or U11921 (N_11921,N_11761,N_11615);
and U11922 (N_11922,N_11685,N_11771);
and U11923 (N_11923,N_11756,N_11743);
nor U11924 (N_11924,N_11710,N_11657);
xnor U11925 (N_11925,N_11746,N_11659);
nand U11926 (N_11926,N_11669,N_11772);
nor U11927 (N_11927,N_11637,N_11719);
and U11928 (N_11928,N_11685,N_11647);
nand U11929 (N_11929,N_11766,N_11709);
or U11930 (N_11930,N_11755,N_11625);
nor U11931 (N_11931,N_11705,N_11784);
or U11932 (N_11932,N_11715,N_11603);
or U11933 (N_11933,N_11707,N_11706);
and U11934 (N_11934,N_11612,N_11662);
or U11935 (N_11935,N_11780,N_11616);
nor U11936 (N_11936,N_11638,N_11616);
nand U11937 (N_11937,N_11640,N_11683);
nand U11938 (N_11938,N_11767,N_11742);
or U11939 (N_11939,N_11648,N_11673);
and U11940 (N_11940,N_11643,N_11737);
nor U11941 (N_11941,N_11628,N_11752);
or U11942 (N_11942,N_11713,N_11774);
xor U11943 (N_11943,N_11623,N_11761);
nor U11944 (N_11944,N_11795,N_11684);
xor U11945 (N_11945,N_11614,N_11611);
or U11946 (N_11946,N_11617,N_11638);
xor U11947 (N_11947,N_11643,N_11686);
or U11948 (N_11948,N_11716,N_11793);
nor U11949 (N_11949,N_11630,N_11680);
nand U11950 (N_11950,N_11727,N_11771);
xnor U11951 (N_11951,N_11654,N_11665);
nor U11952 (N_11952,N_11704,N_11668);
xnor U11953 (N_11953,N_11665,N_11726);
or U11954 (N_11954,N_11624,N_11700);
nand U11955 (N_11955,N_11617,N_11674);
xnor U11956 (N_11956,N_11693,N_11610);
xor U11957 (N_11957,N_11716,N_11633);
nor U11958 (N_11958,N_11641,N_11745);
nand U11959 (N_11959,N_11676,N_11641);
or U11960 (N_11960,N_11620,N_11743);
nor U11961 (N_11961,N_11654,N_11786);
nand U11962 (N_11962,N_11704,N_11628);
and U11963 (N_11963,N_11776,N_11642);
nor U11964 (N_11964,N_11666,N_11728);
nor U11965 (N_11965,N_11602,N_11615);
or U11966 (N_11966,N_11624,N_11796);
and U11967 (N_11967,N_11637,N_11796);
and U11968 (N_11968,N_11684,N_11738);
nand U11969 (N_11969,N_11736,N_11727);
or U11970 (N_11970,N_11793,N_11711);
nand U11971 (N_11971,N_11770,N_11632);
nor U11972 (N_11972,N_11795,N_11617);
xor U11973 (N_11973,N_11758,N_11620);
nor U11974 (N_11974,N_11694,N_11757);
or U11975 (N_11975,N_11701,N_11703);
nor U11976 (N_11976,N_11680,N_11762);
and U11977 (N_11977,N_11769,N_11676);
nor U11978 (N_11978,N_11635,N_11609);
nand U11979 (N_11979,N_11617,N_11759);
or U11980 (N_11980,N_11762,N_11771);
and U11981 (N_11981,N_11659,N_11709);
nand U11982 (N_11982,N_11675,N_11747);
nor U11983 (N_11983,N_11715,N_11769);
and U11984 (N_11984,N_11734,N_11621);
and U11985 (N_11985,N_11629,N_11696);
xnor U11986 (N_11986,N_11680,N_11726);
and U11987 (N_11987,N_11617,N_11753);
nand U11988 (N_11988,N_11687,N_11725);
xor U11989 (N_11989,N_11745,N_11741);
and U11990 (N_11990,N_11609,N_11662);
nor U11991 (N_11991,N_11690,N_11778);
or U11992 (N_11992,N_11631,N_11611);
nand U11993 (N_11993,N_11715,N_11600);
or U11994 (N_11994,N_11711,N_11695);
and U11995 (N_11995,N_11777,N_11627);
nor U11996 (N_11996,N_11700,N_11726);
nor U11997 (N_11997,N_11674,N_11701);
or U11998 (N_11998,N_11759,N_11652);
nor U11999 (N_11999,N_11784,N_11679);
xor U12000 (N_12000,N_11882,N_11844);
xor U12001 (N_12001,N_11933,N_11902);
xnor U12002 (N_12002,N_11818,N_11929);
nand U12003 (N_12003,N_11889,N_11891);
nand U12004 (N_12004,N_11941,N_11864);
nor U12005 (N_12005,N_11953,N_11972);
nor U12006 (N_12006,N_11861,N_11813);
nor U12007 (N_12007,N_11855,N_11955);
nor U12008 (N_12008,N_11870,N_11804);
nand U12009 (N_12009,N_11912,N_11852);
xor U12010 (N_12010,N_11971,N_11934);
or U12011 (N_12011,N_11998,N_11997);
nor U12012 (N_12012,N_11905,N_11806);
and U12013 (N_12013,N_11879,N_11896);
nand U12014 (N_12014,N_11915,N_11826);
xor U12015 (N_12015,N_11936,N_11932);
nor U12016 (N_12016,N_11994,N_11858);
xor U12017 (N_12017,N_11880,N_11982);
or U12018 (N_12018,N_11974,N_11989);
or U12019 (N_12019,N_11931,N_11970);
xor U12020 (N_12020,N_11916,N_11837);
or U12021 (N_12021,N_11897,N_11845);
nand U12022 (N_12022,N_11963,N_11860);
nor U12023 (N_12023,N_11903,N_11962);
nor U12024 (N_12024,N_11839,N_11831);
and U12025 (N_12025,N_11959,N_11978);
nor U12026 (N_12026,N_11807,N_11884);
xnor U12027 (N_12027,N_11908,N_11842);
nor U12028 (N_12028,N_11899,N_11816);
and U12029 (N_12029,N_11850,N_11853);
and U12030 (N_12030,N_11872,N_11995);
xor U12031 (N_12031,N_11980,N_11838);
and U12032 (N_12032,N_11814,N_11895);
nand U12033 (N_12033,N_11877,N_11996);
nand U12034 (N_12034,N_11938,N_11928);
xnor U12035 (N_12035,N_11825,N_11886);
xnor U12036 (N_12036,N_11913,N_11848);
nor U12037 (N_12037,N_11836,N_11904);
or U12038 (N_12038,N_11830,N_11801);
and U12039 (N_12039,N_11987,N_11948);
xor U12040 (N_12040,N_11986,N_11817);
or U12041 (N_12041,N_11820,N_11910);
nor U12042 (N_12042,N_11992,N_11883);
and U12043 (N_12043,N_11927,N_11835);
nor U12044 (N_12044,N_11893,N_11869);
or U12045 (N_12045,N_11873,N_11939);
nand U12046 (N_12046,N_11863,N_11800);
or U12047 (N_12047,N_11815,N_11828);
and U12048 (N_12048,N_11944,N_11930);
nand U12049 (N_12049,N_11876,N_11832);
xnor U12050 (N_12050,N_11950,N_11991);
and U12051 (N_12051,N_11921,N_11866);
xnor U12052 (N_12052,N_11984,N_11874);
or U12053 (N_12053,N_11849,N_11964);
or U12054 (N_12054,N_11812,N_11956);
nor U12055 (N_12055,N_11900,N_11990);
or U12056 (N_12056,N_11810,N_11957);
nand U12057 (N_12057,N_11887,N_11966);
nand U12058 (N_12058,N_11951,N_11942);
nor U12059 (N_12059,N_11811,N_11985);
nor U12060 (N_12060,N_11859,N_11829);
or U12061 (N_12061,N_11824,N_11952);
and U12062 (N_12062,N_11922,N_11803);
nor U12063 (N_12063,N_11923,N_11925);
nor U12064 (N_12064,N_11958,N_11988);
xnor U12065 (N_12065,N_11937,N_11878);
xor U12066 (N_12066,N_11965,N_11833);
and U12067 (N_12067,N_11917,N_11805);
nor U12068 (N_12068,N_11975,N_11862);
nor U12069 (N_12069,N_11808,N_11940);
xor U12070 (N_12070,N_11868,N_11834);
and U12071 (N_12071,N_11841,N_11907);
and U12072 (N_12072,N_11840,N_11802);
xnor U12073 (N_12073,N_11949,N_11976);
xor U12074 (N_12074,N_11892,N_11935);
nor U12075 (N_12075,N_11911,N_11926);
or U12076 (N_12076,N_11885,N_11827);
or U12077 (N_12077,N_11945,N_11865);
nand U12078 (N_12078,N_11888,N_11918);
and U12079 (N_12079,N_11822,N_11857);
and U12080 (N_12080,N_11909,N_11983);
xnor U12081 (N_12081,N_11809,N_11969);
nor U12082 (N_12082,N_11901,N_11960);
and U12083 (N_12083,N_11973,N_11920);
nand U12084 (N_12084,N_11890,N_11894);
or U12085 (N_12085,N_11914,N_11819);
and U12086 (N_12086,N_11854,N_11967);
or U12087 (N_12087,N_11856,N_11977);
nand U12088 (N_12088,N_11999,N_11871);
and U12089 (N_12089,N_11821,N_11875);
nand U12090 (N_12090,N_11924,N_11979);
xnor U12091 (N_12091,N_11943,N_11993);
and U12092 (N_12092,N_11898,N_11919);
xnor U12093 (N_12093,N_11823,N_11881);
xor U12094 (N_12094,N_11947,N_11846);
xor U12095 (N_12095,N_11867,N_11954);
nand U12096 (N_12096,N_11946,N_11961);
nand U12097 (N_12097,N_11981,N_11968);
xnor U12098 (N_12098,N_11843,N_11847);
and U12099 (N_12099,N_11906,N_11851);
and U12100 (N_12100,N_11953,N_11811);
nor U12101 (N_12101,N_11839,N_11822);
or U12102 (N_12102,N_11989,N_11821);
and U12103 (N_12103,N_11858,N_11901);
nand U12104 (N_12104,N_11891,N_11902);
and U12105 (N_12105,N_11836,N_11859);
or U12106 (N_12106,N_11908,N_11838);
xor U12107 (N_12107,N_11978,N_11808);
xor U12108 (N_12108,N_11980,N_11920);
nor U12109 (N_12109,N_11999,N_11864);
xor U12110 (N_12110,N_11913,N_11903);
or U12111 (N_12111,N_11889,N_11943);
nand U12112 (N_12112,N_11832,N_11985);
xnor U12113 (N_12113,N_11954,N_11914);
nor U12114 (N_12114,N_11925,N_11998);
xor U12115 (N_12115,N_11853,N_11910);
and U12116 (N_12116,N_11938,N_11959);
nor U12117 (N_12117,N_11983,N_11978);
xor U12118 (N_12118,N_11948,N_11922);
nor U12119 (N_12119,N_11846,N_11987);
or U12120 (N_12120,N_11904,N_11978);
and U12121 (N_12121,N_11888,N_11949);
nand U12122 (N_12122,N_11833,N_11815);
nor U12123 (N_12123,N_11856,N_11927);
xnor U12124 (N_12124,N_11978,N_11927);
nor U12125 (N_12125,N_11814,N_11931);
nand U12126 (N_12126,N_11954,N_11830);
nor U12127 (N_12127,N_11857,N_11927);
nand U12128 (N_12128,N_11980,N_11819);
and U12129 (N_12129,N_11926,N_11836);
nor U12130 (N_12130,N_11953,N_11963);
or U12131 (N_12131,N_11869,N_11905);
or U12132 (N_12132,N_11822,N_11937);
xnor U12133 (N_12133,N_11961,N_11890);
and U12134 (N_12134,N_11839,N_11832);
xnor U12135 (N_12135,N_11948,N_11927);
nor U12136 (N_12136,N_11910,N_11971);
nand U12137 (N_12137,N_11890,N_11906);
or U12138 (N_12138,N_11842,N_11855);
or U12139 (N_12139,N_11872,N_11964);
nand U12140 (N_12140,N_11817,N_11815);
nor U12141 (N_12141,N_11931,N_11831);
or U12142 (N_12142,N_11923,N_11936);
xor U12143 (N_12143,N_11892,N_11967);
xor U12144 (N_12144,N_11869,N_11979);
nand U12145 (N_12145,N_11837,N_11809);
nor U12146 (N_12146,N_11871,N_11835);
nor U12147 (N_12147,N_11908,N_11933);
xor U12148 (N_12148,N_11865,N_11825);
or U12149 (N_12149,N_11983,N_11880);
and U12150 (N_12150,N_11820,N_11911);
xor U12151 (N_12151,N_11987,N_11999);
or U12152 (N_12152,N_11866,N_11868);
and U12153 (N_12153,N_11863,N_11958);
nand U12154 (N_12154,N_11946,N_11860);
nand U12155 (N_12155,N_11968,N_11861);
nand U12156 (N_12156,N_11807,N_11890);
nor U12157 (N_12157,N_11868,N_11910);
and U12158 (N_12158,N_11953,N_11875);
xor U12159 (N_12159,N_11982,N_11893);
nor U12160 (N_12160,N_11988,N_11979);
and U12161 (N_12161,N_11964,N_11929);
nand U12162 (N_12162,N_11834,N_11920);
xor U12163 (N_12163,N_11868,N_11874);
nand U12164 (N_12164,N_11997,N_11866);
xor U12165 (N_12165,N_11933,N_11954);
and U12166 (N_12166,N_11856,N_11844);
and U12167 (N_12167,N_11811,N_11851);
xor U12168 (N_12168,N_11889,N_11952);
nand U12169 (N_12169,N_11972,N_11901);
or U12170 (N_12170,N_11985,N_11821);
xnor U12171 (N_12171,N_11984,N_11989);
xnor U12172 (N_12172,N_11802,N_11851);
nand U12173 (N_12173,N_11885,N_11914);
and U12174 (N_12174,N_11863,N_11917);
xor U12175 (N_12175,N_11970,N_11874);
and U12176 (N_12176,N_11904,N_11906);
nor U12177 (N_12177,N_11923,N_11894);
or U12178 (N_12178,N_11851,N_11866);
nand U12179 (N_12179,N_11994,N_11805);
and U12180 (N_12180,N_11956,N_11850);
or U12181 (N_12181,N_11985,N_11953);
nand U12182 (N_12182,N_11840,N_11862);
nor U12183 (N_12183,N_11965,N_11968);
and U12184 (N_12184,N_11951,N_11908);
nand U12185 (N_12185,N_11934,N_11983);
nor U12186 (N_12186,N_11938,N_11996);
xor U12187 (N_12187,N_11888,N_11908);
or U12188 (N_12188,N_11800,N_11804);
and U12189 (N_12189,N_11834,N_11975);
nor U12190 (N_12190,N_11832,N_11992);
and U12191 (N_12191,N_11869,N_11810);
and U12192 (N_12192,N_11896,N_11897);
and U12193 (N_12193,N_11977,N_11921);
xnor U12194 (N_12194,N_11826,N_11805);
xor U12195 (N_12195,N_11930,N_11895);
xor U12196 (N_12196,N_11841,N_11873);
nand U12197 (N_12197,N_11918,N_11903);
and U12198 (N_12198,N_11808,N_11831);
xnor U12199 (N_12199,N_11979,N_11822);
nand U12200 (N_12200,N_12149,N_12182);
and U12201 (N_12201,N_12067,N_12110);
nor U12202 (N_12202,N_12001,N_12195);
and U12203 (N_12203,N_12011,N_12117);
xnor U12204 (N_12204,N_12034,N_12090);
and U12205 (N_12205,N_12026,N_12124);
xor U12206 (N_12206,N_12078,N_12093);
xnor U12207 (N_12207,N_12048,N_12062);
xor U12208 (N_12208,N_12092,N_12105);
nand U12209 (N_12209,N_12169,N_12072);
nor U12210 (N_12210,N_12033,N_12080);
nand U12211 (N_12211,N_12100,N_12155);
nor U12212 (N_12212,N_12097,N_12039);
nor U12213 (N_12213,N_12133,N_12015);
or U12214 (N_12214,N_12004,N_12139);
xor U12215 (N_12215,N_12042,N_12055);
nor U12216 (N_12216,N_12088,N_12160);
xnor U12217 (N_12217,N_12016,N_12141);
and U12218 (N_12218,N_12157,N_12059);
or U12219 (N_12219,N_12057,N_12103);
and U12220 (N_12220,N_12044,N_12051);
nand U12221 (N_12221,N_12198,N_12163);
and U12222 (N_12222,N_12115,N_12021);
and U12223 (N_12223,N_12158,N_12084);
or U12224 (N_12224,N_12165,N_12036);
nand U12225 (N_12225,N_12164,N_12168);
and U12226 (N_12226,N_12031,N_12068);
and U12227 (N_12227,N_12076,N_12102);
nand U12228 (N_12228,N_12058,N_12003);
or U12229 (N_12229,N_12142,N_12073);
or U12230 (N_12230,N_12153,N_12049);
xnor U12231 (N_12231,N_12152,N_12188);
xor U12232 (N_12232,N_12178,N_12006);
nand U12233 (N_12233,N_12052,N_12099);
and U12234 (N_12234,N_12010,N_12104);
and U12235 (N_12235,N_12056,N_12184);
xnor U12236 (N_12236,N_12122,N_12009);
and U12237 (N_12237,N_12060,N_12189);
xor U12238 (N_12238,N_12079,N_12043);
nand U12239 (N_12239,N_12070,N_12064);
xor U12240 (N_12240,N_12180,N_12166);
nor U12241 (N_12241,N_12196,N_12111);
or U12242 (N_12242,N_12082,N_12173);
or U12243 (N_12243,N_12130,N_12136);
xor U12244 (N_12244,N_12063,N_12022);
and U12245 (N_12245,N_12192,N_12172);
and U12246 (N_12246,N_12114,N_12179);
and U12247 (N_12247,N_12131,N_12077);
nand U12248 (N_12248,N_12037,N_12095);
xnor U12249 (N_12249,N_12191,N_12113);
nor U12250 (N_12250,N_12125,N_12050);
nand U12251 (N_12251,N_12140,N_12106);
nor U12252 (N_12252,N_12197,N_12190);
and U12253 (N_12253,N_12002,N_12177);
xnor U12254 (N_12254,N_12066,N_12089);
nor U12255 (N_12255,N_12032,N_12135);
nand U12256 (N_12256,N_12129,N_12098);
and U12257 (N_12257,N_12096,N_12176);
nand U12258 (N_12258,N_12012,N_12126);
and U12259 (N_12259,N_12187,N_12101);
nand U12260 (N_12260,N_12083,N_12154);
xnor U12261 (N_12261,N_12123,N_12005);
or U12262 (N_12262,N_12150,N_12161);
nand U12263 (N_12263,N_12053,N_12132);
xor U12264 (N_12264,N_12019,N_12171);
or U12265 (N_12265,N_12075,N_12054);
xnor U12266 (N_12266,N_12027,N_12199);
xor U12267 (N_12267,N_12030,N_12108);
nand U12268 (N_12268,N_12038,N_12074);
xnor U12269 (N_12269,N_12156,N_12091);
nand U12270 (N_12270,N_12047,N_12109);
xor U12271 (N_12271,N_12146,N_12183);
nand U12272 (N_12272,N_12065,N_12008);
nand U12273 (N_12273,N_12167,N_12120);
or U12274 (N_12274,N_12061,N_12085);
xor U12275 (N_12275,N_12025,N_12000);
xor U12276 (N_12276,N_12181,N_12134);
xor U12277 (N_12277,N_12069,N_12045);
xor U12278 (N_12278,N_12071,N_12194);
nor U12279 (N_12279,N_12121,N_12023);
nand U12280 (N_12280,N_12143,N_12040);
nand U12281 (N_12281,N_12107,N_12175);
xnor U12282 (N_12282,N_12193,N_12013);
xor U12283 (N_12283,N_12170,N_12094);
and U12284 (N_12284,N_12128,N_12186);
and U12285 (N_12285,N_12116,N_12162);
nor U12286 (N_12286,N_12112,N_12028);
xor U12287 (N_12287,N_12138,N_12118);
and U12288 (N_12288,N_12029,N_12137);
or U12289 (N_12289,N_12147,N_12087);
or U12290 (N_12290,N_12127,N_12024);
nand U12291 (N_12291,N_12185,N_12041);
and U12292 (N_12292,N_12020,N_12081);
nand U12293 (N_12293,N_12017,N_12014);
xor U12294 (N_12294,N_12046,N_12159);
or U12295 (N_12295,N_12144,N_12148);
and U12296 (N_12296,N_12035,N_12007);
nand U12297 (N_12297,N_12145,N_12086);
xor U12298 (N_12298,N_12018,N_12151);
nor U12299 (N_12299,N_12174,N_12119);
nand U12300 (N_12300,N_12153,N_12005);
xor U12301 (N_12301,N_12059,N_12087);
nand U12302 (N_12302,N_12150,N_12115);
or U12303 (N_12303,N_12078,N_12166);
and U12304 (N_12304,N_12048,N_12179);
or U12305 (N_12305,N_12163,N_12130);
or U12306 (N_12306,N_12078,N_12086);
nand U12307 (N_12307,N_12051,N_12092);
or U12308 (N_12308,N_12112,N_12191);
and U12309 (N_12309,N_12054,N_12062);
nand U12310 (N_12310,N_12143,N_12071);
xor U12311 (N_12311,N_12190,N_12029);
xnor U12312 (N_12312,N_12112,N_12150);
nand U12313 (N_12313,N_12074,N_12088);
and U12314 (N_12314,N_12175,N_12046);
or U12315 (N_12315,N_12017,N_12110);
nor U12316 (N_12316,N_12169,N_12166);
xnor U12317 (N_12317,N_12011,N_12046);
xor U12318 (N_12318,N_12062,N_12149);
and U12319 (N_12319,N_12052,N_12122);
nor U12320 (N_12320,N_12081,N_12199);
xnor U12321 (N_12321,N_12133,N_12151);
or U12322 (N_12322,N_12021,N_12087);
nand U12323 (N_12323,N_12077,N_12093);
or U12324 (N_12324,N_12062,N_12129);
or U12325 (N_12325,N_12134,N_12192);
and U12326 (N_12326,N_12141,N_12168);
xnor U12327 (N_12327,N_12165,N_12153);
xor U12328 (N_12328,N_12061,N_12157);
and U12329 (N_12329,N_12067,N_12142);
nand U12330 (N_12330,N_12057,N_12114);
xnor U12331 (N_12331,N_12152,N_12047);
xnor U12332 (N_12332,N_12199,N_12192);
or U12333 (N_12333,N_12066,N_12125);
xnor U12334 (N_12334,N_12027,N_12104);
xnor U12335 (N_12335,N_12079,N_12021);
nand U12336 (N_12336,N_12011,N_12148);
nand U12337 (N_12337,N_12186,N_12076);
nand U12338 (N_12338,N_12141,N_12043);
xor U12339 (N_12339,N_12130,N_12190);
xor U12340 (N_12340,N_12089,N_12108);
or U12341 (N_12341,N_12148,N_12195);
nand U12342 (N_12342,N_12022,N_12047);
xnor U12343 (N_12343,N_12108,N_12175);
or U12344 (N_12344,N_12118,N_12097);
or U12345 (N_12345,N_12197,N_12154);
nor U12346 (N_12346,N_12081,N_12032);
xor U12347 (N_12347,N_12096,N_12138);
or U12348 (N_12348,N_12063,N_12080);
nand U12349 (N_12349,N_12065,N_12125);
and U12350 (N_12350,N_12096,N_12137);
nand U12351 (N_12351,N_12189,N_12086);
nand U12352 (N_12352,N_12048,N_12088);
or U12353 (N_12353,N_12140,N_12086);
nand U12354 (N_12354,N_12082,N_12098);
or U12355 (N_12355,N_12100,N_12193);
nor U12356 (N_12356,N_12081,N_12179);
nor U12357 (N_12357,N_12034,N_12078);
nor U12358 (N_12358,N_12147,N_12090);
nor U12359 (N_12359,N_12133,N_12191);
nor U12360 (N_12360,N_12129,N_12134);
and U12361 (N_12361,N_12037,N_12147);
or U12362 (N_12362,N_12108,N_12196);
nor U12363 (N_12363,N_12139,N_12037);
nor U12364 (N_12364,N_12040,N_12160);
and U12365 (N_12365,N_12039,N_12076);
and U12366 (N_12366,N_12172,N_12058);
xor U12367 (N_12367,N_12184,N_12032);
xnor U12368 (N_12368,N_12031,N_12109);
nand U12369 (N_12369,N_12168,N_12098);
xnor U12370 (N_12370,N_12196,N_12193);
xor U12371 (N_12371,N_12143,N_12094);
or U12372 (N_12372,N_12076,N_12013);
nor U12373 (N_12373,N_12128,N_12000);
and U12374 (N_12374,N_12184,N_12052);
nor U12375 (N_12375,N_12170,N_12186);
or U12376 (N_12376,N_12082,N_12106);
nand U12377 (N_12377,N_12159,N_12199);
nand U12378 (N_12378,N_12001,N_12164);
nand U12379 (N_12379,N_12089,N_12088);
nand U12380 (N_12380,N_12089,N_12046);
nand U12381 (N_12381,N_12017,N_12156);
nor U12382 (N_12382,N_12070,N_12131);
and U12383 (N_12383,N_12075,N_12066);
xnor U12384 (N_12384,N_12191,N_12101);
and U12385 (N_12385,N_12132,N_12072);
xnor U12386 (N_12386,N_12053,N_12168);
and U12387 (N_12387,N_12005,N_12128);
xor U12388 (N_12388,N_12006,N_12079);
nor U12389 (N_12389,N_12061,N_12108);
and U12390 (N_12390,N_12118,N_12079);
and U12391 (N_12391,N_12026,N_12052);
and U12392 (N_12392,N_12035,N_12071);
nor U12393 (N_12393,N_12096,N_12058);
xnor U12394 (N_12394,N_12045,N_12046);
or U12395 (N_12395,N_12070,N_12162);
nor U12396 (N_12396,N_12191,N_12081);
nand U12397 (N_12397,N_12098,N_12160);
and U12398 (N_12398,N_12035,N_12185);
nor U12399 (N_12399,N_12010,N_12038);
nand U12400 (N_12400,N_12203,N_12347);
xnor U12401 (N_12401,N_12229,N_12285);
and U12402 (N_12402,N_12294,N_12386);
nor U12403 (N_12403,N_12221,N_12371);
or U12404 (N_12404,N_12308,N_12339);
xor U12405 (N_12405,N_12303,N_12206);
or U12406 (N_12406,N_12233,N_12209);
or U12407 (N_12407,N_12291,N_12251);
or U12408 (N_12408,N_12354,N_12397);
nor U12409 (N_12409,N_12337,N_12280);
nand U12410 (N_12410,N_12292,N_12321);
xnor U12411 (N_12411,N_12326,N_12227);
nor U12412 (N_12412,N_12387,N_12356);
and U12413 (N_12413,N_12330,N_12357);
and U12414 (N_12414,N_12200,N_12346);
nand U12415 (N_12415,N_12317,N_12241);
xnor U12416 (N_12416,N_12263,N_12245);
nor U12417 (N_12417,N_12376,N_12299);
nor U12418 (N_12418,N_12364,N_12304);
or U12419 (N_12419,N_12231,N_12293);
xor U12420 (N_12420,N_12319,N_12223);
xor U12421 (N_12421,N_12323,N_12313);
or U12422 (N_12422,N_12315,N_12302);
nor U12423 (N_12423,N_12272,N_12248);
and U12424 (N_12424,N_12208,N_12342);
xnor U12425 (N_12425,N_12246,N_12320);
nor U12426 (N_12426,N_12290,N_12214);
or U12427 (N_12427,N_12332,N_12380);
and U12428 (N_12428,N_12382,N_12384);
xnor U12429 (N_12429,N_12211,N_12205);
or U12430 (N_12430,N_12295,N_12394);
xor U12431 (N_12431,N_12361,N_12358);
or U12432 (N_12432,N_12363,N_12232);
xor U12433 (N_12433,N_12207,N_12276);
xor U12434 (N_12434,N_12212,N_12262);
and U12435 (N_12435,N_12254,N_12389);
and U12436 (N_12436,N_12353,N_12228);
xor U12437 (N_12437,N_12238,N_12340);
and U12438 (N_12438,N_12213,N_12278);
or U12439 (N_12439,N_12283,N_12217);
xnor U12440 (N_12440,N_12219,N_12311);
xnor U12441 (N_12441,N_12268,N_12242);
xor U12442 (N_12442,N_12256,N_12329);
xnor U12443 (N_12443,N_12383,N_12252);
and U12444 (N_12444,N_12398,N_12350);
xnor U12445 (N_12445,N_12343,N_12282);
nor U12446 (N_12446,N_12348,N_12391);
nand U12447 (N_12447,N_12370,N_12388);
xnor U12448 (N_12448,N_12352,N_12393);
or U12449 (N_12449,N_12325,N_12239);
nor U12450 (N_12450,N_12267,N_12255);
nand U12451 (N_12451,N_12235,N_12333);
or U12452 (N_12452,N_12344,N_12345);
nor U12453 (N_12453,N_12234,N_12274);
or U12454 (N_12454,N_12281,N_12296);
and U12455 (N_12455,N_12368,N_12271);
nand U12456 (N_12456,N_12275,N_12374);
xnor U12457 (N_12457,N_12265,N_12286);
and U12458 (N_12458,N_12369,N_12381);
and U12459 (N_12459,N_12253,N_12301);
xor U12460 (N_12460,N_12392,N_12367);
xnor U12461 (N_12461,N_12316,N_12270);
or U12462 (N_12462,N_12355,N_12215);
or U12463 (N_12463,N_12377,N_12249);
xnor U12464 (N_12464,N_12372,N_12322);
nand U12465 (N_12465,N_12360,N_12247);
nand U12466 (N_12466,N_12266,N_12269);
or U12467 (N_12467,N_12351,N_12396);
nand U12468 (N_12468,N_12297,N_12264);
nor U12469 (N_12469,N_12279,N_12305);
xnor U12470 (N_12470,N_12273,N_12366);
and U12471 (N_12471,N_12373,N_12258);
and U12472 (N_12472,N_12257,N_12314);
xnor U12473 (N_12473,N_12220,N_12335);
xor U12474 (N_12474,N_12287,N_12338);
xor U12475 (N_12475,N_12378,N_12244);
xnor U12476 (N_12476,N_12390,N_12201);
or U12477 (N_12477,N_12327,N_12218);
and U12478 (N_12478,N_12222,N_12226);
xnor U12479 (N_12479,N_12243,N_12395);
nor U12480 (N_12480,N_12284,N_12230);
and U12481 (N_12481,N_12375,N_12341);
nand U12482 (N_12482,N_12204,N_12328);
and U12483 (N_12483,N_12362,N_12312);
nor U12484 (N_12484,N_12236,N_12216);
xnor U12485 (N_12485,N_12250,N_12306);
and U12486 (N_12486,N_12288,N_12225);
nand U12487 (N_12487,N_12260,N_12309);
nand U12488 (N_12488,N_12334,N_12379);
nand U12489 (N_12489,N_12359,N_12300);
nand U12490 (N_12490,N_12224,N_12210);
nor U12491 (N_12491,N_12237,N_12399);
nand U12492 (N_12492,N_12261,N_12318);
xnor U12493 (N_12493,N_12331,N_12259);
xor U12494 (N_12494,N_12240,N_12277);
or U12495 (N_12495,N_12289,N_12385);
and U12496 (N_12496,N_12349,N_12298);
xor U12497 (N_12497,N_12202,N_12365);
nand U12498 (N_12498,N_12324,N_12336);
nor U12499 (N_12499,N_12307,N_12310);
or U12500 (N_12500,N_12351,N_12264);
and U12501 (N_12501,N_12277,N_12347);
nand U12502 (N_12502,N_12277,N_12262);
and U12503 (N_12503,N_12387,N_12319);
nor U12504 (N_12504,N_12336,N_12300);
and U12505 (N_12505,N_12245,N_12364);
xnor U12506 (N_12506,N_12384,N_12372);
nor U12507 (N_12507,N_12361,N_12281);
and U12508 (N_12508,N_12209,N_12242);
and U12509 (N_12509,N_12275,N_12350);
xor U12510 (N_12510,N_12360,N_12380);
nand U12511 (N_12511,N_12373,N_12294);
xnor U12512 (N_12512,N_12340,N_12309);
xor U12513 (N_12513,N_12282,N_12363);
or U12514 (N_12514,N_12228,N_12217);
nor U12515 (N_12515,N_12261,N_12249);
nand U12516 (N_12516,N_12252,N_12216);
and U12517 (N_12517,N_12297,N_12353);
xor U12518 (N_12518,N_12227,N_12228);
and U12519 (N_12519,N_12249,N_12322);
and U12520 (N_12520,N_12258,N_12370);
and U12521 (N_12521,N_12371,N_12313);
nor U12522 (N_12522,N_12381,N_12366);
and U12523 (N_12523,N_12340,N_12307);
xor U12524 (N_12524,N_12356,N_12338);
nor U12525 (N_12525,N_12282,N_12339);
xor U12526 (N_12526,N_12329,N_12247);
nor U12527 (N_12527,N_12368,N_12213);
or U12528 (N_12528,N_12295,N_12313);
nor U12529 (N_12529,N_12298,N_12342);
and U12530 (N_12530,N_12376,N_12324);
xnor U12531 (N_12531,N_12210,N_12204);
or U12532 (N_12532,N_12289,N_12323);
xnor U12533 (N_12533,N_12311,N_12376);
or U12534 (N_12534,N_12326,N_12234);
xnor U12535 (N_12535,N_12211,N_12269);
xor U12536 (N_12536,N_12269,N_12341);
or U12537 (N_12537,N_12312,N_12341);
xnor U12538 (N_12538,N_12374,N_12236);
or U12539 (N_12539,N_12368,N_12319);
nor U12540 (N_12540,N_12343,N_12337);
and U12541 (N_12541,N_12376,N_12338);
or U12542 (N_12542,N_12352,N_12376);
or U12543 (N_12543,N_12222,N_12238);
or U12544 (N_12544,N_12280,N_12278);
or U12545 (N_12545,N_12336,N_12367);
or U12546 (N_12546,N_12359,N_12241);
nor U12547 (N_12547,N_12389,N_12226);
nor U12548 (N_12548,N_12383,N_12304);
xnor U12549 (N_12549,N_12226,N_12397);
and U12550 (N_12550,N_12328,N_12252);
xnor U12551 (N_12551,N_12372,N_12320);
or U12552 (N_12552,N_12227,N_12328);
nand U12553 (N_12553,N_12205,N_12343);
xor U12554 (N_12554,N_12282,N_12289);
nor U12555 (N_12555,N_12274,N_12363);
and U12556 (N_12556,N_12295,N_12260);
and U12557 (N_12557,N_12258,N_12226);
or U12558 (N_12558,N_12345,N_12395);
nor U12559 (N_12559,N_12348,N_12397);
and U12560 (N_12560,N_12263,N_12237);
xnor U12561 (N_12561,N_12289,N_12397);
xnor U12562 (N_12562,N_12266,N_12394);
and U12563 (N_12563,N_12331,N_12249);
or U12564 (N_12564,N_12301,N_12232);
nor U12565 (N_12565,N_12329,N_12239);
and U12566 (N_12566,N_12209,N_12320);
or U12567 (N_12567,N_12394,N_12339);
and U12568 (N_12568,N_12237,N_12246);
xor U12569 (N_12569,N_12274,N_12243);
and U12570 (N_12570,N_12342,N_12393);
nand U12571 (N_12571,N_12305,N_12351);
or U12572 (N_12572,N_12368,N_12389);
or U12573 (N_12573,N_12281,N_12327);
or U12574 (N_12574,N_12306,N_12243);
xnor U12575 (N_12575,N_12342,N_12233);
nor U12576 (N_12576,N_12245,N_12372);
and U12577 (N_12577,N_12242,N_12355);
nor U12578 (N_12578,N_12247,N_12333);
or U12579 (N_12579,N_12289,N_12279);
or U12580 (N_12580,N_12210,N_12306);
and U12581 (N_12581,N_12220,N_12306);
nor U12582 (N_12582,N_12380,N_12216);
xnor U12583 (N_12583,N_12308,N_12388);
or U12584 (N_12584,N_12210,N_12268);
nand U12585 (N_12585,N_12335,N_12380);
or U12586 (N_12586,N_12241,N_12295);
xor U12587 (N_12587,N_12376,N_12218);
nor U12588 (N_12588,N_12332,N_12251);
or U12589 (N_12589,N_12338,N_12224);
or U12590 (N_12590,N_12398,N_12202);
xor U12591 (N_12591,N_12331,N_12301);
nor U12592 (N_12592,N_12394,N_12345);
nor U12593 (N_12593,N_12312,N_12204);
nand U12594 (N_12594,N_12258,N_12280);
xnor U12595 (N_12595,N_12382,N_12220);
nor U12596 (N_12596,N_12349,N_12254);
and U12597 (N_12597,N_12334,N_12360);
xor U12598 (N_12598,N_12249,N_12209);
or U12599 (N_12599,N_12205,N_12326);
xnor U12600 (N_12600,N_12440,N_12486);
xnor U12601 (N_12601,N_12566,N_12434);
nand U12602 (N_12602,N_12436,N_12586);
or U12603 (N_12603,N_12521,N_12468);
or U12604 (N_12604,N_12430,N_12494);
nand U12605 (N_12605,N_12504,N_12551);
nand U12606 (N_12606,N_12533,N_12456);
nor U12607 (N_12607,N_12444,N_12499);
nor U12608 (N_12608,N_12505,N_12588);
xor U12609 (N_12609,N_12488,N_12482);
xnor U12610 (N_12610,N_12577,N_12584);
nor U12611 (N_12611,N_12596,N_12403);
nand U12612 (N_12612,N_12570,N_12498);
xor U12613 (N_12613,N_12483,N_12565);
xor U12614 (N_12614,N_12490,N_12473);
and U12615 (N_12615,N_12414,N_12575);
nor U12616 (N_12616,N_12464,N_12540);
or U12617 (N_12617,N_12478,N_12441);
or U12618 (N_12618,N_12510,N_12526);
nand U12619 (N_12619,N_12511,N_12453);
or U12620 (N_12620,N_12530,N_12563);
xnor U12621 (N_12621,N_12466,N_12479);
and U12622 (N_12622,N_12474,N_12514);
or U12623 (N_12623,N_12567,N_12472);
nand U12624 (N_12624,N_12568,N_12542);
nor U12625 (N_12625,N_12493,N_12562);
nor U12626 (N_12626,N_12475,N_12500);
or U12627 (N_12627,N_12572,N_12432);
and U12628 (N_12628,N_12413,N_12491);
and U12629 (N_12629,N_12412,N_12406);
and U12630 (N_12630,N_12560,N_12506);
or U12631 (N_12631,N_12467,N_12594);
nor U12632 (N_12632,N_12576,N_12582);
xnor U12633 (N_12633,N_12546,N_12559);
nor U12634 (N_12634,N_12503,N_12547);
xnor U12635 (N_12635,N_12548,N_12536);
and U12636 (N_12636,N_12497,N_12435);
and U12637 (N_12637,N_12543,N_12442);
nand U12638 (N_12638,N_12408,N_12420);
nor U12639 (N_12639,N_12476,N_12445);
nor U12640 (N_12640,N_12539,N_12553);
and U12641 (N_12641,N_12534,N_12524);
nand U12642 (N_12642,N_12465,N_12522);
or U12643 (N_12643,N_12496,N_12424);
nor U12644 (N_12644,N_12580,N_12470);
xor U12645 (N_12645,N_12404,N_12452);
nor U12646 (N_12646,N_12583,N_12592);
and U12647 (N_12647,N_12571,N_12449);
or U12648 (N_12648,N_12581,N_12431);
and U12649 (N_12649,N_12528,N_12595);
nor U12650 (N_12650,N_12425,N_12574);
nor U12651 (N_12651,N_12438,N_12558);
nor U12652 (N_12652,N_12512,N_12455);
or U12653 (N_12653,N_12489,N_12450);
xor U12654 (N_12654,N_12597,N_12411);
and U12655 (N_12655,N_12421,N_12516);
and U12656 (N_12656,N_12532,N_12599);
and U12657 (N_12657,N_12459,N_12417);
xnor U12658 (N_12658,N_12477,N_12587);
or U12659 (N_12659,N_12419,N_12518);
and U12660 (N_12660,N_12537,N_12561);
xnor U12661 (N_12661,N_12578,N_12585);
or U12662 (N_12662,N_12429,N_12550);
and U12663 (N_12663,N_12555,N_12422);
xnor U12664 (N_12664,N_12531,N_12400);
or U12665 (N_12665,N_12525,N_12485);
and U12666 (N_12666,N_12454,N_12437);
or U12667 (N_12667,N_12527,N_12469);
xor U12668 (N_12668,N_12535,N_12593);
and U12669 (N_12669,N_12507,N_12589);
nor U12670 (N_12670,N_12463,N_12579);
xnor U12671 (N_12671,N_12538,N_12502);
nor U12672 (N_12672,N_12428,N_12443);
nor U12673 (N_12673,N_12448,N_12509);
or U12674 (N_12674,N_12515,N_12549);
and U12675 (N_12675,N_12405,N_12544);
nor U12676 (N_12676,N_12554,N_12492);
nand U12677 (N_12677,N_12426,N_12591);
xnor U12678 (N_12678,N_12402,N_12520);
nand U12679 (N_12679,N_12458,N_12541);
or U12680 (N_12680,N_12461,N_12401);
or U12681 (N_12681,N_12556,N_12484);
nand U12682 (N_12682,N_12590,N_12598);
or U12683 (N_12683,N_12487,N_12407);
xor U12684 (N_12684,N_12508,N_12415);
or U12685 (N_12685,N_12471,N_12557);
nor U12686 (N_12686,N_12439,N_12427);
nor U12687 (N_12687,N_12501,N_12573);
nor U12688 (N_12688,N_12418,N_12529);
xor U12689 (N_12689,N_12552,N_12460);
nor U12690 (N_12690,N_12446,N_12517);
or U12691 (N_12691,N_12447,N_12513);
or U12692 (N_12692,N_12564,N_12433);
or U12693 (N_12693,N_12480,N_12519);
nand U12694 (N_12694,N_12523,N_12410);
or U12695 (N_12695,N_12451,N_12545);
nand U12696 (N_12696,N_12423,N_12495);
and U12697 (N_12697,N_12416,N_12409);
nand U12698 (N_12698,N_12569,N_12457);
nor U12699 (N_12699,N_12462,N_12481);
xor U12700 (N_12700,N_12448,N_12521);
xor U12701 (N_12701,N_12573,N_12489);
or U12702 (N_12702,N_12450,N_12477);
nor U12703 (N_12703,N_12421,N_12414);
nand U12704 (N_12704,N_12513,N_12449);
and U12705 (N_12705,N_12484,N_12412);
and U12706 (N_12706,N_12525,N_12591);
and U12707 (N_12707,N_12451,N_12535);
and U12708 (N_12708,N_12584,N_12422);
nand U12709 (N_12709,N_12522,N_12421);
nand U12710 (N_12710,N_12439,N_12476);
and U12711 (N_12711,N_12527,N_12483);
or U12712 (N_12712,N_12543,N_12445);
and U12713 (N_12713,N_12491,N_12415);
nand U12714 (N_12714,N_12447,N_12589);
or U12715 (N_12715,N_12543,N_12538);
nand U12716 (N_12716,N_12550,N_12463);
xor U12717 (N_12717,N_12554,N_12480);
nand U12718 (N_12718,N_12488,N_12475);
nand U12719 (N_12719,N_12450,N_12434);
nand U12720 (N_12720,N_12486,N_12476);
or U12721 (N_12721,N_12552,N_12479);
or U12722 (N_12722,N_12554,N_12442);
nor U12723 (N_12723,N_12439,N_12567);
and U12724 (N_12724,N_12469,N_12466);
nand U12725 (N_12725,N_12463,N_12519);
or U12726 (N_12726,N_12413,N_12545);
or U12727 (N_12727,N_12581,N_12567);
or U12728 (N_12728,N_12573,N_12520);
and U12729 (N_12729,N_12501,N_12420);
nor U12730 (N_12730,N_12444,N_12597);
nand U12731 (N_12731,N_12545,N_12508);
and U12732 (N_12732,N_12447,N_12500);
xor U12733 (N_12733,N_12508,N_12479);
or U12734 (N_12734,N_12400,N_12537);
nor U12735 (N_12735,N_12599,N_12566);
and U12736 (N_12736,N_12548,N_12497);
nor U12737 (N_12737,N_12434,N_12569);
nand U12738 (N_12738,N_12487,N_12511);
and U12739 (N_12739,N_12471,N_12444);
xnor U12740 (N_12740,N_12468,N_12479);
and U12741 (N_12741,N_12510,N_12422);
and U12742 (N_12742,N_12453,N_12430);
and U12743 (N_12743,N_12544,N_12515);
or U12744 (N_12744,N_12458,N_12570);
or U12745 (N_12745,N_12560,N_12539);
nand U12746 (N_12746,N_12580,N_12416);
xnor U12747 (N_12747,N_12513,N_12476);
or U12748 (N_12748,N_12461,N_12453);
nand U12749 (N_12749,N_12411,N_12529);
and U12750 (N_12750,N_12574,N_12583);
nand U12751 (N_12751,N_12570,N_12561);
or U12752 (N_12752,N_12400,N_12502);
xnor U12753 (N_12753,N_12532,N_12593);
or U12754 (N_12754,N_12574,N_12482);
and U12755 (N_12755,N_12499,N_12542);
or U12756 (N_12756,N_12540,N_12413);
or U12757 (N_12757,N_12568,N_12587);
nor U12758 (N_12758,N_12509,N_12553);
xor U12759 (N_12759,N_12474,N_12545);
xnor U12760 (N_12760,N_12579,N_12408);
nor U12761 (N_12761,N_12428,N_12466);
nor U12762 (N_12762,N_12554,N_12454);
and U12763 (N_12763,N_12418,N_12432);
nand U12764 (N_12764,N_12434,N_12523);
nand U12765 (N_12765,N_12470,N_12592);
or U12766 (N_12766,N_12583,N_12438);
xnor U12767 (N_12767,N_12458,N_12480);
nand U12768 (N_12768,N_12589,N_12584);
nand U12769 (N_12769,N_12503,N_12475);
xnor U12770 (N_12770,N_12576,N_12431);
xnor U12771 (N_12771,N_12543,N_12456);
nand U12772 (N_12772,N_12438,N_12453);
or U12773 (N_12773,N_12535,N_12463);
and U12774 (N_12774,N_12523,N_12532);
xor U12775 (N_12775,N_12524,N_12414);
or U12776 (N_12776,N_12571,N_12529);
and U12777 (N_12777,N_12541,N_12446);
nand U12778 (N_12778,N_12508,N_12482);
nand U12779 (N_12779,N_12522,N_12456);
nand U12780 (N_12780,N_12414,N_12528);
nor U12781 (N_12781,N_12435,N_12446);
nor U12782 (N_12782,N_12522,N_12523);
or U12783 (N_12783,N_12475,N_12508);
nand U12784 (N_12784,N_12411,N_12579);
xnor U12785 (N_12785,N_12429,N_12557);
or U12786 (N_12786,N_12472,N_12576);
and U12787 (N_12787,N_12465,N_12446);
or U12788 (N_12788,N_12579,N_12533);
nor U12789 (N_12789,N_12413,N_12456);
and U12790 (N_12790,N_12588,N_12461);
nand U12791 (N_12791,N_12590,N_12531);
or U12792 (N_12792,N_12453,N_12544);
or U12793 (N_12793,N_12544,N_12530);
nand U12794 (N_12794,N_12541,N_12410);
nand U12795 (N_12795,N_12458,N_12550);
and U12796 (N_12796,N_12568,N_12470);
nand U12797 (N_12797,N_12598,N_12445);
or U12798 (N_12798,N_12494,N_12596);
nor U12799 (N_12799,N_12546,N_12545);
and U12800 (N_12800,N_12634,N_12682);
or U12801 (N_12801,N_12605,N_12629);
or U12802 (N_12802,N_12707,N_12606);
or U12803 (N_12803,N_12701,N_12735);
and U12804 (N_12804,N_12759,N_12748);
xor U12805 (N_12805,N_12774,N_12658);
xnor U12806 (N_12806,N_12795,N_12616);
and U12807 (N_12807,N_12739,N_12790);
and U12808 (N_12808,N_12676,N_12679);
and U12809 (N_12809,N_12639,N_12665);
nor U12810 (N_12810,N_12675,N_12785);
or U12811 (N_12811,N_12733,N_12696);
nand U12812 (N_12812,N_12650,N_12670);
nor U12813 (N_12813,N_12793,N_12652);
nand U12814 (N_12814,N_12776,N_12613);
nand U12815 (N_12815,N_12602,N_12746);
or U12816 (N_12816,N_12643,N_12697);
nor U12817 (N_12817,N_12621,N_12797);
and U12818 (N_12818,N_12757,N_12778);
nor U12819 (N_12819,N_12612,N_12725);
and U12820 (N_12820,N_12702,N_12720);
nor U12821 (N_12821,N_12749,N_12711);
xnor U12822 (N_12822,N_12705,N_12763);
and U12823 (N_12823,N_12728,N_12719);
and U12824 (N_12824,N_12627,N_12635);
nand U12825 (N_12825,N_12661,N_12775);
and U12826 (N_12826,N_12656,N_12729);
xnor U12827 (N_12827,N_12773,N_12727);
nand U12828 (N_12828,N_12770,N_12768);
nor U12829 (N_12829,N_12710,N_12767);
or U12830 (N_12830,N_12653,N_12717);
nor U12831 (N_12831,N_12709,N_12601);
xnor U12832 (N_12832,N_12622,N_12743);
nor U12833 (N_12833,N_12692,N_12742);
xnor U12834 (N_12834,N_12654,N_12754);
xor U12835 (N_12835,N_12772,N_12794);
and U12836 (N_12836,N_12608,N_12699);
and U12837 (N_12837,N_12764,N_12698);
nand U12838 (N_12838,N_12642,N_12747);
xor U12839 (N_12839,N_12731,N_12766);
and U12840 (N_12840,N_12668,N_12657);
or U12841 (N_12841,N_12781,N_12730);
nor U12842 (N_12842,N_12726,N_12648);
nor U12843 (N_12843,N_12721,N_12760);
nand U12844 (N_12844,N_12600,N_12734);
nor U12845 (N_12845,N_12761,N_12779);
nand U12846 (N_12846,N_12674,N_12647);
nand U12847 (N_12847,N_12684,N_12644);
or U12848 (N_12848,N_12689,N_12669);
or U12849 (N_12849,N_12628,N_12737);
and U12850 (N_12850,N_12736,N_12706);
or U12851 (N_12851,N_12625,N_12704);
nand U12852 (N_12852,N_12751,N_12798);
nand U12853 (N_12853,N_12712,N_12695);
or U12854 (N_12854,N_12617,N_12789);
and U12855 (N_12855,N_12630,N_12660);
or U12856 (N_12856,N_12756,N_12672);
or U12857 (N_12857,N_12700,N_12690);
xor U12858 (N_12858,N_12620,N_12755);
and U12859 (N_12859,N_12791,N_12681);
xnor U12860 (N_12860,N_12632,N_12752);
xor U12861 (N_12861,N_12687,N_12640);
and U12862 (N_12862,N_12671,N_12666);
or U12863 (N_12863,N_12765,N_12744);
nand U12864 (N_12864,N_12784,N_12633);
nand U12865 (N_12865,N_12750,N_12673);
nor U12866 (N_12866,N_12718,N_12745);
nor U12867 (N_12867,N_12685,N_12615);
nor U12868 (N_12868,N_12655,N_12607);
nand U12869 (N_12869,N_12792,N_12771);
nor U12870 (N_12870,N_12663,N_12799);
nor U12871 (N_12871,N_12610,N_12762);
xor U12872 (N_12872,N_12740,N_12780);
xnor U12873 (N_12873,N_12667,N_12623);
xor U12874 (N_12874,N_12604,N_12787);
and U12875 (N_12875,N_12626,N_12686);
nor U12876 (N_12876,N_12732,N_12651);
nand U12877 (N_12877,N_12738,N_12715);
or U12878 (N_12878,N_12769,N_12724);
nand U12879 (N_12879,N_12624,N_12796);
or U12880 (N_12880,N_12788,N_12691);
nor U12881 (N_12881,N_12614,N_12645);
xor U12882 (N_12882,N_12693,N_12708);
nand U12883 (N_12883,N_12637,N_12619);
xnor U12884 (N_12884,N_12723,N_12680);
and U12885 (N_12885,N_12664,N_12683);
and U12886 (N_12886,N_12741,N_12758);
nand U12887 (N_12887,N_12659,N_12649);
nor U12888 (N_12888,N_12611,N_12694);
or U12889 (N_12889,N_12716,N_12777);
and U12890 (N_12890,N_12786,N_12646);
or U12891 (N_12891,N_12641,N_12722);
nand U12892 (N_12892,N_12713,N_12714);
nand U12893 (N_12893,N_12662,N_12753);
and U12894 (N_12894,N_12703,N_12609);
or U12895 (N_12895,N_12636,N_12631);
nor U12896 (N_12896,N_12783,N_12677);
xnor U12897 (N_12897,N_12782,N_12638);
nand U12898 (N_12898,N_12603,N_12688);
and U12899 (N_12899,N_12618,N_12678);
or U12900 (N_12900,N_12612,N_12687);
and U12901 (N_12901,N_12689,N_12769);
nor U12902 (N_12902,N_12716,N_12749);
nand U12903 (N_12903,N_12680,N_12699);
or U12904 (N_12904,N_12771,N_12615);
or U12905 (N_12905,N_12675,N_12767);
xnor U12906 (N_12906,N_12660,N_12770);
or U12907 (N_12907,N_12600,N_12664);
nand U12908 (N_12908,N_12710,N_12640);
and U12909 (N_12909,N_12683,N_12734);
nand U12910 (N_12910,N_12752,N_12711);
nand U12911 (N_12911,N_12705,N_12773);
and U12912 (N_12912,N_12765,N_12725);
nand U12913 (N_12913,N_12744,N_12715);
and U12914 (N_12914,N_12669,N_12716);
nand U12915 (N_12915,N_12767,N_12666);
nor U12916 (N_12916,N_12714,N_12672);
or U12917 (N_12917,N_12704,N_12684);
xor U12918 (N_12918,N_12793,N_12663);
or U12919 (N_12919,N_12746,N_12794);
xor U12920 (N_12920,N_12739,N_12706);
or U12921 (N_12921,N_12676,N_12693);
or U12922 (N_12922,N_12677,N_12644);
xor U12923 (N_12923,N_12729,N_12628);
xor U12924 (N_12924,N_12661,N_12672);
or U12925 (N_12925,N_12759,N_12694);
nor U12926 (N_12926,N_12613,N_12649);
and U12927 (N_12927,N_12744,N_12655);
xnor U12928 (N_12928,N_12680,N_12636);
xnor U12929 (N_12929,N_12712,N_12789);
nor U12930 (N_12930,N_12632,N_12666);
nand U12931 (N_12931,N_12738,N_12720);
and U12932 (N_12932,N_12603,N_12709);
or U12933 (N_12933,N_12627,N_12676);
xnor U12934 (N_12934,N_12785,N_12793);
nor U12935 (N_12935,N_12655,N_12634);
and U12936 (N_12936,N_12760,N_12798);
and U12937 (N_12937,N_12653,N_12654);
nor U12938 (N_12938,N_12752,N_12740);
nor U12939 (N_12939,N_12675,N_12691);
or U12940 (N_12940,N_12672,N_12716);
xor U12941 (N_12941,N_12688,N_12734);
xor U12942 (N_12942,N_12745,N_12630);
and U12943 (N_12943,N_12789,N_12630);
xnor U12944 (N_12944,N_12625,N_12784);
nand U12945 (N_12945,N_12603,N_12626);
nor U12946 (N_12946,N_12600,N_12724);
xor U12947 (N_12947,N_12660,N_12730);
nor U12948 (N_12948,N_12606,N_12790);
xnor U12949 (N_12949,N_12713,N_12696);
xnor U12950 (N_12950,N_12695,N_12788);
xnor U12951 (N_12951,N_12754,N_12687);
or U12952 (N_12952,N_12670,N_12633);
and U12953 (N_12953,N_12643,N_12637);
nor U12954 (N_12954,N_12641,N_12644);
nor U12955 (N_12955,N_12660,N_12782);
and U12956 (N_12956,N_12665,N_12780);
nor U12957 (N_12957,N_12657,N_12735);
and U12958 (N_12958,N_12720,N_12661);
nor U12959 (N_12959,N_12636,N_12691);
xnor U12960 (N_12960,N_12628,N_12614);
or U12961 (N_12961,N_12679,N_12605);
nand U12962 (N_12962,N_12661,N_12691);
nand U12963 (N_12963,N_12614,N_12706);
nor U12964 (N_12964,N_12624,N_12684);
xor U12965 (N_12965,N_12644,N_12797);
or U12966 (N_12966,N_12670,N_12635);
nor U12967 (N_12967,N_12689,N_12712);
and U12968 (N_12968,N_12636,N_12793);
nand U12969 (N_12969,N_12722,N_12755);
or U12970 (N_12970,N_12608,N_12683);
or U12971 (N_12971,N_12615,N_12710);
nor U12972 (N_12972,N_12673,N_12677);
nand U12973 (N_12973,N_12663,N_12642);
nor U12974 (N_12974,N_12791,N_12734);
or U12975 (N_12975,N_12706,N_12613);
xnor U12976 (N_12976,N_12698,N_12618);
and U12977 (N_12977,N_12643,N_12752);
nand U12978 (N_12978,N_12655,N_12769);
nand U12979 (N_12979,N_12673,N_12634);
or U12980 (N_12980,N_12780,N_12646);
or U12981 (N_12981,N_12772,N_12669);
or U12982 (N_12982,N_12621,N_12713);
xor U12983 (N_12983,N_12799,N_12678);
or U12984 (N_12984,N_12787,N_12775);
or U12985 (N_12985,N_12752,N_12658);
xnor U12986 (N_12986,N_12633,N_12678);
xor U12987 (N_12987,N_12749,N_12718);
nor U12988 (N_12988,N_12648,N_12683);
nor U12989 (N_12989,N_12621,N_12616);
nand U12990 (N_12990,N_12658,N_12702);
and U12991 (N_12991,N_12685,N_12787);
nor U12992 (N_12992,N_12779,N_12747);
xnor U12993 (N_12993,N_12767,N_12798);
xor U12994 (N_12994,N_12783,N_12738);
and U12995 (N_12995,N_12798,N_12678);
and U12996 (N_12996,N_12703,N_12732);
nand U12997 (N_12997,N_12773,N_12605);
and U12998 (N_12998,N_12785,N_12627);
or U12999 (N_12999,N_12764,N_12737);
xnor U13000 (N_13000,N_12973,N_12894);
nor U13001 (N_13001,N_12898,N_12999);
or U13002 (N_13002,N_12819,N_12873);
nand U13003 (N_13003,N_12804,N_12826);
nand U13004 (N_13004,N_12904,N_12803);
nor U13005 (N_13005,N_12981,N_12972);
nand U13006 (N_13006,N_12996,N_12947);
or U13007 (N_13007,N_12812,N_12860);
or U13008 (N_13008,N_12946,N_12995);
or U13009 (N_13009,N_12839,N_12871);
xnor U13010 (N_13010,N_12895,N_12950);
nand U13011 (N_13011,N_12892,N_12887);
or U13012 (N_13012,N_12901,N_12859);
or U13013 (N_13013,N_12925,N_12915);
nand U13014 (N_13014,N_12858,N_12814);
or U13015 (N_13015,N_12921,N_12962);
nand U13016 (N_13016,N_12936,N_12922);
xor U13017 (N_13017,N_12847,N_12951);
and U13018 (N_13018,N_12878,N_12868);
nor U13019 (N_13019,N_12993,N_12820);
or U13020 (N_13020,N_12834,N_12931);
or U13021 (N_13021,N_12919,N_12802);
nor U13022 (N_13022,N_12968,N_12940);
nor U13023 (N_13023,N_12982,N_12825);
and U13024 (N_13024,N_12964,N_12903);
and U13025 (N_13025,N_12914,N_12817);
xor U13026 (N_13026,N_12920,N_12877);
xnor U13027 (N_13027,N_12850,N_12913);
nand U13028 (N_13028,N_12998,N_12835);
xor U13029 (N_13029,N_12805,N_12852);
or U13030 (N_13030,N_12876,N_12935);
and U13031 (N_13031,N_12836,N_12821);
nand U13032 (N_13032,N_12864,N_12910);
or U13033 (N_13033,N_12917,N_12815);
xnor U13034 (N_13034,N_12854,N_12987);
and U13035 (N_13035,N_12843,N_12807);
nor U13036 (N_13036,N_12944,N_12879);
and U13037 (N_13037,N_12959,N_12934);
or U13038 (N_13038,N_12923,N_12984);
or U13039 (N_13039,N_12977,N_12908);
and U13040 (N_13040,N_12924,N_12853);
and U13041 (N_13041,N_12927,N_12845);
nor U13042 (N_13042,N_12960,N_12828);
xnor U13043 (N_13043,N_12969,N_12886);
nand U13044 (N_13044,N_12943,N_12875);
or U13045 (N_13045,N_12967,N_12811);
and U13046 (N_13046,N_12952,N_12884);
or U13047 (N_13047,N_12906,N_12856);
xor U13048 (N_13048,N_12932,N_12938);
and U13049 (N_13049,N_12928,N_12963);
xor U13050 (N_13050,N_12989,N_12986);
nor U13051 (N_13051,N_12861,N_12941);
or U13052 (N_13052,N_12958,N_12844);
nor U13053 (N_13053,N_12902,N_12867);
or U13054 (N_13054,N_12900,N_12907);
xnor U13055 (N_13055,N_12916,N_12889);
nor U13056 (N_13056,N_12945,N_12918);
xnor U13057 (N_13057,N_12890,N_12991);
or U13058 (N_13058,N_12824,N_12905);
and U13059 (N_13059,N_12942,N_12840);
nor U13060 (N_13060,N_12830,N_12897);
or U13061 (N_13061,N_12975,N_12863);
nor U13062 (N_13062,N_12983,N_12809);
nand U13063 (N_13063,N_12926,N_12976);
xor U13064 (N_13064,N_12971,N_12985);
and U13065 (N_13065,N_12893,N_12988);
nand U13066 (N_13066,N_12891,N_12833);
xnor U13067 (N_13067,N_12888,N_12930);
or U13068 (N_13068,N_12937,N_12956);
nor U13069 (N_13069,N_12829,N_12912);
nand U13070 (N_13070,N_12979,N_12911);
xor U13071 (N_13071,N_12831,N_12955);
nand U13072 (N_13072,N_12992,N_12869);
nor U13073 (N_13073,N_12949,N_12827);
or U13074 (N_13074,N_12848,N_12881);
or U13075 (N_13075,N_12865,N_12841);
or U13076 (N_13076,N_12806,N_12896);
nor U13077 (N_13077,N_12980,N_12899);
or U13078 (N_13078,N_12933,N_12823);
nor U13079 (N_13079,N_12872,N_12965);
nor U13080 (N_13080,N_12882,N_12990);
xnor U13081 (N_13081,N_12961,N_12801);
nand U13082 (N_13082,N_12832,N_12810);
xnor U13083 (N_13083,N_12978,N_12885);
xor U13084 (N_13084,N_12966,N_12866);
or U13085 (N_13085,N_12883,N_12837);
nor U13086 (N_13086,N_12855,N_12870);
nor U13087 (N_13087,N_12857,N_12808);
xnor U13088 (N_13088,N_12997,N_12874);
nand U13089 (N_13089,N_12957,N_12851);
xor U13090 (N_13090,N_12846,N_12880);
nor U13091 (N_13091,N_12929,N_12842);
nand U13092 (N_13092,N_12909,N_12953);
xor U13093 (N_13093,N_12818,N_12822);
or U13094 (N_13094,N_12994,N_12800);
and U13095 (N_13095,N_12813,N_12939);
nor U13096 (N_13096,N_12970,N_12838);
or U13097 (N_13097,N_12954,N_12948);
nand U13098 (N_13098,N_12862,N_12849);
nor U13099 (N_13099,N_12816,N_12974);
nor U13100 (N_13100,N_12832,N_12941);
or U13101 (N_13101,N_12806,N_12909);
nand U13102 (N_13102,N_12966,N_12996);
and U13103 (N_13103,N_12993,N_12848);
xnor U13104 (N_13104,N_12806,N_12874);
and U13105 (N_13105,N_12838,N_12902);
nand U13106 (N_13106,N_12942,N_12828);
and U13107 (N_13107,N_12970,N_12864);
and U13108 (N_13108,N_12808,N_12992);
nor U13109 (N_13109,N_12835,N_12873);
nor U13110 (N_13110,N_12905,N_12912);
or U13111 (N_13111,N_12960,N_12987);
and U13112 (N_13112,N_12847,N_12882);
nor U13113 (N_13113,N_12842,N_12889);
xnor U13114 (N_13114,N_12827,N_12864);
or U13115 (N_13115,N_12929,N_12882);
or U13116 (N_13116,N_12972,N_12956);
xor U13117 (N_13117,N_12924,N_12824);
nand U13118 (N_13118,N_12920,N_12858);
or U13119 (N_13119,N_12844,N_12839);
xor U13120 (N_13120,N_12844,N_12823);
xor U13121 (N_13121,N_12984,N_12840);
or U13122 (N_13122,N_12886,N_12883);
and U13123 (N_13123,N_12964,N_12980);
nor U13124 (N_13124,N_12971,N_12836);
nor U13125 (N_13125,N_12959,N_12970);
and U13126 (N_13126,N_12882,N_12986);
or U13127 (N_13127,N_12848,N_12906);
xnor U13128 (N_13128,N_12946,N_12987);
xnor U13129 (N_13129,N_12991,N_12830);
and U13130 (N_13130,N_12859,N_12858);
and U13131 (N_13131,N_12985,N_12837);
nand U13132 (N_13132,N_12868,N_12836);
nand U13133 (N_13133,N_12937,N_12856);
nor U13134 (N_13134,N_12831,N_12990);
nor U13135 (N_13135,N_12868,N_12810);
or U13136 (N_13136,N_12983,N_12925);
or U13137 (N_13137,N_12829,N_12852);
or U13138 (N_13138,N_12953,N_12883);
xor U13139 (N_13139,N_12906,N_12973);
nor U13140 (N_13140,N_12862,N_12926);
and U13141 (N_13141,N_12988,N_12856);
or U13142 (N_13142,N_12907,N_12885);
nand U13143 (N_13143,N_12893,N_12815);
xnor U13144 (N_13144,N_12966,N_12995);
or U13145 (N_13145,N_12889,N_12920);
nor U13146 (N_13146,N_12906,N_12975);
and U13147 (N_13147,N_12966,N_12889);
or U13148 (N_13148,N_12903,N_12949);
xor U13149 (N_13149,N_12981,N_12915);
and U13150 (N_13150,N_12841,N_12896);
and U13151 (N_13151,N_12999,N_12936);
and U13152 (N_13152,N_12837,N_12838);
nor U13153 (N_13153,N_12874,N_12998);
or U13154 (N_13154,N_12822,N_12979);
xnor U13155 (N_13155,N_12968,N_12986);
or U13156 (N_13156,N_12819,N_12883);
or U13157 (N_13157,N_12957,N_12974);
nand U13158 (N_13158,N_12940,N_12866);
nor U13159 (N_13159,N_12917,N_12842);
or U13160 (N_13160,N_12839,N_12916);
xor U13161 (N_13161,N_12992,N_12856);
or U13162 (N_13162,N_12948,N_12971);
xor U13163 (N_13163,N_12941,N_12882);
and U13164 (N_13164,N_12989,N_12985);
or U13165 (N_13165,N_12848,N_12869);
nand U13166 (N_13166,N_12871,N_12834);
or U13167 (N_13167,N_12987,N_12967);
and U13168 (N_13168,N_12951,N_12880);
nand U13169 (N_13169,N_12861,N_12955);
xor U13170 (N_13170,N_12874,N_12832);
or U13171 (N_13171,N_12876,N_12968);
nor U13172 (N_13172,N_12816,N_12893);
and U13173 (N_13173,N_12959,N_12810);
and U13174 (N_13174,N_12814,N_12806);
or U13175 (N_13175,N_12894,N_12842);
nor U13176 (N_13176,N_12945,N_12806);
or U13177 (N_13177,N_12897,N_12851);
or U13178 (N_13178,N_12866,N_12899);
xor U13179 (N_13179,N_12825,N_12905);
nor U13180 (N_13180,N_12938,N_12889);
nor U13181 (N_13181,N_12862,N_12901);
xor U13182 (N_13182,N_12867,N_12943);
nand U13183 (N_13183,N_12936,N_12879);
and U13184 (N_13184,N_12888,N_12865);
nand U13185 (N_13185,N_12975,N_12917);
xnor U13186 (N_13186,N_12807,N_12815);
xor U13187 (N_13187,N_12860,N_12914);
nor U13188 (N_13188,N_12886,N_12811);
or U13189 (N_13189,N_12846,N_12964);
nand U13190 (N_13190,N_12838,N_12859);
nor U13191 (N_13191,N_12884,N_12969);
or U13192 (N_13192,N_12905,N_12931);
xor U13193 (N_13193,N_12873,N_12800);
nand U13194 (N_13194,N_12800,N_12911);
and U13195 (N_13195,N_12960,N_12817);
nor U13196 (N_13196,N_12949,N_12857);
nor U13197 (N_13197,N_12815,N_12872);
nor U13198 (N_13198,N_12905,N_12867);
and U13199 (N_13199,N_12998,N_12936);
and U13200 (N_13200,N_13142,N_13026);
nand U13201 (N_13201,N_13076,N_13048);
and U13202 (N_13202,N_13133,N_13006);
nand U13203 (N_13203,N_13135,N_13122);
nand U13204 (N_13204,N_13139,N_13127);
or U13205 (N_13205,N_13096,N_13137);
nor U13206 (N_13206,N_13020,N_13054);
and U13207 (N_13207,N_13077,N_13179);
xnor U13208 (N_13208,N_13154,N_13047);
or U13209 (N_13209,N_13007,N_13126);
and U13210 (N_13210,N_13101,N_13088);
nand U13211 (N_13211,N_13140,N_13146);
xor U13212 (N_13212,N_13198,N_13195);
nand U13213 (N_13213,N_13175,N_13163);
and U13214 (N_13214,N_13005,N_13090);
or U13215 (N_13215,N_13173,N_13015);
nor U13216 (N_13216,N_13080,N_13189);
nand U13217 (N_13217,N_13089,N_13143);
xor U13218 (N_13218,N_13147,N_13196);
and U13219 (N_13219,N_13068,N_13036);
nand U13220 (N_13220,N_13045,N_13069);
nor U13221 (N_13221,N_13149,N_13031);
nor U13222 (N_13222,N_13170,N_13115);
or U13223 (N_13223,N_13168,N_13158);
or U13224 (N_13224,N_13191,N_13114);
xnor U13225 (N_13225,N_13125,N_13060);
xor U13226 (N_13226,N_13017,N_13013);
nand U13227 (N_13227,N_13177,N_13082);
nor U13228 (N_13228,N_13197,N_13092);
xor U13229 (N_13229,N_13042,N_13009);
nor U13230 (N_13230,N_13072,N_13112);
nand U13231 (N_13231,N_13156,N_13152);
nand U13232 (N_13232,N_13117,N_13128);
nand U13233 (N_13233,N_13171,N_13008);
xor U13234 (N_13234,N_13085,N_13178);
nand U13235 (N_13235,N_13065,N_13040);
and U13236 (N_13236,N_13110,N_13098);
and U13237 (N_13237,N_13169,N_13130);
or U13238 (N_13238,N_13190,N_13049);
nand U13239 (N_13239,N_13061,N_13136);
nor U13240 (N_13240,N_13134,N_13186);
xnor U13241 (N_13241,N_13056,N_13001);
xnor U13242 (N_13242,N_13018,N_13183);
xnor U13243 (N_13243,N_13148,N_13162);
or U13244 (N_13244,N_13039,N_13166);
nand U13245 (N_13245,N_13097,N_13079);
nand U13246 (N_13246,N_13046,N_13035);
nand U13247 (N_13247,N_13103,N_13120);
nor U13248 (N_13248,N_13037,N_13022);
or U13249 (N_13249,N_13145,N_13073);
or U13250 (N_13250,N_13074,N_13144);
nor U13251 (N_13251,N_13104,N_13172);
nand U13252 (N_13252,N_13066,N_13093);
or U13253 (N_13253,N_13113,N_13021);
xnor U13254 (N_13254,N_13107,N_13188);
xor U13255 (N_13255,N_13185,N_13019);
or U13256 (N_13256,N_13192,N_13083);
xor U13257 (N_13257,N_13161,N_13062);
and U13258 (N_13258,N_13091,N_13153);
and U13259 (N_13259,N_13105,N_13164);
nor U13260 (N_13260,N_13086,N_13160);
nand U13261 (N_13261,N_13029,N_13123);
and U13262 (N_13262,N_13027,N_13051);
nand U13263 (N_13263,N_13155,N_13067);
and U13264 (N_13264,N_13057,N_13167);
xnor U13265 (N_13265,N_13004,N_13011);
and U13266 (N_13266,N_13010,N_13059);
nor U13267 (N_13267,N_13071,N_13102);
nor U13268 (N_13268,N_13034,N_13180);
xnor U13269 (N_13269,N_13070,N_13014);
nor U13270 (N_13270,N_13041,N_13050);
xnor U13271 (N_13271,N_13028,N_13087);
xnor U13272 (N_13272,N_13199,N_13094);
and U13273 (N_13273,N_13174,N_13095);
nor U13274 (N_13274,N_13150,N_13032);
xor U13275 (N_13275,N_13184,N_13012);
nand U13276 (N_13276,N_13182,N_13159);
nand U13277 (N_13277,N_13165,N_13100);
xor U13278 (N_13278,N_13058,N_13081);
nor U13279 (N_13279,N_13024,N_13002);
xnor U13280 (N_13280,N_13118,N_13109);
nor U13281 (N_13281,N_13084,N_13078);
nand U13282 (N_13282,N_13193,N_13025);
or U13283 (N_13283,N_13003,N_13016);
nor U13284 (N_13284,N_13124,N_13055);
nand U13285 (N_13285,N_13063,N_13030);
nand U13286 (N_13286,N_13000,N_13038);
nor U13287 (N_13287,N_13157,N_13052);
and U13288 (N_13288,N_13194,N_13064);
xnor U13289 (N_13289,N_13151,N_13129);
nand U13290 (N_13290,N_13043,N_13044);
xnor U13291 (N_13291,N_13176,N_13106);
nand U13292 (N_13292,N_13181,N_13141);
nand U13293 (N_13293,N_13119,N_13111);
nand U13294 (N_13294,N_13132,N_13023);
or U13295 (N_13295,N_13121,N_13053);
xnor U13296 (N_13296,N_13131,N_13033);
nor U13297 (N_13297,N_13099,N_13187);
and U13298 (N_13298,N_13075,N_13116);
and U13299 (N_13299,N_13138,N_13108);
nand U13300 (N_13300,N_13024,N_13158);
or U13301 (N_13301,N_13174,N_13031);
and U13302 (N_13302,N_13104,N_13023);
xor U13303 (N_13303,N_13090,N_13158);
nor U13304 (N_13304,N_13157,N_13082);
and U13305 (N_13305,N_13148,N_13080);
xor U13306 (N_13306,N_13070,N_13085);
or U13307 (N_13307,N_13088,N_13095);
or U13308 (N_13308,N_13119,N_13151);
nor U13309 (N_13309,N_13127,N_13132);
or U13310 (N_13310,N_13046,N_13122);
nor U13311 (N_13311,N_13140,N_13083);
or U13312 (N_13312,N_13004,N_13179);
nor U13313 (N_13313,N_13050,N_13063);
nor U13314 (N_13314,N_13075,N_13055);
xnor U13315 (N_13315,N_13074,N_13187);
and U13316 (N_13316,N_13086,N_13051);
and U13317 (N_13317,N_13168,N_13172);
or U13318 (N_13318,N_13071,N_13158);
nand U13319 (N_13319,N_13074,N_13062);
nor U13320 (N_13320,N_13027,N_13064);
and U13321 (N_13321,N_13139,N_13115);
or U13322 (N_13322,N_13032,N_13005);
nand U13323 (N_13323,N_13000,N_13127);
and U13324 (N_13324,N_13101,N_13023);
or U13325 (N_13325,N_13075,N_13113);
and U13326 (N_13326,N_13000,N_13083);
nand U13327 (N_13327,N_13039,N_13125);
nor U13328 (N_13328,N_13001,N_13177);
or U13329 (N_13329,N_13060,N_13064);
xnor U13330 (N_13330,N_13094,N_13047);
xor U13331 (N_13331,N_13030,N_13038);
xor U13332 (N_13332,N_13133,N_13065);
xor U13333 (N_13333,N_13021,N_13071);
and U13334 (N_13334,N_13009,N_13121);
nand U13335 (N_13335,N_13136,N_13049);
xnor U13336 (N_13336,N_13000,N_13157);
or U13337 (N_13337,N_13030,N_13108);
nor U13338 (N_13338,N_13138,N_13117);
and U13339 (N_13339,N_13005,N_13080);
xnor U13340 (N_13340,N_13086,N_13059);
xnor U13341 (N_13341,N_13028,N_13142);
nor U13342 (N_13342,N_13023,N_13009);
xnor U13343 (N_13343,N_13161,N_13074);
or U13344 (N_13344,N_13035,N_13006);
xnor U13345 (N_13345,N_13145,N_13028);
xor U13346 (N_13346,N_13129,N_13058);
nand U13347 (N_13347,N_13154,N_13091);
and U13348 (N_13348,N_13024,N_13090);
nor U13349 (N_13349,N_13030,N_13090);
nor U13350 (N_13350,N_13139,N_13164);
or U13351 (N_13351,N_13161,N_13075);
or U13352 (N_13352,N_13166,N_13038);
nand U13353 (N_13353,N_13074,N_13124);
xor U13354 (N_13354,N_13030,N_13036);
nand U13355 (N_13355,N_13006,N_13040);
and U13356 (N_13356,N_13032,N_13182);
nand U13357 (N_13357,N_13083,N_13079);
xnor U13358 (N_13358,N_13100,N_13090);
nor U13359 (N_13359,N_13176,N_13099);
or U13360 (N_13360,N_13001,N_13180);
nand U13361 (N_13361,N_13076,N_13119);
xnor U13362 (N_13362,N_13105,N_13095);
xnor U13363 (N_13363,N_13165,N_13091);
and U13364 (N_13364,N_13159,N_13003);
nand U13365 (N_13365,N_13119,N_13051);
nor U13366 (N_13366,N_13177,N_13003);
nor U13367 (N_13367,N_13164,N_13067);
and U13368 (N_13368,N_13069,N_13164);
nand U13369 (N_13369,N_13004,N_13056);
or U13370 (N_13370,N_13156,N_13135);
or U13371 (N_13371,N_13197,N_13105);
nor U13372 (N_13372,N_13152,N_13002);
xnor U13373 (N_13373,N_13113,N_13006);
nand U13374 (N_13374,N_13108,N_13118);
xnor U13375 (N_13375,N_13043,N_13098);
xnor U13376 (N_13376,N_13019,N_13076);
nand U13377 (N_13377,N_13048,N_13103);
nand U13378 (N_13378,N_13112,N_13132);
or U13379 (N_13379,N_13037,N_13034);
or U13380 (N_13380,N_13166,N_13187);
xnor U13381 (N_13381,N_13185,N_13166);
or U13382 (N_13382,N_13024,N_13017);
and U13383 (N_13383,N_13033,N_13186);
xnor U13384 (N_13384,N_13074,N_13181);
xor U13385 (N_13385,N_13055,N_13169);
and U13386 (N_13386,N_13182,N_13188);
nand U13387 (N_13387,N_13029,N_13171);
nor U13388 (N_13388,N_13040,N_13094);
and U13389 (N_13389,N_13132,N_13104);
or U13390 (N_13390,N_13079,N_13055);
or U13391 (N_13391,N_13149,N_13111);
or U13392 (N_13392,N_13181,N_13190);
nand U13393 (N_13393,N_13060,N_13158);
nor U13394 (N_13394,N_13015,N_13192);
xnor U13395 (N_13395,N_13154,N_13017);
and U13396 (N_13396,N_13080,N_13104);
or U13397 (N_13397,N_13192,N_13001);
nor U13398 (N_13398,N_13081,N_13095);
and U13399 (N_13399,N_13109,N_13079);
or U13400 (N_13400,N_13317,N_13368);
xnor U13401 (N_13401,N_13216,N_13325);
nor U13402 (N_13402,N_13246,N_13241);
nor U13403 (N_13403,N_13383,N_13310);
nand U13404 (N_13404,N_13367,N_13307);
xor U13405 (N_13405,N_13303,N_13256);
nor U13406 (N_13406,N_13386,N_13362);
nor U13407 (N_13407,N_13334,N_13312);
or U13408 (N_13408,N_13295,N_13373);
xnor U13409 (N_13409,N_13332,N_13215);
nor U13410 (N_13410,N_13337,N_13340);
nor U13411 (N_13411,N_13287,N_13327);
nand U13412 (N_13412,N_13296,N_13207);
nor U13413 (N_13413,N_13231,N_13277);
and U13414 (N_13414,N_13224,N_13397);
or U13415 (N_13415,N_13262,N_13249);
nand U13416 (N_13416,N_13283,N_13343);
xnor U13417 (N_13417,N_13242,N_13211);
xor U13418 (N_13418,N_13350,N_13311);
and U13419 (N_13419,N_13274,N_13391);
nor U13420 (N_13420,N_13267,N_13285);
nand U13421 (N_13421,N_13387,N_13225);
and U13422 (N_13422,N_13230,N_13218);
xnor U13423 (N_13423,N_13339,N_13348);
or U13424 (N_13424,N_13321,N_13361);
xor U13425 (N_13425,N_13320,N_13359);
xnor U13426 (N_13426,N_13237,N_13375);
nand U13427 (N_13427,N_13390,N_13306);
and U13428 (N_13428,N_13253,N_13229);
nor U13429 (N_13429,N_13294,N_13245);
xor U13430 (N_13430,N_13379,N_13324);
or U13431 (N_13431,N_13369,N_13289);
or U13432 (N_13432,N_13202,N_13243);
or U13433 (N_13433,N_13316,N_13200);
and U13434 (N_13434,N_13349,N_13292);
or U13435 (N_13435,N_13214,N_13352);
xnor U13436 (N_13436,N_13353,N_13268);
nor U13437 (N_13437,N_13270,N_13220);
and U13438 (N_13438,N_13318,N_13331);
and U13439 (N_13439,N_13389,N_13226);
or U13440 (N_13440,N_13354,N_13210);
and U13441 (N_13441,N_13399,N_13261);
xnor U13442 (N_13442,N_13222,N_13258);
or U13443 (N_13443,N_13264,N_13382);
nand U13444 (N_13444,N_13356,N_13278);
nor U13445 (N_13445,N_13206,N_13263);
and U13446 (N_13446,N_13288,N_13205);
nor U13447 (N_13447,N_13333,N_13300);
nor U13448 (N_13448,N_13232,N_13279);
or U13449 (N_13449,N_13217,N_13355);
nand U13450 (N_13450,N_13384,N_13255);
and U13451 (N_13451,N_13351,N_13336);
and U13452 (N_13452,N_13203,N_13234);
nand U13453 (N_13453,N_13271,N_13315);
xor U13454 (N_13454,N_13358,N_13266);
xnor U13455 (N_13455,N_13260,N_13378);
or U13456 (N_13456,N_13385,N_13304);
nor U13457 (N_13457,N_13265,N_13366);
or U13458 (N_13458,N_13236,N_13290);
nor U13459 (N_13459,N_13344,N_13395);
and U13460 (N_13460,N_13301,N_13342);
nor U13461 (N_13461,N_13281,N_13212);
and U13462 (N_13462,N_13338,N_13370);
nand U13463 (N_13463,N_13345,N_13305);
nand U13464 (N_13464,N_13250,N_13347);
or U13465 (N_13465,N_13322,N_13233);
xnor U13466 (N_13466,N_13326,N_13377);
and U13467 (N_13467,N_13357,N_13364);
nor U13468 (N_13468,N_13394,N_13371);
and U13469 (N_13469,N_13247,N_13213);
nor U13470 (N_13470,N_13393,N_13269);
or U13471 (N_13471,N_13313,N_13376);
nor U13472 (N_13472,N_13341,N_13223);
or U13473 (N_13473,N_13240,N_13314);
or U13474 (N_13474,N_13208,N_13280);
or U13475 (N_13475,N_13286,N_13209);
nand U13476 (N_13476,N_13204,N_13330);
xor U13477 (N_13477,N_13259,N_13392);
xnor U13478 (N_13478,N_13282,N_13299);
xnor U13479 (N_13479,N_13238,N_13360);
nand U13480 (N_13480,N_13380,N_13276);
and U13481 (N_13481,N_13219,N_13248);
nor U13482 (N_13482,N_13346,N_13398);
and U13483 (N_13483,N_13388,N_13365);
and U13484 (N_13484,N_13323,N_13335);
nand U13485 (N_13485,N_13201,N_13329);
and U13486 (N_13486,N_13291,N_13244);
nand U13487 (N_13487,N_13275,N_13293);
and U13488 (N_13488,N_13235,N_13257);
nor U13489 (N_13489,N_13374,N_13273);
nor U13490 (N_13490,N_13272,N_13363);
and U13491 (N_13491,N_13251,N_13228);
xnor U13492 (N_13492,N_13298,N_13254);
nand U13493 (N_13493,N_13381,N_13227);
and U13494 (N_13494,N_13309,N_13328);
nor U13495 (N_13495,N_13252,N_13319);
nand U13496 (N_13496,N_13302,N_13221);
nor U13497 (N_13497,N_13297,N_13239);
or U13498 (N_13498,N_13396,N_13372);
and U13499 (N_13499,N_13284,N_13308);
nor U13500 (N_13500,N_13205,N_13289);
nor U13501 (N_13501,N_13383,N_13219);
or U13502 (N_13502,N_13315,N_13237);
nand U13503 (N_13503,N_13217,N_13398);
or U13504 (N_13504,N_13205,N_13245);
nand U13505 (N_13505,N_13340,N_13325);
and U13506 (N_13506,N_13201,N_13236);
nand U13507 (N_13507,N_13351,N_13330);
and U13508 (N_13508,N_13287,N_13285);
nand U13509 (N_13509,N_13368,N_13384);
or U13510 (N_13510,N_13246,N_13249);
and U13511 (N_13511,N_13348,N_13289);
and U13512 (N_13512,N_13288,N_13312);
or U13513 (N_13513,N_13274,N_13319);
xor U13514 (N_13514,N_13204,N_13248);
nand U13515 (N_13515,N_13386,N_13389);
or U13516 (N_13516,N_13324,N_13250);
and U13517 (N_13517,N_13222,N_13294);
and U13518 (N_13518,N_13342,N_13250);
nand U13519 (N_13519,N_13386,N_13244);
or U13520 (N_13520,N_13255,N_13207);
xor U13521 (N_13521,N_13390,N_13277);
xnor U13522 (N_13522,N_13294,N_13395);
xnor U13523 (N_13523,N_13348,N_13312);
nor U13524 (N_13524,N_13391,N_13345);
nor U13525 (N_13525,N_13334,N_13372);
nor U13526 (N_13526,N_13216,N_13203);
xnor U13527 (N_13527,N_13261,N_13379);
or U13528 (N_13528,N_13205,N_13298);
and U13529 (N_13529,N_13378,N_13294);
nand U13530 (N_13530,N_13261,N_13220);
xnor U13531 (N_13531,N_13312,N_13215);
and U13532 (N_13532,N_13344,N_13276);
nand U13533 (N_13533,N_13346,N_13367);
xor U13534 (N_13534,N_13227,N_13277);
nor U13535 (N_13535,N_13276,N_13361);
nor U13536 (N_13536,N_13318,N_13359);
and U13537 (N_13537,N_13303,N_13366);
or U13538 (N_13538,N_13310,N_13268);
and U13539 (N_13539,N_13385,N_13257);
xnor U13540 (N_13540,N_13239,N_13397);
nand U13541 (N_13541,N_13304,N_13273);
nor U13542 (N_13542,N_13389,N_13359);
nand U13543 (N_13543,N_13267,N_13380);
and U13544 (N_13544,N_13340,N_13324);
xor U13545 (N_13545,N_13296,N_13232);
nand U13546 (N_13546,N_13362,N_13397);
and U13547 (N_13547,N_13289,N_13381);
nand U13548 (N_13548,N_13220,N_13228);
or U13549 (N_13549,N_13285,N_13218);
or U13550 (N_13550,N_13350,N_13240);
and U13551 (N_13551,N_13288,N_13328);
nor U13552 (N_13552,N_13246,N_13372);
nand U13553 (N_13553,N_13385,N_13315);
nand U13554 (N_13554,N_13234,N_13201);
or U13555 (N_13555,N_13367,N_13296);
xor U13556 (N_13556,N_13383,N_13361);
nand U13557 (N_13557,N_13295,N_13374);
nand U13558 (N_13558,N_13356,N_13354);
xnor U13559 (N_13559,N_13201,N_13332);
and U13560 (N_13560,N_13233,N_13324);
xor U13561 (N_13561,N_13340,N_13358);
nor U13562 (N_13562,N_13273,N_13313);
or U13563 (N_13563,N_13347,N_13358);
xor U13564 (N_13564,N_13301,N_13333);
or U13565 (N_13565,N_13294,N_13260);
or U13566 (N_13566,N_13244,N_13376);
nand U13567 (N_13567,N_13315,N_13369);
nand U13568 (N_13568,N_13358,N_13333);
nand U13569 (N_13569,N_13288,N_13391);
and U13570 (N_13570,N_13369,N_13205);
xnor U13571 (N_13571,N_13293,N_13224);
nor U13572 (N_13572,N_13209,N_13329);
or U13573 (N_13573,N_13390,N_13218);
or U13574 (N_13574,N_13242,N_13308);
xor U13575 (N_13575,N_13248,N_13388);
or U13576 (N_13576,N_13300,N_13251);
and U13577 (N_13577,N_13262,N_13390);
nor U13578 (N_13578,N_13375,N_13253);
or U13579 (N_13579,N_13370,N_13288);
and U13580 (N_13580,N_13258,N_13251);
or U13581 (N_13581,N_13226,N_13310);
and U13582 (N_13582,N_13262,N_13394);
xor U13583 (N_13583,N_13307,N_13253);
xor U13584 (N_13584,N_13256,N_13352);
xnor U13585 (N_13585,N_13344,N_13327);
nor U13586 (N_13586,N_13264,N_13272);
and U13587 (N_13587,N_13237,N_13383);
nor U13588 (N_13588,N_13226,N_13319);
and U13589 (N_13589,N_13396,N_13348);
nor U13590 (N_13590,N_13253,N_13342);
nand U13591 (N_13591,N_13202,N_13349);
nand U13592 (N_13592,N_13216,N_13213);
nor U13593 (N_13593,N_13273,N_13382);
nand U13594 (N_13594,N_13202,N_13311);
and U13595 (N_13595,N_13381,N_13269);
or U13596 (N_13596,N_13349,N_13216);
nand U13597 (N_13597,N_13205,N_13376);
and U13598 (N_13598,N_13241,N_13373);
and U13599 (N_13599,N_13233,N_13265);
nor U13600 (N_13600,N_13538,N_13578);
xor U13601 (N_13601,N_13424,N_13589);
and U13602 (N_13602,N_13440,N_13497);
nand U13603 (N_13603,N_13452,N_13571);
nand U13604 (N_13604,N_13433,N_13413);
xor U13605 (N_13605,N_13597,N_13556);
nor U13606 (N_13606,N_13435,N_13521);
nor U13607 (N_13607,N_13446,N_13490);
nor U13608 (N_13608,N_13463,N_13590);
nor U13609 (N_13609,N_13476,N_13515);
nor U13610 (N_13610,N_13557,N_13544);
nor U13611 (N_13611,N_13583,N_13401);
xnor U13612 (N_13612,N_13430,N_13454);
or U13613 (N_13613,N_13466,N_13488);
and U13614 (N_13614,N_13530,N_13576);
and U13615 (N_13615,N_13457,N_13568);
xnor U13616 (N_13616,N_13451,N_13514);
nor U13617 (N_13617,N_13465,N_13573);
or U13618 (N_13618,N_13560,N_13529);
xor U13619 (N_13619,N_13562,N_13595);
xnor U13620 (N_13620,N_13569,N_13419);
xor U13621 (N_13621,N_13537,N_13484);
nand U13622 (N_13622,N_13408,N_13426);
xor U13623 (N_13623,N_13472,N_13406);
xnor U13624 (N_13624,N_13444,N_13525);
and U13625 (N_13625,N_13539,N_13460);
xnor U13626 (N_13626,N_13405,N_13471);
or U13627 (N_13627,N_13501,N_13438);
xnor U13628 (N_13628,N_13431,N_13459);
or U13629 (N_13629,N_13499,N_13527);
and U13630 (N_13630,N_13554,N_13445);
and U13631 (N_13631,N_13513,N_13547);
nand U13632 (N_13632,N_13494,N_13481);
xor U13633 (N_13633,N_13421,N_13464);
and U13634 (N_13634,N_13453,N_13404);
nor U13635 (N_13635,N_13486,N_13599);
nand U13636 (N_13636,N_13526,N_13516);
xnor U13637 (N_13637,N_13442,N_13534);
xor U13638 (N_13638,N_13553,N_13473);
xor U13639 (N_13639,N_13586,N_13427);
and U13640 (N_13640,N_13585,N_13448);
xnor U13641 (N_13641,N_13443,N_13482);
or U13642 (N_13642,N_13417,N_13407);
nand U13643 (N_13643,N_13412,N_13447);
xnor U13644 (N_13644,N_13559,N_13508);
or U13645 (N_13645,N_13478,N_13594);
nand U13646 (N_13646,N_13450,N_13410);
xor U13647 (N_13647,N_13546,N_13572);
xor U13648 (N_13648,N_13565,N_13498);
xor U13649 (N_13649,N_13532,N_13528);
xnor U13650 (N_13650,N_13496,N_13422);
or U13651 (N_13651,N_13485,N_13536);
nand U13652 (N_13652,N_13533,N_13428);
nor U13653 (N_13653,N_13558,N_13458);
nand U13654 (N_13654,N_13434,N_13581);
or U13655 (N_13655,N_13507,N_13423);
nor U13656 (N_13656,N_13477,N_13480);
nor U13657 (N_13657,N_13475,N_13495);
nand U13658 (N_13658,N_13524,N_13439);
xnor U13659 (N_13659,N_13470,N_13489);
nand U13660 (N_13660,N_13577,N_13414);
nand U13661 (N_13661,N_13567,N_13555);
or U13662 (N_13662,N_13461,N_13520);
or U13663 (N_13663,N_13542,N_13400);
xor U13664 (N_13664,N_13543,N_13449);
nand U13665 (N_13665,N_13598,N_13551);
xor U13666 (N_13666,N_13416,N_13509);
nand U13667 (N_13667,N_13517,N_13580);
and U13668 (N_13668,N_13469,N_13462);
nor U13669 (N_13669,N_13540,N_13411);
or U13670 (N_13670,N_13519,N_13587);
and U13671 (N_13671,N_13561,N_13593);
nor U13672 (N_13672,N_13548,N_13596);
nor U13673 (N_13673,N_13418,N_13491);
nand U13674 (N_13674,N_13582,N_13552);
xor U13675 (N_13675,N_13493,N_13487);
and U13676 (N_13676,N_13584,N_13500);
or U13677 (N_13677,N_13467,N_13510);
nor U13678 (N_13678,N_13506,N_13549);
nor U13679 (N_13679,N_13420,N_13575);
nand U13680 (N_13680,N_13402,N_13574);
nand U13681 (N_13681,N_13436,N_13564);
and U13682 (N_13682,N_13409,N_13492);
nor U13683 (N_13683,N_13579,N_13455);
nor U13684 (N_13684,N_13403,N_13550);
and U13685 (N_13685,N_13502,N_13437);
nor U13686 (N_13686,N_13563,N_13588);
nor U13687 (N_13687,N_13425,N_13591);
nand U13688 (N_13688,N_13518,N_13523);
xnor U13689 (N_13689,N_13503,N_13535);
and U13690 (N_13690,N_13441,N_13483);
nor U13691 (N_13691,N_13468,N_13522);
and U13692 (N_13692,N_13545,N_13474);
xor U13693 (N_13693,N_13432,N_13531);
or U13694 (N_13694,N_13541,N_13456);
nand U13695 (N_13695,N_13511,N_13566);
nand U13696 (N_13696,N_13504,N_13429);
nor U13697 (N_13697,N_13512,N_13570);
nor U13698 (N_13698,N_13479,N_13505);
and U13699 (N_13699,N_13415,N_13592);
or U13700 (N_13700,N_13568,N_13405);
nand U13701 (N_13701,N_13400,N_13417);
or U13702 (N_13702,N_13498,N_13541);
and U13703 (N_13703,N_13406,N_13420);
nand U13704 (N_13704,N_13567,N_13575);
nor U13705 (N_13705,N_13471,N_13577);
xnor U13706 (N_13706,N_13557,N_13483);
or U13707 (N_13707,N_13592,N_13586);
nor U13708 (N_13708,N_13518,N_13461);
nand U13709 (N_13709,N_13452,N_13503);
nand U13710 (N_13710,N_13576,N_13562);
xor U13711 (N_13711,N_13492,N_13581);
nor U13712 (N_13712,N_13517,N_13514);
and U13713 (N_13713,N_13553,N_13561);
or U13714 (N_13714,N_13488,N_13424);
xor U13715 (N_13715,N_13450,N_13540);
nand U13716 (N_13716,N_13432,N_13543);
and U13717 (N_13717,N_13546,N_13581);
nor U13718 (N_13718,N_13519,N_13528);
nand U13719 (N_13719,N_13560,N_13519);
and U13720 (N_13720,N_13402,N_13542);
or U13721 (N_13721,N_13483,N_13417);
and U13722 (N_13722,N_13548,N_13553);
xnor U13723 (N_13723,N_13522,N_13441);
nor U13724 (N_13724,N_13403,N_13522);
or U13725 (N_13725,N_13456,N_13403);
and U13726 (N_13726,N_13595,N_13421);
xor U13727 (N_13727,N_13535,N_13441);
or U13728 (N_13728,N_13565,N_13425);
nor U13729 (N_13729,N_13449,N_13504);
nor U13730 (N_13730,N_13464,N_13439);
or U13731 (N_13731,N_13550,N_13510);
and U13732 (N_13732,N_13496,N_13439);
and U13733 (N_13733,N_13455,N_13578);
nand U13734 (N_13734,N_13568,N_13514);
and U13735 (N_13735,N_13426,N_13547);
xor U13736 (N_13736,N_13525,N_13559);
nand U13737 (N_13737,N_13546,N_13428);
nor U13738 (N_13738,N_13485,N_13593);
xor U13739 (N_13739,N_13485,N_13564);
nand U13740 (N_13740,N_13546,N_13583);
nand U13741 (N_13741,N_13432,N_13476);
or U13742 (N_13742,N_13596,N_13568);
nand U13743 (N_13743,N_13465,N_13410);
nor U13744 (N_13744,N_13409,N_13566);
nor U13745 (N_13745,N_13510,N_13500);
or U13746 (N_13746,N_13467,N_13591);
nand U13747 (N_13747,N_13552,N_13403);
and U13748 (N_13748,N_13521,N_13470);
or U13749 (N_13749,N_13427,N_13409);
nor U13750 (N_13750,N_13566,N_13435);
xnor U13751 (N_13751,N_13526,N_13593);
and U13752 (N_13752,N_13474,N_13528);
nand U13753 (N_13753,N_13582,N_13450);
nor U13754 (N_13754,N_13496,N_13462);
nor U13755 (N_13755,N_13534,N_13490);
nor U13756 (N_13756,N_13557,N_13440);
or U13757 (N_13757,N_13407,N_13552);
and U13758 (N_13758,N_13538,N_13436);
xnor U13759 (N_13759,N_13438,N_13547);
nor U13760 (N_13760,N_13423,N_13561);
nor U13761 (N_13761,N_13418,N_13561);
or U13762 (N_13762,N_13483,N_13425);
or U13763 (N_13763,N_13525,N_13413);
or U13764 (N_13764,N_13400,N_13572);
nand U13765 (N_13765,N_13546,N_13409);
and U13766 (N_13766,N_13549,N_13491);
xor U13767 (N_13767,N_13475,N_13576);
and U13768 (N_13768,N_13567,N_13492);
nand U13769 (N_13769,N_13483,N_13433);
and U13770 (N_13770,N_13460,N_13571);
nand U13771 (N_13771,N_13509,N_13540);
xnor U13772 (N_13772,N_13586,N_13501);
nand U13773 (N_13773,N_13426,N_13463);
nor U13774 (N_13774,N_13535,N_13596);
and U13775 (N_13775,N_13436,N_13595);
nand U13776 (N_13776,N_13412,N_13567);
xnor U13777 (N_13777,N_13580,N_13508);
xnor U13778 (N_13778,N_13537,N_13527);
or U13779 (N_13779,N_13429,N_13410);
or U13780 (N_13780,N_13535,N_13417);
nand U13781 (N_13781,N_13430,N_13511);
nand U13782 (N_13782,N_13464,N_13489);
or U13783 (N_13783,N_13437,N_13410);
nor U13784 (N_13784,N_13424,N_13419);
or U13785 (N_13785,N_13552,N_13579);
or U13786 (N_13786,N_13594,N_13523);
nand U13787 (N_13787,N_13504,N_13513);
xor U13788 (N_13788,N_13496,N_13465);
nor U13789 (N_13789,N_13513,N_13500);
and U13790 (N_13790,N_13586,N_13539);
xor U13791 (N_13791,N_13514,N_13537);
xnor U13792 (N_13792,N_13536,N_13554);
and U13793 (N_13793,N_13550,N_13579);
and U13794 (N_13794,N_13497,N_13498);
xnor U13795 (N_13795,N_13480,N_13437);
nand U13796 (N_13796,N_13488,N_13414);
and U13797 (N_13797,N_13563,N_13435);
xnor U13798 (N_13798,N_13544,N_13571);
or U13799 (N_13799,N_13575,N_13588);
or U13800 (N_13800,N_13642,N_13735);
or U13801 (N_13801,N_13720,N_13668);
or U13802 (N_13802,N_13654,N_13704);
nand U13803 (N_13803,N_13669,N_13758);
nor U13804 (N_13804,N_13759,N_13756);
or U13805 (N_13805,N_13609,N_13635);
nor U13806 (N_13806,N_13763,N_13714);
nor U13807 (N_13807,N_13626,N_13796);
xnor U13808 (N_13808,N_13616,N_13643);
or U13809 (N_13809,N_13760,N_13713);
xor U13810 (N_13810,N_13795,N_13630);
nor U13811 (N_13811,N_13783,N_13683);
xnor U13812 (N_13812,N_13649,N_13749);
and U13813 (N_13813,N_13723,N_13774);
and U13814 (N_13814,N_13753,N_13679);
or U13815 (N_13815,N_13757,N_13606);
and U13816 (N_13816,N_13687,N_13699);
xor U13817 (N_13817,N_13681,N_13694);
nand U13818 (N_13818,N_13733,N_13743);
nor U13819 (N_13819,N_13770,N_13786);
nand U13820 (N_13820,N_13767,N_13631);
nand U13821 (N_13821,N_13691,N_13641);
and U13822 (N_13822,N_13634,N_13744);
or U13823 (N_13823,N_13678,N_13670);
nor U13824 (N_13824,N_13612,N_13793);
xor U13825 (N_13825,N_13705,N_13639);
nand U13826 (N_13826,N_13690,N_13784);
or U13827 (N_13827,N_13703,N_13721);
nor U13828 (N_13828,N_13648,N_13667);
xnor U13829 (N_13829,N_13725,N_13709);
nor U13830 (N_13830,N_13764,N_13628);
xnor U13831 (N_13831,N_13617,N_13696);
or U13832 (N_13832,N_13688,N_13740);
nor U13833 (N_13833,N_13755,N_13772);
xnor U13834 (N_13834,N_13621,N_13775);
and U13835 (N_13835,N_13666,N_13741);
nand U13836 (N_13836,N_13779,N_13600);
nand U13837 (N_13837,N_13636,N_13745);
xnor U13838 (N_13838,N_13640,N_13665);
or U13839 (N_13839,N_13731,N_13653);
or U13840 (N_13840,N_13708,N_13663);
nand U13841 (N_13841,N_13710,N_13718);
and U13842 (N_13842,N_13661,N_13650);
or U13843 (N_13843,N_13790,N_13660);
and U13844 (N_13844,N_13676,N_13798);
or U13845 (N_13845,N_13697,N_13788);
nand U13846 (N_13846,N_13615,N_13673);
xnor U13847 (N_13847,N_13706,N_13777);
nand U13848 (N_13848,N_13656,N_13602);
nor U13849 (N_13849,N_13604,N_13719);
xnor U13850 (N_13850,N_13647,N_13768);
or U13851 (N_13851,N_13657,N_13624);
nand U13852 (N_13852,N_13742,N_13785);
nand U13853 (N_13853,N_13680,N_13682);
xnor U13854 (N_13854,N_13613,N_13717);
and U13855 (N_13855,N_13782,N_13750);
nor U13856 (N_13856,N_13765,N_13662);
nor U13857 (N_13857,N_13693,N_13603);
nor U13858 (N_13858,N_13792,N_13728);
or U13859 (N_13859,N_13701,N_13736);
xnor U13860 (N_13860,N_13689,N_13727);
xnor U13861 (N_13861,N_13737,N_13766);
nand U13862 (N_13862,N_13730,N_13729);
nor U13863 (N_13863,N_13778,N_13776);
xnor U13864 (N_13864,N_13645,N_13791);
nand U13865 (N_13865,N_13752,N_13762);
xnor U13866 (N_13866,N_13726,N_13625);
xor U13867 (N_13867,N_13716,N_13623);
xor U13868 (N_13868,N_13695,N_13747);
or U13869 (N_13869,N_13761,N_13620);
nand U13870 (N_13870,N_13618,N_13651);
xnor U13871 (N_13871,N_13685,N_13732);
and U13872 (N_13872,N_13684,N_13799);
xnor U13873 (N_13873,N_13655,N_13698);
or U13874 (N_13874,N_13658,N_13671);
and U13875 (N_13875,N_13644,N_13734);
and U13876 (N_13876,N_13700,N_13769);
or U13877 (N_13877,N_13773,N_13619);
or U13878 (N_13878,N_13633,N_13611);
xor U13879 (N_13879,N_13797,N_13607);
nand U13880 (N_13880,N_13702,N_13739);
and U13881 (N_13881,N_13692,N_13610);
and U13882 (N_13882,N_13754,N_13605);
nor U13883 (N_13883,N_13686,N_13787);
nand U13884 (N_13884,N_13601,N_13707);
and U13885 (N_13885,N_13622,N_13632);
or U13886 (N_13886,N_13677,N_13652);
xor U13887 (N_13887,N_13675,N_13629);
xnor U13888 (N_13888,N_13748,N_13672);
xor U13889 (N_13889,N_13715,N_13724);
and U13890 (N_13890,N_13746,N_13722);
xor U13891 (N_13891,N_13771,N_13780);
and U13892 (N_13892,N_13646,N_13637);
or U13893 (N_13893,N_13711,N_13614);
nand U13894 (N_13894,N_13712,N_13738);
nor U13895 (N_13895,N_13751,N_13794);
nand U13896 (N_13896,N_13789,N_13627);
nor U13897 (N_13897,N_13638,N_13664);
xor U13898 (N_13898,N_13674,N_13608);
nand U13899 (N_13899,N_13659,N_13781);
nand U13900 (N_13900,N_13785,N_13715);
or U13901 (N_13901,N_13694,N_13604);
nor U13902 (N_13902,N_13730,N_13798);
nand U13903 (N_13903,N_13721,N_13633);
xor U13904 (N_13904,N_13698,N_13779);
nand U13905 (N_13905,N_13771,N_13758);
xor U13906 (N_13906,N_13775,N_13767);
nor U13907 (N_13907,N_13750,N_13703);
xnor U13908 (N_13908,N_13777,N_13687);
or U13909 (N_13909,N_13765,N_13723);
and U13910 (N_13910,N_13712,N_13739);
or U13911 (N_13911,N_13781,N_13754);
or U13912 (N_13912,N_13647,N_13791);
or U13913 (N_13913,N_13784,N_13754);
and U13914 (N_13914,N_13702,N_13687);
and U13915 (N_13915,N_13785,N_13706);
and U13916 (N_13916,N_13638,N_13631);
nor U13917 (N_13917,N_13719,N_13736);
nand U13918 (N_13918,N_13773,N_13655);
nand U13919 (N_13919,N_13601,N_13702);
xnor U13920 (N_13920,N_13759,N_13603);
nor U13921 (N_13921,N_13746,N_13774);
and U13922 (N_13922,N_13707,N_13623);
nor U13923 (N_13923,N_13688,N_13730);
and U13924 (N_13924,N_13697,N_13628);
nand U13925 (N_13925,N_13638,N_13776);
nor U13926 (N_13926,N_13747,N_13775);
xnor U13927 (N_13927,N_13649,N_13753);
nand U13928 (N_13928,N_13642,N_13778);
nand U13929 (N_13929,N_13760,N_13718);
or U13930 (N_13930,N_13648,N_13741);
and U13931 (N_13931,N_13680,N_13739);
and U13932 (N_13932,N_13600,N_13702);
nand U13933 (N_13933,N_13698,N_13675);
and U13934 (N_13934,N_13696,N_13793);
or U13935 (N_13935,N_13641,N_13672);
or U13936 (N_13936,N_13717,N_13718);
nand U13937 (N_13937,N_13738,N_13729);
or U13938 (N_13938,N_13601,N_13694);
nand U13939 (N_13939,N_13756,N_13703);
and U13940 (N_13940,N_13750,N_13689);
or U13941 (N_13941,N_13747,N_13739);
or U13942 (N_13942,N_13707,N_13787);
xnor U13943 (N_13943,N_13756,N_13683);
nor U13944 (N_13944,N_13730,N_13624);
nor U13945 (N_13945,N_13752,N_13626);
xor U13946 (N_13946,N_13725,N_13643);
nand U13947 (N_13947,N_13710,N_13760);
nor U13948 (N_13948,N_13615,N_13657);
xnor U13949 (N_13949,N_13768,N_13635);
and U13950 (N_13950,N_13635,N_13692);
nand U13951 (N_13951,N_13778,N_13616);
or U13952 (N_13952,N_13763,N_13771);
and U13953 (N_13953,N_13644,N_13784);
nand U13954 (N_13954,N_13664,N_13799);
and U13955 (N_13955,N_13778,N_13758);
nor U13956 (N_13956,N_13633,N_13618);
nand U13957 (N_13957,N_13725,N_13733);
xnor U13958 (N_13958,N_13723,N_13750);
nor U13959 (N_13959,N_13733,N_13799);
and U13960 (N_13960,N_13784,N_13692);
nor U13961 (N_13961,N_13681,N_13617);
xnor U13962 (N_13962,N_13739,N_13726);
and U13963 (N_13963,N_13785,N_13795);
and U13964 (N_13964,N_13647,N_13698);
or U13965 (N_13965,N_13669,N_13604);
or U13966 (N_13966,N_13609,N_13713);
and U13967 (N_13967,N_13619,N_13746);
nor U13968 (N_13968,N_13647,N_13765);
and U13969 (N_13969,N_13646,N_13689);
or U13970 (N_13970,N_13676,N_13649);
nand U13971 (N_13971,N_13782,N_13758);
nor U13972 (N_13972,N_13624,N_13711);
xor U13973 (N_13973,N_13720,N_13795);
xor U13974 (N_13974,N_13680,N_13669);
xor U13975 (N_13975,N_13748,N_13738);
nor U13976 (N_13976,N_13626,N_13754);
nor U13977 (N_13977,N_13657,N_13648);
xnor U13978 (N_13978,N_13646,N_13682);
and U13979 (N_13979,N_13670,N_13766);
nand U13980 (N_13980,N_13676,N_13659);
or U13981 (N_13981,N_13692,N_13620);
nand U13982 (N_13982,N_13664,N_13770);
xor U13983 (N_13983,N_13718,N_13627);
nand U13984 (N_13984,N_13756,N_13735);
and U13985 (N_13985,N_13759,N_13783);
xor U13986 (N_13986,N_13795,N_13756);
xor U13987 (N_13987,N_13616,N_13615);
or U13988 (N_13988,N_13702,N_13671);
and U13989 (N_13989,N_13737,N_13616);
or U13990 (N_13990,N_13647,N_13742);
nand U13991 (N_13991,N_13706,N_13789);
and U13992 (N_13992,N_13666,N_13677);
nand U13993 (N_13993,N_13669,N_13797);
nor U13994 (N_13994,N_13692,N_13751);
xor U13995 (N_13995,N_13675,N_13735);
or U13996 (N_13996,N_13715,N_13729);
and U13997 (N_13997,N_13647,N_13651);
nand U13998 (N_13998,N_13793,N_13732);
xnor U13999 (N_13999,N_13792,N_13652);
xor U14000 (N_14000,N_13901,N_13865);
or U14001 (N_14001,N_13899,N_13872);
xor U14002 (N_14002,N_13853,N_13934);
nor U14003 (N_14003,N_13852,N_13832);
xor U14004 (N_14004,N_13906,N_13992);
or U14005 (N_14005,N_13837,N_13953);
xor U14006 (N_14006,N_13845,N_13816);
and U14007 (N_14007,N_13931,N_13846);
nor U14008 (N_14008,N_13891,N_13983);
nor U14009 (N_14009,N_13818,N_13978);
and U14010 (N_14010,N_13909,N_13850);
xor U14011 (N_14011,N_13890,N_13841);
nand U14012 (N_14012,N_13958,N_13952);
nor U14013 (N_14013,N_13888,N_13903);
xor U14014 (N_14014,N_13977,N_13885);
nand U14015 (N_14015,N_13877,N_13919);
xnor U14016 (N_14016,N_13827,N_13811);
or U14017 (N_14017,N_13976,N_13967);
and U14018 (N_14018,N_13951,N_13927);
or U14019 (N_14019,N_13905,N_13942);
xnor U14020 (N_14020,N_13855,N_13889);
nor U14021 (N_14021,N_13883,N_13802);
nor U14022 (N_14022,N_13862,N_13940);
and U14023 (N_14023,N_13821,N_13985);
nand U14024 (N_14024,N_13928,N_13870);
or U14025 (N_14025,N_13950,N_13873);
xor U14026 (N_14026,N_13932,N_13881);
nor U14027 (N_14027,N_13922,N_13972);
or U14028 (N_14028,N_13829,N_13941);
nand U14029 (N_14029,N_13908,N_13948);
and U14030 (N_14030,N_13868,N_13887);
xor U14031 (N_14031,N_13860,N_13939);
xor U14032 (N_14032,N_13954,N_13966);
or U14033 (N_14033,N_13863,N_13858);
xnor U14034 (N_14034,N_13831,N_13902);
or U14035 (N_14035,N_13986,N_13947);
nand U14036 (N_14036,N_13896,N_13938);
xor U14037 (N_14037,N_13982,N_13804);
xor U14038 (N_14038,N_13848,N_13898);
xnor U14039 (N_14039,N_13875,N_13971);
nand U14040 (N_14040,N_13842,N_13955);
nor U14041 (N_14041,N_13936,N_13808);
or U14042 (N_14042,N_13960,N_13973);
or U14043 (N_14043,N_13819,N_13970);
nand U14044 (N_14044,N_13915,N_13921);
xor U14045 (N_14045,N_13805,N_13878);
and U14046 (N_14046,N_13897,N_13913);
nor U14047 (N_14047,N_13814,N_13993);
nor U14048 (N_14048,N_13937,N_13933);
nor U14049 (N_14049,N_13984,N_13824);
and U14050 (N_14050,N_13861,N_13895);
nand U14051 (N_14051,N_13806,N_13989);
nor U14052 (N_14052,N_13810,N_13893);
or U14053 (N_14053,N_13800,N_13988);
nand U14054 (N_14054,N_13946,N_13994);
and U14055 (N_14055,N_13964,N_13990);
nand U14056 (N_14056,N_13894,N_13975);
nand U14057 (N_14057,N_13876,N_13840);
nand U14058 (N_14058,N_13916,N_13833);
or U14059 (N_14059,N_13929,N_13866);
xnor U14060 (N_14060,N_13981,N_13980);
xnor U14061 (N_14061,N_13874,N_13820);
nand U14062 (N_14062,N_13839,N_13854);
or U14063 (N_14063,N_13812,N_13843);
or U14064 (N_14064,N_13807,N_13923);
xor U14065 (N_14065,N_13944,N_13886);
or U14066 (N_14066,N_13892,N_13911);
nand U14067 (N_14067,N_13817,N_13907);
xor U14068 (N_14068,N_13996,N_13864);
xnor U14069 (N_14069,N_13834,N_13949);
and U14070 (N_14070,N_13835,N_13859);
nand U14071 (N_14071,N_13825,N_13847);
or U14072 (N_14072,N_13813,N_13961);
nand U14073 (N_14073,N_13965,N_13904);
nand U14074 (N_14074,N_13822,N_13918);
xnor U14075 (N_14075,N_13849,N_13945);
nor U14076 (N_14076,N_13880,N_13803);
xor U14077 (N_14077,N_13856,N_13914);
nor U14078 (N_14078,N_13884,N_13828);
nand U14079 (N_14079,N_13995,N_13974);
and U14080 (N_14080,N_13838,N_13969);
and U14081 (N_14081,N_13801,N_13963);
nor U14082 (N_14082,N_13943,N_13815);
nor U14083 (N_14083,N_13924,N_13869);
nor U14084 (N_14084,N_13935,N_13823);
nand U14085 (N_14085,N_13987,N_13959);
or U14086 (N_14086,N_13857,N_13809);
nor U14087 (N_14087,N_13998,N_13991);
xnor U14088 (N_14088,N_13879,N_13920);
or U14089 (N_14089,N_13912,N_13956);
xor U14090 (N_14090,N_13851,N_13844);
or U14091 (N_14091,N_13910,N_13968);
and U14092 (N_14092,N_13882,N_13997);
nor U14093 (N_14093,N_13930,N_13867);
and U14094 (N_14094,N_13830,N_13900);
nand U14095 (N_14095,N_13871,N_13926);
and U14096 (N_14096,N_13957,N_13836);
nor U14097 (N_14097,N_13925,N_13979);
and U14098 (N_14098,N_13962,N_13999);
and U14099 (N_14099,N_13917,N_13826);
nor U14100 (N_14100,N_13970,N_13960);
xnor U14101 (N_14101,N_13950,N_13937);
nand U14102 (N_14102,N_13965,N_13860);
and U14103 (N_14103,N_13863,N_13880);
nand U14104 (N_14104,N_13874,N_13818);
and U14105 (N_14105,N_13829,N_13986);
and U14106 (N_14106,N_13848,N_13861);
nor U14107 (N_14107,N_13946,N_13934);
xnor U14108 (N_14108,N_13983,N_13927);
or U14109 (N_14109,N_13864,N_13902);
nand U14110 (N_14110,N_13948,N_13862);
xnor U14111 (N_14111,N_13981,N_13853);
nand U14112 (N_14112,N_13893,N_13920);
nand U14113 (N_14113,N_13845,N_13916);
nor U14114 (N_14114,N_13968,N_13850);
nor U14115 (N_14115,N_13979,N_13848);
xor U14116 (N_14116,N_13868,N_13909);
xnor U14117 (N_14117,N_13865,N_13832);
or U14118 (N_14118,N_13906,N_13893);
nor U14119 (N_14119,N_13869,N_13841);
and U14120 (N_14120,N_13956,N_13960);
nor U14121 (N_14121,N_13998,N_13906);
and U14122 (N_14122,N_13871,N_13979);
nand U14123 (N_14123,N_13961,N_13884);
or U14124 (N_14124,N_13943,N_13930);
and U14125 (N_14125,N_13853,N_13849);
or U14126 (N_14126,N_13979,N_13913);
nand U14127 (N_14127,N_13895,N_13817);
nor U14128 (N_14128,N_13970,N_13813);
xnor U14129 (N_14129,N_13809,N_13994);
or U14130 (N_14130,N_13909,N_13966);
xor U14131 (N_14131,N_13905,N_13936);
and U14132 (N_14132,N_13840,N_13839);
nand U14133 (N_14133,N_13833,N_13858);
or U14134 (N_14134,N_13876,N_13828);
nand U14135 (N_14135,N_13876,N_13947);
xnor U14136 (N_14136,N_13913,N_13867);
or U14137 (N_14137,N_13884,N_13980);
and U14138 (N_14138,N_13901,N_13987);
nand U14139 (N_14139,N_13969,N_13987);
and U14140 (N_14140,N_13964,N_13996);
xnor U14141 (N_14141,N_13888,N_13830);
nand U14142 (N_14142,N_13925,N_13852);
and U14143 (N_14143,N_13870,N_13920);
and U14144 (N_14144,N_13887,N_13905);
or U14145 (N_14145,N_13821,N_13833);
xor U14146 (N_14146,N_13938,N_13966);
nand U14147 (N_14147,N_13866,N_13846);
nor U14148 (N_14148,N_13885,N_13874);
or U14149 (N_14149,N_13995,N_13947);
nand U14150 (N_14150,N_13981,N_13907);
and U14151 (N_14151,N_13998,N_13861);
and U14152 (N_14152,N_13985,N_13978);
or U14153 (N_14153,N_13995,N_13903);
and U14154 (N_14154,N_13938,N_13881);
nand U14155 (N_14155,N_13972,N_13808);
and U14156 (N_14156,N_13880,N_13971);
or U14157 (N_14157,N_13986,N_13845);
nand U14158 (N_14158,N_13824,N_13906);
or U14159 (N_14159,N_13834,N_13922);
nor U14160 (N_14160,N_13994,N_13905);
nand U14161 (N_14161,N_13911,N_13880);
xnor U14162 (N_14162,N_13952,N_13835);
xor U14163 (N_14163,N_13865,N_13984);
and U14164 (N_14164,N_13828,N_13867);
and U14165 (N_14165,N_13818,N_13883);
xor U14166 (N_14166,N_13930,N_13885);
nor U14167 (N_14167,N_13978,N_13871);
or U14168 (N_14168,N_13932,N_13906);
nand U14169 (N_14169,N_13881,N_13866);
or U14170 (N_14170,N_13888,N_13918);
nor U14171 (N_14171,N_13833,N_13826);
xnor U14172 (N_14172,N_13923,N_13990);
or U14173 (N_14173,N_13918,N_13980);
nand U14174 (N_14174,N_13884,N_13908);
and U14175 (N_14175,N_13982,N_13816);
nand U14176 (N_14176,N_13820,N_13814);
or U14177 (N_14177,N_13953,N_13860);
and U14178 (N_14178,N_13832,N_13895);
nand U14179 (N_14179,N_13945,N_13868);
or U14180 (N_14180,N_13979,N_13928);
nor U14181 (N_14181,N_13818,N_13852);
nor U14182 (N_14182,N_13841,N_13919);
and U14183 (N_14183,N_13844,N_13983);
and U14184 (N_14184,N_13944,N_13913);
and U14185 (N_14185,N_13844,N_13901);
nor U14186 (N_14186,N_13944,N_13805);
or U14187 (N_14187,N_13815,N_13962);
or U14188 (N_14188,N_13890,N_13855);
and U14189 (N_14189,N_13831,N_13870);
xor U14190 (N_14190,N_13929,N_13868);
nor U14191 (N_14191,N_13806,N_13816);
nand U14192 (N_14192,N_13922,N_13980);
and U14193 (N_14193,N_13874,N_13894);
nand U14194 (N_14194,N_13871,N_13847);
or U14195 (N_14195,N_13932,N_13851);
or U14196 (N_14196,N_13892,N_13820);
and U14197 (N_14197,N_13954,N_13844);
nand U14198 (N_14198,N_13877,N_13845);
and U14199 (N_14199,N_13951,N_13976);
nand U14200 (N_14200,N_14047,N_14014);
nor U14201 (N_14201,N_14072,N_14076);
nor U14202 (N_14202,N_14163,N_14022);
nand U14203 (N_14203,N_14121,N_14146);
xor U14204 (N_14204,N_14024,N_14050);
nor U14205 (N_14205,N_14130,N_14101);
nor U14206 (N_14206,N_14073,N_14150);
nor U14207 (N_14207,N_14032,N_14185);
and U14208 (N_14208,N_14085,N_14173);
nor U14209 (N_14209,N_14025,N_14001);
and U14210 (N_14210,N_14088,N_14046);
and U14211 (N_14211,N_14000,N_14183);
or U14212 (N_14212,N_14051,N_14133);
nor U14213 (N_14213,N_14069,N_14129);
nor U14214 (N_14214,N_14011,N_14153);
nor U14215 (N_14215,N_14191,N_14174);
nand U14216 (N_14216,N_14197,N_14168);
nor U14217 (N_14217,N_14010,N_14106);
or U14218 (N_14218,N_14145,N_14067);
nor U14219 (N_14219,N_14104,N_14002);
xnor U14220 (N_14220,N_14020,N_14107);
and U14221 (N_14221,N_14157,N_14038);
nor U14222 (N_14222,N_14048,N_14099);
nand U14223 (N_14223,N_14003,N_14086);
or U14224 (N_14224,N_14187,N_14040);
nor U14225 (N_14225,N_14118,N_14125);
and U14226 (N_14226,N_14171,N_14023);
or U14227 (N_14227,N_14136,N_14122);
nor U14228 (N_14228,N_14128,N_14119);
nor U14229 (N_14229,N_14194,N_14195);
xor U14230 (N_14230,N_14190,N_14117);
and U14231 (N_14231,N_14184,N_14031);
or U14232 (N_14232,N_14156,N_14026);
and U14233 (N_14233,N_14054,N_14193);
xor U14234 (N_14234,N_14021,N_14116);
nor U14235 (N_14235,N_14165,N_14009);
and U14236 (N_14236,N_14177,N_14199);
nand U14237 (N_14237,N_14037,N_14029);
nand U14238 (N_14238,N_14115,N_14036);
nand U14239 (N_14239,N_14162,N_14134);
xor U14240 (N_14240,N_14139,N_14148);
nor U14241 (N_14241,N_14112,N_14126);
or U14242 (N_14242,N_14064,N_14071);
or U14243 (N_14243,N_14172,N_14114);
nand U14244 (N_14244,N_14039,N_14044);
or U14245 (N_14245,N_14030,N_14013);
nand U14246 (N_14246,N_14094,N_14063);
nand U14247 (N_14247,N_14075,N_14066);
or U14248 (N_14248,N_14095,N_14097);
nor U14249 (N_14249,N_14070,N_14192);
nand U14250 (N_14250,N_14080,N_14147);
and U14251 (N_14251,N_14181,N_14074);
xor U14252 (N_14252,N_14100,N_14078);
nor U14253 (N_14253,N_14149,N_14028);
nor U14254 (N_14254,N_14062,N_14176);
nor U14255 (N_14255,N_14186,N_14012);
xnor U14256 (N_14256,N_14052,N_14182);
nand U14257 (N_14257,N_14167,N_14019);
nor U14258 (N_14258,N_14016,N_14077);
nor U14259 (N_14259,N_14120,N_14098);
and U14260 (N_14260,N_14060,N_14053);
or U14261 (N_14261,N_14082,N_14198);
or U14262 (N_14262,N_14005,N_14161);
nor U14263 (N_14263,N_14041,N_14035);
or U14264 (N_14264,N_14049,N_14154);
or U14265 (N_14265,N_14151,N_14108);
xor U14266 (N_14266,N_14089,N_14084);
nand U14267 (N_14267,N_14008,N_14152);
or U14268 (N_14268,N_14138,N_14091);
or U14269 (N_14269,N_14141,N_14081);
nor U14270 (N_14270,N_14034,N_14033);
nor U14271 (N_14271,N_14135,N_14043);
nor U14272 (N_14272,N_14158,N_14092);
xor U14273 (N_14273,N_14057,N_14096);
and U14274 (N_14274,N_14175,N_14180);
or U14275 (N_14275,N_14142,N_14061);
xnor U14276 (N_14276,N_14132,N_14166);
xnor U14277 (N_14277,N_14113,N_14164);
and U14278 (N_14278,N_14004,N_14188);
xor U14279 (N_14279,N_14105,N_14087);
or U14280 (N_14280,N_14065,N_14068);
nor U14281 (N_14281,N_14123,N_14110);
and U14282 (N_14282,N_14102,N_14170);
nor U14283 (N_14283,N_14178,N_14055);
nor U14284 (N_14284,N_14169,N_14131);
nand U14285 (N_14285,N_14007,N_14111);
nand U14286 (N_14286,N_14093,N_14006);
nor U14287 (N_14287,N_14090,N_14109);
and U14288 (N_14288,N_14140,N_14056);
and U14289 (N_14289,N_14045,N_14058);
nand U14290 (N_14290,N_14015,N_14127);
nor U14291 (N_14291,N_14042,N_14017);
nand U14292 (N_14292,N_14059,N_14179);
xor U14293 (N_14293,N_14103,N_14159);
nand U14294 (N_14294,N_14124,N_14083);
or U14295 (N_14295,N_14144,N_14027);
and U14296 (N_14296,N_14079,N_14189);
xnor U14297 (N_14297,N_14160,N_14143);
nor U14298 (N_14298,N_14155,N_14196);
and U14299 (N_14299,N_14137,N_14018);
xnor U14300 (N_14300,N_14104,N_14045);
nor U14301 (N_14301,N_14162,N_14190);
nand U14302 (N_14302,N_14073,N_14051);
nor U14303 (N_14303,N_14001,N_14166);
or U14304 (N_14304,N_14163,N_14056);
xnor U14305 (N_14305,N_14001,N_14113);
and U14306 (N_14306,N_14089,N_14109);
nand U14307 (N_14307,N_14011,N_14082);
or U14308 (N_14308,N_14047,N_14124);
nor U14309 (N_14309,N_14196,N_14101);
nand U14310 (N_14310,N_14065,N_14039);
or U14311 (N_14311,N_14166,N_14109);
nand U14312 (N_14312,N_14117,N_14003);
or U14313 (N_14313,N_14055,N_14131);
or U14314 (N_14314,N_14111,N_14017);
or U14315 (N_14315,N_14165,N_14126);
and U14316 (N_14316,N_14130,N_14119);
xor U14317 (N_14317,N_14008,N_14125);
and U14318 (N_14318,N_14172,N_14007);
nand U14319 (N_14319,N_14060,N_14098);
nand U14320 (N_14320,N_14055,N_14154);
or U14321 (N_14321,N_14062,N_14094);
and U14322 (N_14322,N_14095,N_14048);
xor U14323 (N_14323,N_14047,N_14053);
nand U14324 (N_14324,N_14051,N_14137);
or U14325 (N_14325,N_14069,N_14190);
nor U14326 (N_14326,N_14133,N_14007);
nor U14327 (N_14327,N_14005,N_14057);
or U14328 (N_14328,N_14083,N_14126);
nand U14329 (N_14329,N_14051,N_14006);
or U14330 (N_14330,N_14017,N_14027);
and U14331 (N_14331,N_14125,N_14107);
and U14332 (N_14332,N_14188,N_14032);
nand U14333 (N_14333,N_14040,N_14191);
nor U14334 (N_14334,N_14063,N_14187);
nor U14335 (N_14335,N_14077,N_14118);
and U14336 (N_14336,N_14131,N_14058);
or U14337 (N_14337,N_14054,N_14100);
or U14338 (N_14338,N_14090,N_14181);
and U14339 (N_14339,N_14004,N_14181);
nor U14340 (N_14340,N_14089,N_14077);
and U14341 (N_14341,N_14065,N_14058);
nor U14342 (N_14342,N_14063,N_14026);
and U14343 (N_14343,N_14072,N_14001);
or U14344 (N_14344,N_14156,N_14192);
and U14345 (N_14345,N_14082,N_14155);
and U14346 (N_14346,N_14157,N_14071);
nor U14347 (N_14347,N_14011,N_14018);
nor U14348 (N_14348,N_14171,N_14125);
xor U14349 (N_14349,N_14058,N_14028);
and U14350 (N_14350,N_14133,N_14011);
and U14351 (N_14351,N_14123,N_14157);
and U14352 (N_14352,N_14053,N_14001);
nand U14353 (N_14353,N_14140,N_14147);
xor U14354 (N_14354,N_14125,N_14169);
and U14355 (N_14355,N_14063,N_14112);
nor U14356 (N_14356,N_14123,N_14079);
nand U14357 (N_14357,N_14114,N_14134);
and U14358 (N_14358,N_14059,N_14008);
xnor U14359 (N_14359,N_14159,N_14157);
and U14360 (N_14360,N_14070,N_14057);
and U14361 (N_14361,N_14131,N_14033);
or U14362 (N_14362,N_14111,N_14075);
nor U14363 (N_14363,N_14016,N_14124);
and U14364 (N_14364,N_14031,N_14002);
and U14365 (N_14365,N_14128,N_14063);
or U14366 (N_14366,N_14022,N_14183);
xnor U14367 (N_14367,N_14016,N_14038);
xor U14368 (N_14368,N_14178,N_14027);
and U14369 (N_14369,N_14087,N_14155);
nor U14370 (N_14370,N_14193,N_14120);
nor U14371 (N_14371,N_14180,N_14103);
and U14372 (N_14372,N_14019,N_14172);
nand U14373 (N_14373,N_14129,N_14051);
or U14374 (N_14374,N_14010,N_14065);
nor U14375 (N_14375,N_14193,N_14089);
and U14376 (N_14376,N_14133,N_14077);
nand U14377 (N_14377,N_14071,N_14147);
xor U14378 (N_14378,N_14144,N_14158);
nand U14379 (N_14379,N_14036,N_14065);
nand U14380 (N_14380,N_14097,N_14126);
nor U14381 (N_14381,N_14057,N_14090);
and U14382 (N_14382,N_14076,N_14080);
or U14383 (N_14383,N_14014,N_14153);
nor U14384 (N_14384,N_14144,N_14194);
nand U14385 (N_14385,N_14171,N_14135);
xnor U14386 (N_14386,N_14025,N_14184);
nand U14387 (N_14387,N_14015,N_14183);
and U14388 (N_14388,N_14170,N_14119);
nand U14389 (N_14389,N_14022,N_14023);
and U14390 (N_14390,N_14172,N_14000);
nand U14391 (N_14391,N_14094,N_14187);
nand U14392 (N_14392,N_14174,N_14177);
nor U14393 (N_14393,N_14027,N_14015);
nand U14394 (N_14394,N_14189,N_14050);
nand U14395 (N_14395,N_14168,N_14164);
xor U14396 (N_14396,N_14178,N_14053);
or U14397 (N_14397,N_14055,N_14197);
xor U14398 (N_14398,N_14146,N_14140);
nand U14399 (N_14399,N_14023,N_14143);
or U14400 (N_14400,N_14329,N_14376);
or U14401 (N_14401,N_14302,N_14341);
xnor U14402 (N_14402,N_14338,N_14215);
or U14403 (N_14403,N_14210,N_14282);
nand U14404 (N_14404,N_14292,N_14333);
and U14405 (N_14405,N_14253,N_14377);
nor U14406 (N_14406,N_14238,N_14205);
or U14407 (N_14407,N_14315,N_14395);
xor U14408 (N_14408,N_14340,N_14219);
nor U14409 (N_14409,N_14263,N_14311);
xnor U14410 (N_14410,N_14360,N_14204);
nor U14411 (N_14411,N_14339,N_14332);
nand U14412 (N_14412,N_14289,N_14211);
and U14413 (N_14413,N_14391,N_14266);
nand U14414 (N_14414,N_14378,N_14290);
xor U14415 (N_14415,N_14330,N_14288);
nor U14416 (N_14416,N_14264,N_14248);
and U14417 (N_14417,N_14231,N_14303);
nor U14418 (N_14418,N_14304,N_14362);
xor U14419 (N_14419,N_14223,N_14370);
nand U14420 (N_14420,N_14374,N_14269);
or U14421 (N_14421,N_14326,N_14310);
or U14422 (N_14422,N_14232,N_14257);
xor U14423 (N_14423,N_14229,N_14388);
or U14424 (N_14424,N_14389,N_14321);
xnor U14425 (N_14425,N_14261,N_14364);
or U14426 (N_14426,N_14236,N_14274);
nor U14427 (N_14427,N_14312,N_14201);
nand U14428 (N_14428,N_14278,N_14367);
nor U14429 (N_14429,N_14255,N_14213);
or U14430 (N_14430,N_14314,N_14281);
or U14431 (N_14431,N_14291,N_14273);
nand U14432 (N_14432,N_14275,N_14298);
nand U14433 (N_14433,N_14297,N_14383);
nor U14434 (N_14434,N_14368,N_14375);
and U14435 (N_14435,N_14317,N_14235);
or U14436 (N_14436,N_14397,N_14319);
or U14437 (N_14437,N_14347,N_14366);
or U14438 (N_14438,N_14399,N_14202);
or U14439 (N_14439,N_14209,N_14299);
nor U14440 (N_14440,N_14349,N_14203);
nand U14441 (N_14441,N_14252,N_14343);
xnor U14442 (N_14442,N_14277,N_14342);
or U14443 (N_14443,N_14355,N_14286);
nand U14444 (N_14444,N_14337,N_14225);
nor U14445 (N_14445,N_14350,N_14307);
nand U14446 (N_14446,N_14300,N_14301);
nor U14447 (N_14447,N_14363,N_14379);
xnor U14448 (N_14448,N_14331,N_14354);
or U14449 (N_14449,N_14228,N_14243);
and U14450 (N_14450,N_14287,N_14335);
nand U14451 (N_14451,N_14345,N_14320);
or U14452 (N_14452,N_14365,N_14258);
xnor U14453 (N_14453,N_14226,N_14369);
xor U14454 (N_14454,N_14259,N_14272);
nand U14455 (N_14455,N_14230,N_14280);
xor U14456 (N_14456,N_14240,N_14262);
nor U14457 (N_14457,N_14316,N_14295);
xor U14458 (N_14458,N_14305,N_14260);
and U14459 (N_14459,N_14398,N_14309);
and U14460 (N_14460,N_14212,N_14390);
nor U14461 (N_14461,N_14351,N_14271);
nand U14462 (N_14462,N_14250,N_14393);
nand U14463 (N_14463,N_14254,N_14328);
nand U14464 (N_14464,N_14247,N_14256);
or U14465 (N_14465,N_14200,N_14344);
nand U14466 (N_14466,N_14284,N_14352);
nor U14467 (N_14467,N_14270,N_14380);
nor U14468 (N_14468,N_14239,N_14313);
xnor U14469 (N_14469,N_14249,N_14318);
and U14470 (N_14470,N_14265,N_14382);
and U14471 (N_14471,N_14371,N_14387);
nor U14472 (N_14472,N_14306,N_14283);
and U14473 (N_14473,N_14233,N_14386);
xnor U14474 (N_14474,N_14356,N_14206);
or U14475 (N_14475,N_14242,N_14324);
nand U14476 (N_14476,N_14373,N_14267);
nand U14477 (N_14477,N_14336,N_14285);
nor U14478 (N_14478,N_14241,N_14276);
and U14479 (N_14479,N_14218,N_14348);
and U14480 (N_14480,N_14244,N_14308);
or U14481 (N_14481,N_14207,N_14214);
or U14482 (N_14482,N_14334,N_14357);
or U14483 (N_14483,N_14361,N_14372);
nand U14484 (N_14484,N_14293,N_14359);
and U14485 (N_14485,N_14251,N_14392);
xnor U14486 (N_14486,N_14384,N_14222);
xnor U14487 (N_14487,N_14227,N_14217);
nand U14488 (N_14488,N_14245,N_14208);
or U14489 (N_14489,N_14234,N_14327);
xnor U14490 (N_14490,N_14394,N_14381);
and U14491 (N_14491,N_14296,N_14220);
and U14492 (N_14492,N_14246,N_14396);
or U14493 (N_14493,N_14322,N_14323);
nor U14494 (N_14494,N_14325,N_14224);
nor U14495 (N_14495,N_14237,N_14279);
xor U14496 (N_14496,N_14268,N_14385);
xor U14497 (N_14497,N_14358,N_14216);
nor U14498 (N_14498,N_14346,N_14221);
nor U14499 (N_14499,N_14353,N_14294);
nand U14500 (N_14500,N_14235,N_14309);
xnor U14501 (N_14501,N_14292,N_14255);
nor U14502 (N_14502,N_14313,N_14395);
and U14503 (N_14503,N_14240,N_14326);
or U14504 (N_14504,N_14276,N_14291);
nor U14505 (N_14505,N_14302,N_14230);
or U14506 (N_14506,N_14278,N_14314);
nand U14507 (N_14507,N_14264,N_14236);
xor U14508 (N_14508,N_14224,N_14328);
or U14509 (N_14509,N_14201,N_14318);
xor U14510 (N_14510,N_14224,N_14396);
nor U14511 (N_14511,N_14382,N_14219);
nand U14512 (N_14512,N_14347,N_14256);
or U14513 (N_14513,N_14207,N_14206);
and U14514 (N_14514,N_14343,N_14220);
and U14515 (N_14515,N_14300,N_14316);
nor U14516 (N_14516,N_14338,N_14281);
nor U14517 (N_14517,N_14277,N_14399);
nand U14518 (N_14518,N_14330,N_14243);
or U14519 (N_14519,N_14202,N_14241);
or U14520 (N_14520,N_14371,N_14336);
xor U14521 (N_14521,N_14307,N_14343);
nor U14522 (N_14522,N_14370,N_14249);
and U14523 (N_14523,N_14335,N_14376);
or U14524 (N_14524,N_14283,N_14313);
and U14525 (N_14525,N_14203,N_14311);
nor U14526 (N_14526,N_14261,N_14391);
nor U14527 (N_14527,N_14320,N_14352);
xor U14528 (N_14528,N_14317,N_14369);
xor U14529 (N_14529,N_14205,N_14307);
nor U14530 (N_14530,N_14369,N_14242);
nand U14531 (N_14531,N_14397,N_14357);
nor U14532 (N_14532,N_14392,N_14353);
nand U14533 (N_14533,N_14387,N_14293);
or U14534 (N_14534,N_14324,N_14300);
nor U14535 (N_14535,N_14340,N_14317);
xor U14536 (N_14536,N_14309,N_14298);
and U14537 (N_14537,N_14302,N_14244);
nand U14538 (N_14538,N_14297,N_14305);
or U14539 (N_14539,N_14312,N_14317);
xnor U14540 (N_14540,N_14348,N_14342);
nand U14541 (N_14541,N_14273,N_14228);
nand U14542 (N_14542,N_14325,N_14221);
nor U14543 (N_14543,N_14391,N_14263);
and U14544 (N_14544,N_14211,N_14319);
and U14545 (N_14545,N_14290,N_14358);
nand U14546 (N_14546,N_14247,N_14359);
or U14547 (N_14547,N_14330,N_14345);
and U14548 (N_14548,N_14358,N_14228);
or U14549 (N_14549,N_14286,N_14386);
nor U14550 (N_14550,N_14202,N_14233);
nand U14551 (N_14551,N_14382,N_14277);
nor U14552 (N_14552,N_14282,N_14298);
and U14553 (N_14553,N_14378,N_14381);
nor U14554 (N_14554,N_14307,N_14256);
and U14555 (N_14555,N_14255,N_14288);
or U14556 (N_14556,N_14328,N_14260);
nor U14557 (N_14557,N_14332,N_14284);
or U14558 (N_14558,N_14295,N_14370);
nand U14559 (N_14559,N_14291,N_14325);
xnor U14560 (N_14560,N_14333,N_14342);
nor U14561 (N_14561,N_14218,N_14228);
and U14562 (N_14562,N_14322,N_14218);
and U14563 (N_14563,N_14357,N_14237);
and U14564 (N_14564,N_14377,N_14260);
or U14565 (N_14565,N_14352,N_14298);
nand U14566 (N_14566,N_14230,N_14312);
nand U14567 (N_14567,N_14374,N_14369);
and U14568 (N_14568,N_14232,N_14342);
nand U14569 (N_14569,N_14278,N_14271);
nor U14570 (N_14570,N_14240,N_14331);
and U14571 (N_14571,N_14372,N_14397);
xnor U14572 (N_14572,N_14200,N_14332);
xor U14573 (N_14573,N_14330,N_14362);
or U14574 (N_14574,N_14346,N_14211);
and U14575 (N_14575,N_14360,N_14280);
nor U14576 (N_14576,N_14360,N_14346);
and U14577 (N_14577,N_14259,N_14341);
or U14578 (N_14578,N_14384,N_14329);
and U14579 (N_14579,N_14272,N_14276);
nor U14580 (N_14580,N_14248,N_14352);
and U14581 (N_14581,N_14271,N_14366);
nand U14582 (N_14582,N_14356,N_14277);
or U14583 (N_14583,N_14325,N_14269);
and U14584 (N_14584,N_14366,N_14320);
or U14585 (N_14585,N_14339,N_14270);
or U14586 (N_14586,N_14336,N_14276);
and U14587 (N_14587,N_14203,N_14239);
or U14588 (N_14588,N_14232,N_14285);
nor U14589 (N_14589,N_14201,N_14374);
nand U14590 (N_14590,N_14337,N_14328);
xnor U14591 (N_14591,N_14217,N_14388);
nand U14592 (N_14592,N_14344,N_14285);
or U14593 (N_14593,N_14290,N_14368);
and U14594 (N_14594,N_14274,N_14218);
or U14595 (N_14595,N_14322,N_14344);
xor U14596 (N_14596,N_14343,N_14306);
nor U14597 (N_14597,N_14247,N_14250);
xor U14598 (N_14598,N_14356,N_14389);
nand U14599 (N_14599,N_14211,N_14359);
nor U14600 (N_14600,N_14449,N_14400);
nand U14601 (N_14601,N_14438,N_14534);
nor U14602 (N_14602,N_14479,N_14556);
nand U14603 (N_14603,N_14420,N_14467);
nor U14604 (N_14604,N_14464,N_14549);
nand U14605 (N_14605,N_14411,N_14487);
nor U14606 (N_14606,N_14521,N_14440);
nand U14607 (N_14607,N_14514,N_14519);
nand U14608 (N_14608,N_14410,N_14581);
nand U14609 (N_14609,N_14493,N_14558);
or U14610 (N_14610,N_14542,N_14566);
xor U14611 (N_14611,N_14474,N_14555);
or U14612 (N_14612,N_14585,N_14441);
nand U14613 (N_14613,N_14582,N_14481);
or U14614 (N_14614,N_14432,N_14494);
nand U14615 (N_14615,N_14430,N_14475);
and U14616 (N_14616,N_14588,N_14428);
xnor U14617 (N_14617,N_14593,N_14522);
nor U14618 (N_14618,N_14553,N_14431);
nand U14619 (N_14619,N_14482,N_14417);
nor U14620 (N_14620,N_14447,N_14590);
nor U14621 (N_14621,N_14564,N_14586);
nand U14622 (N_14622,N_14540,N_14403);
nor U14623 (N_14623,N_14426,N_14433);
and U14624 (N_14624,N_14473,N_14509);
nand U14625 (N_14625,N_14418,N_14483);
and U14626 (N_14626,N_14520,N_14416);
or U14627 (N_14627,N_14486,N_14414);
nor U14628 (N_14628,N_14453,N_14527);
nand U14629 (N_14629,N_14407,N_14557);
and U14630 (N_14630,N_14543,N_14594);
or U14631 (N_14631,N_14531,N_14434);
nor U14632 (N_14632,N_14471,N_14528);
xor U14633 (N_14633,N_14508,N_14435);
nand U14634 (N_14634,N_14406,N_14450);
xnor U14635 (N_14635,N_14496,N_14423);
xnor U14636 (N_14636,N_14548,N_14415);
nand U14637 (N_14637,N_14589,N_14560);
and U14638 (N_14638,N_14460,N_14462);
nor U14639 (N_14639,N_14525,N_14476);
or U14640 (N_14640,N_14478,N_14529);
or U14641 (N_14641,N_14500,N_14577);
or U14642 (N_14642,N_14584,N_14429);
nand U14643 (N_14643,N_14498,N_14404);
and U14644 (N_14644,N_14468,N_14472);
and U14645 (N_14645,N_14554,N_14569);
nor U14646 (N_14646,N_14545,N_14597);
nand U14647 (N_14647,N_14574,N_14532);
xor U14648 (N_14648,N_14515,N_14541);
or U14649 (N_14649,N_14567,N_14537);
nor U14650 (N_14650,N_14446,N_14413);
nor U14651 (N_14651,N_14511,N_14568);
nor U14652 (N_14652,N_14442,N_14523);
and U14653 (N_14653,N_14533,N_14591);
and U14654 (N_14654,N_14427,N_14562);
nor U14655 (N_14655,N_14492,N_14491);
nor U14656 (N_14656,N_14477,N_14524);
xor U14657 (N_14657,N_14536,N_14485);
nor U14658 (N_14658,N_14439,N_14576);
or U14659 (N_14659,N_14547,N_14490);
and U14660 (N_14660,N_14570,N_14445);
or U14661 (N_14661,N_14437,N_14402);
nand U14662 (N_14662,N_14513,N_14512);
and U14663 (N_14663,N_14510,N_14497);
xnor U14664 (N_14664,N_14495,N_14550);
xnor U14665 (N_14665,N_14405,N_14559);
or U14666 (N_14666,N_14459,N_14458);
nand U14667 (N_14667,N_14573,N_14424);
nor U14668 (N_14668,N_14526,N_14580);
and U14669 (N_14669,N_14565,N_14452);
nand U14670 (N_14670,N_14561,N_14448);
xor U14671 (N_14671,N_14518,N_14401);
nand U14672 (N_14672,N_14501,N_14408);
nand U14673 (N_14673,N_14469,N_14425);
xnor U14674 (N_14674,N_14578,N_14507);
xnor U14675 (N_14675,N_14599,N_14595);
nor U14676 (N_14676,N_14422,N_14546);
and U14677 (N_14677,N_14436,N_14579);
or U14678 (N_14678,N_14502,N_14575);
or U14679 (N_14679,N_14444,N_14457);
xor U14680 (N_14680,N_14596,N_14505);
nor U14681 (N_14681,N_14598,N_14480);
or U14682 (N_14682,N_14504,N_14489);
xnor U14683 (N_14683,N_14443,N_14419);
xor U14684 (N_14684,N_14592,N_14517);
nor U14685 (N_14685,N_14551,N_14461);
or U14686 (N_14686,N_14409,N_14587);
and U14687 (N_14687,N_14456,N_14503);
or U14688 (N_14688,N_14572,N_14516);
xnor U14689 (N_14689,N_14539,N_14535);
and U14690 (N_14690,N_14465,N_14544);
and U14691 (N_14691,N_14455,N_14470);
xor U14692 (N_14692,N_14563,N_14451);
or U14693 (N_14693,N_14499,N_14488);
and U14694 (N_14694,N_14538,N_14466);
or U14695 (N_14695,N_14530,N_14421);
nand U14696 (N_14696,N_14506,N_14463);
or U14697 (N_14697,N_14571,N_14412);
nand U14698 (N_14698,N_14454,N_14484);
xnor U14699 (N_14699,N_14583,N_14552);
and U14700 (N_14700,N_14571,N_14497);
nor U14701 (N_14701,N_14553,N_14543);
xnor U14702 (N_14702,N_14550,N_14424);
nor U14703 (N_14703,N_14504,N_14422);
and U14704 (N_14704,N_14402,N_14424);
or U14705 (N_14705,N_14415,N_14457);
xnor U14706 (N_14706,N_14538,N_14429);
nand U14707 (N_14707,N_14486,N_14543);
xnor U14708 (N_14708,N_14562,N_14546);
xor U14709 (N_14709,N_14478,N_14597);
and U14710 (N_14710,N_14432,N_14590);
nor U14711 (N_14711,N_14450,N_14401);
xor U14712 (N_14712,N_14421,N_14532);
xnor U14713 (N_14713,N_14462,N_14533);
or U14714 (N_14714,N_14576,N_14585);
or U14715 (N_14715,N_14539,N_14465);
xnor U14716 (N_14716,N_14516,N_14410);
and U14717 (N_14717,N_14436,N_14502);
xor U14718 (N_14718,N_14476,N_14582);
xor U14719 (N_14719,N_14599,N_14439);
and U14720 (N_14720,N_14422,N_14551);
nand U14721 (N_14721,N_14499,N_14574);
xnor U14722 (N_14722,N_14517,N_14463);
and U14723 (N_14723,N_14572,N_14411);
nand U14724 (N_14724,N_14421,N_14524);
nor U14725 (N_14725,N_14476,N_14429);
nor U14726 (N_14726,N_14427,N_14526);
and U14727 (N_14727,N_14425,N_14480);
and U14728 (N_14728,N_14527,N_14578);
nor U14729 (N_14729,N_14524,N_14434);
nor U14730 (N_14730,N_14432,N_14516);
nor U14731 (N_14731,N_14533,N_14486);
xnor U14732 (N_14732,N_14493,N_14509);
nand U14733 (N_14733,N_14514,N_14447);
nand U14734 (N_14734,N_14417,N_14458);
xnor U14735 (N_14735,N_14555,N_14464);
xnor U14736 (N_14736,N_14443,N_14487);
nand U14737 (N_14737,N_14400,N_14421);
nor U14738 (N_14738,N_14505,N_14494);
nor U14739 (N_14739,N_14512,N_14558);
or U14740 (N_14740,N_14464,N_14504);
and U14741 (N_14741,N_14570,N_14488);
xor U14742 (N_14742,N_14411,N_14433);
and U14743 (N_14743,N_14573,N_14578);
nor U14744 (N_14744,N_14414,N_14509);
or U14745 (N_14745,N_14445,N_14487);
nand U14746 (N_14746,N_14473,N_14472);
and U14747 (N_14747,N_14569,N_14547);
or U14748 (N_14748,N_14490,N_14446);
and U14749 (N_14749,N_14442,N_14448);
nor U14750 (N_14750,N_14462,N_14514);
or U14751 (N_14751,N_14531,N_14508);
nor U14752 (N_14752,N_14576,N_14544);
nor U14753 (N_14753,N_14432,N_14490);
xor U14754 (N_14754,N_14470,N_14416);
nand U14755 (N_14755,N_14520,N_14421);
nand U14756 (N_14756,N_14499,N_14565);
xor U14757 (N_14757,N_14485,N_14547);
nor U14758 (N_14758,N_14571,N_14513);
or U14759 (N_14759,N_14506,N_14528);
nand U14760 (N_14760,N_14564,N_14581);
nor U14761 (N_14761,N_14423,N_14540);
nand U14762 (N_14762,N_14416,N_14598);
and U14763 (N_14763,N_14469,N_14548);
and U14764 (N_14764,N_14517,N_14491);
or U14765 (N_14765,N_14567,N_14581);
xor U14766 (N_14766,N_14572,N_14458);
nand U14767 (N_14767,N_14419,N_14459);
nor U14768 (N_14768,N_14424,N_14585);
and U14769 (N_14769,N_14542,N_14589);
nand U14770 (N_14770,N_14590,N_14478);
and U14771 (N_14771,N_14413,N_14455);
nor U14772 (N_14772,N_14513,N_14523);
xor U14773 (N_14773,N_14403,N_14572);
nand U14774 (N_14774,N_14421,N_14568);
or U14775 (N_14775,N_14555,N_14556);
and U14776 (N_14776,N_14432,N_14483);
nor U14777 (N_14777,N_14570,N_14547);
nor U14778 (N_14778,N_14591,N_14574);
xnor U14779 (N_14779,N_14451,N_14491);
nand U14780 (N_14780,N_14556,N_14558);
nand U14781 (N_14781,N_14534,N_14531);
xor U14782 (N_14782,N_14458,N_14560);
nand U14783 (N_14783,N_14476,N_14488);
nand U14784 (N_14784,N_14591,N_14537);
and U14785 (N_14785,N_14539,N_14592);
or U14786 (N_14786,N_14430,N_14417);
xnor U14787 (N_14787,N_14527,N_14427);
nor U14788 (N_14788,N_14586,N_14465);
xor U14789 (N_14789,N_14435,N_14449);
and U14790 (N_14790,N_14455,N_14438);
nor U14791 (N_14791,N_14561,N_14454);
xnor U14792 (N_14792,N_14445,N_14545);
and U14793 (N_14793,N_14532,N_14514);
and U14794 (N_14794,N_14418,N_14404);
and U14795 (N_14795,N_14484,N_14542);
nand U14796 (N_14796,N_14542,N_14517);
and U14797 (N_14797,N_14549,N_14405);
or U14798 (N_14798,N_14446,N_14570);
and U14799 (N_14799,N_14553,N_14591);
and U14800 (N_14800,N_14608,N_14773);
or U14801 (N_14801,N_14691,N_14718);
nor U14802 (N_14802,N_14749,N_14689);
or U14803 (N_14803,N_14686,N_14673);
xor U14804 (N_14804,N_14699,N_14603);
nand U14805 (N_14805,N_14756,N_14634);
xor U14806 (N_14806,N_14627,N_14740);
xnor U14807 (N_14807,N_14703,N_14776);
nand U14808 (N_14808,N_14650,N_14625);
or U14809 (N_14809,N_14794,N_14619);
nor U14810 (N_14810,N_14713,N_14640);
nor U14811 (N_14811,N_14693,N_14618);
nor U14812 (N_14812,N_14628,N_14624);
xnor U14813 (N_14813,N_14787,N_14796);
or U14814 (N_14814,N_14760,N_14626);
xor U14815 (N_14815,N_14651,N_14681);
or U14816 (N_14816,N_14623,N_14652);
or U14817 (N_14817,N_14731,N_14637);
nand U14818 (N_14818,N_14751,N_14752);
nor U14819 (N_14819,N_14738,N_14757);
and U14820 (N_14820,N_14677,N_14670);
nand U14821 (N_14821,N_14679,N_14607);
and U14822 (N_14822,N_14744,N_14600);
nand U14823 (N_14823,N_14768,N_14636);
nor U14824 (N_14824,N_14741,N_14659);
nor U14825 (N_14825,N_14784,N_14641);
nor U14826 (N_14826,N_14780,N_14754);
xor U14827 (N_14827,N_14667,N_14606);
and U14828 (N_14828,N_14622,N_14615);
xnor U14829 (N_14829,N_14633,N_14632);
nand U14830 (N_14830,N_14669,N_14655);
nand U14831 (N_14831,N_14629,N_14705);
nor U14832 (N_14832,N_14702,N_14662);
or U14833 (N_14833,N_14671,N_14621);
and U14834 (N_14834,N_14609,N_14658);
xor U14835 (N_14835,N_14732,N_14704);
xnor U14836 (N_14836,N_14770,N_14674);
and U14837 (N_14837,N_14762,N_14721);
nand U14838 (N_14838,N_14646,N_14714);
nor U14839 (N_14839,N_14730,N_14727);
and U14840 (N_14840,N_14715,N_14672);
or U14841 (N_14841,N_14778,N_14734);
and U14842 (N_14842,N_14680,N_14635);
and U14843 (N_14843,N_14775,N_14765);
xnor U14844 (N_14844,N_14645,N_14663);
or U14845 (N_14845,N_14767,N_14706);
and U14846 (N_14846,N_14642,N_14725);
and U14847 (N_14847,N_14638,N_14648);
nand U14848 (N_14848,N_14722,N_14656);
nor U14849 (N_14849,N_14736,N_14712);
xor U14850 (N_14850,N_14654,N_14610);
nor U14851 (N_14851,N_14747,N_14789);
xor U14852 (N_14852,N_14717,N_14755);
nand U14853 (N_14853,N_14708,N_14783);
nor U14854 (N_14854,N_14664,N_14720);
and U14855 (N_14855,N_14798,N_14675);
or U14856 (N_14856,N_14737,N_14716);
nor U14857 (N_14857,N_14742,N_14695);
and U14858 (N_14858,N_14792,N_14631);
nand U14859 (N_14859,N_14657,N_14753);
xor U14860 (N_14860,N_14639,N_14769);
or U14861 (N_14861,N_14779,N_14684);
nand U14862 (N_14862,N_14795,N_14660);
and U14863 (N_14863,N_14698,N_14649);
or U14864 (N_14864,N_14647,N_14682);
nor U14865 (N_14865,N_14678,N_14766);
nor U14866 (N_14866,N_14764,N_14685);
nand U14867 (N_14867,N_14611,N_14643);
or U14868 (N_14868,N_14797,N_14791);
nor U14869 (N_14869,N_14701,N_14602);
xnor U14870 (N_14870,N_14666,N_14772);
nand U14871 (N_14871,N_14735,N_14758);
nor U14872 (N_14872,N_14692,N_14771);
xor U14873 (N_14873,N_14687,N_14745);
and U14874 (N_14874,N_14733,N_14750);
xnor U14875 (N_14875,N_14788,N_14700);
and U14876 (N_14876,N_14694,N_14653);
nand U14877 (N_14877,N_14729,N_14616);
and U14878 (N_14878,N_14739,N_14799);
and U14879 (N_14879,N_14707,N_14763);
or U14880 (N_14880,N_14785,N_14761);
or U14881 (N_14881,N_14724,N_14746);
xnor U14882 (N_14882,N_14604,N_14697);
and U14883 (N_14883,N_14696,N_14710);
or U14884 (N_14884,N_14728,N_14759);
or U14885 (N_14885,N_14612,N_14774);
nand U14886 (N_14886,N_14743,N_14782);
or U14887 (N_14887,N_14661,N_14690);
or U14888 (N_14888,N_14683,N_14781);
nand U14889 (N_14889,N_14676,N_14605);
nor U14890 (N_14890,N_14665,N_14630);
nor U14891 (N_14891,N_14711,N_14777);
nor U14892 (N_14892,N_14709,N_14644);
or U14893 (N_14893,N_14614,N_14719);
and U14894 (N_14894,N_14793,N_14688);
nor U14895 (N_14895,N_14748,N_14613);
xor U14896 (N_14896,N_14668,N_14601);
nor U14897 (N_14897,N_14786,N_14620);
or U14898 (N_14898,N_14726,N_14790);
or U14899 (N_14899,N_14617,N_14723);
or U14900 (N_14900,N_14602,N_14759);
xor U14901 (N_14901,N_14781,N_14610);
nand U14902 (N_14902,N_14769,N_14743);
or U14903 (N_14903,N_14633,N_14685);
nor U14904 (N_14904,N_14758,N_14757);
xor U14905 (N_14905,N_14622,N_14799);
nand U14906 (N_14906,N_14791,N_14650);
nor U14907 (N_14907,N_14702,N_14632);
nand U14908 (N_14908,N_14655,N_14657);
nor U14909 (N_14909,N_14678,N_14693);
nor U14910 (N_14910,N_14778,N_14718);
or U14911 (N_14911,N_14622,N_14651);
and U14912 (N_14912,N_14672,N_14651);
xor U14913 (N_14913,N_14663,N_14667);
nor U14914 (N_14914,N_14678,N_14703);
xnor U14915 (N_14915,N_14779,N_14750);
and U14916 (N_14916,N_14775,N_14617);
or U14917 (N_14917,N_14672,N_14676);
nand U14918 (N_14918,N_14684,N_14693);
or U14919 (N_14919,N_14630,N_14639);
nand U14920 (N_14920,N_14679,N_14664);
xor U14921 (N_14921,N_14717,N_14690);
and U14922 (N_14922,N_14694,N_14639);
xnor U14923 (N_14923,N_14705,N_14780);
nand U14924 (N_14924,N_14697,N_14660);
nand U14925 (N_14925,N_14722,N_14768);
and U14926 (N_14926,N_14715,N_14792);
nor U14927 (N_14927,N_14675,N_14785);
or U14928 (N_14928,N_14796,N_14795);
xor U14929 (N_14929,N_14601,N_14786);
nand U14930 (N_14930,N_14741,N_14631);
xor U14931 (N_14931,N_14610,N_14602);
and U14932 (N_14932,N_14759,N_14650);
nor U14933 (N_14933,N_14714,N_14661);
or U14934 (N_14934,N_14617,N_14741);
nor U14935 (N_14935,N_14722,N_14653);
or U14936 (N_14936,N_14701,N_14618);
nand U14937 (N_14937,N_14739,N_14607);
nor U14938 (N_14938,N_14788,N_14718);
or U14939 (N_14939,N_14776,N_14718);
and U14940 (N_14940,N_14680,N_14722);
nand U14941 (N_14941,N_14663,N_14746);
and U14942 (N_14942,N_14661,N_14682);
or U14943 (N_14943,N_14674,N_14709);
and U14944 (N_14944,N_14690,N_14767);
nor U14945 (N_14945,N_14608,N_14779);
and U14946 (N_14946,N_14671,N_14614);
and U14947 (N_14947,N_14645,N_14782);
xnor U14948 (N_14948,N_14746,N_14720);
nand U14949 (N_14949,N_14690,N_14730);
and U14950 (N_14950,N_14627,N_14739);
nor U14951 (N_14951,N_14746,N_14752);
or U14952 (N_14952,N_14614,N_14705);
nor U14953 (N_14953,N_14675,N_14710);
nor U14954 (N_14954,N_14606,N_14761);
and U14955 (N_14955,N_14750,N_14773);
xnor U14956 (N_14956,N_14747,N_14601);
xor U14957 (N_14957,N_14732,N_14652);
or U14958 (N_14958,N_14641,N_14750);
or U14959 (N_14959,N_14601,N_14607);
nor U14960 (N_14960,N_14785,N_14799);
and U14961 (N_14961,N_14729,N_14766);
nand U14962 (N_14962,N_14754,N_14704);
xor U14963 (N_14963,N_14772,N_14718);
or U14964 (N_14964,N_14635,N_14777);
xnor U14965 (N_14965,N_14665,N_14788);
xnor U14966 (N_14966,N_14705,N_14764);
nor U14967 (N_14967,N_14783,N_14771);
or U14968 (N_14968,N_14789,N_14648);
or U14969 (N_14969,N_14684,N_14695);
and U14970 (N_14970,N_14739,N_14727);
nand U14971 (N_14971,N_14637,N_14704);
nor U14972 (N_14972,N_14631,N_14659);
nor U14973 (N_14973,N_14703,N_14793);
nor U14974 (N_14974,N_14627,N_14625);
or U14975 (N_14975,N_14747,N_14672);
nand U14976 (N_14976,N_14665,N_14620);
xor U14977 (N_14977,N_14785,N_14611);
nand U14978 (N_14978,N_14712,N_14691);
and U14979 (N_14979,N_14714,N_14716);
xor U14980 (N_14980,N_14700,N_14732);
or U14981 (N_14981,N_14605,N_14642);
nand U14982 (N_14982,N_14626,N_14757);
nand U14983 (N_14983,N_14734,N_14789);
and U14984 (N_14984,N_14617,N_14735);
or U14985 (N_14985,N_14629,N_14653);
and U14986 (N_14986,N_14648,N_14735);
or U14987 (N_14987,N_14747,N_14696);
nor U14988 (N_14988,N_14771,N_14622);
and U14989 (N_14989,N_14608,N_14689);
nand U14990 (N_14990,N_14648,N_14624);
nand U14991 (N_14991,N_14656,N_14611);
nor U14992 (N_14992,N_14705,N_14634);
and U14993 (N_14993,N_14704,N_14722);
nor U14994 (N_14994,N_14665,N_14695);
and U14995 (N_14995,N_14758,N_14643);
nor U14996 (N_14996,N_14622,N_14789);
nand U14997 (N_14997,N_14772,N_14777);
xnor U14998 (N_14998,N_14608,N_14644);
nand U14999 (N_14999,N_14612,N_14716);
xnor U15000 (N_15000,N_14841,N_14958);
xnor U15001 (N_15001,N_14902,N_14827);
or U15002 (N_15002,N_14897,N_14952);
nand U15003 (N_15003,N_14853,N_14901);
nor U15004 (N_15004,N_14870,N_14935);
nand U15005 (N_15005,N_14984,N_14999);
nand U15006 (N_15006,N_14890,N_14925);
or U15007 (N_15007,N_14954,N_14851);
nor U15008 (N_15008,N_14863,N_14820);
or U15009 (N_15009,N_14943,N_14904);
or U15010 (N_15010,N_14873,N_14932);
nand U15011 (N_15011,N_14927,N_14881);
and U15012 (N_15012,N_14941,N_14970);
or U15013 (N_15013,N_14973,N_14911);
xnor U15014 (N_15014,N_14854,N_14822);
xor U15015 (N_15015,N_14899,N_14916);
xnor U15016 (N_15016,N_14974,N_14907);
nand U15017 (N_15017,N_14956,N_14805);
or U15018 (N_15018,N_14814,N_14844);
nor U15019 (N_15019,N_14919,N_14836);
nand U15020 (N_15020,N_14823,N_14884);
nor U15021 (N_15021,N_14903,N_14843);
and U15022 (N_15022,N_14846,N_14977);
nand U15023 (N_15023,N_14839,N_14869);
and U15024 (N_15024,N_14883,N_14990);
nor U15025 (N_15025,N_14963,N_14898);
and U15026 (N_15026,N_14921,N_14871);
or U15027 (N_15027,N_14972,N_14803);
and U15028 (N_15028,N_14910,N_14924);
nand U15029 (N_15029,N_14891,N_14939);
and U15030 (N_15030,N_14808,N_14842);
nand U15031 (N_15031,N_14961,N_14857);
nor U15032 (N_15032,N_14962,N_14892);
nand U15033 (N_15033,N_14926,N_14874);
nand U15034 (N_15034,N_14950,N_14845);
or U15035 (N_15035,N_14860,N_14937);
or U15036 (N_15036,N_14802,N_14989);
and U15037 (N_15037,N_14893,N_14872);
and U15038 (N_15038,N_14896,N_14988);
or U15039 (N_15039,N_14942,N_14982);
nor U15040 (N_15040,N_14966,N_14983);
or U15041 (N_15041,N_14900,N_14965);
or U15042 (N_15042,N_14929,N_14964);
or U15043 (N_15043,N_14824,N_14960);
and U15044 (N_15044,N_14905,N_14848);
and U15045 (N_15045,N_14914,N_14809);
xor U15046 (N_15046,N_14980,N_14850);
xor U15047 (N_15047,N_14922,N_14852);
and U15048 (N_15048,N_14951,N_14826);
nor U15049 (N_15049,N_14959,N_14878);
and U15050 (N_15050,N_14913,N_14815);
and U15051 (N_15051,N_14855,N_14993);
or U15052 (N_15052,N_14934,N_14923);
and U15053 (N_15053,N_14948,N_14976);
and U15054 (N_15054,N_14800,N_14995);
or U15055 (N_15055,N_14830,N_14981);
or U15056 (N_15056,N_14831,N_14997);
nand U15057 (N_15057,N_14940,N_14945);
or U15058 (N_15058,N_14864,N_14877);
and U15059 (N_15059,N_14986,N_14979);
nor U15060 (N_15060,N_14996,N_14985);
xor U15061 (N_15061,N_14859,N_14968);
xnor U15062 (N_15062,N_14832,N_14933);
xnor U15063 (N_15063,N_14807,N_14856);
xnor U15064 (N_15064,N_14862,N_14969);
nor U15065 (N_15065,N_14817,N_14806);
or U15066 (N_15066,N_14947,N_14888);
or U15067 (N_15067,N_14840,N_14917);
xor U15068 (N_15068,N_14931,N_14812);
xnor U15069 (N_15069,N_14920,N_14955);
and U15070 (N_15070,N_14825,N_14894);
nand U15071 (N_15071,N_14975,N_14810);
or U15072 (N_15072,N_14882,N_14938);
and U15073 (N_15073,N_14879,N_14944);
or U15074 (N_15074,N_14849,N_14994);
nor U15075 (N_15075,N_14978,N_14885);
nand U15076 (N_15076,N_14835,N_14967);
and U15077 (N_15077,N_14928,N_14909);
nand U15078 (N_15078,N_14837,N_14946);
or U15079 (N_15079,N_14953,N_14838);
nand U15080 (N_15080,N_14912,N_14887);
xor U15081 (N_15081,N_14987,N_14936);
and U15082 (N_15082,N_14918,N_14876);
xnor U15083 (N_15083,N_14828,N_14801);
nor U15084 (N_15084,N_14833,N_14971);
nor U15085 (N_15085,N_14861,N_14819);
or U15086 (N_15086,N_14847,N_14991);
and U15087 (N_15087,N_14865,N_14811);
or U15088 (N_15088,N_14818,N_14804);
nand U15089 (N_15089,N_14868,N_14998);
and U15090 (N_15090,N_14930,N_14866);
and U15091 (N_15091,N_14886,N_14992);
xnor U15092 (N_15092,N_14949,N_14908);
nor U15093 (N_15093,N_14915,N_14957);
nor U15094 (N_15094,N_14867,N_14875);
nor U15095 (N_15095,N_14889,N_14834);
or U15096 (N_15096,N_14813,N_14821);
xor U15097 (N_15097,N_14816,N_14895);
and U15098 (N_15098,N_14858,N_14829);
and U15099 (N_15099,N_14906,N_14880);
and U15100 (N_15100,N_14959,N_14901);
nor U15101 (N_15101,N_14854,N_14920);
nand U15102 (N_15102,N_14872,N_14863);
xor U15103 (N_15103,N_14881,N_14869);
nor U15104 (N_15104,N_14832,N_14978);
xor U15105 (N_15105,N_14991,N_14908);
and U15106 (N_15106,N_14948,N_14926);
and U15107 (N_15107,N_14825,N_14994);
or U15108 (N_15108,N_14800,N_14919);
nand U15109 (N_15109,N_14810,N_14808);
or U15110 (N_15110,N_14972,N_14810);
nand U15111 (N_15111,N_14927,N_14848);
nor U15112 (N_15112,N_14987,N_14845);
nand U15113 (N_15113,N_14890,N_14834);
and U15114 (N_15114,N_14911,N_14853);
or U15115 (N_15115,N_14990,N_14970);
nand U15116 (N_15116,N_14973,N_14937);
or U15117 (N_15117,N_14884,N_14864);
or U15118 (N_15118,N_14924,N_14935);
and U15119 (N_15119,N_14862,N_14990);
and U15120 (N_15120,N_14857,N_14858);
nand U15121 (N_15121,N_14910,N_14813);
or U15122 (N_15122,N_14831,N_14898);
and U15123 (N_15123,N_14990,N_14859);
and U15124 (N_15124,N_14835,N_14959);
or U15125 (N_15125,N_14892,N_14988);
nand U15126 (N_15126,N_14934,N_14999);
nand U15127 (N_15127,N_14932,N_14855);
xnor U15128 (N_15128,N_14820,N_14988);
nor U15129 (N_15129,N_14835,N_14861);
or U15130 (N_15130,N_14967,N_14881);
and U15131 (N_15131,N_14990,N_14820);
xor U15132 (N_15132,N_14993,N_14863);
or U15133 (N_15133,N_14907,N_14886);
nand U15134 (N_15134,N_14922,N_14817);
nor U15135 (N_15135,N_14933,N_14942);
and U15136 (N_15136,N_14847,N_14984);
nor U15137 (N_15137,N_14854,N_14894);
nor U15138 (N_15138,N_14832,N_14961);
nand U15139 (N_15139,N_14964,N_14890);
nand U15140 (N_15140,N_14820,N_14811);
nor U15141 (N_15141,N_14937,N_14931);
xor U15142 (N_15142,N_14941,N_14912);
nand U15143 (N_15143,N_14878,N_14949);
nand U15144 (N_15144,N_14852,N_14990);
xor U15145 (N_15145,N_14959,N_14902);
and U15146 (N_15146,N_14955,N_14950);
and U15147 (N_15147,N_14902,N_14873);
xnor U15148 (N_15148,N_14951,N_14827);
and U15149 (N_15149,N_14906,N_14876);
nor U15150 (N_15150,N_14883,N_14907);
or U15151 (N_15151,N_14846,N_14829);
xnor U15152 (N_15152,N_14940,N_14907);
or U15153 (N_15153,N_14905,N_14835);
nand U15154 (N_15154,N_14920,N_14928);
or U15155 (N_15155,N_14965,N_14916);
and U15156 (N_15156,N_14882,N_14866);
nor U15157 (N_15157,N_14924,N_14824);
xnor U15158 (N_15158,N_14862,N_14908);
xnor U15159 (N_15159,N_14810,N_14809);
and U15160 (N_15160,N_14873,N_14874);
or U15161 (N_15161,N_14848,N_14886);
nor U15162 (N_15162,N_14826,N_14974);
nor U15163 (N_15163,N_14898,N_14952);
or U15164 (N_15164,N_14955,N_14853);
nor U15165 (N_15165,N_14825,N_14835);
xnor U15166 (N_15166,N_14898,N_14846);
or U15167 (N_15167,N_14921,N_14840);
or U15168 (N_15168,N_14951,N_14933);
nand U15169 (N_15169,N_14814,N_14837);
and U15170 (N_15170,N_14934,N_14899);
and U15171 (N_15171,N_14998,N_14824);
nor U15172 (N_15172,N_14946,N_14880);
and U15173 (N_15173,N_14869,N_14930);
nor U15174 (N_15174,N_14908,N_14939);
and U15175 (N_15175,N_14847,N_14833);
and U15176 (N_15176,N_14842,N_14846);
nor U15177 (N_15177,N_14941,N_14930);
or U15178 (N_15178,N_14869,N_14975);
nand U15179 (N_15179,N_14881,N_14959);
nand U15180 (N_15180,N_14852,N_14841);
nor U15181 (N_15181,N_14828,N_14963);
xnor U15182 (N_15182,N_14841,N_14987);
nand U15183 (N_15183,N_14933,N_14969);
and U15184 (N_15184,N_14956,N_14889);
or U15185 (N_15185,N_14985,N_14801);
or U15186 (N_15186,N_14965,N_14818);
nor U15187 (N_15187,N_14985,N_14942);
nand U15188 (N_15188,N_14851,N_14928);
or U15189 (N_15189,N_14812,N_14960);
or U15190 (N_15190,N_14915,N_14889);
and U15191 (N_15191,N_14824,N_14922);
or U15192 (N_15192,N_14950,N_14866);
and U15193 (N_15193,N_14801,N_14891);
nand U15194 (N_15194,N_14980,N_14989);
nor U15195 (N_15195,N_14823,N_14932);
xnor U15196 (N_15196,N_14927,N_14803);
nand U15197 (N_15197,N_14983,N_14918);
xor U15198 (N_15198,N_14947,N_14869);
or U15199 (N_15199,N_14862,N_14967);
or U15200 (N_15200,N_15170,N_15019);
or U15201 (N_15201,N_15110,N_15142);
and U15202 (N_15202,N_15109,N_15063);
nand U15203 (N_15203,N_15197,N_15052);
nor U15204 (N_15204,N_15030,N_15140);
xnor U15205 (N_15205,N_15027,N_15047);
and U15206 (N_15206,N_15088,N_15022);
and U15207 (N_15207,N_15023,N_15137);
and U15208 (N_15208,N_15112,N_15134);
nor U15209 (N_15209,N_15072,N_15188);
and U15210 (N_15210,N_15059,N_15199);
or U15211 (N_15211,N_15163,N_15165);
xnor U15212 (N_15212,N_15120,N_15174);
xor U15213 (N_15213,N_15070,N_15107);
or U15214 (N_15214,N_15066,N_15103);
and U15215 (N_15215,N_15092,N_15003);
or U15216 (N_15216,N_15155,N_15051);
or U15217 (N_15217,N_15100,N_15099);
xor U15218 (N_15218,N_15039,N_15020);
nand U15219 (N_15219,N_15184,N_15021);
or U15220 (N_15220,N_15113,N_15074);
nor U15221 (N_15221,N_15016,N_15053);
nor U15222 (N_15222,N_15090,N_15015);
nand U15223 (N_15223,N_15156,N_15012);
and U15224 (N_15224,N_15196,N_15179);
xnor U15225 (N_15225,N_15175,N_15158);
or U15226 (N_15226,N_15093,N_15116);
or U15227 (N_15227,N_15044,N_15191);
xor U15228 (N_15228,N_15193,N_15118);
nor U15229 (N_15229,N_15075,N_15036);
nand U15230 (N_15230,N_15011,N_15106);
and U15231 (N_15231,N_15166,N_15041);
nand U15232 (N_15232,N_15058,N_15181);
nor U15233 (N_15233,N_15061,N_15128);
nand U15234 (N_15234,N_15117,N_15172);
or U15235 (N_15235,N_15190,N_15178);
or U15236 (N_15236,N_15055,N_15121);
nand U15237 (N_15237,N_15101,N_15152);
xor U15238 (N_15238,N_15133,N_15013);
nor U15239 (N_15239,N_15042,N_15160);
nor U15240 (N_15240,N_15162,N_15089);
xnor U15241 (N_15241,N_15000,N_15054);
nor U15242 (N_15242,N_15008,N_15138);
and U15243 (N_15243,N_15048,N_15076);
or U15244 (N_15244,N_15043,N_15168);
nor U15245 (N_15245,N_15146,N_15087);
xnor U15246 (N_15246,N_15176,N_15182);
or U15247 (N_15247,N_15071,N_15028);
nor U15248 (N_15248,N_15131,N_15010);
xnor U15249 (N_15249,N_15167,N_15198);
and U15250 (N_15250,N_15111,N_15035);
nand U15251 (N_15251,N_15119,N_15079);
nand U15252 (N_15252,N_15057,N_15145);
nand U15253 (N_15253,N_15129,N_15060);
and U15254 (N_15254,N_15122,N_15127);
nor U15255 (N_15255,N_15002,N_15144);
and U15256 (N_15256,N_15115,N_15132);
or U15257 (N_15257,N_15130,N_15154);
xor U15258 (N_15258,N_15045,N_15081);
nand U15259 (N_15259,N_15073,N_15091);
nand U15260 (N_15260,N_15067,N_15077);
xor U15261 (N_15261,N_15171,N_15046);
nor U15262 (N_15262,N_15147,N_15150);
nor U15263 (N_15263,N_15157,N_15148);
xor U15264 (N_15264,N_15114,N_15095);
nand U15265 (N_15265,N_15141,N_15124);
nor U15266 (N_15266,N_15040,N_15149);
and U15267 (N_15267,N_15136,N_15125);
and U15268 (N_15268,N_15031,N_15173);
xnor U15269 (N_15269,N_15104,N_15065);
xnor U15270 (N_15270,N_15084,N_15180);
nor U15271 (N_15271,N_15068,N_15062);
nor U15272 (N_15272,N_15082,N_15034);
nand U15273 (N_15273,N_15151,N_15183);
xnor U15274 (N_15274,N_15050,N_15018);
or U15275 (N_15275,N_15085,N_15161);
nand U15276 (N_15276,N_15126,N_15194);
xnor U15277 (N_15277,N_15164,N_15169);
or U15278 (N_15278,N_15096,N_15192);
and U15279 (N_15279,N_15009,N_15038);
nand U15280 (N_15280,N_15004,N_15105);
xor U15281 (N_15281,N_15185,N_15069);
nand U15282 (N_15282,N_15083,N_15187);
xnor U15283 (N_15283,N_15032,N_15049);
xor U15284 (N_15284,N_15123,N_15029);
or U15285 (N_15285,N_15195,N_15186);
nor U15286 (N_15286,N_15177,N_15005);
xnor U15287 (N_15287,N_15153,N_15086);
and U15288 (N_15288,N_15014,N_15080);
xor U15289 (N_15289,N_15026,N_15006);
nand U15290 (N_15290,N_15024,N_15135);
and U15291 (N_15291,N_15064,N_15033);
and U15292 (N_15292,N_15159,N_15001);
nor U15293 (N_15293,N_15143,N_15017);
nand U15294 (N_15294,N_15025,N_15102);
and U15295 (N_15295,N_15056,N_15037);
or U15296 (N_15296,N_15094,N_15098);
nor U15297 (N_15297,N_15078,N_15139);
xnor U15298 (N_15298,N_15108,N_15097);
nand U15299 (N_15299,N_15189,N_15007);
or U15300 (N_15300,N_15092,N_15040);
xnor U15301 (N_15301,N_15084,N_15098);
xnor U15302 (N_15302,N_15136,N_15074);
xnor U15303 (N_15303,N_15026,N_15043);
nand U15304 (N_15304,N_15101,N_15039);
nor U15305 (N_15305,N_15003,N_15150);
xor U15306 (N_15306,N_15167,N_15020);
nand U15307 (N_15307,N_15142,N_15140);
xnor U15308 (N_15308,N_15044,N_15179);
nor U15309 (N_15309,N_15090,N_15105);
xor U15310 (N_15310,N_15179,N_15066);
nor U15311 (N_15311,N_15069,N_15068);
or U15312 (N_15312,N_15003,N_15000);
xnor U15313 (N_15313,N_15099,N_15190);
nand U15314 (N_15314,N_15085,N_15032);
and U15315 (N_15315,N_15168,N_15152);
and U15316 (N_15316,N_15031,N_15102);
xnor U15317 (N_15317,N_15102,N_15128);
or U15318 (N_15318,N_15019,N_15067);
or U15319 (N_15319,N_15150,N_15030);
nor U15320 (N_15320,N_15184,N_15000);
nor U15321 (N_15321,N_15159,N_15144);
and U15322 (N_15322,N_15063,N_15191);
nor U15323 (N_15323,N_15094,N_15141);
and U15324 (N_15324,N_15091,N_15148);
nand U15325 (N_15325,N_15156,N_15120);
or U15326 (N_15326,N_15197,N_15063);
or U15327 (N_15327,N_15153,N_15171);
or U15328 (N_15328,N_15195,N_15158);
nand U15329 (N_15329,N_15035,N_15144);
or U15330 (N_15330,N_15130,N_15134);
or U15331 (N_15331,N_15080,N_15180);
xor U15332 (N_15332,N_15118,N_15013);
or U15333 (N_15333,N_15110,N_15020);
and U15334 (N_15334,N_15091,N_15160);
xor U15335 (N_15335,N_15010,N_15050);
or U15336 (N_15336,N_15046,N_15109);
nor U15337 (N_15337,N_15165,N_15159);
nor U15338 (N_15338,N_15049,N_15050);
nand U15339 (N_15339,N_15052,N_15037);
nand U15340 (N_15340,N_15119,N_15073);
nor U15341 (N_15341,N_15061,N_15043);
nor U15342 (N_15342,N_15056,N_15044);
or U15343 (N_15343,N_15115,N_15167);
or U15344 (N_15344,N_15065,N_15169);
nand U15345 (N_15345,N_15170,N_15146);
nand U15346 (N_15346,N_15055,N_15089);
xnor U15347 (N_15347,N_15036,N_15060);
or U15348 (N_15348,N_15130,N_15014);
nor U15349 (N_15349,N_15045,N_15086);
or U15350 (N_15350,N_15020,N_15139);
xor U15351 (N_15351,N_15172,N_15163);
or U15352 (N_15352,N_15055,N_15103);
xnor U15353 (N_15353,N_15083,N_15199);
and U15354 (N_15354,N_15132,N_15059);
nand U15355 (N_15355,N_15130,N_15149);
and U15356 (N_15356,N_15051,N_15142);
or U15357 (N_15357,N_15029,N_15004);
or U15358 (N_15358,N_15056,N_15153);
xor U15359 (N_15359,N_15001,N_15196);
or U15360 (N_15360,N_15179,N_15026);
xnor U15361 (N_15361,N_15060,N_15031);
or U15362 (N_15362,N_15054,N_15123);
or U15363 (N_15363,N_15067,N_15098);
nand U15364 (N_15364,N_15129,N_15080);
xor U15365 (N_15365,N_15005,N_15007);
or U15366 (N_15366,N_15196,N_15109);
or U15367 (N_15367,N_15084,N_15005);
nand U15368 (N_15368,N_15106,N_15120);
or U15369 (N_15369,N_15015,N_15166);
xor U15370 (N_15370,N_15065,N_15010);
nor U15371 (N_15371,N_15199,N_15167);
or U15372 (N_15372,N_15062,N_15063);
nor U15373 (N_15373,N_15137,N_15026);
and U15374 (N_15374,N_15136,N_15111);
or U15375 (N_15375,N_15058,N_15021);
nor U15376 (N_15376,N_15001,N_15145);
nor U15377 (N_15377,N_15121,N_15109);
nand U15378 (N_15378,N_15192,N_15029);
nand U15379 (N_15379,N_15183,N_15077);
xnor U15380 (N_15380,N_15073,N_15063);
or U15381 (N_15381,N_15177,N_15129);
or U15382 (N_15382,N_15180,N_15149);
nand U15383 (N_15383,N_15124,N_15024);
nand U15384 (N_15384,N_15141,N_15097);
nand U15385 (N_15385,N_15088,N_15025);
nor U15386 (N_15386,N_15154,N_15085);
xnor U15387 (N_15387,N_15051,N_15112);
xnor U15388 (N_15388,N_15036,N_15178);
nand U15389 (N_15389,N_15006,N_15104);
nor U15390 (N_15390,N_15090,N_15185);
nand U15391 (N_15391,N_15052,N_15103);
and U15392 (N_15392,N_15061,N_15052);
nand U15393 (N_15393,N_15159,N_15077);
nor U15394 (N_15394,N_15183,N_15026);
nor U15395 (N_15395,N_15077,N_15143);
and U15396 (N_15396,N_15067,N_15102);
or U15397 (N_15397,N_15016,N_15146);
or U15398 (N_15398,N_15007,N_15112);
nand U15399 (N_15399,N_15105,N_15054);
and U15400 (N_15400,N_15229,N_15212);
xor U15401 (N_15401,N_15386,N_15323);
nand U15402 (N_15402,N_15363,N_15217);
xnor U15403 (N_15403,N_15384,N_15326);
xnor U15404 (N_15404,N_15367,N_15218);
nand U15405 (N_15405,N_15224,N_15279);
xnor U15406 (N_15406,N_15364,N_15298);
and U15407 (N_15407,N_15357,N_15373);
or U15408 (N_15408,N_15230,N_15377);
nor U15409 (N_15409,N_15390,N_15392);
or U15410 (N_15410,N_15352,N_15330);
xor U15411 (N_15411,N_15382,N_15374);
nor U15412 (N_15412,N_15248,N_15278);
or U15413 (N_15413,N_15255,N_15341);
or U15414 (N_15414,N_15308,N_15253);
nor U15415 (N_15415,N_15245,N_15237);
xor U15416 (N_15416,N_15287,N_15295);
nand U15417 (N_15417,N_15397,N_15360);
and U15418 (N_15418,N_15284,N_15346);
xnor U15419 (N_15419,N_15370,N_15344);
and U15420 (N_15420,N_15203,N_15399);
nor U15421 (N_15421,N_15291,N_15316);
and U15422 (N_15422,N_15236,N_15281);
nor U15423 (N_15423,N_15283,N_15350);
and U15424 (N_15424,N_15368,N_15322);
xnor U15425 (N_15425,N_15312,N_15396);
nand U15426 (N_15426,N_15294,N_15301);
nand U15427 (N_15427,N_15307,N_15302);
nand U15428 (N_15428,N_15246,N_15223);
nand U15429 (N_15429,N_15336,N_15338);
nand U15430 (N_15430,N_15268,N_15208);
and U15431 (N_15431,N_15258,N_15369);
nand U15432 (N_15432,N_15226,N_15297);
or U15433 (N_15433,N_15269,N_15277);
xnor U15434 (N_15434,N_15242,N_15264);
and U15435 (N_15435,N_15398,N_15347);
nor U15436 (N_15436,N_15228,N_15262);
and U15437 (N_15437,N_15249,N_15211);
nor U15438 (N_15438,N_15285,N_15356);
or U15439 (N_15439,N_15256,N_15250);
xor U15440 (N_15440,N_15328,N_15247);
nor U15441 (N_15441,N_15270,N_15342);
xnor U15442 (N_15442,N_15310,N_15251);
xnor U15443 (N_15443,N_15381,N_15355);
and U15444 (N_15444,N_15309,N_15303);
xor U15445 (N_15445,N_15319,N_15235);
nor U15446 (N_15446,N_15239,N_15379);
nor U15447 (N_15447,N_15361,N_15266);
xnor U15448 (N_15448,N_15257,N_15314);
and U15449 (N_15449,N_15315,N_15339);
xnor U15450 (N_15450,N_15371,N_15219);
xnor U15451 (N_15451,N_15206,N_15231);
or U15452 (N_15452,N_15221,N_15387);
xnor U15453 (N_15453,N_15252,N_15207);
xor U15454 (N_15454,N_15343,N_15271);
or U15455 (N_15455,N_15289,N_15380);
nor U15456 (N_15456,N_15359,N_15273);
nor U15457 (N_15457,N_15225,N_15227);
and U15458 (N_15458,N_15332,N_15276);
and U15459 (N_15459,N_15337,N_15378);
nor U15460 (N_15460,N_15331,N_15304);
or U15461 (N_15461,N_15299,N_15259);
or U15462 (N_15462,N_15317,N_15324);
xor U15463 (N_15463,N_15274,N_15202);
and U15464 (N_15464,N_15348,N_15376);
and U15465 (N_15465,N_15290,N_15366);
and U15466 (N_15466,N_15267,N_15325);
xor U15467 (N_15467,N_15389,N_15209);
nor U15468 (N_15468,N_15313,N_15234);
or U15469 (N_15469,N_15254,N_15393);
and U15470 (N_15470,N_15300,N_15210);
and U15471 (N_15471,N_15349,N_15244);
xor U15472 (N_15472,N_15306,N_15201);
or U15473 (N_15473,N_15220,N_15305);
xnor U15474 (N_15474,N_15334,N_15385);
or U15475 (N_15475,N_15205,N_15200);
xor U15476 (N_15476,N_15265,N_15272);
and U15477 (N_15477,N_15329,N_15240);
and U15478 (N_15478,N_15280,N_15375);
nor U15479 (N_15479,N_15288,N_15320);
and U15480 (N_15480,N_15362,N_15232);
xnor U15481 (N_15481,N_15353,N_15275);
nor U15482 (N_15482,N_15213,N_15215);
or U15483 (N_15483,N_15394,N_15383);
nor U15484 (N_15484,N_15318,N_15261);
nand U15485 (N_15485,N_15327,N_15351);
xor U15486 (N_15486,N_15293,N_15358);
nand U15487 (N_15487,N_15311,N_15372);
nor U15488 (N_15488,N_15243,N_15391);
xor U15489 (N_15489,N_15241,N_15233);
and U15490 (N_15490,N_15388,N_15214);
and U15491 (N_15491,N_15222,N_15292);
nor U15492 (N_15492,N_15340,N_15263);
and U15493 (N_15493,N_15204,N_15296);
xnor U15494 (N_15494,N_15238,N_15333);
nand U15495 (N_15495,N_15395,N_15354);
nand U15496 (N_15496,N_15335,N_15365);
or U15497 (N_15497,N_15260,N_15286);
or U15498 (N_15498,N_15216,N_15345);
or U15499 (N_15499,N_15282,N_15321);
nor U15500 (N_15500,N_15231,N_15326);
xnor U15501 (N_15501,N_15287,N_15368);
xor U15502 (N_15502,N_15382,N_15310);
or U15503 (N_15503,N_15334,N_15328);
nor U15504 (N_15504,N_15356,N_15277);
and U15505 (N_15505,N_15233,N_15318);
or U15506 (N_15506,N_15222,N_15340);
and U15507 (N_15507,N_15262,N_15378);
nor U15508 (N_15508,N_15318,N_15292);
xnor U15509 (N_15509,N_15300,N_15272);
and U15510 (N_15510,N_15335,N_15258);
or U15511 (N_15511,N_15362,N_15271);
and U15512 (N_15512,N_15398,N_15200);
nor U15513 (N_15513,N_15269,N_15298);
xor U15514 (N_15514,N_15383,N_15399);
xor U15515 (N_15515,N_15257,N_15325);
nor U15516 (N_15516,N_15278,N_15219);
nor U15517 (N_15517,N_15276,N_15396);
or U15518 (N_15518,N_15306,N_15267);
xor U15519 (N_15519,N_15278,N_15271);
nand U15520 (N_15520,N_15392,N_15209);
xor U15521 (N_15521,N_15243,N_15397);
or U15522 (N_15522,N_15203,N_15225);
or U15523 (N_15523,N_15335,N_15227);
nand U15524 (N_15524,N_15389,N_15335);
and U15525 (N_15525,N_15233,N_15243);
xor U15526 (N_15526,N_15344,N_15271);
and U15527 (N_15527,N_15329,N_15226);
xor U15528 (N_15528,N_15296,N_15241);
nor U15529 (N_15529,N_15317,N_15282);
and U15530 (N_15530,N_15275,N_15311);
nand U15531 (N_15531,N_15315,N_15344);
and U15532 (N_15532,N_15221,N_15365);
or U15533 (N_15533,N_15260,N_15372);
or U15534 (N_15534,N_15280,N_15350);
xor U15535 (N_15535,N_15244,N_15250);
nor U15536 (N_15536,N_15237,N_15256);
nand U15537 (N_15537,N_15294,N_15206);
xnor U15538 (N_15538,N_15255,N_15376);
nor U15539 (N_15539,N_15202,N_15281);
nor U15540 (N_15540,N_15247,N_15310);
nand U15541 (N_15541,N_15366,N_15339);
and U15542 (N_15542,N_15266,N_15321);
xnor U15543 (N_15543,N_15208,N_15352);
xor U15544 (N_15544,N_15370,N_15233);
and U15545 (N_15545,N_15343,N_15288);
nand U15546 (N_15546,N_15307,N_15350);
nand U15547 (N_15547,N_15309,N_15254);
nor U15548 (N_15548,N_15246,N_15304);
or U15549 (N_15549,N_15207,N_15258);
nand U15550 (N_15550,N_15231,N_15214);
nand U15551 (N_15551,N_15323,N_15367);
nor U15552 (N_15552,N_15319,N_15329);
or U15553 (N_15553,N_15397,N_15258);
nand U15554 (N_15554,N_15219,N_15314);
nor U15555 (N_15555,N_15336,N_15237);
and U15556 (N_15556,N_15299,N_15372);
and U15557 (N_15557,N_15339,N_15301);
and U15558 (N_15558,N_15363,N_15399);
and U15559 (N_15559,N_15278,N_15221);
nor U15560 (N_15560,N_15279,N_15238);
or U15561 (N_15561,N_15321,N_15261);
and U15562 (N_15562,N_15259,N_15258);
or U15563 (N_15563,N_15280,N_15246);
nor U15564 (N_15564,N_15230,N_15235);
nor U15565 (N_15565,N_15246,N_15342);
and U15566 (N_15566,N_15367,N_15330);
xor U15567 (N_15567,N_15254,N_15370);
nor U15568 (N_15568,N_15293,N_15225);
xor U15569 (N_15569,N_15273,N_15348);
nand U15570 (N_15570,N_15292,N_15201);
nor U15571 (N_15571,N_15243,N_15205);
and U15572 (N_15572,N_15284,N_15368);
nor U15573 (N_15573,N_15358,N_15226);
nor U15574 (N_15574,N_15397,N_15280);
or U15575 (N_15575,N_15244,N_15293);
and U15576 (N_15576,N_15339,N_15227);
and U15577 (N_15577,N_15211,N_15355);
xor U15578 (N_15578,N_15398,N_15266);
xor U15579 (N_15579,N_15304,N_15295);
or U15580 (N_15580,N_15263,N_15328);
nor U15581 (N_15581,N_15262,N_15270);
nor U15582 (N_15582,N_15313,N_15360);
and U15583 (N_15583,N_15261,N_15395);
nor U15584 (N_15584,N_15234,N_15381);
nand U15585 (N_15585,N_15303,N_15250);
xnor U15586 (N_15586,N_15382,N_15207);
nor U15587 (N_15587,N_15257,N_15315);
nand U15588 (N_15588,N_15308,N_15292);
nand U15589 (N_15589,N_15392,N_15372);
nor U15590 (N_15590,N_15393,N_15224);
xor U15591 (N_15591,N_15233,N_15258);
xor U15592 (N_15592,N_15315,N_15290);
or U15593 (N_15593,N_15304,N_15334);
xnor U15594 (N_15594,N_15377,N_15340);
or U15595 (N_15595,N_15280,N_15364);
and U15596 (N_15596,N_15260,N_15205);
nand U15597 (N_15597,N_15294,N_15320);
nor U15598 (N_15598,N_15362,N_15370);
nor U15599 (N_15599,N_15325,N_15252);
nand U15600 (N_15600,N_15560,N_15455);
or U15601 (N_15601,N_15512,N_15553);
nor U15602 (N_15602,N_15400,N_15456);
xnor U15603 (N_15603,N_15579,N_15569);
nor U15604 (N_15604,N_15424,N_15416);
nor U15605 (N_15605,N_15449,N_15502);
or U15606 (N_15606,N_15493,N_15530);
nand U15607 (N_15607,N_15529,N_15482);
or U15608 (N_15608,N_15419,N_15426);
and U15609 (N_15609,N_15459,N_15490);
or U15610 (N_15610,N_15511,N_15433);
or U15611 (N_15611,N_15495,N_15436);
nand U15612 (N_15612,N_15581,N_15578);
xor U15613 (N_15613,N_15427,N_15582);
nand U15614 (N_15614,N_15531,N_15498);
nand U15615 (N_15615,N_15404,N_15527);
and U15616 (N_15616,N_15516,N_15522);
nand U15617 (N_15617,N_15478,N_15407);
nand U15618 (N_15618,N_15559,N_15472);
nor U15619 (N_15619,N_15470,N_15571);
or U15620 (N_15620,N_15585,N_15491);
xor U15621 (N_15621,N_15451,N_15519);
nand U15622 (N_15622,N_15570,N_15575);
or U15623 (N_15623,N_15467,N_15486);
and U15624 (N_15624,N_15515,N_15461);
or U15625 (N_15625,N_15437,N_15454);
nor U15626 (N_15626,N_15580,N_15558);
xnor U15627 (N_15627,N_15548,N_15521);
nor U15628 (N_15628,N_15588,N_15457);
nand U15629 (N_15629,N_15532,N_15441);
nand U15630 (N_15630,N_15450,N_15574);
xnor U15631 (N_15631,N_15566,N_15576);
xor U15632 (N_15632,N_15541,N_15497);
and U15633 (N_15633,N_15465,N_15425);
and U15634 (N_15634,N_15520,N_15410);
nand U15635 (N_15635,N_15483,N_15460);
nand U15636 (N_15636,N_15492,N_15594);
nand U15637 (N_15637,N_15434,N_15533);
nand U15638 (N_15638,N_15438,N_15552);
or U15639 (N_15639,N_15535,N_15453);
nor U15640 (N_15640,N_15543,N_15408);
and U15641 (N_15641,N_15444,N_15406);
xnor U15642 (N_15642,N_15513,N_15431);
nand U15643 (N_15643,N_15510,N_15485);
nor U15644 (N_15644,N_15555,N_15557);
nand U15645 (N_15645,N_15432,N_15471);
xor U15646 (N_15646,N_15489,N_15468);
xor U15647 (N_15647,N_15411,N_15445);
or U15648 (N_15648,N_15554,N_15443);
or U15649 (N_15649,N_15479,N_15561);
xor U15650 (N_15650,N_15429,N_15415);
and U15651 (N_15651,N_15423,N_15544);
or U15652 (N_15652,N_15549,N_15583);
or U15653 (N_15653,N_15592,N_15573);
xor U15654 (N_15654,N_15568,N_15525);
xnor U15655 (N_15655,N_15420,N_15589);
xnor U15656 (N_15656,N_15538,N_15517);
nand U15657 (N_15657,N_15542,N_15442);
nand U15658 (N_15658,N_15546,N_15545);
or U15659 (N_15659,N_15524,N_15440);
nand U15660 (N_15660,N_15547,N_15473);
nor U15661 (N_15661,N_15403,N_15550);
nor U15662 (N_15662,N_15508,N_15556);
or U15663 (N_15663,N_15474,N_15500);
xnor U15664 (N_15664,N_15480,N_15452);
or U15665 (N_15665,N_15476,N_15540);
and U15666 (N_15666,N_15439,N_15597);
and U15667 (N_15667,N_15430,N_15598);
and U15668 (N_15668,N_15428,N_15496);
xnor U15669 (N_15669,N_15596,N_15477);
nand U15670 (N_15670,N_15593,N_15528);
or U15671 (N_15671,N_15504,N_15447);
and U15672 (N_15672,N_15501,N_15494);
and U15673 (N_15673,N_15507,N_15536);
and U15674 (N_15674,N_15462,N_15551);
or U15675 (N_15675,N_15421,N_15503);
nor U15676 (N_15676,N_15417,N_15402);
nand U15677 (N_15677,N_15475,N_15401);
xor U15678 (N_15678,N_15506,N_15572);
xnor U15679 (N_15679,N_15564,N_15405);
and U15680 (N_15680,N_15488,N_15469);
xor U15681 (N_15681,N_15487,N_15565);
or U15682 (N_15682,N_15563,N_15458);
or U15683 (N_15683,N_15418,N_15481);
xnor U15684 (N_15684,N_15584,N_15586);
nor U15685 (N_15685,N_15448,N_15414);
xnor U15686 (N_15686,N_15413,N_15422);
xnor U15687 (N_15687,N_15446,N_15539);
nor U15688 (N_15688,N_15587,N_15412);
nor U15689 (N_15689,N_15526,N_15537);
nor U15690 (N_15690,N_15577,N_15463);
or U15691 (N_15691,N_15523,N_15499);
or U15692 (N_15692,N_15595,N_15534);
and U15693 (N_15693,N_15509,N_15505);
nor U15694 (N_15694,N_15562,N_15466);
or U15695 (N_15695,N_15518,N_15409);
or U15696 (N_15696,N_15464,N_15484);
and U15697 (N_15697,N_15591,N_15590);
xor U15698 (N_15698,N_15567,N_15435);
xnor U15699 (N_15699,N_15599,N_15514);
nor U15700 (N_15700,N_15461,N_15403);
and U15701 (N_15701,N_15546,N_15493);
or U15702 (N_15702,N_15466,N_15515);
and U15703 (N_15703,N_15415,N_15568);
xor U15704 (N_15704,N_15434,N_15475);
and U15705 (N_15705,N_15511,N_15538);
nor U15706 (N_15706,N_15480,N_15532);
and U15707 (N_15707,N_15480,N_15570);
xor U15708 (N_15708,N_15464,N_15445);
nand U15709 (N_15709,N_15425,N_15458);
xor U15710 (N_15710,N_15572,N_15403);
or U15711 (N_15711,N_15484,N_15493);
xor U15712 (N_15712,N_15422,N_15489);
and U15713 (N_15713,N_15425,N_15483);
nor U15714 (N_15714,N_15572,N_15526);
and U15715 (N_15715,N_15454,N_15547);
or U15716 (N_15716,N_15452,N_15506);
and U15717 (N_15717,N_15529,N_15525);
or U15718 (N_15718,N_15424,N_15474);
or U15719 (N_15719,N_15451,N_15508);
or U15720 (N_15720,N_15534,N_15416);
nand U15721 (N_15721,N_15545,N_15477);
or U15722 (N_15722,N_15494,N_15542);
nor U15723 (N_15723,N_15508,N_15541);
and U15724 (N_15724,N_15594,N_15579);
nand U15725 (N_15725,N_15579,N_15599);
and U15726 (N_15726,N_15511,N_15524);
nand U15727 (N_15727,N_15413,N_15580);
xor U15728 (N_15728,N_15483,N_15519);
xnor U15729 (N_15729,N_15460,N_15502);
nand U15730 (N_15730,N_15443,N_15424);
xnor U15731 (N_15731,N_15597,N_15590);
or U15732 (N_15732,N_15598,N_15418);
nand U15733 (N_15733,N_15416,N_15430);
xnor U15734 (N_15734,N_15540,N_15595);
nor U15735 (N_15735,N_15438,N_15509);
nand U15736 (N_15736,N_15529,N_15522);
xnor U15737 (N_15737,N_15574,N_15456);
nand U15738 (N_15738,N_15507,N_15418);
or U15739 (N_15739,N_15578,N_15549);
or U15740 (N_15740,N_15456,N_15409);
xnor U15741 (N_15741,N_15556,N_15473);
or U15742 (N_15742,N_15474,N_15579);
or U15743 (N_15743,N_15453,N_15532);
nor U15744 (N_15744,N_15499,N_15406);
xor U15745 (N_15745,N_15418,N_15531);
and U15746 (N_15746,N_15415,N_15580);
or U15747 (N_15747,N_15527,N_15542);
or U15748 (N_15748,N_15548,N_15435);
or U15749 (N_15749,N_15559,N_15534);
or U15750 (N_15750,N_15569,N_15462);
and U15751 (N_15751,N_15561,N_15419);
nor U15752 (N_15752,N_15490,N_15528);
xnor U15753 (N_15753,N_15527,N_15410);
xnor U15754 (N_15754,N_15419,N_15498);
nand U15755 (N_15755,N_15548,N_15426);
nand U15756 (N_15756,N_15419,N_15432);
and U15757 (N_15757,N_15550,N_15475);
and U15758 (N_15758,N_15426,N_15405);
nor U15759 (N_15759,N_15505,N_15451);
xnor U15760 (N_15760,N_15503,N_15490);
or U15761 (N_15761,N_15524,N_15536);
and U15762 (N_15762,N_15552,N_15529);
xnor U15763 (N_15763,N_15593,N_15595);
or U15764 (N_15764,N_15507,N_15484);
nand U15765 (N_15765,N_15531,N_15448);
nor U15766 (N_15766,N_15575,N_15511);
xor U15767 (N_15767,N_15577,N_15495);
and U15768 (N_15768,N_15579,N_15446);
xnor U15769 (N_15769,N_15476,N_15524);
xnor U15770 (N_15770,N_15564,N_15569);
xor U15771 (N_15771,N_15424,N_15558);
or U15772 (N_15772,N_15584,N_15589);
and U15773 (N_15773,N_15593,N_15432);
nand U15774 (N_15774,N_15478,N_15450);
and U15775 (N_15775,N_15450,N_15429);
nor U15776 (N_15776,N_15417,N_15565);
and U15777 (N_15777,N_15483,N_15445);
and U15778 (N_15778,N_15457,N_15533);
and U15779 (N_15779,N_15401,N_15491);
nand U15780 (N_15780,N_15471,N_15586);
or U15781 (N_15781,N_15406,N_15584);
and U15782 (N_15782,N_15524,N_15456);
xor U15783 (N_15783,N_15532,N_15589);
nand U15784 (N_15784,N_15450,N_15498);
nor U15785 (N_15785,N_15595,N_15424);
nand U15786 (N_15786,N_15468,N_15511);
xnor U15787 (N_15787,N_15452,N_15456);
xor U15788 (N_15788,N_15512,N_15527);
nand U15789 (N_15789,N_15446,N_15417);
or U15790 (N_15790,N_15588,N_15470);
xor U15791 (N_15791,N_15426,N_15587);
or U15792 (N_15792,N_15582,N_15416);
nand U15793 (N_15793,N_15479,N_15508);
nand U15794 (N_15794,N_15409,N_15543);
or U15795 (N_15795,N_15510,N_15443);
nor U15796 (N_15796,N_15433,N_15534);
xnor U15797 (N_15797,N_15547,N_15478);
nor U15798 (N_15798,N_15518,N_15584);
xor U15799 (N_15799,N_15462,N_15505);
nor U15800 (N_15800,N_15712,N_15633);
xor U15801 (N_15801,N_15685,N_15619);
and U15802 (N_15802,N_15665,N_15602);
xor U15803 (N_15803,N_15744,N_15770);
xor U15804 (N_15804,N_15773,N_15715);
nor U15805 (N_15805,N_15664,N_15796);
or U15806 (N_15806,N_15655,N_15640);
nand U15807 (N_15807,N_15694,N_15720);
or U15808 (N_15808,N_15647,N_15784);
and U15809 (N_15809,N_15684,N_15696);
nor U15810 (N_15810,N_15794,N_15658);
and U15811 (N_15811,N_15753,N_15624);
nand U15812 (N_15812,N_15682,N_15700);
nor U15813 (N_15813,N_15644,N_15754);
and U15814 (N_15814,N_15738,N_15785);
and U15815 (N_15815,N_15673,N_15764);
nor U15816 (N_15816,N_15639,N_15630);
xnor U15817 (N_15817,N_15675,N_15710);
nor U15818 (N_15818,N_15618,N_15615);
nand U15819 (N_15819,N_15637,N_15656);
or U15820 (N_15820,N_15654,N_15726);
nand U15821 (N_15821,N_15628,N_15760);
xnor U15822 (N_15822,N_15670,N_15740);
nand U15823 (N_15823,N_15689,N_15652);
or U15824 (N_15824,N_15632,N_15739);
or U15825 (N_15825,N_15677,N_15612);
xnor U15826 (N_15826,N_15613,N_15716);
and U15827 (N_15827,N_15638,N_15749);
or U15828 (N_15828,N_15728,N_15713);
xnor U15829 (N_15829,N_15606,N_15707);
or U15830 (N_15830,N_15705,N_15769);
or U15831 (N_15831,N_15798,N_15610);
or U15832 (N_15832,N_15625,N_15787);
or U15833 (N_15833,N_15724,N_15741);
and U15834 (N_15834,N_15751,N_15695);
or U15835 (N_15835,N_15631,N_15708);
xor U15836 (N_15836,N_15605,N_15608);
nand U15837 (N_15837,N_15737,N_15663);
and U15838 (N_15838,N_15763,N_15641);
nand U15839 (N_15839,N_15635,N_15697);
nor U15840 (N_15840,N_15748,N_15681);
and U15841 (N_15841,N_15761,N_15725);
xnor U15842 (N_15842,N_15723,N_15603);
and U15843 (N_15843,N_15623,N_15793);
nand U15844 (N_15844,N_15674,N_15776);
and U15845 (N_15845,N_15733,N_15651);
and U15846 (N_15846,N_15686,N_15750);
xnor U15847 (N_15847,N_15780,N_15621);
xnor U15848 (N_15848,N_15722,N_15601);
and U15849 (N_15849,N_15693,N_15611);
or U15850 (N_15850,N_15718,N_15777);
or U15851 (N_15851,N_15704,N_15795);
and U15852 (N_15852,N_15735,N_15616);
nand U15853 (N_15853,N_15600,N_15775);
xor U15854 (N_15854,N_15634,N_15701);
nand U15855 (N_15855,N_15755,N_15756);
and U15856 (N_15856,N_15782,N_15702);
or U15857 (N_15857,N_15669,N_15699);
nor U15858 (N_15858,N_15709,N_15779);
or U15859 (N_15859,N_15786,N_15768);
or U15860 (N_15860,N_15730,N_15729);
nor U15861 (N_15861,N_15711,N_15643);
nor U15862 (N_15862,N_15609,N_15736);
nand U15863 (N_15863,N_15672,N_15745);
or U15864 (N_15864,N_15648,N_15752);
xnor U15865 (N_15865,N_15683,N_15662);
nand U15866 (N_15866,N_15771,N_15614);
xor U15867 (N_15867,N_15774,N_15690);
and U15868 (N_15868,N_15671,N_15783);
nor U15869 (N_15869,N_15646,N_15692);
and U15870 (N_15870,N_15679,N_15667);
xor U15871 (N_15871,N_15765,N_15680);
nand U15872 (N_15872,N_15742,N_15649);
and U15873 (N_15873,N_15691,N_15719);
or U15874 (N_15874,N_15792,N_15627);
and U15875 (N_15875,N_15698,N_15688);
xor U15876 (N_15876,N_15636,N_15687);
xnor U15877 (N_15877,N_15799,N_15660);
and U15878 (N_15878,N_15620,N_15789);
and U15879 (N_15879,N_15790,N_15617);
xor U15880 (N_15880,N_15746,N_15767);
xor U15881 (N_15881,N_15759,N_15743);
and U15882 (N_15882,N_15781,N_15659);
and U15883 (N_15883,N_15778,N_15731);
nand U15884 (N_15884,N_15714,N_15653);
and U15885 (N_15885,N_15747,N_15668);
and U15886 (N_15886,N_15629,N_15706);
or U15887 (N_15887,N_15734,N_15642);
and U15888 (N_15888,N_15666,N_15604);
nand U15889 (N_15889,N_15622,N_15650);
nor U15890 (N_15890,N_15661,N_15766);
nor U15891 (N_15891,N_15758,N_15732);
nor U15892 (N_15892,N_15762,N_15607);
nand U15893 (N_15893,N_15717,N_15727);
xor U15894 (N_15894,N_15703,N_15797);
nand U15895 (N_15895,N_15721,N_15626);
nand U15896 (N_15896,N_15676,N_15757);
or U15897 (N_15897,N_15772,N_15645);
nand U15898 (N_15898,N_15788,N_15791);
xnor U15899 (N_15899,N_15657,N_15678);
xor U15900 (N_15900,N_15721,N_15633);
and U15901 (N_15901,N_15647,N_15648);
and U15902 (N_15902,N_15648,N_15715);
or U15903 (N_15903,N_15796,N_15729);
nand U15904 (N_15904,N_15796,N_15763);
nor U15905 (N_15905,N_15792,N_15685);
nor U15906 (N_15906,N_15759,N_15756);
or U15907 (N_15907,N_15711,N_15772);
or U15908 (N_15908,N_15725,N_15673);
or U15909 (N_15909,N_15689,N_15609);
or U15910 (N_15910,N_15751,N_15705);
nand U15911 (N_15911,N_15737,N_15791);
nor U15912 (N_15912,N_15678,N_15734);
and U15913 (N_15913,N_15615,N_15772);
nor U15914 (N_15914,N_15705,N_15771);
xnor U15915 (N_15915,N_15675,N_15643);
nand U15916 (N_15916,N_15697,N_15791);
or U15917 (N_15917,N_15694,N_15741);
nor U15918 (N_15918,N_15725,N_15764);
or U15919 (N_15919,N_15797,N_15679);
or U15920 (N_15920,N_15675,N_15770);
nor U15921 (N_15921,N_15749,N_15681);
and U15922 (N_15922,N_15781,N_15778);
or U15923 (N_15923,N_15725,N_15707);
nand U15924 (N_15924,N_15753,N_15639);
nand U15925 (N_15925,N_15730,N_15614);
nor U15926 (N_15926,N_15729,N_15768);
nor U15927 (N_15927,N_15748,N_15764);
and U15928 (N_15928,N_15641,N_15734);
and U15929 (N_15929,N_15788,N_15798);
nor U15930 (N_15930,N_15638,N_15609);
and U15931 (N_15931,N_15614,N_15622);
nor U15932 (N_15932,N_15639,N_15688);
and U15933 (N_15933,N_15771,N_15673);
nor U15934 (N_15934,N_15683,N_15745);
or U15935 (N_15935,N_15678,N_15768);
nor U15936 (N_15936,N_15755,N_15784);
nor U15937 (N_15937,N_15715,N_15788);
nor U15938 (N_15938,N_15749,N_15675);
nand U15939 (N_15939,N_15664,N_15702);
nor U15940 (N_15940,N_15732,N_15606);
xor U15941 (N_15941,N_15779,N_15730);
nand U15942 (N_15942,N_15730,N_15667);
xnor U15943 (N_15943,N_15761,N_15730);
and U15944 (N_15944,N_15799,N_15680);
and U15945 (N_15945,N_15775,N_15686);
and U15946 (N_15946,N_15745,N_15772);
xnor U15947 (N_15947,N_15787,N_15674);
nor U15948 (N_15948,N_15627,N_15794);
and U15949 (N_15949,N_15601,N_15672);
nand U15950 (N_15950,N_15797,N_15620);
nor U15951 (N_15951,N_15604,N_15709);
nor U15952 (N_15952,N_15622,N_15652);
nand U15953 (N_15953,N_15614,N_15729);
nor U15954 (N_15954,N_15608,N_15629);
nand U15955 (N_15955,N_15767,N_15764);
nand U15956 (N_15956,N_15688,N_15701);
or U15957 (N_15957,N_15625,N_15756);
xnor U15958 (N_15958,N_15604,N_15694);
and U15959 (N_15959,N_15601,N_15762);
and U15960 (N_15960,N_15709,N_15637);
or U15961 (N_15961,N_15684,N_15767);
nand U15962 (N_15962,N_15748,N_15635);
nor U15963 (N_15963,N_15710,N_15618);
and U15964 (N_15964,N_15764,N_15688);
and U15965 (N_15965,N_15617,N_15685);
or U15966 (N_15966,N_15714,N_15636);
and U15967 (N_15967,N_15637,N_15739);
nor U15968 (N_15968,N_15731,N_15759);
nor U15969 (N_15969,N_15624,N_15629);
and U15970 (N_15970,N_15724,N_15701);
xnor U15971 (N_15971,N_15636,N_15779);
and U15972 (N_15972,N_15747,N_15670);
nand U15973 (N_15973,N_15664,N_15691);
and U15974 (N_15974,N_15610,N_15667);
xnor U15975 (N_15975,N_15679,N_15632);
xor U15976 (N_15976,N_15626,N_15718);
xnor U15977 (N_15977,N_15739,N_15772);
nand U15978 (N_15978,N_15681,N_15703);
and U15979 (N_15979,N_15787,N_15733);
and U15980 (N_15980,N_15611,N_15601);
xnor U15981 (N_15981,N_15792,N_15760);
nand U15982 (N_15982,N_15773,N_15675);
nor U15983 (N_15983,N_15670,N_15648);
or U15984 (N_15984,N_15757,N_15692);
nor U15985 (N_15985,N_15769,N_15683);
and U15986 (N_15986,N_15623,N_15736);
and U15987 (N_15987,N_15659,N_15690);
nor U15988 (N_15988,N_15767,N_15662);
nand U15989 (N_15989,N_15798,N_15694);
and U15990 (N_15990,N_15685,N_15689);
nor U15991 (N_15991,N_15650,N_15748);
or U15992 (N_15992,N_15773,N_15749);
or U15993 (N_15993,N_15700,N_15633);
xor U15994 (N_15994,N_15737,N_15627);
xnor U15995 (N_15995,N_15661,N_15703);
and U15996 (N_15996,N_15746,N_15634);
nand U15997 (N_15997,N_15649,N_15646);
nand U15998 (N_15998,N_15741,N_15791);
xnor U15999 (N_15999,N_15777,N_15696);
and U16000 (N_16000,N_15830,N_15837);
xnor U16001 (N_16001,N_15907,N_15871);
nand U16002 (N_16002,N_15923,N_15851);
and U16003 (N_16003,N_15939,N_15865);
or U16004 (N_16004,N_15850,N_15960);
xnor U16005 (N_16005,N_15818,N_15946);
and U16006 (N_16006,N_15944,N_15981);
or U16007 (N_16007,N_15872,N_15812);
nor U16008 (N_16008,N_15930,N_15902);
or U16009 (N_16009,N_15969,N_15876);
and U16010 (N_16010,N_15973,N_15974);
or U16011 (N_16011,N_15994,N_15880);
xor U16012 (N_16012,N_15950,N_15942);
nor U16013 (N_16013,N_15893,N_15881);
or U16014 (N_16014,N_15966,N_15977);
xor U16015 (N_16015,N_15829,N_15801);
xor U16016 (N_16016,N_15873,N_15862);
nand U16017 (N_16017,N_15932,N_15962);
nand U16018 (N_16018,N_15856,N_15898);
nor U16019 (N_16019,N_15916,N_15903);
nor U16020 (N_16020,N_15941,N_15938);
nor U16021 (N_16021,N_15984,N_15913);
nand U16022 (N_16022,N_15885,N_15918);
xnor U16023 (N_16023,N_15852,N_15847);
xor U16024 (N_16024,N_15816,N_15956);
and U16025 (N_16025,N_15925,N_15912);
or U16026 (N_16026,N_15919,N_15922);
and U16027 (N_16027,N_15814,N_15874);
nand U16028 (N_16028,N_15866,N_15965);
xor U16029 (N_16029,N_15943,N_15935);
and U16030 (N_16030,N_15905,N_15979);
nand U16031 (N_16031,N_15917,N_15858);
xor U16032 (N_16032,N_15955,N_15890);
and U16033 (N_16033,N_15998,N_15929);
and U16034 (N_16034,N_15958,N_15800);
xor U16035 (N_16035,N_15824,N_15968);
xnor U16036 (N_16036,N_15883,N_15914);
or U16037 (N_16037,N_15805,N_15831);
nor U16038 (N_16038,N_15864,N_15859);
and U16039 (N_16039,N_15803,N_15886);
and U16040 (N_16040,N_15843,N_15853);
nor U16041 (N_16041,N_15827,N_15924);
and U16042 (N_16042,N_15909,N_15991);
nor U16043 (N_16043,N_15867,N_15823);
or U16044 (N_16044,N_15848,N_15804);
or U16045 (N_16045,N_15936,N_15934);
nand U16046 (N_16046,N_15910,N_15992);
and U16047 (N_16047,N_15838,N_15808);
and U16048 (N_16048,N_15959,N_15986);
xnor U16049 (N_16049,N_15817,N_15811);
nor U16050 (N_16050,N_15953,N_15826);
nand U16051 (N_16051,N_15840,N_15888);
xor U16052 (N_16052,N_15849,N_15967);
nor U16053 (N_16053,N_15815,N_15892);
or U16054 (N_16054,N_15882,N_15988);
nor U16055 (N_16055,N_15860,N_15904);
and U16056 (N_16056,N_15920,N_15945);
xnor U16057 (N_16057,N_15832,N_15855);
or U16058 (N_16058,N_15825,N_15940);
and U16059 (N_16059,N_15870,N_15861);
and U16060 (N_16060,N_15900,N_15927);
nor U16061 (N_16061,N_15822,N_15963);
nor U16062 (N_16062,N_15810,N_15921);
nand U16063 (N_16063,N_15901,N_15947);
and U16064 (N_16064,N_15971,N_15896);
or U16065 (N_16065,N_15990,N_15996);
nand U16066 (N_16066,N_15928,N_15985);
and U16067 (N_16067,N_15915,N_15836);
or U16068 (N_16068,N_15839,N_15908);
xor U16069 (N_16069,N_15887,N_15869);
xor U16070 (N_16070,N_15933,N_15813);
nor U16071 (N_16071,N_15884,N_15807);
nor U16072 (N_16072,N_15951,N_15978);
nor U16073 (N_16073,N_15879,N_15989);
nor U16074 (N_16074,N_15983,N_15957);
and U16075 (N_16075,N_15819,N_15976);
and U16076 (N_16076,N_15999,N_15954);
nand U16077 (N_16077,N_15806,N_15821);
nor U16078 (N_16078,N_15995,N_15982);
nand U16079 (N_16079,N_15961,N_15937);
nand U16080 (N_16080,N_15854,N_15868);
and U16081 (N_16081,N_15802,N_15970);
xor U16082 (N_16082,N_15842,N_15845);
xor U16083 (N_16083,N_15975,N_15911);
nand U16084 (N_16084,N_15895,N_15875);
nand U16085 (N_16085,N_15972,N_15844);
nand U16086 (N_16086,N_15809,N_15993);
xor U16087 (N_16087,N_15891,N_15877);
and U16088 (N_16088,N_15926,N_15820);
nand U16089 (N_16089,N_15964,N_15906);
nand U16090 (N_16090,N_15931,N_15949);
and U16091 (N_16091,N_15846,N_15899);
nor U16092 (N_16092,N_15980,N_15997);
and U16093 (N_16093,N_15863,N_15835);
xor U16094 (N_16094,N_15878,N_15897);
nor U16095 (N_16095,N_15841,N_15857);
or U16096 (N_16096,N_15987,N_15828);
nor U16097 (N_16097,N_15948,N_15833);
and U16098 (N_16098,N_15952,N_15834);
nand U16099 (N_16099,N_15894,N_15889);
and U16100 (N_16100,N_15919,N_15891);
nor U16101 (N_16101,N_15917,N_15887);
nor U16102 (N_16102,N_15906,N_15847);
or U16103 (N_16103,N_15978,N_15918);
nor U16104 (N_16104,N_15842,N_15964);
or U16105 (N_16105,N_15848,N_15956);
and U16106 (N_16106,N_15905,N_15939);
and U16107 (N_16107,N_15904,N_15932);
or U16108 (N_16108,N_15942,N_15978);
or U16109 (N_16109,N_15992,N_15946);
xnor U16110 (N_16110,N_15870,N_15857);
and U16111 (N_16111,N_15874,N_15907);
nor U16112 (N_16112,N_15961,N_15928);
or U16113 (N_16113,N_15852,N_15950);
and U16114 (N_16114,N_15841,N_15869);
or U16115 (N_16115,N_15803,N_15903);
and U16116 (N_16116,N_15928,N_15875);
nor U16117 (N_16117,N_15984,N_15804);
and U16118 (N_16118,N_15970,N_15921);
nand U16119 (N_16119,N_15982,N_15948);
xnor U16120 (N_16120,N_15893,N_15967);
or U16121 (N_16121,N_15876,N_15891);
nand U16122 (N_16122,N_15940,N_15979);
nand U16123 (N_16123,N_15945,N_15904);
xnor U16124 (N_16124,N_15949,N_15806);
and U16125 (N_16125,N_15995,N_15998);
xor U16126 (N_16126,N_15808,N_15801);
and U16127 (N_16127,N_15852,N_15849);
xor U16128 (N_16128,N_15956,N_15961);
nand U16129 (N_16129,N_15966,N_15954);
xnor U16130 (N_16130,N_15947,N_15845);
nor U16131 (N_16131,N_15907,N_15939);
or U16132 (N_16132,N_15803,N_15909);
nor U16133 (N_16133,N_15975,N_15822);
xor U16134 (N_16134,N_15970,N_15900);
and U16135 (N_16135,N_15949,N_15887);
nor U16136 (N_16136,N_15972,N_15990);
xor U16137 (N_16137,N_15945,N_15883);
xor U16138 (N_16138,N_15848,N_15849);
xnor U16139 (N_16139,N_15924,N_15908);
and U16140 (N_16140,N_15991,N_15836);
nor U16141 (N_16141,N_15913,N_15840);
and U16142 (N_16142,N_15866,N_15942);
nor U16143 (N_16143,N_15968,N_15850);
nor U16144 (N_16144,N_15917,N_15808);
xor U16145 (N_16145,N_15994,N_15935);
or U16146 (N_16146,N_15892,N_15839);
or U16147 (N_16147,N_15888,N_15858);
and U16148 (N_16148,N_15895,N_15811);
and U16149 (N_16149,N_15803,N_15913);
xor U16150 (N_16150,N_15859,N_15850);
and U16151 (N_16151,N_15823,N_15900);
xor U16152 (N_16152,N_15984,N_15850);
xnor U16153 (N_16153,N_15914,N_15989);
xor U16154 (N_16154,N_15915,N_15952);
and U16155 (N_16155,N_15939,N_15888);
nor U16156 (N_16156,N_15955,N_15832);
or U16157 (N_16157,N_15957,N_15854);
xnor U16158 (N_16158,N_15830,N_15841);
nor U16159 (N_16159,N_15923,N_15951);
nor U16160 (N_16160,N_15913,N_15938);
xor U16161 (N_16161,N_15979,N_15887);
and U16162 (N_16162,N_15844,N_15948);
xnor U16163 (N_16163,N_15922,N_15802);
and U16164 (N_16164,N_15862,N_15998);
nand U16165 (N_16165,N_15997,N_15856);
nor U16166 (N_16166,N_15882,N_15980);
xnor U16167 (N_16167,N_15815,N_15988);
and U16168 (N_16168,N_15880,N_15911);
nor U16169 (N_16169,N_15892,N_15989);
nor U16170 (N_16170,N_15836,N_15939);
or U16171 (N_16171,N_15862,N_15861);
nand U16172 (N_16172,N_15853,N_15913);
nor U16173 (N_16173,N_15970,N_15832);
xor U16174 (N_16174,N_15980,N_15861);
and U16175 (N_16175,N_15857,N_15988);
or U16176 (N_16176,N_15844,N_15864);
nor U16177 (N_16177,N_15986,N_15979);
or U16178 (N_16178,N_15854,N_15948);
and U16179 (N_16179,N_15964,N_15894);
nor U16180 (N_16180,N_15824,N_15882);
and U16181 (N_16181,N_15821,N_15980);
nor U16182 (N_16182,N_15902,N_15844);
nor U16183 (N_16183,N_15894,N_15829);
or U16184 (N_16184,N_15889,N_15911);
xor U16185 (N_16185,N_15951,N_15820);
xnor U16186 (N_16186,N_15910,N_15864);
or U16187 (N_16187,N_15949,N_15995);
nor U16188 (N_16188,N_15926,N_15810);
or U16189 (N_16189,N_15827,N_15889);
or U16190 (N_16190,N_15911,N_15976);
nor U16191 (N_16191,N_15901,N_15848);
and U16192 (N_16192,N_15906,N_15815);
or U16193 (N_16193,N_15969,N_15873);
or U16194 (N_16194,N_15942,N_15882);
xnor U16195 (N_16195,N_15908,N_15946);
nor U16196 (N_16196,N_15865,N_15967);
xnor U16197 (N_16197,N_15837,N_15970);
and U16198 (N_16198,N_15816,N_15890);
and U16199 (N_16199,N_15813,N_15980);
xor U16200 (N_16200,N_16166,N_16003);
xnor U16201 (N_16201,N_16050,N_16095);
xor U16202 (N_16202,N_16026,N_16079);
and U16203 (N_16203,N_16182,N_16129);
xnor U16204 (N_16204,N_16048,N_16187);
xnor U16205 (N_16205,N_16165,N_16043);
xnor U16206 (N_16206,N_16100,N_16186);
xor U16207 (N_16207,N_16034,N_16124);
xor U16208 (N_16208,N_16075,N_16069);
xor U16209 (N_16209,N_16022,N_16140);
nand U16210 (N_16210,N_16099,N_16052);
xnor U16211 (N_16211,N_16198,N_16110);
or U16212 (N_16212,N_16035,N_16059);
nand U16213 (N_16213,N_16102,N_16020);
nand U16214 (N_16214,N_16018,N_16001);
and U16215 (N_16215,N_16096,N_16162);
nand U16216 (N_16216,N_16009,N_16112);
xnor U16217 (N_16217,N_16146,N_16178);
nor U16218 (N_16218,N_16062,N_16177);
xnor U16219 (N_16219,N_16184,N_16155);
xor U16220 (N_16220,N_16065,N_16194);
and U16221 (N_16221,N_16131,N_16080);
xor U16222 (N_16222,N_16078,N_16040);
nand U16223 (N_16223,N_16141,N_16119);
and U16224 (N_16224,N_16006,N_16137);
nand U16225 (N_16225,N_16180,N_16169);
xnor U16226 (N_16226,N_16084,N_16054);
nand U16227 (N_16227,N_16172,N_16197);
and U16228 (N_16228,N_16067,N_16150);
nor U16229 (N_16229,N_16163,N_16045);
or U16230 (N_16230,N_16111,N_16170);
xnor U16231 (N_16231,N_16028,N_16127);
xnor U16232 (N_16232,N_16053,N_16188);
or U16233 (N_16233,N_16107,N_16036);
or U16234 (N_16234,N_16193,N_16176);
nand U16235 (N_16235,N_16021,N_16083);
xor U16236 (N_16236,N_16046,N_16049);
nand U16237 (N_16237,N_16098,N_16060);
or U16238 (N_16238,N_16118,N_16148);
nor U16239 (N_16239,N_16159,N_16016);
and U16240 (N_16240,N_16130,N_16000);
or U16241 (N_16241,N_16076,N_16012);
xnor U16242 (N_16242,N_16106,N_16025);
or U16243 (N_16243,N_16081,N_16144);
and U16244 (N_16244,N_16072,N_16047);
nor U16245 (N_16245,N_16175,N_16063);
nor U16246 (N_16246,N_16199,N_16073);
nor U16247 (N_16247,N_16070,N_16038);
nor U16248 (N_16248,N_16168,N_16024);
or U16249 (N_16249,N_16190,N_16173);
or U16250 (N_16250,N_16074,N_16090);
or U16251 (N_16251,N_16115,N_16174);
nand U16252 (N_16252,N_16088,N_16134);
nor U16253 (N_16253,N_16030,N_16031);
or U16254 (N_16254,N_16160,N_16103);
or U16255 (N_16255,N_16122,N_16109);
nand U16256 (N_16256,N_16116,N_16123);
nor U16257 (N_16257,N_16002,N_16153);
or U16258 (N_16258,N_16139,N_16077);
and U16259 (N_16259,N_16108,N_16051);
xor U16260 (N_16260,N_16013,N_16126);
and U16261 (N_16261,N_16056,N_16014);
and U16262 (N_16262,N_16149,N_16089);
nor U16263 (N_16263,N_16185,N_16086);
and U16264 (N_16264,N_16179,N_16183);
or U16265 (N_16265,N_16041,N_16181);
and U16266 (N_16266,N_16057,N_16097);
nor U16267 (N_16267,N_16101,N_16147);
nor U16268 (N_16268,N_16019,N_16064);
or U16269 (N_16269,N_16113,N_16133);
and U16270 (N_16270,N_16082,N_16058);
xor U16271 (N_16271,N_16042,N_16128);
nor U16272 (N_16272,N_16071,N_16032);
nor U16273 (N_16273,N_16120,N_16037);
and U16274 (N_16274,N_16061,N_16151);
and U16275 (N_16275,N_16117,N_16145);
and U16276 (N_16276,N_16093,N_16004);
nor U16277 (N_16277,N_16010,N_16005);
and U16278 (N_16278,N_16007,N_16152);
or U16279 (N_16279,N_16135,N_16138);
nor U16280 (N_16280,N_16017,N_16068);
or U16281 (N_16281,N_16121,N_16055);
nand U16282 (N_16282,N_16171,N_16189);
and U16283 (N_16283,N_16164,N_16008);
xor U16284 (N_16284,N_16192,N_16011);
and U16285 (N_16285,N_16114,N_16015);
xor U16286 (N_16286,N_16154,N_16039);
and U16287 (N_16287,N_16158,N_16161);
and U16288 (N_16288,N_16136,N_16094);
nand U16289 (N_16289,N_16143,N_16023);
and U16290 (N_16290,N_16092,N_16091);
xnor U16291 (N_16291,N_16033,N_16044);
and U16292 (N_16292,N_16105,N_16125);
and U16293 (N_16293,N_16027,N_16196);
and U16294 (N_16294,N_16029,N_16195);
and U16295 (N_16295,N_16066,N_16191);
and U16296 (N_16296,N_16085,N_16132);
nor U16297 (N_16297,N_16104,N_16087);
nand U16298 (N_16298,N_16142,N_16157);
nand U16299 (N_16299,N_16156,N_16167);
xnor U16300 (N_16300,N_16101,N_16002);
or U16301 (N_16301,N_16022,N_16133);
nand U16302 (N_16302,N_16014,N_16086);
xor U16303 (N_16303,N_16175,N_16112);
nand U16304 (N_16304,N_16186,N_16060);
nor U16305 (N_16305,N_16081,N_16008);
nand U16306 (N_16306,N_16011,N_16065);
xnor U16307 (N_16307,N_16152,N_16146);
xor U16308 (N_16308,N_16156,N_16057);
or U16309 (N_16309,N_16019,N_16025);
xnor U16310 (N_16310,N_16022,N_16112);
or U16311 (N_16311,N_16016,N_16144);
and U16312 (N_16312,N_16033,N_16019);
nand U16313 (N_16313,N_16147,N_16174);
nand U16314 (N_16314,N_16164,N_16026);
and U16315 (N_16315,N_16161,N_16037);
nor U16316 (N_16316,N_16134,N_16032);
or U16317 (N_16317,N_16128,N_16147);
or U16318 (N_16318,N_16055,N_16085);
and U16319 (N_16319,N_16072,N_16068);
nand U16320 (N_16320,N_16152,N_16144);
or U16321 (N_16321,N_16150,N_16078);
xnor U16322 (N_16322,N_16021,N_16065);
xor U16323 (N_16323,N_16159,N_16187);
xor U16324 (N_16324,N_16076,N_16039);
and U16325 (N_16325,N_16185,N_16071);
nor U16326 (N_16326,N_16095,N_16147);
nor U16327 (N_16327,N_16070,N_16172);
nor U16328 (N_16328,N_16084,N_16006);
nand U16329 (N_16329,N_16061,N_16183);
or U16330 (N_16330,N_16142,N_16097);
or U16331 (N_16331,N_16015,N_16073);
nor U16332 (N_16332,N_16047,N_16013);
and U16333 (N_16333,N_16063,N_16192);
nor U16334 (N_16334,N_16161,N_16142);
xor U16335 (N_16335,N_16085,N_16020);
xnor U16336 (N_16336,N_16123,N_16094);
xor U16337 (N_16337,N_16167,N_16160);
xor U16338 (N_16338,N_16158,N_16018);
and U16339 (N_16339,N_16033,N_16143);
xor U16340 (N_16340,N_16047,N_16010);
or U16341 (N_16341,N_16020,N_16094);
xor U16342 (N_16342,N_16060,N_16084);
nand U16343 (N_16343,N_16140,N_16165);
and U16344 (N_16344,N_16144,N_16063);
and U16345 (N_16345,N_16076,N_16173);
or U16346 (N_16346,N_16191,N_16171);
and U16347 (N_16347,N_16060,N_16040);
nand U16348 (N_16348,N_16055,N_16041);
nor U16349 (N_16349,N_16044,N_16053);
xnor U16350 (N_16350,N_16158,N_16020);
nand U16351 (N_16351,N_16152,N_16035);
xnor U16352 (N_16352,N_16054,N_16157);
and U16353 (N_16353,N_16066,N_16055);
nor U16354 (N_16354,N_16019,N_16090);
nand U16355 (N_16355,N_16091,N_16036);
xor U16356 (N_16356,N_16147,N_16003);
or U16357 (N_16357,N_16052,N_16034);
and U16358 (N_16358,N_16168,N_16103);
nor U16359 (N_16359,N_16035,N_16184);
xor U16360 (N_16360,N_16108,N_16041);
nor U16361 (N_16361,N_16188,N_16063);
nor U16362 (N_16362,N_16045,N_16172);
nand U16363 (N_16363,N_16146,N_16064);
and U16364 (N_16364,N_16121,N_16175);
xnor U16365 (N_16365,N_16197,N_16029);
and U16366 (N_16366,N_16189,N_16175);
nand U16367 (N_16367,N_16005,N_16166);
nand U16368 (N_16368,N_16042,N_16120);
or U16369 (N_16369,N_16005,N_16157);
nor U16370 (N_16370,N_16167,N_16084);
or U16371 (N_16371,N_16140,N_16085);
or U16372 (N_16372,N_16163,N_16190);
and U16373 (N_16373,N_16026,N_16017);
xnor U16374 (N_16374,N_16072,N_16064);
nand U16375 (N_16375,N_16148,N_16094);
nand U16376 (N_16376,N_16008,N_16089);
or U16377 (N_16377,N_16138,N_16075);
and U16378 (N_16378,N_16085,N_16056);
or U16379 (N_16379,N_16037,N_16094);
and U16380 (N_16380,N_16048,N_16002);
or U16381 (N_16381,N_16173,N_16162);
nor U16382 (N_16382,N_16085,N_16007);
nand U16383 (N_16383,N_16126,N_16186);
xor U16384 (N_16384,N_16169,N_16152);
xnor U16385 (N_16385,N_16168,N_16007);
nand U16386 (N_16386,N_16128,N_16064);
nor U16387 (N_16387,N_16186,N_16055);
or U16388 (N_16388,N_16039,N_16117);
and U16389 (N_16389,N_16043,N_16143);
xnor U16390 (N_16390,N_16094,N_16096);
and U16391 (N_16391,N_16160,N_16178);
nor U16392 (N_16392,N_16003,N_16087);
and U16393 (N_16393,N_16154,N_16081);
nand U16394 (N_16394,N_16042,N_16022);
and U16395 (N_16395,N_16125,N_16189);
nand U16396 (N_16396,N_16042,N_16196);
or U16397 (N_16397,N_16097,N_16092);
or U16398 (N_16398,N_16002,N_16051);
nand U16399 (N_16399,N_16068,N_16055);
xor U16400 (N_16400,N_16352,N_16340);
or U16401 (N_16401,N_16383,N_16376);
nand U16402 (N_16402,N_16368,N_16274);
and U16403 (N_16403,N_16338,N_16325);
or U16404 (N_16404,N_16247,N_16281);
xor U16405 (N_16405,N_16307,N_16280);
nand U16406 (N_16406,N_16333,N_16387);
xnor U16407 (N_16407,N_16201,N_16283);
xor U16408 (N_16408,N_16207,N_16299);
or U16409 (N_16409,N_16379,N_16298);
xnor U16410 (N_16410,N_16222,N_16301);
xor U16411 (N_16411,N_16339,N_16311);
or U16412 (N_16412,N_16388,N_16219);
nand U16413 (N_16413,N_16305,N_16221);
or U16414 (N_16414,N_16334,N_16269);
xnor U16415 (N_16415,N_16364,N_16258);
nor U16416 (N_16416,N_16277,N_16202);
or U16417 (N_16417,N_16239,N_16291);
xnor U16418 (N_16418,N_16211,N_16342);
xnor U16419 (N_16419,N_16275,N_16341);
or U16420 (N_16420,N_16245,N_16214);
or U16421 (N_16421,N_16223,N_16204);
xor U16422 (N_16422,N_16208,N_16396);
nand U16423 (N_16423,N_16357,N_16385);
and U16424 (N_16424,N_16365,N_16308);
and U16425 (N_16425,N_16351,N_16215);
xnor U16426 (N_16426,N_16398,N_16251);
or U16427 (N_16427,N_16366,N_16246);
and U16428 (N_16428,N_16248,N_16389);
and U16429 (N_16429,N_16256,N_16312);
nand U16430 (N_16430,N_16267,N_16288);
or U16431 (N_16431,N_16271,N_16331);
nand U16432 (N_16432,N_16330,N_16300);
nand U16433 (N_16433,N_16345,N_16290);
and U16434 (N_16434,N_16336,N_16217);
or U16435 (N_16435,N_16350,N_16209);
or U16436 (N_16436,N_16260,N_16354);
or U16437 (N_16437,N_16272,N_16380);
and U16438 (N_16438,N_16335,N_16319);
nor U16439 (N_16439,N_16367,N_16273);
or U16440 (N_16440,N_16250,N_16268);
xor U16441 (N_16441,N_16287,N_16241);
nand U16442 (N_16442,N_16295,N_16276);
and U16443 (N_16443,N_16372,N_16393);
or U16444 (N_16444,N_16369,N_16332);
nand U16445 (N_16445,N_16284,N_16285);
xor U16446 (N_16446,N_16254,N_16234);
or U16447 (N_16447,N_16306,N_16390);
and U16448 (N_16448,N_16228,N_16375);
and U16449 (N_16449,N_16203,N_16294);
nand U16450 (N_16450,N_16293,N_16259);
nand U16451 (N_16451,N_16264,N_16310);
xnor U16452 (N_16452,N_16252,N_16328);
or U16453 (N_16453,N_16329,N_16244);
xnor U16454 (N_16454,N_16218,N_16282);
and U16455 (N_16455,N_16317,N_16270);
and U16456 (N_16456,N_16303,N_16313);
xnor U16457 (N_16457,N_16216,N_16316);
nor U16458 (N_16458,N_16337,N_16381);
xnor U16459 (N_16459,N_16257,N_16286);
or U16460 (N_16460,N_16324,N_16394);
nand U16461 (N_16461,N_16384,N_16240);
nand U16462 (N_16462,N_16348,N_16263);
xnor U16463 (N_16463,N_16349,N_16382);
or U16464 (N_16464,N_16253,N_16326);
and U16465 (N_16465,N_16210,N_16353);
nor U16466 (N_16466,N_16289,N_16370);
xnor U16467 (N_16467,N_16360,N_16297);
and U16468 (N_16468,N_16231,N_16315);
nand U16469 (N_16469,N_16279,N_16206);
nand U16470 (N_16470,N_16397,N_16361);
and U16471 (N_16471,N_16318,N_16236);
and U16472 (N_16472,N_16321,N_16224);
nor U16473 (N_16473,N_16230,N_16386);
or U16474 (N_16474,N_16304,N_16255);
xnor U16475 (N_16475,N_16378,N_16226);
xnor U16476 (N_16476,N_16359,N_16261);
nor U16477 (N_16477,N_16212,N_16265);
and U16478 (N_16478,N_16322,N_16220);
nor U16479 (N_16479,N_16302,N_16343);
nand U16480 (N_16480,N_16320,N_16344);
or U16481 (N_16481,N_16227,N_16249);
nor U16482 (N_16482,N_16395,N_16356);
or U16483 (N_16483,N_16374,N_16278);
and U16484 (N_16484,N_16233,N_16235);
nand U16485 (N_16485,N_16346,N_16363);
or U16486 (N_16486,N_16296,N_16242);
and U16487 (N_16487,N_16200,N_16347);
nor U16488 (N_16488,N_16213,N_16205);
nand U16489 (N_16489,N_16229,N_16225);
and U16490 (N_16490,N_16327,N_16362);
nor U16491 (N_16491,N_16243,N_16262);
or U16492 (N_16492,N_16399,N_16355);
nor U16493 (N_16493,N_16237,N_16373);
and U16494 (N_16494,N_16266,N_16377);
and U16495 (N_16495,N_16292,N_16314);
nand U16496 (N_16496,N_16391,N_16238);
xnor U16497 (N_16497,N_16323,N_16371);
nor U16498 (N_16498,N_16392,N_16309);
nor U16499 (N_16499,N_16358,N_16232);
nand U16500 (N_16500,N_16238,N_16388);
and U16501 (N_16501,N_16248,N_16293);
nand U16502 (N_16502,N_16279,N_16356);
nor U16503 (N_16503,N_16309,N_16332);
or U16504 (N_16504,N_16348,N_16371);
xnor U16505 (N_16505,N_16308,N_16288);
nand U16506 (N_16506,N_16355,N_16269);
nand U16507 (N_16507,N_16275,N_16280);
xnor U16508 (N_16508,N_16351,N_16333);
and U16509 (N_16509,N_16214,N_16211);
and U16510 (N_16510,N_16288,N_16382);
and U16511 (N_16511,N_16248,N_16276);
xnor U16512 (N_16512,N_16324,N_16237);
nand U16513 (N_16513,N_16303,N_16264);
or U16514 (N_16514,N_16242,N_16243);
or U16515 (N_16515,N_16359,N_16272);
or U16516 (N_16516,N_16383,N_16388);
or U16517 (N_16517,N_16293,N_16268);
xnor U16518 (N_16518,N_16381,N_16299);
xnor U16519 (N_16519,N_16222,N_16217);
xnor U16520 (N_16520,N_16313,N_16384);
nand U16521 (N_16521,N_16361,N_16237);
nor U16522 (N_16522,N_16268,N_16281);
and U16523 (N_16523,N_16391,N_16263);
and U16524 (N_16524,N_16251,N_16359);
nand U16525 (N_16525,N_16308,N_16228);
or U16526 (N_16526,N_16263,N_16279);
or U16527 (N_16527,N_16278,N_16321);
xnor U16528 (N_16528,N_16299,N_16264);
and U16529 (N_16529,N_16343,N_16231);
or U16530 (N_16530,N_16290,N_16217);
or U16531 (N_16531,N_16304,N_16240);
and U16532 (N_16532,N_16276,N_16292);
nand U16533 (N_16533,N_16340,N_16250);
nand U16534 (N_16534,N_16240,N_16234);
nand U16535 (N_16535,N_16322,N_16341);
xor U16536 (N_16536,N_16348,N_16271);
and U16537 (N_16537,N_16297,N_16311);
xnor U16538 (N_16538,N_16364,N_16368);
and U16539 (N_16539,N_16226,N_16247);
nand U16540 (N_16540,N_16217,N_16398);
xor U16541 (N_16541,N_16382,N_16389);
xor U16542 (N_16542,N_16215,N_16309);
xnor U16543 (N_16543,N_16246,N_16342);
and U16544 (N_16544,N_16247,N_16219);
xnor U16545 (N_16545,N_16269,N_16386);
nor U16546 (N_16546,N_16240,N_16238);
and U16547 (N_16547,N_16357,N_16376);
nand U16548 (N_16548,N_16289,N_16327);
or U16549 (N_16549,N_16365,N_16228);
and U16550 (N_16550,N_16265,N_16237);
and U16551 (N_16551,N_16272,N_16250);
nor U16552 (N_16552,N_16260,N_16357);
and U16553 (N_16553,N_16316,N_16237);
nor U16554 (N_16554,N_16331,N_16299);
nand U16555 (N_16555,N_16239,N_16296);
xor U16556 (N_16556,N_16256,N_16221);
or U16557 (N_16557,N_16217,N_16390);
nor U16558 (N_16558,N_16285,N_16363);
nor U16559 (N_16559,N_16302,N_16370);
xnor U16560 (N_16560,N_16212,N_16213);
and U16561 (N_16561,N_16318,N_16311);
nor U16562 (N_16562,N_16392,N_16278);
nand U16563 (N_16563,N_16235,N_16263);
xor U16564 (N_16564,N_16386,N_16299);
and U16565 (N_16565,N_16266,N_16228);
xnor U16566 (N_16566,N_16344,N_16337);
and U16567 (N_16567,N_16217,N_16369);
or U16568 (N_16568,N_16290,N_16274);
and U16569 (N_16569,N_16327,N_16358);
or U16570 (N_16570,N_16220,N_16225);
and U16571 (N_16571,N_16336,N_16314);
xnor U16572 (N_16572,N_16259,N_16200);
nor U16573 (N_16573,N_16330,N_16399);
xnor U16574 (N_16574,N_16315,N_16297);
nand U16575 (N_16575,N_16327,N_16369);
or U16576 (N_16576,N_16327,N_16231);
nor U16577 (N_16577,N_16340,N_16301);
or U16578 (N_16578,N_16213,N_16372);
nand U16579 (N_16579,N_16249,N_16243);
nor U16580 (N_16580,N_16260,N_16252);
xor U16581 (N_16581,N_16281,N_16228);
or U16582 (N_16582,N_16308,N_16304);
or U16583 (N_16583,N_16299,N_16382);
nand U16584 (N_16584,N_16352,N_16365);
nand U16585 (N_16585,N_16333,N_16314);
or U16586 (N_16586,N_16355,N_16379);
or U16587 (N_16587,N_16215,N_16211);
nand U16588 (N_16588,N_16235,N_16391);
nand U16589 (N_16589,N_16346,N_16204);
nor U16590 (N_16590,N_16362,N_16231);
xor U16591 (N_16591,N_16375,N_16339);
or U16592 (N_16592,N_16222,N_16280);
or U16593 (N_16593,N_16397,N_16240);
nor U16594 (N_16594,N_16295,N_16297);
and U16595 (N_16595,N_16307,N_16322);
nand U16596 (N_16596,N_16370,N_16358);
nor U16597 (N_16597,N_16256,N_16384);
nand U16598 (N_16598,N_16319,N_16234);
xor U16599 (N_16599,N_16273,N_16279);
and U16600 (N_16600,N_16532,N_16458);
xnor U16601 (N_16601,N_16508,N_16538);
nand U16602 (N_16602,N_16580,N_16541);
and U16603 (N_16603,N_16554,N_16450);
or U16604 (N_16604,N_16475,N_16403);
xor U16605 (N_16605,N_16457,N_16534);
and U16606 (N_16606,N_16527,N_16407);
xor U16607 (N_16607,N_16524,N_16591);
nor U16608 (N_16608,N_16451,N_16424);
nand U16609 (N_16609,N_16582,N_16455);
nor U16610 (N_16610,N_16565,N_16509);
nor U16611 (N_16611,N_16492,N_16537);
and U16612 (N_16612,N_16506,N_16493);
xor U16613 (N_16613,N_16526,N_16523);
or U16614 (N_16614,N_16406,N_16401);
or U16615 (N_16615,N_16445,N_16415);
nor U16616 (N_16616,N_16471,N_16469);
xnor U16617 (N_16617,N_16483,N_16474);
xor U16618 (N_16618,N_16557,N_16564);
xnor U16619 (N_16619,N_16426,N_16536);
or U16620 (N_16620,N_16413,N_16411);
and U16621 (N_16621,N_16468,N_16405);
nand U16622 (N_16622,N_16545,N_16590);
nand U16623 (N_16623,N_16431,N_16593);
and U16624 (N_16624,N_16497,N_16423);
nor U16625 (N_16625,N_16435,N_16404);
and U16626 (N_16626,N_16425,N_16438);
and U16627 (N_16627,N_16546,N_16560);
xor U16628 (N_16628,N_16465,N_16454);
xnor U16629 (N_16629,N_16491,N_16495);
and U16630 (N_16630,N_16486,N_16409);
nor U16631 (N_16631,N_16459,N_16592);
nand U16632 (N_16632,N_16446,N_16449);
xor U16633 (N_16633,N_16539,N_16470);
or U16634 (N_16634,N_16430,N_16441);
or U16635 (N_16635,N_16453,N_16562);
or U16636 (N_16636,N_16416,N_16584);
or U16637 (N_16637,N_16595,N_16583);
xor U16638 (N_16638,N_16442,N_16480);
or U16639 (N_16639,N_16520,N_16428);
xor U16640 (N_16640,N_16500,N_16596);
nand U16641 (N_16641,N_16598,N_16587);
nor U16642 (N_16642,N_16577,N_16440);
or U16643 (N_16643,N_16414,N_16549);
and U16644 (N_16644,N_16512,N_16568);
xnor U16645 (N_16645,N_16575,N_16408);
xor U16646 (N_16646,N_16586,N_16597);
nand U16647 (N_16647,N_16427,N_16533);
and U16648 (N_16648,N_16507,N_16420);
nand U16649 (N_16649,N_16462,N_16437);
nor U16650 (N_16650,N_16410,N_16429);
and U16651 (N_16651,N_16467,N_16511);
nor U16652 (N_16652,N_16515,N_16400);
xor U16653 (N_16653,N_16553,N_16481);
and U16654 (N_16654,N_16556,N_16552);
nand U16655 (N_16655,N_16517,N_16436);
nand U16656 (N_16656,N_16518,N_16589);
nand U16657 (N_16657,N_16514,N_16448);
nand U16658 (N_16658,N_16461,N_16558);
and U16659 (N_16659,N_16463,N_16447);
xnor U16660 (N_16660,N_16529,N_16528);
and U16661 (N_16661,N_16525,N_16464);
nand U16662 (N_16662,N_16460,N_16485);
and U16663 (N_16663,N_16513,N_16466);
and U16664 (N_16664,N_16519,N_16540);
and U16665 (N_16665,N_16418,N_16402);
nor U16666 (N_16666,N_16588,N_16531);
and U16667 (N_16667,N_16574,N_16547);
nor U16668 (N_16668,N_16473,N_16421);
xor U16669 (N_16669,N_16548,N_16570);
and U16670 (N_16670,N_16422,N_16510);
nand U16671 (N_16671,N_16444,N_16555);
nand U16672 (N_16672,N_16478,N_16521);
nand U16673 (N_16673,N_16550,N_16571);
and U16674 (N_16674,N_16503,N_16522);
and U16675 (N_16675,N_16579,N_16496);
xor U16676 (N_16676,N_16559,N_16412);
nor U16677 (N_16677,N_16419,N_16504);
or U16678 (N_16678,N_16578,N_16487);
or U16679 (N_16679,N_16499,N_16498);
nand U16680 (N_16680,N_16542,N_16566);
or U16681 (N_16681,N_16585,N_16572);
nand U16682 (N_16682,N_16432,N_16452);
nand U16683 (N_16683,N_16456,N_16434);
or U16684 (N_16684,N_16494,N_16482);
and U16685 (N_16685,N_16569,N_16476);
and U16686 (N_16686,N_16489,N_16479);
xor U16687 (N_16687,N_16439,N_16544);
or U16688 (N_16688,N_16484,N_16573);
nand U16689 (N_16689,N_16551,N_16563);
or U16690 (N_16690,N_16516,N_16477);
or U16691 (N_16691,N_16561,N_16581);
xor U16692 (N_16692,N_16443,N_16599);
or U16693 (N_16693,N_16472,N_16501);
and U16694 (N_16694,N_16417,N_16594);
or U16695 (N_16695,N_16543,N_16502);
nand U16696 (N_16696,N_16490,N_16567);
nor U16697 (N_16697,N_16576,N_16505);
or U16698 (N_16698,N_16530,N_16535);
nor U16699 (N_16699,N_16433,N_16488);
and U16700 (N_16700,N_16498,N_16446);
and U16701 (N_16701,N_16530,N_16408);
or U16702 (N_16702,N_16418,N_16451);
xor U16703 (N_16703,N_16437,N_16448);
or U16704 (N_16704,N_16559,N_16406);
or U16705 (N_16705,N_16569,N_16500);
or U16706 (N_16706,N_16452,N_16513);
xor U16707 (N_16707,N_16488,N_16506);
or U16708 (N_16708,N_16544,N_16499);
and U16709 (N_16709,N_16585,N_16468);
nand U16710 (N_16710,N_16442,N_16571);
or U16711 (N_16711,N_16536,N_16575);
nor U16712 (N_16712,N_16456,N_16439);
or U16713 (N_16713,N_16421,N_16519);
xnor U16714 (N_16714,N_16529,N_16499);
and U16715 (N_16715,N_16583,N_16581);
or U16716 (N_16716,N_16564,N_16470);
or U16717 (N_16717,N_16550,N_16560);
or U16718 (N_16718,N_16537,N_16552);
and U16719 (N_16719,N_16519,N_16593);
xor U16720 (N_16720,N_16424,N_16469);
xnor U16721 (N_16721,N_16539,N_16452);
xor U16722 (N_16722,N_16449,N_16584);
nor U16723 (N_16723,N_16441,N_16489);
or U16724 (N_16724,N_16472,N_16475);
xor U16725 (N_16725,N_16588,N_16475);
and U16726 (N_16726,N_16437,N_16472);
xor U16727 (N_16727,N_16553,N_16556);
and U16728 (N_16728,N_16499,N_16419);
xnor U16729 (N_16729,N_16450,N_16425);
nor U16730 (N_16730,N_16529,N_16455);
and U16731 (N_16731,N_16467,N_16403);
nand U16732 (N_16732,N_16506,N_16542);
nand U16733 (N_16733,N_16570,N_16474);
or U16734 (N_16734,N_16491,N_16454);
nor U16735 (N_16735,N_16566,N_16400);
nand U16736 (N_16736,N_16470,N_16452);
and U16737 (N_16737,N_16480,N_16581);
and U16738 (N_16738,N_16446,N_16587);
nand U16739 (N_16739,N_16457,N_16566);
nand U16740 (N_16740,N_16427,N_16582);
nor U16741 (N_16741,N_16545,N_16418);
or U16742 (N_16742,N_16460,N_16478);
nand U16743 (N_16743,N_16531,N_16537);
and U16744 (N_16744,N_16599,N_16584);
or U16745 (N_16745,N_16585,N_16591);
or U16746 (N_16746,N_16409,N_16480);
xnor U16747 (N_16747,N_16407,N_16478);
nor U16748 (N_16748,N_16412,N_16534);
nor U16749 (N_16749,N_16445,N_16426);
and U16750 (N_16750,N_16425,N_16573);
nor U16751 (N_16751,N_16427,N_16472);
and U16752 (N_16752,N_16532,N_16412);
xor U16753 (N_16753,N_16449,N_16461);
nor U16754 (N_16754,N_16598,N_16548);
nor U16755 (N_16755,N_16498,N_16415);
or U16756 (N_16756,N_16542,N_16475);
and U16757 (N_16757,N_16518,N_16473);
nor U16758 (N_16758,N_16573,N_16465);
and U16759 (N_16759,N_16572,N_16569);
nand U16760 (N_16760,N_16553,N_16499);
nor U16761 (N_16761,N_16544,N_16446);
nand U16762 (N_16762,N_16505,N_16425);
nand U16763 (N_16763,N_16469,N_16530);
nand U16764 (N_16764,N_16476,N_16506);
nor U16765 (N_16765,N_16417,N_16455);
nand U16766 (N_16766,N_16501,N_16583);
xor U16767 (N_16767,N_16403,N_16411);
xnor U16768 (N_16768,N_16564,N_16597);
and U16769 (N_16769,N_16521,N_16570);
xnor U16770 (N_16770,N_16585,N_16553);
nor U16771 (N_16771,N_16551,N_16448);
and U16772 (N_16772,N_16448,N_16428);
and U16773 (N_16773,N_16550,N_16528);
and U16774 (N_16774,N_16422,N_16433);
or U16775 (N_16775,N_16579,N_16540);
and U16776 (N_16776,N_16579,N_16577);
or U16777 (N_16777,N_16495,N_16572);
or U16778 (N_16778,N_16562,N_16511);
nand U16779 (N_16779,N_16487,N_16545);
xor U16780 (N_16780,N_16546,N_16587);
or U16781 (N_16781,N_16573,N_16444);
xor U16782 (N_16782,N_16401,N_16597);
and U16783 (N_16783,N_16515,N_16443);
nor U16784 (N_16784,N_16423,N_16430);
xnor U16785 (N_16785,N_16573,N_16593);
and U16786 (N_16786,N_16523,N_16539);
nand U16787 (N_16787,N_16519,N_16416);
or U16788 (N_16788,N_16511,N_16546);
nor U16789 (N_16789,N_16568,N_16456);
nand U16790 (N_16790,N_16509,N_16530);
xnor U16791 (N_16791,N_16518,N_16586);
or U16792 (N_16792,N_16519,N_16435);
nand U16793 (N_16793,N_16482,N_16486);
nand U16794 (N_16794,N_16487,N_16565);
nor U16795 (N_16795,N_16539,N_16473);
or U16796 (N_16796,N_16461,N_16467);
nor U16797 (N_16797,N_16504,N_16563);
xnor U16798 (N_16798,N_16580,N_16508);
nand U16799 (N_16799,N_16486,N_16570);
nor U16800 (N_16800,N_16797,N_16736);
nor U16801 (N_16801,N_16633,N_16704);
nand U16802 (N_16802,N_16627,N_16787);
or U16803 (N_16803,N_16756,N_16640);
or U16804 (N_16804,N_16680,N_16688);
nand U16805 (N_16805,N_16631,N_16632);
and U16806 (N_16806,N_16600,N_16603);
nand U16807 (N_16807,N_16690,N_16724);
nand U16808 (N_16808,N_16618,N_16611);
nor U16809 (N_16809,N_16612,N_16749);
or U16810 (N_16810,N_16773,N_16671);
nand U16811 (N_16811,N_16654,N_16616);
or U16812 (N_16812,N_16685,N_16694);
and U16813 (N_16813,N_16684,N_16652);
or U16814 (N_16814,N_16635,N_16614);
nand U16815 (N_16815,N_16657,N_16795);
nor U16816 (N_16816,N_16769,N_16759);
nor U16817 (N_16817,N_16630,N_16605);
nor U16818 (N_16818,N_16659,N_16711);
and U16819 (N_16819,N_16698,N_16753);
and U16820 (N_16820,N_16726,N_16757);
nand U16821 (N_16821,N_16661,N_16799);
or U16822 (N_16822,N_16709,N_16766);
xnor U16823 (N_16823,N_16682,N_16708);
nand U16824 (N_16824,N_16697,N_16707);
xor U16825 (N_16825,N_16744,N_16721);
and U16826 (N_16826,N_16676,N_16686);
nand U16827 (N_16827,N_16731,N_16642);
and U16828 (N_16828,N_16663,N_16705);
nor U16829 (N_16829,N_16628,N_16734);
and U16830 (N_16830,N_16762,N_16728);
nor U16831 (N_16831,N_16702,N_16788);
xnor U16832 (N_16832,N_16645,N_16715);
and U16833 (N_16833,N_16717,N_16778);
xor U16834 (N_16834,N_16729,N_16718);
or U16835 (N_16835,N_16782,N_16752);
xnor U16836 (N_16836,N_16667,N_16783);
or U16837 (N_16837,N_16660,N_16754);
nand U16838 (N_16838,N_16735,N_16687);
and U16839 (N_16839,N_16789,N_16621);
xor U16840 (N_16840,N_16626,N_16784);
nor U16841 (N_16841,N_16674,N_16706);
or U16842 (N_16842,N_16779,N_16609);
and U16843 (N_16843,N_16748,N_16741);
or U16844 (N_16844,N_16641,N_16745);
nor U16845 (N_16845,N_16768,N_16622);
or U16846 (N_16846,N_16722,N_16791);
and U16847 (N_16847,N_16774,N_16740);
nor U16848 (N_16848,N_16777,N_16747);
xnor U16849 (N_16849,N_16655,N_16607);
xor U16850 (N_16850,N_16683,N_16672);
and U16851 (N_16851,N_16796,N_16712);
and U16852 (N_16852,N_16700,N_16647);
xor U16853 (N_16853,N_16691,N_16629);
or U16854 (N_16854,N_16695,N_16623);
xnor U16855 (N_16855,N_16798,N_16613);
nor U16856 (N_16856,N_16606,N_16742);
nor U16857 (N_16857,N_16716,N_16692);
nand U16858 (N_16858,N_16601,N_16637);
xnor U16859 (N_16859,N_16602,N_16701);
xnor U16860 (N_16860,N_16689,N_16758);
nor U16861 (N_16861,N_16764,N_16604);
nor U16862 (N_16862,N_16790,N_16678);
and U16863 (N_16863,N_16649,N_16737);
nand U16864 (N_16864,N_16666,N_16634);
nand U16865 (N_16865,N_16639,N_16670);
xor U16866 (N_16866,N_16608,N_16703);
or U16867 (N_16867,N_16765,N_16794);
nor U16868 (N_16868,N_16620,N_16679);
or U16869 (N_16869,N_16693,N_16786);
and U16870 (N_16870,N_16710,N_16732);
xor U16871 (N_16871,N_16760,N_16719);
and U16872 (N_16872,N_16699,N_16733);
or U16873 (N_16873,N_16669,N_16668);
or U16874 (N_16874,N_16776,N_16624);
nand U16875 (N_16875,N_16761,N_16648);
and U16876 (N_16876,N_16725,N_16644);
xor U16877 (N_16877,N_16739,N_16767);
xnor U16878 (N_16878,N_16780,N_16743);
nand U16879 (N_16879,N_16793,N_16755);
xor U16880 (N_16880,N_16673,N_16650);
nand U16881 (N_16881,N_16730,N_16615);
nor U16882 (N_16882,N_16625,N_16638);
or U16883 (N_16883,N_16646,N_16770);
nand U16884 (N_16884,N_16636,N_16696);
and U16885 (N_16885,N_16751,N_16675);
xor U16886 (N_16886,N_16651,N_16775);
or U16887 (N_16887,N_16658,N_16714);
nor U16888 (N_16888,N_16723,N_16785);
xor U16889 (N_16889,N_16763,N_16617);
nand U16890 (N_16890,N_16664,N_16656);
and U16891 (N_16891,N_16750,N_16643);
nand U16892 (N_16892,N_16746,N_16781);
nor U16893 (N_16893,N_16610,N_16665);
or U16894 (N_16894,N_16720,N_16619);
or U16895 (N_16895,N_16677,N_16681);
or U16896 (N_16896,N_16792,N_16653);
xnor U16897 (N_16897,N_16662,N_16771);
nor U16898 (N_16898,N_16772,N_16738);
and U16899 (N_16899,N_16713,N_16727);
and U16900 (N_16900,N_16699,N_16694);
nor U16901 (N_16901,N_16766,N_16646);
or U16902 (N_16902,N_16770,N_16609);
or U16903 (N_16903,N_16718,N_16692);
nor U16904 (N_16904,N_16724,N_16709);
nand U16905 (N_16905,N_16761,N_16685);
nand U16906 (N_16906,N_16657,N_16735);
and U16907 (N_16907,N_16714,N_16688);
nand U16908 (N_16908,N_16701,N_16726);
xor U16909 (N_16909,N_16662,N_16664);
nand U16910 (N_16910,N_16722,N_16723);
nand U16911 (N_16911,N_16640,N_16681);
nand U16912 (N_16912,N_16784,N_16705);
or U16913 (N_16913,N_16609,N_16641);
nand U16914 (N_16914,N_16716,N_16654);
xor U16915 (N_16915,N_16658,N_16706);
nand U16916 (N_16916,N_16667,N_16655);
nand U16917 (N_16917,N_16703,N_16705);
or U16918 (N_16918,N_16642,N_16646);
nor U16919 (N_16919,N_16616,N_16637);
or U16920 (N_16920,N_16710,N_16737);
nand U16921 (N_16921,N_16692,N_16683);
and U16922 (N_16922,N_16641,N_16634);
or U16923 (N_16923,N_16791,N_16631);
or U16924 (N_16924,N_16741,N_16755);
nor U16925 (N_16925,N_16690,N_16714);
and U16926 (N_16926,N_16648,N_16611);
nor U16927 (N_16927,N_16755,N_16724);
or U16928 (N_16928,N_16667,N_16712);
nor U16929 (N_16929,N_16684,N_16750);
nor U16930 (N_16930,N_16699,N_16749);
xor U16931 (N_16931,N_16649,N_16724);
nor U16932 (N_16932,N_16790,N_16658);
and U16933 (N_16933,N_16743,N_16756);
nor U16934 (N_16934,N_16646,N_16600);
nand U16935 (N_16935,N_16775,N_16665);
xnor U16936 (N_16936,N_16664,N_16685);
and U16937 (N_16937,N_16691,N_16797);
nand U16938 (N_16938,N_16683,N_16678);
xnor U16939 (N_16939,N_16609,N_16785);
xor U16940 (N_16940,N_16612,N_16667);
xnor U16941 (N_16941,N_16774,N_16647);
or U16942 (N_16942,N_16664,N_16643);
nand U16943 (N_16943,N_16658,N_16730);
xor U16944 (N_16944,N_16757,N_16609);
nor U16945 (N_16945,N_16632,N_16628);
and U16946 (N_16946,N_16693,N_16758);
xnor U16947 (N_16947,N_16730,N_16742);
and U16948 (N_16948,N_16786,N_16739);
or U16949 (N_16949,N_16705,N_16769);
xor U16950 (N_16950,N_16605,N_16609);
nor U16951 (N_16951,N_16645,N_16743);
xnor U16952 (N_16952,N_16749,N_16641);
xnor U16953 (N_16953,N_16763,N_16651);
xnor U16954 (N_16954,N_16611,N_16717);
or U16955 (N_16955,N_16714,N_16760);
nand U16956 (N_16956,N_16623,N_16645);
or U16957 (N_16957,N_16730,N_16639);
nor U16958 (N_16958,N_16772,N_16671);
xor U16959 (N_16959,N_16726,N_16640);
nor U16960 (N_16960,N_16722,N_16703);
nand U16961 (N_16961,N_16602,N_16761);
nand U16962 (N_16962,N_16775,N_16779);
nand U16963 (N_16963,N_16741,N_16693);
and U16964 (N_16964,N_16652,N_16779);
xor U16965 (N_16965,N_16708,N_16729);
nor U16966 (N_16966,N_16610,N_16637);
nand U16967 (N_16967,N_16714,N_16731);
nor U16968 (N_16968,N_16761,N_16764);
xor U16969 (N_16969,N_16659,N_16634);
nand U16970 (N_16970,N_16695,N_16716);
nor U16971 (N_16971,N_16785,N_16643);
and U16972 (N_16972,N_16642,N_16778);
xor U16973 (N_16973,N_16685,N_16627);
xor U16974 (N_16974,N_16731,N_16704);
xnor U16975 (N_16975,N_16707,N_16676);
and U16976 (N_16976,N_16660,N_16603);
nand U16977 (N_16977,N_16779,N_16729);
or U16978 (N_16978,N_16651,N_16718);
nor U16979 (N_16979,N_16709,N_16644);
xor U16980 (N_16980,N_16735,N_16644);
nor U16981 (N_16981,N_16656,N_16737);
or U16982 (N_16982,N_16744,N_16777);
and U16983 (N_16983,N_16601,N_16684);
xnor U16984 (N_16984,N_16679,N_16753);
or U16985 (N_16985,N_16687,N_16705);
xor U16986 (N_16986,N_16645,N_16643);
xnor U16987 (N_16987,N_16674,N_16764);
or U16988 (N_16988,N_16673,N_16707);
xnor U16989 (N_16989,N_16667,N_16652);
and U16990 (N_16990,N_16765,N_16777);
and U16991 (N_16991,N_16644,N_16742);
and U16992 (N_16992,N_16685,N_16746);
and U16993 (N_16993,N_16663,N_16798);
or U16994 (N_16994,N_16677,N_16679);
nor U16995 (N_16995,N_16723,N_16728);
and U16996 (N_16996,N_16746,N_16710);
nor U16997 (N_16997,N_16748,N_16653);
and U16998 (N_16998,N_16746,N_16632);
xnor U16999 (N_16999,N_16786,N_16738);
xnor U17000 (N_17000,N_16894,N_16860);
xor U17001 (N_17001,N_16806,N_16858);
nand U17002 (N_17002,N_16856,N_16804);
xor U17003 (N_17003,N_16924,N_16938);
or U17004 (N_17004,N_16971,N_16957);
and U17005 (N_17005,N_16961,N_16829);
or U17006 (N_17006,N_16948,N_16819);
and U17007 (N_17007,N_16964,N_16901);
nand U17008 (N_17008,N_16807,N_16976);
nand U17009 (N_17009,N_16913,N_16881);
or U17010 (N_17010,N_16968,N_16851);
nand U17011 (N_17011,N_16973,N_16911);
or U17012 (N_17012,N_16930,N_16842);
nand U17013 (N_17013,N_16996,N_16833);
xor U17014 (N_17014,N_16910,N_16945);
xor U17015 (N_17015,N_16823,N_16831);
and U17016 (N_17016,N_16850,N_16951);
or U17017 (N_17017,N_16918,N_16905);
and U17018 (N_17018,N_16917,N_16977);
nand U17019 (N_17019,N_16962,N_16970);
nand U17020 (N_17020,N_16869,N_16998);
or U17021 (N_17021,N_16866,N_16954);
nand U17022 (N_17022,N_16812,N_16999);
and U17023 (N_17023,N_16947,N_16893);
and U17024 (N_17024,N_16934,N_16890);
and U17025 (N_17025,N_16800,N_16848);
or U17026 (N_17026,N_16925,N_16939);
nor U17027 (N_17027,N_16963,N_16845);
xor U17028 (N_17028,N_16814,N_16808);
nand U17029 (N_17029,N_16825,N_16928);
nand U17030 (N_17030,N_16914,N_16955);
or U17031 (N_17031,N_16892,N_16997);
nand U17032 (N_17032,N_16986,N_16820);
nand U17033 (N_17033,N_16878,N_16984);
nor U17034 (N_17034,N_16896,N_16927);
nor U17035 (N_17035,N_16975,N_16940);
or U17036 (N_17036,N_16809,N_16959);
and U17037 (N_17037,N_16841,N_16906);
nand U17038 (N_17038,N_16982,N_16871);
or U17039 (N_17039,N_16832,N_16838);
xor U17040 (N_17040,N_16815,N_16822);
nand U17041 (N_17041,N_16840,N_16980);
or U17042 (N_17042,N_16872,N_16895);
nor U17043 (N_17043,N_16880,N_16852);
xor U17044 (N_17044,N_16836,N_16958);
and U17045 (N_17045,N_16988,N_16891);
and U17046 (N_17046,N_16943,N_16803);
or U17047 (N_17047,N_16916,N_16817);
xnor U17048 (N_17048,N_16952,N_16932);
and U17049 (N_17049,N_16972,N_16992);
nand U17050 (N_17050,N_16846,N_16879);
or U17051 (N_17051,N_16920,N_16867);
nor U17052 (N_17052,N_16985,N_16859);
nand U17053 (N_17053,N_16864,N_16912);
or U17054 (N_17054,N_16885,N_16801);
nand U17055 (N_17055,N_16853,N_16889);
nand U17056 (N_17056,N_16983,N_16995);
and U17057 (N_17057,N_16941,N_16811);
nor U17058 (N_17058,N_16991,N_16994);
xor U17059 (N_17059,N_16802,N_16979);
xor U17060 (N_17060,N_16843,N_16870);
xnor U17061 (N_17061,N_16899,N_16826);
xor U17062 (N_17062,N_16950,N_16931);
and U17063 (N_17063,N_16873,N_16944);
xnor U17064 (N_17064,N_16839,N_16989);
nor U17065 (N_17065,N_16909,N_16960);
and U17066 (N_17066,N_16847,N_16902);
and U17067 (N_17067,N_16821,N_16877);
and U17068 (N_17068,N_16816,N_16921);
nor U17069 (N_17069,N_16861,N_16908);
nand U17070 (N_17070,N_16868,N_16903);
or U17071 (N_17071,N_16897,N_16923);
and U17072 (N_17072,N_16966,N_16907);
nor U17073 (N_17073,N_16887,N_16933);
nor U17074 (N_17074,N_16956,N_16990);
xnor U17075 (N_17075,N_16965,N_16844);
nand U17076 (N_17076,N_16883,N_16863);
nor U17077 (N_17077,N_16874,N_16993);
nor U17078 (N_17078,N_16810,N_16942);
nor U17079 (N_17079,N_16827,N_16935);
xnor U17080 (N_17080,N_16818,N_16849);
nor U17081 (N_17081,N_16884,N_16898);
or U17082 (N_17082,N_16919,N_16835);
xor U17083 (N_17083,N_16876,N_16824);
or U17084 (N_17084,N_16969,N_16882);
xnor U17085 (N_17085,N_16937,N_16830);
xor U17086 (N_17086,N_16949,N_16862);
xnor U17087 (N_17087,N_16854,N_16987);
xor U17088 (N_17088,N_16805,N_16855);
and U17089 (N_17089,N_16929,N_16981);
xnor U17090 (N_17090,N_16837,N_16926);
nand U17091 (N_17091,N_16875,N_16978);
nor U17092 (N_17092,N_16936,N_16953);
or U17093 (N_17093,N_16886,N_16915);
nand U17094 (N_17094,N_16857,N_16828);
nand U17095 (N_17095,N_16922,N_16813);
nand U17096 (N_17096,N_16900,N_16974);
nand U17097 (N_17097,N_16946,N_16834);
xnor U17098 (N_17098,N_16904,N_16967);
xor U17099 (N_17099,N_16888,N_16865);
nand U17100 (N_17100,N_16847,N_16836);
nor U17101 (N_17101,N_16952,N_16865);
xor U17102 (N_17102,N_16970,N_16895);
nand U17103 (N_17103,N_16999,N_16937);
and U17104 (N_17104,N_16842,N_16873);
xnor U17105 (N_17105,N_16832,N_16943);
and U17106 (N_17106,N_16953,N_16966);
and U17107 (N_17107,N_16979,N_16871);
nand U17108 (N_17108,N_16988,N_16859);
and U17109 (N_17109,N_16975,N_16858);
or U17110 (N_17110,N_16944,N_16916);
nand U17111 (N_17111,N_16958,N_16866);
or U17112 (N_17112,N_16966,N_16806);
xnor U17113 (N_17113,N_16924,N_16845);
nor U17114 (N_17114,N_16930,N_16823);
and U17115 (N_17115,N_16959,N_16982);
nor U17116 (N_17116,N_16836,N_16942);
xor U17117 (N_17117,N_16900,N_16967);
and U17118 (N_17118,N_16851,N_16821);
and U17119 (N_17119,N_16994,N_16837);
nand U17120 (N_17120,N_16997,N_16942);
xnor U17121 (N_17121,N_16863,N_16966);
nor U17122 (N_17122,N_16858,N_16964);
and U17123 (N_17123,N_16834,N_16838);
xor U17124 (N_17124,N_16828,N_16968);
and U17125 (N_17125,N_16914,N_16942);
xnor U17126 (N_17126,N_16850,N_16906);
or U17127 (N_17127,N_16885,N_16959);
or U17128 (N_17128,N_16883,N_16881);
nand U17129 (N_17129,N_16890,N_16800);
nand U17130 (N_17130,N_16978,N_16902);
nand U17131 (N_17131,N_16802,N_16916);
nor U17132 (N_17132,N_16869,N_16966);
or U17133 (N_17133,N_16841,N_16805);
or U17134 (N_17134,N_16839,N_16834);
or U17135 (N_17135,N_16921,N_16932);
and U17136 (N_17136,N_16851,N_16933);
nor U17137 (N_17137,N_16905,N_16927);
nand U17138 (N_17138,N_16854,N_16802);
or U17139 (N_17139,N_16964,N_16874);
or U17140 (N_17140,N_16949,N_16885);
and U17141 (N_17141,N_16916,N_16825);
nor U17142 (N_17142,N_16902,N_16883);
xor U17143 (N_17143,N_16816,N_16913);
and U17144 (N_17144,N_16948,N_16824);
xor U17145 (N_17145,N_16890,N_16879);
nor U17146 (N_17146,N_16882,N_16936);
nor U17147 (N_17147,N_16845,N_16855);
or U17148 (N_17148,N_16847,N_16892);
nand U17149 (N_17149,N_16820,N_16936);
xor U17150 (N_17150,N_16913,N_16898);
and U17151 (N_17151,N_16904,N_16947);
nand U17152 (N_17152,N_16962,N_16923);
xnor U17153 (N_17153,N_16847,N_16801);
nor U17154 (N_17154,N_16951,N_16893);
nand U17155 (N_17155,N_16859,N_16931);
xor U17156 (N_17156,N_16845,N_16951);
nor U17157 (N_17157,N_16824,N_16905);
xnor U17158 (N_17158,N_16820,N_16867);
nor U17159 (N_17159,N_16902,N_16996);
or U17160 (N_17160,N_16875,N_16995);
nand U17161 (N_17161,N_16994,N_16946);
nand U17162 (N_17162,N_16960,N_16827);
nor U17163 (N_17163,N_16909,N_16976);
nor U17164 (N_17164,N_16907,N_16965);
nor U17165 (N_17165,N_16853,N_16833);
and U17166 (N_17166,N_16965,N_16841);
xnor U17167 (N_17167,N_16989,N_16837);
nand U17168 (N_17168,N_16806,N_16877);
nor U17169 (N_17169,N_16923,N_16860);
nor U17170 (N_17170,N_16802,N_16849);
nor U17171 (N_17171,N_16869,N_16968);
and U17172 (N_17172,N_16903,N_16901);
and U17173 (N_17173,N_16840,N_16841);
and U17174 (N_17174,N_16909,N_16856);
or U17175 (N_17175,N_16984,N_16939);
xor U17176 (N_17176,N_16981,N_16853);
nand U17177 (N_17177,N_16874,N_16881);
xor U17178 (N_17178,N_16975,N_16931);
nand U17179 (N_17179,N_16936,N_16871);
nor U17180 (N_17180,N_16991,N_16855);
nor U17181 (N_17181,N_16866,N_16975);
nand U17182 (N_17182,N_16967,N_16910);
nand U17183 (N_17183,N_16944,N_16930);
and U17184 (N_17184,N_16962,N_16842);
or U17185 (N_17185,N_16988,N_16870);
nor U17186 (N_17186,N_16863,N_16905);
and U17187 (N_17187,N_16825,N_16814);
xor U17188 (N_17188,N_16863,N_16972);
nor U17189 (N_17189,N_16881,N_16814);
nand U17190 (N_17190,N_16878,N_16910);
nand U17191 (N_17191,N_16949,N_16829);
nor U17192 (N_17192,N_16927,N_16968);
and U17193 (N_17193,N_16918,N_16901);
and U17194 (N_17194,N_16888,N_16920);
xor U17195 (N_17195,N_16962,N_16831);
or U17196 (N_17196,N_16876,N_16883);
or U17197 (N_17197,N_16974,N_16806);
nor U17198 (N_17198,N_16803,N_16940);
nor U17199 (N_17199,N_16986,N_16980);
or U17200 (N_17200,N_17166,N_17107);
or U17201 (N_17201,N_17079,N_17196);
nand U17202 (N_17202,N_17130,N_17119);
or U17203 (N_17203,N_17188,N_17164);
xor U17204 (N_17204,N_17105,N_17123);
and U17205 (N_17205,N_17121,N_17090);
nand U17206 (N_17206,N_17135,N_17124);
and U17207 (N_17207,N_17026,N_17020);
or U17208 (N_17208,N_17093,N_17138);
or U17209 (N_17209,N_17070,N_17127);
and U17210 (N_17210,N_17142,N_17055);
nor U17211 (N_17211,N_17024,N_17167);
nand U17212 (N_17212,N_17106,N_17193);
or U17213 (N_17213,N_17038,N_17081);
nand U17214 (N_17214,N_17054,N_17080);
and U17215 (N_17215,N_17157,N_17012);
xor U17216 (N_17216,N_17045,N_17047);
nand U17217 (N_17217,N_17061,N_17134);
or U17218 (N_17218,N_17066,N_17027);
nor U17219 (N_17219,N_17168,N_17013);
and U17220 (N_17220,N_17153,N_17062);
or U17221 (N_17221,N_17161,N_17109);
xor U17222 (N_17222,N_17056,N_17165);
xnor U17223 (N_17223,N_17190,N_17139);
xor U17224 (N_17224,N_17098,N_17175);
xor U17225 (N_17225,N_17001,N_17178);
or U17226 (N_17226,N_17091,N_17085);
or U17227 (N_17227,N_17100,N_17075);
or U17228 (N_17228,N_17143,N_17008);
xnor U17229 (N_17229,N_17073,N_17156);
xnor U17230 (N_17230,N_17071,N_17154);
nor U17231 (N_17231,N_17034,N_17010);
nand U17232 (N_17232,N_17177,N_17197);
xor U17233 (N_17233,N_17078,N_17144);
or U17234 (N_17234,N_17040,N_17069);
xnor U17235 (N_17235,N_17112,N_17043);
or U17236 (N_17236,N_17033,N_17087);
xnor U17237 (N_17237,N_17060,N_17067);
or U17238 (N_17238,N_17160,N_17110);
and U17239 (N_17239,N_17111,N_17115);
or U17240 (N_17240,N_17184,N_17152);
and U17241 (N_17241,N_17016,N_17006);
nor U17242 (N_17242,N_17023,N_17037);
or U17243 (N_17243,N_17129,N_17159);
xor U17244 (N_17244,N_17031,N_17132);
and U17245 (N_17245,N_17120,N_17053);
or U17246 (N_17246,N_17131,N_17064);
and U17247 (N_17247,N_17113,N_17051);
or U17248 (N_17248,N_17074,N_17155);
nor U17249 (N_17249,N_17048,N_17147);
or U17250 (N_17250,N_17097,N_17007);
nor U17251 (N_17251,N_17171,N_17095);
and U17252 (N_17252,N_17005,N_17102);
or U17253 (N_17253,N_17189,N_17174);
nand U17254 (N_17254,N_17015,N_17163);
nand U17255 (N_17255,N_17028,N_17068);
nand U17256 (N_17256,N_17185,N_17141);
or U17257 (N_17257,N_17199,N_17052);
and U17258 (N_17258,N_17150,N_17019);
and U17259 (N_17259,N_17088,N_17137);
nor U17260 (N_17260,N_17004,N_17118);
and U17261 (N_17261,N_17140,N_17181);
nor U17262 (N_17262,N_17072,N_17101);
nor U17263 (N_17263,N_17186,N_17114);
nor U17264 (N_17264,N_17036,N_17032);
and U17265 (N_17265,N_17116,N_17059);
xor U17266 (N_17266,N_17162,N_17044);
or U17267 (N_17267,N_17050,N_17099);
nor U17268 (N_17268,N_17022,N_17018);
xnor U17269 (N_17269,N_17146,N_17176);
xor U17270 (N_17270,N_17041,N_17092);
or U17271 (N_17271,N_17003,N_17002);
xor U17272 (N_17272,N_17082,N_17096);
nand U17273 (N_17273,N_17117,N_17145);
and U17274 (N_17274,N_17057,N_17058);
xnor U17275 (N_17275,N_17133,N_17046);
xor U17276 (N_17276,N_17094,N_17084);
or U17277 (N_17277,N_17182,N_17187);
nor U17278 (N_17278,N_17014,N_17029);
or U17279 (N_17279,N_17025,N_17170);
nor U17280 (N_17280,N_17042,N_17049);
nand U17281 (N_17281,N_17035,N_17030);
or U17282 (N_17282,N_17000,N_17148);
or U17283 (N_17283,N_17017,N_17172);
nand U17284 (N_17284,N_17136,N_17076);
nand U17285 (N_17285,N_17128,N_17009);
nand U17286 (N_17286,N_17149,N_17183);
nand U17287 (N_17287,N_17039,N_17065);
nor U17288 (N_17288,N_17198,N_17180);
and U17289 (N_17289,N_17011,N_17195);
xor U17290 (N_17290,N_17191,N_17077);
xnor U17291 (N_17291,N_17089,N_17126);
or U17292 (N_17292,N_17108,N_17021);
or U17293 (N_17293,N_17158,N_17194);
or U17294 (N_17294,N_17125,N_17179);
nor U17295 (N_17295,N_17169,N_17063);
nor U17296 (N_17296,N_17086,N_17103);
xor U17297 (N_17297,N_17192,N_17104);
xor U17298 (N_17298,N_17151,N_17173);
and U17299 (N_17299,N_17083,N_17122);
and U17300 (N_17300,N_17078,N_17188);
nor U17301 (N_17301,N_17066,N_17019);
or U17302 (N_17302,N_17185,N_17023);
and U17303 (N_17303,N_17106,N_17039);
xor U17304 (N_17304,N_17165,N_17130);
xor U17305 (N_17305,N_17109,N_17103);
nor U17306 (N_17306,N_17043,N_17034);
xor U17307 (N_17307,N_17159,N_17141);
nor U17308 (N_17308,N_17184,N_17165);
or U17309 (N_17309,N_17041,N_17068);
xor U17310 (N_17310,N_17108,N_17128);
nor U17311 (N_17311,N_17122,N_17103);
nor U17312 (N_17312,N_17135,N_17046);
xor U17313 (N_17313,N_17145,N_17049);
nor U17314 (N_17314,N_17074,N_17001);
and U17315 (N_17315,N_17041,N_17013);
and U17316 (N_17316,N_17099,N_17074);
and U17317 (N_17317,N_17138,N_17143);
nand U17318 (N_17318,N_17194,N_17135);
and U17319 (N_17319,N_17082,N_17195);
nor U17320 (N_17320,N_17073,N_17001);
xnor U17321 (N_17321,N_17112,N_17110);
or U17322 (N_17322,N_17092,N_17195);
nor U17323 (N_17323,N_17111,N_17171);
and U17324 (N_17324,N_17178,N_17152);
nor U17325 (N_17325,N_17177,N_17067);
nor U17326 (N_17326,N_17108,N_17058);
xnor U17327 (N_17327,N_17017,N_17083);
nand U17328 (N_17328,N_17179,N_17184);
and U17329 (N_17329,N_17120,N_17079);
xnor U17330 (N_17330,N_17045,N_17053);
xor U17331 (N_17331,N_17142,N_17010);
or U17332 (N_17332,N_17197,N_17045);
nor U17333 (N_17333,N_17005,N_17112);
nand U17334 (N_17334,N_17152,N_17086);
xnor U17335 (N_17335,N_17150,N_17001);
or U17336 (N_17336,N_17184,N_17079);
xor U17337 (N_17337,N_17058,N_17052);
nand U17338 (N_17338,N_17087,N_17047);
nor U17339 (N_17339,N_17174,N_17111);
xnor U17340 (N_17340,N_17083,N_17185);
and U17341 (N_17341,N_17080,N_17030);
nand U17342 (N_17342,N_17188,N_17170);
and U17343 (N_17343,N_17084,N_17000);
nand U17344 (N_17344,N_17113,N_17160);
nand U17345 (N_17345,N_17088,N_17180);
xnor U17346 (N_17346,N_17153,N_17163);
nand U17347 (N_17347,N_17086,N_17066);
and U17348 (N_17348,N_17004,N_17166);
xnor U17349 (N_17349,N_17184,N_17167);
or U17350 (N_17350,N_17131,N_17018);
or U17351 (N_17351,N_17035,N_17012);
nand U17352 (N_17352,N_17075,N_17179);
and U17353 (N_17353,N_17189,N_17086);
or U17354 (N_17354,N_17017,N_17152);
or U17355 (N_17355,N_17104,N_17026);
and U17356 (N_17356,N_17138,N_17051);
xnor U17357 (N_17357,N_17189,N_17092);
nor U17358 (N_17358,N_17130,N_17173);
nand U17359 (N_17359,N_17188,N_17070);
and U17360 (N_17360,N_17102,N_17194);
nor U17361 (N_17361,N_17057,N_17076);
xnor U17362 (N_17362,N_17106,N_17036);
and U17363 (N_17363,N_17161,N_17187);
nor U17364 (N_17364,N_17017,N_17023);
and U17365 (N_17365,N_17185,N_17159);
nand U17366 (N_17366,N_17103,N_17102);
and U17367 (N_17367,N_17101,N_17074);
xor U17368 (N_17368,N_17194,N_17059);
and U17369 (N_17369,N_17065,N_17014);
or U17370 (N_17370,N_17179,N_17113);
nor U17371 (N_17371,N_17188,N_17084);
xnor U17372 (N_17372,N_17016,N_17115);
nand U17373 (N_17373,N_17145,N_17191);
or U17374 (N_17374,N_17050,N_17075);
nor U17375 (N_17375,N_17171,N_17130);
nor U17376 (N_17376,N_17113,N_17029);
nand U17377 (N_17377,N_17019,N_17073);
nand U17378 (N_17378,N_17093,N_17043);
nor U17379 (N_17379,N_17150,N_17195);
and U17380 (N_17380,N_17167,N_17037);
or U17381 (N_17381,N_17061,N_17172);
nor U17382 (N_17382,N_17012,N_17188);
or U17383 (N_17383,N_17121,N_17174);
xor U17384 (N_17384,N_17084,N_17085);
nand U17385 (N_17385,N_17034,N_17038);
xnor U17386 (N_17386,N_17171,N_17173);
and U17387 (N_17387,N_17108,N_17130);
xor U17388 (N_17388,N_17198,N_17187);
or U17389 (N_17389,N_17029,N_17184);
nand U17390 (N_17390,N_17073,N_17003);
nor U17391 (N_17391,N_17014,N_17159);
and U17392 (N_17392,N_17018,N_17142);
and U17393 (N_17393,N_17044,N_17114);
or U17394 (N_17394,N_17157,N_17010);
xor U17395 (N_17395,N_17179,N_17010);
or U17396 (N_17396,N_17108,N_17094);
or U17397 (N_17397,N_17041,N_17104);
nand U17398 (N_17398,N_17057,N_17124);
nor U17399 (N_17399,N_17121,N_17085);
or U17400 (N_17400,N_17243,N_17311);
nand U17401 (N_17401,N_17202,N_17397);
nor U17402 (N_17402,N_17246,N_17223);
nor U17403 (N_17403,N_17391,N_17285);
or U17404 (N_17404,N_17253,N_17324);
nand U17405 (N_17405,N_17353,N_17388);
and U17406 (N_17406,N_17333,N_17350);
nor U17407 (N_17407,N_17277,N_17357);
nand U17408 (N_17408,N_17205,N_17245);
xnor U17409 (N_17409,N_17371,N_17234);
xnor U17410 (N_17410,N_17326,N_17259);
xor U17411 (N_17411,N_17295,N_17222);
xor U17412 (N_17412,N_17332,N_17384);
nor U17413 (N_17413,N_17323,N_17375);
or U17414 (N_17414,N_17322,N_17329);
and U17415 (N_17415,N_17352,N_17211);
nor U17416 (N_17416,N_17225,N_17301);
and U17417 (N_17417,N_17292,N_17242);
or U17418 (N_17418,N_17283,N_17341);
nand U17419 (N_17419,N_17227,N_17201);
xnor U17420 (N_17420,N_17248,N_17380);
and U17421 (N_17421,N_17215,N_17304);
and U17422 (N_17422,N_17263,N_17256);
or U17423 (N_17423,N_17296,N_17280);
xnor U17424 (N_17424,N_17385,N_17254);
xor U17425 (N_17425,N_17374,N_17214);
and U17426 (N_17426,N_17340,N_17233);
xnor U17427 (N_17427,N_17349,N_17290);
nand U17428 (N_17428,N_17210,N_17393);
or U17429 (N_17429,N_17230,N_17203);
nand U17430 (N_17430,N_17213,N_17212);
nor U17431 (N_17431,N_17276,N_17273);
nand U17432 (N_17432,N_17370,N_17232);
nor U17433 (N_17433,N_17221,N_17217);
or U17434 (N_17434,N_17267,N_17330);
xnor U17435 (N_17435,N_17297,N_17251);
or U17436 (N_17436,N_17342,N_17313);
nor U17437 (N_17437,N_17284,N_17351);
and U17438 (N_17438,N_17338,N_17339);
nand U17439 (N_17439,N_17300,N_17231);
and U17440 (N_17440,N_17207,N_17237);
or U17441 (N_17441,N_17265,N_17200);
xnor U17442 (N_17442,N_17373,N_17383);
xnor U17443 (N_17443,N_17318,N_17281);
and U17444 (N_17444,N_17268,N_17319);
or U17445 (N_17445,N_17278,N_17238);
and U17446 (N_17446,N_17316,N_17365);
xnor U17447 (N_17447,N_17347,N_17293);
nor U17448 (N_17448,N_17379,N_17275);
nand U17449 (N_17449,N_17274,N_17343);
and U17450 (N_17450,N_17307,N_17264);
nand U17451 (N_17451,N_17291,N_17286);
nor U17452 (N_17452,N_17239,N_17229);
and U17453 (N_17453,N_17315,N_17261);
xnor U17454 (N_17454,N_17369,N_17204);
and U17455 (N_17455,N_17255,N_17389);
and U17456 (N_17456,N_17390,N_17216);
or U17457 (N_17457,N_17226,N_17219);
nand U17458 (N_17458,N_17348,N_17364);
and U17459 (N_17459,N_17327,N_17247);
nor U17460 (N_17460,N_17312,N_17337);
nor U17461 (N_17461,N_17335,N_17208);
or U17462 (N_17462,N_17331,N_17310);
nand U17463 (N_17463,N_17314,N_17320);
nor U17464 (N_17464,N_17334,N_17382);
xor U17465 (N_17465,N_17354,N_17321);
nand U17466 (N_17466,N_17303,N_17363);
nor U17467 (N_17467,N_17252,N_17308);
nand U17468 (N_17468,N_17386,N_17346);
nor U17469 (N_17469,N_17269,N_17366);
and U17470 (N_17470,N_17240,N_17355);
nor U17471 (N_17471,N_17362,N_17361);
or U17472 (N_17472,N_17396,N_17317);
xor U17473 (N_17473,N_17209,N_17395);
nor U17474 (N_17474,N_17294,N_17241);
or U17475 (N_17475,N_17378,N_17289);
xnor U17476 (N_17476,N_17262,N_17398);
and U17477 (N_17477,N_17360,N_17367);
or U17478 (N_17478,N_17270,N_17271);
xnor U17479 (N_17479,N_17356,N_17266);
nand U17480 (N_17480,N_17260,N_17387);
nand U17481 (N_17481,N_17358,N_17306);
nand U17482 (N_17482,N_17372,N_17381);
or U17483 (N_17483,N_17392,N_17250);
or U17484 (N_17484,N_17279,N_17359);
xor U17485 (N_17485,N_17328,N_17228);
xnor U17486 (N_17486,N_17218,N_17345);
and U17487 (N_17487,N_17220,N_17272);
or U17488 (N_17488,N_17305,N_17377);
or U17489 (N_17489,N_17288,N_17282);
nor U17490 (N_17490,N_17206,N_17249);
and U17491 (N_17491,N_17344,N_17298);
xnor U17492 (N_17492,N_17236,N_17258);
or U17493 (N_17493,N_17368,N_17336);
or U17494 (N_17494,N_17376,N_17302);
nand U17495 (N_17495,N_17287,N_17325);
nand U17496 (N_17496,N_17299,N_17394);
xor U17497 (N_17497,N_17224,N_17244);
and U17498 (N_17498,N_17399,N_17257);
xnor U17499 (N_17499,N_17309,N_17235);
and U17500 (N_17500,N_17286,N_17303);
nand U17501 (N_17501,N_17309,N_17231);
nor U17502 (N_17502,N_17394,N_17371);
nand U17503 (N_17503,N_17357,N_17231);
nand U17504 (N_17504,N_17365,N_17241);
nand U17505 (N_17505,N_17298,N_17288);
nor U17506 (N_17506,N_17387,N_17297);
nand U17507 (N_17507,N_17398,N_17249);
nor U17508 (N_17508,N_17275,N_17383);
or U17509 (N_17509,N_17369,N_17340);
or U17510 (N_17510,N_17368,N_17323);
xor U17511 (N_17511,N_17296,N_17382);
or U17512 (N_17512,N_17328,N_17334);
nand U17513 (N_17513,N_17324,N_17223);
or U17514 (N_17514,N_17361,N_17318);
nor U17515 (N_17515,N_17211,N_17372);
and U17516 (N_17516,N_17317,N_17300);
or U17517 (N_17517,N_17343,N_17394);
xor U17518 (N_17518,N_17222,N_17320);
xnor U17519 (N_17519,N_17321,N_17255);
nor U17520 (N_17520,N_17207,N_17206);
and U17521 (N_17521,N_17380,N_17250);
or U17522 (N_17522,N_17235,N_17355);
xnor U17523 (N_17523,N_17269,N_17263);
xnor U17524 (N_17524,N_17248,N_17302);
nor U17525 (N_17525,N_17277,N_17327);
nand U17526 (N_17526,N_17350,N_17281);
xor U17527 (N_17527,N_17274,N_17285);
xnor U17528 (N_17528,N_17379,N_17207);
nand U17529 (N_17529,N_17374,N_17336);
xnor U17530 (N_17530,N_17345,N_17268);
and U17531 (N_17531,N_17214,N_17332);
or U17532 (N_17532,N_17206,N_17277);
xnor U17533 (N_17533,N_17220,N_17306);
or U17534 (N_17534,N_17205,N_17202);
xnor U17535 (N_17535,N_17343,N_17334);
and U17536 (N_17536,N_17245,N_17378);
and U17537 (N_17537,N_17233,N_17331);
and U17538 (N_17538,N_17384,N_17238);
nand U17539 (N_17539,N_17263,N_17206);
nor U17540 (N_17540,N_17246,N_17208);
nor U17541 (N_17541,N_17392,N_17399);
nand U17542 (N_17542,N_17210,N_17364);
nor U17543 (N_17543,N_17285,N_17330);
and U17544 (N_17544,N_17375,N_17342);
xor U17545 (N_17545,N_17258,N_17329);
xor U17546 (N_17546,N_17283,N_17348);
nor U17547 (N_17547,N_17312,N_17353);
nand U17548 (N_17548,N_17250,N_17340);
xor U17549 (N_17549,N_17362,N_17373);
and U17550 (N_17550,N_17361,N_17232);
nand U17551 (N_17551,N_17377,N_17391);
and U17552 (N_17552,N_17301,N_17305);
xor U17553 (N_17553,N_17204,N_17282);
and U17554 (N_17554,N_17271,N_17243);
nand U17555 (N_17555,N_17244,N_17245);
nor U17556 (N_17556,N_17316,N_17345);
or U17557 (N_17557,N_17282,N_17285);
nor U17558 (N_17558,N_17276,N_17256);
xnor U17559 (N_17559,N_17258,N_17266);
xor U17560 (N_17560,N_17348,N_17222);
xnor U17561 (N_17561,N_17252,N_17229);
nand U17562 (N_17562,N_17218,N_17334);
nor U17563 (N_17563,N_17347,N_17370);
and U17564 (N_17564,N_17292,N_17293);
xor U17565 (N_17565,N_17381,N_17362);
nor U17566 (N_17566,N_17231,N_17312);
and U17567 (N_17567,N_17201,N_17388);
nand U17568 (N_17568,N_17238,N_17229);
xor U17569 (N_17569,N_17330,N_17324);
nand U17570 (N_17570,N_17294,N_17375);
xor U17571 (N_17571,N_17224,N_17293);
or U17572 (N_17572,N_17216,N_17237);
nand U17573 (N_17573,N_17254,N_17395);
nor U17574 (N_17574,N_17282,N_17373);
xor U17575 (N_17575,N_17353,N_17316);
and U17576 (N_17576,N_17273,N_17226);
and U17577 (N_17577,N_17335,N_17398);
and U17578 (N_17578,N_17398,N_17362);
nor U17579 (N_17579,N_17317,N_17202);
or U17580 (N_17580,N_17397,N_17306);
or U17581 (N_17581,N_17229,N_17328);
nand U17582 (N_17582,N_17348,N_17334);
nand U17583 (N_17583,N_17361,N_17252);
xor U17584 (N_17584,N_17261,N_17361);
nor U17585 (N_17585,N_17216,N_17305);
nand U17586 (N_17586,N_17360,N_17382);
or U17587 (N_17587,N_17242,N_17342);
nor U17588 (N_17588,N_17286,N_17360);
xnor U17589 (N_17589,N_17300,N_17299);
xnor U17590 (N_17590,N_17325,N_17237);
xnor U17591 (N_17591,N_17219,N_17356);
and U17592 (N_17592,N_17398,N_17353);
nor U17593 (N_17593,N_17375,N_17387);
and U17594 (N_17594,N_17248,N_17282);
or U17595 (N_17595,N_17335,N_17291);
nor U17596 (N_17596,N_17296,N_17257);
and U17597 (N_17597,N_17304,N_17305);
xnor U17598 (N_17598,N_17336,N_17356);
nand U17599 (N_17599,N_17327,N_17275);
nand U17600 (N_17600,N_17432,N_17482);
xor U17601 (N_17601,N_17586,N_17504);
and U17602 (N_17602,N_17594,N_17506);
or U17603 (N_17603,N_17404,N_17477);
xnor U17604 (N_17604,N_17540,N_17592);
and U17605 (N_17605,N_17416,N_17565);
and U17606 (N_17606,N_17508,N_17555);
or U17607 (N_17607,N_17403,N_17434);
nor U17608 (N_17608,N_17431,N_17512);
or U17609 (N_17609,N_17402,N_17409);
nor U17610 (N_17610,N_17478,N_17552);
and U17611 (N_17611,N_17491,N_17421);
or U17612 (N_17612,N_17442,N_17449);
and U17613 (N_17613,N_17501,N_17452);
nor U17614 (N_17614,N_17572,N_17588);
nor U17615 (N_17615,N_17472,N_17426);
nor U17616 (N_17616,N_17514,N_17439);
xnor U17617 (N_17617,N_17430,N_17495);
and U17618 (N_17618,N_17479,N_17503);
nand U17619 (N_17619,N_17548,N_17597);
nor U17620 (N_17620,N_17575,N_17521);
nor U17621 (N_17621,N_17566,N_17515);
nand U17622 (N_17622,N_17529,N_17446);
or U17623 (N_17623,N_17558,N_17599);
nor U17624 (N_17624,N_17496,N_17522);
and U17625 (N_17625,N_17530,N_17440);
xnor U17626 (N_17626,N_17465,N_17445);
nand U17627 (N_17627,N_17528,N_17436);
nand U17628 (N_17628,N_17435,N_17535);
and U17629 (N_17629,N_17595,N_17580);
nor U17630 (N_17630,N_17450,N_17505);
and U17631 (N_17631,N_17502,N_17533);
or U17632 (N_17632,N_17507,N_17571);
and U17633 (N_17633,N_17547,N_17562);
or U17634 (N_17634,N_17511,N_17466);
nor U17635 (N_17635,N_17567,N_17494);
nand U17636 (N_17636,N_17422,N_17527);
xor U17637 (N_17637,N_17583,N_17568);
or U17638 (N_17638,N_17587,N_17519);
and U17639 (N_17639,N_17490,N_17489);
or U17640 (N_17640,N_17516,N_17590);
and U17641 (N_17641,N_17543,N_17554);
nor U17642 (N_17642,N_17523,N_17471);
xnor U17643 (N_17643,N_17582,N_17425);
or U17644 (N_17644,N_17444,N_17531);
nor U17645 (N_17645,N_17557,N_17589);
nand U17646 (N_17646,N_17406,N_17560);
nor U17647 (N_17647,N_17553,N_17526);
xor U17648 (N_17648,N_17492,N_17462);
or U17649 (N_17649,N_17578,N_17424);
nor U17650 (N_17650,N_17574,N_17497);
or U17651 (N_17651,N_17591,N_17420);
and U17652 (N_17652,N_17538,N_17429);
xnor U17653 (N_17653,N_17455,N_17541);
xor U17654 (N_17654,N_17412,N_17484);
or U17655 (N_17655,N_17534,N_17469);
nor U17656 (N_17656,N_17532,N_17563);
or U17657 (N_17657,N_17498,N_17573);
xnor U17658 (N_17658,N_17546,N_17447);
nand U17659 (N_17659,N_17411,N_17500);
nand U17660 (N_17660,N_17517,N_17437);
or U17661 (N_17661,N_17438,N_17537);
nand U17662 (N_17662,N_17458,N_17414);
nand U17663 (N_17663,N_17577,N_17467);
or U17664 (N_17664,N_17451,N_17464);
or U17665 (N_17665,N_17487,N_17585);
or U17666 (N_17666,N_17542,N_17570);
nor U17667 (N_17667,N_17417,N_17441);
xor U17668 (N_17668,N_17569,N_17493);
xnor U17669 (N_17669,N_17486,N_17423);
xor U17670 (N_17670,N_17524,N_17483);
nor U17671 (N_17671,N_17470,N_17456);
or U17672 (N_17672,N_17549,N_17457);
xor U17673 (N_17673,N_17481,N_17405);
and U17674 (N_17674,N_17485,N_17453);
xnor U17675 (N_17675,N_17556,N_17539);
or U17676 (N_17676,N_17475,N_17550);
nand U17677 (N_17677,N_17443,N_17520);
nor U17678 (N_17678,N_17480,N_17561);
or U17679 (N_17679,N_17415,N_17459);
nand U17680 (N_17680,N_17545,N_17448);
or U17681 (N_17681,N_17473,N_17581);
nor U17682 (N_17682,N_17513,N_17401);
nand U17683 (N_17683,N_17463,N_17418);
xor U17684 (N_17684,N_17536,N_17407);
nand U17685 (N_17685,N_17400,N_17584);
nand U17686 (N_17686,N_17410,N_17525);
xor U17687 (N_17687,N_17596,N_17576);
nor U17688 (N_17688,N_17510,N_17551);
nand U17689 (N_17689,N_17544,N_17433);
nand U17690 (N_17690,N_17598,N_17427);
nor U17691 (N_17691,N_17461,N_17559);
and U17692 (N_17692,N_17454,N_17419);
or U17693 (N_17693,N_17488,N_17593);
nor U17694 (N_17694,N_17564,N_17509);
nand U17695 (N_17695,N_17460,N_17428);
nor U17696 (N_17696,N_17468,N_17408);
nand U17697 (N_17697,N_17413,N_17518);
xor U17698 (N_17698,N_17476,N_17499);
xnor U17699 (N_17699,N_17474,N_17579);
xnor U17700 (N_17700,N_17557,N_17540);
nor U17701 (N_17701,N_17450,N_17575);
nor U17702 (N_17702,N_17405,N_17514);
or U17703 (N_17703,N_17595,N_17471);
xnor U17704 (N_17704,N_17513,N_17483);
and U17705 (N_17705,N_17414,N_17460);
and U17706 (N_17706,N_17576,N_17516);
xnor U17707 (N_17707,N_17476,N_17430);
and U17708 (N_17708,N_17501,N_17426);
nor U17709 (N_17709,N_17489,N_17534);
nor U17710 (N_17710,N_17598,N_17447);
and U17711 (N_17711,N_17435,N_17584);
or U17712 (N_17712,N_17585,N_17418);
or U17713 (N_17713,N_17522,N_17404);
or U17714 (N_17714,N_17408,N_17557);
or U17715 (N_17715,N_17574,N_17468);
nor U17716 (N_17716,N_17416,N_17403);
and U17717 (N_17717,N_17503,N_17554);
and U17718 (N_17718,N_17455,N_17473);
and U17719 (N_17719,N_17491,N_17532);
and U17720 (N_17720,N_17474,N_17537);
nor U17721 (N_17721,N_17478,N_17437);
or U17722 (N_17722,N_17526,N_17536);
or U17723 (N_17723,N_17579,N_17595);
nor U17724 (N_17724,N_17556,N_17472);
xor U17725 (N_17725,N_17457,N_17497);
nor U17726 (N_17726,N_17509,N_17491);
nand U17727 (N_17727,N_17508,N_17452);
or U17728 (N_17728,N_17553,N_17515);
nor U17729 (N_17729,N_17433,N_17446);
xnor U17730 (N_17730,N_17421,N_17534);
or U17731 (N_17731,N_17445,N_17488);
nor U17732 (N_17732,N_17592,N_17558);
and U17733 (N_17733,N_17596,N_17439);
and U17734 (N_17734,N_17455,N_17463);
nand U17735 (N_17735,N_17582,N_17501);
or U17736 (N_17736,N_17517,N_17435);
or U17737 (N_17737,N_17478,N_17549);
xnor U17738 (N_17738,N_17524,N_17427);
nand U17739 (N_17739,N_17472,N_17432);
and U17740 (N_17740,N_17429,N_17500);
nor U17741 (N_17741,N_17527,N_17523);
and U17742 (N_17742,N_17554,N_17456);
xnor U17743 (N_17743,N_17417,N_17550);
nor U17744 (N_17744,N_17568,N_17559);
nor U17745 (N_17745,N_17401,N_17432);
xor U17746 (N_17746,N_17489,N_17512);
xor U17747 (N_17747,N_17530,N_17529);
xor U17748 (N_17748,N_17454,N_17453);
nor U17749 (N_17749,N_17518,N_17415);
nor U17750 (N_17750,N_17472,N_17478);
nand U17751 (N_17751,N_17444,N_17593);
xor U17752 (N_17752,N_17508,N_17445);
and U17753 (N_17753,N_17416,N_17462);
nand U17754 (N_17754,N_17508,N_17540);
nor U17755 (N_17755,N_17437,N_17549);
nand U17756 (N_17756,N_17520,N_17414);
and U17757 (N_17757,N_17403,N_17471);
and U17758 (N_17758,N_17577,N_17472);
and U17759 (N_17759,N_17452,N_17486);
and U17760 (N_17760,N_17591,N_17538);
nand U17761 (N_17761,N_17467,N_17455);
xnor U17762 (N_17762,N_17581,N_17422);
xnor U17763 (N_17763,N_17531,N_17519);
and U17764 (N_17764,N_17447,N_17406);
xor U17765 (N_17765,N_17557,N_17566);
nor U17766 (N_17766,N_17401,N_17596);
or U17767 (N_17767,N_17420,N_17544);
or U17768 (N_17768,N_17416,N_17400);
nor U17769 (N_17769,N_17588,N_17579);
and U17770 (N_17770,N_17550,N_17431);
nand U17771 (N_17771,N_17476,N_17535);
nand U17772 (N_17772,N_17428,N_17528);
nor U17773 (N_17773,N_17533,N_17559);
nor U17774 (N_17774,N_17439,N_17478);
nor U17775 (N_17775,N_17521,N_17504);
nor U17776 (N_17776,N_17534,N_17448);
and U17777 (N_17777,N_17597,N_17523);
and U17778 (N_17778,N_17585,N_17552);
nor U17779 (N_17779,N_17495,N_17477);
nand U17780 (N_17780,N_17439,N_17457);
and U17781 (N_17781,N_17538,N_17417);
or U17782 (N_17782,N_17586,N_17555);
nor U17783 (N_17783,N_17488,N_17416);
nor U17784 (N_17784,N_17512,N_17569);
xnor U17785 (N_17785,N_17581,N_17442);
nor U17786 (N_17786,N_17527,N_17489);
or U17787 (N_17787,N_17465,N_17536);
and U17788 (N_17788,N_17512,N_17416);
nor U17789 (N_17789,N_17413,N_17489);
xor U17790 (N_17790,N_17487,N_17565);
and U17791 (N_17791,N_17400,N_17532);
nand U17792 (N_17792,N_17449,N_17495);
nand U17793 (N_17793,N_17519,N_17530);
or U17794 (N_17794,N_17494,N_17551);
or U17795 (N_17795,N_17521,N_17513);
xnor U17796 (N_17796,N_17408,N_17528);
xnor U17797 (N_17797,N_17520,N_17441);
and U17798 (N_17798,N_17591,N_17559);
nor U17799 (N_17799,N_17579,N_17530);
nand U17800 (N_17800,N_17731,N_17770);
xnor U17801 (N_17801,N_17654,N_17638);
xor U17802 (N_17802,N_17613,N_17675);
or U17803 (N_17803,N_17671,N_17703);
nand U17804 (N_17804,N_17680,N_17683);
nor U17805 (N_17805,N_17601,N_17711);
nand U17806 (N_17806,N_17724,N_17635);
nor U17807 (N_17807,N_17689,N_17722);
and U17808 (N_17808,N_17655,N_17740);
xor U17809 (N_17809,N_17645,N_17648);
or U17810 (N_17810,N_17764,N_17789);
xor U17811 (N_17811,N_17614,N_17743);
nand U17812 (N_17812,N_17765,N_17716);
and U17813 (N_17813,N_17610,N_17657);
and U17814 (N_17814,N_17618,N_17647);
or U17815 (N_17815,N_17785,N_17757);
nor U17816 (N_17816,N_17799,N_17726);
or U17817 (N_17817,N_17631,N_17600);
or U17818 (N_17818,N_17728,N_17623);
or U17819 (N_17819,N_17761,N_17663);
and U17820 (N_17820,N_17606,N_17611);
and U17821 (N_17821,N_17777,N_17685);
nand U17822 (N_17822,N_17696,N_17609);
xnor U17823 (N_17823,N_17629,N_17730);
xnor U17824 (N_17824,N_17619,N_17630);
xnor U17825 (N_17825,N_17769,N_17732);
nor U17826 (N_17826,N_17616,N_17786);
nor U17827 (N_17827,N_17708,N_17646);
xor U17828 (N_17828,N_17604,N_17725);
and U17829 (N_17829,N_17632,N_17795);
and U17830 (N_17830,N_17694,N_17690);
nor U17831 (N_17831,N_17713,N_17622);
nand U17832 (N_17832,N_17603,N_17617);
nand U17833 (N_17833,N_17612,N_17698);
nor U17834 (N_17834,N_17684,N_17772);
xor U17835 (N_17835,N_17776,N_17624);
or U17836 (N_17836,N_17741,N_17715);
xnor U17837 (N_17837,N_17733,N_17681);
or U17838 (N_17838,N_17707,N_17723);
nor U17839 (N_17839,N_17644,N_17710);
nor U17840 (N_17840,N_17780,N_17634);
or U17841 (N_17841,N_17759,N_17650);
xor U17842 (N_17842,N_17674,N_17742);
and U17843 (N_17843,N_17665,N_17745);
nor U17844 (N_17844,N_17760,N_17709);
nor U17845 (N_17845,N_17771,N_17737);
and U17846 (N_17846,N_17640,N_17784);
or U17847 (N_17847,N_17643,N_17686);
nor U17848 (N_17848,N_17693,N_17717);
or U17849 (N_17849,N_17798,N_17656);
and U17850 (N_17850,N_17704,N_17697);
xor U17851 (N_17851,N_17747,N_17651);
nor U17852 (N_17852,N_17779,N_17721);
or U17853 (N_17853,N_17749,N_17636);
and U17854 (N_17854,N_17662,N_17660);
nor U17855 (N_17855,N_17790,N_17627);
xnor U17856 (N_17856,N_17667,N_17673);
nand U17857 (N_17857,N_17677,N_17748);
and U17858 (N_17858,N_17608,N_17672);
nand U17859 (N_17859,N_17637,N_17746);
and U17860 (N_17860,N_17735,N_17718);
nor U17861 (N_17861,N_17767,N_17706);
nand U17862 (N_17862,N_17739,N_17705);
xor U17863 (N_17863,N_17628,N_17688);
nand U17864 (N_17864,N_17756,N_17676);
nor U17865 (N_17865,N_17797,N_17775);
and U17866 (N_17866,N_17758,N_17699);
and U17867 (N_17867,N_17702,N_17620);
or U17868 (N_17868,N_17679,N_17744);
or U17869 (N_17869,N_17727,N_17763);
nor U17870 (N_17870,N_17762,N_17602);
or U17871 (N_17871,N_17753,N_17787);
nor U17872 (N_17872,N_17720,N_17649);
nor U17873 (N_17873,N_17773,N_17712);
nor U17874 (N_17874,N_17621,N_17642);
nand U17875 (N_17875,N_17729,N_17670);
nand U17876 (N_17876,N_17669,N_17754);
or U17877 (N_17877,N_17752,N_17625);
and U17878 (N_17878,N_17666,N_17751);
xnor U17879 (N_17879,N_17641,N_17714);
xnor U17880 (N_17880,N_17788,N_17783);
xnor U17881 (N_17881,N_17778,N_17653);
and U17882 (N_17882,N_17701,N_17652);
nor U17883 (N_17883,N_17678,N_17793);
or U17884 (N_17884,N_17659,N_17792);
and U17885 (N_17885,N_17796,N_17605);
xnor U17886 (N_17886,N_17633,N_17700);
nand U17887 (N_17887,N_17695,N_17687);
or U17888 (N_17888,N_17781,N_17661);
xnor U17889 (N_17889,N_17794,N_17734);
and U17890 (N_17890,N_17774,N_17766);
or U17891 (N_17891,N_17692,N_17639);
nand U17892 (N_17892,N_17607,N_17738);
or U17893 (N_17893,N_17664,N_17736);
or U17894 (N_17894,N_17691,N_17750);
or U17895 (N_17895,N_17755,N_17791);
nor U17896 (N_17896,N_17768,N_17719);
nand U17897 (N_17897,N_17658,N_17626);
or U17898 (N_17898,N_17782,N_17668);
xor U17899 (N_17899,N_17615,N_17682);
and U17900 (N_17900,N_17620,N_17667);
nand U17901 (N_17901,N_17694,N_17677);
nor U17902 (N_17902,N_17643,N_17672);
xnor U17903 (N_17903,N_17796,N_17687);
or U17904 (N_17904,N_17751,N_17693);
and U17905 (N_17905,N_17760,N_17790);
nor U17906 (N_17906,N_17706,N_17635);
nand U17907 (N_17907,N_17652,N_17753);
nand U17908 (N_17908,N_17664,N_17721);
nor U17909 (N_17909,N_17634,N_17686);
or U17910 (N_17910,N_17642,N_17654);
nor U17911 (N_17911,N_17726,N_17719);
or U17912 (N_17912,N_17757,N_17795);
or U17913 (N_17913,N_17726,N_17783);
and U17914 (N_17914,N_17739,N_17685);
nor U17915 (N_17915,N_17779,N_17685);
nand U17916 (N_17916,N_17637,N_17620);
nor U17917 (N_17917,N_17700,N_17749);
nor U17918 (N_17918,N_17603,N_17751);
xnor U17919 (N_17919,N_17623,N_17670);
nand U17920 (N_17920,N_17633,N_17636);
nor U17921 (N_17921,N_17767,N_17778);
nor U17922 (N_17922,N_17630,N_17621);
or U17923 (N_17923,N_17760,N_17770);
and U17924 (N_17924,N_17788,N_17743);
xor U17925 (N_17925,N_17745,N_17631);
nor U17926 (N_17926,N_17688,N_17619);
or U17927 (N_17927,N_17712,N_17731);
and U17928 (N_17928,N_17678,N_17668);
or U17929 (N_17929,N_17758,N_17658);
and U17930 (N_17930,N_17698,N_17736);
and U17931 (N_17931,N_17693,N_17786);
xor U17932 (N_17932,N_17651,N_17748);
and U17933 (N_17933,N_17693,N_17646);
and U17934 (N_17934,N_17725,N_17763);
and U17935 (N_17935,N_17720,N_17659);
nor U17936 (N_17936,N_17609,N_17743);
nor U17937 (N_17937,N_17746,N_17695);
nand U17938 (N_17938,N_17715,N_17722);
xor U17939 (N_17939,N_17675,N_17656);
nor U17940 (N_17940,N_17740,N_17742);
xor U17941 (N_17941,N_17644,N_17709);
and U17942 (N_17942,N_17764,N_17702);
xnor U17943 (N_17943,N_17725,N_17745);
or U17944 (N_17944,N_17724,N_17714);
nand U17945 (N_17945,N_17786,N_17623);
xor U17946 (N_17946,N_17600,N_17793);
nor U17947 (N_17947,N_17646,N_17601);
nand U17948 (N_17948,N_17646,N_17714);
nand U17949 (N_17949,N_17780,N_17686);
xor U17950 (N_17950,N_17763,N_17728);
nor U17951 (N_17951,N_17750,N_17757);
and U17952 (N_17952,N_17667,N_17738);
or U17953 (N_17953,N_17778,N_17647);
and U17954 (N_17954,N_17789,N_17734);
xor U17955 (N_17955,N_17665,N_17742);
and U17956 (N_17956,N_17608,N_17761);
xor U17957 (N_17957,N_17678,N_17720);
and U17958 (N_17958,N_17747,N_17676);
or U17959 (N_17959,N_17697,N_17789);
xnor U17960 (N_17960,N_17694,N_17608);
xor U17961 (N_17961,N_17710,N_17625);
nand U17962 (N_17962,N_17691,N_17705);
nor U17963 (N_17963,N_17782,N_17677);
and U17964 (N_17964,N_17788,N_17675);
or U17965 (N_17965,N_17745,N_17673);
or U17966 (N_17966,N_17601,N_17730);
and U17967 (N_17967,N_17753,N_17609);
nand U17968 (N_17968,N_17737,N_17697);
xnor U17969 (N_17969,N_17754,N_17797);
or U17970 (N_17970,N_17680,N_17686);
and U17971 (N_17971,N_17761,N_17609);
or U17972 (N_17972,N_17695,N_17664);
or U17973 (N_17973,N_17652,N_17671);
or U17974 (N_17974,N_17642,N_17691);
or U17975 (N_17975,N_17690,N_17763);
nor U17976 (N_17976,N_17798,N_17785);
nor U17977 (N_17977,N_17608,N_17639);
xnor U17978 (N_17978,N_17659,N_17641);
xnor U17979 (N_17979,N_17622,N_17767);
or U17980 (N_17980,N_17669,N_17708);
or U17981 (N_17981,N_17602,N_17725);
xor U17982 (N_17982,N_17661,N_17675);
nor U17983 (N_17983,N_17724,N_17766);
nor U17984 (N_17984,N_17600,N_17740);
or U17985 (N_17985,N_17676,N_17626);
or U17986 (N_17986,N_17606,N_17748);
nand U17987 (N_17987,N_17746,N_17608);
xnor U17988 (N_17988,N_17736,N_17682);
or U17989 (N_17989,N_17672,N_17634);
and U17990 (N_17990,N_17784,N_17797);
nand U17991 (N_17991,N_17785,N_17614);
nor U17992 (N_17992,N_17639,N_17791);
and U17993 (N_17993,N_17663,N_17696);
nor U17994 (N_17994,N_17627,N_17658);
and U17995 (N_17995,N_17601,N_17794);
or U17996 (N_17996,N_17772,N_17663);
nand U17997 (N_17997,N_17770,N_17626);
and U17998 (N_17998,N_17696,N_17680);
nor U17999 (N_17999,N_17639,N_17744);
nor U18000 (N_18000,N_17837,N_17805);
and U18001 (N_18001,N_17952,N_17991);
xnor U18002 (N_18002,N_17932,N_17943);
xnor U18003 (N_18003,N_17843,N_17841);
nand U18004 (N_18004,N_17978,N_17910);
nor U18005 (N_18005,N_17875,N_17891);
and U18006 (N_18006,N_17819,N_17925);
xnor U18007 (N_18007,N_17851,N_17833);
xnor U18008 (N_18008,N_17913,N_17901);
or U18009 (N_18009,N_17849,N_17844);
and U18010 (N_18010,N_17908,N_17989);
nand U18011 (N_18011,N_17890,N_17965);
nand U18012 (N_18012,N_17867,N_17853);
and U18013 (N_18013,N_17802,N_17800);
xor U18014 (N_18014,N_17815,N_17895);
or U18015 (N_18015,N_17812,N_17927);
xnor U18016 (N_18016,N_17821,N_17956);
nor U18017 (N_18017,N_17856,N_17988);
or U18018 (N_18018,N_17971,N_17840);
nand U18019 (N_18019,N_17823,N_17864);
nor U18020 (N_18020,N_17889,N_17961);
nand U18021 (N_18021,N_17898,N_17811);
nor U18022 (N_18022,N_17945,N_17957);
and U18023 (N_18023,N_17974,N_17935);
or U18024 (N_18024,N_17924,N_17869);
or U18025 (N_18025,N_17854,N_17983);
or U18026 (N_18026,N_17832,N_17999);
xnor U18027 (N_18027,N_17948,N_17827);
xor U18028 (N_18028,N_17966,N_17953);
and U18029 (N_18029,N_17907,N_17941);
nand U18030 (N_18030,N_17868,N_17960);
and U18031 (N_18031,N_17846,N_17919);
xor U18032 (N_18032,N_17922,N_17835);
and U18033 (N_18033,N_17831,N_17929);
or U18034 (N_18034,N_17950,N_17994);
nor U18035 (N_18035,N_17939,N_17986);
nand U18036 (N_18036,N_17958,N_17933);
nand U18037 (N_18037,N_17938,N_17860);
nor U18038 (N_18038,N_17972,N_17914);
or U18039 (N_18039,N_17818,N_17918);
and U18040 (N_18040,N_17987,N_17970);
nand U18041 (N_18041,N_17981,N_17976);
and U18042 (N_18042,N_17985,N_17858);
nor U18043 (N_18043,N_17877,N_17872);
xor U18044 (N_18044,N_17816,N_17848);
xnor U18045 (N_18045,N_17904,N_17855);
and U18046 (N_18046,N_17969,N_17885);
nand U18047 (N_18047,N_17923,N_17900);
xor U18048 (N_18048,N_17921,N_17808);
and U18049 (N_18049,N_17830,N_17825);
or U18050 (N_18050,N_17906,N_17937);
or U18051 (N_18051,N_17884,N_17809);
or U18052 (N_18052,N_17964,N_17916);
xnor U18053 (N_18053,N_17909,N_17862);
nor U18054 (N_18054,N_17955,N_17917);
xnor U18055 (N_18055,N_17920,N_17828);
nor U18056 (N_18056,N_17801,N_17888);
nor U18057 (N_18057,N_17949,N_17820);
nor U18058 (N_18058,N_17947,N_17813);
and U18059 (N_18059,N_17984,N_17866);
and U18060 (N_18060,N_17881,N_17824);
xnor U18061 (N_18061,N_17940,N_17993);
nor U18062 (N_18062,N_17804,N_17963);
xnor U18063 (N_18063,N_17876,N_17807);
nor U18064 (N_18064,N_17954,N_17902);
and U18065 (N_18065,N_17834,N_17903);
and U18066 (N_18066,N_17896,N_17861);
nor U18067 (N_18067,N_17962,N_17814);
nand U18068 (N_18068,N_17817,N_17865);
nand U18069 (N_18069,N_17873,N_17951);
nor U18070 (N_18070,N_17915,N_17930);
nor U18071 (N_18071,N_17822,N_17911);
and U18072 (N_18072,N_17803,N_17845);
nor U18073 (N_18073,N_17894,N_17806);
and U18074 (N_18074,N_17975,N_17878);
nand U18075 (N_18075,N_17998,N_17946);
nand U18076 (N_18076,N_17944,N_17859);
or U18077 (N_18077,N_17863,N_17931);
xnor U18078 (N_18078,N_17839,N_17942);
nand U18079 (N_18079,N_17871,N_17967);
and U18080 (N_18080,N_17842,N_17979);
xor U18081 (N_18081,N_17934,N_17899);
or U18082 (N_18082,N_17977,N_17829);
nor U18083 (N_18083,N_17912,N_17874);
nor U18084 (N_18084,N_17968,N_17973);
nor U18085 (N_18085,N_17857,N_17980);
or U18086 (N_18086,N_17847,N_17992);
and U18087 (N_18087,N_17850,N_17982);
nor U18088 (N_18088,N_17886,N_17810);
or U18089 (N_18089,N_17995,N_17836);
xor U18090 (N_18090,N_17926,N_17870);
nor U18091 (N_18091,N_17838,N_17905);
xnor U18092 (N_18092,N_17996,N_17959);
nor U18093 (N_18093,N_17826,N_17879);
or U18094 (N_18094,N_17997,N_17892);
nand U18095 (N_18095,N_17852,N_17990);
xnor U18096 (N_18096,N_17880,N_17882);
or U18097 (N_18097,N_17936,N_17887);
or U18098 (N_18098,N_17883,N_17893);
nor U18099 (N_18099,N_17897,N_17928);
xor U18100 (N_18100,N_17914,N_17870);
and U18101 (N_18101,N_17871,N_17989);
or U18102 (N_18102,N_17811,N_17909);
xnor U18103 (N_18103,N_17973,N_17864);
xnor U18104 (N_18104,N_17846,N_17860);
nor U18105 (N_18105,N_17878,N_17943);
nand U18106 (N_18106,N_17875,N_17895);
xor U18107 (N_18107,N_17998,N_17916);
nor U18108 (N_18108,N_17898,N_17896);
or U18109 (N_18109,N_17913,N_17882);
nor U18110 (N_18110,N_17814,N_17832);
or U18111 (N_18111,N_17953,N_17875);
nand U18112 (N_18112,N_17997,N_17903);
nor U18113 (N_18113,N_17979,N_17990);
nor U18114 (N_18114,N_17960,N_17896);
and U18115 (N_18115,N_17977,N_17990);
nor U18116 (N_18116,N_17882,N_17812);
and U18117 (N_18117,N_17999,N_17844);
or U18118 (N_18118,N_17934,N_17952);
nor U18119 (N_18119,N_17820,N_17950);
xor U18120 (N_18120,N_17869,N_17875);
and U18121 (N_18121,N_17985,N_17903);
and U18122 (N_18122,N_17947,N_17885);
or U18123 (N_18123,N_17952,N_17818);
or U18124 (N_18124,N_17875,N_17847);
nor U18125 (N_18125,N_17965,N_17836);
nor U18126 (N_18126,N_17823,N_17869);
nand U18127 (N_18127,N_17861,N_17970);
nor U18128 (N_18128,N_17980,N_17911);
or U18129 (N_18129,N_17985,N_17866);
or U18130 (N_18130,N_17809,N_17955);
xnor U18131 (N_18131,N_17948,N_17976);
nand U18132 (N_18132,N_17880,N_17908);
or U18133 (N_18133,N_17941,N_17802);
and U18134 (N_18134,N_17874,N_17883);
xnor U18135 (N_18135,N_17919,N_17963);
xor U18136 (N_18136,N_17921,N_17879);
nand U18137 (N_18137,N_17903,N_17929);
nand U18138 (N_18138,N_17848,N_17961);
nor U18139 (N_18139,N_17820,N_17804);
nor U18140 (N_18140,N_17806,N_17801);
nand U18141 (N_18141,N_17883,N_17865);
and U18142 (N_18142,N_17945,N_17975);
nor U18143 (N_18143,N_17887,N_17972);
nand U18144 (N_18144,N_17917,N_17996);
and U18145 (N_18145,N_17931,N_17854);
nand U18146 (N_18146,N_17900,N_17884);
nor U18147 (N_18147,N_17915,N_17852);
nor U18148 (N_18148,N_17980,N_17919);
xor U18149 (N_18149,N_17893,N_17882);
xor U18150 (N_18150,N_17832,N_17825);
or U18151 (N_18151,N_17835,N_17969);
xnor U18152 (N_18152,N_17912,N_17831);
and U18153 (N_18153,N_17944,N_17924);
xor U18154 (N_18154,N_17898,N_17954);
or U18155 (N_18155,N_17863,N_17977);
and U18156 (N_18156,N_17925,N_17995);
or U18157 (N_18157,N_17844,N_17878);
xor U18158 (N_18158,N_17903,N_17889);
nor U18159 (N_18159,N_17820,N_17879);
nor U18160 (N_18160,N_17844,N_17915);
or U18161 (N_18161,N_17954,N_17877);
and U18162 (N_18162,N_17809,N_17816);
nand U18163 (N_18163,N_17886,N_17873);
nor U18164 (N_18164,N_17895,N_17835);
nand U18165 (N_18165,N_17972,N_17966);
xnor U18166 (N_18166,N_17874,N_17877);
xnor U18167 (N_18167,N_17949,N_17804);
and U18168 (N_18168,N_17928,N_17830);
xor U18169 (N_18169,N_17887,N_17997);
or U18170 (N_18170,N_17851,N_17919);
xnor U18171 (N_18171,N_17889,N_17872);
xnor U18172 (N_18172,N_17853,N_17933);
nor U18173 (N_18173,N_17947,N_17990);
and U18174 (N_18174,N_17839,N_17987);
or U18175 (N_18175,N_17946,N_17995);
and U18176 (N_18176,N_17969,N_17967);
nand U18177 (N_18177,N_17972,N_17950);
xor U18178 (N_18178,N_17898,N_17876);
nand U18179 (N_18179,N_17999,N_17873);
nand U18180 (N_18180,N_17869,N_17874);
or U18181 (N_18181,N_17888,N_17916);
and U18182 (N_18182,N_17856,N_17995);
nor U18183 (N_18183,N_17894,N_17902);
or U18184 (N_18184,N_17876,N_17877);
nand U18185 (N_18185,N_17932,N_17897);
nor U18186 (N_18186,N_17912,N_17867);
or U18187 (N_18187,N_17848,N_17900);
and U18188 (N_18188,N_17952,N_17979);
or U18189 (N_18189,N_17983,N_17914);
and U18190 (N_18190,N_17900,N_17821);
nor U18191 (N_18191,N_17991,N_17880);
nor U18192 (N_18192,N_17869,N_17980);
nand U18193 (N_18193,N_17974,N_17851);
nor U18194 (N_18194,N_17960,N_17938);
and U18195 (N_18195,N_17909,N_17889);
and U18196 (N_18196,N_17803,N_17967);
nor U18197 (N_18197,N_17817,N_17931);
nor U18198 (N_18198,N_17934,N_17903);
or U18199 (N_18199,N_17913,N_17922);
or U18200 (N_18200,N_18099,N_18026);
xor U18201 (N_18201,N_18098,N_18162);
or U18202 (N_18202,N_18007,N_18020);
and U18203 (N_18203,N_18143,N_18130);
or U18204 (N_18204,N_18166,N_18083);
and U18205 (N_18205,N_18041,N_18113);
and U18206 (N_18206,N_18015,N_18031);
and U18207 (N_18207,N_18006,N_18068);
xor U18208 (N_18208,N_18088,N_18025);
xnor U18209 (N_18209,N_18037,N_18071);
and U18210 (N_18210,N_18029,N_18091);
nand U18211 (N_18211,N_18182,N_18049);
and U18212 (N_18212,N_18161,N_18180);
nor U18213 (N_18213,N_18198,N_18138);
xnor U18214 (N_18214,N_18123,N_18133);
xor U18215 (N_18215,N_18171,N_18117);
or U18216 (N_18216,N_18170,N_18040);
xnor U18217 (N_18217,N_18178,N_18104);
nand U18218 (N_18218,N_18154,N_18080);
nand U18219 (N_18219,N_18101,N_18121);
nor U18220 (N_18220,N_18012,N_18066);
nand U18221 (N_18221,N_18036,N_18057);
xor U18222 (N_18222,N_18077,N_18158);
or U18223 (N_18223,N_18194,N_18100);
nor U18224 (N_18224,N_18055,N_18022);
or U18225 (N_18225,N_18129,N_18043);
or U18226 (N_18226,N_18052,N_18188);
xor U18227 (N_18227,N_18039,N_18109);
nor U18228 (N_18228,N_18134,N_18106);
xnor U18229 (N_18229,N_18008,N_18081);
xor U18230 (N_18230,N_18092,N_18142);
and U18231 (N_18231,N_18046,N_18136);
nor U18232 (N_18232,N_18061,N_18027);
xor U18233 (N_18233,N_18184,N_18102);
and U18234 (N_18234,N_18195,N_18060);
nand U18235 (N_18235,N_18003,N_18193);
and U18236 (N_18236,N_18132,N_18079);
or U18237 (N_18237,N_18119,N_18089);
xor U18238 (N_18238,N_18084,N_18176);
nor U18239 (N_18239,N_18173,N_18145);
xnor U18240 (N_18240,N_18144,N_18017);
nand U18241 (N_18241,N_18141,N_18028);
xor U18242 (N_18242,N_18108,N_18126);
and U18243 (N_18243,N_18069,N_18019);
nor U18244 (N_18244,N_18118,N_18192);
xor U18245 (N_18245,N_18107,N_18160);
nor U18246 (N_18246,N_18151,N_18186);
or U18247 (N_18247,N_18063,N_18018);
or U18248 (N_18248,N_18078,N_18085);
nor U18249 (N_18249,N_18190,N_18168);
nand U18250 (N_18250,N_18010,N_18103);
nand U18251 (N_18251,N_18164,N_18169);
nand U18252 (N_18252,N_18059,N_18075);
and U18253 (N_18253,N_18038,N_18074);
or U18254 (N_18254,N_18096,N_18053);
xor U18255 (N_18255,N_18013,N_18140);
xor U18256 (N_18256,N_18112,N_18120);
xnor U18257 (N_18257,N_18070,N_18127);
or U18258 (N_18258,N_18067,N_18016);
and U18259 (N_18259,N_18175,N_18115);
and U18260 (N_18260,N_18086,N_18034);
or U18261 (N_18261,N_18148,N_18187);
and U18262 (N_18262,N_18087,N_18177);
nand U18263 (N_18263,N_18035,N_18163);
and U18264 (N_18264,N_18023,N_18149);
and U18265 (N_18265,N_18111,N_18181);
xor U18266 (N_18266,N_18153,N_18073);
xnor U18267 (N_18267,N_18097,N_18122);
xnor U18268 (N_18268,N_18128,N_18054);
nor U18269 (N_18269,N_18045,N_18090);
and U18270 (N_18270,N_18021,N_18095);
nor U18271 (N_18271,N_18155,N_18065);
or U18272 (N_18272,N_18179,N_18014);
nand U18273 (N_18273,N_18183,N_18048);
nand U18274 (N_18274,N_18137,N_18146);
and U18275 (N_18275,N_18165,N_18047);
xnor U18276 (N_18276,N_18139,N_18185);
nand U18277 (N_18277,N_18033,N_18110);
or U18278 (N_18278,N_18094,N_18116);
nor U18279 (N_18279,N_18135,N_18032);
xor U18280 (N_18280,N_18114,N_18072);
nor U18281 (N_18281,N_18011,N_18001);
and U18282 (N_18282,N_18159,N_18189);
or U18283 (N_18283,N_18062,N_18147);
nand U18284 (N_18284,N_18042,N_18030);
and U18285 (N_18285,N_18002,N_18191);
and U18286 (N_18286,N_18004,N_18125);
nand U18287 (N_18287,N_18058,N_18005);
xnor U18288 (N_18288,N_18082,N_18076);
and U18289 (N_18289,N_18197,N_18093);
nor U18290 (N_18290,N_18124,N_18167);
and U18291 (N_18291,N_18000,N_18131);
nand U18292 (N_18292,N_18024,N_18174);
nand U18293 (N_18293,N_18051,N_18044);
xor U18294 (N_18294,N_18050,N_18105);
and U18295 (N_18295,N_18156,N_18056);
nor U18296 (N_18296,N_18150,N_18199);
and U18297 (N_18297,N_18064,N_18152);
and U18298 (N_18298,N_18009,N_18172);
xor U18299 (N_18299,N_18196,N_18157);
nand U18300 (N_18300,N_18024,N_18113);
and U18301 (N_18301,N_18017,N_18154);
and U18302 (N_18302,N_18073,N_18048);
or U18303 (N_18303,N_18036,N_18157);
and U18304 (N_18304,N_18098,N_18029);
xor U18305 (N_18305,N_18119,N_18160);
nor U18306 (N_18306,N_18040,N_18076);
nand U18307 (N_18307,N_18157,N_18071);
nor U18308 (N_18308,N_18129,N_18150);
or U18309 (N_18309,N_18042,N_18051);
and U18310 (N_18310,N_18119,N_18028);
nand U18311 (N_18311,N_18142,N_18103);
and U18312 (N_18312,N_18162,N_18070);
nand U18313 (N_18313,N_18121,N_18043);
nand U18314 (N_18314,N_18048,N_18120);
nand U18315 (N_18315,N_18002,N_18198);
or U18316 (N_18316,N_18171,N_18068);
nand U18317 (N_18317,N_18063,N_18107);
nor U18318 (N_18318,N_18151,N_18023);
or U18319 (N_18319,N_18026,N_18096);
xor U18320 (N_18320,N_18051,N_18011);
nor U18321 (N_18321,N_18078,N_18172);
and U18322 (N_18322,N_18186,N_18120);
nand U18323 (N_18323,N_18183,N_18079);
nand U18324 (N_18324,N_18047,N_18036);
and U18325 (N_18325,N_18046,N_18070);
nor U18326 (N_18326,N_18073,N_18090);
xor U18327 (N_18327,N_18122,N_18054);
nand U18328 (N_18328,N_18024,N_18007);
nand U18329 (N_18329,N_18079,N_18146);
or U18330 (N_18330,N_18162,N_18016);
or U18331 (N_18331,N_18116,N_18071);
or U18332 (N_18332,N_18174,N_18095);
nand U18333 (N_18333,N_18001,N_18162);
nor U18334 (N_18334,N_18194,N_18175);
xor U18335 (N_18335,N_18042,N_18025);
xor U18336 (N_18336,N_18100,N_18108);
and U18337 (N_18337,N_18064,N_18083);
and U18338 (N_18338,N_18147,N_18073);
xor U18339 (N_18339,N_18115,N_18075);
xnor U18340 (N_18340,N_18140,N_18026);
or U18341 (N_18341,N_18102,N_18070);
or U18342 (N_18342,N_18111,N_18034);
nand U18343 (N_18343,N_18140,N_18185);
or U18344 (N_18344,N_18041,N_18007);
and U18345 (N_18345,N_18016,N_18155);
xor U18346 (N_18346,N_18177,N_18113);
xnor U18347 (N_18347,N_18051,N_18029);
nor U18348 (N_18348,N_18124,N_18079);
nand U18349 (N_18349,N_18165,N_18087);
xnor U18350 (N_18350,N_18073,N_18171);
nand U18351 (N_18351,N_18045,N_18102);
nand U18352 (N_18352,N_18021,N_18068);
nor U18353 (N_18353,N_18125,N_18049);
xor U18354 (N_18354,N_18135,N_18098);
nand U18355 (N_18355,N_18121,N_18133);
or U18356 (N_18356,N_18199,N_18126);
xor U18357 (N_18357,N_18185,N_18131);
nand U18358 (N_18358,N_18055,N_18097);
or U18359 (N_18359,N_18176,N_18014);
or U18360 (N_18360,N_18199,N_18130);
xnor U18361 (N_18361,N_18127,N_18010);
xnor U18362 (N_18362,N_18149,N_18130);
xor U18363 (N_18363,N_18133,N_18052);
and U18364 (N_18364,N_18073,N_18113);
and U18365 (N_18365,N_18012,N_18111);
or U18366 (N_18366,N_18188,N_18123);
xnor U18367 (N_18367,N_18174,N_18140);
and U18368 (N_18368,N_18049,N_18122);
or U18369 (N_18369,N_18019,N_18095);
or U18370 (N_18370,N_18077,N_18112);
xor U18371 (N_18371,N_18075,N_18025);
nor U18372 (N_18372,N_18157,N_18011);
xnor U18373 (N_18373,N_18090,N_18024);
nand U18374 (N_18374,N_18080,N_18164);
nand U18375 (N_18375,N_18126,N_18015);
and U18376 (N_18376,N_18083,N_18031);
xnor U18377 (N_18377,N_18030,N_18141);
or U18378 (N_18378,N_18078,N_18179);
nor U18379 (N_18379,N_18029,N_18133);
or U18380 (N_18380,N_18150,N_18044);
and U18381 (N_18381,N_18060,N_18141);
or U18382 (N_18382,N_18097,N_18032);
nor U18383 (N_18383,N_18005,N_18067);
nand U18384 (N_18384,N_18064,N_18173);
xnor U18385 (N_18385,N_18094,N_18059);
xnor U18386 (N_18386,N_18105,N_18022);
xor U18387 (N_18387,N_18119,N_18166);
and U18388 (N_18388,N_18054,N_18010);
nand U18389 (N_18389,N_18065,N_18166);
nor U18390 (N_18390,N_18169,N_18142);
nand U18391 (N_18391,N_18076,N_18136);
and U18392 (N_18392,N_18138,N_18101);
xor U18393 (N_18393,N_18068,N_18017);
xnor U18394 (N_18394,N_18036,N_18030);
and U18395 (N_18395,N_18093,N_18063);
xor U18396 (N_18396,N_18043,N_18051);
or U18397 (N_18397,N_18129,N_18178);
nor U18398 (N_18398,N_18110,N_18041);
nand U18399 (N_18399,N_18055,N_18153);
nand U18400 (N_18400,N_18272,N_18372);
nor U18401 (N_18401,N_18223,N_18390);
nor U18402 (N_18402,N_18391,N_18363);
nor U18403 (N_18403,N_18276,N_18203);
or U18404 (N_18404,N_18233,N_18224);
or U18405 (N_18405,N_18333,N_18282);
nand U18406 (N_18406,N_18273,N_18231);
and U18407 (N_18407,N_18318,N_18321);
nand U18408 (N_18408,N_18266,N_18214);
or U18409 (N_18409,N_18348,N_18341);
xor U18410 (N_18410,N_18210,N_18376);
nand U18411 (N_18411,N_18327,N_18325);
nor U18412 (N_18412,N_18384,N_18297);
nor U18413 (N_18413,N_18225,N_18388);
nor U18414 (N_18414,N_18259,N_18213);
or U18415 (N_18415,N_18251,N_18370);
xor U18416 (N_18416,N_18356,N_18238);
and U18417 (N_18417,N_18398,N_18389);
nor U18418 (N_18418,N_18248,N_18209);
nor U18419 (N_18419,N_18366,N_18395);
nor U18420 (N_18420,N_18293,N_18367);
nand U18421 (N_18421,N_18201,N_18287);
and U18422 (N_18422,N_18328,N_18230);
or U18423 (N_18423,N_18355,N_18295);
xor U18424 (N_18424,N_18305,N_18334);
nor U18425 (N_18425,N_18234,N_18313);
or U18426 (N_18426,N_18221,N_18397);
nand U18427 (N_18427,N_18378,N_18267);
or U18428 (N_18428,N_18284,N_18368);
nand U18429 (N_18429,N_18340,N_18314);
or U18430 (N_18430,N_18311,N_18336);
or U18431 (N_18431,N_18301,N_18208);
and U18432 (N_18432,N_18360,N_18365);
nand U18433 (N_18433,N_18300,N_18315);
or U18434 (N_18434,N_18204,N_18324);
nor U18435 (N_18435,N_18382,N_18394);
xor U18436 (N_18436,N_18241,N_18337);
xnor U18437 (N_18437,N_18250,N_18218);
or U18438 (N_18438,N_18329,N_18257);
nor U18439 (N_18439,N_18226,N_18335);
or U18440 (N_18440,N_18255,N_18383);
nor U18441 (N_18441,N_18339,N_18264);
xnor U18442 (N_18442,N_18288,N_18346);
and U18443 (N_18443,N_18386,N_18338);
and U18444 (N_18444,N_18359,N_18269);
nor U18445 (N_18445,N_18285,N_18309);
or U18446 (N_18446,N_18281,N_18399);
nand U18447 (N_18447,N_18396,N_18275);
or U18448 (N_18448,N_18242,N_18229);
nor U18449 (N_18449,N_18278,N_18350);
xnor U18450 (N_18450,N_18371,N_18317);
nor U18451 (N_18451,N_18361,N_18271);
nand U18452 (N_18452,N_18215,N_18243);
xor U18453 (N_18453,N_18216,N_18246);
nor U18454 (N_18454,N_18320,N_18244);
or U18455 (N_18455,N_18319,N_18274);
or U18456 (N_18456,N_18358,N_18298);
nor U18457 (N_18457,N_18268,N_18393);
nand U18458 (N_18458,N_18377,N_18380);
nand U18459 (N_18459,N_18239,N_18387);
or U18460 (N_18460,N_18322,N_18258);
nor U18461 (N_18461,N_18374,N_18369);
nand U18462 (N_18462,N_18392,N_18375);
nor U18463 (N_18463,N_18228,N_18294);
and U18464 (N_18464,N_18263,N_18283);
xor U18465 (N_18465,N_18235,N_18362);
nand U18466 (N_18466,N_18323,N_18306);
and U18467 (N_18467,N_18240,N_18200);
or U18468 (N_18468,N_18227,N_18307);
xor U18469 (N_18469,N_18217,N_18220);
nand U18470 (N_18470,N_18260,N_18351);
xor U18471 (N_18471,N_18253,N_18211);
or U18472 (N_18472,N_18353,N_18357);
or U18473 (N_18473,N_18349,N_18286);
nor U18474 (N_18474,N_18379,N_18202);
nand U18475 (N_18475,N_18206,N_18247);
nor U18476 (N_18476,N_18381,N_18332);
nor U18477 (N_18477,N_18302,N_18245);
or U18478 (N_18478,N_18343,N_18347);
or U18479 (N_18479,N_18385,N_18265);
and U18480 (N_18480,N_18232,N_18261);
or U18481 (N_18481,N_18316,N_18212);
xor U18482 (N_18482,N_18262,N_18331);
xnor U18483 (N_18483,N_18277,N_18303);
or U18484 (N_18484,N_18312,N_18289);
nand U18485 (N_18485,N_18344,N_18252);
nand U18486 (N_18486,N_18219,N_18304);
nand U18487 (N_18487,N_18291,N_18364);
or U18488 (N_18488,N_18292,N_18270);
or U18489 (N_18489,N_18254,N_18205);
nand U18490 (N_18490,N_18310,N_18256);
and U18491 (N_18491,N_18296,N_18330);
nand U18492 (N_18492,N_18308,N_18342);
xor U18493 (N_18493,N_18280,N_18352);
nand U18494 (N_18494,N_18222,N_18373);
xnor U18495 (N_18495,N_18354,N_18299);
and U18496 (N_18496,N_18236,N_18345);
and U18497 (N_18497,N_18237,N_18290);
nand U18498 (N_18498,N_18249,N_18207);
and U18499 (N_18499,N_18326,N_18279);
nor U18500 (N_18500,N_18375,N_18315);
and U18501 (N_18501,N_18269,N_18289);
nor U18502 (N_18502,N_18228,N_18252);
nand U18503 (N_18503,N_18268,N_18219);
and U18504 (N_18504,N_18306,N_18313);
or U18505 (N_18505,N_18229,N_18396);
nand U18506 (N_18506,N_18390,N_18249);
and U18507 (N_18507,N_18238,N_18361);
xnor U18508 (N_18508,N_18266,N_18211);
and U18509 (N_18509,N_18333,N_18313);
or U18510 (N_18510,N_18344,N_18294);
or U18511 (N_18511,N_18330,N_18390);
and U18512 (N_18512,N_18337,N_18397);
nor U18513 (N_18513,N_18327,N_18349);
xor U18514 (N_18514,N_18320,N_18300);
nand U18515 (N_18515,N_18277,N_18245);
or U18516 (N_18516,N_18389,N_18292);
xor U18517 (N_18517,N_18342,N_18385);
nand U18518 (N_18518,N_18398,N_18234);
or U18519 (N_18519,N_18348,N_18275);
nor U18520 (N_18520,N_18378,N_18294);
nor U18521 (N_18521,N_18205,N_18328);
xor U18522 (N_18522,N_18202,N_18304);
nor U18523 (N_18523,N_18298,N_18364);
or U18524 (N_18524,N_18250,N_18262);
and U18525 (N_18525,N_18343,N_18271);
nor U18526 (N_18526,N_18276,N_18208);
xnor U18527 (N_18527,N_18242,N_18318);
and U18528 (N_18528,N_18217,N_18280);
nor U18529 (N_18529,N_18233,N_18346);
nor U18530 (N_18530,N_18217,N_18317);
xnor U18531 (N_18531,N_18252,N_18237);
xnor U18532 (N_18532,N_18201,N_18241);
and U18533 (N_18533,N_18301,N_18346);
xnor U18534 (N_18534,N_18316,N_18211);
nor U18535 (N_18535,N_18204,N_18318);
nand U18536 (N_18536,N_18297,N_18212);
or U18537 (N_18537,N_18256,N_18349);
xor U18538 (N_18538,N_18219,N_18388);
nor U18539 (N_18539,N_18280,N_18242);
nor U18540 (N_18540,N_18235,N_18366);
or U18541 (N_18541,N_18391,N_18285);
nand U18542 (N_18542,N_18307,N_18363);
xor U18543 (N_18543,N_18237,N_18371);
nor U18544 (N_18544,N_18222,N_18250);
or U18545 (N_18545,N_18371,N_18324);
or U18546 (N_18546,N_18209,N_18238);
xor U18547 (N_18547,N_18274,N_18330);
nand U18548 (N_18548,N_18380,N_18244);
nor U18549 (N_18549,N_18359,N_18286);
or U18550 (N_18550,N_18262,N_18364);
and U18551 (N_18551,N_18217,N_18225);
or U18552 (N_18552,N_18278,N_18225);
or U18553 (N_18553,N_18306,N_18387);
nor U18554 (N_18554,N_18267,N_18287);
xnor U18555 (N_18555,N_18214,N_18293);
and U18556 (N_18556,N_18289,N_18287);
nor U18557 (N_18557,N_18312,N_18262);
or U18558 (N_18558,N_18318,N_18251);
nor U18559 (N_18559,N_18317,N_18343);
nor U18560 (N_18560,N_18235,N_18303);
xnor U18561 (N_18561,N_18349,N_18281);
xnor U18562 (N_18562,N_18329,N_18391);
or U18563 (N_18563,N_18348,N_18393);
and U18564 (N_18564,N_18205,N_18308);
xnor U18565 (N_18565,N_18348,N_18304);
nor U18566 (N_18566,N_18334,N_18349);
or U18567 (N_18567,N_18360,N_18212);
and U18568 (N_18568,N_18249,N_18369);
xor U18569 (N_18569,N_18226,N_18395);
and U18570 (N_18570,N_18337,N_18389);
nor U18571 (N_18571,N_18362,N_18366);
or U18572 (N_18572,N_18234,N_18351);
nand U18573 (N_18573,N_18228,N_18236);
and U18574 (N_18574,N_18306,N_18354);
xor U18575 (N_18575,N_18311,N_18293);
xor U18576 (N_18576,N_18334,N_18336);
xor U18577 (N_18577,N_18303,N_18314);
xnor U18578 (N_18578,N_18250,N_18318);
nand U18579 (N_18579,N_18289,N_18300);
and U18580 (N_18580,N_18280,N_18213);
and U18581 (N_18581,N_18314,N_18296);
or U18582 (N_18582,N_18273,N_18369);
nand U18583 (N_18583,N_18376,N_18299);
and U18584 (N_18584,N_18396,N_18291);
xnor U18585 (N_18585,N_18363,N_18296);
xor U18586 (N_18586,N_18212,N_18266);
or U18587 (N_18587,N_18252,N_18334);
nand U18588 (N_18588,N_18256,N_18278);
or U18589 (N_18589,N_18245,N_18391);
or U18590 (N_18590,N_18238,N_18350);
xnor U18591 (N_18591,N_18343,N_18335);
or U18592 (N_18592,N_18383,N_18397);
or U18593 (N_18593,N_18295,N_18300);
xor U18594 (N_18594,N_18285,N_18306);
nor U18595 (N_18595,N_18398,N_18202);
xor U18596 (N_18596,N_18394,N_18232);
nand U18597 (N_18597,N_18300,N_18379);
or U18598 (N_18598,N_18225,N_18254);
nor U18599 (N_18599,N_18341,N_18316);
or U18600 (N_18600,N_18405,N_18574);
and U18601 (N_18601,N_18453,N_18422);
or U18602 (N_18602,N_18463,N_18417);
nand U18603 (N_18603,N_18497,N_18506);
nor U18604 (N_18604,N_18476,N_18424);
xor U18605 (N_18605,N_18530,N_18498);
xnor U18606 (N_18606,N_18598,N_18467);
nand U18607 (N_18607,N_18559,N_18544);
or U18608 (N_18608,N_18520,N_18557);
and U18609 (N_18609,N_18505,N_18564);
or U18610 (N_18610,N_18481,N_18510);
nor U18611 (N_18611,N_18529,N_18408);
nand U18612 (N_18612,N_18435,N_18438);
or U18613 (N_18613,N_18522,N_18567);
xnor U18614 (N_18614,N_18434,N_18579);
and U18615 (N_18615,N_18508,N_18430);
xor U18616 (N_18616,N_18409,N_18445);
or U18617 (N_18617,N_18493,N_18555);
or U18618 (N_18618,N_18480,N_18406);
nor U18619 (N_18619,N_18575,N_18479);
and U18620 (N_18620,N_18410,N_18490);
and U18621 (N_18621,N_18553,N_18440);
and U18622 (N_18622,N_18441,N_18412);
nand U18623 (N_18623,N_18419,N_18538);
xor U18624 (N_18624,N_18540,N_18526);
and U18625 (N_18625,N_18446,N_18584);
nand U18626 (N_18626,N_18489,N_18403);
xnor U18627 (N_18627,N_18569,N_18411);
nor U18628 (N_18628,N_18556,N_18460);
xor U18629 (N_18629,N_18546,N_18459);
nand U18630 (N_18630,N_18429,N_18433);
nor U18631 (N_18631,N_18562,N_18491);
xnor U18632 (N_18632,N_18452,N_18531);
nor U18633 (N_18633,N_18561,N_18503);
or U18634 (N_18634,N_18487,N_18488);
nand U18635 (N_18635,N_18478,N_18416);
nor U18636 (N_18636,N_18499,N_18472);
nand U18637 (N_18637,N_18418,N_18532);
xor U18638 (N_18638,N_18473,N_18402);
or U18639 (N_18639,N_18448,N_18485);
nand U18640 (N_18640,N_18523,N_18527);
nor U18641 (N_18641,N_18577,N_18566);
nand U18642 (N_18642,N_18494,N_18492);
nand U18643 (N_18643,N_18507,N_18449);
xnor U18644 (N_18644,N_18587,N_18437);
xnor U18645 (N_18645,N_18436,N_18570);
and U18646 (N_18646,N_18426,N_18590);
nand U18647 (N_18647,N_18413,N_18458);
xor U18648 (N_18648,N_18420,N_18533);
and U18649 (N_18649,N_18568,N_18461);
nor U18650 (N_18650,N_18558,N_18582);
and U18651 (N_18651,N_18486,N_18576);
nor U18652 (N_18652,N_18571,N_18443);
nand U18653 (N_18653,N_18444,N_18469);
or U18654 (N_18654,N_18552,N_18578);
nand U18655 (N_18655,N_18509,N_18442);
nor U18656 (N_18656,N_18462,N_18547);
xor U18657 (N_18657,N_18513,N_18548);
or U18658 (N_18658,N_18536,N_18549);
nand U18659 (N_18659,N_18421,N_18495);
nor U18660 (N_18660,N_18427,N_18496);
xor U18661 (N_18661,N_18514,N_18439);
nor U18662 (N_18662,N_18432,N_18482);
xnor U18663 (N_18663,N_18596,N_18560);
or U18664 (N_18664,N_18518,N_18534);
nor U18665 (N_18665,N_18551,N_18572);
nand U18666 (N_18666,N_18414,N_18470);
and U18667 (N_18667,N_18539,N_18565);
or U18668 (N_18668,N_18484,N_18519);
and U18669 (N_18669,N_18428,N_18521);
xor U18670 (N_18670,N_18474,N_18591);
nand U18671 (N_18671,N_18589,N_18588);
nor U18672 (N_18672,N_18599,N_18466);
nand U18673 (N_18673,N_18457,N_18554);
and U18674 (N_18674,N_18525,N_18512);
nor U18675 (N_18675,N_18580,N_18454);
and U18676 (N_18676,N_18550,N_18573);
xnor U18677 (N_18677,N_18545,N_18447);
xor U18678 (N_18678,N_18415,N_18592);
nor U18679 (N_18679,N_18468,N_18404);
or U18680 (N_18680,N_18593,N_18431);
or U18681 (N_18681,N_18537,N_18535);
nand U18682 (N_18682,N_18594,N_18501);
nor U18683 (N_18683,N_18504,N_18502);
nor U18684 (N_18684,N_18516,N_18423);
nand U18685 (N_18685,N_18563,N_18528);
or U18686 (N_18686,N_18585,N_18483);
or U18687 (N_18687,N_18400,N_18542);
or U18688 (N_18688,N_18451,N_18541);
and U18689 (N_18689,N_18586,N_18425);
or U18690 (N_18690,N_18511,N_18471);
and U18691 (N_18691,N_18455,N_18407);
or U18692 (N_18692,N_18456,N_18583);
nand U18693 (N_18693,N_18524,N_18450);
and U18694 (N_18694,N_18597,N_18595);
nand U18695 (N_18695,N_18500,N_18464);
nor U18696 (N_18696,N_18515,N_18477);
and U18697 (N_18697,N_18465,N_18401);
nand U18698 (N_18698,N_18581,N_18475);
nor U18699 (N_18699,N_18517,N_18543);
nand U18700 (N_18700,N_18513,N_18599);
xor U18701 (N_18701,N_18404,N_18412);
or U18702 (N_18702,N_18562,N_18417);
xnor U18703 (N_18703,N_18455,N_18446);
nor U18704 (N_18704,N_18401,N_18472);
xor U18705 (N_18705,N_18557,N_18494);
or U18706 (N_18706,N_18543,N_18586);
nand U18707 (N_18707,N_18506,N_18487);
and U18708 (N_18708,N_18470,N_18437);
and U18709 (N_18709,N_18579,N_18457);
and U18710 (N_18710,N_18530,N_18543);
nor U18711 (N_18711,N_18403,N_18590);
nor U18712 (N_18712,N_18502,N_18461);
nor U18713 (N_18713,N_18406,N_18437);
and U18714 (N_18714,N_18486,N_18511);
nor U18715 (N_18715,N_18596,N_18404);
or U18716 (N_18716,N_18429,N_18523);
xnor U18717 (N_18717,N_18462,N_18587);
and U18718 (N_18718,N_18514,N_18547);
nand U18719 (N_18719,N_18524,N_18554);
or U18720 (N_18720,N_18465,N_18504);
nor U18721 (N_18721,N_18478,N_18451);
and U18722 (N_18722,N_18592,N_18491);
or U18723 (N_18723,N_18547,N_18401);
nor U18724 (N_18724,N_18457,N_18469);
and U18725 (N_18725,N_18444,N_18530);
and U18726 (N_18726,N_18431,N_18568);
and U18727 (N_18727,N_18445,N_18599);
nand U18728 (N_18728,N_18446,N_18539);
nor U18729 (N_18729,N_18595,N_18547);
or U18730 (N_18730,N_18444,N_18517);
nand U18731 (N_18731,N_18598,N_18509);
and U18732 (N_18732,N_18459,N_18498);
nor U18733 (N_18733,N_18453,N_18483);
or U18734 (N_18734,N_18447,N_18554);
nand U18735 (N_18735,N_18412,N_18540);
xnor U18736 (N_18736,N_18417,N_18428);
nor U18737 (N_18737,N_18427,N_18598);
nor U18738 (N_18738,N_18523,N_18598);
nand U18739 (N_18739,N_18543,N_18553);
nor U18740 (N_18740,N_18452,N_18446);
xor U18741 (N_18741,N_18415,N_18521);
nor U18742 (N_18742,N_18578,N_18422);
nor U18743 (N_18743,N_18557,N_18411);
nor U18744 (N_18744,N_18575,N_18572);
or U18745 (N_18745,N_18586,N_18443);
nand U18746 (N_18746,N_18477,N_18415);
nand U18747 (N_18747,N_18429,N_18478);
or U18748 (N_18748,N_18420,N_18522);
or U18749 (N_18749,N_18542,N_18509);
nor U18750 (N_18750,N_18572,N_18545);
or U18751 (N_18751,N_18466,N_18579);
and U18752 (N_18752,N_18441,N_18403);
nand U18753 (N_18753,N_18409,N_18511);
or U18754 (N_18754,N_18537,N_18418);
nor U18755 (N_18755,N_18442,N_18421);
or U18756 (N_18756,N_18402,N_18564);
nand U18757 (N_18757,N_18421,N_18552);
and U18758 (N_18758,N_18564,N_18504);
xnor U18759 (N_18759,N_18524,N_18432);
nor U18760 (N_18760,N_18400,N_18512);
or U18761 (N_18761,N_18591,N_18414);
xnor U18762 (N_18762,N_18427,N_18452);
xor U18763 (N_18763,N_18587,N_18478);
and U18764 (N_18764,N_18469,N_18441);
nor U18765 (N_18765,N_18418,N_18447);
nor U18766 (N_18766,N_18503,N_18566);
or U18767 (N_18767,N_18410,N_18452);
nand U18768 (N_18768,N_18564,N_18560);
nand U18769 (N_18769,N_18585,N_18567);
nand U18770 (N_18770,N_18496,N_18411);
nand U18771 (N_18771,N_18494,N_18536);
or U18772 (N_18772,N_18492,N_18466);
nand U18773 (N_18773,N_18476,N_18540);
nor U18774 (N_18774,N_18466,N_18441);
nor U18775 (N_18775,N_18404,N_18415);
nand U18776 (N_18776,N_18460,N_18402);
or U18777 (N_18777,N_18588,N_18474);
xnor U18778 (N_18778,N_18519,N_18564);
nor U18779 (N_18779,N_18560,N_18513);
xnor U18780 (N_18780,N_18426,N_18506);
and U18781 (N_18781,N_18475,N_18524);
or U18782 (N_18782,N_18502,N_18457);
nand U18783 (N_18783,N_18514,N_18420);
and U18784 (N_18784,N_18588,N_18515);
or U18785 (N_18785,N_18474,N_18461);
and U18786 (N_18786,N_18452,N_18467);
or U18787 (N_18787,N_18573,N_18487);
nor U18788 (N_18788,N_18472,N_18404);
and U18789 (N_18789,N_18490,N_18531);
nand U18790 (N_18790,N_18472,N_18508);
nand U18791 (N_18791,N_18536,N_18533);
xnor U18792 (N_18792,N_18553,N_18510);
nand U18793 (N_18793,N_18469,N_18563);
nor U18794 (N_18794,N_18545,N_18594);
nand U18795 (N_18795,N_18448,N_18576);
and U18796 (N_18796,N_18401,N_18548);
or U18797 (N_18797,N_18458,N_18462);
xor U18798 (N_18798,N_18483,N_18578);
xor U18799 (N_18799,N_18554,N_18588);
nand U18800 (N_18800,N_18616,N_18708);
nand U18801 (N_18801,N_18697,N_18700);
xnor U18802 (N_18802,N_18711,N_18732);
nor U18803 (N_18803,N_18726,N_18679);
nor U18804 (N_18804,N_18799,N_18767);
nor U18805 (N_18805,N_18724,N_18770);
and U18806 (N_18806,N_18672,N_18626);
nand U18807 (N_18807,N_18783,N_18788);
or U18808 (N_18808,N_18641,N_18787);
nand U18809 (N_18809,N_18763,N_18753);
nand U18810 (N_18810,N_18747,N_18655);
nand U18811 (N_18811,N_18646,N_18678);
nor U18812 (N_18812,N_18682,N_18683);
and U18813 (N_18813,N_18650,N_18656);
or U18814 (N_18814,N_18612,N_18781);
xnor U18815 (N_18815,N_18756,N_18660);
or U18816 (N_18816,N_18659,N_18628);
and U18817 (N_18817,N_18714,N_18796);
xor U18818 (N_18818,N_18617,N_18765);
and U18819 (N_18819,N_18699,N_18666);
nand U18820 (N_18820,N_18772,N_18762);
or U18821 (N_18821,N_18644,N_18603);
or U18822 (N_18822,N_18631,N_18627);
xor U18823 (N_18823,N_18635,N_18786);
nor U18824 (N_18824,N_18642,N_18661);
nor U18825 (N_18825,N_18748,N_18733);
nor U18826 (N_18826,N_18709,N_18601);
nand U18827 (N_18827,N_18632,N_18743);
xnor U18828 (N_18828,N_18725,N_18730);
nand U18829 (N_18829,N_18618,N_18658);
nor U18830 (N_18830,N_18744,N_18671);
or U18831 (N_18831,N_18773,N_18737);
or U18832 (N_18832,N_18701,N_18761);
or U18833 (N_18833,N_18611,N_18653);
nor U18834 (N_18834,N_18705,N_18774);
or U18835 (N_18835,N_18685,N_18689);
nor U18836 (N_18836,N_18621,N_18794);
nand U18837 (N_18837,N_18639,N_18624);
xnor U18838 (N_18838,N_18633,N_18649);
and U18839 (N_18839,N_18604,N_18674);
and U18840 (N_18840,N_18637,N_18681);
nand U18841 (N_18841,N_18759,N_18790);
or U18842 (N_18842,N_18749,N_18793);
nand U18843 (N_18843,N_18746,N_18605);
or U18844 (N_18844,N_18771,N_18703);
or U18845 (N_18845,N_18782,N_18694);
and U18846 (N_18846,N_18692,N_18610);
nor U18847 (N_18847,N_18664,N_18643);
xnor U18848 (N_18848,N_18630,N_18677);
xnor U18849 (N_18849,N_18652,N_18760);
nand U18850 (N_18850,N_18758,N_18663);
or U18851 (N_18851,N_18795,N_18702);
or U18852 (N_18852,N_18775,N_18625);
and U18853 (N_18853,N_18607,N_18693);
or U18854 (N_18854,N_18729,N_18784);
xor U18855 (N_18855,N_18719,N_18704);
and U18856 (N_18856,N_18602,N_18738);
nand U18857 (N_18857,N_18609,N_18686);
or U18858 (N_18858,N_18640,N_18721);
xor U18859 (N_18859,N_18766,N_18741);
nor U18860 (N_18860,N_18722,N_18675);
nand U18861 (N_18861,N_18614,N_18657);
nor U18862 (N_18862,N_18769,N_18669);
and U18863 (N_18863,N_18739,N_18716);
xnor U18864 (N_18864,N_18620,N_18713);
nor U18865 (N_18865,N_18622,N_18751);
and U18866 (N_18866,N_18791,N_18740);
nor U18867 (N_18867,N_18670,N_18667);
or U18868 (N_18868,N_18684,N_18715);
nor U18869 (N_18869,N_18613,N_18710);
or U18870 (N_18870,N_18690,N_18785);
nor U18871 (N_18871,N_18688,N_18735);
nor U18872 (N_18872,N_18745,N_18731);
or U18873 (N_18873,N_18734,N_18757);
or U18874 (N_18874,N_18755,N_18768);
or U18875 (N_18875,N_18673,N_18615);
and U18876 (N_18876,N_18623,N_18636);
nand U18877 (N_18877,N_18654,N_18712);
and U18878 (N_18878,N_18750,N_18723);
or U18879 (N_18879,N_18728,N_18647);
or U18880 (N_18880,N_18600,N_18776);
nor U18881 (N_18881,N_18778,N_18645);
nand U18882 (N_18882,N_18720,N_18752);
xnor U18883 (N_18883,N_18662,N_18789);
xnor U18884 (N_18884,N_18717,N_18718);
nand U18885 (N_18885,N_18676,N_18706);
nand U18886 (N_18886,N_18754,N_18619);
or U18887 (N_18887,N_18691,N_18696);
nand U18888 (N_18888,N_18742,N_18797);
xor U18889 (N_18889,N_18777,N_18680);
nor U18890 (N_18890,N_18780,N_18665);
and U18891 (N_18891,N_18695,N_18608);
or U18892 (N_18892,N_18727,N_18698);
nor U18893 (N_18893,N_18638,N_18798);
or U18894 (N_18894,N_18651,N_18648);
and U18895 (N_18895,N_18779,N_18687);
or U18896 (N_18896,N_18634,N_18668);
or U18897 (N_18897,N_18792,N_18606);
and U18898 (N_18898,N_18629,N_18707);
or U18899 (N_18899,N_18736,N_18764);
nor U18900 (N_18900,N_18714,N_18611);
nand U18901 (N_18901,N_18756,N_18681);
xor U18902 (N_18902,N_18656,N_18666);
and U18903 (N_18903,N_18792,N_18603);
nor U18904 (N_18904,N_18612,N_18613);
or U18905 (N_18905,N_18646,N_18633);
or U18906 (N_18906,N_18651,N_18786);
xor U18907 (N_18907,N_18622,N_18691);
nor U18908 (N_18908,N_18726,N_18687);
nand U18909 (N_18909,N_18625,N_18635);
or U18910 (N_18910,N_18704,N_18709);
and U18911 (N_18911,N_18792,N_18679);
and U18912 (N_18912,N_18685,N_18714);
or U18913 (N_18913,N_18654,N_18758);
nor U18914 (N_18914,N_18668,N_18726);
nand U18915 (N_18915,N_18621,N_18776);
xor U18916 (N_18916,N_18774,N_18736);
or U18917 (N_18917,N_18664,N_18699);
or U18918 (N_18918,N_18785,N_18642);
xor U18919 (N_18919,N_18624,N_18603);
nand U18920 (N_18920,N_18708,N_18746);
nor U18921 (N_18921,N_18604,N_18693);
xnor U18922 (N_18922,N_18651,N_18603);
nand U18923 (N_18923,N_18708,N_18771);
or U18924 (N_18924,N_18606,N_18604);
nor U18925 (N_18925,N_18644,N_18647);
xor U18926 (N_18926,N_18762,N_18780);
and U18927 (N_18927,N_18757,N_18750);
nand U18928 (N_18928,N_18704,N_18609);
xnor U18929 (N_18929,N_18752,N_18738);
or U18930 (N_18930,N_18751,N_18799);
nand U18931 (N_18931,N_18734,N_18788);
or U18932 (N_18932,N_18616,N_18601);
and U18933 (N_18933,N_18641,N_18773);
xnor U18934 (N_18934,N_18696,N_18714);
xnor U18935 (N_18935,N_18629,N_18719);
and U18936 (N_18936,N_18636,N_18754);
or U18937 (N_18937,N_18636,N_18779);
and U18938 (N_18938,N_18686,N_18665);
nand U18939 (N_18939,N_18712,N_18777);
nor U18940 (N_18940,N_18788,N_18667);
nor U18941 (N_18941,N_18627,N_18713);
xor U18942 (N_18942,N_18727,N_18670);
or U18943 (N_18943,N_18647,N_18785);
and U18944 (N_18944,N_18748,N_18786);
xor U18945 (N_18945,N_18778,N_18794);
xnor U18946 (N_18946,N_18773,N_18695);
xnor U18947 (N_18947,N_18755,N_18675);
nand U18948 (N_18948,N_18669,N_18645);
xnor U18949 (N_18949,N_18688,N_18601);
xnor U18950 (N_18950,N_18714,N_18703);
nand U18951 (N_18951,N_18759,N_18721);
nand U18952 (N_18952,N_18686,N_18751);
nand U18953 (N_18953,N_18623,N_18738);
nor U18954 (N_18954,N_18621,N_18639);
and U18955 (N_18955,N_18785,N_18605);
nand U18956 (N_18956,N_18667,N_18741);
nand U18957 (N_18957,N_18745,N_18631);
nand U18958 (N_18958,N_18746,N_18637);
or U18959 (N_18959,N_18644,N_18783);
nor U18960 (N_18960,N_18646,N_18628);
nand U18961 (N_18961,N_18724,N_18658);
nor U18962 (N_18962,N_18759,N_18736);
or U18963 (N_18963,N_18661,N_18600);
nor U18964 (N_18964,N_18738,N_18605);
nor U18965 (N_18965,N_18650,N_18661);
and U18966 (N_18966,N_18669,N_18608);
and U18967 (N_18967,N_18710,N_18781);
and U18968 (N_18968,N_18758,N_18640);
and U18969 (N_18969,N_18692,N_18670);
nand U18970 (N_18970,N_18644,N_18774);
and U18971 (N_18971,N_18638,N_18776);
nand U18972 (N_18972,N_18620,N_18778);
nand U18973 (N_18973,N_18755,N_18719);
nor U18974 (N_18974,N_18747,N_18765);
xor U18975 (N_18975,N_18728,N_18763);
nor U18976 (N_18976,N_18754,N_18739);
nand U18977 (N_18977,N_18769,N_18742);
nor U18978 (N_18978,N_18601,N_18762);
nand U18979 (N_18979,N_18795,N_18739);
xor U18980 (N_18980,N_18745,N_18787);
nand U18981 (N_18981,N_18681,N_18761);
or U18982 (N_18982,N_18769,N_18661);
xnor U18983 (N_18983,N_18754,N_18753);
xnor U18984 (N_18984,N_18711,N_18738);
nor U18985 (N_18985,N_18660,N_18638);
or U18986 (N_18986,N_18728,N_18627);
xor U18987 (N_18987,N_18605,N_18731);
nor U18988 (N_18988,N_18639,N_18636);
nand U18989 (N_18989,N_18680,N_18644);
or U18990 (N_18990,N_18680,N_18735);
nor U18991 (N_18991,N_18716,N_18730);
xor U18992 (N_18992,N_18740,N_18647);
and U18993 (N_18993,N_18770,N_18783);
nor U18994 (N_18994,N_18639,N_18654);
or U18995 (N_18995,N_18659,N_18740);
nor U18996 (N_18996,N_18774,N_18749);
xnor U18997 (N_18997,N_18614,N_18725);
and U18998 (N_18998,N_18671,N_18765);
nand U18999 (N_18999,N_18667,N_18646);
or U19000 (N_19000,N_18811,N_18907);
or U19001 (N_19001,N_18965,N_18903);
nand U19002 (N_19002,N_18967,N_18867);
nor U19003 (N_19003,N_18917,N_18912);
nor U19004 (N_19004,N_18897,N_18821);
and U19005 (N_19005,N_18944,N_18801);
or U19006 (N_19006,N_18849,N_18941);
xor U19007 (N_19007,N_18991,N_18943);
nand U19008 (N_19008,N_18893,N_18972);
nand U19009 (N_19009,N_18839,N_18922);
or U19010 (N_19010,N_18854,N_18950);
or U19011 (N_19011,N_18892,N_18885);
or U19012 (N_19012,N_18833,N_18868);
xor U19013 (N_19013,N_18986,N_18840);
or U19014 (N_19014,N_18895,N_18876);
nor U19015 (N_19015,N_18843,N_18880);
nand U19016 (N_19016,N_18938,N_18992);
nor U19017 (N_19017,N_18915,N_18805);
xnor U19018 (N_19018,N_18988,N_18810);
xnor U19019 (N_19019,N_18926,N_18858);
xor U19020 (N_19020,N_18989,N_18931);
xor U19021 (N_19021,N_18924,N_18990);
or U19022 (N_19022,N_18934,N_18960);
nand U19023 (N_19023,N_18873,N_18818);
nand U19024 (N_19024,N_18957,N_18969);
and U19025 (N_19025,N_18827,N_18890);
nand U19026 (N_19026,N_18975,N_18879);
nand U19027 (N_19027,N_18898,N_18951);
or U19028 (N_19028,N_18901,N_18993);
or U19029 (N_19029,N_18942,N_18812);
nor U19030 (N_19030,N_18883,N_18930);
nand U19031 (N_19031,N_18819,N_18828);
and U19032 (N_19032,N_18998,N_18856);
nand U19033 (N_19033,N_18981,N_18923);
nor U19034 (N_19034,N_18886,N_18863);
xor U19035 (N_19035,N_18822,N_18888);
and U19036 (N_19036,N_18997,N_18846);
or U19037 (N_19037,N_18947,N_18838);
and U19038 (N_19038,N_18980,N_18881);
or U19039 (N_19039,N_18921,N_18877);
nor U19040 (N_19040,N_18932,N_18808);
nand U19041 (N_19041,N_18829,N_18826);
or U19042 (N_19042,N_18933,N_18896);
xor U19043 (N_19043,N_18911,N_18948);
nor U19044 (N_19044,N_18977,N_18936);
or U19045 (N_19045,N_18985,N_18968);
xnor U19046 (N_19046,N_18929,N_18804);
nor U19047 (N_19047,N_18800,N_18900);
xnor U19048 (N_19048,N_18952,N_18954);
and U19049 (N_19049,N_18994,N_18832);
and U19050 (N_19050,N_18853,N_18995);
xor U19051 (N_19051,N_18953,N_18955);
nor U19052 (N_19052,N_18872,N_18874);
nor U19053 (N_19053,N_18966,N_18920);
and U19054 (N_19054,N_18802,N_18831);
or U19055 (N_19055,N_18889,N_18987);
or U19056 (N_19056,N_18940,N_18816);
and U19057 (N_19057,N_18959,N_18852);
or U19058 (N_19058,N_18904,N_18891);
nor U19059 (N_19059,N_18857,N_18847);
xor U19060 (N_19060,N_18806,N_18803);
and U19061 (N_19061,N_18916,N_18961);
xnor U19062 (N_19062,N_18970,N_18860);
nor U19063 (N_19063,N_18958,N_18913);
nand U19064 (N_19064,N_18820,N_18884);
or U19065 (N_19065,N_18864,N_18830);
nand U19066 (N_19066,N_18871,N_18869);
xor U19067 (N_19067,N_18928,N_18841);
nand U19068 (N_19068,N_18855,N_18973);
nand U19069 (N_19069,N_18949,N_18927);
and U19070 (N_19070,N_18946,N_18848);
nand U19071 (N_19071,N_18996,N_18862);
nand U19072 (N_19072,N_18962,N_18807);
or U19073 (N_19073,N_18935,N_18964);
or U19074 (N_19074,N_18963,N_18937);
nor U19075 (N_19075,N_18925,N_18882);
nor U19076 (N_19076,N_18910,N_18851);
nand U19077 (N_19077,N_18999,N_18899);
or U19078 (N_19078,N_18984,N_18905);
nand U19079 (N_19079,N_18837,N_18866);
xnor U19080 (N_19080,N_18894,N_18814);
and U19081 (N_19081,N_18983,N_18979);
nor U19082 (N_19082,N_18971,N_18909);
xor U19083 (N_19083,N_18813,N_18974);
nor U19084 (N_19084,N_18825,N_18914);
nor U19085 (N_19085,N_18836,N_18842);
xor U19086 (N_19086,N_18956,N_18824);
xor U19087 (N_19087,N_18906,N_18870);
nand U19088 (N_19088,N_18919,N_18865);
and U19089 (N_19089,N_18878,N_18887);
or U19090 (N_19090,N_18861,N_18902);
nand U19091 (N_19091,N_18817,N_18945);
nand U19092 (N_19092,N_18834,N_18859);
xnor U19093 (N_19093,N_18845,N_18844);
and U19094 (N_19094,N_18918,N_18823);
or U19095 (N_19095,N_18835,N_18850);
and U19096 (N_19096,N_18809,N_18908);
nor U19097 (N_19097,N_18875,N_18976);
nand U19098 (N_19098,N_18978,N_18982);
or U19099 (N_19099,N_18939,N_18815);
nor U19100 (N_19100,N_18919,N_18821);
nor U19101 (N_19101,N_18981,N_18870);
xnor U19102 (N_19102,N_18925,N_18946);
or U19103 (N_19103,N_18930,N_18984);
and U19104 (N_19104,N_18875,N_18924);
xor U19105 (N_19105,N_18996,N_18942);
nand U19106 (N_19106,N_18823,N_18945);
nor U19107 (N_19107,N_18828,N_18802);
and U19108 (N_19108,N_18912,N_18992);
nor U19109 (N_19109,N_18921,N_18894);
xor U19110 (N_19110,N_18966,N_18940);
and U19111 (N_19111,N_18958,N_18808);
and U19112 (N_19112,N_18979,N_18995);
or U19113 (N_19113,N_18919,N_18976);
xor U19114 (N_19114,N_18841,N_18882);
and U19115 (N_19115,N_18809,N_18822);
and U19116 (N_19116,N_18910,N_18883);
xor U19117 (N_19117,N_18804,N_18828);
and U19118 (N_19118,N_18824,N_18919);
or U19119 (N_19119,N_18959,N_18937);
or U19120 (N_19120,N_18903,N_18988);
nor U19121 (N_19121,N_18813,N_18906);
and U19122 (N_19122,N_18837,N_18828);
and U19123 (N_19123,N_18935,N_18891);
and U19124 (N_19124,N_18870,N_18803);
or U19125 (N_19125,N_18909,N_18885);
or U19126 (N_19126,N_18845,N_18962);
or U19127 (N_19127,N_18952,N_18992);
nand U19128 (N_19128,N_18922,N_18817);
or U19129 (N_19129,N_18871,N_18865);
or U19130 (N_19130,N_18813,N_18951);
or U19131 (N_19131,N_18945,N_18991);
nand U19132 (N_19132,N_18846,N_18886);
nand U19133 (N_19133,N_18914,N_18871);
nor U19134 (N_19134,N_18825,N_18950);
and U19135 (N_19135,N_18910,N_18958);
nor U19136 (N_19136,N_18905,N_18869);
xnor U19137 (N_19137,N_18992,N_18893);
nor U19138 (N_19138,N_18940,N_18838);
nor U19139 (N_19139,N_18975,N_18827);
or U19140 (N_19140,N_18904,N_18981);
nor U19141 (N_19141,N_18805,N_18833);
xor U19142 (N_19142,N_18963,N_18813);
nand U19143 (N_19143,N_18855,N_18834);
xnor U19144 (N_19144,N_18887,N_18826);
and U19145 (N_19145,N_18992,N_18993);
and U19146 (N_19146,N_18916,N_18931);
or U19147 (N_19147,N_18857,N_18862);
nand U19148 (N_19148,N_18926,N_18836);
nor U19149 (N_19149,N_18885,N_18954);
xnor U19150 (N_19150,N_18932,N_18903);
xor U19151 (N_19151,N_18926,N_18820);
and U19152 (N_19152,N_18927,N_18983);
nand U19153 (N_19153,N_18948,N_18947);
nor U19154 (N_19154,N_18890,N_18864);
or U19155 (N_19155,N_18907,N_18881);
and U19156 (N_19156,N_18927,N_18836);
nor U19157 (N_19157,N_18965,N_18856);
nand U19158 (N_19158,N_18977,N_18815);
nand U19159 (N_19159,N_18945,N_18881);
nor U19160 (N_19160,N_18812,N_18995);
or U19161 (N_19161,N_18964,N_18958);
and U19162 (N_19162,N_18891,N_18850);
nor U19163 (N_19163,N_18865,N_18902);
or U19164 (N_19164,N_18853,N_18945);
xnor U19165 (N_19165,N_18806,N_18872);
and U19166 (N_19166,N_18876,N_18905);
and U19167 (N_19167,N_18939,N_18800);
nand U19168 (N_19168,N_18851,N_18888);
xor U19169 (N_19169,N_18963,N_18962);
and U19170 (N_19170,N_18854,N_18828);
nand U19171 (N_19171,N_18932,N_18837);
xor U19172 (N_19172,N_18959,N_18995);
or U19173 (N_19173,N_18866,N_18808);
xor U19174 (N_19174,N_18831,N_18957);
xnor U19175 (N_19175,N_18891,N_18920);
nand U19176 (N_19176,N_18945,N_18937);
or U19177 (N_19177,N_18801,N_18941);
or U19178 (N_19178,N_18989,N_18982);
or U19179 (N_19179,N_18870,N_18905);
nor U19180 (N_19180,N_18926,N_18956);
and U19181 (N_19181,N_18931,N_18938);
xnor U19182 (N_19182,N_18935,N_18920);
or U19183 (N_19183,N_18898,N_18964);
or U19184 (N_19184,N_18995,N_18878);
and U19185 (N_19185,N_18968,N_18972);
nor U19186 (N_19186,N_18821,N_18875);
nor U19187 (N_19187,N_18806,N_18853);
or U19188 (N_19188,N_18903,N_18951);
nor U19189 (N_19189,N_18811,N_18993);
or U19190 (N_19190,N_18909,N_18804);
or U19191 (N_19191,N_18974,N_18923);
nand U19192 (N_19192,N_18930,N_18906);
nor U19193 (N_19193,N_18964,N_18902);
or U19194 (N_19194,N_18930,N_18854);
nand U19195 (N_19195,N_18911,N_18997);
xnor U19196 (N_19196,N_18810,N_18998);
xor U19197 (N_19197,N_18813,N_18867);
nor U19198 (N_19198,N_18827,N_18957);
and U19199 (N_19199,N_18950,N_18858);
and U19200 (N_19200,N_19101,N_19097);
nor U19201 (N_19201,N_19107,N_19109);
xnor U19202 (N_19202,N_19060,N_19159);
or U19203 (N_19203,N_19055,N_19195);
or U19204 (N_19204,N_19182,N_19175);
nor U19205 (N_19205,N_19147,N_19019);
nand U19206 (N_19206,N_19098,N_19164);
or U19207 (N_19207,N_19002,N_19193);
xor U19208 (N_19208,N_19000,N_19033);
xnor U19209 (N_19209,N_19199,N_19194);
nor U19210 (N_19210,N_19054,N_19128);
and U19211 (N_19211,N_19025,N_19158);
or U19212 (N_19212,N_19137,N_19058);
and U19213 (N_19213,N_19040,N_19047);
nor U19214 (N_19214,N_19048,N_19134);
or U19215 (N_19215,N_19118,N_19069);
or U19216 (N_19216,N_19073,N_19132);
xor U19217 (N_19217,N_19150,N_19045);
and U19218 (N_19218,N_19029,N_19123);
xor U19219 (N_19219,N_19115,N_19064);
and U19220 (N_19220,N_19140,N_19066);
nor U19221 (N_19221,N_19136,N_19076);
nand U19222 (N_19222,N_19053,N_19014);
nand U19223 (N_19223,N_19056,N_19100);
nor U19224 (N_19224,N_19078,N_19007);
nor U19225 (N_19225,N_19166,N_19027);
nor U19226 (N_19226,N_19028,N_19016);
or U19227 (N_19227,N_19125,N_19050);
nand U19228 (N_19228,N_19059,N_19034);
nand U19229 (N_19229,N_19142,N_19011);
or U19230 (N_19230,N_19077,N_19186);
nor U19231 (N_19231,N_19157,N_19030);
or U19232 (N_19232,N_19152,N_19013);
and U19233 (N_19233,N_19044,N_19149);
xnor U19234 (N_19234,N_19088,N_19165);
nand U19235 (N_19235,N_19163,N_19075);
xnor U19236 (N_19236,N_19018,N_19169);
or U19237 (N_19237,N_19096,N_19192);
nor U19238 (N_19238,N_19086,N_19092);
and U19239 (N_19239,N_19198,N_19119);
nand U19240 (N_19240,N_19188,N_19015);
xnor U19241 (N_19241,N_19067,N_19191);
xnor U19242 (N_19242,N_19084,N_19057);
and U19243 (N_19243,N_19181,N_19174);
and U19244 (N_19244,N_19037,N_19062);
or U19245 (N_19245,N_19072,N_19139);
and U19246 (N_19246,N_19068,N_19083);
or U19247 (N_19247,N_19184,N_19041);
xnor U19248 (N_19248,N_19117,N_19120);
nand U19249 (N_19249,N_19110,N_19154);
and U19250 (N_19250,N_19035,N_19005);
or U19251 (N_19251,N_19144,N_19176);
or U19252 (N_19252,N_19189,N_19049);
xnor U19253 (N_19253,N_19099,N_19116);
or U19254 (N_19254,N_19087,N_19168);
or U19255 (N_19255,N_19008,N_19113);
xor U19256 (N_19256,N_19010,N_19180);
xnor U19257 (N_19257,N_19051,N_19052);
nand U19258 (N_19258,N_19197,N_19093);
or U19259 (N_19259,N_19124,N_19036);
nand U19260 (N_19260,N_19187,N_19082);
nand U19261 (N_19261,N_19039,N_19170);
nand U19262 (N_19262,N_19183,N_19004);
and U19263 (N_19263,N_19003,N_19009);
nand U19264 (N_19264,N_19114,N_19079);
xnor U19265 (N_19265,N_19141,N_19090);
and U19266 (N_19266,N_19063,N_19190);
xor U19267 (N_19267,N_19094,N_19111);
nor U19268 (N_19268,N_19177,N_19017);
nor U19269 (N_19269,N_19085,N_19091);
nor U19270 (N_19270,N_19167,N_19104);
and U19271 (N_19271,N_19185,N_19026);
xnor U19272 (N_19272,N_19106,N_19126);
and U19273 (N_19273,N_19074,N_19061);
xnor U19274 (N_19274,N_19133,N_19130);
nor U19275 (N_19275,N_19095,N_19138);
nand U19276 (N_19276,N_19179,N_19131);
or U19277 (N_19277,N_19032,N_19122);
xnor U19278 (N_19278,N_19038,N_19171);
or U19279 (N_19279,N_19155,N_19020);
nor U19280 (N_19280,N_19108,N_19151);
or U19281 (N_19281,N_19143,N_19178);
or U19282 (N_19282,N_19156,N_19112);
xor U19283 (N_19283,N_19162,N_19001);
nand U19284 (N_19284,N_19006,N_19146);
nor U19285 (N_19285,N_19089,N_19135);
xnor U19286 (N_19286,N_19071,N_19105);
nor U19287 (N_19287,N_19103,N_19196);
and U19288 (N_19288,N_19129,N_19021);
and U19289 (N_19289,N_19042,N_19127);
and U19290 (N_19290,N_19024,N_19022);
nand U19291 (N_19291,N_19081,N_19172);
nand U19292 (N_19292,N_19148,N_19023);
xor U19293 (N_19293,N_19043,N_19145);
and U19294 (N_19294,N_19102,N_19161);
nand U19295 (N_19295,N_19121,N_19031);
or U19296 (N_19296,N_19160,N_19065);
or U19297 (N_19297,N_19080,N_19070);
nand U19298 (N_19298,N_19173,N_19153);
nand U19299 (N_19299,N_19046,N_19012);
nor U19300 (N_19300,N_19054,N_19075);
nand U19301 (N_19301,N_19135,N_19022);
nand U19302 (N_19302,N_19122,N_19188);
or U19303 (N_19303,N_19006,N_19118);
nor U19304 (N_19304,N_19030,N_19193);
nand U19305 (N_19305,N_19141,N_19048);
xor U19306 (N_19306,N_19076,N_19089);
and U19307 (N_19307,N_19094,N_19108);
or U19308 (N_19308,N_19191,N_19035);
xor U19309 (N_19309,N_19077,N_19146);
nor U19310 (N_19310,N_19055,N_19102);
nor U19311 (N_19311,N_19034,N_19058);
xor U19312 (N_19312,N_19070,N_19193);
nand U19313 (N_19313,N_19009,N_19148);
and U19314 (N_19314,N_19103,N_19069);
and U19315 (N_19315,N_19149,N_19170);
nand U19316 (N_19316,N_19002,N_19020);
nand U19317 (N_19317,N_19070,N_19176);
xnor U19318 (N_19318,N_19184,N_19044);
nor U19319 (N_19319,N_19036,N_19004);
xnor U19320 (N_19320,N_19132,N_19053);
nand U19321 (N_19321,N_19198,N_19036);
and U19322 (N_19322,N_19064,N_19088);
nand U19323 (N_19323,N_19199,N_19043);
nor U19324 (N_19324,N_19123,N_19151);
nor U19325 (N_19325,N_19163,N_19118);
or U19326 (N_19326,N_19067,N_19163);
and U19327 (N_19327,N_19111,N_19149);
or U19328 (N_19328,N_19045,N_19133);
and U19329 (N_19329,N_19084,N_19193);
or U19330 (N_19330,N_19129,N_19060);
and U19331 (N_19331,N_19026,N_19197);
nor U19332 (N_19332,N_19150,N_19120);
and U19333 (N_19333,N_19111,N_19176);
and U19334 (N_19334,N_19141,N_19190);
or U19335 (N_19335,N_19124,N_19177);
or U19336 (N_19336,N_19107,N_19091);
nor U19337 (N_19337,N_19051,N_19115);
nand U19338 (N_19338,N_19108,N_19002);
xnor U19339 (N_19339,N_19002,N_19029);
nand U19340 (N_19340,N_19035,N_19105);
or U19341 (N_19341,N_19153,N_19047);
and U19342 (N_19342,N_19112,N_19002);
or U19343 (N_19343,N_19070,N_19015);
nor U19344 (N_19344,N_19028,N_19114);
and U19345 (N_19345,N_19169,N_19094);
or U19346 (N_19346,N_19082,N_19111);
and U19347 (N_19347,N_19030,N_19008);
nor U19348 (N_19348,N_19135,N_19006);
or U19349 (N_19349,N_19056,N_19111);
and U19350 (N_19350,N_19032,N_19066);
nor U19351 (N_19351,N_19114,N_19145);
and U19352 (N_19352,N_19073,N_19122);
xor U19353 (N_19353,N_19104,N_19108);
nand U19354 (N_19354,N_19044,N_19083);
and U19355 (N_19355,N_19042,N_19086);
nand U19356 (N_19356,N_19029,N_19158);
nor U19357 (N_19357,N_19028,N_19090);
or U19358 (N_19358,N_19072,N_19063);
or U19359 (N_19359,N_19117,N_19016);
and U19360 (N_19360,N_19019,N_19101);
or U19361 (N_19361,N_19074,N_19137);
and U19362 (N_19362,N_19139,N_19043);
xor U19363 (N_19363,N_19114,N_19105);
and U19364 (N_19364,N_19061,N_19048);
nand U19365 (N_19365,N_19090,N_19053);
nor U19366 (N_19366,N_19181,N_19124);
nand U19367 (N_19367,N_19046,N_19010);
xor U19368 (N_19368,N_19063,N_19145);
xor U19369 (N_19369,N_19001,N_19134);
nand U19370 (N_19370,N_19167,N_19125);
nand U19371 (N_19371,N_19148,N_19112);
nand U19372 (N_19372,N_19184,N_19159);
xnor U19373 (N_19373,N_19046,N_19187);
nand U19374 (N_19374,N_19098,N_19125);
nor U19375 (N_19375,N_19017,N_19013);
or U19376 (N_19376,N_19166,N_19037);
and U19377 (N_19377,N_19027,N_19109);
or U19378 (N_19378,N_19023,N_19062);
or U19379 (N_19379,N_19170,N_19063);
nand U19380 (N_19380,N_19194,N_19032);
and U19381 (N_19381,N_19043,N_19026);
and U19382 (N_19382,N_19160,N_19028);
and U19383 (N_19383,N_19175,N_19147);
and U19384 (N_19384,N_19091,N_19147);
nor U19385 (N_19385,N_19039,N_19120);
xor U19386 (N_19386,N_19078,N_19103);
nand U19387 (N_19387,N_19019,N_19146);
or U19388 (N_19388,N_19179,N_19074);
nand U19389 (N_19389,N_19139,N_19171);
xnor U19390 (N_19390,N_19037,N_19010);
and U19391 (N_19391,N_19130,N_19015);
and U19392 (N_19392,N_19114,N_19092);
and U19393 (N_19393,N_19089,N_19144);
nand U19394 (N_19394,N_19107,N_19124);
nor U19395 (N_19395,N_19015,N_19195);
and U19396 (N_19396,N_19117,N_19097);
nand U19397 (N_19397,N_19086,N_19197);
nor U19398 (N_19398,N_19154,N_19044);
nand U19399 (N_19399,N_19157,N_19072);
nand U19400 (N_19400,N_19313,N_19286);
nor U19401 (N_19401,N_19222,N_19256);
nand U19402 (N_19402,N_19228,N_19387);
xor U19403 (N_19403,N_19365,N_19224);
xnor U19404 (N_19404,N_19221,N_19367);
or U19405 (N_19405,N_19237,N_19219);
xor U19406 (N_19406,N_19346,N_19381);
nor U19407 (N_19407,N_19333,N_19382);
and U19408 (N_19408,N_19397,N_19218);
and U19409 (N_19409,N_19220,N_19312);
nand U19410 (N_19410,N_19372,N_19244);
nor U19411 (N_19411,N_19285,N_19206);
nor U19412 (N_19412,N_19262,N_19388);
or U19413 (N_19413,N_19385,N_19287);
xnor U19414 (N_19414,N_19263,N_19343);
or U19415 (N_19415,N_19317,N_19309);
xnor U19416 (N_19416,N_19215,N_19281);
xnor U19417 (N_19417,N_19214,N_19230);
or U19418 (N_19418,N_19362,N_19366);
nand U19419 (N_19419,N_19339,N_19208);
nor U19420 (N_19420,N_19245,N_19261);
xor U19421 (N_19421,N_19269,N_19352);
nor U19422 (N_19422,N_19384,N_19297);
nand U19423 (N_19423,N_19279,N_19329);
xnor U19424 (N_19424,N_19351,N_19247);
nand U19425 (N_19425,N_19307,N_19373);
and U19426 (N_19426,N_19341,N_19389);
and U19427 (N_19427,N_19283,N_19310);
nor U19428 (N_19428,N_19213,N_19315);
xnor U19429 (N_19429,N_19212,N_19254);
xor U19430 (N_19430,N_19340,N_19334);
and U19431 (N_19431,N_19327,N_19396);
nor U19432 (N_19432,N_19233,N_19235);
nor U19433 (N_19433,N_19209,N_19326);
and U19434 (N_19434,N_19399,N_19350);
and U19435 (N_19435,N_19332,N_19304);
nand U19436 (N_19436,N_19328,N_19272);
and U19437 (N_19437,N_19330,N_19395);
nand U19438 (N_19438,N_19318,N_19374);
nor U19439 (N_19439,N_19303,N_19299);
nand U19440 (N_19440,N_19282,N_19386);
xor U19441 (N_19441,N_19205,N_19323);
and U19442 (N_19442,N_19277,N_19398);
nor U19443 (N_19443,N_19391,N_19360);
nor U19444 (N_19444,N_19377,N_19308);
and U19445 (N_19445,N_19241,N_19371);
and U19446 (N_19446,N_19324,N_19336);
nand U19447 (N_19447,N_19246,N_19335);
nor U19448 (N_19448,N_19204,N_19364);
and U19449 (N_19449,N_19289,N_19311);
or U19450 (N_19450,N_19216,N_19240);
nor U19451 (N_19451,N_19376,N_19211);
nand U19452 (N_19452,N_19257,N_19268);
or U19453 (N_19453,N_19255,N_19363);
and U19454 (N_19454,N_19345,N_19202);
and U19455 (N_19455,N_19242,N_19280);
and U19456 (N_19456,N_19319,N_19349);
nor U19457 (N_19457,N_19200,N_19270);
xor U19458 (N_19458,N_19260,N_19347);
nor U19459 (N_19459,N_19267,N_19316);
nand U19460 (N_19460,N_19232,N_19293);
xnor U19461 (N_19461,N_19288,N_19253);
or U19462 (N_19462,N_19207,N_19203);
xnor U19463 (N_19463,N_19301,N_19251);
or U19464 (N_19464,N_19306,N_19383);
and U19465 (N_19465,N_19201,N_19266);
xor U19466 (N_19466,N_19264,N_19338);
nand U19467 (N_19467,N_19325,N_19356);
xor U19468 (N_19468,N_19295,N_19357);
nor U19469 (N_19469,N_19231,N_19210);
nand U19470 (N_19470,N_19348,N_19234);
nor U19471 (N_19471,N_19358,N_19226);
xnor U19472 (N_19472,N_19322,N_19342);
nand U19473 (N_19473,N_19380,N_19271);
nand U19474 (N_19474,N_19331,N_19393);
nor U19475 (N_19475,N_19298,N_19278);
or U19476 (N_19476,N_19248,N_19225);
nand U19477 (N_19477,N_19274,N_19392);
or U19478 (N_19478,N_19300,N_19249);
nor U19479 (N_19479,N_19223,N_19259);
and U19480 (N_19480,N_19292,N_19337);
nor U19481 (N_19481,N_19229,N_19361);
or U19482 (N_19482,N_19321,N_19217);
and U19483 (N_19483,N_19344,N_19305);
and U19484 (N_19484,N_19276,N_19375);
and U19485 (N_19485,N_19284,N_19353);
xor U19486 (N_19486,N_19368,N_19243);
or U19487 (N_19487,N_19290,N_19291);
nand U19488 (N_19488,N_19252,N_19354);
xnor U19489 (N_19489,N_19320,N_19355);
or U19490 (N_19490,N_19294,N_19227);
xnor U19491 (N_19491,N_19370,N_19302);
and U19492 (N_19492,N_19314,N_19273);
and U19493 (N_19493,N_19369,N_19378);
xnor U19494 (N_19494,N_19265,N_19390);
nand U19495 (N_19495,N_19359,N_19236);
nand U19496 (N_19496,N_19239,N_19379);
nand U19497 (N_19497,N_19296,N_19258);
nand U19498 (N_19498,N_19250,N_19275);
xnor U19499 (N_19499,N_19238,N_19394);
nor U19500 (N_19500,N_19231,N_19385);
or U19501 (N_19501,N_19282,N_19264);
nand U19502 (N_19502,N_19262,N_19354);
xor U19503 (N_19503,N_19242,N_19357);
and U19504 (N_19504,N_19392,N_19355);
or U19505 (N_19505,N_19309,N_19221);
xor U19506 (N_19506,N_19334,N_19365);
nand U19507 (N_19507,N_19322,N_19291);
nand U19508 (N_19508,N_19297,N_19393);
nand U19509 (N_19509,N_19282,N_19208);
xor U19510 (N_19510,N_19240,N_19360);
xnor U19511 (N_19511,N_19342,N_19369);
xnor U19512 (N_19512,N_19231,N_19214);
nor U19513 (N_19513,N_19396,N_19306);
and U19514 (N_19514,N_19384,N_19222);
or U19515 (N_19515,N_19256,N_19321);
and U19516 (N_19516,N_19210,N_19223);
and U19517 (N_19517,N_19276,N_19367);
nand U19518 (N_19518,N_19372,N_19397);
nand U19519 (N_19519,N_19250,N_19320);
and U19520 (N_19520,N_19254,N_19290);
and U19521 (N_19521,N_19382,N_19271);
or U19522 (N_19522,N_19338,N_19234);
and U19523 (N_19523,N_19339,N_19397);
xor U19524 (N_19524,N_19313,N_19363);
nor U19525 (N_19525,N_19252,N_19264);
and U19526 (N_19526,N_19318,N_19308);
nor U19527 (N_19527,N_19219,N_19302);
nand U19528 (N_19528,N_19316,N_19327);
xor U19529 (N_19529,N_19281,N_19375);
xnor U19530 (N_19530,N_19352,N_19243);
or U19531 (N_19531,N_19253,N_19254);
and U19532 (N_19532,N_19356,N_19226);
or U19533 (N_19533,N_19307,N_19323);
and U19534 (N_19534,N_19304,N_19293);
and U19535 (N_19535,N_19390,N_19329);
and U19536 (N_19536,N_19278,N_19295);
and U19537 (N_19537,N_19217,N_19326);
or U19538 (N_19538,N_19370,N_19235);
or U19539 (N_19539,N_19357,N_19330);
and U19540 (N_19540,N_19325,N_19309);
nor U19541 (N_19541,N_19230,N_19350);
or U19542 (N_19542,N_19285,N_19231);
or U19543 (N_19543,N_19243,N_19317);
nor U19544 (N_19544,N_19321,N_19272);
nand U19545 (N_19545,N_19385,N_19213);
nor U19546 (N_19546,N_19200,N_19379);
or U19547 (N_19547,N_19208,N_19318);
nor U19548 (N_19548,N_19282,N_19238);
xnor U19549 (N_19549,N_19229,N_19299);
xor U19550 (N_19550,N_19273,N_19260);
xor U19551 (N_19551,N_19384,N_19315);
nand U19552 (N_19552,N_19323,N_19249);
nor U19553 (N_19553,N_19333,N_19242);
and U19554 (N_19554,N_19312,N_19291);
and U19555 (N_19555,N_19359,N_19283);
nand U19556 (N_19556,N_19352,N_19256);
nand U19557 (N_19557,N_19216,N_19377);
nor U19558 (N_19558,N_19214,N_19247);
or U19559 (N_19559,N_19336,N_19247);
nor U19560 (N_19560,N_19272,N_19390);
nor U19561 (N_19561,N_19208,N_19247);
xnor U19562 (N_19562,N_19355,N_19372);
nor U19563 (N_19563,N_19215,N_19256);
and U19564 (N_19564,N_19341,N_19216);
and U19565 (N_19565,N_19220,N_19259);
or U19566 (N_19566,N_19263,N_19354);
and U19567 (N_19567,N_19239,N_19371);
nor U19568 (N_19568,N_19379,N_19259);
and U19569 (N_19569,N_19361,N_19336);
and U19570 (N_19570,N_19372,N_19292);
xnor U19571 (N_19571,N_19319,N_19288);
nand U19572 (N_19572,N_19264,N_19383);
xnor U19573 (N_19573,N_19247,N_19233);
xnor U19574 (N_19574,N_19383,N_19273);
nand U19575 (N_19575,N_19315,N_19379);
and U19576 (N_19576,N_19374,N_19329);
or U19577 (N_19577,N_19279,N_19270);
and U19578 (N_19578,N_19247,N_19341);
nand U19579 (N_19579,N_19321,N_19368);
nor U19580 (N_19580,N_19345,N_19237);
nand U19581 (N_19581,N_19331,N_19334);
nand U19582 (N_19582,N_19208,N_19244);
xnor U19583 (N_19583,N_19354,N_19397);
and U19584 (N_19584,N_19324,N_19268);
or U19585 (N_19585,N_19211,N_19251);
nor U19586 (N_19586,N_19342,N_19373);
nand U19587 (N_19587,N_19321,N_19386);
or U19588 (N_19588,N_19305,N_19215);
xnor U19589 (N_19589,N_19251,N_19349);
nor U19590 (N_19590,N_19282,N_19227);
or U19591 (N_19591,N_19313,N_19347);
nor U19592 (N_19592,N_19267,N_19388);
or U19593 (N_19593,N_19293,N_19313);
nor U19594 (N_19594,N_19351,N_19230);
or U19595 (N_19595,N_19229,N_19274);
or U19596 (N_19596,N_19367,N_19252);
nor U19597 (N_19597,N_19357,N_19249);
xnor U19598 (N_19598,N_19203,N_19397);
or U19599 (N_19599,N_19281,N_19351);
or U19600 (N_19600,N_19554,N_19436);
and U19601 (N_19601,N_19502,N_19401);
or U19602 (N_19602,N_19570,N_19548);
nand U19603 (N_19603,N_19578,N_19531);
and U19604 (N_19604,N_19525,N_19439);
nor U19605 (N_19605,N_19585,N_19566);
and U19606 (N_19606,N_19595,N_19455);
nand U19607 (N_19607,N_19416,N_19581);
or U19608 (N_19608,N_19557,N_19438);
xor U19609 (N_19609,N_19434,N_19582);
nor U19610 (N_19610,N_19500,N_19551);
xnor U19611 (N_19611,N_19547,N_19543);
nand U19612 (N_19612,N_19404,N_19597);
nand U19613 (N_19613,N_19486,N_19481);
and U19614 (N_19614,N_19411,N_19428);
and U19615 (N_19615,N_19544,N_19587);
and U19616 (N_19616,N_19424,N_19476);
and U19617 (N_19617,N_19599,N_19556);
or U19618 (N_19618,N_19496,N_19508);
nor U19619 (N_19619,N_19490,N_19425);
and U19620 (N_19620,N_19560,N_19541);
nand U19621 (N_19621,N_19452,N_19563);
nand U19622 (N_19622,N_19503,N_19586);
nand U19623 (N_19623,N_19528,N_19464);
nand U19624 (N_19624,N_19542,N_19433);
and U19625 (N_19625,N_19406,N_19461);
nand U19626 (N_19626,N_19443,N_19475);
xor U19627 (N_19627,N_19492,N_19545);
and U19628 (N_19628,N_19407,N_19419);
and U19629 (N_19629,N_19482,N_19524);
nand U19630 (N_19630,N_19400,N_19403);
and U19631 (N_19631,N_19555,N_19479);
or U19632 (N_19632,N_19409,N_19571);
or U19633 (N_19633,N_19483,N_19565);
nor U19634 (N_19634,N_19501,N_19539);
nor U19635 (N_19635,N_19512,N_19444);
xor U19636 (N_19636,N_19511,N_19460);
and U19637 (N_19637,N_19523,N_19598);
nand U19638 (N_19638,N_19580,N_19450);
or U19639 (N_19639,N_19402,N_19510);
or U19640 (N_19640,N_19442,N_19575);
or U19641 (N_19641,N_19579,N_19453);
nor U19642 (N_19642,N_19474,N_19536);
xor U19643 (N_19643,N_19499,N_19538);
xor U19644 (N_19644,N_19408,N_19412);
nand U19645 (N_19645,N_19505,N_19413);
nand U19646 (N_19646,N_19430,N_19520);
xnor U19647 (N_19647,N_19540,N_19447);
and U19648 (N_19648,N_19445,N_19488);
nor U19649 (N_19649,N_19515,N_19405);
nor U19650 (N_19650,N_19569,N_19534);
and U19651 (N_19651,N_19417,N_19590);
or U19652 (N_19652,N_19494,N_19509);
and U19653 (N_19653,N_19414,N_19584);
or U19654 (N_19654,N_19521,N_19415);
and U19655 (N_19655,N_19431,N_19574);
xnor U19656 (N_19656,N_19507,N_19550);
nor U19657 (N_19657,N_19418,N_19420);
and U19658 (N_19658,N_19456,N_19589);
nand U19659 (N_19659,N_19459,N_19532);
xnor U19660 (N_19660,N_19546,N_19469);
nor U19661 (N_19661,N_19498,N_19465);
xnor U19662 (N_19662,N_19593,N_19427);
nand U19663 (N_19663,N_19463,N_19491);
nor U19664 (N_19664,N_19559,N_19468);
and U19665 (N_19665,N_19567,N_19564);
xnor U19666 (N_19666,N_19596,N_19526);
or U19667 (N_19667,N_19583,N_19485);
nand U19668 (N_19668,N_19487,N_19529);
and U19669 (N_19669,N_19517,N_19519);
nand U19670 (N_19670,N_19467,N_19588);
or U19671 (N_19671,N_19426,N_19489);
nand U19672 (N_19672,N_19423,N_19535);
nor U19673 (N_19673,N_19440,N_19594);
or U19674 (N_19674,N_19449,N_19454);
and U19675 (N_19675,N_19495,N_19533);
nand U19676 (N_19676,N_19527,N_19576);
xnor U19677 (N_19677,N_19561,N_19516);
nand U19678 (N_19678,N_19421,N_19522);
xnor U19679 (N_19679,N_19429,N_19506);
nand U19680 (N_19680,N_19549,N_19473);
nand U19681 (N_19681,N_19472,N_19466);
xnor U19682 (N_19682,N_19514,N_19537);
and U19683 (N_19683,N_19553,N_19441);
xor U19684 (N_19684,N_19591,N_19458);
or U19685 (N_19685,N_19470,N_19432);
and U19686 (N_19686,N_19462,N_19504);
nand U19687 (N_19687,N_19530,N_19577);
or U19688 (N_19688,N_19477,N_19562);
or U19689 (N_19689,N_19446,N_19572);
xor U19690 (N_19690,N_19410,N_19457);
xnor U19691 (N_19691,N_19573,N_19513);
or U19692 (N_19692,N_19451,N_19480);
nand U19693 (N_19693,N_19471,N_19435);
xnor U19694 (N_19694,N_19592,N_19478);
and U19695 (N_19695,N_19497,N_19568);
nand U19696 (N_19696,N_19437,N_19448);
nor U19697 (N_19697,N_19552,N_19484);
or U19698 (N_19698,N_19493,N_19518);
nand U19699 (N_19699,N_19558,N_19422);
and U19700 (N_19700,N_19475,N_19480);
nor U19701 (N_19701,N_19431,N_19587);
and U19702 (N_19702,N_19449,N_19430);
nand U19703 (N_19703,N_19574,N_19568);
xor U19704 (N_19704,N_19536,N_19599);
or U19705 (N_19705,N_19565,N_19596);
nor U19706 (N_19706,N_19549,N_19563);
nand U19707 (N_19707,N_19449,N_19555);
xor U19708 (N_19708,N_19477,N_19513);
or U19709 (N_19709,N_19529,N_19533);
xnor U19710 (N_19710,N_19484,N_19536);
or U19711 (N_19711,N_19453,N_19409);
nand U19712 (N_19712,N_19442,N_19574);
nand U19713 (N_19713,N_19517,N_19583);
or U19714 (N_19714,N_19515,N_19580);
xnor U19715 (N_19715,N_19419,N_19464);
nor U19716 (N_19716,N_19470,N_19469);
and U19717 (N_19717,N_19441,N_19401);
and U19718 (N_19718,N_19589,N_19524);
xor U19719 (N_19719,N_19425,N_19575);
nor U19720 (N_19720,N_19590,N_19543);
or U19721 (N_19721,N_19477,N_19585);
nor U19722 (N_19722,N_19420,N_19487);
nor U19723 (N_19723,N_19484,N_19578);
nor U19724 (N_19724,N_19529,N_19559);
xnor U19725 (N_19725,N_19414,N_19494);
or U19726 (N_19726,N_19460,N_19538);
nor U19727 (N_19727,N_19430,N_19494);
xor U19728 (N_19728,N_19554,N_19494);
or U19729 (N_19729,N_19596,N_19443);
or U19730 (N_19730,N_19457,N_19517);
nor U19731 (N_19731,N_19577,N_19411);
or U19732 (N_19732,N_19434,N_19544);
nor U19733 (N_19733,N_19533,N_19488);
or U19734 (N_19734,N_19575,N_19471);
and U19735 (N_19735,N_19436,N_19576);
nor U19736 (N_19736,N_19542,N_19480);
and U19737 (N_19737,N_19549,N_19409);
xor U19738 (N_19738,N_19509,N_19468);
xnor U19739 (N_19739,N_19549,N_19450);
and U19740 (N_19740,N_19440,N_19533);
xnor U19741 (N_19741,N_19411,N_19552);
xor U19742 (N_19742,N_19501,N_19574);
or U19743 (N_19743,N_19546,N_19587);
xor U19744 (N_19744,N_19517,N_19471);
nand U19745 (N_19745,N_19522,N_19572);
nor U19746 (N_19746,N_19577,N_19462);
or U19747 (N_19747,N_19597,N_19414);
nand U19748 (N_19748,N_19491,N_19468);
or U19749 (N_19749,N_19527,N_19489);
or U19750 (N_19750,N_19467,N_19412);
xnor U19751 (N_19751,N_19460,N_19578);
xor U19752 (N_19752,N_19561,N_19526);
or U19753 (N_19753,N_19555,N_19455);
or U19754 (N_19754,N_19523,N_19436);
or U19755 (N_19755,N_19427,N_19445);
nand U19756 (N_19756,N_19552,N_19579);
nor U19757 (N_19757,N_19475,N_19560);
xor U19758 (N_19758,N_19438,N_19564);
and U19759 (N_19759,N_19500,N_19513);
and U19760 (N_19760,N_19426,N_19507);
or U19761 (N_19761,N_19528,N_19500);
xnor U19762 (N_19762,N_19454,N_19583);
nor U19763 (N_19763,N_19528,N_19486);
or U19764 (N_19764,N_19461,N_19504);
or U19765 (N_19765,N_19413,N_19548);
or U19766 (N_19766,N_19493,N_19405);
nor U19767 (N_19767,N_19449,N_19509);
or U19768 (N_19768,N_19407,N_19577);
or U19769 (N_19769,N_19550,N_19514);
and U19770 (N_19770,N_19474,N_19589);
or U19771 (N_19771,N_19539,N_19434);
and U19772 (N_19772,N_19405,N_19514);
and U19773 (N_19773,N_19444,N_19482);
nand U19774 (N_19774,N_19508,N_19542);
xor U19775 (N_19775,N_19471,N_19436);
and U19776 (N_19776,N_19584,N_19549);
xor U19777 (N_19777,N_19468,N_19454);
or U19778 (N_19778,N_19558,N_19580);
xnor U19779 (N_19779,N_19580,N_19485);
nand U19780 (N_19780,N_19443,N_19577);
and U19781 (N_19781,N_19517,N_19480);
nor U19782 (N_19782,N_19585,N_19581);
nor U19783 (N_19783,N_19525,N_19499);
nand U19784 (N_19784,N_19474,N_19596);
nor U19785 (N_19785,N_19457,N_19475);
or U19786 (N_19786,N_19525,N_19514);
or U19787 (N_19787,N_19581,N_19463);
nor U19788 (N_19788,N_19529,N_19485);
nor U19789 (N_19789,N_19437,N_19563);
nand U19790 (N_19790,N_19463,N_19554);
nor U19791 (N_19791,N_19581,N_19406);
or U19792 (N_19792,N_19405,N_19580);
or U19793 (N_19793,N_19512,N_19445);
or U19794 (N_19794,N_19514,N_19433);
xor U19795 (N_19795,N_19580,N_19442);
xnor U19796 (N_19796,N_19443,N_19529);
and U19797 (N_19797,N_19415,N_19419);
nor U19798 (N_19798,N_19520,N_19579);
nand U19799 (N_19799,N_19454,N_19473);
and U19800 (N_19800,N_19667,N_19728);
nand U19801 (N_19801,N_19738,N_19633);
nand U19802 (N_19802,N_19699,N_19772);
xnor U19803 (N_19803,N_19692,N_19736);
nand U19804 (N_19804,N_19670,N_19799);
nand U19805 (N_19805,N_19601,N_19602);
xor U19806 (N_19806,N_19747,N_19631);
nor U19807 (N_19807,N_19744,N_19698);
or U19808 (N_19808,N_19794,N_19659);
xor U19809 (N_19809,N_19748,N_19608);
and U19810 (N_19810,N_19788,N_19790);
nand U19811 (N_19811,N_19739,N_19662);
nand U19812 (N_19812,N_19796,N_19664);
nor U19813 (N_19813,N_19716,N_19792);
or U19814 (N_19814,N_19787,N_19672);
and U19815 (N_19815,N_19759,N_19785);
nor U19816 (N_19816,N_19732,N_19720);
and U19817 (N_19817,N_19690,N_19719);
nand U19818 (N_19818,N_19758,N_19705);
nand U19819 (N_19819,N_19707,N_19613);
or U19820 (N_19820,N_19714,N_19756);
nand U19821 (N_19821,N_19770,N_19789);
and U19822 (N_19822,N_19773,N_19786);
and U19823 (N_19823,N_19767,N_19763);
and U19824 (N_19824,N_19777,N_19614);
and U19825 (N_19825,N_19686,N_19691);
or U19826 (N_19826,N_19679,N_19771);
nand U19827 (N_19827,N_19766,N_19656);
nor U19828 (N_19828,N_19685,N_19626);
xor U19829 (N_19829,N_19717,N_19625);
or U19830 (N_19830,N_19791,N_19635);
and U19831 (N_19831,N_19652,N_19702);
and U19832 (N_19832,N_19798,N_19693);
nand U19833 (N_19833,N_19768,N_19715);
xor U19834 (N_19834,N_19610,N_19774);
nand U19835 (N_19835,N_19761,N_19751);
nand U19836 (N_19836,N_19629,N_19755);
and U19837 (N_19837,N_19673,N_19658);
xor U19838 (N_19838,N_19764,N_19666);
xor U19839 (N_19839,N_19797,N_19710);
xnor U19840 (N_19840,N_19653,N_19703);
and U19841 (N_19841,N_19754,N_19655);
and U19842 (N_19842,N_19776,N_19628);
xnor U19843 (N_19843,N_19600,N_19606);
nor U19844 (N_19844,N_19731,N_19654);
or U19845 (N_19845,N_19639,N_19750);
nand U19846 (N_19846,N_19603,N_19607);
nand U19847 (N_19847,N_19795,N_19627);
xor U19848 (N_19848,N_19638,N_19641);
nand U19849 (N_19849,N_19650,N_19780);
xor U19850 (N_19850,N_19649,N_19630);
nand U19851 (N_19851,N_19682,N_19783);
and U19852 (N_19852,N_19793,N_19697);
or U19853 (N_19853,N_19746,N_19676);
nand U19854 (N_19854,N_19733,N_19651);
nor U19855 (N_19855,N_19713,N_19604);
and U19856 (N_19856,N_19729,N_19752);
xnor U19857 (N_19857,N_19619,N_19660);
and U19858 (N_19858,N_19678,N_19760);
nor U19859 (N_19859,N_19645,N_19712);
nand U19860 (N_19860,N_19727,N_19680);
nor U19861 (N_19861,N_19643,N_19632);
nor U19862 (N_19862,N_19701,N_19779);
xor U19863 (N_19863,N_19674,N_19784);
xnor U19864 (N_19864,N_19735,N_19725);
nor U19865 (N_19865,N_19743,N_19623);
xor U19866 (N_19866,N_19708,N_19694);
nor U19867 (N_19867,N_19669,N_19657);
nor U19868 (N_19868,N_19737,N_19637);
nor U19869 (N_19869,N_19778,N_19683);
nor U19870 (N_19870,N_19769,N_19688);
and U19871 (N_19871,N_19695,N_19681);
xor U19872 (N_19872,N_19616,N_19668);
or U19873 (N_19873,N_19782,N_19700);
xor U19874 (N_19874,N_19711,N_19765);
or U19875 (N_19875,N_19696,N_19734);
and U19876 (N_19876,N_19661,N_19742);
or U19877 (N_19877,N_19724,N_19675);
nor U19878 (N_19878,N_19726,N_19636);
xnor U19879 (N_19879,N_19706,N_19644);
nand U19880 (N_19880,N_19611,N_19721);
nor U19881 (N_19881,N_19687,N_19689);
xnor U19882 (N_19882,N_19745,N_19762);
nand U19883 (N_19883,N_19722,N_19640);
and U19884 (N_19884,N_19753,N_19634);
nand U19885 (N_19885,N_19618,N_19757);
and U19886 (N_19886,N_19740,N_19749);
and U19887 (N_19887,N_19609,N_19647);
nand U19888 (N_19888,N_19615,N_19677);
xnor U19889 (N_19889,N_19612,N_19730);
xor U19890 (N_19890,N_19704,N_19663);
and U19891 (N_19891,N_19621,N_19646);
and U19892 (N_19892,N_19622,N_19718);
or U19893 (N_19893,N_19620,N_19723);
or U19894 (N_19894,N_19781,N_19741);
and U19895 (N_19895,N_19671,N_19684);
and U19896 (N_19896,N_19617,N_19775);
or U19897 (N_19897,N_19665,N_19642);
and U19898 (N_19898,N_19709,N_19605);
xor U19899 (N_19899,N_19648,N_19624);
xor U19900 (N_19900,N_19763,N_19609);
xor U19901 (N_19901,N_19797,N_19777);
nor U19902 (N_19902,N_19611,N_19650);
nand U19903 (N_19903,N_19668,N_19729);
nor U19904 (N_19904,N_19710,N_19642);
nand U19905 (N_19905,N_19612,N_19611);
or U19906 (N_19906,N_19717,N_19610);
or U19907 (N_19907,N_19787,N_19798);
nor U19908 (N_19908,N_19643,N_19759);
or U19909 (N_19909,N_19764,N_19609);
nor U19910 (N_19910,N_19797,N_19654);
nor U19911 (N_19911,N_19746,N_19708);
xnor U19912 (N_19912,N_19652,N_19712);
and U19913 (N_19913,N_19763,N_19652);
or U19914 (N_19914,N_19606,N_19757);
nor U19915 (N_19915,N_19627,N_19738);
nand U19916 (N_19916,N_19634,N_19681);
nor U19917 (N_19917,N_19686,N_19651);
nand U19918 (N_19918,N_19742,N_19613);
nand U19919 (N_19919,N_19668,N_19667);
nor U19920 (N_19920,N_19762,N_19679);
and U19921 (N_19921,N_19660,N_19659);
nor U19922 (N_19922,N_19786,N_19746);
or U19923 (N_19923,N_19724,N_19608);
xnor U19924 (N_19924,N_19677,N_19623);
xnor U19925 (N_19925,N_19710,N_19681);
and U19926 (N_19926,N_19705,N_19772);
or U19927 (N_19927,N_19784,N_19778);
nand U19928 (N_19928,N_19700,N_19783);
nand U19929 (N_19929,N_19697,N_19658);
nor U19930 (N_19930,N_19744,N_19770);
and U19931 (N_19931,N_19723,N_19767);
or U19932 (N_19932,N_19758,N_19747);
nor U19933 (N_19933,N_19694,N_19754);
nor U19934 (N_19934,N_19633,N_19674);
and U19935 (N_19935,N_19624,N_19770);
and U19936 (N_19936,N_19620,N_19631);
or U19937 (N_19937,N_19668,N_19653);
nor U19938 (N_19938,N_19607,N_19797);
xnor U19939 (N_19939,N_19780,N_19782);
xnor U19940 (N_19940,N_19643,N_19687);
nor U19941 (N_19941,N_19676,N_19661);
xnor U19942 (N_19942,N_19613,N_19773);
or U19943 (N_19943,N_19631,N_19642);
nand U19944 (N_19944,N_19699,N_19794);
xnor U19945 (N_19945,N_19720,N_19666);
and U19946 (N_19946,N_19698,N_19621);
nand U19947 (N_19947,N_19621,N_19637);
xor U19948 (N_19948,N_19755,N_19686);
or U19949 (N_19949,N_19634,N_19617);
nand U19950 (N_19950,N_19645,N_19707);
nor U19951 (N_19951,N_19627,N_19765);
nand U19952 (N_19952,N_19610,N_19622);
xnor U19953 (N_19953,N_19785,N_19755);
nand U19954 (N_19954,N_19765,N_19652);
xnor U19955 (N_19955,N_19653,N_19600);
nor U19956 (N_19956,N_19752,N_19619);
xnor U19957 (N_19957,N_19648,N_19691);
and U19958 (N_19958,N_19775,N_19654);
and U19959 (N_19959,N_19746,N_19618);
nor U19960 (N_19960,N_19711,N_19710);
xnor U19961 (N_19961,N_19746,N_19740);
or U19962 (N_19962,N_19777,N_19666);
or U19963 (N_19963,N_19679,N_19631);
nor U19964 (N_19964,N_19607,N_19753);
and U19965 (N_19965,N_19781,N_19788);
xnor U19966 (N_19966,N_19700,N_19723);
or U19967 (N_19967,N_19716,N_19708);
or U19968 (N_19968,N_19641,N_19693);
or U19969 (N_19969,N_19704,N_19785);
and U19970 (N_19970,N_19622,N_19761);
and U19971 (N_19971,N_19637,N_19706);
and U19972 (N_19972,N_19690,N_19710);
or U19973 (N_19973,N_19693,N_19752);
nor U19974 (N_19974,N_19685,N_19763);
nand U19975 (N_19975,N_19767,N_19697);
and U19976 (N_19976,N_19687,N_19739);
nor U19977 (N_19977,N_19777,N_19602);
and U19978 (N_19978,N_19799,N_19755);
and U19979 (N_19979,N_19685,N_19724);
and U19980 (N_19980,N_19676,N_19791);
or U19981 (N_19981,N_19619,N_19615);
xnor U19982 (N_19982,N_19736,N_19784);
nor U19983 (N_19983,N_19763,N_19728);
or U19984 (N_19984,N_19612,N_19789);
or U19985 (N_19985,N_19771,N_19737);
and U19986 (N_19986,N_19675,N_19690);
or U19987 (N_19987,N_19651,N_19670);
nor U19988 (N_19988,N_19653,N_19773);
xor U19989 (N_19989,N_19623,N_19733);
or U19990 (N_19990,N_19779,N_19744);
nand U19991 (N_19991,N_19631,N_19734);
and U19992 (N_19992,N_19771,N_19685);
nand U19993 (N_19993,N_19618,N_19689);
xnor U19994 (N_19994,N_19714,N_19799);
nor U19995 (N_19995,N_19716,N_19799);
or U19996 (N_19996,N_19678,N_19672);
xnor U19997 (N_19997,N_19749,N_19772);
nor U19998 (N_19998,N_19627,N_19617);
or U19999 (N_19999,N_19752,N_19742);
nand U20000 (N_20000,N_19909,N_19947);
xnor U20001 (N_20001,N_19844,N_19891);
nor U20002 (N_20002,N_19881,N_19828);
nor U20003 (N_20003,N_19916,N_19813);
xnor U20004 (N_20004,N_19923,N_19900);
nand U20005 (N_20005,N_19806,N_19904);
nor U20006 (N_20006,N_19808,N_19972);
xnor U20007 (N_20007,N_19886,N_19819);
nand U20008 (N_20008,N_19832,N_19801);
nor U20009 (N_20009,N_19931,N_19982);
and U20010 (N_20010,N_19902,N_19905);
or U20011 (N_20011,N_19892,N_19889);
nand U20012 (N_20012,N_19814,N_19864);
and U20013 (N_20013,N_19994,N_19876);
or U20014 (N_20014,N_19924,N_19897);
xnor U20015 (N_20015,N_19885,N_19937);
and U20016 (N_20016,N_19936,N_19996);
and U20017 (N_20017,N_19861,N_19811);
and U20018 (N_20018,N_19848,N_19835);
and U20019 (N_20019,N_19884,N_19855);
or U20020 (N_20020,N_19988,N_19875);
xnor U20021 (N_20021,N_19986,N_19925);
or U20022 (N_20022,N_19944,N_19860);
and U20023 (N_20023,N_19825,N_19997);
xnor U20024 (N_20024,N_19852,N_19822);
and U20025 (N_20025,N_19846,N_19817);
and U20026 (N_20026,N_19823,N_19973);
xor U20027 (N_20027,N_19950,N_19847);
or U20028 (N_20028,N_19922,N_19815);
xor U20029 (N_20029,N_19901,N_19887);
or U20030 (N_20030,N_19995,N_19841);
nand U20031 (N_20031,N_19963,N_19839);
and U20032 (N_20032,N_19927,N_19976);
xnor U20033 (N_20033,N_19890,N_19962);
and U20034 (N_20034,N_19859,N_19858);
nor U20035 (N_20035,N_19809,N_19940);
nand U20036 (N_20036,N_19802,N_19998);
and U20037 (N_20037,N_19974,N_19810);
nand U20038 (N_20038,N_19805,N_19863);
xor U20039 (N_20039,N_19975,N_19966);
or U20040 (N_20040,N_19894,N_19834);
nand U20041 (N_20041,N_19867,N_19932);
xor U20042 (N_20042,N_19993,N_19935);
or U20043 (N_20043,N_19969,N_19898);
nor U20044 (N_20044,N_19870,N_19915);
nand U20045 (N_20045,N_19911,N_19948);
nor U20046 (N_20046,N_19930,N_19866);
xnor U20047 (N_20047,N_19964,N_19987);
or U20048 (N_20048,N_19939,N_19960);
nand U20049 (N_20049,N_19919,N_19967);
nor U20050 (N_20050,N_19807,N_19913);
and U20051 (N_20051,N_19854,N_19903);
nand U20052 (N_20052,N_19955,N_19882);
or U20053 (N_20053,N_19906,N_19945);
xnor U20054 (N_20054,N_19949,N_19990);
nor U20055 (N_20055,N_19929,N_19880);
and U20056 (N_20056,N_19812,N_19838);
nor U20057 (N_20057,N_19943,N_19979);
or U20058 (N_20058,N_19833,N_19845);
nand U20059 (N_20059,N_19831,N_19840);
and U20060 (N_20060,N_19871,N_19954);
and U20061 (N_20061,N_19893,N_19873);
nor U20062 (N_20062,N_19907,N_19952);
xor U20063 (N_20063,N_19992,N_19872);
nor U20064 (N_20064,N_19843,N_19978);
nor U20065 (N_20065,N_19991,N_19946);
nand U20066 (N_20066,N_19938,N_19984);
or U20067 (N_20067,N_19957,N_19917);
nand U20068 (N_20068,N_19829,N_19951);
nor U20069 (N_20069,N_19856,N_19956);
nor U20070 (N_20070,N_19816,N_19977);
and U20071 (N_20071,N_19908,N_19899);
or U20072 (N_20072,N_19820,N_19953);
or U20073 (N_20073,N_19983,N_19826);
nor U20074 (N_20074,N_19961,N_19970);
nand U20075 (N_20075,N_19910,N_19865);
and U20076 (N_20076,N_19942,N_19980);
xor U20077 (N_20077,N_19968,N_19862);
nor U20078 (N_20078,N_19934,N_19883);
nor U20079 (N_20079,N_19896,N_19804);
and U20080 (N_20080,N_19971,N_19850);
or U20081 (N_20081,N_19895,N_19868);
nand U20082 (N_20082,N_19959,N_19989);
xnor U20083 (N_20083,N_19941,N_19933);
nand U20084 (N_20084,N_19912,N_19821);
and U20085 (N_20085,N_19877,N_19824);
xor U20086 (N_20086,N_19800,N_19879);
xor U20087 (N_20087,N_19928,N_19965);
nor U20088 (N_20088,N_19921,N_19857);
and U20089 (N_20089,N_19874,N_19985);
nand U20090 (N_20090,N_19920,N_19926);
xor U20091 (N_20091,N_19914,N_19818);
nand U20092 (N_20092,N_19999,N_19849);
and U20093 (N_20093,N_19853,N_19830);
xnor U20094 (N_20094,N_19869,N_19958);
or U20095 (N_20095,N_19803,N_19837);
nor U20096 (N_20096,N_19851,N_19888);
nand U20097 (N_20097,N_19878,N_19981);
xor U20098 (N_20098,N_19842,N_19827);
xor U20099 (N_20099,N_19918,N_19836);
nor U20100 (N_20100,N_19965,N_19918);
nor U20101 (N_20101,N_19944,N_19834);
or U20102 (N_20102,N_19999,N_19837);
or U20103 (N_20103,N_19955,N_19858);
or U20104 (N_20104,N_19998,N_19801);
or U20105 (N_20105,N_19825,N_19930);
nand U20106 (N_20106,N_19961,N_19915);
nand U20107 (N_20107,N_19850,N_19883);
nand U20108 (N_20108,N_19994,N_19855);
xor U20109 (N_20109,N_19954,N_19967);
nand U20110 (N_20110,N_19840,N_19908);
or U20111 (N_20111,N_19891,N_19886);
nand U20112 (N_20112,N_19985,N_19881);
xor U20113 (N_20113,N_19802,N_19845);
and U20114 (N_20114,N_19965,N_19980);
xnor U20115 (N_20115,N_19819,N_19806);
xor U20116 (N_20116,N_19943,N_19969);
and U20117 (N_20117,N_19853,N_19848);
or U20118 (N_20118,N_19887,N_19867);
and U20119 (N_20119,N_19970,N_19893);
and U20120 (N_20120,N_19967,N_19871);
xor U20121 (N_20121,N_19879,N_19969);
xor U20122 (N_20122,N_19973,N_19956);
and U20123 (N_20123,N_19812,N_19805);
nand U20124 (N_20124,N_19895,N_19911);
nand U20125 (N_20125,N_19855,N_19892);
nand U20126 (N_20126,N_19856,N_19877);
and U20127 (N_20127,N_19910,N_19878);
or U20128 (N_20128,N_19948,N_19873);
xnor U20129 (N_20129,N_19996,N_19940);
and U20130 (N_20130,N_19852,N_19914);
and U20131 (N_20131,N_19925,N_19898);
and U20132 (N_20132,N_19985,N_19840);
and U20133 (N_20133,N_19973,N_19853);
nand U20134 (N_20134,N_19858,N_19868);
nand U20135 (N_20135,N_19856,N_19805);
nand U20136 (N_20136,N_19947,N_19959);
and U20137 (N_20137,N_19815,N_19928);
or U20138 (N_20138,N_19820,N_19893);
xnor U20139 (N_20139,N_19902,N_19932);
and U20140 (N_20140,N_19838,N_19859);
nand U20141 (N_20141,N_19966,N_19803);
nand U20142 (N_20142,N_19818,N_19904);
nor U20143 (N_20143,N_19964,N_19836);
or U20144 (N_20144,N_19851,N_19838);
and U20145 (N_20145,N_19946,N_19804);
or U20146 (N_20146,N_19991,N_19951);
nand U20147 (N_20147,N_19964,N_19848);
nor U20148 (N_20148,N_19909,N_19990);
nor U20149 (N_20149,N_19828,N_19984);
nor U20150 (N_20150,N_19879,N_19955);
xor U20151 (N_20151,N_19814,N_19872);
and U20152 (N_20152,N_19803,N_19833);
nand U20153 (N_20153,N_19931,N_19938);
xor U20154 (N_20154,N_19853,N_19842);
and U20155 (N_20155,N_19883,N_19955);
nand U20156 (N_20156,N_19990,N_19824);
nand U20157 (N_20157,N_19985,N_19810);
or U20158 (N_20158,N_19989,N_19832);
xor U20159 (N_20159,N_19971,N_19928);
or U20160 (N_20160,N_19806,N_19816);
and U20161 (N_20161,N_19911,N_19921);
nand U20162 (N_20162,N_19905,N_19840);
xor U20163 (N_20163,N_19948,N_19999);
or U20164 (N_20164,N_19822,N_19892);
nand U20165 (N_20165,N_19854,N_19910);
nand U20166 (N_20166,N_19892,N_19819);
or U20167 (N_20167,N_19988,N_19876);
nand U20168 (N_20168,N_19895,N_19848);
and U20169 (N_20169,N_19876,N_19949);
or U20170 (N_20170,N_19884,N_19868);
or U20171 (N_20171,N_19991,N_19954);
nand U20172 (N_20172,N_19892,N_19881);
nor U20173 (N_20173,N_19895,N_19983);
nand U20174 (N_20174,N_19865,N_19974);
or U20175 (N_20175,N_19941,N_19970);
nand U20176 (N_20176,N_19976,N_19914);
nor U20177 (N_20177,N_19985,N_19804);
and U20178 (N_20178,N_19974,N_19801);
nand U20179 (N_20179,N_19893,N_19824);
nand U20180 (N_20180,N_19818,N_19958);
nor U20181 (N_20181,N_19927,N_19890);
and U20182 (N_20182,N_19945,N_19827);
or U20183 (N_20183,N_19867,N_19996);
nor U20184 (N_20184,N_19878,N_19976);
xnor U20185 (N_20185,N_19828,N_19912);
xnor U20186 (N_20186,N_19932,N_19904);
xnor U20187 (N_20187,N_19857,N_19854);
and U20188 (N_20188,N_19918,N_19806);
nand U20189 (N_20189,N_19843,N_19800);
nand U20190 (N_20190,N_19891,N_19955);
nand U20191 (N_20191,N_19925,N_19957);
xor U20192 (N_20192,N_19840,N_19830);
nand U20193 (N_20193,N_19991,N_19892);
nor U20194 (N_20194,N_19832,N_19869);
and U20195 (N_20195,N_19871,N_19939);
and U20196 (N_20196,N_19888,N_19927);
nand U20197 (N_20197,N_19944,N_19853);
nor U20198 (N_20198,N_19842,N_19850);
and U20199 (N_20199,N_19891,N_19925);
xor U20200 (N_20200,N_20027,N_20093);
xor U20201 (N_20201,N_20085,N_20113);
and U20202 (N_20202,N_20187,N_20028);
xor U20203 (N_20203,N_20007,N_20185);
nand U20204 (N_20204,N_20173,N_20106);
xor U20205 (N_20205,N_20174,N_20096);
xor U20206 (N_20206,N_20108,N_20146);
and U20207 (N_20207,N_20188,N_20039);
or U20208 (N_20208,N_20014,N_20165);
nand U20209 (N_20209,N_20004,N_20018);
xnor U20210 (N_20210,N_20143,N_20012);
or U20211 (N_20211,N_20129,N_20088);
xnor U20212 (N_20212,N_20192,N_20139);
or U20213 (N_20213,N_20194,N_20172);
nor U20214 (N_20214,N_20000,N_20030);
and U20215 (N_20215,N_20057,N_20074);
xnor U20216 (N_20216,N_20116,N_20111);
nand U20217 (N_20217,N_20066,N_20145);
xor U20218 (N_20218,N_20011,N_20024);
and U20219 (N_20219,N_20046,N_20163);
nand U20220 (N_20220,N_20026,N_20043);
nor U20221 (N_20221,N_20151,N_20086);
or U20222 (N_20222,N_20156,N_20084);
or U20223 (N_20223,N_20047,N_20032);
or U20224 (N_20224,N_20054,N_20197);
nor U20225 (N_20225,N_20040,N_20102);
nand U20226 (N_20226,N_20128,N_20193);
and U20227 (N_20227,N_20112,N_20051);
nand U20228 (N_20228,N_20157,N_20005);
and U20229 (N_20229,N_20065,N_20060);
nor U20230 (N_20230,N_20050,N_20137);
or U20231 (N_20231,N_20067,N_20147);
nand U20232 (N_20232,N_20130,N_20037);
nor U20233 (N_20233,N_20160,N_20003);
nand U20234 (N_20234,N_20059,N_20080);
nand U20235 (N_20235,N_20182,N_20158);
nand U20236 (N_20236,N_20083,N_20062);
nand U20237 (N_20237,N_20091,N_20183);
nor U20238 (N_20238,N_20199,N_20117);
nand U20239 (N_20239,N_20115,N_20053);
or U20240 (N_20240,N_20195,N_20041);
nand U20241 (N_20241,N_20019,N_20070);
and U20242 (N_20242,N_20015,N_20022);
nand U20243 (N_20243,N_20101,N_20035);
xnor U20244 (N_20244,N_20056,N_20140);
nand U20245 (N_20245,N_20097,N_20034);
nand U20246 (N_20246,N_20103,N_20119);
xor U20247 (N_20247,N_20114,N_20016);
nand U20248 (N_20248,N_20122,N_20186);
and U20249 (N_20249,N_20073,N_20105);
nor U20250 (N_20250,N_20121,N_20107);
xor U20251 (N_20251,N_20077,N_20082);
and U20252 (N_20252,N_20033,N_20095);
or U20253 (N_20253,N_20132,N_20152);
nor U20254 (N_20254,N_20079,N_20166);
xor U20255 (N_20255,N_20010,N_20150);
and U20256 (N_20256,N_20153,N_20081);
nor U20257 (N_20257,N_20094,N_20090);
and U20258 (N_20258,N_20008,N_20155);
nand U20259 (N_20259,N_20161,N_20148);
and U20260 (N_20260,N_20100,N_20089);
nand U20261 (N_20261,N_20196,N_20049);
xor U20262 (N_20262,N_20029,N_20017);
and U20263 (N_20263,N_20123,N_20178);
xnor U20264 (N_20264,N_20167,N_20052);
xor U20265 (N_20265,N_20009,N_20044);
or U20266 (N_20266,N_20078,N_20075);
xor U20267 (N_20267,N_20098,N_20063);
xnor U20268 (N_20268,N_20164,N_20141);
xnor U20269 (N_20269,N_20092,N_20198);
or U20270 (N_20270,N_20124,N_20135);
xor U20271 (N_20271,N_20175,N_20149);
nor U20272 (N_20272,N_20072,N_20020);
nor U20273 (N_20273,N_20177,N_20013);
and U20274 (N_20274,N_20099,N_20021);
xor U20275 (N_20275,N_20058,N_20179);
xor U20276 (N_20276,N_20064,N_20038);
and U20277 (N_20277,N_20162,N_20159);
nor U20278 (N_20278,N_20069,N_20087);
xor U20279 (N_20279,N_20170,N_20042);
nor U20280 (N_20280,N_20184,N_20071);
nor U20281 (N_20281,N_20104,N_20120);
nand U20282 (N_20282,N_20138,N_20036);
xnor U20283 (N_20283,N_20110,N_20133);
or U20284 (N_20284,N_20181,N_20125);
xnor U20285 (N_20285,N_20025,N_20144);
and U20286 (N_20286,N_20127,N_20176);
nor U20287 (N_20287,N_20031,N_20191);
xnor U20288 (N_20288,N_20134,N_20171);
and U20289 (N_20289,N_20118,N_20190);
nor U20290 (N_20290,N_20169,N_20109);
or U20291 (N_20291,N_20154,N_20168);
and U20292 (N_20292,N_20189,N_20180);
and U20293 (N_20293,N_20048,N_20023);
or U20294 (N_20294,N_20142,N_20068);
nand U20295 (N_20295,N_20076,N_20006);
xnor U20296 (N_20296,N_20061,N_20136);
nand U20297 (N_20297,N_20001,N_20055);
nor U20298 (N_20298,N_20045,N_20126);
or U20299 (N_20299,N_20131,N_20002);
xor U20300 (N_20300,N_20082,N_20014);
xnor U20301 (N_20301,N_20184,N_20116);
xor U20302 (N_20302,N_20128,N_20040);
nand U20303 (N_20303,N_20086,N_20159);
nand U20304 (N_20304,N_20014,N_20068);
and U20305 (N_20305,N_20030,N_20115);
nand U20306 (N_20306,N_20003,N_20185);
or U20307 (N_20307,N_20022,N_20160);
and U20308 (N_20308,N_20009,N_20004);
xnor U20309 (N_20309,N_20060,N_20111);
nand U20310 (N_20310,N_20115,N_20098);
xnor U20311 (N_20311,N_20030,N_20001);
and U20312 (N_20312,N_20017,N_20044);
or U20313 (N_20313,N_20142,N_20037);
xnor U20314 (N_20314,N_20002,N_20095);
nand U20315 (N_20315,N_20047,N_20056);
nor U20316 (N_20316,N_20121,N_20130);
or U20317 (N_20317,N_20043,N_20024);
or U20318 (N_20318,N_20083,N_20180);
xor U20319 (N_20319,N_20153,N_20056);
nor U20320 (N_20320,N_20169,N_20057);
nor U20321 (N_20321,N_20102,N_20005);
nor U20322 (N_20322,N_20183,N_20194);
or U20323 (N_20323,N_20133,N_20033);
nand U20324 (N_20324,N_20147,N_20045);
nor U20325 (N_20325,N_20057,N_20141);
nor U20326 (N_20326,N_20137,N_20153);
xor U20327 (N_20327,N_20092,N_20077);
xnor U20328 (N_20328,N_20011,N_20088);
xor U20329 (N_20329,N_20092,N_20171);
nand U20330 (N_20330,N_20124,N_20034);
xnor U20331 (N_20331,N_20191,N_20128);
nand U20332 (N_20332,N_20180,N_20153);
nor U20333 (N_20333,N_20063,N_20005);
or U20334 (N_20334,N_20059,N_20155);
nor U20335 (N_20335,N_20121,N_20015);
nand U20336 (N_20336,N_20092,N_20101);
nor U20337 (N_20337,N_20039,N_20003);
nor U20338 (N_20338,N_20026,N_20184);
and U20339 (N_20339,N_20091,N_20119);
nand U20340 (N_20340,N_20081,N_20043);
nand U20341 (N_20341,N_20168,N_20084);
nand U20342 (N_20342,N_20024,N_20041);
nor U20343 (N_20343,N_20078,N_20048);
nor U20344 (N_20344,N_20195,N_20070);
nand U20345 (N_20345,N_20165,N_20136);
nor U20346 (N_20346,N_20054,N_20048);
or U20347 (N_20347,N_20084,N_20105);
or U20348 (N_20348,N_20065,N_20091);
nor U20349 (N_20349,N_20123,N_20152);
or U20350 (N_20350,N_20176,N_20111);
nand U20351 (N_20351,N_20111,N_20047);
nor U20352 (N_20352,N_20092,N_20074);
xnor U20353 (N_20353,N_20067,N_20092);
and U20354 (N_20354,N_20182,N_20010);
nor U20355 (N_20355,N_20173,N_20067);
nand U20356 (N_20356,N_20136,N_20187);
nor U20357 (N_20357,N_20000,N_20011);
xnor U20358 (N_20358,N_20090,N_20038);
nor U20359 (N_20359,N_20173,N_20076);
nand U20360 (N_20360,N_20031,N_20047);
or U20361 (N_20361,N_20126,N_20147);
xnor U20362 (N_20362,N_20161,N_20129);
xor U20363 (N_20363,N_20049,N_20122);
and U20364 (N_20364,N_20186,N_20133);
nor U20365 (N_20365,N_20030,N_20034);
nor U20366 (N_20366,N_20037,N_20107);
xor U20367 (N_20367,N_20198,N_20105);
nor U20368 (N_20368,N_20094,N_20053);
nor U20369 (N_20369,N_20035,N_20111);
nand U20370 (N_20370,N_20082,N_20013);
and U20371 (N_20371,N_20163,N_20007);
and U20372 (N_20372,N_20156,N_20007);
or U20373 (N_20373,N_20142,N_20130);
nand U20374 (N_20374,N_20078,N_20015);
xnor U20375 (N_20375,N_20118,N_20016);
xnor U20376 (N_20376,N_20131,N_20140);
or U20377 (N_20377,N_20040,N_20046);
nor U20378 (N_20378,N_20186,N_20028);
and U20379 (N_20379,N_20033,N_20193);
or U20380 (N_20380,N_20079,N_20099);
nand U20381 (N_20381,N_20193,N_20159);
nor U20382 (N_20382,N_20109,N_20082);
nand U20383 (N_20383,N_20161,N_20133);
and U20384 (N_20384,N_20198,N_20038);
or U20385 (N_20385,N_20175,N_20001);
or U20386 (N_20386,N_20118,N_20113);
or U20387 (N_20387,N_20120,N_20128);
or U20388 (N_20388,N_20179,N_20193);
or U20389 (N_20389,N_20198,N_20123);
nor U20390 (N_20390,N_20196,N_20022);
and U20391 (N_20391,N_20041,N_20180);
and U20392 (N_20392,N_20166,N_20043);
and U20393 (N_20393,N_20004,N_20190);
and U20394 (N_20394,N_20048,N_20173);
and U20395 (N_20395,N_20180,N_20057);
nand U20396 (N_20396,N_20095,N_20091);
and U20397 (N_20397,N_20067,N_20195);
nor U20398 (N_20398,N_20009,N_20096);
nand U20399 (N_20399,N_20092,N_20119);
nor U20400 (N_20400,N_20241,N_20348);
and U20401 (N_20401,N_20253,N_20215);
and U20402 (N_20402,N_20293,N_20302);
xnor U20403 (N_20403,N_20266,N_20347);
nand U20404 (N_20404,N_20396,N_20259);
nand U20405 (N_20405,N_20272,N_20342);
and U20406 (N_20406,N_20256,N_20352);
nand U20407 (N_20407,N_20242,N_20225);
nor U20408 (N_20408,N_20207,N_20235);
nand U20409 (N_20409,N_20267,N_20280);
nor U20410 (N_20410,N_20249,N_20287);
nand U20411 (N_20411,N_20254,N_20209);
nand U20412 (N_20412,N_20260,N_20344);
nand U20413 (N_20413,N_20323,N_20319);
xor U20414 (N_20414,N_20214,N_20245);
xnor U20415 (N_20415,N_20271,N_20376);
xor U20416 (N_20416,N_20247,N_20273);
nand U20417 (N_20417,N_20246,N_20202);
nand U20418 (N_20418,N_20313,N_20368);
or U20419 (N_20419,N_20336,N_20284);
nand U20420 (N_20420,N_20372,N_20219);
xnor U20421 (N_20421,N_20311,N_20375);
xor U20422 (N_20422,N_20262,N_20232);
and U20423 (N_20423,N_20335,N_20310);
and U20424 (N_20424,N_20222,N_20330);
nand U20425 (N_20425,N_20286,N_20334);
and U20426 (N_20426,N_20393,N_20371);
xnor U20427 (N_20427,N_20263,N_20357);
xnor U20428 (N_20428,N_20381,N_20298);
nor U20429 (N_20429,N_20331,N_20353);
nand U20430 (N_20430,N_20360,N_20261);
nor U20431 (N_20431,N_20324,N_20201);
or U20432 (N_20432,N_20355,N_20339);
nand U20433 (N_20433,N_20274,N_20210);
or U20434 (N_20434,N_20237,N_20304);
nand U20435 (N_20435,N_20397,N_20359);
and U20436 (N_20436,N_20248,N_20350);
or U20437 (N_20437,N_20268,N_20392);
nor U20438 (N_20438,N_20373,N_20328);
nand U20439 (N_20439,N_20299,N_20307);
xnor U20440 (N_20440,N_20233,N_20205);
and U20441 (N_20441,N_20289,N_20203);
or U20442 (N_20442,N_20270,N_20231);
xor U20443 (N_20443,N_20291,N_20206);
or U20444 (N_20444,N_20282,N_20356);
xor U20445 (N_20445,N_20258,N_20227);
nand U20446 (N_20446,N_20275,N_20220);
xor U20447 (N_20447,N_20309,N_20301);
and U20448 (N_20448,N_20251,N_20312);
nor U20449 (N_20449,N_20322,N_20243);
nand U20450 (N_20450,N_20252,N_20305);
or U20451 (N_20451,N_20361,N_20306);
nor U20452 (N_20452,N_20370,N_20308);
nand U20453 (N_20453,N_20395,N_20386);
and U20454 (N_20454,N_20234,N_20379);
and U20455 (N_20455,N_20390,N_20238);
nor U20456 (N_20456,N_20388,N_20223);
xnor U20457 (N_20457,N_20389,N_20367);
nor U20458 (N_20458,N_20387,N_20358);
or U20459 (N_20459,N_20281,N_20314);
or U20460 (N_20460,N_20224,N_20277);
xnor U20461 (N_20461,N_20211,N_20349);
and U20462 (N_20462,N_20333,N_20226);
xor U20463 (N_20463,N_20384,N_20217);
nand U20464 (N_20464,N_20303,N_20327);
xnor U20465 (N_20465,N_20383,N_20200);
and U20466 (N_20466,N_20332,N_20338);
and U20467 (N_20467,N_20369,N_20212);
xnor U20468 (N_20468,N_20340,N_20264);
nand U20469 (N_20469,N_20318,N_20297);
nand U20470 (N_20470,N_20363,N_20399);
xor U20471 (N_20471,N_20391,N_20276);
nand U20472 (N_20472,N_20257,N_20204);
or U20473 (N_20473,N_20278,N_20230);
xnor U20474 (N_20474,N_20343,N_20398);
or U20475 (N_20475,N_20240,N_20296);
xnor U20476 (N_20476,N_20351,N_20283);
and U20477 (N_20477,N_20315,N_20326);
xnor U20478 (N_20478,N_20385,N_20229);
nand U20479 (N_20479,N_20354,N_20269);
xnor U20480 (N_20480,N_20294,N_20364);
and U20481 (N_20481,N_20341,N_20228);
nand U20482 (N_20482,N_20279,N_20295);
nand U20483 (N_20483,N_20329,N_20320);
or U20484 (N_20484,N_20244,N_20365);
and U20485 (N_20485,N_20346,N_20325);
or U20486 (N_20486,N_20250,N_20377);
and U20487 (N_20487,N_20362,N_20317);
nor U20488 (N_20488,N_20265,N_20321);
xnor U20489 (N_20489,N_20218,N_20213);
or U20490 (N_20490,N_20316,N_20366);
nor U20491 (N_20491,N_20236,N_20382);
nand U20492 (N_20492,N_20292,N_20239);
or U20493 (N_20493,N_20290,N_20255);
nor U20494 (N_20494,N_20380,N_20374);
and U20495 (N_20495,N_20208,N_20337);
nand U20496 (N_20496,N_20394,N_20378);
or U20497 (N_20497,N_20216,N_20300);
xor U20498 (N_20498,N_20285,N_20288);
nand U20499 (N_20499,N_20345,N_20221);
and U20500 (N_20500,N_20315,N_20289);
or U20501 (N_20501,N_20390,N_20307);
nor U20502 (N_20502,N_20267,N_20255);
nor U20503 (N_20503,N_20227,N_20231);
and U20504 (N_20504,N_20314,N_20349);
nor U20505 (N_20505,N_20380,N_20334);
xnor U20506 (N_20506,N_20347,N_20225);
and U20507 (N_20507,N_20373,N_20298);
or U20508 (N_20508,N_20369,N_20239);
nor U20509 (N_20509,N_20264,N_20358);
xor U20510 (N_20510,N_20283,N_20353);
nand U20511 (N_20511,N_20349,N_20346);
nor U20512 (N_20512,N_20378,N_20239);
or U20513 (N_20513,N_20389,N_20293);
nor U20514 (N_20514,N_20377,N_20205);
nand U20515 (N_20515,N_20207,N_20245);
and U20516 (N_20516,N_20388,N_20236);
xor U20517 (N_20517,N_20318,N_20398);
nand U20518 (N_20518,N_20364,N_20261);
xor U20519 (N_20519,N_20213,N_20369);
or U20520 (N_20520,N_20274,N_20306);
and U20521 (N_20521,N_20329,N_20243);
or U20522 (N_20522,N_20300,N_20246);
xor U20523 (N_20523,N_20296,N_20290);
or U20524 (N_20524,N_20284,N_20303);
or U20525 (N_20525,N_20339,N_20236);
xnor U20526 (N_20526,N_20239,N_20350);
nor U20527 (N_20527,N_20233,N_20281);
xor U20528 (N_20528,N_20280,N_20294);
and U20529 (N_20529,N_20278,N_20284);
and U20530 (N_20530,N_20215,N_20226);
xor U20531 (N_20531,N_20272,N_20341);
and U20532 (N_20532,N_20386,N_20334);
or U20533 (N_20533,N_20337,N_20349);
or U20534 (N_20534,N_20203,N_20246);
nor U20535 (N_20535,N_20301,N_20294);
nand U20536 (N_20536,N_20387,N_20231);
nand U20537 (N_20537,N_20265,N_20304);
xor U20538 (N_20538,N_20375,N_20240);
or U20539 (N_20539,N_20398,N_20394);
nand U20540 (N_20540,N_20320,N_20394);
xor U20541 (N_20541,N_20394,N_20344);
nor U20542 (N_20542,N_20281,N_20224);
or U20543 (N_20543,N_20322,N_20309);
nor U20544 (N_20544,N_20253,N_20388);
nand U20545 (N_20545,N_20259,N_20291);
nor U20546 (N_20546,N_20297,N_20329);
and U20547 (N_20547,N_20346,N_20311);
or U20548 (N_20548,N_20206,N_20226);
xor U20549 (N_20549,N_20233,N_20390);
and U20550 (N_20550,N_20287,N_20261);
and U20551 (N_20551,N_20304,N_20339);
and U20552 (N_20552,N_20321,N_20287);
and U20553 (N_20553,N_20246,N_20354);
xnor U20554 (N_20554,N_20260,N_20395);
nor U20555 (N_20555,N_20333,N_20327);
xnor U20556 (N_20556,N_20218,N_20311);
xor U20557 (N_20557,N_20392,N_20337);
nand U20558 (N_20558,N_20339,N_20263);
or U20559 (N_20559,N_20341,N_20370);
or U20560 (N_20560,N_20279,N_20243);
nor U20561 (N_20561,N_20270,N_20235);
nand U20562 (N_20562,N_20311,N_20255);
xor U20563 (N_20563,N_20207,N_20396);
nand U20564 (N_20564,N_20322,N_20374);
or U20565 (N_20565,N_20296,N_20279);
xnor U20566 (N_20566,N_20261,N_20398);
or U20567 (N_20567,N_20334,N_20307);
or U20568 (N_20568,N_20338,N_20399);
nor U20569 (N_20569,N_20305,N_20360);
nand U20570 (N_20570,N_20397,N_20285);
or U20571 (N_20571,N_20261,N_20208);
and U20572 (N_20572,N_20384,N_20245);
nor U20573 (N_20573,N_20335,N_20246);
nor U20574 (N_20574,N_20283,N_20204);
xnor U20575 (N_20575,N_20303,N_20357);
and U20576 (N_20576,N_20294,N_20354);
and U20577 (N_20577,N_20206,N_20371);
or U20578 (N_20578,N_20304,N_20358);
xnor U20579 (N_20579,N_20213,N_20240);
nand U20580 (N_20580,N_20302,N_20227);
nand U20581 (N_20581,N_20377,N_20376);
nor U20582 (N_20582,N_20302,N_20226);
xnor U20583 (N_20583,N_20254,N_20369);
nand U20584 (N_20584,N_20250,N_20274);
nand U20585 (N_20585,N_20359,N_20313);
nor U20586 (N_20586,N_20202,N_20319);
nand U20587 (N_20587,N_20224,N_20324);
and U20588 (N_20588,N_20324,N_20281);
nand U20589 (N_20589,N_20270,N_20287);
nor U20590 (N_20590,N_20215,N_20390);
and U20591 (N_20591,N_20317,N_20336);
nand U20592 (N_20592,N_20296,N_20242);
xnor U20593 (N_20593,N_20249,N_20256);
or U20594 (N_20594,N_20284,N_20222);
nor U20595 (N_20595,N_20340,N_20220);
and U20596 (N_20596,N_20322,N_20202);
and U20597 (N_20597,N_20371,N_20239);
nand U20598 (N_20598,N_20321,N_20372);
nor U20599 (N_20599,N_20283,N_20361);
nor U20600 (N_20600,N_20428,N_20491);
nor U20601 (N_20601,N_20499,N_20543);
and U20602 (N_20602,N_20571,N_20475);
or U20603 (N_20603,N_20411,N_20546);
xnor U20604 (N_20604,N_20541,N_20525);
and U20605 (N_20605,N_20501,N_20568);
and U20606 (N_20606,N_20412,N_20540);
or U20607 (N_20607,N_20415,N_20544);
or U20608 (N_20608,N_20576,N_20417);
nor U20609 (N_20609,N_20514,N_20515);
and U20610 (N_20610,N_20523,N_20551);
xnor U20611 (N_20611,N_20587,N_20457);
or U20612 (N_20612,N_20574,N_20472);
or U20613 (N_20613,N_20529,N_20463);
xor U20614 (N_20614,N_20488,N_20410);
and U20615 (N_20615,N_20512,N_20466);
nand U20616 (N_20616,N_20583,N_20596);
and U20617 (N_20617,N_20430,N_20450);
xnor U20618 (N_20618,N_20593,N_20500);
and U20619 (N_20619,N_20555,N_20504);
xor U20620 (N_20620,N_20449,N_20545);
nand U20621 (N_20621,N_20460,N_20401);
or U20622 (N_20622,N_20444,N_20482);
xor U20623 (N_20623,N_20425,N_20526);
nand U20624 (N_20624,N_20517,N_20524);
and U20625 (N_20625,N_20521,N_20573);
nor U20626 (N_20626,N_20542,N_20554);
and U20627 (N_20627,N_20427,N_20508);
nor U20628 (N_20628,N_20575,N_20424);
or U20629 (N_20629,N_20563,N_20516);
nor U20630 (N_20630,N_20589,N_20539);
xor U20631 (N_20631,N_20564,N_20433);
nor U20632 (N_20632,N_20513,N_20431);
nand U20633 (N_20633,N_20465,N_20458);
or U20634 (N_20634,N_20439,N_20558);
nand U20635 (N_20635,N_20537,N_20552);
nand U20636 (N_20636,N_20532,N_20440);
xor U20637 (N_20637,N_20414,N_20476);
and U20638 (N_20638,N_20469,N_20549);
nand U20639 (N_20639,N_20435,N_20464);
nor U20640 (N_20640,N_20467,N_20538);
xnor U20641 (N_20641,N_20556,N_20487);
and U20642 (N_20642,N_20586,N_20506);
and U20643 (N_20643,N_20403,N_20502);
or U20644 (N_20644,N_20400,N_20420);
or U20645 (N_20645,N_20599,N_20520);
xor U20646 (N_20646,N_20530,N_20489);
nor U20647 (N_20647,N_20598,N_20509);
nand U20648 (N_20648,N_20561,N_20584);
xnor U20649 (N_20649,N_20479,N_20461);
nand U20650 (N_20650,N_20594,N_20591);
nand U20651 (N_20651,N_20592,N_20579);
nand U20652 (N_20652,N_20547,N_20493);
xor U20653 (N_20653,N_20503,N_20477);
xnor U20654 (N_20654,N_20455,N_20498);
or U20655 (N_20655,N_20405,N_20562);
nand U20656 (N_20656,N_20505,N_20447);
and U20657 (N_20657,N_20557,N_20580);
xor U20658 (N_20658,N_20566,N_20408);
nor U20659 (N_20659,N_20585,N_20409);
nor U20660 (N_20660,N_20507,N_20456);
xor U20661 (N_20661,N_20485,N_20470);
or U20662 (N_20662,N_20553,N_20535);
or U20663 (N_20663,N_20445,N_20490);
nand U20664 (N_20664,N_20581,N_20478);
nand U20665 (N_20665,N_20416,N_20550);
nor U20666 (N_20666,N_20423,N_20441);
nor U20667 (N_20667,N_20448,N_20459);
xnor U20668 (N_20668,N_20406,N_20595);
nor U20669 (N_20669,N_20510,N_20436);
nand U20670 (N_20670,N_20492,N_20531);
or U20671 (N_20671,N_20486,N_20453);
or U20672 (N_20672,N_20597,N_20511);
and U20673 (N_20673,N_20468,N_20588);
and U20674 (N_20674,N_20590,N_20548);
nor U20675 (N_20675,N_20527,N_20481);
nand U20676 (N_20676,N_20522,N_20421);
xnor U20677 (N_20677,N_20434,N_20572);
nor U20678 (N_20678,N_20438,N_20569);
xnor U20679 (N_20679,N_20426,N_20446);
nor U20680 (N_20680,N_20565,N_20437);
or U20681 (N_20681,N_20443,N_20533);
or U20682 (N_20682,N_20484,N_20474);
nor U20683 (N_20683,N_20432,N_20418);
or U20684 (N_20684,N_20494,N_20496);
xor U20685 (N_20685,N_20536,N_20407);
nor U20686 (N_20686,N_20567,N_20559);
and U20687 (N_20687,N_20402,N_20519);
or U20688 (N_20688,N_20413,N_20429);
nand U20689 (N_20689,N_20497,N_20462);
nand U20690 (N_20690,N_20473,N_20451);
or U20691 (N_20691,N_20404,N_20471);
nor U20692 (N_20692,N_20560,N_20480);
and U20693 (N_20693,N_20528,N_20518);
nor U20694 (N_20694,N_20422,N_20419);
nand U20695 (N_20695,N_20582,N_20534);
xnor U20696 (N_20696,N_20452,N_20442);
nand U20697 (N_20697,N_20454,N_20577);
xnor U20698 (N_20698,N_20483,N_20495);
nor U20699 (N_20699,N_20578,N_20570);
or U20700 (N_20700,N_20440,N_20579);
and U20701 (N_20701,N_20571,N_20483);
or U20702 (N_20702,N_20549,N_20587);
or U20703 (N_20703,N_20420,N_20443);
xnor U20704 (N_20704,N_20555,N_20547);
and U20705 (N_20705,N_20483,N_20579);
nand U20706 (N_20706,N_20483,N_20400);
nand U20707 (N_20707,N_20552,N_20490);
nand U20708 (N_20708,N_20414,N_20568);
xnor U20709 (N_20709,N_20488,N_20481);
nor U20710 (N_20710,N_20559,N_20581);
xor U20711 (N_20711,N_20565,N_20459);
nand U20712 (N_20712,N_20461,N_20553);
and U20713 (N_20713,N_20480,N_20532);
nor U20714 (N_20714,N_20410,N_20455);
nand U20715 (N_20715,N_20424,N_20551);
nand U20716 (N_20716,N_20580,N_20587);
and U20717 (N_20717,N_20534,N_20476);
or U20718 (N_20718,N_20400,N_20458);
and U20719 (N_20719,N_20479,N_20536);
nand U20720 (N_20720,N_20464,N_20584);
nor U20721 (N_20721,N_20529,N_20503);
nand U20722 (N_20722,N_20568,N_20563);
nand U20723 (N_20723,N_20493,N_20511);
xor U20724 (N_20724,N_20495,N_20503);
nand U20725 (N_20725,N_20497,N_20460);
xnor U20726 (N_20726,N_20510,N_20573);
nand U20727 (N_20727,N_20446,N_20449);
or U20728 (N_20728,N_20520,N_20466);
nor U20729 (N_20729,N_20591,N_20472);
or U20730 (N_20730,N_20548,N_20535);
or U20731 (N_20731,N_20504,N_20523);
nor U20732 (N_20732,N_20442,N_20415);
nor U20733 (N_20733,N_20597,N_20426);
nor U20734 (N_20734,N_20419,N_20553);
xor U20735 (N_20735,N_20404,N_20528);
or U20736 (N_20736,N_20429,N_20494);
and U20737 (N_20737,N_20525,N_20446);
nand U20738 (N_20738,N_20466,N_20498);
nand U20739 (N_20739,N_20422,N_20464);
or U20740 (N_20740,N_20561,N_20585);
or U20741 (N_20741,N_20598,N_20421);
nor U20742 (N_20742,N_20563,N_20508);
nor U20743 (N_20743,N_20573,N_20508);
nor U20744 (N_20744,N_20440,N_20500);
xor U20745 (N_20745,N_20546,N_20558);
or U20746 (N_20746,N_20499,N_20599);
nor U20747 (N_20747,N_20507,N_20524);
nand U20748 (N_20748,N_20594,N_20457);
nand U20749 (N_20749,N_20547,N_20436);
or U20750 (N_20750,N_20512,N_20449);
and U20751 (N_20751,N_20444,N_20450);
xor U20752 (N_20752,N_20587,N_20551);
nor U20753 (N_20753,N_20410,N_20465);
nand U20754 (N_20754,N_20436,N_20558);
xnor U20755 (N_20755,N_20516,N_20411);
nor U20756 (N_20756,N_20404,N_20507);
nor U20757 (N_20757,N_20468,N_20509);
nor U20758 (N_20758,N_20505,N_20546);
nand U20759 (N_20759,N_20444,N_20543);
or U20760 (N_20760,N_20574,N_20439);
xor U20761 (N_20761,N_20494,N_20591);
or U20762 (N_20762,N_20529,N_20431);
and U20763 (N_20763,N_20582,N_20486);
nor U20764 (N_20764,N_20405,N_20517);
nand U20765 (N_20765,N_20549,N_20523);
xnor U20766 (N_20766,N_20577,N_20487);
nand U20767 (N_20767,N_20539,N_20529);
xor U20768 (N_20768,N_20475,N_20458);
xor U20769 (N_20769,N_20472,N_20558);
xor U20770 (N_20770,N_20425,N_20411);
or U20771 (N_20771,N_20513,N_20521);
nand U20772 (N_20772,N_20419,N_20540);
or U20773 (N_20773,N_20457,N_20515);
and U20774 (N_20774,N_20527,N_20407);
and U20775 (N_20775,N_20487,N_20483);
or U20776 (N_20776,N_20447,N_20523);
nand U20777 (N_20777,N_20472,N_20594);
xnor U20778 (N_20778,N_20531,N_20529);
nor U20779 (N_20779,N_20419,N_20520);
and U20780 (N_20780,N_20401,N_20524);
xor U20781 (N_20781,N_20529,N_20497);
or U20782 (N_20782,N_20475,N_20478);
or U20783 (N_20783,N_20453,N_20543);
or U20784 (N_20784,N_20557,N_20401);
xor U20785 (N_20785,N_20463,N_20485);
and U20786 (N_20786,N_20520,N_20534);
nor U20787 (N_20787,N_20487,N_20492);
xor U20788 (N_20788,N_20421,N_20478);
nor U20789 (N_20789,N_20499,N_20587);
xor U20790 (N_20790,N_20432,N_20578);
nor U20791 (N_20791,N_20576,N_20589);
nor U20792 (N_20792,N_20432,N_20589);
xnor U20793 (N_20793,N_20567,N_20475);
xnor U20794 (N_20794,N_20515,N_20464);
or U20795 (N_20795,N_20467,N_20419);
xor U20796 (N_20796,N_20458,N_20505);
and U20797 (N_20797,N_20527,N_20543);
xor U20798 (N_20798,N_20582,N_20405);
nand U20799 (N_20799,N_20428,N_20516);
xnor U20800 (N_20800,N_20705,N_20666);
or U20801 (N_20801,N_20786,N_20613);
nor U20802 (N_20802,N_20731,N_20650);
xor U20803 (N_20803,N_20732,N_20778);
nand U20804 (N_20804,N_20695,N_20750);
and U20805 (N_20805,N_20684,N_20764);
xor U20806 (N_20806,N_20604,N_20672);
nor U20807 (N_20807,N_20641,N_20626);
xnor U20808 (N_20808,N_20678,N_20692);
xnor U20809 (N_20809,N_20729,N_20708);
xor U20810 (N_20810,N_20675,N_20785);
xor U20811 (N_20811,N_20796,N_20671);
nand U20812 (N_20812,N_20746,N_20691);
and U20813 (N_20813,N_20709,N_20611);
nor U20814 (N_20814,N_20605,N_20667);
nand U20815 (N_20815,N_20752,N_20735);
xnor U20816 (N_20816,N_20733,N_20624);
nor U20817 (N_20817,N_20619,N_20730);
xnor U20818 (N_20818,N_20794,N_20724);
nor U20819 (N_20819,N_20797,N_20700);
and U20820 (N_20820,N_20656,N_20767);
xnor U20821 (N_20821,N_20620,N_20647);
xor U20822 (N_20822,N_20789,N_20637);
and U20823 (N_20823,N_20645,N_20682);
nor U20824 (N_20824,N_20761,N_20640);
and U20825 (N_20825,N_20759,N_20721);
nor U20826 (N_20826,N_20725,N_20639);
xnor U20827 (N_20827,N_20670,N_20755);
xor U20828 (N_20828,N_20630,N_20792);
nand U20829 (N_20829,N_20701,N_20710);
and U20830 (N_20830,N_20696,N_20616);
xnor U20831 (N_20831,N_20689,N_20726);
or U20832 (N_20832,N_20791,N_20737);
and U20833 (N_20833,N_20783,N_20775);
or U20834 (N_20834,N_20683,N_20743);
or U20835 (N_20835,N_20679,N_20782);
nor U20836 (N_20836,N_20722,N_20627);
nor U20837 (N_20837,N_20623,N_20749);
nor U20838 (N_20838,N_20606,N_20713);
xor U20839 (N_20839,N_20658,N_20720);
and U20840 (N_20840,N_20669,N_20612);
and U20841 (N_20841,N_20603,N_20772);
nor U20842 (N_20842,N_20742,N_20712);
or U20843 (N_20843,N_20771,N_20768);
and U20844 (N_20844,N_20662,N_20781);
nand U20845 (N_20845,N_20677,N_20763);
nand U20846 (N_20846,N_20688,N_20681);
or U20847 (N_20847,N_20719,N_20685);
and U20848 (N_20848,N_20625,N_20715);
nor U20849 (N_20849,N_20655,N_20757);
xnor U20850 (N_20850,N_20601,N_20795);
xnor U20851 (N_20851,N_20673,N_20762);
xor U20852 (N_20852,N_20697,N_20774);
or U20853 (N_20853,N_20635,N_20674);
xor U20854 (N_20854,N_20646,N_20615);
nand U20855 (N_20855,N_20621,N_20659);
and U20856 (N_20856,N_20738,N_20788);
nand U20857 (N_20857,N_20717,N_20664);
nand U20858 (N_20858,N_20660,N_20642);
or U20859 (N_20859,N_20756,N_20634);
and U20860 (N_20860,N_20663,N_20610);
or U20861 (N_20861,N_20607,N_20628);
nor U20862 (N_20862,N_20614,N_20693);
nor U20863 (N_20863,N_20734,N_20633);
xor U20864 (N_20864,N_20636,N_20736);
xor U20865 (N_20865,N_20758,N_20779);
xor U20866 (N_20866,N_20790,N_20770);
nor U20867 (N_20867,N_20609,N_20754);
xnor U20868 (N_20868,N_20744,N_20657);
or U20869 (N_20869,N_20643,N_20784);
and U20870 (N_20870,N_20780,N_20769);
xor U20871 (N_20871,N_20787,N_20748);
nand U20872 (N_20872,N_20653,N_20649);
nand U20873 (N_20873,N_20723,N_20694);
and U20874 (N_20874,N_20728,N_20706);
xnor U20875 (N_20875,N_20698,N_20798);
nand U20876 (N_20876,N_20766,N_20680);
and U20877 (N_20877,N_20648,N_20714);
nor U20878 (N_20878,N_20765,N_20711);
and U20879 (N_20879,N_20751,N_20707);
xor U20880 (N_20880,N_20652,N_20661);
xor U20881 (N_20881,N_20686,N_20760);
nand U20882 (N_20882,N_20777,N_20676);
and U20883 (N_20883,N_20716,N_20665);
or U20884 (N_20884,N_20608,N_20718);
xor U20885 (N_20885,N_20741,N_20687);
xor U20886 (N_20886,N_20753,N_20617);
xor U20887 (N_20887,N_20702,N_20773);
xnor U20888 (N_20888,N_20651,N_20747);
nor U20889 (N_20889,N_20776,N_20727);
or U20890 (N_20890,N_20602,N_20632);
nor U20891 (N_20891,N_20799,N_20740);
nor U20892 (N_20892,N_20600,N_20793);
nor U20893 (N_20893,N_20644,N_20618);
or U20894 (N_20894,N_20703,N_20638);
nor U20895 (N_20895,N_20622,N_20690);
xnor U20896 (N_20896,N_20745,N_20654);
xor U20897 (N_20897,N_20631,N_20704);
and U20898 (N_20898,N_20739,N_20668);
or U20899 (N_20899,N_20629,N_20699);
xnor U20900 (N_20900,N_20790,N_20684);
nor U20901 (N_20901,N_20622,N_20730);
nand U20902 (N_20902,N_20752,N_20634);
or U20903 (N_20903,N_20675,N_20703);
and U20904 (N_20904,N_20672,N_20612);
nor U20905 (N_20905,N_20759,N_20765);
xor U20906 (N_20906,N_20746,N_20677);
nand U20907 (N_20907,N_20777,N_20607);
xnor U20908 (N_20908,N_20736,N_20758);
nor U20909 (N_20909,N_20666,N_20748);
or U20910 (N_20910,N_20615,N_20693);
nor U20911 (N_20911,N_20665,N_20770);
nand U20912 (N_20912,N_20652,N_20746);
nor U20913 (N_20913,N_20777,N_20707);
nand U20914 (N_20914,N_20726,N_20749);
or U20915 (N_20915,N_20735,N_20685);
or U20916 (N_20916,N_20642,N_20619);
xor U20917 (N_20917,N_20760,N_20630);
or U20918 (N_20918,N_20725,N_20606);
nand U20919 (N_20919,N_20664,N_20683);
or U20920 (N_20920,N_20783,N_20689);
nand U20921 (N_20921,N_20751,N_20758);
or U20922 (N_20922,N_20620,N_20744);
xor U20923 (N_20923,N_20654,N_20731);
xor U20924 (N_20924,N_20628,N_20692);
nand U20925 (N_20925,N_20730,N_20663);
or U20926 (N_20926,N_20700,N_20641);
nand U20927 (N_20927,N_20609,N_20696);
xnor U20928 (N_20928,N_20752,N_20766);
xnor U20929 (N_20929,N_20692,N_20657);
nand U20930 (N_20930,N_20640,N_20789);
and U20931 (N_20931,N_20654,N_20625);
nand U20932 (N_20932,N_20627,N_20774);
xnor U20933 (N_20933,N_20675,N_20782);
xor U20934 (N_20934,N_20732,N_20622);
and U20935 (N_20935,N_20649,N_20757);
or U20936 (N_20936,N_20755,N_20619);
and U20937 (N_20937,N_20754,N_20730);
or U20938 (N_20938,N_20725,N_20636);
nand U20939 (N_20939,N_20774,N_20764);
nor U20940 (N_20940,N_20627,N_20688);
or U20941 (N_20941,N_20609,N_20660);
nor U20942 (N_20942,N_20705,N_20699);
xnor U20943 (N_20943,N_20729,N_20746);
or U20944 (N_20944,N_20740,N_20758);
nand U20945 (N_20945,N_20671,N_20731);
nand U20946 (N_20946,N_20752,N_20739);
and U20947 (N_20947,N_20754,N_20729);
and U20948 (N_20948,N_20638,N_20734);
nor U20949 (N_20949,N_20752,N_20603);
xnor U20950 (N_20950,N_20621,N_20701);
or U20951 (N_20951,N_20758,N_20793);
xor U20952 (N_20952,N_20773,N_20616);
nor U20953 (N_20953,N_20796,N_20743);
nor U20954 (N_20954,N_20642,N_20615);
or U20955 (N_20955,N_20629,N_20622);
or U20956 (N_20956,N_20704,N_20638);
xor U20957 (N_20957,N_20661,N_20771);
nor U20958 (N_20958,N_20707,N_20621);
nor U20959 (N_20959,N_20642,N_20694);
nand U20960 (N_20960,N_20722,N_20787);
nand U20961 (N_20961,N_20770,N_20742);
xnor U20962 (N_20962,N_20785,N_20623);
and U20963 (N_20963,N_20724,N_20676);
nand U20964 (N_20964,N_20707,N_20781);
or U20965 (N_20965,N_20717,N_20686);
nand U20966 (N_20966,N_20772,N_20766);
nor U20967 (N_20967,N_20631,N_20693);
xnor U20968 (N_20968,N_20777,N_20615);
or U20969 (N_20969,N_20744,N_20637);
xor U20970 (N_20970,N_20682,N_20635);
nand U20971 (N_20971,N_20698,N_20739);
xnor U20972 (N_20972,N_20757,N_20666);
nand U20973 (N_20973,N_20663,N_20637);
nor U20974 (N_20974,N_20770,N_20694);
or U20975 (N_20975,N_20628,N_20797);
nand U20976 (N_20976,N_20712,N_20703);
nand U20977 (N_20977,N_20792,N_20677);
and U20978 (N_20978,N_20603,N_20736);
nor U20979 (N_20979,N_20707,N_20656);
xnor U20980 (N_20980,N_20701,N_20742);
and U20981 (N_20981,N_20601,N_20645);
nand U20982 (N_20982,N_20676,N_20741);
and U20983 (N_20983,N_20786,N_20728);
nor U20984 (N_20984,N_20715,N_20699);
and U20985 (N_20985,N_20774,N_20682);
nand U20986 (N_20986,N_20705,N_20720);
nand U20987 (N_20987,N_20768,N_20699);
xnor U20988 (N_20988,N_20754,N_20601);
nor U20989 (N_20989,N_20765,N_20671);
or U20990 (N_20990,N_20769,N_20659);
nand U20991 (N_20991,N_20729,N_20780);
and U20992 (N_20992,N_20639,N_20767);
nand U20993 (N_20993,N_20612,N_20745);
and U20994 (N_20994,N_20624,N_20619);
nor U20995 (N_20995,N_20699,N_20612);
xnor U20996 (N_20996,N_20711,N_20710);
nand U20997 (N_20997,N_20696,N_20701);
nand U20998 (N_20998,N_20637,N_20661);
xor U20999 (N_20999,N_20660,N_20752);
nor U21000 (N_21000,N_20886,N_20889);
nand U21001 (N_21001,N_20860,N_20985);
or U21002 (N_21002,N_20915,N_20897);
or U21003 (N_21003,N_20996,N_20937);
xor U21004 (N_21004,N_20977,N_20972);
or U21005 (N_21005,N_20984,N_20999);
nand U21006 (N_21006,N_20846,N_20938);
and U21007 (N_21007,N_20830,N_20819);
xor U21008 (N_21008,N_20918,N_20837);
nor U21009 (N_21009,N_20894,N_20914);
or U21010 (N_21010,N_20932,N_20913);
and U21011 (N_21011,N_20929,N_20962);
xnor U21012 (N_21012,N_20815,N_20992);
and U21013 (N_21013,N_20821,N_20858);
or U21014 (N_21014,N_20947,N_20877);
and U21015 (N_21015,N_20850,N_20901);
xnor U21016 (N_21016,N_20880,N_20824);
nand U21017 (N_21017,N_20807,N_20919);
or U21018 (N_21018,N_20958,N_20998);
and U21019 (N_21019,N_20853,N_20935);
or U21020 (N_21020,N_20867,N_20873);
nor U21021 (N_21021,N_20957,N_20809);
xor U21022 (N_21022,N_20812,N_20896);
nor U21023 (N_21023,N_20836,N_20834);
nand U21024 (N_21024,N_20995,N_20875);
or U21025 (N_21025,N_20816,N_20944);
or U21026 (N_21026,N_20868,N_20856);
or U21027 (N_21027,N_20951,N_20909);
nand U21028 (N_21028,N_20903,N_20843);
or U21029 (N_21029,N_20804,N_20931);
nand U21030 (N_21030,N_20863,N_20803);
xor U21031 (N_21031,N_20943,N_20939);
and U21032 (N_21032,N_20952,N_20832);
or U21033 (N_21033,N_20801,N_20974);
or U21034 (N_21034,N_20851,N_20982);
and U21035 (N_21035,N_20916,N_20805);
and U21036 (N_21036,N_20861,N_20912);
nand U21037 (N_21037,N_20956,N_20891);
nor U21038 (N_21038,N_20970,N_20988);
nand U21039 (N_21039,N_20862,N_20906);
xnor U21040 (N_21040,N_20884,N_20855);
xnor U21041 (N_21041,N_20849,N_20930);
nand U21042 (N_21042,N_20993,N_20865);
xnor U21043 (N_21043,N_20898,N_20927);
nand U21044 (N_21044,N_20847,N_20892);
nor U21045 (N_21045,N_20840,N_20802);
or U21046 (N_21046,N_20831,N_20978);
nand U21047 (N_21047,N_20902,N_20888);
and U21048 (N_21048,N_20808,N_20818);
or U21049 (N_21049,N_20997,N_20961);
and U21050 (N_21050,N_20965,N_20959);
xnor U21051 (N_21051,N_20940,N_20835);
xor U21052 (N_21052,N_20968,N_20981);
and U21053 (N_21053,N_20866,N_20922);
and U21054 (N_21054,N_20991,N_20989);
and U21055 (N_21055,N_20800,N_20920);
xnor U21056 (N_21056,N_20826,N_20990);
nand U21057 (N_21057,N_20882,N_20852);
xor U21058 (N_21058,N_20883,N_20828);
nand U21059 (N_21059,N_20841,N_20949);
nor U21060 (N_21060,N_20885,N_20859);
nand U21061 (N_21061,N_20833,N_20872);
nor U21062 (N_21062,N_20954,N_20946);
nor U21063 (N_21063,N_20923,N_20945);
xnor U21064 (N_21064,N_20910,N_20864);
nand U21065 (N_21065,N_20829,N_20911);
xor U21066 (N_21066,N_20994,N_20806);
nand U21067 (N_21067,N_20844,N_20924);
nor U21068 (N_21068,N_20960,N_20973);
xor U21069 (N_21069,N_20870,N_20823);
and U21070 (N_21070,N_20893,N_20905);
and U21071 (N_21071,N_20890,N_20857);
and U21072 (N_21072,N_20975,N_20917);
xnor U21073 (N_21073,N_20934,N_20810);
nand U21074 (N_21074,N_20936,N_20876);
xor U21075 (N_21075,N_20848,N_20955);
nand U21076 (N_21076,N_20842,N_20969);
or U21077 (N_21077,N_20887,N_20854);
and U21078 (N_21078,N_20869,N_20813);
nor U21079 (N_21079,N_20948,N_20921);
nand U21080 (N_21080,N_20879,N_20971);
xnor U21081 (N_21081,N_20964,N_20950);
and U21082 (N_21082,N_20926,N_20908);
and U21083 (N_21083,N_20986,N_20942);
and U21084 (N_21084,N_20874,N_20928);
xor U21085 (N_21085,N_20817,N_20933);
or U21086 (N_21086,N_20900,N_20976);
xor U21087 (N_21087,N_20979,N_20904);
or U21088 (N_21088,N_20983,N_20881);
xnor U21089 (N_21089,N_20825,N_20966);
nor U21090 (N_21090,N_20838,N_20907);
or U21091 (N_21091,N_20980,N_20925);
and U21092 (N_21092,N_20987,N_20878);
xnor U21093 (N_21093,N_20963,N_20820);
or U21094 (N_21094,N_20871,N_20839);
nor U21095 (N_21095,N_20953,N_20822);
nand U21096 (N_21096,N_20967,N_20941);
nor U21097 (N_21097,N_20827,N_20895);
or U21098 (N_21098,N_20899,N_20814);
nor U21099 (N_21099,N_20845,N_20811);
nor U21100 (N_21100,N_20990,N_20885);
xor U21101 (N_21101,N_20888,N_20920);
nor U21102 (N_21102,N_20979,N_20860);
xnor U21103 (N_21103,N_20995,N_20990);
xor U21104 (N_21104,N_20902,N_20970);
or U21105 (N_21105,N_20803,N_20917);
and U21106 (N_21106,N_20850,N_20868);
and U21107 (N_21107,N_20898,N_20955);
nor U21108 (N_21108,N_20912,N_20844);
nor U21109 (N_21109,N_20948,N_20832);
and U21110 (N_21110,N_20982,N_20949);
nor U21111 (N_21111,N_20833,N_20982);
nand U21112 (N_21112,N_20857,N_20925);
or U21113 (N_21113,N_20819,N_20805);
nor U21114 (N_21114,N_20940,N_20806);
nor U21115 (N_21115,N_20992,N_20915);
xor U21116 (N_21116,N_20829,N_20805);
xor U21117 (N_21117,N_20817,N_20922);
nand U21118 (N_21118,N_20879,N_20952);
and U21119 (N_21119,N_20975,N_20978);
or U21120 (N_21120,N_20800,N_20898);
xor U21121 (N_21121,N_20929,N_20914);
and U21122 (N_21122,N_20816,N_20998);
xor U21123 (N_21123,N_20882,N_20833);
or U21124 (N_21124,N_20998,N_20900);
or U21125 (N_21125,N_20942,N_20872);
nor U21126 (N_21126,N_20953,N_20885);
xor U21127 (N_21127,N_20984,N_20991);
nor U21128 (N_21128,N_20871,N_20883);
xor U21129 (N_21129,N_20947,N_20885);
nor U21130 (N_21130,N_20895,N_20853);
nand U21131 (N_21131,N_20968,N_20835);
and U21132 (N_21132,N_20956,N_20993);
and U21133 (N_21133,N_20995,N_20844);
or U21134 (N_21134,N_20880,N_20826);
nor U21135 (N_21135,N_20962,N_20857);
nor U21136 (N_21136,N_20831,N_20926);
xor U21137 (N_21137,N_20903,N_20933);
nand U21138 (N_21138,N_20924,N_20984);
nand U21139 (N_21139,N_20883,N_20951);
nand U21140 (N_21140,N_20806,N_20891);
and U21141 (N_21141,N_20928,N_20941);
nor U21142 (N_21142,N_20969,N_20960);
nand U21143 (N_21143,N_20953,N_20851);
and U21144 (N_21144,N_20932,N_20833);
or U21145 (N_21145,N_20904,N_20942);
or U21146 (N_21146,N_20976,N_20872);
or U21147 (N_21147,N_20888,N_20974);
nor U21148 (N_21148,N_20888,N_20864);
xor U21149 (N_21149,N_20804,N_20834);
nor U21150 (N_21150,N_20834,N_20827);
xor U21151 (N_21151,N_20977,N_20839);
and U21152 (N_21152,N_20937,N_20936);
nor U21153 (N_21153,N_20829,N_20881);
nor U21154 (N_21154,N_20937,N_20891);
nor U21155 (N_21155,N_20986,N_20821);
or U21156 (N_21156,N_20977,N_20958);
or U21157 (N_21157,N_20999,N_20818);
or U21158 (N_21158,N_20952,N_20918);
nand U21159 (N_21159,N_20954,N_20903);
xnor U21160 (N_21160,N_20975,N_20966);
or U21161 (N_21161,N_20873,N_20866);
and U21162 (N_21162,N_20989,N_20887);
or U21163 (N_21163,N_20962,N_20918);
xnor U21164 (N_21164,N_20847,N_20897);
and U21165 (N_21165,N_20954,N_20803);
and U21166 (N_21166,N_20947,N_20861);
and U21167 (N_21167,N_20913,N_20819);
xnor U21168 (N_21168,N_20901,N_20897);
nand U21169 (N_21169,N_20959,N_20832);
nand U21170 (N_21170,N_20949,N_20968);
or U21171 (N_21171,N_20941,N_20867);
and U21172 (N_21172,N_20948,N_20899);
and U21173 (N_21173,N_20804,N_20864);
xor U21174 (N_21174,N_20954,N_20929);
nor U21175 (N_21175,N_20884,N_20906);
nand U21176 (N_21176,N_20943,N_20966);
nor U21177 (N_21177,N_20956,N_20965);
nand U21178 (N_21178,N_20843,N_20868);
or U21179 (N_21179,N_20969,N_20847);
nand U21180 (N_21180,N_20919,N_20933);
nand U21181 (N_21181,N_20820,N_20917);
or U21182 (N_21182,N_20800,N_20974);
and U21183 (N_21183,N_20853,N_20979);
nand U21184 (N_21184,N_20865,N_20942);
nor U21185 (N_21185,N_20996,N_20949);
nand U21186 (N_21186,N_20967,N_20993);
nand U21187 (N_21187,N_20809,N_20984);
nor U21188 (N_21188,N_20995,N_20952);
or U21189 (N_21189,N_20866,N_20924);
and U21190 (N_21190,N_20994,N_20865);
nor U21191 (N_21191,N_20869,N_20987);
nor U21192 (N_21192,N_20853,N_20974);
nand U21193 (N_21193,N_20867,N_20959);
nand U21194 (N_21194,N_20999,N_20859);
or U21195 (N_21195,N_20901,N_20997);
xnor U21196 (N_21196,N_20967,N_20942);
or U21197 (N_21197,N_20981,N_20918);
and U21198 (N_21198,N_20952,N_20915);
and U21199 (N_21199,N_20987,N_20875);
and U21200 (N_21200,N_21197,N_21186);
xnor U21201 (N_21201,N_21137,N_21038);
xnor U21202 (N_21202,N_21127,N_21098);
nand U21203 (N_21203,N_21088,N_21108);
or U21204 (N_21204,N_21151,N_21181);
xor U21205 (N_21205,N_21077,N_21100);
or U21206 (N_21206,N_21189,N_21168);
or U21207 (N_21207,N_21183,N_21152);
nand U21208 (N_21208,N_21075,N_21136);
nand U21209 (N_21209,N_21061,N_21033);
or U21210 (N_21210,N_21079,N_21138);
nor U21211 (N_21211,N_21162,N_21103);
and U21212 (N_21212,N_21132,N_21032);
xnor U21213 (N_21213,N_21121,N_21131);
xor U21214 (N_21214,N_21135,N_21196);
and U21215 (N_21215,N_21052,N_21110);
and U21216 (N_21216,N_21027,N_21064);
and U21217 (N_21217,N_21195,N_21089);
and U21218 (N_21218,N_21024,N_21040);
and U21219 (N_21219,N_21099,N_21170);
xnor U21220 (N_21220,N_21199,N_21072);
or U21221 (N_21221,N_21120,N_21028);
or U21222 (N_21222,N_21109,N_21125);
or U21223 (N_21223,N_21182,N_21045);
or U21224 (N_21224,N_21080,N_21043);
or U21225 (N_21225,N_21046,N_21025);
nand U21226 (N_21226,N_21093,N_21063);
xnor U21227 (N_21227,N_21022,N_21185);
nand U21228 (N_21228,N_21115,N_21047);
or U21229 (N_21229,N_21164,N_21154);
and U21230 (N_21230,N_21039,N_21113);
nor U21231 (N_21231,N_21056,N_21163);
nand U21232 (N_21232,N_21020,N_21086);
xnor U21233 (N_21233,N_21034,N_21076);
nand U21234 (N_21234,N_21101,N_21190);
nand U21235 (N_21235,N_21074,N_21092);
nand U21236 (N_21236,N_21083,N_21096);
or U21237 (N_21237,N_21147,N_21078);
xnor U21238 (N_21238,N_21161,N_21065);
nor U21239 (N_21239,N_21014,N_21019);
nand U21240 (N_21240,N_21126,N_21174);
xor U21241 (N_21241,N_21130,N_21010);
nor U21242 (N_21242,N_21134,N_21143);
xor U21243 (N_21243,N_21193,N_21128);
nand U21244 (N_21244,N_21165,N_21012);
and U21245 (N_21245,N_21084,N_21102);
nor U21246 (N_21246,N_21142,N_21104);
xor U21247 (N_21247,N_21119,N_21026);
nor U21248 (N_21248,N_21166,N_21018);
nor U21249 (N_21249,N_21123,N_21017);
nor U21250 (N_21250,N_21058,N_21000);
xor U21251 (N_21251,N_21037,N_21050);
nor U21252 (N_21252,N_21107,N_21062);
nand U21253 (N_21253,N_21031,N_21124);
xor U21254 (N_21254,N_21175,N_21179);
or U21255 (N_21255,N_21071,N_21009);
xnor U21256 (N_21256,N_21188,N_21060);
and U21257 (N_21257,N_21003,N_21011);
or U21258 (N_21258,N_21035,N_21157);
xnor U21259 (N_21259,N_21048,N_21111);
or U21260 (N_21260,N_21081,N_21067);
nor U21261 (N_21261,N_21148,N_21149);
or U21262 (N_21262,N_21005,N_21095);
and U21263 (N_21263,N_21187,N_21153);
and U21264 (N_21264,N_21070,N_21159);
and U21265 (N_21265,N_21097,N_21091);
and U21266 (N_21266,N_21044,N_21007);
and U21267 (N_21267,N_21041,N_21090);
nand U21268 (N_21268,N_21051,N_21169);
nor U21269 (N_21269,N_21150,N_21192);
or U21270 (N_21270,N_21172,N_21114);
nand U21271 (N_21271,N_21144,N_21105);
or U21272 (N_21272,N_21085,N_21069);
or U21273 (N_21273,N_21054,N_21140);
nand U21274 (N_21274,N_21156,N_21118);
xnor U21275 (N_21275,N_21049,N_21176);
nor U21276 (N_21276,N_21194,N_21015);
nand U21277 (N_21277,N_21006,N_21133);
or U21278 (N_21278,N_21198,N_21029);
xnor U21279 (N_21279,N_21059,N_21001);
nand U21280 (N_21280,N_21117,N_21167);
xor U21281 (N_21281,N_21030,N_21002);
nand U21282 (N_21282,N_21139,N_21146);
xnor U21283 (N_21283,N_21013,N_21094);
nor U21284 (N_21284,N_21082,N_21145);
or U21285 (N_21285,N_21106,N_21155);
xnor U21286 (N_21286,N_21129,N_21180);
nand U21287 (N_21287,N_21116,N_21055);
and U21288 (N_21288,N_21073,N_21008);
xnor U21289 (N_21289,N_21066,N_21004);
nand U21290 (N_21290,N_21184,N_21122);
or U21291 (N_21291,N_21191,N_21171);
nand U21292 (N_21292,N_21042,N_21021);
xnor U21293 (N_21293,N_21112,N_21023);
or U21294 (N_21294,N_21158,N_21087);
xnor U21295 (N_21295,N_21141,N_21016);
nand U21296 (N_21296,N_21057,N_21178);
xnor U21297 (N_21297,N_21160,N_21068);
nand U21298 (N_21298,N_21173,N_21053);
nor U21299 (N_21299,N_21036,N_21177);
nand U21300 (N_21300,N_21108,N_21105);
and U21301 (N_21301,N_21096,N_21100);
and U21302 (N_21302,N_21149,N_21155);
nor U21303 (N_21303,N_21130,N_21009);
and U21304 (N_21304,N_21029,N_21183);
xor U21305 (N_21305,N_21037,N_21092);
or U21306 (N_21306,N_21161,N_21007);
nor U21307 (N_21307,N_21089,N_21154);
or U21308 (N_21308,N_21105,N_21124);
xor U21309 (N_21309,N_21138,N_21165);
and U21310 (N_21310,N_21004,N_21040);
nor U21311 (N_21311,N_21156,N_21080);
nor U21312 (N_21312,N_21194,N_21053);
nand U21313 (N_21313,N_21071,N_21040);
nor U21314 (N_21314,N_21148,N_21033);
and U21315 (N_21315,N_21142,N_21091);
or U21316 (N_21316,N_21139,N_21101);
xor U21317 (N_21317,N_21016,N_21125);
nand U21318 (N_21318,N_21126,N_21108);
nand U21319 (N_21319,N_21135,N_21084);
or U21320 (N_21320,N_21055,N_21050);
nor U21321 (N_21321,N_21010,N_21140);
or U21322 (N_21322,N_21038,N_21162);
nor U21323 (N_21323,N_21027,N_21130);
or U21324 (N_21324,N_21146,N_21129);
nor U21325 (N_21325,N_21176,N_21041);
nand U21326 (N_21326,N_21084,N_21187);
and U21327 (N_21327,N_21156,N_21185);
xor U21328 (N_21328,N_21137,N_21128);
or U21329 (N_21329,N_21013,N_21049);
nor U21330 (N_21330,N_21014,N_21176);
and U21331 (N_21331,N_21045,N_21147);
and U21332 (N_21332,N_21028,N_21068);
or U21333 (N_21333,N_21096,N_21147);
or U21334 (N_21334,N_21011,N_21179);
or U21335 (N_21335,N_21018,N_21105);
and U21336 (N_21336,N_21198,N_21126);
nand U21337 (N_21337,N_21005,N_21181);
nand U21338 (N_21338,N_21114,N_21152);
xnor U21339 (N_21339,N_21095,N_21070);
or U21340 (N_21340,N_21193,N_21160);
xor U21341 (N_21341,N_21040,N_21006);
and U21342 (N_21342,N_21178,N_21187);
nor U21343 (N_21343,N_21187,N_21132);
or U21344 (N_21344,N_21043,N_21022);
xnor U21345 (N_21345,N_21121,N_21024);
or U21346 (N_21346,N_21090,N_21143);
or U21347 (N_21347,N_21043,N_21077);
nand U21348 (N_21348,N_21035,N_21085);
and U21349 (N_21349,N_21039,N_21037);
nor U21350 (N_21350,N_21047,N_21192);
xnor U21351 (N_21351,N_21067,N_21136);
and U21352 (N_21352,N_21136,N_21102);
xnor U21353 (N_21353,N_21086,N_21189);
nor U21354 (N_21354,N_21027,N_21175);
xnor U21355 (N_21355,N_21045,N_21037);
nand U21356 (N_21356,N_21191,N_21064);
nor U21357 (N_21357,N_21032,N_21165);
or U21358 (N_21358,N_21129,N_21026);
nand U21359 (N_21359,N_21158,N_21093);
nor U21360 (N_21360,N_21040,N_21194);
nand U21361 (N_21361,N_21027,N_21108);
xor U21362 (N_21362,N_21020,N_21012);
nand U21363 (N_21363,N_21069,N_21048);
xnor U21364 (N_21364,N_21069,N_21151);
and U21365 (N_21365,N_21194,N_21043);
or U21366 (N_21366,N_21101,N_21089);
or U21367 (N_21367,N_21180,N_21156);
or U21368 (N_21368,N_21165,N_21075);
nand U21369 (N_21369,N_21151,N_21003);
nor U21370 (N_21370,N_21124,N_21101);
nand U21371 (N_21371,N_21055,N_21074);
xor U21372 (N_21372,N_21038,N_21091);
and U21373 (N_21373,N_21075,N_21057);
xnor U21374 (N_21374,N_21082,N_21054);
nand U21375 (N_21375,N_21016,N_21159);
nand U21376 (N_21376,N_21175,N_21154);
nand U21377 (N_21377,N_21007,N_21122);
xnor U21378 (N_21378,N_21176,N_21135);
and U21379 (N_21379,N_21018,N_21179);
and U21380 (N_21380,N_21114,N_21194);
and U21381 (N_21381,N_21082,N_21105);
nand U21382 (N_21382,N_21137,N_21086);
nand U21383 (N_21383,N_21069,N_21119);
nor U21384 (N_21384,N_21145,N_21197);
xnor U21385 (N_21385,N_21131,N_21001);
nand U21386 (N_21386,N_21077,N_21168);
nand U21387 (N_21387,N_21114,N_21077);
and U21388 (N_21388,N_21083,N_21057);
xnor U21389 (N_21389,N_21074,N_21068);
xor U21390 (N_21390,N_21057,N_21150);
and U21391 (N_21391,N_21007,N_21116);
nand U21392 (N_21392,N_21014,N_21149);
or U21393 (N_21393,N_21018,N_21178);
and U21394 (N_21394,N_21183,N_21134);
nor U21395 (N_21395,N_21155,N_21091);
or U21396 (N_21396,N_21008,N_21179);
xnor U21397 (N_21397,N_21084,N_21005);
and U21398 (N_21398,N_21174,N_21003);
nor U21399 (N_21399,N_21012,N_21068);
and U21400 (N_21400,N_21348,N_21238);
and U21401 (N_21401,N_21253,N_21295);
xor U21402 (N_21402,N_21379,N_21377);
and U21403 (N_21403,N_21311,N_21209);
xor U21404 (N_21404,N_21359,N_21251);
nor U21405 (N_21405,N_21213,N_21387);
nand U21406 (N_21406,N_21307,N_21200);
and U21407 (N_21407,N_21331,N_21284);
nand U21408 (N_21408,N_21220,N_21246);
nand U21409 (N_21409,N_21369,N_21273);
nor U21410 (N_21410,N_21279,N_21249);
and U21411 (N_21411,N_21399,N_21393);
nor U21412 (N_21412,N_21226,N_21340);
nor U21413 (N_21413,N_21292,N_21293);
or U21414 (N_21414,N_21208,N_21385);
or U21415 (N_21415,N_21265,N_21243);
and U21416 (N_21416,N_21262,N_21276);
nor U21417 (N_21417,N_21383,N_21366);
nand U21418 (N_21418,N_21303,N_21339);
or U21419 (N_21419,N_21352,N_21321);
xnor U21420 (N_21420,N_21228,N_21334);
and U21421 (N_21421,N_21298,N_21290);
xor U21422 (N_21422,N_21313,N_21382);
or U21423 (N_21423,N_21223,N_21304);
nand U21424 (N_21424,N_21349,N_21212);
nor U21425 (N_21425,N_21329,N_21288);
xor U21426 (N_21426,N_21363,N_21332);
or U21427 (N_21427,N_21232,N_21322);
and U21428 (N_21428,N_21234,N_21373);
or U21429 (N_21429,N_21204,N_21309);
and U21430 (N_21430,N_21218,N_21239);
nand U21431 (N_21431,N_21299,N_21241);
or U21432 (N_21432,N_21378,N_21353);
nand U21433 (N_21433,N_21355,N_21229);
xnor U21434 (N_21434,N_21328,N_21222);
xor U21435 (N_21435,N_21207,N_21381);
nor U21436 (N_21436,N_21274,N_21255);
or U21437 (N_21437,N_21296,N_21354);
nand U21438 (N_21438,N_21257,N_21390);
nand U21439 (N_21439,N_21275,N_21240);
or U21440 (N_21440,N_21283,N_21286);
nor U21441 (N_21441,N_21395,N_21269);
and U21442 (N_21442,N_21326,N_21384);
xnor U21443 (N_21443,N_21314,N_21398);
nor U21444 (N_21444,N_21345,N_21291);
nand U21445 (N_21445,N_21225,N_21396);
or U21446 (N_21446,N_21260,N_21256);
or U21447 (N_21447,N_21277,N_21245);
nand U21448 (N_21448,N_21315,N_21259);
or U21449 (N_21449,N_21203,N_21319);
and U21450 (N_21450,N_21372,N_21221);
nor U21451 (N_21451,N_21394,N_21310);
nand U21452 (N_21452,N_21312,N_21210);
nand U21453 (N_21453,N_21282,N_21327);
or U21454 (N_21454,N_21306,N_21356);
nand U21455 (N_21455,N_21237,N_21272);
nand U21456 (N_21456,N_21337,N_21280);
nand U21457 (N_21457,N_21201,N_21324);
xnor U21458 (N_21458,N_21323,N_21357);
nand U21459 (N_21459,N_21294,N_21285);
and U21460 (N_21460,N_21347,N_21344);
and U21461 (N_21461,N_21270,N_21287);
nand U21462 (N_21462,N_21250,N_21278);
and U21463 (N_21463,N_21342,N_21367);
xor U21464 (N_21464,N_21230,N_21330);
or U21465 (N_21465,N_21302,N_21317);
xnor U21466 (N_21466,N_21267,N_21271);
and U21467 (N_21467,N_21215,N_21219);
xor U21468 (N_21468,N_21325,N_21380);
and U21469 (N_21469,N_21397,N_21289);
nor U21470 (N_21470,N_21333,N_21214);
nor U21471 (N_21471,N_21346,N_21268);
and U21472 (N_21472,N_21391,N_21266);
and U21473 (N_21473,N_21248,N_21335);
xor U21474 (N_21474,N_21318,N_21336);
and U21475 (N_21475,N_21308,N_21368);
and U21476 (N_21476,N_21361,N_21343);
nor U21477 (N_21477,N_21300,N_21264);
nand U21478 (N_21478,N_21224,N_21236);
nor U21479 (N_21479,N_21358,N_21297);
or U21480 (N_21480,N_21388,N_21301);
nor U21481 (N_21481,N_21261,N_21376);
nand U21482 (N_21482,N_21216,N_21371);
nor U21483 (N_21483,N_21254,N_21247);
and U21484 (N_21484,N_21235,N_21341);
or U21485 (N_21485,N_21392,N_21211);
and U21486 (N_21486,N_21205,N_21374);
xor U21487 (N_21487,N_21362,N_21365);
and U21488 (N_21488,N_21305,N_21217);
nand U21489 (N_21489,N_21252,N_21227);
nand U21490 (N_21490,N_21370,N_21375);
nor U21491 (N_21491,N_21360,N_21281);
or U21492 (N_21492,N_21389,N_21242);
xor U21493 (N_21493,N_21320,N_21233);
and U21494 (N_21494,N_21338,N_21202);
and U21495 (N_21495,N_21350,N_21231);
nor U21496 (N_21496,N_21386,N_21244);
and U21497 (N_21497,N_21316,N_21206);
nand U21498 (N_21498,N_21263,N_21364);
and U21499 (N_21499,N_21351,N_21258);
and U21500 (N_21500,N_21346,N_21389);
and U21501 (N_21501,N_21242,N_21359);
nor U21502 (N_21502,N_21228,N_21205);
xor U21503 (N_21503,N_21258,N_21293);
and U21504 (N_21504,N_21362,N_21298);
nor U21505 (N_21505,N_21361,N_21306);
xnor U21506 (N_21506,N_21324,N_21203);
nand U21507 (N_21507,N_21319,N_21363);
xor U21508 (N_21508,N_21337,N_21263);
and U21509 (N_21509,N_21230,N_21379);
nand U21510 (N_21510,N_21353,N_21375);
xor U21511 (N_21511,N_21327,N_21370);
xor U21512 (N_21512,N_21359,N_21245);
nor U21513 (N_21513,N_21324,N_21307);
and U21514 (N_21514,N_21229,N_21209);
or U21515 (N_21515,N_21281,N_21367);
and U21516 (N_21516,N_21317,N_21288);
xnor U21517 (N_21517,N_21211,N_21274);
nand U21518 (N_21518,N_21243,N_21239);
or U21519 (N_21519,N_21313,N_21396);
nor U21520 (N_21520,N_21253,N_21240);
or U21521 (N_21521,N_21226,N_21362);
or U21522 (N_21522,N_21263,N_21339);
or U21523 (N_21523,N_21397,N_21311);
xor U21524 (N_21524,N_21388,N_21265);
nand U21525 (N_21525,N_21315,N_21253);
nor U21526 (N_21526,N_21358,N_21331);
nand U21527 (N_21527,N_21289,N_21228);
or U21528 (N_21528,N_21214,N_21241);
or U21529 (N_21529,N_21265,N_21228);
xor U21530 (N_21530,N_21313,N_21218);
and U21531 (N_21531,N_21377,N_21256);
nand U21532 (N_21532,N_21367,N_21226);
nor U21533 (N_21533,N_21281,N_21208);
nand U21534 (N_21534,N_21398,N_21258);
nand U21535 (N_21535,N_21399,N_21302);
nor U21536 (N_21536,N_21351,N_21277);
nor U21537 (N_21537,N_21320,N_21246);
xor U21538 (N_21538,N_21263,N_21204);
and U21539 (N_21539,N_21387,N_21365);
and U21540 (N_21540,N_21252,N_21272);
nand U21541 (N_21541,N_21397,N_21318);
xnor U21542 (N_21542,N_21295,N_21354);
nand U21543 (N_21543,N_21394,N_21344);
or U21544 (N_21544,N_21301,N_21302);
xor U21545 (N_21545,N_21384,N_21204);
and U21546 (N_21546,N_21300,N_21357);
nand U21547 (N_21547,N_21274,N_21387);
or U21548 (N_21548,N_21268,N_21361);
xor U21549 (N_21549,N_21272,N_21314);
nor U21550 (N_21550,N_21381,N_21332);
xnor U21551 (N_21551,N_21266,N_21214);
nor U21552 (N_21552,N_21351,N_21355);
or U21553 (N_21553,N_21363,N_21381);
and U21554 (N_21554,N_21372,N_21338);
nor U21555 (N_21555,N_21328,N_21300);
or U21556 (N_21556,N_21217,N_21383);
nand U21557 (N_21557,N_21362,N_21356);
xor U21558 (N_21558,N_21366,N_21260);
nor U21559 (N_21559,N_21241,N_21217);
xnor U21560 (N_21560,N_21276,N_21341);
xor U21561 (N_21561,N_21392,N_21397);
nor U21562 (N_21562,N_21226,N_21314);
and U21563 (N_21563,N_21230,N_21267);
or U21564 (N_21564,N_21203,N_21391);
nor U21565 (N_21565,N_21282,N_21372);
and U21566 (N_21566,N_21356,N_21234);
and U21567 (N_21567,N_21209,N_21241);
xnor U21568 (N_21568,N_21399,N_21232);
nand U21569 (N_21569,N_21295,N_21272);
xnor U21570 (N_21570,N_21270,N_21323);
nor U21571 (N_21571,N_21297,N_21375);
nor U21572 (N_21572,N_21317,N_21240);
xor U21573 (N_21573,N_21256,N_21391);
or U21574 (N_21574,N_21285,N_21398);
nor U21575 (N_21575,N_21364,N_21299);
xor U21576 (N_21576,N_21294,N_21375);
nor U21577 (N_21577,N_21325,N_21226);
xor U21578 (N_21578,N_21322,N_21284);
nand U21579 (N_21579,N_21240,N_21291);
nor U21580 (N_21580,N_21231,N_21308);
nor U21581 (N_21581,N_21333,N_21308);
xor U21582 (N_21582,N_21366,N_21326);
and U21583 (N_21583,N_21384,N_21317);
nor U21584 (N_21584,N_21200,N_21380);
nor U21585 (N_21585,N_21205,N_21301);
and U21586 (N_21586,N_21310,N_21253);
nor U21587 (N_21587,N_21301,N_21357);
xor U21588 (N_21588,N_21273,N_21321);
and U21589 (N_21589,N_21361,N_21308);
or U21590 (N_21590,N_21204,N_21331);
nand U21591 (N_21591,N_21319,N_21381);
xnor U21592 (N_21592,N_21202,N_21342);
nor U21593 (N_21593,N_21362,N_21264);
and U21594 (N_21594,N_21251,N_21325);
nor U21595 (N_21595,N_21353,N_21329);
or U21596 (N_21596,N_21341,N_21364);
or U21597 (N_21597,N_21284,N_21249);
and U21598 (N_21598,N_21381,N_21289);
nand U21599 (N_21599,N_21245,N_21230);
nor U21600 (N_21600,N_21555,N_21432);
or U21601 (N_21601,N_21485,N_21576);
xnor U21602 (N_21602,N_21490,N_21530);
xor U21603 (N_21603,N_21428,N_21435);
and U21604 (N_21604,N_21588,N_21481);
nand U21605 (N_21605,N_21492,N_21478);
nand U21606 (N_21606,N_21438,N_21529);
nor U21607 (N_21607,N_21532,N_21427);
xnor U21608 (N_21608,N_21519,N_21509);
or U21609 (N_21609,N_21513,N_21512);
xnor U21610 (N_21610,N_21520,N_21568);
nand U21611 (N_21611,N_21420,N_21467);
nand U21612 (N_21612,N_21452,N_21543);
nand U21613 (N_21613,N_21589,N_21521);
and U21614 (N_21614,N_21422,N_21417);
and U21615 (N_21615,N_21590,N_21510);
nand U21616 (N_21616,N_21415,N_21592);
nor U21617 (N_21617,N_21430,N_21462);
and U21618 (N_21618,N_21461,N_21595);
and U21619 (N_21619,N_21434,N_21571);
or U21620 (N_21620,N_21561,N_21491);
or U21621 (N_21621,N_21414,N_21448);
and U21622 (N_21622,N_21525,N_21507);
or U21623 (N_21623,N_21538,N_21409);
nor U21624 (N_21624,N_21559,N_21431);
or U21625 (N_21625,N_21488,N_21468);
nand U21626 (N_21626,N_21551,N_21522);
xor U21627 (N_21627,N_21433,N_21524);
xnor U21628 (N_21628,N_21426,N_21483);
nor U21629 (N_21629,N_21552,N_21572);
nor U21630 (N_21630,N_21472,N_21556);
nor U21631 (N_21631,N_21449,N_21496);
nand U21632 (N_21632,N_21464,N_21407);
or U21633 (N_21633,N_21436,N_21503);
and U21634 (N_21634,N_21587,N_21563);
and U21635 (N_21635,N_21564,N_21515);
and U21636 (N_21636,N_21534,N_21540);
or U21637 (N_21637,N_21402,N_21403);
or U21638 (N_21638,N_21498,N_21575);
or U21639 (N_21639,N_21593,N_21470);
and U21640 (N_21640,N_21514,N_21406);
or U21641 (N_21641,N_21501,N_21482);
xor U21642 (N_21642,N_21526,N_21594);
nand U21643 (N_21643,N_21458,N_21446);
or U21644 (N_21644,N_21505,N_21545);
nor U21645 (N_21645,N_21421,N_21573);
nor U21646 (N_21646,N_21574,N_21447);
and U21647 (N_21647,N_21566,N_21480);
and U21648 (N_21648,N_21580,N_21598);
and U21649 (N_21649,N_21456,N_21484);
or U21650 (N_21650,N_21475,N_21554);
and U21651 (N_21651,N_21533,N_21504);
xor U21652 (N_21652,N_21547,N_21453);
nand U21653 (N_21653,N_21429,N_21550);
nor U21654 (N_21654,N_21549,N_21455);
or U21655 (N_21655,N_21579,N_21599);
and U21656 (N_21656,N_21451,N_21546);
xor U21657 (N_21657,N_21493,N_21445);
and U21658 (N_21658,N_21401,N_21591);
nor U21659 (N_21659,N_21404,N_21528);
or U21660 (N_21660,N_21466,N_21539);
and U21661 (N_21661,N_21405,N_21500);
and U21662 (N_21662,N_21518,N_21494);
xnor U21663 (N_21663,N_21584,N_21531);
nor U21664 (N_21664,N_21544,N_21450);
nand U21665 (N_21665,N_21585,N_21410);
nor U21666 (N_21666,N_21437,N_21558);
and U21667 (N_21667,N_21440,N_21567);
nand U21668 (N_21668,N_21516,N_21460);
nor U21669 (N_21669,N_21562,N_21497);
or U21670 (N_21670,N_21418,N_21471);
nand U21671 (N_21671,N_21444,N_21413);
or U21672 (N_21672,N_21583,N_21557);
and U21673 (N_21673,N_21535,N_21473);
xor U21674 (N_21674,N_21465,N_21477);
and U21675 (N_21675,N_21577,N_21495);
nor U21676 (N_21676,N_21586,N_21411);
and U21677 (N_21677,N_21474,N_21578);
and U21678 (N_21678,N_21487,N_21469);
or U21679 (N_21679,N_21419,N_21548);
or U21680 (N_21680,N_21560,N_21442);
nand U21681 (N_21681,N_21424,N_21523);
nor U21682 (N_21682,N_21408,N_21536);
nor U21683 (N_21683,N_21457,N_21506);
and U21684 (N_21684,N_21412,N_21541);
nor U21685 (N_21685,N_21570,N_21486);
xor U21686 (N_21686,N_21581,N_21569);
xor U21687 (N_21687,N_21443,N_21553);
and U21688 (N_21688,N_21565,N_21454);
or U21689 (N_21689,N_21463,N_21425);
xnor U21690 (N_21690,N_21459,N_21439);
and U21691 (N_21691,N_21479,N_21502);
nor U21692 (N_21692,N_21489,N_21416);
nor U21693 (N_21693,N_21441,N_21511);
and U21694 (N_21694,N_21537,N_21582);
xnor U21695 (N_21695,N_21423,N_21476);
and U21696 (N_21696,N_21597,N_21542);
and U21697 (N_21697,N_21400,N_21596);
nand U21698 (N_21698,N_21499,N_21527);
and U21699 (N_21699,N_21508,N_21517);
xnor U21700 (N_21700,N_21448,N_21416);
xnor U21701 (N_21701,N_21585,N_21568);
xor U21702 (N_21702,N_21478,N_21449);
xnor U21703 (N_21703,N_21410,N_21411);
nor U21704 (N_21704,N_21547,N_21408);
nor U21705 (N_21705,N_21492,N_21475);
xnor U21706 (N_21706,N_21554,N_21463);
or U21707 (N_21707,N_21469,N_21546);
nand U21708 (N_21708,N_21457,N_21585);
and U21709 (N_21709,N_21434,N_21535);
nand U21710 (N_21710,N_21428,N_21560);
nand U21711 (N_21711,N_21431,N_21573);
and U21712 (N_21712,N_21550,N_21446);
or U21713 (N_21713,N_21508,N_21458);
xor U21714 (N_21714,N_21420,N_21530);
nor U21715 (N_21715,N_21559,N_21543);
or U21716 (N_21716,N_21525,N_21475);
or U21717 (N_21717,N_21502,N_21431);
xnor U21718 (N_21718,N_21481,N_21446);
nor U21719 (N_21719,N_21551,N_21418);
or U21720 (N_21720,N_21406,N_21458);
nor U21721 (N_21721,N_21453,N_21488);
and U21722 (N_21722,N_21500,N_21437);
and U21723 (N_21723,N_21504,N_21472);
nand U21724 (N_21724,N_21563,N_21564);
nor U21725 (N_21725,N_21411,N_21488);
nand U21726 (N_21726,N_21531,N_21481);
and U21727 (N_21727,N_21450,N_21502);
and U21728 (N_21728,N_21408,N_21569);
nor U21729 (N_21729,N_21502,N_21456);
xnor U21730 (N_21730,N_21404,N_21491);
nor U21731 (N_21731,N_21499,N_21539);
nand U21732 (N_21732,N_21574,N_21477);
nor U21733 (N_21733,N_21535,N_21445);
nand U21734 (N_21734,N_21433,N_21454);
xnor U21735 (N_21735,N_21577,N_21439);
and U21736 (N_21736,N_21468,N_21514);
nand U21737 (N_21737,N_21435,N_21507);
nor U21738 (N_21738,N_21499,N_21522);
and U21739 (N_21739,N_21507,N_21422);
xnor U21740 (N_21740,N_21532,N_21498);
or U21741 (N_21741,N_21542,N_21599);
and U21742 (N_21742,N_21460,N_21555);
xnor U21743 (N_21743,N_21486,N_21469);
nand U21744 (N_21744,N_21538,N_21598);
xnor U21745 (N_21745,N_21519,N_21518);
and U21746 (N_21746,N_21410,N_21404);
nand U21747 (N_21747,N_21533,N_21459);
nand U21748 (N_21748,N_21406,N_21476);
nor U21749 (N_21749,N_21489,N_21507);
xor U21750 (N_21750,N_21423,N_21467);
xor U21751 (N_21751,N_21521,N_21431);
nor U21752 (N_21752,N_21518,N_21581);
xor U21753 (N_21753,N_21459,N_21535);
nand U21754 (N_21754,N_21595,N_21487);
nand U21755 (N_21755,N_21468,N_21446);
xnor U21756 (N_21756,N_21463,N_21440);
nand U21757 (N_21757,N_21433,N_21534);
nand U21758 (N_21758,N_21427,N_21562);
or U21759 (N_21759,N_21595,N_21490);
xor U21760 (N_21760,N_21543,N_21571);
nor U21761 (N_21761,N_21450,N_21556);
xnor U21762 (N_21762,N_21528,N_21538);
xnor U21763 (N_21763,N_21512,N_21434);
nand U21764 (N_21764,N_21482,N_21567);
and U21765 (N_21765,N_21570,N_21455);
or U21766 (N_21766,N_21544,N_21501);
and U21767 (N_21767,N_21572,N_21568);
nor U21768 (N_21768,N_21437,N_21429);
nand U21769 (N_21769,N_21428,N_21437);
and U21770 (N_21770,N_21498,N_21493);
and U21771 (N_21771,N_21418,N_21459);
nor U21772 (N_21772,N_21551,N_21544);
xor U21773 (N_21773,N_21562,N_21442);
nor U21774 (N_21774,N_21449,N_21425);
and U21775 (N_21775,N_21438,N_21599);
xor U21776 (N_21776,N_21444,N_21530);
nand U21777 (N_21777,N_21578,N_21574);
nor U21778 (N_21778,N_21471,N_21597);
nand U21779 (N_21779,N_21506,N_21549);
nand U21780 (N_21780,N_21523,N_21564);
or U21781 (N_21781,N_21445,N_21450);
nor U21782 (N_21782,N_21502,N_21495);
nand U21783 (N_21783,N_21422,N_21493);
nand U21784 (N_21784,N_21569,N_21527);
xnor U21785 (N_21785,N_21523,N_21556);
xnor U21786 (N_21786,N_21431,N_21519);
or U21787 (N_21787,N_21594,N_21515);
and U21788 (N_21788,N_21552,N_21487);
nor U21789 (N_21789,N_21591,N_21595);
xor U21790 (N_21790,N_21456,N_21592);
or U21791 (N_21791,N_21534,N_21422);
or U21792 (N_21792,N_21454,N_21463);
or U21793 (N_21793,N_21431,N_21510);
nor U21794 (N_21794,N_21582,N_21563);
nor U21795 (N_21795,N_21418,N_21408);
xor U21796 (N_21796,N_21504,N_21576);
and U21797 (N_21797,N_21400,N_21460);
and U21798 (N_21798,N_21480,N_21553);
or U21799 (N_21799,N_21423,N_21487);
and U21800 (N_21800,N_21608,N_21699);
and U21801 (N_21801,N_21635,N_21636);
nand U21802 (N_21802,N_21642,N_21655);
or U21803 (N_21803,N_21613,N_21738);
and U21804 (N_21804,N_21612,N_21764);
nor U21805 (N_21805,N_21639,N_21785);
xnor U21806 (N_21806,N_21763,N_21783);
nand U21807 (N_21807,N_21634,N_21615);
and U21808 (N_21808,N_21669,N_21739);
xnor U21809 (N_21809,N_21743,N_21653);
nor U21810 (N_21810,N_21605,N_21792);
nor U21811 (N_21811,N_21771,N_21647);
xor U21812 (N_21812,N_21694,N_21777);
nand U21813 (N_21813,N_21787,N_21791);
nand U21814 (N_21814,N_21610,N_21640);
nand U21815 (N_21815,N_21600,N_21652);
xor U21816 (N_21816,N_21650,N_21759);
nor U21817 (N_21817,N_21724,N_21799);
and U21818 (N_21818,N_21670,N_21621);
nor U21819 (N_21819,N_21625,N_21609);
nor U21820 (N_21820,N_21614,N_21618);
nand U21821 (N_21821,N_21775,N_21681);
nor U21822 (N_21822,N_21638,N_21797);
or U21823 (N_21823,N_21692,N_21667);
xor U21824 (N_21824,N_21637,N_21794);
nor U21825 (N_21825,N_21668,N_21644);
nand U21826 (N_21826,N_21672,N_21690);
and U21827 (N_21827,N_21740,N_21781);
and U21828 (N_21828,N_21676,N_21732);
or U21829 (N_21829,N_21796,N_21633);
nand U21830 (N_21830,N_21627,N_21616);
nand U21831 (N_21831,N_21760,N_21623);
and U21832 (N_21832,N_21719,N_21604);
nor U21833 (N_21833,N_21720,N_21680);
nor U21834 (N_21834,N_21671,N_21712);
xor U21835 (N_21835,N_21659,N_21651);
nor U21836 (N_21836,N_21749,N_21761);
nor U21837 (N_21837,N_21663,N_21751);
or U21838 (N_21838,N_21767,N_21766);
xor U21839 (N_21839,N_21774,N_21730);
or U21840 (N_21840,N_21688,N_21722);
and U21841 (N_21841,N_21687,N_21649);
xor U21842 (N_21842,N_21619,N_21714);
nor U21843 (N_21843,N_21717,N_21675);
nand U21844 (N_21844,N_21603,N_21683);
nand U21845 (N_21845,N_21744,N_21757);
and U21846 (N_21846,N_21753,N_21602);
xor U21847 (N_21847,N_21691,N_21700);
nor U21848 (N_21848,N_21735,N_21752);
nor U21849 (N_21849,N_21762,N_21657);
nand U21850 (N_21850,N_21708,N_21678);
nor U21851 (N_21851,N_21745,N_21758);
nor U21852 (N_21852,N_21679,N_21772);
nand U21853 (N_21853,N_21734,N_21696);
nand U21854 (N_21854,N_21628,N_21666);
and U21855 (N_21855,N_21790,N_21756);
or U21856 (N_21856,N_21674,N_21742);
and U21857 (N_21857,N_21755,N_21773);
xnor U21858 (N_21858,N_21711,N_21728);
nor U21859 (N_21859,N_21782,N_21664);
and U21860 (N_21860,N_21737,N_21632);
and U21861 (N_21861,N_21654,N_21780);
nand U21862 (N_21862,N_21754,N_21779);
xnor U21863 (N_21863,N_21709,N_21656);
nor U21864 (N_21864,N_21697,N_21765);
nand U21865 (N_21865,N_21715,N_21705);
nand U21866 (N_21866,N_21622,N_21631);
nand U21867 (N_21867,N_21710,N_21768);
nand U21868 (N_21868,N_21641,N_21698);
or U21869 (N_21869,N_21727,N_21741);
nor U21870 (N_21870,N_21786,N_21789);
nand U21871 (N_21871,N_21601,N_21723);
xnor U21872 (N_21872,N_21731,N_21630);
or U21873 (N_21873,N_21665,N_21685);
nor U21874 (N_21874,N_21686,N_21660);
nor U21875 (N_21875,N_21701,N_21798);
nor U21876 (N_21876,N_21646,N_21684);
xnor U21877 (N_21877,N_21788,N_21725);
nand U21878 (N_21878,N_21606,N_21702);
or U21879 (N_21879,N_21695,N_21645);
nor U21880 (N_21880,N_21648,N_21750);
and U21881 (N_21881,N_21617,N_21778);
nor U21882 (N_21882,N_21682,N_21770);
and U21883 (N_21883,N_21776,N_21673);
xnor U21884 (N_21884,N_21624,N_21661);
and U21885 (N_21885,N_21726,N_21747);
nand U21886 (N_21886,N_21607,N_21643);
xnor U21887 (N_21887,N_21748,N_21706);
nand U21888 (N_21888,N_21693,N_21713);
nand U21889 (N_21889,N_21677,N_21721);
nor U21890 (N_21890,N_21795,N_21746);
nor U21891 (N_21891,N_21703,N_21793);
or U21892 (N_21892,N_21662,N_21626);
or U21893 (N_21893,N_21769,N_21784);
nand U21894 (N_21894,N_21733,N_21707);
nor U21895 (N_21895,N_21736,N_21658);
and U21896 (N_21896,N_21716,N_21704);
and U21897 (N_21897,N_21620,N_21729);
or U21898 (N_21898,N_21629,N_21611);
and U21899 (N_21899,N_21718,N_21689);
or U21900 (N_21900,N_21742,N_21732);
nor U21901 (N_21901,N_21631,N_21792);
nor U21902 (N_21902,N_21780,N_21656);
or U21903 (N_21903,N_21688,N_21663);
or U21904 (N_21904,N_21664,N_21777);
or U21905 (N_21905,N_21674,N_21616);
or U21906 (N_21906,N_21732,N_21792);
and U21907 (N_21907,N_21746,N_21786);
xor U21908 (N_21908,N_21674,N_21769);
xnor U21909 (N_21909,N_21766,N_21707);
nor U21910 (N_21910,N_21638,N_21635);
nand U21911 (N_21911,N_21622,N_21762);
nor U21912 (N_21912,N_21787,N_21662);
xor U21913 (N_21913,N_21650,N_21742);
nand U21914 (N_21914,N_21668,N_21671);
xor U21915 (N_21915,N_21667,N_21795);
nand U21916 (N_21916,N_21743,N_21727);
and U21917 (N_21917,N_21744,N_21737);
nand U21918 (N_21918,N_21685,N_21698);
xor U21919 (N_21919,N_21787,N_21764);
nand U21920 (N_21920,N_21727,N_21677);
and U21921 (N_21921,N_21733,N_21621);
and U21922 (N_21922,N_21780,N_21742);
or U21923 (N_21923,N_21608,N_21701);
or U21924 (N_21924,N_21641,N_21730);
nand U21925 (N_21925,N_21761,N_21644);
or U21926 (N_21926,N_21680,N_21746);
and U21927 (N_21927,N_21620,N_21652);
nor U21928 (N_21928,N_21647,N_21658);
nor U21929 (N_21929,N_21685,N_21736);
nor U21930 (N_21930,N_21665,N_21758);
nand U21931 (N_21931,N_21765,N_21756);
nor U21932 (N_21932,N_21794,N_21670);
or U21933 (N_21933,N_21798,N_21733);
nand U21934 (N_21934,N_21661,N_21758);
nand U21935 (N_21935,N_21601,N_21638);
xnor U21936 (N_21936,N_21669,N_21695);
or U21937 (N_21937,N_21720,N_21730);
or U21938 (N_21938,N_21783,N_21797);
xnor U21939 (N_21939,N_21726,N_21789);
nor U21940 (N_21940,N_21634,N_21690);
or U21941 (N_21941,N_21683,N_21623);
and U21942 (N_21942,N_21709,N_21620);
nand U21943 (N_21943,N_21760,N_21639);
xnor U21944 (N_21944,N_21772,N_21788);
or U21945 (N_21945,N_21614,N_21694);
nand U21946 (N_21946,N_21607,N_21670);
nor U21947 (N_21947,N_21662,N_21617);
xnor U21948 (N_21948,N_21674,N_21789);
xor U21949 (N_21949,N_21678,N_21737);
nand U21950 (N_21950,N_21669,N_21725);
or U21951 (N_21951,N_21610,N_21663);
or U21952 (N_21952,N_21687,N_21619);
or U21953 (N_21953,N_21662,N_21710);
nand U21954 (N_21954,N_21783,N_21717);
xor U21955 (N_21955,N_21760,N_21797);
and U21956 (N_21956,N_21700,N_21684);
nand U21957 (N_21957,N_21690,N_21669);
nand U21958 (N_21958,N_21600,N_21727);
or U21959 (N_21959,N_21780,N_21729);
nor U21960 (N_21960,N_21776,N_21797);
and U21961 (N_21961,N_21640,N_21655);
or U21962 (N_21962,N_21633,N_21600);
nand U21963 (N_21963,N_21775,N_21718);
and U21964 (N_21964,N_21666,N_21649);
nor U21965 (N_21965,N_21727,N_21606);
xor U21966 (N_21966,N_21799,N_21707);
nand U21967 (N_21967,N_21633,N_21765);
and U21968 (N_21968,N_21689,N_21638);
xnor U21969 (N_21969,N_21720,N_21603);
nand U21970 (N_21970,N_21655,N_21622);
or U21971 (N_21971,N_21782,N_21759);
xor U21972 (N_21972,N_21727,N_21751);
and U21973 (N_21973,N_21740,N_21649);
or U21974 (N_21974,N_21732,N_21756);
and U21975 (N_21975,N_21760,N_21675);
nand U21976 (N_21976,N_21608,N_21698);
nand U21977 (N_21977,N_21791,N_21669);
and U21978 (N_21978,N_21711,N_21616);
and U21979 (N_21979,N_21653,N_21629);
nor U21980 (N_21980,N_21661,N_21785);
and U21981 (N_21981,N_21692,N_21683);
nand U21982 (N_21982,N_21700,N_21731);
or U21983 (N_21983,N_21740,N_21787);
xnor U21984 (N_21984,N_21795,N_21610);
or U21985 (N_21985,N_21744,N_21739);
or U21986 (N_21986,N_21783,N_21612);
xor U21987 (N_21987,N_21654,N_21610);
nor U21988 (N_21988,N_21674,N_21734);
and U21989 (N_21989,N_21618,N_21725);
and U21990 (N_21990,N_21771,N_21635);
nor U21991 (N_21991,N_21719,N_21710);
nand U21992 (N_21992,N_21627,N_21748);
nand U21993 (N_21993,N_21737,N_21714);
nand U21994 (N_21994,N_21747,N_21727);
nor U21995 (N_21995,N_21780,N_21796);
xnor U21996 (N_21996,N_21618,N_21720);
nor U21997 (N_21997,N_21754,N_21656);
or U21998 (N_21998,N_21722,N_21750);
and U21999 (N_21999,N_21606,N_21751);
or U22000 (N_22000,N_21947,N_21943);
nand U22001 (N_22001,N_21824,N_21832);
xor U22002 (N_22002,N_21816,N_21940);
xor U22003 (N_22003,N_21804,N_21830);
or U22004 (N_22004,N_21931,N_21838);
nand U22005 (N_22005,N_21886,N_21911);
xnor U22006 (N_22006,N_21957,N_21989);
nand U22007 (N_22007,N_21892,N_21977);
and U22008 (N_22008,N_21800,N_21981);
nand U22009 (N_22009,N_21811,N_21949);
or U22010 (N_22010,N_21803,N_21910);
or U22011 (N_22011,N_21983,N_21999);
xor U22012 (N_22012,N_21859,N_21982);
xor U22013 (N_22013,N_21987,N_21965);
xor U22014 (N_22014,N_21812,N_21821);
xor U22015 (N_22015,N_21845,N_21935);
and U22016 (N_22016,N_21878,N_21835);
xnor U22017 (N_22017,N_21933,N_21847);
and U22018 (N_22018,N_21921,N_21958);
nor U22019 (N_22019,N_21915,N_21819);
nor U22020 (N_22020,N_21988,N_21902);
xnor U22021 (N_22021,N_21936,N_21869);
nor U22022 (N_22022,N_21844,N_21946);
nor U22023 (N_22023,N_21896,N_21927);
nor U22024 (N_22024,N_21833,N_21818);
xnor U22025 (N_22025,N_21950,N_21928);
nand U22026 (N_22026,N_21840,N_21926);
and U22027 (N_22027,N_21961,N_21836);
nand U22028 (N_22028,N_21937,N_21942);
nor U22029 (N_22029,N_21850,N_21805);
and U22030 (N_22030,N_21891,N_21817);
nand U22031 (N_22031,N_21848,N_21909);
nand U22032 (N_22032,N_21953,N_21938);
or U22033 (N_22033,N_21898,N_21901);
nand U22034 (N_22034,N_21806,N_21932);
and U22035 (N_22035,N_21808,N_21994);
nor U22036 (N_22036,N_21908,N_21913);
nand U22037 (N_22037,N_21841,N_21876);
xnor U22038 (N_22038,N_21956,N_21975);
nor U22039 (N_22039,N_21858,N_21944);
nand U22040 (N_22040,N_21941,N_21846);
nand U22041 (N_22041,N_21864,N_21925);
nor U22042 (N_22042,N_21951,N_21813);
and U22043 (N_22043,N_21882,N_21801);
or U22044 (N_22044,N_21861,N_21923);
nand U22045 (N_22045,N_21877,N_21873);
or U22046 (N_22046,N_21952,N_21964);
nor U22047 (N_22047,N_21826,N_21945);
nor U22048 (N_22048,N_21885,N_21920);
or U22049 (N_22049,N_21829,N_21810);
xnor U22050 (N_22050,N_21972,N_21979);
xor U22051 (N_22051,N_21969,N_21916);
nor U22052 (N_22052,N_21906,N_21971);
xnor U22053 (N_22053,N_21860,N_21894);
and U22054 (N_22054,N_21871,N_21867);
nor U22055 (N_22055,N_21884,N_21856);
nand U22056 (N_22056,N_21880,N_21863);
or U22057 (N_22057,N_21831,N_21966);
and U22058 (N_22058,N_21888,N_21984);
or U22059 (N_22059,N_21889,N_21967);
xor U22060 (N_22060,N_21874,N_21897);
xor U22061 (N_22061,N_21934,N_21973);
xor U22062 (N_22062,N_21960,N_21990);
nor U22063 (N_22063,N_21955,N_21842);
xnor U22064 (N_22064,N_21907,N_21929);
nand U22065 (N_22065,N_21822,N_21959);
nor U22066 (N_22066,N_21839,N_21852);
or U22067 (N_22067,N_21881,N_21922);
or U22068 (N_22068,N_21980,N_21887);
or U22069 (N_22069,N_21954,N_21974);
xnor U22070 (N_22070,N_21998,N_21924);
and U22071 (N_22071,N_21904,N_21828);
nand U22072 (N_22072,N_21823,N_21963);
or U22073 (N_22073,N_21995,N_21978);
and U22074 (N_22074,N_21948,N_21890);
xnor U22075 (N_22075,N_21837,N_21993);
or U22076 (N_22076,N_21872,N_21814);
and U22077 (N_22077,N_21807,N_21883);
xor U22078 (N_22078,N_21985,N_21996);
xnor U22079 (N_22079,N_21855,N_21893);
xnor U22080 (N_22080,N_21968,N_21970);
nand U22081 (N_22081,N_21976,N_21912);
nor U22082 (N_22082,N_21930,N_21851);
nor U22083 (N_22083,N_21802,N_21905);
xor U22084 (N_22084,N_21986,N_21809);
or U22085 (N_22085,N_21815,N_21939);
or U22086 (N_22086,N_21919,N_21857);
nand U22087 (N_22087,N_21875,N_21903);
and U22088 (N_22088,N_21820,N_21917);
or U22089 (N_22089,N_21865,N_21827);
nor U22090 (N_22090,N_21991,N_21997);
nor U22091 (N_22091,N_21962,N_21868);
or U22092 (N_22092,N_21899,N_21918);
xnor U22093 (N_22093,N_21870,N_21914);
nand U22094 (N_22094,N_21895,N_21900);
nor U22095 (N_22095,N_21849,N_21866);
or U22096 (N_22096,N_21992,N_21834);
and U22097 (N_22097,N_21862,N_21843);
nand U22098 (N_22098,N_21879,N_21854);
nand U22099 (N_22099,N_21853,N_21825);
xnor U22100 (N_22100,N_21885,N_21990);
or U22101 (N_22101,N_21982,N_21920);
xor U22102 (N_22102,N_21845,N_21934);
or U22103 (N_22103,N_21954,N_21934);
and U22104 (N_22104,N_21852,N_21892);
or U22105 (N_22105,N_21891,N_21877);
and U22106 (N_22106,N_21873,N_21847);
nor U22107 (N_22107,N_21983,N_21941);
nand U22108 (N_22108,N_21826,N_21806);
xnor U22109 (N_22109,N_21860,N_21819);
nand U22110 (N_22110,N_21864,N_21886);
xor U22111 (N_22111,N_21921,N_21936);
nand U22112 (N_22112,N_21856,N_21855);
nand U22113 (N_22113,N_21941,N_21935);
nand U22114 (N_22114,N_21955,N_21855);
nor U22115 (N_22115,N_21922,N_21939);
and U22116 (N_22116,N_21836,N_21889);
and U22117 (N_22117,N_21859,N_21867);
nand U22118 (N_22118,N_21981,N_21851);
and U22119 (N_22119,N_21921,N_21866);
nand U22120 (N_22120,N_21811,N_21894);
or U22121 (N_22121,N_21847,N_21913);
xnor U22122 (N_22122,N_21900,N_21825);
xor U22123 (N_22123,N_21809,N_21803);
nand U22124 (N_22124,N_21890,N_21995);
nor U22125 (N_22125,N_21923,N_21849);
xor U22126 (N_22126,N_21904,N_21932);
and U22127 (N_22127,N_21815,N_21965);
nand U22128 (N_22128,N_21832,N_21837);
nand U22129 (N_22129,N_21831,N_21990);
xor U22130 (N_22130,N_21824,N_21882);
nor U22131 (N_22131,N_21935,N_21947);
xor U22132 (N_22132,N_21987,N_21938);
or U22133 (N_22133,N_21839,N_21886);
xor U22134 (N_22134,N_21866,N_21868);
and U22135 (N_22135,N_21982,N_21838);
nand U22136 (N_22136,N_21800,N_21995);
and U22137 (N_22137,N_21910,N_21854);
xnor U22138 (N_22138,N_21884,N_21979);
and U22139 (N_22139,N_21875,N_21915);
or U22140 (N_22140,N_21893,N_21962);
nor U22141 (N_22141,N_21946,N_21918);
nor U22142 (N_22142,N_21801,N_21812);
nand U22143 (N_22143,N_21845,N_21932);
or U22144 (N_22144,N_21905,N_21909);
xor U22145 (N_22145,N_21994,N_21845);
nor U22146 (N_22146,N_21886,N_21804);
or U22147 (N_22147,N_21907,N_21988);
or U22148 (N_22148,N_21913,N_21969);
nor U22149 (N_22149,N_21899,N_21942);
nand U22150 (N_22150,N_21837,N_21800);
nor U22151 (N_22151,N_21801,N_21804);
and U22152 (N_22152,N_21913,N_21924);
and U22153 (N_22153,N_21996,N_21987);
xnor U22154 (N_22154,N_21839,N_21851);
and U22155 (N_22155,N_21945,N_21845);
xor U22156 (N_22156,N_21803,N_21802);
nor U22157 (N_22157,N_21814,N_21801);
and U22158 (N_22158,N_21985,N_21839);
xor U22159 (N_22159,N_21890,N_21805);
and U22160 (N_22160,N_21870,N_21826);
xnor U22161 (N_22161,N_21896,N_21809);
or U22162 (N_22162,N_21883,N_21996);
nand U22163 (N_22163,N_21852,N_21936);
or U22164 (N_22164,N_21830,N_21822);
xor U22165 (N_22165,N_21975,N_21835);
or U22166 (N_22166,N_21952,N_21836);
nand U22167 (N_22167,N_21909,N_21899);
xor U22168 (N_22168,N_21804,N_21858);
and U22169 (N_22169,N_21917,N_21972);
nor U22170 (N_22170,N_21900,N_21995);
nor U22171 (N_22171,N_21911,N_21919);
nor U22172 (N_22172,N_21841,N_21933);
nand U22173 (N_22173,N_21866,N_21896);
nand U22174 (N_22174,N_21963,N_21958);
and U22175 (N_22175,N_21870,N_21921);
or U22176 (N_22176,N_21808,N_21805);
xnor U22177 (N_22177,N_21816,N_21915);
nand U22178 (N_22178,N_21986,N_21816);
or U22179 (N_22179,N_21833,N_21920);
xnor U22180 (N_22180,N_21808,N_21885);
nand U22181 (N_22181,N_21812,N_21986);
nand U22182 (N_22182,N_21821,N_21838);
nor U22183 (N_22183,N_21819,N_21974);
or U22184 (N_22184,N_21907,N_21919);
nor U22185 (N_22185,N_21837,N_21848);
nand U22186 (N_22186,N_21818,N_21884);
or U22187 (N_22187,N_21942,N_21806);
and U22188 (N_22188,N_21961,N_21828);
nand U22189 (N_22189,N_21997,N_21895);
or U22190 (N_22190,N_21953,N_21896);
nor U22191 (N_22191,N_21841,N_21925);
xnor U22192 (N_22192,N_21975,N_21912);
nor U22193 (N_22193,N_21864,N_21842);
or U22194 (N_22194,N_21985,N_21906);
nor U22195 (N_22195,N_21812,N_21803);
or U22196 (N_22196,N_21889,N_21876);
or U22197 (N_22197,N_21941,N_21866);
xor U22198 (N_22198,N_21835,N_21890);
nand U22199 (N_22199,N_21864,N_21803);
nand U22200 (N_22200,N_22184,N_22121);
or U22201 (N_22201,N_22165,N_22152);
nor U22202 (N_22202,N_22197,N_22007);
or U22203 (N_22203,N_22014,N_22168);
and U22204 (N_22204,N_22053,N_22067);
nor U22205 (N_22205,N_22015,N_22162);
or U22206 (N_22206,N_22179,N_22084);
nand U22207 (N_22207,N_22194,N_22122);
or U22208 (N_22208,N_22086,N_22127);
xnor U22209 (N_22209,N_22113,N_22029);
nor U22210 (N_22210,N_22042,N_22140);
xor U22211 (N_22211,N_22006,N_22104);
xor U22212 (N_22212,N_22188,N_22022);
nor U22213 (N_22213,N_22148,N_22021);
nor U22214 (N_22214,N_22112,N_22093);
nand U22215 (N_22215,N_22091,N_22125);
and U22216 (N_22216,N_22128,N_22085);
nor U22217 (N_22217,N_22008,N_22002);
or U22218 (N_22218,N_22126,N_22024);
or U22219 (N_22219,N_22176,N_22108);
and U22220 (N_22220,N_22100,N_22186);
nand U22221 (N_22221,N_22039,N_22132);
xor U22222 (N_22222,N_22060,N_22033);
and U22223 (N_22223,N_22041,N_22163);
nand U22224 (N_22224,N_22123,N_22096);
and U22225 (N_22225,N_22032,N_22065);
nand U22226 (N_22226,N_22134,N_22105);
nand U22227 (N_22227,N_22023,N_22054);
or U22228 (N_22228,N_22063,N_22185);
or U22229 (N_22229,N_22069,N_22156);
nor U22230 (N_22230,N_22017,N_22097);
xor U22231 (N_22231,N_22145,N_22079);
nand U22232 (N_22232,N_22161,N_22103);
or U22233 (N_22233,N_22057,N_22115);
nor U22234 (N_22234,N_22013,N_22001);
xnor U22235 (N_22235,N_22130,N_22195);
xor U22236 (N_22236,N_22048,N_22052);
nand U22237 (N_22237,N_22199,N_22011);
and U22238 (N_22238,N_22026,N_22173);
or U22239 (N_22239,N_22095,N_22167);
or U22240 (N_22240,N_22004,N_22154);
nor U22241 (N_22241,N_22030,N_22120);
or U22242 (N_22242,N_22019,N_22193);
nor U22243 (N_22243,N_22102,N_22119);
nor U22244 (N_22244,N_22070,N_22092);
or U22245 (N_22245,N_22150,N_22110);
xnor U22246 (N_22246,N_22071,N_22078);
xor U22247 (N_22247,N_22009,N_22137);
nor U22248 (N_22248,N_22056,N_22076);
or U22249 (N_22249,N_22175,N_22083);
or U22250 (N_22250,N_22050,N_22038);
or U22251 (N_22251,N_22062,N_22135);
nand U22252 (N_22252,N_22081,N_22020);
xnor U22253 (N_22253,N_22045,N_22068);
nor U22254 (N_22254,N_22025,N_22046);
nand U22255 (N_22255,N_22090,N_22101);
nor U22256 (N_22256,N_22158,N_22133);
nand U22257 (N_22257,N_22143,N_22170);
and U22258 (N_22258,N_22171,N_22088);
xnor U22259 (N_22259,N_22149,N_22160);
or U22260 (N_22260,N_22178,N_22016);
nand U22261 (N_22261,N_22166,N_22099);
or U22262 (N_22262,N_22155,N_22000);
nor U22263 (N_22263,N_22124,N_22172);
and U22264 (N_22264,N_22077,N_22035);
nand U22265 (N_22265,N_22191,N_22182);
nand U22266 (N_22266,N_22159,N_22040);
xnor U22267 (N_22267,N_22144,N_22141);
and U22268 (N_22268,N_22037,N_22051);
xor U22269 (N_22269,N_22131,N_22157);
and U22270 (N_22270,N_22198,N_22177);
or U22271 (N_22271,N_22073,N_22018);
nand U22272 (N_22272,N_22146,N_22036);
nor U22273 (N_22273,N_22082,N_22196);
or U22274 (N_22274,N_22044,N_22005);
xnor U22275 (N_22275,N_22012,N_22003);
or U22276 (N_22276,N_22055,N_22080);
or U22277 (N_22277,N_22129,N_22010);
nor U22278 (N_22278,N_22031,N_22138);
nand U22279 (N_22279,N_22181,N_22075);
and U22280 (N_22280,N_22049,N_22066);
nor U22281 (N_22281,N_22072,N_22190);
xnor U22282 (N_22282,N_22058,N_22189);
xor U22283 (N_22283,N_22169,N_22117);
nand U22284 (N_22284,N_22142,N_22074);
and U22285 (N_22285,N_22192,N_22187);
or U22286 (N_22286,N_22139,N_22027);
nand U22287 (N_22287,N_22153,N_22047);
xor U22288 (N_22288,N_22147,N_22109);
nor U22289 (N_22289,N_22028,N_22151);
or U22290 (N_22290,N_22034,N_22116);
or U22291 (N_22291,N_22136,N_22064);
xnor U22292 (N_22292,N_22043,N_22164);
xnor U22293 (N_22293,N_22087,N_22114);
and U22294 (N_22294,N_22059,N_22180);
xnor U22295 (N_22295,N_22118,N_22107);
and U22296 (N_22296,N_22106,N_22061);
and U22297 (N_22297,N_22174,N_22183);
nand U22298 (N_22298,N_22111,N_22089);
xnor U22299 (N_22299,N_22098,N_22094);
and U22300 (N_22300,N_22031,N_22038);
or U22301 (N_22301,N_22046,N_22067);
or U22302 (N_22302,N_22120,N_22036);
and U22303 (N_22303,N_22080,N_22034);
nand U22304 (N_22304,N_22069,N_22178);
or U22305 (N_22305,N_22078,N_22018);
nor U22306 (N_22306,N_22047,N_22003);
and U22307 (N_22307,N_22124,N_22151);
xnor U22308 (N_22308,N_22182,N_22072);
and U22309 (N_22309,N_22178,N_22145);
and U22310 (N_22310,N_22097,N_22199);
nor U22311 (N_22311,N_22089,N_22025);
and U22312 (N_22312,N_22066,N_22080);
nand U22313 (N_22313,N_22175,N_22052);
nor U22314 (N_22314,N_22080,N_22120);
nand U22315 (N_22315,N_22076,N_22080);
or U22316 (N_22316,N_22134,N_22167);
nand U22317 (N_22317,N_22123,N_22159);
or U22318 (N_22318,N_22072,N_22103);
nand U22319 (N_22319,N_22113,N_22041);
nand U22320 (N_22320,N_22103,N_22159);
nor U22321 (N_22321,N_22092,N_22083);
nor U22322 (N_22322,N_22019,N_22163);
nor U22323 (N_22323,N_22006,N_22109);
or U22324 (N_22324,N_22077,N_22126);
and U22325 (N_22325,N_22084,N_22068);
xor U22326 (N_22326,N_22193,N_22047);
or U22327 (N_22327,N_22019,N_22104);
nand U22328 (N_22328,N_22135,N_22021);
nand U22329 (N_22329,N_22140,N_22011);
or U22330 (N_22330,N_22175,N_22192);
nand U22331 (N_22331,N_22176,N_22097);
nor U22332 (N_22332,N_22172,N_22159);
or U22333 (N_22333,N_22143,N_22168);
nand U22334 (N_22334,N_22175,N_22190);
nand U22335 (N_22335,N_22078,N_22041);
or U22336 (N_22336,N_22147,N_22115);
nand U22337 (N_22337,N_22015,N_22053);
xnor U22338 (N_22338,N_22170,N_22180);
nand U22339 (N_22339,N_22126,N_22134);
or U22340 (N_22340,N_22177,N_22110);
xnor U22341 (N_22341,N_22120,N_22044);
and U22342 (N_22342,N_22080,N_22033);
nand U22343 (N_22343,N_22192,N_22137);
nand U22344 (N_22344,N_22042,N_22037);
and U22345 (N_22345,N_22069,N_22028);
and U22346 (N_22346,N_22101,N_22117);
or U22347 (N_22347,N_22061,N_22139);
or U22348 (N_22348,N_22165,N_22138);
xor U22349 (N_22349,N_22116,N_22168);
nand U22350 (N_22350,N_22057,N_22130);
xnor U22351 (N_22351,N_22059,N_22124);
xor U22352 (N_22352,N_22061,N_22123);
nand U22353 (N_22353,N_22028,N_22008);
nand U22354 (N_22354,N_22169,N_22127);
nor U22355 (N_22355,N_22112,N_22168);
nand U22356 (N_22356,N_22068,N_22035);
xor U22357 (N_22357,N_22193,N_22132);
or U22358 (N_22358,N_22126,N_22130);
nor U22359 (N_22359,N_22114,N_22069);
or U22360 (N_22360,N_22019,N_22102);
xor U22361 (N_22361,N_22117,N_22073);
nand U22362 (N_22362,N_22041,N_22016);
xnor U22363 (N_22363,N_22123,N_22104);
nand U22364 (N_22364,N_22092,N_22062);
or U22365 (N_22365,N_22096,N_22074);
or U22366 (N_22366,N_22115,N_22042);
xor U22367 (N_22367,N_22108,N_22180);
nand U22368 (N_22368,N_22112,N_22068);
and U22369 (N_22369,N_22132,N_22027);
and U22370 (N_22370,N_22161,N_22157);
or U22371 (N_22371,N_22107,N_22160);
and U22372 (N_22372,N_22138,N_22030);
or U22373 (N_22373,N_22076,N_22178);
xnor U22374 (N_22374,N_22097,N_22121);
or U22375 (N_22375,N_22120,N_22049);
xor U22376 (N_22376,N_22191,N_22198);
nor U22377 (N_22377,N_22197,N_22098);
and U22378 (N_22378,N_22053,N_22176);
nor U22379 (N_22379,N_22082,N_22060);
nand U22380 (N_22380,N_22161,N_22069);
nor U22381 (N_22381,N_22045,N_22165);
nand U22382 (N_22382,N_22182,N_22050);
or U22383 (N_22383,N_22166,N_22138);
nor U22384 (N_22384,N_22000,N_22083);
or U22385 (N_22385,N_22128,N_22050);
nor U22386 (N_22386,N_22172,N_22049);
nor U22387 (N_22387,N_22180,N_22177);
or U22388 (N_22388,N_22023,N_22062);
or U22389 (N_22389,N_22085,N_22193);
nand U22390 (N_22390,N_22096,N_22000);
nor U22391 (N_22391,N_22150,N_22158);
xor U22392 (N_22392,N_22017,N_22079);
nor U22393 (N_22393,N_22167,N_22112);
xor U22394 (N_22394,N_22173,N_22191);
or U22395 (N_22395,N_22154,N_22069);
xor U22396 (N_22396,N_22036,N_22016);
or U22397 (N_22397,N_22146,N_22144);
and U22398 (N_22398,N_22128,N_22095);
nand U22399 (N_22399,N_22093,N_22151);
xnor U22400 (N_22400,N_22226,N_22273);
nand U22401 (N_22401,N_22380,N_22271);
and U22402 (N_22402,N_22312,N_22229);
and U22403 (N_22403,N_22336,N_22393);
xnor U22404 (N_22404,N_22359,N_22227);
xnor U22405 (N_22405,N_22364,N_22213);
nand U22406 (N_22406,N_22201,N_22315);
nand U22407 (N_22407,N_22398,N_22269);
xnor U22408 (N_22408,N_22339,N_22261);
or U22409 (N_22409,N_22371,N_22238);
or U22410 (N_22410,N_22381,N_22333);
and U22411 (N_22411,N_22251,N_22275);
or U22412 (N_22412,N_22215,N_22375);
xnor U22413 (N_22413,N_22242,N_22321);
xnor U22414 (N_22414,N_22262,N_22386);
xor U22415 (N_22415,N_22248,N_22383);
nand U22416 (N_22416,N_22302,N_22326);
xnor U22417 (N_22417,N_22303,N_22353);
and U22418 (N_22418,N_22214,N_22350);
or U22419 (N_22419,N_22284,N_22361);
or U22420 (N_22420,N_22255,N_22246);
or U22421 (N_22421,N_22205,N_22268);
nand U22422 (N_22422,N_22338,N_22372);
xnor U22423 (N_22423,N_22320,N_22387);
xor U22424 (N_22424,N_22200,N_22349);
or U22425 (N_22425,N_22343,N_22210);
or U22426 (N_22426,N_22222,N_22342);
or U22427 (N_22427,N_22347,N_22344);
or U22428 (N_22428,N_22270,N_22234);
nor U22429 (N_22429,N_22239,N_22236);
or U22430 (N_22430,N_22216,N_22392);
xor U22431 (N_22431,N_22310,N_22305);
and U22432 (N_22432,N_22249,N_22385);
or U22433 (N_22433,N_22357,N_22265);
xor U22434 (N_22434,N_22294,N_22382);
and U22435 (N_22435,N_22340,N_22292);
or U22436 (N_22436,N_22328,N_22219);
nand U22437 (N_22437,N_22396,N_22301);
and U22438 (N_22438,N_22244,N_22289);
nor U22439 (N_22439,N_22224,N_22272);
nand U22440 (N_22440,N_22352,N_22264);
and U22441 (N_22441,N_22241,N_22212);
and U22442 (N_22442,N_22220,N_22299);
nor U22443 (N_22443,N_22274,N_22278);
xor U22444 (N_22444,N_22287,N_22388);
and U22445 (N_22445,N_22324,N_22280);
and U22446 (N_22446,N_22247,N_22360);
and U22447 (N_22447,N_22285,N_22293);
and U22448 (N_22448,N_22308,N_22311);
or U22449 (N_22449,N_22317,N_22369);
nand U22450 (N_22450,N_22276,N_22304);
and U22451 (N_22451,N_22290,N_22218);
and U22452 (N_22452,N_22363,N_22313);
nand U22453 (N_22453,N_22346,N_22245);
or U22454 (N_22454,N_22228,N_22348);
nand U22455 (N_22455,N_22243,N_22399);
and U22456 (N_22456,N_22252,N_22327);
and U22457 (N_22457,N_22331,N_22377);
xor U22458 (N_22458,N_22300,N_22230);
and U22459 (N_22459,N_22306,N_22281);
or U22460 (N_22460,N_22345,N_22354);
nor U22461 (N_22461,N_22221,N_22291);
xnor U22462 (N_22462,N_22233,N_22368);
xnor U22463 (N_22463,N_22297,N_22329);
xor U22464 (N_22464,N_22267,N_22250);
or U22465 (N_22465,N_22325,N_22266);
or U22466 (N_22466,N_22235,N_22254);
and U22467 (N_22467,N_22330,N_22295);
and U22468 (N_22468,N_22394,N_22322);
nor U22469 (N_22469,N_22365,N_22367);
nand U22470 (N_22470,N_22288,N_22370);
nor U22471 (N_22471,N_22277,N_22207);
or U22472 (N_22472,N_22356,N_22296);
xnor U22473 (N_22473,N_22217,N_22257);
or U22474 (N_22474,N_22378,N_22323);
xnor U22475 (N_22475,N_22366,N_22223);
nor U22476 (N_22476,N_22351,N_22314);
xor U22477 (N_22477,N_22253,N_22390);
xor U22478 (N_22478,N_22358,N_22231);
nand U22479 (N_22479,N_22211,N_22286);
nand U22480 (N_22480,N_22355,N_22208);
or U22481 (N_22481,N_22332,N_22373);
and U22482 (N_22482,N_22391,N_22202);
nor U22483 (N_22483,N_22283,N_22384);
nand U22484 (N_22484,N_22376,N_22309);
and U22485 (N_22485,N_22379,N_22225);
and U22486 (N_22486,N_22362,N_22318);
and U22487 (N_22487,N_22307,N_22259);
nand U22488 (N_22488,N_22256,N_22334);
nor U22489 (N_22489,N_22335,N_22206);
nor U22490 (N_22490,N_22374,N_22341);
xor U22491 (N_22491,N_22232,N_22237);
or U22492 (N_22492,N_22240,N_22395);
nor U22493 (N_22493,N_22298,N_22319);
xnor U22494 (N_22494,N_22316,N_22260);
nand U22495 (N_22495,N_22203,N_22209);
nor U22496 (N_22496,N_22282,N_22204);
and U22497 (N_22497,N_22389,N_22397);
nand U22498 (N_22498,N_22258,N_22279);
nor U22499 (N_22499,N_22337,N_22263);
xnor U22500 (N_22500,N_22291,N_22255);
and U22501 (N_22501,N_22391,N_22302);
and U22502 (N_22502,N_22320,N_22318);
nor U22503 (N_22503,N_22359,N_22332);
or U22504 (N_22504,N_22264,N_22261);
and U22505 (N_22505,N_22309,N_22255);
nand U22506 (N_22506,N_22340,N_22309);
xnor U22507 (N_22507,N_22258,N_22223);
and U22508 (N_22508,N_22384,N_22274);
and U22509 (N_22509,N_22372,N_22238);
and U22510 (N_22510,N_22279,N_22200);
xnor U22511 (N_22511,N_22306,N_22297);
nand U22512 (N_22512,N_22272,N_22255);
nor U22513 (N_22513,N_22258,N_22206);
nand U22514 (N_22514,N_22388,N_22259);
nor U22515 (N_22515,N_22224,N_22241);
nand U22516 (N_22516,N_22324,N_22349);
nor U22517 (N_22517,N_22248,N_22341);
or U22518 (N_22518,N_22268,N_22267);
nand U22519 (N_22519,N_22327,N_22341);
nor U22520 (N_22520,N_22376,N_22275);
or U22521 (N_22521,N_22331,N_22210);
nor U22522 (N_22522,N_22354,N_22235);
and U22523 (N_22523,N_22333,N_22390);
xor U22524 (N_22524,N_22274,N_22202);
xor U22525 (N_22525,N_22201,N_22289);
or U22526 (N_22526,N_22201,N_22374);
nand U22527 (N_22527,N_22239,N_22351);
nand U22528 (N_22528,N_22341,N_22202);
xor U22529 (N_22529,N_22250,N_22380);
xor U22530 (N_22530,N_22278,N_22225);
nand U22531 (N_22531,N_22360,N_22396);
nand U22532 (N_22532,N_22346,N_22283);
or U22533 (N_22533,N_22266,N_22267);
or U22534 (N_22534,N_22236,N_22354);
and U22535 (N_22535,N_22367,N_22338);
and U22536 (N_22536,N_22281,N_22254);
xor U22537 (N_22537,N_22397,N_22347);
nor U22538 (N_22538,N_22330,N_22259);
xor U22539 (N_22539,N_22298,N_22367);
or U22540 (N_22540,N_22348,N_22220);
xor U22541 (N_22541,N_22247,N_22272);
nor U22542 (N_22542,N_22265,N_22260);
or U22543 (N_22543,N_22342,N_22210);
nand U22544 (N_22544,N_22360,N_22386);
nand U22545 (N_22545,N_22293,N_22214);
nor U22546 (N_22546,N_22311,N_22313);
and U22547 (N_22547,N_22228,N_22302);
and U22548 (N_22548,N_22252,N_22251);
nand U22549 (N_22549,N_22311,N_22345);
or U22550 (N_22550,N_22270,N_22238);
xnor U22551 (N_22551,N_22218,N_22211);
or U22552 (N_22552,N_22287,N_22248);
or U22553 (N_22553,N_22251,N_22201);
or U22554 (N_22554,N_22346,N_22291);
and U22555 (N_22555,N_22200,N_22328);
nand U22556 (N_22556,N_22371,N_22320);
or U22557 (N_22557,N_22315,N_22297);
or U22558 (N_22558,N_22254,N_22237);
or U22559 (N_22559,N_22222,N_22299);
nand U22560 (N_22560,N_22313,N_22319);
xor U22561 (N_22561,N_22382,N_22299);
xnor U22562 (N_22562,N_22365,N_22300);
nor U22563 (N_22563,N_22209,N_22292);
or U22564 (N_22564,N_22332,N_22253);
nor U22565 (N_22565,N_22211,N_22358);
and U22566 (N_22566,N_22295,N_22347);
xnor U22567 (N_22567,N_22352,N_22231);
or U22568 (N_22568,N_22353,N_22252);
xnor U22569 (N_22569,N_22244,N_22397);
nand U22570 (N_22570,N_22358,N_22345);
nand U22571 (N_22571,N_22239,N_22278);
nor U22572 (N_22572,N_22229,N_22357);
nand U22573 (N_22573,N_22210,N_22361);
xnor U22574 (N_22574,N_22242,N_22341);
xor U22575 (N_22575,N_22373,N_22256);
and U22576 (N_22576,N_22221,N_22264);
nand U22577 (N_22577,N_22280,N_22238);
xor U22578 (N_22578,N_22356,N_22312);
nor U22579 (N_22579,N_22215,N_22388);
or U22580 (N_22580,N_22327,N_22305);
nor U22581 (N_22581,N_22230,N_22352);
and U22582 (N_22582,N_22262,N_22348);
nand U22583 (N_22583,N_22239,N_22363);
nor U22584 (N_22584,N_22386,N_22246);
nor U22585 (N_22585,N_22268,N_22311);
and U22586 (N_22586,N_22231,N_22378);
and U22587 (N_22587,N_22359,N_22204);
xor U22588 (N_22588,N_22291,N_22309);
or U22589 (N_22589,N_22274,N_22345);
nor U22590 (N_22590,N_22337,N_22230);
and U22591 (N_22591,N_22309,N_22293);
and U22592 (N_22592,N_22385,N_22319);
or U22593 (N_22593,N_22225,N_22366);
and U22594 (N_22594,N_22208,N_22267);
or U22595 (N_22595,N_22245,N_22310);
nor U22596 (N_22596,N_22328,N_22238);
xnor U22597 (N_22597,N_22289,N_22372);
nand U22598 (N_22598,N_22216,N_22205);
and U22599 (N_22599,N_22271,N_22384);
and U22600 (N_22600,N_22581,N_22431);
or U22601 (N_22601,N_22489,N_22514);
nand U22602 (N_22602,N_22418,N_22504);
nor U22603 (N_22603,N_22521,N_22511);
and U22604 (N_22604,N_22530,N_22410);
or U22605 (N_22605,N_22500,N_22553);
nor U22606 (N_22606,N_22474,N_22417);
nor U22607 (N_22607,N_22580,N_22437);
nor U22608 (N_22608,N_22536,N_22493);
and U22609 (N_22609,N_22481,N_22430);
xor U22610 (N_22610,N_22546,N_22549);
nor U22611 (N_22611,N_22448,N_22557);
and U22612 (N_22612,N_22591,N_22475);
xnor U22613 (N_22613,N_22544,N_22455);
nand U22614 (N_22614,N_22473,N_22406);
nand U22615 (N_22615,N_22534,N_22477);
nor U22616 (N_22616,N_22458,N_22421);
and U22617 (N_22617,N_22495,N_22434);
xnor U22618 (N_22618,N_22563,N_22450);
nand U22619 (N_22619,N_22586,N_22401);
nor U22620 (N_22620,N_22497,N_22569);
nor U22621 (N_22621,N_22415,N_22433);
xor U22622 (N_22622,N_22516,N_22505);
xnor U22623 (N_22623,N_22496,N_22540);
or U22624 (N_22624,N_22484,N_22507);
and U22625 (N_22625,N_22574,N_22427);
nand U22626 (N_22626,N_22508,N_22598);
nor U22627 (N_22627,N_22487,N_22518);
xor U22628 (N_22628,N_22400,N_22411);
nor U22629 (N_22629,N_22560,N_22593);
and U22630 (N_22630,N_22567,N_22552);
xor U22631 (N_22631,N_22550,N_22439);
nor U22632 (N_22632,N_22525,N_22463);
or U22633 (N_22633,N_22583,N_22568);
nand U22634 (N_22634,N_22443,N_22470);
xor U22635 (N_22635,N_22498,N_22419);
nand U22636 (N_22636,N_22412,N_22528);
nor U22637 (N_22637,N_22403,N_22526);
nor U22638 (N_22638,N_22482,N_22539);
nor U22639 (N_22639,N_22579,N_22467);
and U22640 (N_22640,N_22457,N_22499);
nor U22641 (N_22641,N_22587,N_22423);
and U22642 (N_22642,N_22416,N_22420);
nor U22643 (N_22643,N_22413,N_22483);
nand U22644 (N_22644,N_22545,N_22543);
xnor U22645 (N_22645,N_22466,N_22519);
xor U22646 (N_22646,N_22527,N_22541);
or U22647 (N_22647,N_22537,N_22509);
nor U22648 (N_22648,N_22575,N_22566);
nor U22649 (N_22649,N_22438,N_22436);
and U22650 (N_22650,N_22594,N_22452);
nor U22651 (N_22651,N_22456,N_22488);
nand U22652 (N_22652,N_22513,N_22572);
xor U22653 (N_22653,N_22460,N_22565);
and U22654 (N_22654,N_22409,N_22429);
nand U22655 (N_22655,N_22564,N_22590);
xnor U22656 (N_22656,N_22465,N_22551);
nor U22657 (N_22657,N_22554,N_22480);
nand U22658 (N_22658,N_22555,N_22445);
xor U22659 (N_22659,N_22556,N_22512);
nor U22660 (N_22660,N_22548,N_22503);
or U22661 (N_22661,N_22506,N_22428);
and U22662 (N_22662,N_22589,N_22592);
and U22663 (N_22663,N_22405,N_22449);
and U22664 (N_22664,N_22490,N_22464);
and U22665 (N_22665,N_22462,N_22529);
and U22666 (N_22666,N_22432,N_22542);
xor U22667 (N_22667,N_22559,N_22441);
nor U22668 (N_22668,N_22478,N_22578);
nor U22669 (N_22669,N_22533,N_22585);
and U22670 (N_22670,N_22453,N_22494);
nor U22671 (N_22671,N_22435,N_22576);
xor U22672 (N_22672,N_22468,N_22531);
or U22673 (N_22673,N_22520,N_22524);
or U22674 (N_22674,N_22486,N_22532);
xnor U22675 (N_22675,N_22502,N_22454);
and U22676 (N_22676,N_22588,N_22561);
or U22677 (N_22677,N_22407,N_22510);
nand U22678 (N_22678,N_22426,N_22461);
and U22679 (N_22679,N_22476,N_22491);
nand U22680 (N_22680,N_22547,N_22492);
and U22681 (N_22681,N_22562,N_22523);
xnor U22682 (N_22682,N_22408,N_22517);
or U22683 (N_22683,N_22597,N_22515);
nor U22684 (N_22684,N_22571,N_22599);
nor U22685 (N_22685,N_22471,N_22573);
and U22686 (N_22686,N_22425,N_22442);
or U22687 (N_22687,N_22485,N_22522);
xor U22688 (N_22688,N_22440,N_22446);
nand U22689 (N_22689,N_22451,N_22459);
and U22690 (N_22690,N_22447,N_22501);
nor U22691 (N_22691,N_22472,N_22570);
nor U22692 (N_22692,N_22479,N_22535);
nor U22693 (N_22693,N_22596,N_22538);
xor U22694 (N_22694,N_22577,N_22582);
xor U22695 (N_22695,N_22422,N_22469);
nand U22696 (N_22696,N_22424,N_22402);
xnor U22697 (N_22697,N_22444,N_22414);
and U22698 (N_22698,N_22404,N_22595);
nor U22699 (N_22699,N_22584,N_22558);
and U22700 (N_22700,N_22569,N_22581);
or U22701 (N_22701,N_22563,N_22538);
or U22702 (N_22702,N_22423,N_22549);
nand U22703 (N_22703,N_22541,N_22558);
nor U22704 (N_22704,N_22546,N_22435);
nor U22705 (N_22705,N_22525,N_22443);
or U22706 (N_22706,N_22500,N_22449);
nand U22707 (N_22707,N_22410,N_22403);
or U22708 (N_22708,N_22490,N_22492);
and U22709 (N_22709,N_22568,N_22402);
xor U22710 (N_22710,N_22465,N_22458);
nor U22711 (N_22711,N_22494,N_22486);
nor U22712 (N_22712,N_22580,N_22588);
and U22713 (N_22713,N_22452,N_22469);
xnor U22714 (N_22714,N_22513,N_22432);
and U22715 (N_22715,N_22555,N_22514);
xnor U22716 (N_22716,N_22561,N_22578);
or U22717 (N_22717,N_22550,N_22463);
xor U22718 (N_22718,N_22478,N_22505);
nor U22719 (N_22719,N_22458,N_22423);
and U22720 (N_22720,N_22451,N_22418);
xnor U22721 (N_22721,N_22427,N_22568);
nor U22722 (N_22722,N_22438,N_22517);
and U22723 (N_22723,N_22472,N_22592);
nand U22724 (N_22724,N_22422,N_22429);
xnor U22725 (N_22725,N_22547,N_22401);
nand U22726 (N_22726,N_22499,N_22509);
nor U22727 (N_22727,N_22487,N_22452);
xor U22728 (N_22728,N_22559,N_22522);
xor U22729 (N_22729,N_22432,N_22433);
nand U22730 (N_22730,N_22560,N_22422);
or U22731 (N_22731,N_22558,N_22415);
xnor U22732 (N_22732,N_22561,N_22481);
nor U22733 (N_22733,N_22543,N_22410);
and U22734 (N_22734,N_22578,N_22598);
xnor U22735 (N_22735,N_22421,N_22429);
and U22736 (N_22736,N_22454,N_22440);
xnor U22737 (N_22737,N_22455,N_22461);
xor U22738 (N_22738,N_22493,N_22525);
or U22739 (N_22739,N_22583,N_22573);
xnor U22740 (N_22740,N_22430,N_22495);
nor U22741 (N_22741,N_22552,N_22589);
nand U22742 (N_22742,N_22501,N_22593);
nor U22743 (N_22743,N_22536,N_22538);
xnor U22744 (N_22744,N_22527,N_22535);
or U22745 (N_22745,N_22409,N_22547);
nor U22746 (N_22746,N_22529,N_22508);
nand U22747 (N_22747,N_22515,N_22573);
nand U22748 (N_22748,N_22464,N_22469);
or U22749 (N_22749,N_22446,N_22503);
or U22750 (N_22750,N_22423,N_22576);
xor U22751 (N_22751,N_22505,N_22512);
and U22752 (N_22752,N_22418,N_22478);
and U22753 (N_22753,N_22556,N_22470);
xnor U22754 (N_22754,N_22492,N_22449);
nand U22755 (N_22755,N_22523,N_22569);
or U22756 (N_22756,N_22469,N_22480);
and U22757 (N_22757,N_22558,N_22500);
nand U22758 (N_22758,N_22404,N_22514);
nor U22759 (N_22759,N_22536,N_22482);
and U22760 (N_22760,N_22550,N_22504);
nand U22761 (N_22761,N_22510,N_22456);
and U22762 (N_22762,N_22467,N_22553);
xnor U22763 (N_22763,N_22400,N_22454);
nor U22764 (N_22764,N_22560,N_22467);
xnor U22765 (N_22765,N_22547,N_22497);
nor U22766 (N_22766,N_22592,N_22487);
xnor U22767 (N_22767,N_22466,N_22496);
nor U22768 (N_22768,N_22537,N_22450);
xor U22769 (N_22769,N_22457,N_22407);
and U22770 (N_22770,N_22450,N_22555);
nor U22771 (N_22771,N_22501,N_22479);
nor U22772 (N_22772,N_22570,N_22511);
and U22773 (N_22773,N_22472,N_22555);
nor U22774 (N_22774,N_22594,N_22572);
and U22775 (N_22775,N_22538,N_22406);
and U22776 (N_22776,N_22524,N_22562);
nor U22777 (N_22777,N_22517,N_22533);
nand U22778 (N_22778,N_22523,N_22506);
nand U22779 (N_22779,N_22571,N_22410);
nand U22780 (N_22780,N_22478,N_22544);
nand U22781 (N_22781,N_22504,N_22587);
xor U22782 (N_22782,N_22424,N_22410);
or U22783 (N_22783,N_22590,N_22516);
or U22784 (N_22784,N_22466,N_22594);
nand U22785 (N_22785,N_22471,N_22424);
nand U22786 (N_22786,N_22471,N_22408);
and U22787 (N_22787,N_22486,N_22404);
nor U22788 (N_22788,N_22591,N_22445);
nand U22789 (N_22789,N_22407,N_22461);
xor U22790 (N_22790,N_22428,N_22593);
or U22791 (N_22791,N_22470,N_22435);
xor U22792 (N_22792,N_22578,N_22513);
xor U22793 (N_22793,N_22434,N_22522);
xor U22794 (N_22794,N_22453,N_22484);
or U22795 (N_22795,N_22541,N_22505);
or U22796 (N_22796,N_22457,N_22584);
xnor U22797 (N_22797,N_22426,N_22560);
nand U22798 (N_22798,N_22444,N_22598);
nor U22799 (N_22799,N_22475,N_22493);
nor U22800 (N_22800,N_22618,N_22790);
nand U22801 (N_22801,N_22609,N_22697);
and U22802 (N_22802,N_22757,N_22661);
and U22803 (N_22803,N_22748,N_22674);
and U22804 (N_22804,N_22683,N_22663);
nor U22805 (N_22805,N_22684,N_22787);
and U22806 (N_22806,N_22636,N_22617);
nand U22807 (N_22807,N_22789,N_22729);
xnor U22808 (N_22808,N_22764,N_22677);
or U22809 (N_22809,N_22613,N_22620);
nand U22810 (N_22810,N_22744,N_22666);
nor U22811 (N_22811,N_22640,N_22767);
xor U22812 (N_22812,N_22610,N_22611);
and U22813 (N_22813,N_22777,N_22708);
nor U22814 (N_22814,N_22792,N_22791);
or U22815 (N_22815,N_22711,N_22686);
and U22816 (N_22816,N_22754,N_22793);
or U22817 (N_22817,N_22736,N_22695);
nor U22818 (N_22818,N_22778,N_22654);
nand U22819 (N_22819,N_22702,N_22687);
or U22820 (N_22820,N_22716,N_22662);
and U22821 (N_22821,N_22667,N_22705);
and U22822 (N_22822,N_22615,N_22651);
nand U22823 (N_22823,N_22658,N_22734);
nor U22824 (N_22824,N_22670,N_22723);
xnor U22825 (N_22825,N_22616,N_22626);
nand U22826 (N_22826,N_22632,N_22785);
nor U22827 (N_22827,N_22763,N_22724);
nand U22828 (N_22828,N_22659,N_22760);
nand U22829 (N_22829,N_22621,N_22765);
nand U22830 (N_22830,N_22689,N_22606);
or U22831 (N_22831,N_22707,N_22656);
or U22832 (N_22832,N_22786,N_22650);
nor U22833 (N_22833,N_22741,N_22665);
nor U22834 (N_22834,N_22727,N_22755);
or U22835 (N_22835,N_22795,N_22694);
xnor U22836 (N_22836,N_22739,N_22607);
or U22837 (N_22837,N_22750,N_22699);
or U22838 (N_22838,N_22735,N_22672);
nor U22839 (N_22839,N_22770,N_22655);
nand U22840 (N_22840,N_22649,N_22671);
nand U22841 (N_22841,N_22731,N_22799);
nor U22842 (N_22842,N_22647,N_22718);
nand U22843 (N_22843,N_22660,N_22728);
xnor U22844 (N_22844,N_22706,N_22608);
nor U22845 (N_22845,N_22625,N_22638);
nor U22846 (N_22846,N_22630,N_22779);
or U22847 (N_22847,N_22680,N_22637);
xnor U22848 (N_22848,N_22642,N_22652);
or U22849 (N_22849,N_22641,N_22784);
nand U22850 (N_22850,N_22668,N_22602);
xnor U22851 (N_22851,N_22623,N_22614);
or U22852 (N_22852,N_22752,N_22796);
nor U22853 (N_22853,N_22798,N_22720);
nor U22854 (N_22854,N_22781,N_22710);
and U22855 (N_22855,N_22797,N_22775);
nand U22856 (N_22856,N_22730,N_22693);
and U22857 (N_22857,N_22601,N_22769);
and U22858 (N_22858,N_22624,N_22622);
nand U22859 (N_22859,N_22740,N_22631);
xnor U22860 (N_22860,N_22751,N_22756);
nand U22861 (N_22861,N_22717,N_22773);
nor U22862 (N_22862,N_22761,N_22732);
xor U22863 (N_22863,N_22743,N_22675);
or U22864 (N_22864,N_22762,N_22691);
xor U22865 (N_22865,N_22749,N_22629);
or U22866 (N_22866,N_22628,N_22627);
nand U22867 (N_22867,N_22681,N_22737);
nor U22868 (N_22868,N_22676,N_22692);
or U22869 (N_22869,N_22747,N_22633);
xnor U22870 (N_22870,N_22635,N_22700);
or U22871 (N_22871,N_22772,N_22657);
nor U22872 (N_22872,N_22733,N_22745);
and U22873 (N_22873,N_22771,N_22788);
and U22874 (N_22874,N_22673,N_22709);
xnor U22875 (N_22875,N_22688,N_22653);
and U22876 (N_22876,N_22726,N_22715);
or U22877 (N_22877,N_22669,N_22678);
or U22878 (N_22878,N_22604,N_22738);
nor U22879 (N_22879,N_22648,N_22782);
or U22880 (N_22880,N_22783,N_22643);
or U22881 (N_22881,N_22701,N_22753);
or U22882 (N_22882,N_22758,N_22600);
xor U22883 (N_22883,N_22703,N_22679);
nand U22884 (N_22884,N_22696,N_22704);
nor U22885 (N_22885,N_22768,N_22722);
nor U22886 (N_22886,N_22714,N_22646);
nand U22887 (N_22887,N_22794,N_22690);
nand U22888 (N_22888,N_22774,N_22713);
nor U22889 (N_22889,N_22712,N_22634);
or U22890 (N_22890,N_22605,N_22698);
xor U22891 (N_22891,N_22682,N_22746);
and U22892 (N_22892,N_22719,N_22603);
nand U22893 (N_22893,N_22759,N_22612);
nand U22894 (N_22894,N_22619,N_22780);
nor U22895 (N_22895,N_22742,N_22725);
nor U22896 (N_22896,N_22721,N_22776);
nor U22897 (N_22897,N_22645,N_22766);
or U22898 (N_22898,N_22644,N_22664);
nand U22899 (N_22899,N_22685,N_22639);
and U22900 (N_22900,N_22747,N_22706);
xor U22901 (N_22901,N_22635,N_22627);
and U22902 (N_22902,N_22740,N_22775);
nor U22903 (N_22903,N_22787,N_22796);
and U22904 (N_22904,N_22715,N_22699);
nand U22905 (N_22905,N_22788,N_22762);
xor U22906 (N_22906,N_22773,N_22731);
xnor U22907 (N_22907,N_22620,N_22671);
xnor U22908 (N_22908,N_22768,N_22770);
xnor U22909 (N_22909,N_22657,N_22655);
nand U22910 (N_22910,N_22647,N_22717);
or U22911 (N_22911,N_22733,N_22634);
nand U22912 (N_22912,N_22662,N_22649);
nor U22913 (N_22913,N_22630,N_22706);
nand U22914 (N_22914,N_22758,N_22639);
nand U22915 (N_22915,N_22652,N_22667);
and U22916 (N_22916,N_22777,N_22730);
nor U22917 (N_22917,N_22688,N_22637);
nand U22918 (N_22918,N_22734,N_22711);
and U22919 (N_22919,N_22745,N_22681);
and U22920 (N_22920,N_22661,N_22798);
and U22921 (N_22921,N_22670,N_22644);
nand U22922 (N_22922,N_22654,N_22653);
and U22923 (N_22923,N_22796,N_22665);
or U22924 (N_22924,N_22698,N_22638);
xnor U22925 (N_22925,N_22779,N_22798);
xor U22926 (N_22926,N_22708,N_22726);
or U22927 (N_22927,N_22700,N_22739);
nor U22928 (N_22928,N_22618,N_22695);
xor U22929 (N_22929,N_22615,N_22621);
xor U22930 (N_22930,N_22740,N_22776);
nand U22931 (N_22931,N_22648,N_22739);
xor U22932 (N_22932,N_22640,N_22736);
xor U22933 (N_22933,N_22789,N_22641);
or U22934 (N_22934,N_22655,N_22751);
or U22935 (N_22935,N_22668,N_22761);
xor U22936 (N_22936,N_22611,N_22687);
nor U22937 (N_22937,N_22617,N_22796);
nor U22938 (N_22938,N_22761,N_22679);
and U22939 (N_22939,N_22696,N_22713);
or U22940 (N_22940,N_22627,N_22729);
nand U22941 (N_22941,N_22710,N_22697);
xnor U22942 (N_22942,N_22787,N_22746);
nor U22943 (N_22943,N_22642,N_22777);
and U22944 (N_22944,N_22603,N_22625);
and U22945 (N_22945,N_22706,N_22666);
nor U22946 (N_22946,N_22749,N_22724);
xnor U22947 (N_22947,N_22767,N_22784);
nand U22948 (N_22948,N_22658,N_22793);
and U22949 (N_22949,N_22600,N_22675);
or U22950 (N_22950,N_22748,N_22757);
nor U22951 (N_22951,N_22778,N_22624);
nand U22952 (N_22952,N_22767,N_22756);
or U22953 (N_22953,N_22794,N_22796);
or U22954 (N_22954,N_22736,N_22791);
or U22955 (N_22955,N_22621,N_22711);
and U22956 (N_22956,N_22769,N_22784);
xor U22957 (N_22957,N_22675,N_22797);
or U22958 (N_22958,N_22630,N_22660);
and U22959 (N_22959,N_22654,N_22733);
nand U22960 (N_22960,N_22672,N_22655);
or U22961 (N_22961,N_22786,N_22774);
or U22962 (N_22962,N_22756,N_22660);
nor U22963 (N_22963,N_22763,N_22656);
or U22964 (N_22964,N_22622,N_22772);
and U22965 (N_22965,N_22684,N_22646);
and U22966 (N_22966,N_22698,N_22690);
or U22967 (N_22967,N_22711,N_22791);
nor U22968 (N_22968,N_22611,N_22681);
nand U22969 (N_22969,N_22737,N_22621);
and U22970 (N_22970,N_22638,N_22796);
and U22971 (N_22971,N_22668,N_22720);
nand U22972 (N_22972,N_22735,N_22649);
xor U22973 (N_22973,N_22714,N_22711);
nor U22974 (N_22974,N_22709,N_22779);
and U22975 (N_22975,N_22716,N_22733);
or U22976 (N_22976,N_22626,N_22730);
xnor U22977 (N_22977,N_22776,N_22790);
or U22978 (N_22978,N_22751,N_22757);
nor U22979 (N_22979,N_22750,N_22771);
or U22980 (N_22980,N_22630,N_22736);
or U22981 (N_22981,N_22784,N_22776);
and U22982 (N_22982,N_22694,N_22665);
and U22983 (N_22983,N_22618,N_22720);
and U22984 (N_22984,N_22759,N_22658);
xor U22985 (N_22985,N_22627,N_22649);
and U22986 (N_22986,N_22673,N_22798);
xor U22987 (N_22987,N_22689,N_22675);
and U22988 (N_22988,N_22772,N_22680);
and U22989 (N_22989,N_22753,N_22690);
xor U22990 (N_22990,N_22725,N_22729);
nand U22991 (N_22991,N_22693,N_22794);
or U22992 (N_22992,N_22784,N_22653);
nand U22993 (N_22993,N_22732,N_22603);
xor U22994 (N_22994,N_22644,N_22717);
and U22995 (N_22995,N_22681,N_22666);
xor U22996 (N_22996,N_22764,N_22718);
nand U22997 (N_22997,N_22720,N_22655);
xnor U22998 (N_22998,N_22639,N_22605);
xnor U22999 (N_22999,N_22790,N_22678);
xor U23000 (N_23000,N_22990,N_22999);
or U23001 (N_23001,N_22982,N_22874);
xor U23002 (N_23002,N_22961,N_22923);
nand U23003 (N_23003,N_22965,N_22866);
nor U23004 (N_23004,N_22868,N_22869);
nor U23005 (N_23005,N_22806,N_22996);
xnor U23006 (N_23006,N_22822,N_22831);
nand U23007 (N_23007,N_22964,N_22946);
nand U23008 (N_23008,N_22947,N_22888);
nand U23009 (N_23009,N_22871,N_22944);
and U23010 (N_23010,N_22921,N_22897);
nand U23011 (N_23011,N_22821,N_22854);
nor U23012 (N_23012,N_22889,N_22972);
xor U23013 (N_23013,N_22812,N_22914);
and U23014 (N_23014,N_22814,N_22922);
or U23015 (N_23015,N_22918,N_22895);
and U23016 (N_23016,N_22925,N_22937);
nor U23017 (N_23017,N_22863,N_22911);
and U23018 (N_23018,N_22856,N_22892);
nand U23019 (N_23019,N_22930,N_22837);
xnor U23020 (N_23020,N_22899,N_22977);
xnor U23021 (N_23021,N_22953,N_22875);
nand U23022 (N_23022,N_22830,N_22942);
or U23023 (N_23023,N_22991,N_22893);
nor U23024 (N_23024,N_22915,N_22809);
nor U23025 (N_23025,N_22960,N_22848);
or U23026 (N_23026,N_22872,N_22825);
xnor U23027 (N_23027,N_22917,N_22966);
nor U23028 (N_23028,N_22910,N_22943);
nor U23029 (N_23029,N_22846,N_22912);
and U23030 (N_23030,N_22924,N_22989);
nand U23031 (N_23031,N_22852,N_22802);
xnor U23032 (N_23032,N_22808,N_22933);
nor U23033 (N_23033,N_22968,N_22976);
nand U23034 (N_23034,N_22959,N_22950);
nand U23035 (N_23035,N_22956,N_22967);
xor U23036 (N_23036,N_22867,N_22974);
and U23037 (N_23037,N_22890,N_22804);
nand U23038 (N_23038,N_22980,N_22811);
xnor U23039 (N_23039,N_22979,N_22800);
and U23040 (N_23040,N_22850,N_22948);
or U23041 (N_23041,N_22884,N_22955);
nand U23042 (N_23042,N_22842,N_22987);
xor U23043 (N_23043,N_22908,N_22881);
or U23044 (N_23044,N_22969,N_22834);
xor U23045 (N_23045,N_22823,N_22843);
and U23046 (N_23046,N_22828,N_22876);
and U23047 (N_23047,N_22981,N_22820);
or U23048 (N_23048,N_22882,N_22907);
nor U23049 (N_23049,N_22905,N_22932);
or U23050 (N_23050,N_22975,N_22878);
xor U23051 (N_23051,N_22940,N_22845);
and U23052 (N_23052,N_22819,N_22906);
nand U23053 (N_23053,N_22986,N_22997);
xor U23054 (N_23054,N_22952,N_22807);
nor U23055 (N_23055,N_22826,N_22896);
nand U23056 (N_23056,N_22844,N_22927);
and U23057 (N_23057,N_22886,N_22916);
nor U23058 (N_23058,N_22971,N_22898);
and U23059 (N_23059,N_22902,N_22957);
xnor U23060 (N_23060,N_22929,N_22883);
or U23061 (N_23061,N_22873,N_22861);
nor U23062 (N_23062,N_22855,N_22988);
nand U23063 (N_23063,N_22877,N_22939);
or U23064 (N_23064,N_22926,N_22951);
and U23065 (N_23065,N_22985,N_22909);
xor U23066 (N_23066,N_22813,N_22851);
or U23067 (N_23067,N_22919,N_22865);
nor U23068 (N_23068,N_22803,N_22857);
or U23069 (N_23069,N_22864,N_22903);
xor U23070 (N_23070,N_22836,N_22900);
nand U23071 (N_23071,N_22879,N_22954);
and U23072 (N_23072,N_22853,N_22962);
or U23073 (N_23073,N_22904,N_22860);
or U23074 (N_23074,N_22832,N_22849);
nand U23075 (N_23075,N_22931,N_22949);
and U23076 (N_23076,N_22841,N_22847);
nor U23077 (N_23077,N_22816,N_22862);
and U23078 (N_23078,N_22839,N_22894);
xnor U23079 (N_23079,N_22833,N_22941);
nor U23080 (N_23080,N_22815,N_22994);
nor U23081 (N_23081,N_22936,N_22838);
xnor U23082 (N_23082,N_22978,N_22870);
nor U23083 (N_23083,N_22995,N_22885);
xor U23084 (N_23084,N_22801,N_22993);
nor U23085 (N_23085,N_22998,N_22920);
nor U23086 (N_23086,N_22938,N_22887);
xnor U23087 (N_23087,N_22992,N_22805);
xor U23088 (N_23088,N_22810,N_22934);
and U23089 (N_23089,N_22827,N_22984);
and U23090 (N_23090,N_22858,N_22913);
nand U23091 (N_23091,N_22901,N_22880);
and U23092 (N_23092,N_22935,N_22970);
xor U23093 (N_23093,N_22973,N_22824);
nor U23094 (N_23094,N_22817,N_22928);
nor U23095 (N_23095,N_22963,N_22835);
nor U23096 (N_23096,N_22818,N_22891);
and U23097 (N_23097,N_22859,N_22958);
xor U23098 (N_23098,N_22983,N_22840);
xor U23099 (N_23099,N_22829,N_22945);
nor U23100 (N_23100,N_22964,N_22949);
xor U23101 (N_23101,N_22986,N_22950);
nand U23102 (N_23102,N_22850,N_22957);
or U23103 (N_23103,N_22801,N_22914);
or U23104 (N_23104,N_22825,N_22942);
or U23105 (N_23105,N_22892,N_22919);
xor U23106 (N_23106,N_22981,N_22924);
xnor U23107 (N_23107,N_22956,N_22992);
nand U23108 (N_23108,N_22902,N_22886);
nor U23109 (N_23109,N_22947,N_22990);
nand U23110 (N_23110,N_22813,N_22869);
nand U23111 (N_23111,N_22921,N_22827);
or U23112 (N_23112,N_22843,N_22893);
or U23113 (N_23113,N_22865,N_22965);
and U23114 (N_23114,N_22889,N_22802);
nor U23115 (N_23115,N_22816,N_22876);
xnor U23116 (N_23116,N_22801,N_22809);
and U23117 (N_23117,N_22973,N_22857);
nand U23118 (N_23118,N_22910,N_22896);
xnor U23119 (N_23119,N_22822,N_22941);
and U23120 (N_23120,N_22820,N_22802);
or U23121 (N_23121,N_22976,N_22899);
nand U23122 (N_23122,N_22872,N_22865);
and U23123 (N_23123,N_22976,N_22856);
nor U23124 (N_23124,N_22834,N_22940);
or U23125 (N_23125,N_22891,N_22948);
and U23126 (N_23126,N_22995,N_22825);
nor U23127 (N_23127,N_22966,N_22945);
xor U23128 (N_23128,N_22974,N_22836);
or U23129 (N_23129,N_22917,N_22998);
or U23130 (N_23130,N_22857,N_22819);
nor U23131 (N_23131,N_22913,N_22871);
or U23132 (N_23132,N_22951,N_22879);
or U23133 (N_23133,N_22907,N_22898);
nand U23134 (N_23134,N_22862,N_22845);
nor U23135 (N_23135,N_22878,N_22921);
and U23136 (N_23136,N_22926,N_22946);
nand U23137 (N_23137,N_22854,N_22987);
or U23138 (N_23138,N_22841,N_22851);
nor U23139 (N_23139,N_22885,N_22920);
or U23140 (N_23140,N_22887,N_22818);
nor U23141 (N_23141,N_22914,N_22963);
nor U23142 (N_23142,N_22910,N_22804);
and U23143 (N_23143,N_22826,N_22939);
and U23144 (N_23144,N_22880,N_22864);
xor U23145 (N_23145,N_22886,N_22905);
and U23146 (N_23146,N_22804,N_22805);
xor U23147 (N_23147,N_22820,N_22827);
or U23148 (N_23148,N_22996,N_22947);
nand U23149 (N_23149,N_22861,N_22898);
or U23150 (N_23150,N_22813,N_22992);
xor U23151 (N_23151,N_22921,N_22982);
and U23152 (N_23152,N_22874,N_22914);
xnor U23153 (N_23153,N_22916,N_22866);
xnor U23154 (N_23154,N_22887,N_22868);
or U23155 (N_23155,N_22889,N_22839);
nand U23156 (N_23156,N_22855,N_22948);
nand U23157 (N_23157,N_22980,N_22824);
or U23158 (N_23158,N_22848,N_22863);
and U23159 (N_23159,N_22958,N_22931);
xnor U23160 (N_23160,N_22899,N_22891);
and U23161 (N_23161,N_22935,N_22942);
nor U23162 (N_23162,N_22890,N_22913);
nand U23163 (N_23163,N_22894,N_22907);
and U23164 (N_23164,N_22934,N_22870);
xor U23165 (N_23165,N_22803,N_22828);
nand U23166 (N_23166,N_22975,N_22856);
xnor U23167 (N_23167,N_22962,N_22825);
nand U23168 (N_23168,N_22962,N_22991);
nand U23169 (N_23169,N_22804,N_22823);
and U23170 (N_23170,N_22993,N_22841);
nor U23171 (N_23171,N_22931,N_22882);
or U23172 (N_23172,N_22827,N_22925);
xnor U23173 (N_23173,N_22874,N_22995);
and U23174 (N_23174,N_22933,N_22966);
xnor U23175 (N_23175,N_22945,N_22801);
nor U23176 (N_23176,N_22882,N_22820);
nor U23177 (N_23177,N_22845,N_22826);
or U23178 (N_23178,N_22846,N_22886);
nand U23179 (N_23179,N_22999,N_22894);
xor U23180 (N_23180,N_22913,N_22852);
nand U23181 (N_23181,N_22914,N_22966);
and U23182 (N_23182,N_22938,N_22985);
and U23183 (N_23183,N_22827,N_22956);
and U23184 (N_23184,N_22944,N_22881);
nor U23185 (N_23185,N_22938,N_22835);
and U23186 (N_23186,N_22966,N_22809);
xnor U23187 (N_23187,N_22858,N_22814);
or U23188 (N_23188,N_22816,N_22881);
nor U23189 (N_23189,N_22945,N_22865);
or U23190 (N_23190,N_22867,N_22824);
nor U23191 (N_23191,N_22935,N_22806);
nand U23192 (N_23192,N_22971,N_22902);
xor U23193 (N_23193,N_22885,N_22954);
xnor U23194 (N_23194,N_22803,N_22834);
nor U23195 (N_23195,N_22907,N_22923);
or U23196 (N_23196,N_22809,N_22919);
xnor U23197 (N_23197,N_22866,N_22823);
xor U23198 (N_23198,N_22807,N_22845);
nor U23199 (N_23199,N_22870,N_22960);
xnor U23200 (N_23200,N_23130,N_23100);
nand U23201 (N_23201,N_23113,N_23104);
nand U23202 (N_23202,N_23053,N_23154);
xnor U23203 (N_23203,N_23182,N_23106);
nor U23204 (N_23204,N_23138,N_23064);
xnor U23205 (N_23205,N_23176,N_23185);
and U23206 (N_23206,N_23028,N_23110);
nor U23207 (N_23207,N_23036,N_23096);
or U23208 (N_23208,N_23128,N_23139);
and U23209 (N_23209,N_23107,N_23172);
or U23210 (N_23210,N_23180,N_23060);
nand U23211 (N_23211,N_23166,N_23038);
and U23212 (N_23212,N_23194,N_23146);
xor U23213 (N_23213,N_23145,N_23078);
nand U23214 (N_23214,N_23134,N_23167);
and U23215 (N_23215,N_23079,N_23099);
nand U23216 (N_23216,N_23184,N_23118);
or U23217 (N_23217,N_23066,N_23189);
and U23218 (N_23218,N_23168,N_23177);
nor U23219 (N_23219,N_23089,N_23178);
nand U23220 (N_23220,N_23093,N_23121);
and U23221 (N_23221,N_23042,N_23010);
nand U23222 (N_23222,N_23188,N_23050);
or U23223 (N_23223,N_23190,N_23068);
nor U23224 (N_23224,N_23080,N_23020);
nand U23225 (N_23225,N_23158,N_23045);
or U23226 (N_23226,N_23148,N_23087);
or U23227 (N_23227,N_23131,N_23092);
nor U23228 (N_23228,N_23072,N_23102);
and U23229 (N_23229,N_23012,N_23143);
nand U23230 (N_23230,N_23056,N_23127);
xnor U23231 (N_23231,N_23044,N_23009);
or U23232 (N_23232,N_23007,N_23197);
or U23233 (N_23233,N_23062,N_23112);
nand U23234 (N_23234,N_23065,N_23001);
nand U23235 (N_23235,N_23006,N_23005);
or U23236 (N_23236,N_23024,N_23082);
nor U23237 (N_23237,N_23091,N_23126);
xnor U23238 (N_23238,N_23164,N_23047);
nor U23239 (N_23239,N_23141,N_23129);
nand U23240 (N_23240,N_23023,N_23063);
xor U23241 (N_23241,N_23193,N_23156);
and U23242 (N_23242,N_23013,N_23049);
or U23243 (N_23243,N_23187,N_23054);
xnor U23244 (N_23244,N_23097,N_23122);
nand U23245 (N_23245,N_23059,N_23192);
nor U23246 (N_23246,N_23147,N_23155);
and U23247 (N_23247,N_23175,N_23037);
nor U23248 (N_23248,N_23095,N_23090);
and U23249 (N_23249,N_23046,N_23116);
xnor U23250 (N_23250,N_23011,N_23186);
nor U23251 (N_23251,N_23101,N_23033);
or U23252 (N_23252,N_23160,N_23018);
and U23253 (N_23253,N_23161,N_23081);
nor U23254 (N_23254,N_23198,N_23026);
nand U23255 (N_23255,N_23048,N_23008);
xor U23256 (N_23256,N_23016,N_23159);
xnor U23257 (N_23257,N_23051,N_23058);
nand U23258 (N_23258,N_23021,N_23165);
and U23259 (N_23259,N_23070,N_23019);
nand U23260 (N_23260,N_23157,N_23108);
xnor U23261 (N_23261,N_23075,N_23183);
xnor U23262 (N_23262,N_23071,N_23027);
nor U23263 (N_23263,N_23196,N_23031);
or U23264 (N_23264,N_23109,N_23195);
and U23265 (N_23265,N_23140,N_23014);
and U23266 (N_23266,N_23135,N_23083);
and U23267 (N_23267,N_23174,N_23144);
nor U23268 (N_23268,N_23142,N_23114);
nand U23269 (N_23269,N_23133,N_23032);
nand U23270 (N_23270,N_23123,N_23034);
nor U23271 (N_23271,N_23040,N_23136);
or U23272 (N_23272,N_23191,N_23169);
and U23273 (N_23273,N_23022,N_23003);
nor U23274 (N_23274,N_23077,N_23043);
or U23275 (N_23275,N_23055,N_23088);
or U23276 (N_23276,N_23086,N_23041);
or U23277 (N_23277,N_23057,N_23004);
or U23278 (N_23278,N_23171,N_23163);
and U23279 (N_23279,N_23111,N_23067);
nand U23280 (N_23280,N_23125,N_23061);
nor U23281 (N_23281,N_23153,N_23150);
nor U23282 (N_23282,N_23103,N_23173);
xor U23283 (N_23283,N_23035,N_23000);
nor U23284 (N_23284,N_23105,N_23069);
nor U23285 (N_23285,N_23199,N_23015);
nand U23286 (N_23286,N_23152,N_23120);
and U23287 (N_23287,N_23179,N_23039);
xor U23288 (N_23288,N_23132,N_23030);
nor U23289 (N_23289,N_23137,N_23025);
xnor U23290 (N_23290,N_23094,N_23017);
and U23291 (N_23291,N_23115,N_23073);
nor U23292 (N_23292,N_23162,N_23181);
or U23293 (N_23293,N_23117,N_23170);
nor U23294 (N_23294,N_23124,N_23029);
or U23295 (N_23295,N_23074,N_23076);
xnor U23296 (N_23296,N_23002,N_23052);
and U23297 (N_23297,N_23119,N_23098);
or U23298 (N_23298,N_23084,N_23149);
nor U23299 (N_23299,N_23151,N_23085);
xnor U23300 (N_23300,N_23113,N_23176);
xor U23301 (N_23301,N_23064,N_23154);
and U23302 (N_23302,N_23154,N_23130);
nand U23303 (N_23303,N_23105,N_23113);
xor U23304 (N_23304,N_23130,N_23192);
xor U23305 (N_23305,N_23030,N_23158);
and U23306 (N_23306,N_23115,N_23067);
nor U23307 (N_23307,N_23197,N_23121);
or U23308 (N_23308,N_23103,N_23158);
or U23309 (N_23309,N_23187,N_23113);
nand U23310 (N_23310,N_23085,N_23179);
or U23311 (N_23311,N_23030,N_23078);
nand U23312 (N_23312,N_23102,N_23026);
and U23313 (N_23313,N_23002,N_23168);
or U23314 (N_23314,N_23051,N_23007);
nand U23315 (N_23315,N_23025,N_23034);
or U23316 (N_23316,N_23071,N_23040);
or U23317 (N_23317,N_23087,N_23138);
or U23318 (N_23318,N_23003,N_23036);
nand U23319 (N_23319,N_23082,N_23016);
nand U23320 (N_23320,N_23049,N_23115);
and U23321 (N_23321,N_23040,N_23189);
or U23322 (N_23322,N_23021,N_23116);
or U23323 (N_23323,N_23007,N_23196);
and U23324 (N_23324,N_23081,N_23020);
and U23325 (N_23325,N_23103,N_23165);
and U23326 (N_23326,N_23017,N_23179);
nor U23327 (N_23327,N_23109,N_23077);
xnor U23328 (N_23328,N_23043,N_23039);
nor U23329 (N_23329,N_23015,N_23192);
nor U23330 (N_23330,N_23079,N_23182);
and U23331 (N_23331,N_23072,N_23131);
nor U23332 (N_23332,N_23098,N_23006);
xnor U23333 (N_23333,N_23168,N_23179);
or U23334 (N_23334,N_23110,N_23109);
xor U23335 (N_23335,N_23179,N_23045);
xnor U23336 (N_23336,N_23170,N_23168);
xor U23337 (N_23337,N_23042,N_23007);
nand U23338 (N_23338,N_23096,N_23130);
or U23339 (N_23339,N_23014,N_23127);
or U23340 (N_23340,N_23061,N_23082);
xor U23341 (N_23341,N_23165,N_23038);
nand U23342 (N_23342,N_23090,N_23138);
and U23343 (N_23343,N_23028,N_23112);
xor U23344 (N_23344,N_23034,N_23183);
nand U23345 (N_23345,N_23006,N_23136);
nand U23346 (N_23346,N_23162,N_23066);
or U23347 (N_23347,N_23061,N_23058);
nor U23348 (N_23348,N_23025,N_23005);
or U23349 (N_23349,N_23196,N_23038);
nor U23350 (N_23350,N_23100,N_23166);
or U23351 (N_23351,N_23152,N_23015);
nand U23352 (N_23352,N_23112,N_23012);
and U23353 (N_23353,N_23101,N_23035);
nand U23354 (N_23354,N_23006,N_23198);
nand U23355 (N_23355,N_23039,N_23001);
nand U23356 (N_23356,N_23137,N_23118);
and U23357 (N_23357,N_23179,N_23073);
and U23358 (N_23358,N_23195,N_23003);
and U23359 (N_23359,N_23019,N_23066);
nand U23360 (N_23360,N_23039,N_23076);
nor U23361 (N_23361,N_23088,N_23076);
nor U23362 (N_23362,N_23164,N_23009);
nand U23363 (N_23363,N_23160,N_23023);
nand U23364 (N_23364,N_23027,N_23099);
xor U23365 (N_23365,N_23184,N_23173);
nor U23366 (N_23366,N_23172,N_23096);
xnor U23367 (N_23367,N_23095,N_23028);
xor U23368 (N_23368,N_23003,N_23118);
or U23369 (N_23369,N_23078,N_23090);
nor U23370 (N_23370,N_23188,N_23021);
and U23371 (N_23371,N_23040,N_23070);
or U23372 (N_23372,N_23172,N_23114);
nor U23373 (N_23373,N_23076,N_23165);
and U23374 (N_23374,N_23030,N_23106);
nor U23375 (N_23375,N_23160,N_23170);
or U23376 (N_23376,N_23140,N_23085);
nand U23377 (N_23377,N_23105,N_23047);
xor U23378 (N_23378,N_23109,N_23098);
nand U23379 (N_23379,N_23148,N_23081);
xor U23380 (N_23380,N_23147,N_23130);
xor U23381 (N_23381,N_23089,N_23012);
nand U23382 (N_23382,N_23110,N_23088);
nor U23383 (N_23383,N_23100,N_23174);
or U23384 (N_23384,N_23180,N_23005);
nand U23385 (N_23385,N_23139,N_23083);
xnor U23386 (N_23386,N_23118,N_23067);
or U23387 (N_23387,N_23147,N_23128);
xnor U23388 (N_23388,N_23025,N_23042);
or U23389 (N_23389,N_23121,N_23185);
nand U23390 (N_23390,N_23157,N_23011);
and U23391 (N_23391,N_23196,N_23070);
and U23392 (N_23392,N_23052,N_23115);
and U23393 (N_23393,N_23180,N_23104);
nor U23394 (N_23394,N_23001,N_23041);
and U23395 (N_23395,N_23071,N_23180);
xnor U23396 (N_23396,N_23153,N_23163);
nor U23397 (N_23397,N_23176,N_23169);
nor U23398 (N_23398,N_23174,N_23160);
nand U23399 (N_23399,N_23149,N_23009);
or U23400 (N_23400,N_23386,N_23352);
and U23401 (N_23401,N_23369,N_23270);
or U23402 (N_23402,N_23327,N_23227);
or U23403 (N_23403,N_23371,N_23334);
nor U23404 (N_23404,N_23296,N_23230);
nand U23405 (N_23405,N_23228,N_23220);
nand U23406 (N_23406,N_23246,N_23316);
or U23407 (N_23407,N_23251,N_23289);
or U23408 (N_23408,N_23350,N_23257);
or U23409 (N_23409,N_23259,N_23254);
nand U23410 (N_23410,N_23272,N_23384);
nand U23411 (N_23411,N_23356,N_23203);
and U23412 (N_23412,N_23382,N_23313);
or U23413 (N_23413,N_23359,N_23312);
xnor U23414 (N_23414,N_23311,N_23361);
and U23415 (N_23415,N_23391,N_23200);
nand U23416 (N_23416,N_23233,N_23280);
nand U23417 (N_23417,N_23201,N_23278);
or U23418 (N_23418,N_23217,N_23247);
or U23419 (N_23419,N_23263,N_23380);
xnor U23420 (N_23420,N_23210,N_23378);
nand U23421 (N_23421,N_23224,N_23301);
xnor U23422 (N_23422,N_23261,N_23277);
or U23423 (N_23423,N_23331,N_23337);
nand U23424 (N_23424,N_23234,N_23357);
xor U23425 (N_23425,N_23349,N_23381);
or U23426 (N_23426,N_23319,N_23281);
nand U23427 (N_23427,N_23387,N_23205);
nand U23428 (N_23428,N_23245,N_23256);
xnor U23429 (N_23429,N_23336,N_23379);
and U23430 (N_23430,N_23383,N_23239);
nand U23431 (N_23431,N_23339,N_23358);
xor U23432 (N_23432,N_23354,N_23287);
or U23433 (N_23433,N_23290,N_23335);
nand U23434 (N_23434,N_23322,N_23218);
or U23435 (N_23435,N_23252,N_23330);
and U23436 (N_23436,N_23286,N_23271);
xor U23437 (N_23437,N_23208,N_23345);
and U23438 (N_23438,N_23388,N_23211);
xor U23439 (N_23439,N_23212,N_23395);
nand U23440 (N_23440,N_23275,N_23238);
xnor U23441 (N_23441,N_23207,N_23206);
nand U23442 (N_23442,N_23393,N_23372);
and U23443 (N_23443,N_23225,N_23340);
nor U23444 (N_23444,N_23276,N_23294);
or U23445 (N_23445,N_23293,N_23202);
or U23446 (N_23446,N_23324,N_23344);
nand U23447 (N_23447,N_23266,N_23204);
nand U23448 (N_23448,N_23332,N_23273);
nor U23449 (N_23449,N_23355,N_23338);
xor U23450 (N_23450,N_23363,N_23267);
nor U23451 (N_23451,N_23248,N_23346);
and U23452 (N_23452,N_23250,N_23295);
nand U23453 (N_23453,N_23236,N_23329);
xor U23454 (N_23454,N_23374,N_23365);
or U23455 (N_23455,N_23285,N_23341);
nor U23456 (N_23456,N_23398,N_23223);
or U23457 (N_23457,N_23221,N_23244);
xnor U23458 (N_23458,N_23308,N_23370);
nor U23459 (N_23459,N_23325,N_23368);
or U23460 (N_23460,N_23307,N_23328);
nor U23461 (N_23461,N_23399,N_23343);
xnor U23462 (N_23462,N_23347,N_23282);
nand U23463 (N_23463,N_23213,N_23314);
and U23464 (N_23464,N_23269,N_23255);
nor U23465 (N_23465,N_23373,N_23229);
and U23466 (N_23466,N_23226,N_23351);
xor U23467 (N_23467,N_23231,N_23243);
and U23468 (N_23468,N_23377,N_23375);
nor U23469 (N_23469,N_23279,N_23367);
nor U23470 (N_23470,N_23333,N_23326);
nor U23471 (N_23471,N_23249,N_23241);
or U23472 (N_23472,N_23253,N_23235);
or U23473 (N_23473,N_23303,N_23315);
nand U23474 (N_23474,N_23306,N_23215);
nor U23475 (N_23475,N_23321,N_23304);
nor U23476 (N_23476,N_23390,N_23288);
xor U23477 (N_23477,N_23300,N_23362);
and U23478 (N_23478,N_23222,N_23317);
nand U23479 (N_23479,N_23284,N_23342);
or U23480 (N_23480,N_23360,N_23214);
nand U23481 (N_23481,N_23240,N_23298);
and U23482 (N_23482,N_23291,N_23397);
xnor U23483 (N_23483,N_23262,N_23265);
nand U23484 (N_23484,N_23323,N_23242);
or U23485 (N_23485,N_23394,N_23309);
or U23486 (N_23486,N_23364,N_23389);
xor U23487 (N_23487,N_23353,N_23219);
and U23488 (N_23488,N_23237,N_23318);
and U23489 (N_23489,N_23396,N_23268);
nor U23490 (N_23490,N_23299,N_23292);
nor U23491 (N_23491,N_23258,N_23216);
or U23492 (N_23492,N_23320,N_23297);
and U23493 (N_23493,N_23348,N_23283);
xor U23494 (N_23494,N_23392,N_23310);
and U23495 (N_23495,N_23302,N_23305);
and U23496 (N_23496,N_23366,N_23274);
xor U23497 (N_23497,N_23232,N_23264);
xor U23498 (N_23498,N_23385,N_23209);
nor U23499 (N_23499,N_23376,N_23260);
nor U23500 (N_23500,N_23266,N_23290);
or U23501 (N_23501,N_23223,N_23225);
nor U23502 (N_23502,N_23370,N_23286);
nand U23503 (N_23503,N_23364,N_23264);
and U23504 (N_23504,N_23244,N_23236);
or U23505 (N_23505,N_23249,N_23243);
xnor U23506 (N_23506,N_23304,N_23241);
xor U23507 (N_23507,N_23241,N_23334);
nand U23508 (N_23508,N_23361,N_23226);
xor U23509 (N_23509,N_23332,N_23381);
or U23510 (N_23510,N_23287,N_23262);
and U23511 (N_23511,N_23331,N_23286);
and U23512 (N_23512,N_23324,N_23386);
xnor U23513 (N_23513,N_23328,N_23375);
nand U23514 (N_23514,N_23375,N_23204);
or U23515 (N_23515,N_23363,N_23265);
nand U23516 (N_23516,N_23293,N_23391);
nand U23517 (N_23517,N_23347,N_23321);
nor U23518 (N_23518,N_23321,N_23269);
nor U23519 (N_23519,N_23285,N_23277);
or U23520 (N_23520,N_23207,N_23345);
xnor U23521 (N_23521,N_23314,N_23352);
xor U23522 (N_23522,N_23226,N_23207);
nand U23523 (N_23523,N_23331,N_23306);
or U23524 (N_23524,N_23301,N_23334);
nand U23525 (N_23525,N_23225,N_23248);
nand U23526 (N_23526,N_23204,N_23283);
xor U23527 (N_23527,N_23361,N_23360);
xor U23528 (N_23528,N_23293,N_23237);
nand U23529 (N_23529,N_23335,N_23362);
xor U23530 (N_23530,N_23387,N_23259);
nand U23531 (N_23531,N_23323,N_23300);
nand U23532 (N_23532,N_23279,N_23294);
and U23533 (N_23533,N_23214,N_23228);
or U23534 (N_23534,N_23233,N_23265);
or U23535 (N_23535,N_23216,N_23208);
or U23536 (N_23536,N_23278,N_23295);
nor U23537 (N_23537,N_23222,N_23266);
xnor U23538 (N_23538,N_23369,N_23233);
and U23539 (N_23539,N_23388,N_23260);
and U23540 (N_23540,N_23250,N_23315);
or U23541 (N_23541,N_23304,N_23224);
and U23542 (N_23542,N_23276,N_23217);
or U23543 (N_23543,N_23200,N_23369);
nor U23544 (N_23544,N_23348,N_23278);
and U23545 (N_23545,N_23327,N_23201);
and U23546 (N_23546,N_23244,N_23374);
and U23547 (N_23547,N_23242,N_23284);
nor U23548 (N_23548,N_23252,N_23202);
nand U23549 (N_23549,N_23385,N_23353);
xor U23550 (N_23550,N_23275,N_23206);
nand U23551 (N_23551,N_23224,N_23391);
and U23552 (N_23552,N_23224,N_23261);
xnor U23553 (N_23553,N_23362,N_23314);
xnor U23554 (N_23554,N_23370,N_23357);
xor U23555 (N_23555,N_23213,N_23384);
xnor U23556 (N_23556,N_23341,N_23377);
xnor U23557 (N_23557,N_23247,N_23331);
and U23558 (N_23558,N_23206,N_23254);
nor U23559 (N_23559,N_23300,N_23369);
or U23560 (N_23560,N_23276,N_23227);
nand U23561 (N_23561,N_23265,N_23220);
xor U23562 (N_23562,N_23244,N_23227);
xor U23563 (N_23563,N_23341,N_23364);
xor U23564 (N_23564,N_23204,N_23370);
or U23565 (N_23565,N_23264,N_23200);
nor U23566 (N_23566,N_23319,N_23248);
and U23567 (N_23567,N_23382,N_23280);
or U23568 (N_23568,N_23326,N_23300);
xor U23569 (N_23569,N_23217,N_23379);
xor U23570 (N_23570,N_23371,N_23265);
and U23571 (N_23571,N_23349,N_23236);
and U23572 (N_23572,N_23273,N_23345);
nor U23573 (N_23573,N_23234,N_23379);
or U23574 (N_23574,N_23276,N_23259);
and U23575 (N_23575,N_23303,N_23214);
and U23576 (N_23576,N_23392,N_23379);
xor U23577 (N_23577,N_23337,N_23355);
or U23578 (N_23578,N_23380,N_23211);
nor U23579 (N_23579,N_23204,N_23300);
nand U23580 (N_23580,N_23384,N_23266);
nor U23581 (N_23581,N_23272,N_23289);
nand U23582 (N_23582,N_23280,N_23372);
xnor U23583 (N_23583,N_23243,N_23363);
xnor U23584 (N_23584,N_23229,N_23262);
nand U23585 (N_23585,N_23221,N_23289);
or U23586 (N_23586,N_23389,N_23336);
xnor U23587 (N_23587,N_23251,N_23288);
nand U23588 (N_23588,N_23366,N_23363);
nor U23589 (N_23589,N_23325,N_23233);
xor U23590 (N_23590,N_23230,N_23343);
nand U23591 (N_23591,N_23289,N_23385);
nand U23592 (N_23592,N_23377,N_23239);
and U23593 (N_23593,N_23343,N_23200);
xnor U23594 (N_23594,N_23357,N_23204);
and U23595 (N_23595,N_23372,N_23282);
or U23596 (N_23596,N_23360,N_23345);
xnor U23597 (N_23597,N_23312,N_23322);
nor U23598 (N_23598,N_23229,N_23336);
or U23599 (N_23599,N_23247,N_23229);
xnor U23600 (N_23600,N_23431,N_23570);
xor U23601 (N_23601,N_23509,N_23413);
xor U23602 (N_23602,N_23411,N_23457);
and U23603 (N_23603,N_23502,N_23586);
or U23604 (N_23604,N_23451,N_23418);
or U23605 (N_23605,N_23430,N_23475);
nor U23606 (N_23606,N_23404,N_23565);
nor U23607 (N_23607,N_23455,N_23529);
nor U23608 (N_23608,N_23452,N_23467);
xor U23609 (N_23609,N_23463,N_23528);
or U23610 (N_23610,N_23567,N_23426);
nor U23611 (N_23611,N_23414,N_23523);
nand U23612 (N_23612,N_23585,N_23563);
and U23613 (N_23613,N_23532,N_23485);
nand U23614 (N_23614,N_23416,N_23560);
and U23615 (N_23615,N_23590,N_23425);
or U23616 (N_23616,N_23423,N_23427);
nand U23617 (N_23617,N_23556,N_23544);
or U23618 (N_23618,N_23496,N_23526);
or U23619 (N_23619,N_23410,N_23437);
nor U23620 (N_23620,N_23534,N_23454);
nor U23621 (N_23621,N_23512,N_23491);
nor U23622 (N_23622,N_23549,N_23595);
nor U23623 (N_23623,N_23494,N_23504);
and U23624 (N_23624,N_23486,N_23447);
nand U23625 (N_23625,N_23478,N_23555);
xnor U23626 (N_23626,N_23472,N_23568);
and U23627 (N_23627,N_23546,N_23522);
nor U23628 (N_23628,N_23453,N_23539);
xor U23629 (N_23629,N_23434,N_23547);
xor U23630 (N_23630,N_23446,N_23481);
nor U23631 (N_23631,N_23442,N_23541);
nand U23632 (N_23632,N_23444,N_23507);
and U23633 (N_23633,N_23591,N_23543);
nor U23634 (N_23634,N_23422,N_23436);
nor U23635 (N_23635,N_23592,N_23476);
nor U23636 (N_23636,N_23510,N_23545);
nor U23637 (N_23637,N_23443,N_23593);
and U23638 (N_23638,N_23530,N_23578);
nand U23639 (N_23639,N_23503,N_23515);
and U23640 (N_23640,N_23493,N_23465);
xor U23641 (N_23641,N_23456,N_23401);
nand U23642 (N_23642,N_23571,N_23459);
and U23643 (N_23643,N_23407,N_23484);
or U23644 (N_23644,N_23524,N_23561);
xor U23645 (N_23645,N_23582,N_23458);
xnor U23646 (N_23646,N_23554,N_23576);
and U23647 (N_23647,N_23462,N_23506);
xnor U23648 (N_23648,N_23428,N_23400);
nor U23649 (N_23649,N_23473,N_23406);
nand U23650 (N_23650,N_23559,N_23588);
nand U23651 (N_23651,N_23402,N_23552);
nor U23652 (N_23652,N_23572,N_23489);
or U23653 (N_23653,N_23490,N_23516);
or U23654 (N_23654,N_23538,N_23533);
and U23655 (N_23655,N_23548,N_23566);
and U23656 (N_23656,N_23558,N_23421);
or U23657 (N_23657,N_23517,N_23470);
and U23658 (N_23658,N_23403,N_23450);
nor U23659 (N_23659,N_23508,N_23540);
xor U23660 (N_23660,N_23488,N_23464);
xor U23661 (N_23661,N_23580,N_23574);
nand U23662 (N_23662,N_23468,N_23520);
or U23663 (N_23663,N_23519,N_23594);
xnor U23664 (N_23664,N_23477,N_23492);
and U23665 (N_23665,N_23439,N_23438);
or U23666 (N_23666,N_23500,N_23527);
nor U23667 (N_23667,N_23495,N_23584);
nand U23668 (N_23668,N_23483,N_23579);
xor U23669 (N_23669,N_23461,N_23435);
nand U23670 (N_23670,N_23564,N_23497);
or U23671 (N_23671,N_23408,N_23531);
or U23672 (N_23672,N_23424,N_23525);
or U23673 (N_23673,N_23599,N_23445);
and U23674 (N_23674,N_23537,N_23535);
and U23675 (N_23675,N_23513,N_23511);
xor U23676 (N_23676,N_23419,N_23405);
nor U23677 (N_23677,N_23432,N_23448);
nor U23678 (N_23678,N_23440,N_23553);
xnor U23679 (N_23679,N_23521,N_23460);
xnor U23680 (N_23680,N_23589,N_23542);
nor U23681 (N_23681,N_23596,N_23597);
nand U23682 (N_23682,N_23518,N_23420);
nor U23683 (N_23683,N_23536,N_23581);
or U23684 (N_23684,N_23429,N_23412);
nor U23685 (N_23685,N_23409,N_23550);
and U23686 (N_23686,N_23449,N_23577);
nor U23687 (N_23687,N_23487,N_23469);
xor U23688 (N_23688,N_23562,N_23498);
or U23689 (N_23689,N_23415,N_23501);
or U23690 (N_23690,N_23557,N_23569);
nor U23691 (N_23691,N_23583,N_23499);
nand U23692 (N_23692,N_23573,N_23514);
nand U23693 (N_23693,N_23474,N_23480);
nand U23694 (N_23694,N_23471,N_23441);
or U23695 (N_23695,N_23482,N_23598);
xor U23696 (N_23696,N_23466,N_23587);
or U23697 (N_23697,N_23505,N_23417);
nand U23698 (N_23698,N_23551,N_23479);
nand U23699 (N_23699,N_23575,N_23433);
and U23700 (N_23700,N_23560,N_23520);
or U23701 (N_23701,N_23515,N_23553);
and U23702 (N_23702,N_23523,N_23570);
and U23703 (N_23703,N_23479,N_23515);
xor U23704 (N_23704,N_23581,N_23516);
or U23705 (N_23705,N_23489,N_23494);
and U23706 (N_23706,N_23515,N_23451);
nand U23707 (N_23707,N_23403,N_23485);
xnor U23708 (N_23708,N_23567,N_23434);
and U23709 (N_23709,N_23475,N_23445);
xnor U23710 (N_23710,N_23466,N_23592);
nand U23711 (N_23711,N_23465,N_23548);
xor U23712 (N_23712,N_23453,N_23452);
nor U23713 (N_23713,N_23504,N_23585);
and U23714 (N_23714,N_23489,N_23490);
xnor U23715 (N_23715,N_23569,N_23475);
nand U23716 (N_23716,N_23460,N_23530);
or U23717 (N_23717,N_23565,N_23489);
or U23718 (N_23718,N_23480,N_23590);
nor U23719 (N_23719,N_23597,N_23593);
or U23720 (N_23720,N_23518,N_23563);
nand U23721 (N_23721,N_23426,N_23497);
and U23722 (N_23722,N_23406,N_23408);
and U23723 (N_23723,N_23571,N_23400);
xnor U23724 (N_23724,N_23590,N_23500);
nand U23725 (N_23725,N_23443,N_23563);
nor U23726 (N_23726,N_23449,N_23580);
and U23727 (N_23727,N_23419,N_23572);
nand U23728 (N_23728,N_23502,N_23408);
and U23729 (N_23729,N_23576,N_23592);
nand U23730 (N_23730,N_23531,N_23433);
and U23731 (N_23731,N_23486,N_23549);
or U23732 (N_23732,N_23440,N_23525);
or U23733 (N_23733,N_23448,N_23592);
nand U23734 (N_23734,N_23460,N_23579);
xnor U23735 (N_23735,N_23533,N_23510);
nor U23736 (N_23736,N_23441,N_23458);
xor U23737 (N_23737,N_23558,N_23516);
or U23738 (N_23738,N_23577,N_23494);
and U23739 (N_23739,N_23499,N_23465);
nand U23740 (N_23740,N_23525,N_23589);
xnor U23741 (N_23741,N_23488,N_23462);
and U23742 (N_23742,N_23450,N_23436);
or U23743 (N_23743,N_23492,N_23415);
nor U23744 (N_23744,N_23501,N_23528);
and U23745 (N_23745,N_23481,N_23585);
nor U23746 (N_23746,N_23449,N_23533);
xnor U23747 (N_23747,N_23588,N_23454);
or U23748 (N_23748,N_23571,N_23449);
or U23749 (N_23749,N_23449,N_23425);
nor U23750 (N_23750,N_23442,N_23551);
nand U23751 (N_23751,N_23465,N_23439);
nor U23752 (N_23752,N_23499,N_23507);
nand U23753 (N_23753,N_23479,N_23423);
and U23754 (N_23754,N_23569,N_23478);
or U23755 (N_23755,N_23510,N_23582);
xor U23756 (N_23756,N_23580,N_23521);
and U23757 (N_23757,N_23531,N_23567);
and U23758 (N_23758,N_23437,N_23540);
nand U23759 (N_23759,N_23463,N_23572);
and U23760 (N_23760,N_23498,N_23424);
or U23761 (N_23761,N_23422,N_23424);
nand U23762 (N_23762,N_23466,N_23590);
nor U23763 (N_23763,N_23551,N_23410);
xnor U23764 (N_23764,N_23595,N_23427);
nor U23765 (N_23765,N_23497,N_23507);
nand U23766 (N_23766,N_23492,N_23430);
and U23767 (N_23767,N_23525,N_23404);
xor U23768 (N_23768,N_23514,N_23577);
nand U23769 (N_23769,N_23549,N_23565);
nand U23770 (N_23770,N_23508,N_23482);
xor U23771 (N_23771,N_23525,N_23537);
xor U23772 (N_23772,N_23415,N_23499);
nand U23773 (N_23773,N_23551,N_23449);
nand U23774 (N_23774,N_23443,N_23578);
or U23775 (N_23775,N_23487,N_23545);
and U23776 (N_23776,N_23461,N_23471);
xor U23777 (N_23777,N_23575,N_23459);
xor U23778 (N_23778,N_23522,N_23425);
nor U23779 (N_23779,N_23445,N_23490);
and U23780 (N_23780,N_23432,N_23487);
and U23781 (N_23781,N_23526,N_23439);
and U23782 (N_23782,N_23495,N_23462);
xnor U23783 (N_23783,N_23510,N_23570);
or U23784 (N_23784,N_23567,N_23404);
or U23785 (N_23785,N_23408,N_23581);
nand U23786 (N_23786,N_23510,N_23550);
nand U23787 (N_23787,N_23436,N_23459);
nand U23788 (N_23788,N_23559,N_23503);
or U23789 (N_23789,N_23469,N_23405);
or U23790 (N_23790,N_23575,N_23442);
nor U23791 (N_23791,N_23436,N_23578);
and U23792 (N_23792,N_23557,N_23541);
xnor U23793 (N_23793,N_23401,N_23530);
xnor U23794 (N_23794,N_23595,N_23409);
or U23795 (N_23795,N_23531,N_23513);
or U23796 (N_23796,N_23575,N_23443);
nand U23797 (N_23797,N_23526,N_23499);
xnor U23798 (N_23798,N_23550,N_23513);
or U23799 (N_23799,N_23445,N_23579);
nor U23800 (N_23800,N_23633,N_23747);
nand U23801 (N_23801,N_23705,N_23613);
and U23802 (N_23802,N_23664,N_23715);
nor U23803 (N_23803,N_23791,N_23762);
or U23804 (N_23804,N_23711,N_23646);
and U23805 (N_23805,N_23757,N_23778);
or U23806 (N_23806,N_23656,N_23730);
nor U23807 (N_23807,N_23652,N_23643);
nand U23808 (N_23808,N_23692,N_23752);
nand U23809 (N_23809,N_23693,N_23708);
and U23810 (N_23810,N_23668,N_23707);
xnor U23811 (N_23811,N_23663,N_23623);
or U23812 (N_23812,N_23769,N_23601);
and U23813 (N_23813,N_23777,N_23756);
or U23814 (N_23814,N_23694,N_23661);
or U23815 (N_23815,N_23699,N_23726);
or U23816 (N_23816,N_23712,N_23700);
xor U23817 (N_23817,N_23758,N_23706);
and U23818 (N_23818,N_23654,N_23689);
and U23819 (N_23819,N_23723,N_23716);
or U23820 (N_23820,N_23790,N_23625);
nor U23821 (N_23821,N_23722,N_23690);
nand U23822 (N_23822,N_23767,N_23657);
or U23823 (N_23823,N_23640,N_23627);
and U23824 (N_23824,N_23717,N_23616);
nor U23825 (N_23825,N_23610,N_23660);
nor U23826 (N_23826,N_23638,N_23776);
or U23827 (N_23827,N_23766,N_23788);
xor U23828 (N_23828,N_23658,N_23732);
nand U23829 (N_23829,N_23780,N_23600);
and U23830 (N_23830,N_23754,N_23686);
and U23831 (N_23831,N_23739,N_23650);
nand U23832 (N_23832,N_23795,N_23743);
nand U23833 (N_23833,N_23615,N_23630);
nor U23834 (N_23834,N_23786,N_23796);
nand U23835 (N_23835,N_23751,N_23704);
or U23836 (N_23836,N_23644,N_23683);
nor U23837 (N_23837,N_23634,N_23682);
or U23838 (N_23838,N_23685,N_23679);
nand U23839 (N_23839,N_23608,N_23612);
xor U23840 (N_23840,N_23669,N_23617);
nor U23841 (N_23841,N_23763,N_23742);
nand U23842 (N_23842,N_23621,N_23622);
xnor U23843 (N_23843,N_23714,N_23659);
xnor U23844 (N_23844,N_23604,N_23798);
and U23845 (N_23845,N_23701,N_23727);
nor U23846 (N_23846,N_23632,N_23680);
or U23847 (N_23847,N_23635,N_23792);
nor U23848 (N_23848,N_23748,N_23768);
nand U23849 (N_23849,N_23611,N_23698);
or U23850 (N_23850,N_23741,N_23606);
or U23851 (N_23851,N_23744,N_23785);
and U23852 (N_23852,N_23603,N_23740);
nor U23853 (N_23853,N_23696,N_23728);
or U23854 (N_23854,N_23651,N_23746);
xnor U23855 (N_23855,N_23653,N_23691);
nand U23856 (N_23856,N_23670,N_23662);
and U23857 (N_23857,N_23614,N_23789);
and U23858 (N_23858,N_23667,N_23710);
and U23859 (N_23859,N_23733,N_23772);
nor U23860 (N_23860,N_23794,N_23695);
xnor U23861 (N_23861,N_23721,N_23775);
nand U23862 (N_23862,N_23645,N_23703);
or U23863 (N_23863,N_23771,N_23677);
nor U23864 (N_23864,N_23799,N_23782);
nor U23865 (N_23865,N_23750,N_23639);
and U23866 (N_23866,N_23647,N_23773);
xor U23867 (N_23867,N_23655,N_23760);
and U23868 (N_23868,N_23781,N_23678);
and U23869 (N_23869,N_23618,N_23675);
or U23870 (N_23870,N_23620,N_23783);
and U23871 (N_23871,N_23672,N_23605);
xnor U23872 (N_23872,N_23665,N_23697);
xnor U23873 (N_23873,N_23666,N_23641);
xor U23874 (N_23874,N_23749,N_23734);
nand U23875 (N_23875,N_23718,N_23629);
or U23876 (N_23876,N_23779,N_23628);
nor U23877 (N_23877,N_23671,N_23607);
nor U23878 (N_23878,N_23753,N_23761);
nor U23879 (N_23879,N_23736,N_23745);
xnor U23880 (N_23880,N_23725,N_23764);
or U23881 (N_23881,N_23702,N_23713);
xor U23882 (N_23882,N_23637,N_23684);
or U23883 (N_23883,N_23793,N_23649);
and U23884 (N_23884,N_23674,N_23774);
and U23885 (N_23885,N_23648,N_23735);
and U23886 (N_23886,N_23784,N_23642);
nor U23887 (N_23887,N_23737,N_23676);
or U23888 (N_23888,N_23765,N_23729);
xnor U23889 (N_23889,N_23631,N_23624);
nand U23890 (N_23890,N_23759,N_23719);
nor U23891 (N_23891,N_23681,N_23770);
and U23892 (N_23892,N_23731,N_23797);
nand U23893 (N_23893,N_23738,N_23687);
nor U23894 (N_23894,N_23787,N_23609);
nor U23895 (N_23895,N_23720,N_23636);
xnor U23896 (N_23896,N_23673,N_23724);
xnor U23897 (N_23897,N_23619,N_23709);
xor U23898 (N_23898,N_23688,N_23602);
nor U23899 (N_23899,N_23755,N_23626);
xnor U23900 (N_23900,N_23761,N_23651);
or U23901 (N_23901,N_23723,N_23747);
and U23902 (N_23902,N_23740,N_23636);
nand U23903 (N_23903,N_23731,N_23633);
nand U23904 (N_23904,N_23678,N_23732);
nand U23905 (N_23905,N_23707,N_23736);
nor U23906 (N_23906,N_23749,N_23628);
nand U23907 (N_23907,N_23656,N_23625);
or U23908 (N_23908,N_23767,N_23678);
and U23909 (N_23909,N_23767,N_23736);
and U23910 (N_23910,N_23710,N_23644);
nor U23911 (N_23911,N_23700,N_23685);
or U23912 (N_23912,N_23757,N_23632);
nor U23913 (N_23913,N_23602,N_23742);
and U23914 (N_23914,N_23784,N_23694);
or U23915 (N_23915,N_23753,N_23697);
nand U23916 (N_23916,N_23630,N_23739);
and U23917 (N_23917,N_23695,N_23680);
xor U23918 (N_23918,N_23686,N_23646);
xnor U23919 (N_23919,N_23635,N_23620);
nand U23920 (N_23920,N_23687,N_23752);
nand U23921 (N_23921,N_23617,N_23722);
xnor U23922 (N_23922,N_23621,N_23648);
nor U23923 (N_23923,N_23782,N_23746);
or U23924 (N_23924,N_23668,N_23617);
xnor U23925 (N_23925,N_23605,N_23794);
nand U23926 (N_23926,N_23647,N_23775);
and U23927 (N_23927,N_23620,N_23679);
and U23928 (N_23928,N_23673,N_23689);
and U23929 (N_23929,N_23662,N_23747);
xnor U23930 (N_23930,N_23753,N_23737);
nand U23931 (N_23931,N_23655,N_23634);
xor U23932 (N_23932,N_23651,N_23618);
or U23933 (N_23933,N_23718,N_23686);
and U23934 (N_23934,N_23621,N_23752);
or U23935 (N_23935,N_23717,N_23721);
nand U23936 (N_23936,N_23798,N_23765);
or U23937 (N_23937,N_23764,N_23698);
and U23938 (N_23938,N_23761,N_23656);
nor U23939 (N_23939,N_23702,N_23680);
or U23940 (N_23940,N_23692,N_23718);
nor U23941 (N_23941,N_23601,N_23668);
nor U23942 (N_23942,N_23712,N_23755);
and U23943 (N_23943,N_23669,N_23631);
and U23944 (N_23944,N_23643,N_23694);
or U23945 (N_23945,N_23646,N_23621);
xnor U23946 (N_23946,N_23768,N_23636);
or U23947 (N_23947,N_23799,N_23747);
nand U23948 (N_23948,N_23731,N_23652);
xnor U23949 (N_23949,N_23616,N_23755);
nor U23950 (N_23950,N_23733,N_23796);
or U23951 (N_23951,N_23758,N_23686);
nor U23952 (N_23952,N_23708,N_23776);
and U23953 (N_23953,N_23767,N_23625);
or U23954 (N_23954,N_23703,N_23705);
and U23955 (N_23955,N_23685,N_23619);
nand U23956 (N_23956,N_23687,N_23659);
nor U23957 (N_23957,N_23614,N_23703);
nor U23958 (N_23958,N_23781,N_23771);
nor U23959 (N_23959,N_23653,N_23645);
nor U23960 (N_23960,N_23666,N_23629);
nand U23961 (N_23961,N_23630,N_23643);
nor U23962 (N_23962,N_23772,N_23638);
xor U23963 (N_23963,N_23775,N_23789);
or U23964 (N_23964,N_23620,N_23756);
nor U23965 (N_23965,N_23709,N_23688);
or U23966 (N_23966,N_23759,N_23767);
xor U23967 (N_23967,N_23668,N_23644);
or U23968 (N_23968,N_23611,N_23725);
nor U23969 (N_23969,N_23651,N_23715);
and U23970 (N_23970,N_23776,N_23706);
and U23971 (N_23971,N_23660,N_23705);
nand U23972 (N_23972,N_23790,N_23711);
or U23973 (N_23973,N_23788,N_23609);
nor U23974 (N_23974,N_23764,N_23783);
nor U23975 (N_23975,N_23723,N_23776);
or U23976 (N_23976,N_23683,N_23696);
or U23977 (N_23977,N_23710,N_23662);
nand U23978 (N_23978,N_23762,N_23649);
or U23979 (N_23979,N_23783,N_23794);
nor U23980 (N_23980,N_23787,N_23611);
nand U23981 (N_23981,N_23720,N_23604);
nor U23982 (N_23982,N_23600,N_23793);
or U23983 (N_23983,N_23722,N_23755);
nor U23984 (N_23984,N_23623,N_23755);
or U23985 (N_23985,N_23778,N_23726);
and U23986 (N_23986,N_23704,N_23730);
nand U23987 (N_23987,N_23692,N_23646);
and U23988 (N_23988,N_23770,N_23793);
or U23989 (N_23989,N_23796,N_23790);
and U23990 (N_23990,N_23603,N_23787);
xnor U23991 (N_23991,N_23681,N_23724);
nand U23992 (N_23992,N_23733,N_23664);
or U23993 (N_23993,N_23704,N_23633);
and U23994 (N_23994,N_23616,N_23649);
nor U23995 (N_23995,N_23718,N_23658);
nand U23996 (N_23996,N_23771,N_23696);
or U23997 (N_23997,N_23608,N_23758);
or U23998 (N_23998,N_23670,N_23687);
nand U23999 (N_23999,N_23601,N_23649);
nand U24000 (N_24000,N_23852,N_23820);
and U24001 (N_24001,N_23802,N_23805);
xor U24002 (N_24002,N_23971,N_23981);
and U24003 (N_24003,N_23972,N_23869);
or U24004 (N_24004,N_23834,N_23988);
nand U24005 (N_24005,N_23855,N_23979);
xor U24006 (N_24006,N_23922,N_23843);
nor U24007 (N_24007,N_23806,N_23880);
nand U24008 (N_24008,N_23929,N_23889);
xnor U24009 (N_24009,N_23903,N_23887);
nand U24010 (N_24010,N_23870,N_23910);
nor U24011 (N_24011,N_23914,N_23876);
and U24012 (N_24012,N_23808,N_23909);
or U24013 (N_24013,N_23949,N_23959);
or U24014 (N_24014,N_23882,N_23915);
nor U24015 (N_24015,N_23803,N_23958);
nor U24016 (N_24016,N_23984,N_23968);
xnor U24017 (N_24017,N_23800,N_23995);
and U24018 (N_24018,N_23867,N_23854);
xor U24019 (N_24019,N_23819,N_23895);
nor U24020 (N_24020,N_23899,N_23923);
nor U24021 (N_24021,N_23823,N_23948);
nor U24022 (N_24022,N_23841,N_23935);
xnor U24023 (N_24023,N_23845,N_23828);
and U24024 (N_24024,N_23991,N_23954);
or U24025 (N_24025,N_23875,N_23973);
xor U24026 (N_24026,N_23842,N_23838);
nand U24027 (N_24027,N_23977,N_23985);
nand U24028 (N_24028,N_23893,N_23975);
nand U24029 (N_24029,N_23941,N_23918);
and U24030 (N_24030,N_23898,N_23822);
nand U24031 (N_24031,N_23927,N_23864);
xor U24032 (N_24032,N_23992,N_23886);
or U24033 (N_24033,N_23900,N_23811);
nor U24034 (N_24034,N_23916,N_23964);
nor U24035 (N_24035,N_23976,N_23891);
xnor U24036 (N_24036,N_23969,N_23963);
and U24037 (N_24037,N_23908,N_23860);
nand U24038 (N_24038,N_23919,N_23833);
nor U24039 (N_24039,N_23917,N_23962);
nor U24040 (N_24040,N_23944,N_23846);
or U24041 (N_24041,N_23937,N_23868);
xor U24042 (N_24042,N_23950,N_23814);
xnor U24043 (N_24043,N_23826,N_23844);
xor U24044 (N_24044,N_23990,N_23866);
and U24045 (N_24045,N_23955,N_23982);
nor U24046 (N_24046,N_23983,N_23965);
nand U24047 (N_24047,N_23804,N_23938);
nor U24048 (N_24048,N_23980,N_23871);
xor U24049 (N_24049,N_23809,N_23851);
or U24050 (N_24050,N_23862,N_23815);
nor U24051 (N_24051,N_23863,N_23832);
xor U24052 (N_24052,N_23943,N_23865);
or U24053 (N_24053,N_23890,N_23897);
xor U24054 (N_24054,N_23881,N_23896);
nor U24055 (N_24055,N_23961,N_23997);
and U24056 (N_24056,N_23974,N_23928);
nand U24057 (N_24057,N_23831,N_23966);
and U24058 (N_24058,N_23926,N_23952);
or U24059 (N_24059,N_23970,N_23993);
and U24060 (N_24060,N_23836,N_23840);
and U24061 (N_24061,N_23946,N_23945);
nand U24062 (N_24062,N_23829,N_23932);
nor U24063 (N_24063,N_23861,N_23857);
nor U24064 (N_24064,N_23920,N_23999);
and U24065 (N_24065,N_23807,N_23942);
xor U24066 (N_24066,N_23879,N_23883);
or U24067 (N_24067,N_23878,N_23853);
and U24068 (N_24068,N_23902,N_23872);
or U24069 (N_24069,N_23939,N_23930);
xnor U24070 (N_24070,N_23885,N_23894);
nand U24071 (N_24071,N_23824,N_23818);
and U24072 (N_24072,N_23913,N_23986);
and U24073 (N_24073,N_23934,N_23940);
and U24074 (N_24074,N_23904,N_23956);
or U24075 (N_24075,N_23839,N_23801);
or U24076 (N_24076,N_23936,N_23996);
xor U24077 (N_24077,N_23837,N_23877);
xor U24078 (N_24078,N_23989,N_23957);
and U24079 (N_24079,N_23933,N_23888);
or U24080 (N_24080,N_23827,N_23812);
and U24081 (N_24081,N_23987,N_23912);
and U24082 (N_24082,N_23884,N_23931);
nor U24083 (N_24083,N_23924,N_23911);
or U24084 (N_24084,N_23817,N_23998);
nor U24085 (N_24085,N_23830,N_23813);
and U24086 (N_24086,N_23921,N_23849);
and U24087 (N_24087,N_23848,N_23873);
nand U24088 (N_24088,N_23906,N_23947);
nand U24089 (N_24089,N_23858,N_23978);
and U24090 (N_24090,N_23994,N_23953);
or U24091 (N_24091,N_23825,N_23907);
nor U24092 (N_24092,N_23951,N_23850);
nand U24093 (N_24093,N_23821,N_23892);
xor U24094 (N_24094,N_23847,N_23874);
xnor U24095 (N_24095,N_23859,N_23835);
nand U24096 (N_24096,N_23925,N_23810);
nand U24097 (N_24097,N_23960,N_23816);
or U24098 (N_24098,N_23905,N_23967);
nand U24099 (N_24099,N_23901,N_23856);
and U24100 (N_24100,N_23880,N_23960);
and U24101 (N_24101,N_23825,N_23807);
or U24102 (N_24102,N_23878,N_23914);
or U24103 (N_24103,N_23870,N_23837);
and U24104 (N_24104,N_23836,N_23976);
and U24105 (N_24105,N_23977,N_23949);
xor U24106 (N_24106,N_23939,N_23819);
nand U24107 (N_24107,N_23877,N_23996);
xnor U24108 (N_24108,N_23885,N_23944);
xnor U24109 (N_24109,N_23903,N_23897);
or U24110 (N_24110,N_23830,N_23873);
nand U24111 (N_24111,N_23876,N_23894);
nand U24112 (N_24112,N_23806,N_23996);
or U24113 (N_24113,N_23990,N_23910);
nor U24114 (N_24114,N_23825,N_23951);
xnor U24115 (N_24115,N_23988,N_23835);
and U24116 (N_24116,N_23929,N_23887);
nor U24117 (N_24117,N_23907,N_23999);
xor U24118 (N_24118,N_23972,N_23812);
nand U24119 (N_24119,N_23861,N_23915);
and U24120 (N_24120,N_23965,N_23964);
and U24121 (N_24121,N_23836,N_23923);
and U24122 (N_24122,N_23993,N_23991);
or U24123 (N_24123,N_23878,N_23991);
nor U24124 (N_24124,N_23901,N_23921);
and U24125 (N_24125,N_23802,N_23888);
nand U24126 (N_24126,N_23877,N_23826);
and U24127 (N_24127,N_23985,N_23872);
nand U24128 (N_24128,N_23956,N_23975);
and U24129 (N_24129,N_23858,N_23939);
and U24130 (N_24130,N_23943,N_23873);
and U24131 (N_24131,N_23888,N_23983);
nor U24132 (N_24132,N_23959,N_23941);
nor U24133 (N_24133,N_23808,N_23832);
xor U24134 (N_24134,N_23845,N_23863);
nand U24135 (N_24135,N_23981,N_23939);
nor U24136 (N_24136,N_23919,N_23981);
xnor U24137 (N_24137,N_23933,N_23806);
xnor U24138 (N_24138,N_23932,N_23832);
xnor U24139 (N_24139,N_23954,N_23935);
and U24140 (N_24140,N_23861,N_23887);
nand U24141 (N_24141,N_23831,N_23852);
or U24142 (N_24142,N_23819,N_23838);
or U24143 (N_24143,N_23858,N_23965);
and U24144 (N_24144,N_23846,N_23900);
and U24145 (N_24145,N_23943,N_23886);
nand U24146 (N_24146,N_23930,N_23808);
or U24147 (N_24147,N_23892,N_23844);
nor U24148 (N_24148,N_23849,N_23837);
xnor U24149 (N_24149,N_23884,N_23983);
or U24150 (N_24150,N_23934,N_23985);
xnor U24151 (N_24151,N_23859,N_23850);
nor U24152 (N_24152,N_23878,N_23974);
and U24153 (N_24153,N_23934,N_23978);
or U24154 (N_24154,N_23968,N_23879);
xnor U24155 (N_24155,N_23944,N_23824);
nand U24156 (N_24156,N_23822,N_23846);
nor U24157 (N_24157,N_23842,N_23913);
xnor U24158 (N_24158,N_23969,N_23863);
nor U24159 (N_24159,N_23936,N_23934);
or U24160 (N_24160,N_23961,N_23871);
nand U24161 (N_24161,N_23936,N_23927);
nand U24162 (N_24162,N_23922,N_23906);
nand U24163 (N_24163,N_23958,N_23887);
nor U24164 (N_24164,N_23991,N_23836);
nand U24165 (N_24165,N_23869,N_23802);
and U24166 (N_24166,N_23974,N_23964);
and U24167 (N_24167,N_23853,N_23874);
or U24168 (N_24168,N_23876,N_23849);
nand U24169 (N_24169,N_23857,N_23837);
or U24170 (N_24170,N_23980,N_23827);
nand U24171 (N_24171,N_23857,N_23860);
and U24172 (N_24172,N_23900,N_23804);
nor U24173 (N_24173,N_23979,N_23836);
nor U24174 (N_24174,N_23927,N_23818);
nand U24175 (N_24175,N_23902,N_23838);
nor U24176 (N_24176,N_23903,N_23806);
xnor U24177 (N_24177,N_23952,N_23944);
nor U24178 (N_24178,N_23949,N_23901);
xor U24179 (N_24179,N_23892,N_23867);
nor U24180 (N_24180,N_23968,N_23812);
and U24181 (N_24181,N_23884,N_23835);
xor U24182 (N_24182,N_23825,N_23940);
and U24183 (N_24183,N_23818,N_23890);
or U24184 (N_24184,N_23922,N_23862);
or U24185 (N_24185,N_23931,N_23823);
or U24186 (N_24186,N_23914,N_23854);
xor U24187 (N_24187,N_23814,N_23972);
nor U24188 (N_24188,N_23964,N_23890);
xor U24189 (N_24189,N_23856,N_23820);
nand U24190 (N_24190,N_23912,N_23856);
and U24191 (N_24191,N_23937,N_23925);
nor U24192 (N_24192,N_23855,N_23869);
and U24193 (N_24193,N_23843,N_23887);
xnor U24194 (N_24194,N_23923,N_23964);
and U24195 (N_24195,N_23872,N_23914);
nand U24196 (N_24196,N_23890,N_23945);
xor U24197 (N_24197,N_23996,N_23953);
and U24198 (N_24198,N_23900,N_23859);
nand U24199 (N_24199,N_23807,N_23949);
nand U24200 (N_24200,N_24061,N_24181);
xnor U24201 (N_24201,N_24052,N_24188);
nor U24202 (N_24202,N_24159,N_24079);
nor U24203 (N_24203,N_24161,N_24149);
nor U24204 (N_24204,N_24105,N_24048);
nor U24205 (N_24205,N_24176,N_24186);
or U24206 (N_24206,N_24035,N_24196);
and U24207 (N_24207,N_24021,N_24171);
and U24208 (N_24208,N_24045,N_24099);
and U24209 (N_24209,N_24066,N_24053);
or U24210 (N_24210,N_24123,N_24110);
or U24211 (N_24211,N_24015,N_24025);
and U24212 (N_24212,N_24094,N_24147);
xnor U24213 (N_24213,N_24141,N_24013);
nand U24214 (N_24214,N_24194,N_24116);
or U24215 (N_24215,N_24150,N_24100);
and U24216 (N_24216,N_24151,N_24117);
and U24217 (N_24217,N_24114,N_24104);
xnor U24218 (N_24218,N_24132,N_24006);
xnor U24219 (N_24219,N_24014,N_24042);
nand U24220 (N_24220,N_24070,N_24135);
nand U24221 (N_24221,N_24091,N_24072);
xnor U24222 (N_24222,N_24184,N_24000);
or U24223 (N_24223,N_24074,N_24189);
or U24224 (N_24224,N_24156,N_24098);
or U24225 (N_24225,N_24001,N_24131);
nand U24226 (N_24226,N_24038,N_24122);
xor U24227 (N_24227,N_24043,N_24080);
nor U24228 (N_24228,N_24071,N_24027);
or U24229 (N_24229,N_24033,N_24167);
xnor U24230 (N_24230,N_24054,N_24164);
xnor U24231 (N_24231,N_24160,N_24127);
and U24232 (N_24232,N_24046,N_24102);
or U24233 (N_24233,N_24059,N_24157);
and U24234 (N_24234,N_24008,N_24057);
or U24235 (N_24235,N_24185,N_24170);
and U24236 (N_24236,N_24175,N_24113);
nor U24237 (N_24237,N_24005,N_24111);
nor U24238 (N_24238,N_24019,N_24121);
nor U24239 (N_24239,N_24130,N_24183);
nor U24240 (N_24240,N_24044,N_24140);
and U24241 (N_24241,N_24009,N_24036);
nand U24242 (N_24242,N_24050,N_24115);
or U24243 (N_24243,N_24138,N_24085);
or U24244 (N_24244,N_24067,N_24077);
xnor U24245 (N_24245,N_24190,N_24047);
nor U24246 (N_24246,N_24030,N_24172);
and U24247 (N_24247,N_24010,N_24039);
xnor U24248 (N_24248,N_24073,N_24158);
nand U24249 (N_24249,N_24120,N_24118);
and U24250 (N_24250,N_24058,N_24018);
and U24251 (N_24251,N_24197,N_24020);
and U24252 (N_24252,N_24192,N_24016);
or U24253 (N_24253,N_24040,N_24049);
and U24254 (N_24254,N_24125,N_24112);
nand U24255 (N_24255,N_24092,N_24143);
nand U24256 (N_24256,N_24195,N_24056);
or U24257 (N_24257,N_24101,N_24097);
or U24258 (N_24258,N_24083,N_24075);
xor U24259 (N_24259,N_24153,N_24180);
xor U24260 (N_24260,N_24152,N_24031);
or U24261 (N_24261,N_24133,N_24069);
xor U24262 (N_24262,N_24193,N_24041);
nand U24263 (N_24263,N_24166,N_24088);
and U24264 (N_24264,N_24119,N_24032);
nand U24265 (N_24265,N_24003,N_24068);
and U24266 (N_24266,N_24011,N_24109);
or U24267 (N_24267,N_24144,N_24012);
and U24268 (N_24268,N_24162,N_24136);
nor U24269 (N_24269,N_24002,N_24086);
nor U24270 (N_24270,N_24089,N_24022);
nand U24271 (N_24271,N_24024,N_24169);
nor U24272 (N_24272,N_24023,N_24182);
nor U24273 (N_24273,N_24076,N_24096);
or U24274 (N_24274,N_24173,N_24106);
or U24275 (N_24275,N_24017,N_24163);
nor U24276 (N_24276,N_24065,N_24155);
xor U24277 (N_24277,N_24064,N_24051);
nor U24278 (N_24278,N_24093,N_24062);
or U24279 (N_24279,N_24078,N_24145);
nor U24280 (N_24280,N_24142,N_24126);
nor U24281 (N_24281,N_24103,N_24081);
or U24282 (N_24282,N_24082,N_24187);
xnor U24283 (N_24283,N_24139,N_24191);
and U24284 (N_24284,N_24154,N_24004);
and U24285 (N_24285,N_24198,N_24108);
nor U24286 (N_24286,N_24090,N_24178);
nor U24287 (N_24287,N_24034,N_24177);
nor U24288 (N_24288,N_24137,N_24146);
xnor U24289 (N_24289,N_24095,N_24168);
xor U24290 (N_24290,N_24128,N_24037);
nand U24291 (N_24291,N_24028,N_24134);
nand U24292 (N_24292,N_24107,N_24084);
nor U24293 (N_24293,N_24129,N_24060);
nor U24294 (N_24294,N_24199,N_24165);
or U24295 (N_24295,N_24179,N_24007);
xor U24296 (N_24296,N_24124,N_24174);
xor U24297 (N_24297,N_24055,N_24026);
nor U24298 (N_24298,N_24029,N_24087);
nand U24299 (N_24299,N_24063,N_24148);
and U24300 (N_24300,N_24074,N_24039);
and U24301 (N_24301,N_24145,N_24026);
nor U24302 (N_24302,N_24077,N_24099);
nand U24303 (N_24303,N_24104,N_24035);
and U24304 (N_24304,N_24001,N_24193);
and U24305 (N_24305,N_24134,N_24040);
xor U24306 (N_24306,N_24083,N_24114);
nor U24307 (N_24307,N_24125,N_24078);
xor U24308 (N_24308,N_24074,N_24127);
xor U24309 (N_24309,N_24191,N_24008);
or U24310 (N_24310,N_24000,N_24012);
xor U24311 (N_24311,N_24165,N_24056);
and U24312 (N_24312,N_24164,N_24087);
and U24313 (N_24313,N_24100,N_24059);
or U24314 (N_24314,N_24056,N_24150);
nor U24315 (N_24315,N_24000,N_24033);
nor U24316 (N_24316,N_24122,N_24182);
nand U24317 (N_24317,N_24103,N_24036);
and U24318 (N_24318,N_24166,N_24005);
and U24319 (N_24319,N_24063,N_24032);
nand U24320 (N_24320,N_24127,N_24116);
nor U24321 (N_24321,N_24118,N_24030);
and U24322 (N_24322,N_24108,N_24143);
nand U24323 (N_24323,N_24159,N_24125);
nor U24324 (N_24324,N_24069,N_24192);
nand U24325 (N_24325,N_24038,N_24003);
and U24326 (N_24326,N_24153,N_24122);
nand U24327 (N_24327,N_24148,N_24102);
and U24328 (N_24328,N_24150,N_24133);
xor U24329 (N_24329,N_24060,N_24185);
xor U24330 (N_24330,N_24052,N_24109);
and U24331 (N_24331,N_24014,N_24116);
nor U24332 (N_24332,N_24081,N_24037);
or U24333 (N_24333,N_24070,N_24020);
nand U24334 (N_24334,N_24030,N_24009);
xnor U24335 (N_24335,N_24075,N_24120);
and U24336 (N_24336,N_24141,N_24185);
xor U24337 (N_24337,N_24084,N_24174);
xor U24338 (N_24338,N_24066,N_24127);
or U24339 (N_24339,N_24063,N_24162);
and U24340 (N_24340,N_24167,N_24145);
nand U24341 (N_24341,N_24153,N_24137);
nor U24342 (N_24342,N_24006,N_24041);
xnor U24343 (N_24343,N_24155,N_24173);
xnor U24344 (N_24344,N_24052,N_24004);
nor U24345 (N_24345,N_24090,N_24109);
or U24346 (N_24346,N_24194,N_24107);
or U24347 (N_24347,N_24070,N_24187);
nand U24348 (N_24348,N_24085,N_24143);
or U24349 (N_24349,N_24187,N_24175);
or U24350 (N_24350,N_24069,N_24082);
xor U24351 (N_24351,N_24001,N_24022);
nand U24352 (N_24352,N_24124,N_24197);
nand U24353 (N_24353,N_24118,N_24106);
and U24354 (N_24354,N_24168,N_24045);
nand U24355 (N_24355,N_24049,N_24039);
nor U24356 (N_24356,N_24158,N_24070);
nand U24357 (N_24357,N_24016,N_24140);
nor U24358 (N_24358,N_24107,N_24051);
or U24359 (N_24359,N_24083,N_24044);
and U24360 (N_24360,N_24055,N_24112);
xnor U24361 (N_24361,N_24020,N_24061);
nor U24362 (N_24362,N_24133,N_24197);
xor U24363 (N_24363,N_24014,N_24154);
and U24364 (N_24364,N_24037,N_24118);
and U24365 (N_24365,N_24090,N_24122);
nor U24366 (N_24366,N_24058,N_24131);
nor U24367 (N_24367,N_24084,N_24010);
xor U24368 (N_24368,N_24020,N_24189);
or U24369 (N_24369,N_24173,N_24116);
xnor U24370 (N_24370,N_24037,N_24161);
nor U24371 (N_24371,N_24108,N_24017);
nand U24372 (N_24372,N_24101,N_24024);
nand U24373 (N_24373,N_24065,N_24186);
and U24374 (N_24374,N_24007,N_24011);
or U24375 (N_24375,N_24183,N_24100);
and U24376 (N_24376,N_24155,N_24193);
xor U24377 (N_24377,N_24150,N_24160);
or U24378 (N_24378,N_24025,N_24154);
xor U24379 (N_24379,N_24043,N_24109);
or U24380 (N_24380,N_24016,N_24042);
and U24381 (N_24381,N_24167,N_24107);
and U24382 (N_24382,N_24194,N_24042);
or U24383 (N_24383,N_24099,N_24051);
xor U24384 (N_24384,N_24101,N_24019);
nor U24385 (N_24385,N_24071,N_24051);
or U24386 (N_24386,N_24031,N_24153);
or U24387 (N_24387,N_24010,N_24189);
or U24388 (N_24388,N_24070,N_24047);
nand U24389 (N_24389,N_24172,N_24110);
and U24390 (N_24390,N_24007,N_24054);
and U24391 (N_24391,N_24059,N_24191);
xor U24392 (N_24392,N_24106,N_24011);
xnor U24393 (N_24393,N_24074,N_24017);
xnor U24394 (N_24394,N_24050,N_24116);
nor U24395 (N_24395,N_24155,N_24143);
or U24396 (N_24396,N_24023,N_24049);
nand U24397 (N_24397,N_24146,N_24158);
and U24398 (N_24398,N_24133,N_24014);
xnor U24399 (N_24399,N_24154,N_24054);
xor U24400 (N_24400,N_24230,N_24226);
nor U24401 (N_24401,N_24366,N_24255);
or U24402 (N_24402,N_24283,N_24324);
nand U24403 (N_24403,N_24392,N_24209);
xnor U24404 (N_24404,N_24213,N_24218);
nor U24405 (N_24405,N_24374,N_24269);
xor U24406 (N_24406,N_24381,N_24243);
nand U24407 (N_24407,N_24274,N_24389);
nor U24408 (N_24408,N_24211,N_24205);
nor U24409 (N_24409,N_24309,N_24252);
nor U24410 (N_24410,N_24343,N_24233);
nor U24411 (N_24411,N_24360,N_24383);
xnor U24412 (N_24412,N_24350,N_24308);
nand U24413 (N_24413,N_24282,N_24341);
and U24414 (N_24414,N_24317,N_24271);
nor U24415 (N_24415,N_24272,N_24292);
nor U24416 (N_24416,N_24315,N_24219);
xor U24417 (N_24417,N_24367,N_24259);
nor U24418 (N_24418,N_24200,N_24261);
nor U24419 (N_24419,N_24361,N_24300);
nor U24420 (N_24420,N_24298,N_24260);
nand U24421 (N_24421,N_24352,N_24279);
nand U24422 (N_24422,N_24375,N_24202);
or U24423 (N_24423,N_24286,N_24257);
nor U24424 (N_24424,N_24273,N_24370);
xnor U24425 (N_24425,N_24242,N_24345);
and U24426 (N_24426,N_24301,N_24306);
nor U24427 (N_24427,N_24391,N_24371);
or U24428 (N_24428,N_24234,N_24221);
nand U24429 (N_24429,N_24278,N_24354);
nor U24430 (N_24430,N_24364,N_24241);
xor U24431 (N_24431,N_24319,N_24329);
xor U24432 (N_24432,N_24365,N_24254);
or U24433 (N_24433,N_24339,N_24399);
nor U24434 (N_24434,N_24311,N_24206);
and U24435 (N_24435,N_24380,N_24224);
xnor U24436 (N_24436,N_24227,N_24280);
and U24437 (N_24437,N_24330,N_24372);
or U24438 (N_24438,N_24336,N_24346);
nor U24439 (N_24439,N_24288,N_24244);
and U24440 (N_24440,N_24314,N_24238);
or U24441 (N_24441,N_24325,N_24397);
xnor U24442 (N_24442,N_24373,N_24321);
and U24443 (N_24443,N_24327,N_24398);
and U24444 (N_24444,N_24332,N_24348);
or U24445 (N_24445,N_24338,N_24245);
nor U24446 (N_24446,N_24335,N_24236);
or U24447 (N_24447,N_24291,N_24207);
and U24448 (N_24448,N_24220,N_24203);
nand U24449 (N_24449,N_24276,N_24289);
nor U24450 (N_24450,N_24344,N_24384);
or U24451 (N_24451,N_24310,N_24326);
nor U24452 (N_24452,N_24251,N_24322);
and U24453 (N_24453,N_24379,N_24285);
and U24454 (N_24454,N_24299,N_24353);
xor U24455 (N_24455,N_24217,N_24293);
or U24456 (N_24456,N_24256,N_24253);
or U24457 (N_24457,N_24295,N_24393);
or U24458 (N_24458,N_24305,N_24357);
xor U24459 (N_24459,N_24212,N_24201);
or U24460 (N_24460,N_24376,N_24237);
nor U24461 (N_24461,N_24328,N_24263);
or U24462 (N_24462,N_24359,N_24331);
xor U24463 (N_24463,N_24337,N_24268);
nand U24464 (N_24464,N_24264,N_24318);
xnor U24465 (N_24465,N_24216,N_24231);
nand U24466 (N_24466,N_24262,N_24369);
xor U24467 (N_24467,N_24395,N_24316);
or U24468 (N_24468,N_24229,N_24385);
nor U24469 (N_24469,N_24235,N_24304);
and U24470 (N_24470,N_24232,N_24302);
nor U24471 (N_24471,N_24225,N_24362);
nor U24472 (N_24472,N_24281,N_24284);
xnor U24473 (N_24473,N_24208,N_24275);
and U24474 (N_24474,N_24222,N_24333);
xnor U24475 (N_24475,N_24287,N_24340);
nor U24476 (N_24476,N_24390,N_24266);
nor U24477 (N_24477,N_24215,N_24323);
nor U24478 (N_24478,N_24270,N_24277);
nand U24479 (N_24479,N_24210,N_24358);
xnor U24480 (N_24480,N_24355,N_24246);
nand U24481 (N_24481,N_24297,N_24312);
and U24482 (N_24482,N_24267,N_24307);
xnor U24483 (N_24483,N_24377,N_24349);
nor U24484 (N_24484,N_24265,N_24386);
xor U24485 (N_24485,N_24342,N_24258);
xnor U24486 (N_24486,N_24320,N_24356);
nand U24487 (N_24487,N_24250,N_24290);
nor U24488 (N_24488,N_24396,N_24247);
nor U24489 (N_24489,N_24228,N_24296);
or U24490 (N_24490,N_24347,N_24368);
or U24491 (N_24491,N_24214,N_24334);
nand U24492 (N_24492,N_24388,N_24204);
nand U24493 (N_24493,N_24378,N_24313);
nand U24494 (N_24494,N_24351,N_24363);
and U24495 (N_24495,N_24294,N_24303);
and U24496 (N_24496,N_24387,N_24239);
xor U24497 (N_24497,N_24223,N_24249);
nor U24498 (N_24498,N_24248,N_24240);
nand U24499 (N_24499,N_24394,N_24382);
xor U24500 (N_24500,N_24355,N_24352);
xnor U24501 (N_24501,N_24363,N_24280);
nor U24502 (N_24502,N_24255,N_24398);
or U24503 (N_24503,N_24385,N_24213);
nand U24504 (N_24504,N_24367,N_24327);
and U24505 (N_24505,N_24260,N_24297);
or U24506 (N_24506,N_24233,N_24338);
or U24507 (N_24507,N_24345,N_24228);
nor U24508 (N_24508,N_24328,N_24392);
xnor U24509 (N_24509,N_24204,N_24261);
nor U24510 (N_24510,N_24294,N_24229);
xnor U24511 (N_24511,N_24364,N_24328);
xor U24512 (N_24512,N_24323,N_24212);
or U24513 (N_24513,N_24393,N_24293);
nor U24514 (N_24514,N_24250,N_24324);
xor U24515 (N_24515,N_24259,N_24241);
or U24516 (N_24516,N_24395,N_24296);
or U24517 (N_24517,N_24247,N_24325);
or U24518 (N_24518,N_24290,N_24303);
and U24519 (N_24519,N_24259,N_24253);
and U24520 (N_24520,N_24347,N_24247);
nand U24521 (N_24521,N_24269,N_24317);
xnor U24522 (N_24522,N_24282,N_24356);
and U24523 (N_24523,N_24254,N_24321);
or U24524 (N_24524,N_24326,N_24313);
nor U24525 (N_24525,N_24294,N_24355);
or U24526 (N_24526,N_24384,N_24342);
and U24527 (N_24527,N_24278,N_24201);
xor U24528 (N_24528,N_24333,N_24236);
nor U24529 (N_24529,N_24382,N_24360);
nor U24530 (N_24530,N_24346,N_24246);
nand U24531 (N_24531,N_24264,N_24277);
or U24532 (N_24532,N_24345,N_24243);
and U24533 (N_24533,N_24287,N_24371);
xor U24534 (N_24534,N_24218,N_24227);
nand U24535 (N_24535,N_24322,N_24332);
and U24536 (N_24536,N_24382,N_24355);
xor U24537 (N_24537,N_24242,N_24292);
or U24538 (N_24538,N_24294,N_24250);
or U24539 (N_24539,N_24230,N_24356);
xnor U24540 (N_24540,N_24206,N_24275);
nand U24541 (N_24541,N_24206,N_24219);
nand U24542 (N_24542,N_24335,N_24226);
xor U24543 (N_24543,N_24319,N_24362);
or U24544 (N_24544,N_24211,N_24342);
nand U24545 (N_24545,N_24300,N_24235);
nor U24546 (N_24546,N_24209,N_24270);
or U24547 (N_24547,N_24364,N_24204);
nor U24548 (N_24548,N_24348,N_24356);
and U24549 (N_24549,N_24213,N_24316);
and U24550 (N_24550,N_24323,N_24309);
or U24551 (N_24551,N_24264,N_24350);
nand U24552 (N_24552,N_24221,N_24391);
or U24553 (N_24553,N_24387,N_24313);
nor U24554 (N_24554,N_24335,N_24330);
nand U24555 (N_24555,N_24260,N_24232);
and U24556 (N_24556,N_24226,N_24297);
nor U24557 (N_24557,N_24259,N_24378);
nand U24558 (N_24558,N_24215,N_24201);
nand U24559 (N_24559,N_24334,N_24386);
and U24560 (N_24560,N_24271,N_24200);
or U24561 (N_24561,N_24353,N_24336);
and U24562 (N_24562,N_24294,N_24257);
and U24563 (N_24563,N_24336,N_24298);
nand U24564 (N_24564,N_24308,N_24304);
xnor U24565 (N_24565,N_24320,N_24358);
nor U24566 (N_24566,N_24249,N_24310);
and U24567 (N_24567,N_24227,N_24369);
nand U24568 (N_24568,N_24386,N_24211);
xor U24569 (N_24569,N_24329,N_24333);
nand U24570 (N_24570,N_24249,N_24275);
nor U24571 (N_24571,N_24347,N_24321);
or U24572 (N_24572,N_24355,N_24363);
xor U24573 (N_24573,N_24276,N_24253);
or U24574 (N_24574,N_24269,N_24264);
and U24575 (N_24575,N_24373,N_24222);
nor U24576 (N_24576,N_24208,N_24265);
or U24577 (N_24577,N_24223,N_24356);
and U24578 (N_24578,N_24264,N_24283);
and U24579 (N_24579,N_24397,N_24275);
nand U24580 (N_24580,N_24391,N_24204);
and U24581 (N_24581,N_24284,N_24207);
nand U24582 (N_24582,N_24342,N_24311);
nand U24583 (N_24583,N_24258,N_24384);
and U24584 (N_24584,N_24362,N_24303);
and U24585 (N_24585,N_24293,N_24242);
xor U24586 (N_24586,N_24318,N_24279);
nand U24587 (N_24587,N_24382,N_24215);
xor U24588 (N_24588,N_24398,N_24352);
nor U24589 (N_24589,N_24328,N_24296);
and U24590 (N_24590,N_24380,N_24283);
xnor U24591 (N_24591,N_24333,N_24340);
or U24592 (N_24592,N_24328,N_24289);
or U24593 (N_24593,N_24267,N_24329);
nand U24594 (N_24594,N_24234,N_24240);
or U24595 (N_24595,N_24224,N_24325);
or U24596 (N_24596,N_24325,N_24339);
nand U24597 (N_24597,N_24357,N_24297);
nor U24598 (N_24598,N_24226,N_24264);
nand U24599 (N_24599,N_24345,N_24266);
nand U24600 (N_24600,N_24477,N_24457);
and U24601 (N_24601,N_24416,N_24592);
nor U24602 (N_24602,N_24436,N_24489);
or U24603 (N_24603,N_24556,N_24453);
nor U24604 (N_24604,N_24500,N_24469);
and U24605 (N_24605,N_24428,N_24427);
or U24606 (N_24606,N_24462,N_24466);
xnor U24607 (N_24607,N_24508,N_24467);
nand U24608 (N_24608,N_24440,N_24407);
nor U24609 (N_24609,N_24565,N_24578);
or U24610 (N_24610,N_24465,N_24482);
or U24611 (N_24611,N_24569,N_24415);
or U24612 (N_24612,N_24573,N_24577);
and U24613 (N_24613,N_24456,N_24461);
nand U24614 (N_24614,N_24587,N_24505);
xnor U24615 (N_24615,N_24580,N_24591);
nor U24616 (N_24616,N_24563,N_24514);
xnor U24617 (N_24617,N_24485,N_24417);
or U24618 (N_24618,N_24409,N_24546);
or U24619 (N_24619,N_24481,N_24525);
or U24620 (N_24620,N_24455,N_24483);
nor U24621 (N_24621,N_24451,N_24425);
nor U24622 (N_24622,N_24447,N_24501);
and U24623 (N_24623,N_24438,N_24452);
or U24624 (N_24624,N_24499,N_24444);
xnor U24625 (N_24625,N_24566,N_24424);
or U24626 (N_24626,N_24480,N_24537);
xor U24627 (N_24627,N_24534,N_24490);
nor U24628 (N_24628,N_24423,N_24403);
nand U24629 (N_24629,N_24475,N_24479);
nor U24630 (N_24630,N_24406,N_24402);
xor U24631 (N_24631,N_24596,N_24593);
nor U24632 (N_24632,N_24585,N_24581);
nor U24633 (N_24633,N_24506,N_24512);
xor U24634 (N_24634,N_24530,N_24529);
xnor U24635 (N_24635,N_24478,N_24511);
nand U24636 (N_24636,N_24486,N_24400);
nor U24637 (N_24637,N_24464,N_24401);
or U24638 (N_24638,N_24542,N_24555);
xnor U24639 (N_24639,N_24441,N_24426);
nor U24640 (N_24640,N_24408,N_24437);
or U24641 (N_24641,N_24433,N_24559);
nor U24642 (N_24642,N_24515,N_24448);
and U24643 (N_24643,N_24599,N_24446);
or U24644 (N_24644,N_24421,N_24560);
nor U24645 (N_24645,N_24494,N_24492);
nand U24646 (N_24646,N_24419,N_24549);
nor U24647 (N_24647,N_24589,N_24404);
or U24648 (N_24648,N_24414,N_24450);
nor U24649 (N_24649,N_24422,N_24526);
or U24650 (N_24650,N_24487,N_24459);
nor U24651 (N_24651,N_24502,N_24598);
or U24652 (N_24652,N_24544,N_24420);
or U24653 (N_24653,N_24507,N_24553);
nor U24654 (N_24654,N_24418,N_24568);
nand U24655 (N_24655,N_24552,N_24523);
xnor U24656 (N_24656,N_24583,N_24518);
nand U24657 (N_24657,N_24576,N_24541);
and U24658 (N_24658,N_24509,N_24586);
xnor U24659 (N_24659,N_24538,N_24497);
xnor U24660 (N_24660,N_24533,N_24496);
nand U24661 (N_24661,N_24536,N_24498);
nand U24662 (N_24662,N_24513,N_24431);
nand U24663 (N_24663,N_24524,N_24439);
nand U24664 (N_24664,N_24412,N_24548);
nand U24665 (N_24665,N_24582,N_24442);
or U24666 (N_24666,N_24405,N_24574);
or U24667 (N_24667,N_24491,N_24543);
nand U24668 (N_24668,N_24458,N_24539);
xor U24669 (N_24669,N_24561,N_24460);
xor U24670 (N_24670,N_24504,N_24532);
nor U24671 (N_24671,N_24463,N_24551);
or U24672 (N_24672,N_24519,N_24473);
and U24673 (N_24673,N_24472,N_24476);
nor U24674 (N_24674,N_24567,N_24562);
nor U24675 (N_24675,N_24554,N_24468);
xor U24676 (N_24676,N_24470,N_24547);
or U24677 (N_24677,N_24557,N_24521);
nor U24678 (N_24678,N_24527,N_24410);
nor U24679 (N_24679,N_24474,N_24488);
nor U24680 (N_24680,N_24517,N_24445);
and U24681 (N_24681,N_24495,N_24579);
nor U24682 (N_24682,N_24471,N_24516);
nor U24683 (N_24683,N_24594,N_24413);
xnor U24684 (N_24684,N_24522,N_24429);
nand U24685 (N_24685,N_24595,N_24434);
and U24686 (N_24686,N_24575,N_24570);
nor U24687 (N_24687,N_24503,N_24588);
xnor U24688 (N_24688,N_24449,N_24584);
nor U24689 (N_24689,N_24443,N_24550);
nor U24690 (N_24690,N_24411,N_24571);
or U24691 (N_24691,N_24531,N_24520);
nand U24692 (N_24692,N_24572,N_24564);
xnor U24693 (N_24693,N_24432,N_24597);
or U24694 (N_24694,N_24558,N_24484);
or U24695 (N_24695,N_24430,N_24535);
or U24696 (N_24696,N_24540,N_24510);
nand U24697 (N_24697,N_24528,N_24435);
nand U24698 (N_24698,N_24493,N_24545);
nor U24699 (N_24699,N_24590,N_24454);
nand U24700 (N_24700,N_24424,N_24444);
nor U24701 (N_24701,N_24403,N_24480);
nand U24702 (N_24702,N_24568,N_24456);
and U24703 (N_24703,N_24406,N_24431);
and U24704 (N_24704,N_24454,N_24592);
xnor U24705 (N_24705,N_24410,N_24525);
or U24706 (N_24706,N_24561,N_24568);
and U24707 (N_24707,N_24580,N_24453);
xor U24708 (N_24708,N_24503,N_24526);
or U24709 (N_24709,N_24438,N_24545);
nand U24710 (N_24710,N_24553,N_24401);
nand U24711 (N_24711,N_24437,N_24499);
xnor U24712 (N_24712,N_24493,N_24504);
and U24713 (N_24713,N_24459,N_24492);
xnor U24714 (N_24714,N_24497,N_24569);
nand U24715 (N_24715,N_24575,N_24539);
nand U24716 (N_24716,N_24519,N_24412);
nor U24717 (N_24717,N_24490,N_24594);
nor U24718 (N_24718,N_24562,N_24469);
xor U24719 (N_24719,N_24549,N_24565);
and U24720 (N_24720,N_24439,N_24560);
nand U24721 (N_24721,N_24451,N_24494);
nor U24722 (N_24722,N_24572,N_24550);
nor U24723 (N_24723,N_24526,N_24544);
and U24724 (N_24724,N_24586,N_24416);
and U24725 (N_24725,N_24425,N_24476);
nor U24726 (N_24726,N_24475,N_24495);
or U24727 (N_24727,N_24546,N_24557);
or U24728 (N_24728,N_24510,N_24406);
and U24729 (N_24729,N_24466,N_24485);
nor U24730 (N_24730,N_24438,N_24416);
nor U24731 (N_24731,N_24490,N_24425);
nand U24732 (N_24732,N_24517,N_24473);
nor U24733 (N_24733,N_24511,N_24499);
xnor U24734 (N_24734,N_24590,N_24548);
and U24735 (N_24735,N_24450,N_24516);
nand U24736 (N_24736,N_24417,N_24522);
or U24737 (N_24737,N_24540,N_24439);
or U24738 (N_24738,N_24542,N_24441);
and U24739 (N_24739,N_24564,N_24427);
nor U24740 (N_24740,N_24585,N_24586);
xnor U24741 (N_24741,N_24431,N_24517);
xnor U24742 (N_24742,N_24522,N_24593);
or U24743 (N_24743,N_24488,N_24515);
nand U24744 (N_24744,N_24503,N_24476);
nand U24745 (N_24745,N_24536,N_24575);
or U24746 (N_24746,N_24586,N_24521);
nor U24747 (N_24747,N_24558,N_24402);
or U24748 (N_24748,N_24580,N_24575);
nand U24749 (N_24749,N_24499,N_24578);
and U24750 (N_24750,N_24585,N_24563);
and U24751 (N_24751,N_24594,N_24514);
nor U24752 (N_24752,N_24499,N_24449);
and U24753 (N_24753,N_24569,N_24408);
and U24754 (N_24754,N_24463,N_24424);
nand U24755 (N_24755,N_24552,N_24594);
xor U24756 (N_24756,N_24438,N_24537);
or U24757 (N_24757,N_24508,N_24527);
nand U24758 (N_24758,N_24511,N_24567);
xor U24759 (N_24759,N_24436,N_24431);
nand U24760 (N_24760,N_24436,N_24514);
and U24761 (N_24761,N_24562,N_24479);
and U24762 (N_24762,N_24466,N_24460);
nand U24763 (N_24763,N_24500,N_24527);
xnor U24764 (N_24764,N_24501,N_24517);
xor U24765 (N_24765,N_24532,N_24544);
nor U24766 (N_24766,N_24518,N_24536);
nor U24767 (N_24767,N_24482,N_24437);
nor U24768 (N_24768,N_24505,N_24598);
and U24769 (N_24769,N_24539,N_24442);
xnor U24770 (N_24770,N_24534,N_24543);
or U24771 (N_24771,N_24439,N_24513);
or U24772 (N_24772,N_24539,N_24580);
nand U24773 (N_24773,N_24472,N_24538);
xor U24774 (N_24774,N_24412,N_24460);
nand U24775 (N_24775,N_24564,N_24498);
xnor U24776 (N_24776,N_24466,N_24524);
xor U24777 (N_24777,N_24554,N_24444);
nand U24778 (N_24778,N_24494,N_24413);
nand U24779 (N_24779,N_24460,N_24444);
nor U24780 (N_24780,N_24476,N_24563);
nand U24781 (N_24781,N_24461,N_24450);
nand U24782 (N_24782,N_24510,N_24596);
nand U24783 (N_24783,N_24401,N_24597);
or U24784 (N_24784,N_24533,N_24563);
xor U24785 (N_24785,N_24563,N_24421);
and U24786 (N_24786,N_24501,N_24564);
and U24787 (N_24787,N_24514,N_24405);
nand U24788 (N_24788,N_24525,N_24404);
and U24789 (N_24789,N_24514,N_24535);
nor U24790 (N_24790,N_24548,N_24535);
xnor U24791 (N_24791,N_24482,N_24514);
or U24792 (N_24792,N_24534,N_24595);
nand U24793 (N_24793,N_24411,N_24430);
and U24794 (N_24794,N_24514,N_24537);
nor U24795 (N_24795,N_24566,N_24528);
nand U24796 (N_24796,N_24510,N_24449);
nor U24797 (N_24797,N_24597,N_24531);
xor U24798 (N_24798,N_24452,N_24457);
and U24799 (N_24799,N_24445,N_24496);
nor U24800 (N_24800,N_24624,N_24608);
xor U24801 (N_24801,N_24607,N_24751);
xnor U24802 (N_24802,N_24669,N_24639);
nor U24803 (N_24803,N_24791,N_24655);
or U24804 (N_24804,N_24653,N_24611);
or U24805 (N_24805,N_24780,N_24688);
or U24806 (N_24806,N_24755,N_24619);
and U24807 (N_24807,N_24625,N_24659);
nor U24808 (N_24808,N_24798,N_24760);
and U24809 (N_24809,N_24786,N_24753);
nand U24810 (N_24810,N_24726,N_24649);
nand U24811 (N_24811,N_24642,N_24664);
and U24812 (N_24812,N_24699,N_24735);
or U24813 (N_24813,N_24643,N_24630);
or U24814 (N_24814,N_24762,N_24770);
or U24815 (N_24815,N_24772,N_24779);
and U24816 (N_24816,N_24730,N_24616);
xnor U24817 (N_24817,N_24648,N_24675);
and U24818 (N_24818,N_24636,N_24612);
or U24819 (N_24819,N_24746,N_24765);
nand U24820 (N_24820,N_24787,N_24691);
xnor U24821 (N_24821,N_24628,N_24799);
and U24822 (N_24822,N_24646,N_24759);
or U24823 (N_24823,N_24626,N_24641);
xnor U24824 (N_24824,N_24788,N_24718);
nor U24825 (N_24825,N_24677,N_24623);
nand U24826 (N_24826,N_24614,N_24745);
xnor U24827 (N_24827,N_24738,N_24609);
or U24828 (N_24828,N_24678,N_24661);
and U24829 (N_24829,N_24679,N_24637);
or U24830 (N_24830,N_24701,N_24652);
and U24831 (N_24831,N_24667,N_24671);
nand U24832 (N_24832,N_24681,N_24769);
xnor U24833 (N_24833,N_24632,N_24613);
xor U24834 (N_24834,N_24778,N_24793);
nor U24835 (N_24835,N_24690,N_24721);
nand U24836 (N_24836,N_24668,N_24716);
xor U24837 (N_24837,N_24733,N_24749);
nor U24838 (N_24838,N_24704,N_24672);
and U24839 (N_24839,N_24604,N_24708);
nor U24840 (N_24840,N_24610,N_24727);
and U24841 (N_24841,N_24732,N_24717);
nand U24842 (N_24842,N_24684,N_24794);
nor U24843 (N_24843,N_24693,N_24784);
nor U24844 (N_24844,N_24638,N_24617);
nor U24845 (N_24845,N_24685,N_24777);
nand U24846 (N_24846,N_24647,N_24734);
nand U24847 (N_24847,N_24711,N_24712);
xnor U24848 (N_24848,N_24700,N_24766);
and U24849 (N_24849,N_24694,N_24603);
nor U24850 (N_24850,N_24629,N_24796);
nand U24851 (N_24851,N_24754,N_24742);
nand U24852 (N_24852,N_24650,N_24600);
and U24853 (N_24853,N_24689,N_24767);
nand U24854 (N_24854,N_24605,N_24680);
and U24855 (N_24855,N_24660,N_24670);
xor U24856 (N_24856,N_24776,N_24705);
xnor U24857 (N_24857,N_24601,N_24774);
nand U24858 (N_24858,N_24620,N_24676);
nand U24859 (N_24859,N_24750,N_24710);
nor U24860 (N_24860,N_24768,N_24706);
nand U24861 (N_24861,N_24692,N_24707);
or U24862 (N_24862,N_24702,N_24737);
nor U24863 (N_24863,N_24720,N_24686);
nor U24864 (N_24864,N_24635,N_24622);
and U24865 (N_24865,N_24657,N_24740);
or U24866 (N_24866,N_24665,N_24763);
xor U24867 (N_24867,N_24654,N_24651);
nand U24868 (N_24868,N_24615,N_24773);
or U24869 (N_24869,N_24634,N_24682);
nand U24870 (N_24870,N_24731,N_24656);
and U24871 (N_24871,N_24757,N_24715);
or U24872 (N_24872,N_24709,N_24797);
nand U24873 (N_24873,N_24673,N_24789);
nand U24874 (N_24874,N_24663,N_24747);
nand U24875 (N_24875,N_24739,N_24633);
xnor U24876 (N_24876,N_24743,N_24741);
and U24877 (N_24877,N_24722,N_24645);
nor U24878 (N_24878,N_24736,N_24756);
or U24879 (N_24879,N_24783,N_24781);
or U24880 (N_24880,N_24618,N_24713);
and U24881 (N_24881,N_24698,N_24640);
nand U24882 (N_24882,N_24627,N_24725);
xor U24883 (N_24883,N_24785,N_24795);
nand U24884 (N_24884,N_24696,N_24723);
nand U24885 (N_24885,N_24683,N_24662);
nand U24886 (N_24886,N_24764,N_24790);
nor U24887 (N_24887,N_24687,N_24697);
nor U24888 (N_24888,N_24752,N_24744);
xnor U24889 (N_24889,N_24792,N_24644);
nor U24890 (N_24890,N_24761,N_24729);
xnor U24891 (N_24891,N_24771,N_24606);
nor U24892 (N_24892,N_24703,N_24775);
and U24893 (N_24893,N_24748,N_24758);
and U24894 (N_24894,N_24724,N_24674);
nand U24895 (N_24895,N_24719,N_24621);
or U24896 (N_24896,N_24666,N_24631);
xor U24897 (N_24897,N_24728,N_24695);
nor U24898 (N_24898,N_24602,N_24782);
xnor U24899 (N_24899,N_24714,N_24658);
nor U24900 (N_24900,N_24794,N_24604);
nand U24901 (N_24901,N_24704,N_24713);
nor U24902 (N_24902,N_24749,N_24623);
or U24903 (N_24903,N_24627,N_24799);
xor U24904 (N_24904,N_24727,N_24712);
and U24905 (N_24905,N_24657,N_24669);
nor U24906 (N_24906,N_24754,N_24719);
nand U24907 (N_24907,N_24602,N_24679);
xnor U24908 (N_24908,N_24644,N_24632);
xor U24909 (N_24909,N_24724,N_24766);
or U24910 (N_24910,N_24765,N_24611);
or U24911 (N_24911,N_24699,N_24753);
and U24912 (N_24912,N_24783,N_24717);
and U24913 (N_24913,N_24619,N_24673);
and U24914 (N_24914,N_24649,N_24723);
or U24915 (N_24915,N_24766,N_24628);
nor U24916 (N_24916,N_24724,N_24637);
nor U24917 (N_24917,N_24727,N_24762);
nand U24918 (N_24918,N_24685,N_24654);
nor U24919 (N_24919,N_24666,N_24672);
nand U24920 (N_24920,N_24610,N_24620);
nand U24921 (N_24921,N_24685,N_24687);
nor U24922 (N_24922,N_24633,N_24682);
xor U24923 (N_24923,N_24696,N_24727);
nand U24924 (N_24924,N_24759,N_24772);
xnor U24925 (N_24925,N_24627,N_24695);
and U24926 (N_24926,N_24631,N_24743);
and U24927 (N_24927,N_24731,N_24715);
xor U24928 (N_24928,N_24761,N_24604);
nand U24929 (N_24929,N_24675,N_24758);
or U24930 (N_24930,N_24706,N_24763);
and U24931 (N_24931,N_24720,N_24705);
nand U24932 (N_24932,N_24684,N_24640);
nor U24933 (N_24933,N_24747,N_24692);
and U24934 (N_24934,N_24670,N_24721);
or U24935 (N_24935,N_24782,N_24661);
xor U24936 (N_24936,N_24622,N_24762);
nor U24937 (N_24937,N_24770,N_24735);
xor U24938 (N_24938,N_24719,N_24783);
nor U24939 (N_24939,N_24776,N_24739);
xor U24940 (N_24940,N_24743,N_24687);
xor U24941 (N_24941,N_24636,N_24675);
nor U24942 (N_24942,N_24655,N_24755);
or U24943 (N_24943,N_24600,N_24652);
nor U24944 (N_24944,N_24625,N_24751);
xnor U24945 (N_24945,N_24622,N_24753);
nand U24946 (N_24946,N_24750,N_24727);
xor U24947 (N_24947,N_24720,N_24655);
and U24948 (N_24948,N_24776,N_24687);
and U24949 (N_24949,N_24622,N_24798);
xnor U24950 (N_24950,N_24776,N_24646);
or U24951 (N_24951,N_24604,N_24759);
nand U24952 (N_24952,N_24615,N_24727);
or U24953 (N_24953,N_24643,N_24786);
and U24954 (N_24954,N_24797,N_24621);
or U24955 (N_24955,N_24703,N_24630);
or U24956 (N_24956,N_24768,N_24751);
and U24957 (N_24957,N_24685,N_24610);
xnor U24958 (N_24958,N_24640,N_24602);
xnor U24959 (N_24959,N_24706,N_24699);
or U24960 (N_24960,N_24729,N_24713);
and U24961 (N_24961,N_24698,N_24659);
or U24962 (N_24962,N_24607,N_24773);
nand U24963 (N_24963,N_24717,N_24761);
nor U24964 (N_24964,N_24720,N_24687);
nor U24965 (N_24965,N_24604,N_24744);
and U24966 (N_24966,N_24717,N_24706);
nand U24967 (N_24967,N_24788,N_24725);
or U24968 (N_24968,N_24794,N_24791);
and U24969 (N_24969,N_24706,N_24761);
nand U24970 (N_24970,N_24766,N_24679);
nor U24971 (N_24971,N_24722,N_24743);
xnor U24972 (N_24972,N_24685,N_24639);
nand U24973 (N_24973,N_24728,N_24727);
nand U24974 (N_24974,N_24784,N_24741);
or U24975 (N_24975,N_24683,N_24688);
xor U24976 (N_24976,N_24688,N_24790);
and U24977 (N_24977,N_24650,N_24667);
nor U24978 (N_24978,N_24718,N_24797);
nor U24979 (N_24979,N_24610,N_24779);
and U24980 (N_24980,N_24650,N_24774);
xor U24981 (N_24981,N_24746,N_24650);
or U24982 (N_24982,N_24747,N_24662);
xor U24983 (N_24983,N_24750,N_24611);
nor U24984 (N_24984,N_24684,N_24685);
and U24985 (N_24985,N_24730,N_24690);
or U24986 (N_24986,N_24776,N_24666);
xor U24987 (N_24987,N_24734,N_24664);
and U24988 (N_24988,N_24750,N_24612);
xor U24989 (N_24989,N_24619,N_24603);
nand U24990 (N_24990,N_24611,N_24675);
nor U24991 (N_24991,N_24700,N_24686);
nand U24992 (N_24992,N_24735,N_24642);
xnor U24993 (N_24993,N_24678,N_24658);
nor U24994 (N_24994,N_24645,N_24684);
or U24995 (N_24995,N_24789,N_24639);
or U24996 (N_24996,N_24797,N_24755);
nor U24997 (N_24997,N_24793,N_24685);
nand U24998 (N_24998,N_24699,N_24778);
and U24999 (N_24999,N_24626,N_24757);
and UO_0 (O_0,N_24880,N_24991);
nand UO_1 (O_1,N_24885,N_24959);
nor UO_2 (O_2,N_24839,N_24812);
or UO_3 (O_3,N_24803,N_24939);
nor UO_4 (O_4,N_24845,N_24809);
nand UO_5 (O_5,N_24883,N_24882);
or UO_6 (O_6,N_24844,N_24889);
and UO_7 (O_7,N_24817,N_24971);
nor UO_8 (O_8,N_24895,N_24919);
xor UO_9 (O_9,N_24977,N_24943);
xor UO_10 (O_10,N_24905,N_24923);
or UO_11 (O_11,N_24800,N_24940);
xor UO_12 (O_12,N_24976,N_24820);
or UO_13 (O_13,N_24806,N_24855);
or UO_14 (O_14,N_24887,N_24928);
nand UO_15 (O_15,N_24890,N_24848);
nand UO_16 (O_16,N_24850,N_24818);
and UO_17 (O_17,N_24900,N_24915);
and UO_18 (O_18,N_24810,N_24918);
and UO_19 (O_19,N_24869,N_24938);
xnor UO_20 (O_20,N_24945,N_24909);
or UO_21 (O_21,N_24995,N_24870);
or UO_22 (O_22,N_24875,N_24825);
and UO_23 (O_23,N_24993,N_24886);
nor UO_24 (O_24,N_24912,N_24866);
or UO_25 (O_25,N_24947,N_24951);
and UO_26 (O_26,N_24807,N_24841);
and UO_27 (O_27,N_24907,N_24861);
nand UO_28 (O_28,N_24873,N_24950);
nand UO_29 (O_29,N_24904,N_24893);
xnor UO_30 (O_30,N_24932,N_24933);
nor UO_31 (O_31,N_24980,N_24990);
and UO_32 (O_32,N_24847,N_24836);
nand UO_33 (O_33,N_24966,N_24981);
xnor UO_34 (O_34,N_24901,N_24874);
or UO_35 (O_35,N_24878,N_24862);
nand UO_36 (O_36,N_24996,N_24823);
xnor UO_37 (O_37,N_24804,N_24908);
nor UO_38 (O_38,N_24877,N_24999);
or UO_39 (O_39,N_24979,N_24962);
xor UO_40 (O_40,N_24902,N_24924);
and UO_41 (O_41,N_24840,N_24960);
xnor UO_42 (O_42,N_24838,N_24937);
or UO_43 (O_43,N_24968,N_24984);
nor UO_44 (O_44,N_24987,N_24865);
xnor UO_45 (O_45,N_24973,N_24801);
or UO_46 (O_46,N_24994,N_24916);
or UO_47 (O_47,N_24842,N_24992);
and UO_48 (O_48,N_24811,N_24964);
and UO_49 (O_49,N_24985,N_24974);
or UO_50 (O_50,N_24911,N_24876);
nand UO_51 (O_51,N_24936,N_24802);
or UO_52 (O_52,N_24813,N_24986);
nand UO_53 (O_53,N_24832,N_24961);
and UO_54 (O_54,N_24989,N_24958);
xor UO_55 (O_55,N_24983,N_24891);
or UO_56 (O_56,N_24853,N_24969);
or UO_57 (O_57,N_24881,N_24897);
nand UO_58 (O_58,N_24896,N_24920);
nand UO_59 (O_59,N_24884,N_24982);
xnor UO_60 (O_60,N_24888,N_24944);
or UO_61 (O_61,N_24846,N_24868);
and UO_62 (O_62,N_24879,N_24914);
xnor UO_63 (O_63,N_24814,N_24808);
or UO_64 (O_64,N_24929,N_24835);
xnor UO_65 (O_65,N_24949,N_24921);
nor UO_66 (O_66,N_24826,N_24860);
and UO_67 (O_67,N_24954,N_24952);
xnor UO_68 (O_68,N_24967,N_24833);
nor UO_69 (O_69,N_24871,N_24837);
or UO_70 (O_70,N_24858,N_24828);
nor UO_71 (O_71,N_24824,N_24854);
nand UO_72 (O_72,N_24906,N_24864);
and UO_73 (O_73,N_24934,N_24815);
nor UO_74 (O_74,N_24913,N_24957);
nand UO_75 (O_75,N_24867,N_24998);
nand UO_76 (O_76,N_24852,N_24925);
nor UO_77 (O_77,N_24851,N_24863);
xor UO_78 (O_78,N_24948,N_24859);
xor UO_79 (O_79,N_24946,N_24819);
nor UO_80 (O_80,N_24975,N_24805);
xor UO_81 (O_81,N_24816,N_24917);
xor UO_82 (O_82,N_24972,N_24857);
nor UO_83 (O_83,N_24827,N_24997);
or UO_84 (O_84,N_24953,N_24942);
or UO_85 (O_85,N_24903,N_24963);
and UO_86 (O_86,N_24831,N_24821);
nor UO_87 (O_87,N_24894,N_24956);
or UO_88 (O_88,N_24970,N_24898);
xnor UO_89 (O_89,N_24829,N_24892);
xnor UO_90 (O_90,N_24856,N_24988);
xor UO_91 (O_91,N_24822,N_24926);
nand UO_92 (O_92,N_24830,N_24955);
xnor UO_93 (O_93,N_24922,N_24930);
and UO_94 (O_94,N_24843,N_24899);
nand UO_95 (O_95,N_24931,N_24834);
nor UO_96 (O_96,N_24872,N_24965);
xnor UO_97 (O_97,N_24910,N_24978);
or UO_98 (O_98,N_24935,N_24941);
or UO_99 (O_99,N_24849,N_24927);
nand UO_100 (O_100,N_24992,N_24987);
nand UO_101 (O_101,N_24838,N_24855);
nand UO_102 (O_102,N_24873,N_24846);
nor UO_103 (O_103,N_24878,N_24952);
nand UO_104 (O_104,N_24823,N_24817);
or UO_105 (O_105,N_24907,N_24960);
and UO_106 (O_106,N_24929,N_24902);
and UO_107 (O_107,N_24901,N_24957);
xnor UO_108 (O_108,N_24834,N_24844);
xnor UO_109 (O_109,N_24956,N_24878);
nand UO_110 (O_110,N_24811,N_24876);
or UO_111 (O_111,N_24829,N_24996);
or UO_112 (O_112,N_24863,N_24936);
xor UO_113 (O_113,N_24838,N_24887);
nand UO_114 (O_114,N_24823,N_24818);
and UO_115 (O_115,N_24895,N_24954);
and UO_116 (O_116,N_24983,N_24966);
and UO_117 (O_117,N_24906,N_24820);
nor UO_118 (O_118,N_24947,N_24907);
nor UO_119 (O_119,N_24836,N_24824);
nand UO_120 (O_120,N_24928,N_24884);
xnor UO_121 (O_121,N_24966,N_24852);
xnor UO_122 (O_122,N_24928,N_24925);
xnor UO_123 (O_123,N_24975,N_24991);
nor UO_124 (O_124,N_24996,N_24983);
nor UO_125 (O_125,N_24814,N_24895);
or UO_126 (O_126,N_24842,N_24994);
nor UO_127 (O_127,N_24878,N_24868);
nor UO_128 (O_128,N_24951,N_24888);
nor UO_129 (O_129,N_24915,N_24869);
or UO_130 (O_130,N_24901,N_24895);
nand UO_131 (O_131,N_24977,N_24805);
and UO_132 (O_132,N_24960,N_24978);
nor UO_133 (O_133,N_24974,N_24800);
and UO_134 (O_134,N_24931,N_24826);
and UO_135 (O_135,N_24840,N_24906);
or UO_136 (O_136,N_24976,N_24923);
nor UO_137 (O_137,N_24903,N_24814);
nor UO_138 (O_138,N_24982,N_24973);
xnor UO_139 (O_139,N_24932,N_24992);
xnor UO_140 (O_140,N_24879,N_24897);
or UO_141 (O_141,N_24897,N_24847);
and UO_142 (O_142,N_24940,N_24875);
xnor UO_143 (O_143,N_24840,N_24907);
nor UO_144 (O_144,N_24859,N_24858);
and UO_145 (O_145,N_24813,N_24809);
nor UO_146 (O_146,N_24900,N_24893);
xnor UO_147 (O_147,N_24884,N_24826);
xor UO_148 (O_148,N_24998,N_24950);
nand UO_149 (O_149,N_24847,N_24967);
nor UO_150 (O_150,N_24955,N_24998);
xor UO_151 (O_151,N_24800,N_24997);
and UO_152 (O_152,N_24955,N_24922);
xnor UO_153 (O_153,N_24823,N_24900);
xnor UO_154 (O_154,N_24812,N_24849);
and UO_155 (O_155,N_24962,N_24949);
and UO_156 (O_156,N_24807,N_24991);
or UO_157 (O_157,N_24969,N_24939);
nand UO_158 (O_158,N_24850,N_24943);
nor UO_159 (O_159,N_24944,N_24880);
nor UO_160 (O_160,N_24880,N_24817);
nand UO_161 (O_161,N_24843,N_24983);
and UO_162 (O_162,N_24989,N_24875);
and UO_163 (O_163,N_24910,N_24838);
nor UO_164 (O_164,N_24849,N_24874);
nand UO_165 (O_165,N_24947,N_24835);
nor UO_166 (O_166,N_24980,N_24972);
nor UO_167 (O_167,N_24886,N_24974);
xnor UO_168 (O_168,N_24822,N_24897);
nor UO_169 (O_169,N_24842,N_24857);
and UO_170 (O_170,N_24974,N_24954);
or UO_171 (O_171,N_24857,N_24880);
nor UO_172 (O_172,N_24945,N_24828);
nand UO_173 (O_173,N_24983,N_24872);
xnor UO_174 (O_174,N_24816,N_24885);
xnor UO_175 (O_175,N_24854,N_24934);
xor UO_176 (O_176,N_24865,N_24928);
nand UO_177 (O_177,N_24987,N_24874);
nor UO_178 (O_178,N_24816,N_24967);
or UO_179 (O_179,N_24938,N_24975);
xor UO_180 (O_180,N_24900,N_24952);
xnor UO_181 (O_181,N_24869,N_24855);
xor UO_182 (O_182,N_24936,N_24847);
and UO_183 (O_183,N_24976,N_24882);
xnor UO_184 (O_184,N_24822,N_24827);
or UO_185 (O_185,N_24942,N_24954);
nand UO_186 (O_186,N_24964,N_24842);
or UO_187 (O_187,N_24891,N_24837);
xnor UO_188 (O_188,N_24960,N_24814);
nand UO_189 (O_189,N_24810,N_24817);
nor UO_190 (O_190,N_24967,N_24943);
nor UO_191 (O_191,N_24968,N_24832);
and UO_192 (O_192,N_24801,N_24943);
nand UO_193 (O_193,N_24931,N_24913);
xor UO_194 (O_194,N_24887,N_24810);
nand UO_195 (O_195,N_24867,N_24827);
or UO_196 (O_196,N_24934,N_24851);
or UO_197 (O_197,N_24928,N_24912);
or UO_198 (O_198,N_24907,N_24961);
nand UO_199 (O_199,N_24838,N_24899);
and UO_200 (O_200,N_24818,N_24971);
nor UO_201 (O_201,N_24880,N_24810);
and UO_202 (O_202,N_24918,N_24875);
xnor UO_203 (O_203,N_24936,N_24927);
and UO_204 (O_204,N_24996,N_24843);
nand UO_205 (O_205,N_24939,N_24833);
nor UO_206 (O_206,N_24813,N_24915);
and UO_207 (O_207,N_24923,N_24865);
nand UO_208 (O_208,N_24829,N_24958);
or UO_209 (O_209,N_24837,N_24995);
and UO_210 (O_210,N_24999,N_24906);
nor UO_211 (O_211,N_24818,N_24871);
nor UO_212 (O_212,N_24913,N_24919);
and UO_213 (O_213,N_24919,N_24838);
and UO_214 (O_214,N_24875,N_24976);
or UO_215 (O_215,N_24965,N_24957);
or UO_216 (O_216,N_24821,N_24935);
nand UO_217 (O_217,N_24850,N_24876);
nor UO_218 (O_218,N_24989,N_24998);
xnor UO_219 (O_219,N_24830,N_24963);
and UO_220 (O_220,N_24939,N_24827);
or UO_221 (O_221,N_24990,N_24828);
nor UO_222 (O_222,N_24957,N_24919);
nand UO_223 (O_223,N_24846,N_24943);
and UO_224 (O_224,N_24812,N_24990);
nor UO_225 (O_225,N_24878,N_24924);
xor UO_226 (O_226,N_24850,N_24832);
nand UO_227 (O_227,N_24997,N_24948);
and UO_228 (O_228,N_24951,N_24979);
or UO_229 (O_229,N_24822,N_24983);
or UO_230 (O_230,N_24912,N_24872);
xor UO_231 (O_231,N_24816,N_24978);
and UO_232 (O_232,N_24996,N_24968);
xor UO_233 (O_233,N_24948,N_24923);
xnor UO_234 (O_234,N_24924,N_24850);
xor UO_235 (O_235,N_24960,N_24837);
and UO_236 (O_236,N_24826,N_24952);
nand UO_237 (O_237,N_24875,N_24953);
nor UO_238 (O_238,N_24841,N_24975);
or UO_239 (O_239,N_24975,N_24829);
nor UO_240 (O_240,N_24814,N_24874);
xor UO_241 (O_241,N_24881,N_24808);
nor UO_242 (O_242,N_24974,N_24836);
nand UO_243 (O_243,N_24973,N_24953);
nand UO_244 (O_244,N_24800,N_24893);
nand UO_245 (O_245,N_24929,N_24873);
and UO_246 (O_246,N_24847,N_24803);
and UO_247 (O_247,N_24913,N_24823);
or UO_248 (O_248,N_24865,N_24910);
xnor UO_249 (O_249,N_24887,N_24964);
and UO_250 (O_250,N_24979,N_24845);
nand UO_251 (O_251,N_24990,N_24891);
nor UO_252 (O_252,N_24884,N_24802);
or UO_253 (O_253,N_24946,N_24980);
nor UO_254 (O_254,N_24827,N_24976);
or UO_255 (O_255,N_24990,N_24813);
xnor UO_256 (O_256,N_24819,N_24950);
and UO_257 (O_257,N_24929,N_24928);
nor UO_258 (O_258,N_24892,N_24980);
nand UO_259 (O_259,N_24947,N_24870);
nor UO_260 (O_260,N_24999,N_24886);
or UO_261 (O_261,N_24954,N_24873);
and UO_262 (O_262,N_24841,N_24853);
or UO_263 (O_263,N_24904,N_24933);
xnor UO_264 (O_264,N_24867,N_24877);
nand UO_265 (O_265,N_24987,N_24920);
nand UO_266 (O_266,N_24887,N_24933);
nor UO_267 (O_267,N_24881,N_24907);
or UO_268 (O_268,N_24994,N_24878);
xor UO_269 (O_269,N_24928,N_24829);
and UO_270 (O_270,N_24975,N_24814);
nand UO_271 (O_271,N_24911,N_24906);
and UO_272 (O_272,N_24952,N_24869);
xnor UO_273 (O_273,N_24901,N_24897);
or UO_274 (O_274,N_24835,N_24811);
and UO_275 (O_275,N_24983,N_24809);
nor UO_276 (O_276,N_24898,N_24902);
nor UO_277 (O_277,N_24810,N_24809);
nor UO_278 (O_278,N_24920,N_24820);
nand UO_279 (O_279,N_24929,N_24991);
nand UO_280 (O_280,N_24869,N_24997);
nor UO_281 (O_281,N_24975,N_24863);
or UO_282 (O_282,N_24912,N_24999);
and UO_283 (O_283,N_24995,N_24953);
nand UO_284 (O_284,N_24843,N_24981);
nand UO_285 (O_285,N_24965,N_24930);
or UO_286 (O_286,N_24980,N_24904);
and UO_287 (O_287,N_24827,N_24832);
and UO_288 (O_288,N_24938,N_24968);
xor UO_289 (O_289,N_24839,N_24831);
nand UO_290 (O_290,N_24819,N_24832);
nor UO_291 (O_291,N_24860,N_24844);
nand UO_292 (O_292,N_24868,N_24872);
and UO_293 (O_293,N_24922,N_24986);
nand UO_294 (O_294,N_24842,N_24934);
and UO_295 (O_295,N_24931,N_24857);
nand UO_296 (O_296,N_24907,N_24973);
nand UO_297 (O_297,N_24939,N_24886);
nor UO_298 (O_298,N_24916,N_24975);
and UO_299 (O_299,N_24879,N_24996);
and UO_300 (O_300,N_24999,N_24816);
and UO_301 (O_301,N_24948,N_24973);
or UO_302 (O_302,N_24971,N_24838);
nand UO_303 (O_303,N_24823,N_24989);
or UO_304 (O_304,N_24925,N_24980);
or UO_305 (O_305,N_24931,N_24997);
xnor UO_306 (O_306,N_24835,N_24983);
or UO_307 (O_307,N_24915,N_24986);
nor UO_308 (O_308,N_24927,N_24939);
nor UO_309 (O_309,N_24880,N_24958);
or UO_310 (O_310,N_24845,N_24898);
and UO_311 (O_311,N_24901,N_24835);
nand UO_312 (O_312,N_24957,N_24855);
xnor UO_313 (O_313,N_24865,N_24897);
or UO_314 (O_314,N_24910,N_24862);
or UO_315 (O_315,N_24822,N_24844);
and UO_316 (O_316,N_24973,N_24853);
xor UO_317 (O_317,N_24843,N_24824);
or UO_318 (O_318,N_24870,N_24860);
and UO_319 (O_319,N_24862,N_24877);
and UO_320 (O_320,N_24801,N_24870);
or UO_321 (O_321,N_24889,N_24894);
nor UO_322 (O_322,N_24936,N_24875);
or UO_323 (O_323,N_24979,N_24887);
or UO_324 (O_324,N_24983,N_24933);
nand UO_325 (O_325,N_24854,N_24828);
or UO_326 (O_326,N_24959,N_24892);
nand UO_327 (O_327,N_24834,N_24847);
nand UO_328 (O_328,N_24909,N_24881);
or UO_329 (O_329,N_24916,N_24855);
nor UO_330 (O_330,N_24875,N_24926);
or UO_331 (O_331,N_24900,N_24842);
or UO_332 (O_332,N_24809,N_24818);
nor UO_333 (O_333,N_24931,N_24838);
nand UO_334 (O_334,N_24911,N_24830);
nand UO_335 (O_335,N_24872,N_24902);
nand UO_336 (O_336,N_24925,N_24931);
xor UO_337 (O_337,N_24905,N_24888);
nand UO_338 (O_338,N_24839,N_24832);
xor UO_339 (O_339,N_24922,N_24873);
nor UO_340 (O_340,N_24881,N_24883);
xor UO_341 (O_341,N_24883,N_24886);
xor UO_342 (O_342,N_24967,N_24960);
and UO_343 (O_343,N_24927,N_24989);
and UO_344 (O_344,N_24804,N_24948);
or UO_345 (O_345,N_24939,N_24959);
and UO_346 (O_346,N_24940,N_24976);
nand UO_347 (O_347,N_24910,N_24960);
or UO_348 (O_348,N_24828,N_24846);
nor UO_349 (O_349,N_24817,N_24820);
nor UO_350 (O_350,N_24995,N_24819);
nor UO_351 (O_351,N_24854,N_24865);
nor UO_352 (O_352,N_24937,N_24946);
nor UO_353 (O_353,N_24815,N_24807);
or UO_354 (O_354,N_24918,N_24899);
and UO_355 (O_355,N_24919,N_24971);
xor UO_356 (O_356,N_24967,N_24875);
xnor UO_357 (O_357,N_24994,N_24928);
nor UO_358 (O_358,N_24839,N_24905);
nor UO_359 (O_359,N_24803,N_24890);
nand UO_360 (O_360,N_24915,N_24837);
nand UO_361 (O_361,N_24895,N_24990);
xnor UO_362 (O_362,N_24994,N_24965);
and UO_363 (O_363,N_24877,N_24901);
or UO_364 (O_364,N_24829,N_24801);
nor UO_365 (O_365,N_24849,N_24867);
xor UO_366 (O_366,N_24895,N_24932);
and UO_367 (O_367,N_24957,N_24999);
xnor UO_368 (O_368,N_24995,N_24851);
nor UO_369 (O_369,N_24809,N_24859);
or UO_370 (O_370,N_24915,N_24974);
nor UO_371 (O_371,N_24954,N_24883);
nand UO_372 (O_372,N_24802,N_24870);
nand UO_373 (O_373,N_24918,N_24905);
and UO_374 (O_374,N_24890,N_24877);
xor UO_375 (O_375,N_24862,N_24900);
or UO_376 (O_376,N_24985,N_24881);
nand UO_377 (O_377,N_24892,N_24824);
nand UO_378 (O_378,N_24847,N_24926);
or UO_379 (O_379,N_24860,N_24857);
xnor UO_380 (O_380,N_24828,N_24804);
nor UO_381 (O_381,N_24905,N_24893);
nand UO_382 (O_382,N_24929,N_24838);
and UO_383 (O_383,N_24891,N_24995);
nor UO_384 (O_384,N_24947,N_24812);
nor UO_385 (O_385,N_24824,N_24967);
and UO_386 (O_386,N_24991,N_24936);
nor UO_387 (O_387,N_24928,N_24845);
nor UO_388 (O_388,N_24985,N_24957);
and UO_389 (O_389,N_24819,N_24862);
xor UO_390 (O_390,N_24978,N_24863);
and UO_391 (O_391,N_24827,N_24803);
nand UO_392 (O_392,N_24995,N_24918);
nand UO_393 (O_393,N_24937,N_24909);
and UO_394 (O_394,N_24972,N_24998);
nand UO_395 (O_395,N_24806,N_24931);
or UO_396 (O_396,N_24807,N_24858);
nand UO_397 (O_397,N_24868,N_24860);
or UO_398 (O_398,N_24945,N_24931);
or UO_399 (O_399,N_24953,N_24989);
and UO_400 (O_400,N_24939,N_24838);
xnor UO_401 (O_401,N_24917,N_24886);
nand UO_402 (O_402,N_24894,N_24908);
nand UO_403 (O_403,N_24800,N_24889);
nor UO_404 (O_404,N_24898,N_24999);
or UO_405 (O_405,N_24829,N_24808);
nor UO_406 (O_406,N_24816,N_24813);
nand UO_407 (O_407,N_24914,N_24858);
and UO_408 (O_408,N_24885,N_24838);
xor UO_409 (O_409,N_24942,N_24897);
xor UO_410 (O_410,N_24875,N_24947);
and UO_411 (O_411,N_24919,N_24891);
nand UO_412 (O_412,N_24985,N_24813);
nand UO_413 (O_413,N_24994,N_24849);
nor UO_414 (O_414,N_24854,N_24841);
or UO_415 (O_415,N_24927,N_24825);
or UO_416 (O_416,N_24985,N_24899);
nor UO_417 (O_417,N_24961,N_24941);
xor UO_418 (O_418,N_24815,N_24827);
or UO_419 (O_419,N_24887,N_24823);
or UO_420 (O_420,N_24851,N_24994);
or UO_421 (O_421,N_24899,N_24860);
nor UO_422 (O_422,N_24851,N_24881);
xor UO_423 (O_423,N_24813,N_24856);
or UO_424 (O_424,N_24862,N_24857);
nor UO_425 (O_425,N_24821,N_24825);
nand UO_426 (O_426,N_24813,N_24935);
nand UO_427 (O_427,N_24910,N_24980);
nand UO_428 (O_428,N_24901,N_24984);
nand UO_429 (O_429,N_24951,N_24904);
or UO_430 (O_430,N_24810,N_24884);
nor UO_431 (O_431,N_24959,N_24854);
nor UO_432 (O_432,N_24899,N_24947);
or UO_433 (O_433,N_24881,N_24846);
xor UO_434 (O_434,N_24878,N_24998);
nand UO_435 (O_435,N_24983,N_24838);
xor UO_436 (O_436,N_24888,N_24986);
xnor UO_437 (O_437,N_24880,N_24979);
xor UO_438 (O_438,N_24807,N_24961);
and UO_439 (O_439,N_24918,N_24843);
and UO_440 (O_440,N_24817,N_24938);
and UO_441 (O_441,N_24955,N_24963);
nand UO_442 (O_442,N_24904,N_24828);
or UO_443 (O_443,N_24905,N_24951);
nor UO_444 (O_444,N_24819,N_24912);
xnor UO_445 (O_445,N_24847,N_24877);
nand UO_446 (O_446,N_24866,N_24993);
nand UO_447 (O_447,N_24885,N_24992);
xor UO_448 (O_448,N_24836,N_24912);
nor UO_449 (O_449,N_24982,N_24873);
and UO_450 (O_450,N_24962,N_24871);
xor UO_451 (O_451,N_24992,N_24814);
xnor UO_452 (O_452,N_24808,N_24873);
and UO_453 (O_453,N_24867,N_24930);
and UO_454 (O_454,N_24891,N_24849);
xor UO_455 (O_455,N_24845,N_24983);
or UO_456 (O_456,N_24968,N_24925);
and UO_457 (O_457,N_24815,N_24906);
or UO_458 (O_458,N_24871,N_24945);
nor UO_459 (O_459,N_24989,N_24821);
and UO_460 (O_460,N_24969,N_24958);
nand UO_461 (O_461,N_24860,N_24956);
xor UO_462 (O_462,N_24812,N_24857);
nor UO_463 (O_463,N_24954,N_24898);
nand UO_464 (O_464,N_24825,N_24935);
nor UO_465 (O_465,N_24909,N_24875);
nor UO_466 (O_466,N_24870,N_24997);
or UO_467 (O_467,N_24821,N_24910);
nor UO_468 (O_468,N_24906,N_24932);
xor UO_469 (O_469,N_24919,N_24871);
and UO_470 (O_470,N_24897,N_24925);
xnor UO_471 (O_471,N_24877,N_24955);
or UO_472 (O_472,N_24848,N_24820);
or UO_473 (O_473,N_24909,N_24916);
and UO_474 (O_474,N_24908,N_24821);
xor UO_475 (O_475,N_24823,N_24915);
or UO_476 (O_476,N_24977,N_24958);
xnor UO_477 (O_477,N_24819,N_24969);
xor UO_478 (O_478,N_24899,N_24988);
nor UO_479 (O_479,N_24845,N_24812);
nor UO_480 (O_480,N_24904,N_24936);
or UO_481 (O_481,N_24891,N_24965);
xor UO_482 (O_482,N_24976,N_24819);
nor UO_483 (O_483,N_24975,N_24803);
and UO_484 (O_484,N_24932,N_24824);
or UO_485 (O_485,N_24819,N_24846);
nand UO_486 (O_486,N_24944,N_24997);
nor UO_487 (O_487,N_24910,N_24849);
and UO_488 (O_488,N_24928,N_24957);
and UO_489 (O_489,N_24911,N_24800);
xor UO_490 (O_490,N_24859,N_24926);
or UO_491 (O_491,N_24818,N_24825);
and UO_492 (O_492,N_24920,N_24870);
or UO_493 (O_493,N_24917,N_24929);
nor UO_494 (O_494,N_24897,N_24983);
xor UO_495 (O_495,N_24949,N_24849);
nor UO_496 (O_496,N_24896,N_24900);
nor UO_497 (O_497,N_24997,N_24805);
or UO_498 (O_498,N_24905,N_24907);
or UO_499 (O_499,N_24834,N_24816);
or UO_500 (O_500,N_24966,N_24946);
or UO_501 (O_501,N_24838,N_24818);
nor UO_502 (O_502,N_24990,N_24938);
nand UO_503 (O_503,N_24878,N_24818);
and UO_504 (O_504,N_24891,N_24915);
or UO_505 (O_505,N_24973,N_24869);
nand UO_506 (O_506,N_24868,N_24812);
and UO_507 (O_507,N_24872,N_24808);
nor UO_508 (O_508,N_24837,N_24838);
nand UO_509 (O_509,N_24967,N_24901);
nor UO_510 (O_510,N_24914,N_24809);
nor UO_511 (O_511,N_24999,N_24803);
xor UO_512 (O_512,N_24908,N_24850);
and UO_513 (O_513,N_24920,N_24850);
nor UO_514 (O_514,N_24823,N_24907);
and UO_515 (O_515,N_24927,N_24839);
and UO_516 (O_516,N_24803,N_24962);
and UO_517 (O_517,N_24946,N_24958);
xnor UO_518 (O_518,N_24961,N_24800);
nor UO_519 (O_519,N_24834,N_24924);
and UO_520 (O_520,N_24968,N_24992);
nand UO_521 (O_521,N_24888,N_24893);
and UO_522 (O_522,N_24873,N_24877);
nand UO_523 (O_523,N_24819,N_24884);
nand UO_524 (O_524,N_24821,N_24920);
and UO_525 (O_525,N_24837,N_24944);
and UO_526 (O_526,N_24958,N_24988);
or UO_527 (O_527,N_24884,N_24927);
nand UO_528 (O_528,N_24820,N_24936);
or UO_529 (O_529,N_24947,N_24849);
and UO_530 (O_530,N_24959,N_24860);
or UO_531 (O_531,N_24859,N_24818);
xnor UO_532 (O_532,N_24888,N_24920);
nand UO_533 (O_533,N_24995,N_24854);
or UO_534 (O_534,N_24806,N_24803);
nand UO_535 (O_535,N_24903,N_24862);
xnor UO_536 (O_536,N_24903,N_24857);
or UO_537 (O_537,N_24873,N_24899);
or UO_538 (O_538,N_24948,N_24881);
or UO_539 (O_539,N_24832,N_24835);
or UO_540 (O_540,N_24841,N_24806);
nand UO_541 (O_541,N_24904,N_24907);
nand UO_542 (O_542,N_24988,N_24866);
or UO_543 (O_543,N_24827,N_24919);
and UO_544 (O_544,N_24845,N_24982);
xor UO_545 (O_545,N_24869,N_24947);
xnor UO_546 (O_546,N_24926,N_24918);
nor UO_547 (O_547,N_24863,N_24841);
xnor UO_548 (O_548,N_24953,N_24865);
and UO_549 (O_549,N_24831,N_24893);
xor UO_550 (O_550,N_24975,N_24895);
xnor UO_551 (O_551,N_24983,N_24940);
nor UO_552 (O_552,N_24989,N_24962);
nor UO_553 (O_553,N_24983,N_24952);
or UO_554 (O_554,N_24909,N_24927);
xnor UO_555 (O_555,N_24802,N_24874);
and UO_556 (O_556,N_24931,N_24978);
and UO_557 (O_557,N_24832,N_24946);
or UO_558 (O_558,N_24843,N_24833);
nor UO_559 (O_559,N_24990,N_24998);
nand UO_560 (O_560,N_24987,N_24952);
or UO_561 (O_561,N_24882,N_24867);
xnor UO_562 (O_562,N_24953,N_24906);
xor UO_563 (O_563,N_24960,N_24980);
xnor UO_564 (O_564,N_24960,N_24892);
xnor UO_565 (O_565,N_24840,N_24841);
and UO_566 (O_566,N_24841,N_24870);
xor UO_567 (O_567,N_24875,N_24978);
nor UO_568 (O_568,N_24811,N_24993);
nand UO_569 (O_569,N_24981,N_24900);
xor UO_570 (O_570,N_24870,N_24982);
nand UO_571 (O_571,N_24897,N_24990);
nor UO_572 (O_572,N_24934,N_24942);
or UO_573 (O_573,N_24900,N_24944);
or UO_574 (O_574,N_24885,N_24911);
xnor UO_575 (O_575,N_24889,N_24964);
and UO_576 (O_576,N_24806,N_24914);
or UO_577 (O_577,N_24887,N_24914);
xor UO_578 (O_578,N_24839,N_24968);
nand UO_579 (O_579,N_24831,N_24817);
and UO_580 (O_580,N_24886,N_24833);
nor UO_581 (O_581,N_24966,N_24936);
and UO_582 (O_582,N_24945,N_24917);
or UO_583 (O_583,N_24889,N_24852);
and UO_584 (O_584,N_24941,N_24904);
or UO_585 (O_585,N_24932,N_24936);
nor UO_586 (O_586,N_24926,N_24922);
nand UO_587 (O_587,N_24946,N_24853);
nor UO_588 (O_588,N_24955,N_24986);
nand UO_589 (O_589,N_24985,N_24930);
nor UO_590 (O_590,N_24855,N_24930);
and UO_591 (O_591,N_24989,N_24889);
or UO_592 (O_592,N_24843,N_24943);
nor UO_593 (O_593,N_24875,N_24886);
xnor UO_594 (O_594,N_24997,N_24990);
or UO_595 (O_595,N_24876,N_24996);
or UO_596 (O_596,N_24929,N_24876);
or UO_597 (O_597,N_24907,N_24912);
and UO_598 (O_598,N_24997,N_24837);
xnor UO_599 (O_599,N_24837,N_24868);
nand UO_600 (O_600,N_24997,N_24994);
nor UO_601 (O_601,N_24955,N_24816);
nand UO_602 (O_602,N_24839,N_24819);
nand UO_603 (O_603,N_24927,N_24831);
nor UO_604 (O_604,N_24952,N_24867);
nand UO_605 (O_605,N_24938,N_24998);
nand UO_606 (O_606,N_24835,N_24918);
nand UO_607 (O_607,N_24991,N_24833);
and UO_608 (O_608,N_24881,N_24968);
nor UO_609 (O_609,N_24864,N_24803);
nor UO_610 (O_610,N_24962,N_24996);
xnor UO_611 (O_611,N_24883,N_24949);
and UO_612 (O_612,N_24926,N_24953);
xnor UO_613 (O_613,N_24998,N_24925);
nor UO_614 (O_614,N_24949,N_24955);
nor UO_615 (O_615,N_24883,N_24966);
xor UO_616 (O_616,N_24905,N_24870);
and UO_617 (O_617,N_24824,N_24958);
xor UO_618 (O_618,N_24819,N_24999);
xnor UO_619 (O_619,N_24874,N_24839);
xnor UO_620 (O_620,N_24893,N_24882);
xor UO_621 (O_621,N_24858,N_24819);
or UO_622 (O_622,N_24943,N_24851);
nor UO_623 (O_623,N_24954,N_24820);
xor UO_624 (O_624,N_24905,N_24831);
xnor UO_625 (O_625,N_24854,N_24840);
and UO_626 (O_626,N_24865,N_24964);
nand UO_627 (O_627,N_24902,N_24938);
nor UO_628 (O_628,N_24941,N_24829);
or UO_629 (O_629,N_24995,N_24998);
and UO_630 (O_630,N_24989,N_24852);
nor UO_631 (O_631,N_24943,N_24903);
xnor UO_632 (O_632,N_24955,N_24818);
or UO_633 (O_633,N_24982,N_24843);
and UO_634 (O_634,N_24852,N_24888);
and UO_635 (O_635,N_24888,N_24805);
xnor UO_636 (O_636,N_24979,N_24809);
nor UO_637 (O_637,N_24991,N_24835);
nand UO_638 (O_638,N_24891,N_24873);
xor UO_639 (O_639,N_24934,N_24999);
and UO_640 (O_640,N_24836,N_24879);
xnor UO_641 (O_641,N_24981,N_24974);
nor UO_642 (O_642,N_24847,N_24861);
or UO_643 (O_643,N_24886,N_24823);
xnor UO_644 (O_644,N_24957,N_24932);
nor UO_645 (O_645,N_24826,N_24841);
xnor UO_646 (O_646,N_24940,N_24864);
nand UO_647 (O_647,N_24997,N_24988);
or UO_648 (O_648,N_24877,N_24903);
or UO_649 (O_649,N_24996,N_24902);
or UO_650 (O_650,N_24908,N_24944);
xnor UO_651 (O_651,N_24800,N_24939);
nand UO_652 (O_652,N_24820,N_24837);
nand UO_653 (O_653,N_24866,N_24971);
and UO_654 (O_654,N_24885,N_24972);
nand UO_655 (O_655,N_24936,N_24825);
xnor UO_656 (O_656,N_24852,N_24800);
nand UO_657 (O_657,N_24957,N_24931);
or UO_658 (O_658,N_24986,N_24980);
and UO_659 (O_659,N_24987,N_24853);
nor UO_660 (O_660,N_24909,N_24902);
xnor UO_661 (O_661,N_24863,N_24897);
and UO_662 (O_662,N_24982,N_24911);
nand UO_663 (O_663,N_24992,N_24822);
nand UO_664 (O_664,N_24994,N_24931);
or UO_665 (O_665,N_24933,N_24927);
nand UO_666 (O_666,N_24847,N_24976);
nand UO_667 (O_667,N_24906,N_24877);
or UO_668 (O_668,N_24939,N_24954);
nor UO_669 (O_669,N_24811,N_24847);
and UO_670 (O_670,N_24864,N_24975);
nor UO_671 (O_671,N_24968,N_24911);
or UO_672 (O_672,N_24970,N_24959);
or UO_673 (O_673,N_24874,N_24953);
nand UO_674 (O_674,N_24903,N_24905);
nand UO_675 (O_675,N_24888,N_24820);
nor UO_676 (O_676,N_24808,N_24912);
and UO_677 (O_677,N_24859,N_24895);
nand UO_678 (O_678,N_24849,N_24981);
and UO_679 (O_679,N_24847,N_24988);
or UO_680 (O_680,N_24929,N_24975);
nor UO_681 (O_681,N_24905,N_24815);
or UO_682 (O_682,N_24840,N_24923);
nor UO_683 (O_683,N_24971,N_24823);
xnor UO_684 (O_684,N_24953,N_24815);
or UO_685 (O_685,N_24988,N_24816);
xor UO_686 (O_686,N_24899,N_24809);
nor UO_687 (O_687,N_24851,N_24921);
nand UO_688 (O_688,N_24917,N_24881);
nand UO_689 (O_689,N_24840,N_24801);
or UO_690 (O_690,N_24855,N_24917);
nor UO_691 (O_691,N_24999,N_24895);
and UO_692 (O_692,N_24892,N_24897);
xor UO_693 (O_693,N_24857,N_24993);
nand UO_694 (O_694,N_24858,N_24977);
or UO_695 (O_695,N_24814,N_24908);
xor UO_696 (O_696,N_24825,N_24893);
nand UO_697 (O_697,N_24884,N_24880);
nand UO_698 (O_698,N_24844,N_24805);
or UO_699 (O_699,N_24923,N_24932);
nor UO_700 (O_700,N_24800,N_24970);
or UO_701 (O_701,N_24811,N_24843);
and UO_702 (O_702,N_24896,N_24923);
or UO_703 (O_703,N_24868,N_24905);
and UO_704 (O_704,N_24879,N_24899);
nand UO_705 (O_705,N_24833,N_24926);
or UO_706 (O_706,N_24927,N_24837);
and UO_707 (O_707,N_24830,N_24884);
xor UO_708 (O_708,N_24885,N_24903);
or UO_709 (O_709,N_24833,N_24994);
or UO_710 (O_710,N_24903,N_24878);
nand UO_711 (O_711,N_24857,N_24916);
nand UO_712 (O_712,N_24966,N_24871);
and UO_713 (O_713,N_24965,N_24974);
or UO_714 (O_714,N_24923,N_24940);
nor UO_715 (O_715,N_24977,N_24852);
xor UO_716 (O_716,N_24982,N_24963);
xnor UO_717 (O_717,N_24846,N_24884);
nand UO_718 (O_718,N_24833,N_24921);
or UO_719 (O_719,N_24917,N_24920);
or UO_720 (O_720,N_24836,N_24808);
and UO_721 (O_721,N_24911,N_24899);
nor UO_722 (O_722,N_24914,N_24941);
or UO_723 (O_723,N_24885,N_24918);
nand UO_724 (O_724,N_24852,N_24847);
and UO_725 (O_725,N_24908,N_24812);
nor UO_726 (O_726,N_24900,N_24849);
nor UO_727 (O_727,N_24859,N_24972);
nand UO_728 (O_728,N_24817,N_24809);
nand UO_729 (O_729,N_24939,N_24995);
xnor UO_730 (O_730,N_24904,N_24836);
nor UO_731 (O_731,N_24809,N_24913);
xor UO_732 (O_732,N_24859,N_24894);
nor UO_733 (O_733,N_24986,N_24864);
and UO_734 (O_734,N_24959,N_24829);
nand UO_735 (O_735,N_24829,N_24891);
nor UO_736 (O_736,N_24889,N_24887);
xor UO_737 (O_737,N_24932,N_24901);
or UO_738 (O_738,N_24902,N_24816);
or UO_739 (O_739,N_24868,N_24886);
or UO_740 (O_740,N_24888,N_24864);
and UO_741 (O_741,N_24822,N_24916);
and UO_742 (O_742,N_24887,N_24885);
and UO_743 (O_743,N_24834,N_24872);
nand UO_744 (O_744,N_24896,N_24968);
or UO_745 (O_745,N_24946,N_24940);
nand UO_746 (O_746,N_24987,N_24801);
nand UO_747 (O_747,N_24953,N_24863);
or UO_748 (O_748,N_24947,N_24986);
and UO_749 (O_749,N_24897,N_24827);
or UO_750 (O_750,N_24833,N_24927);
or UO_751 (O_751,N_24869,N_24985);
nand UO_752 (O_752,N_24837,N_24910);
or UO_753 (O_753,N_24968,N_24917);
nand UO_754 (O_754,N_24816,N_24972);
and UO_755 (O_755,N_24858,N_24806);
nand UO_756 (O_756,N_24972,N_24925);
nand UO_757 (O_757,N_24953,N_24984);
nand UO_758 (O_758,N_24854,N_24963);
nand UO_759 (O_759,N_24988,N_24969);
and UO_760 (O_760,N_24983,N_24992);
nor UO_761 (O_761,N_24844,N_24931);
xor UO_762 (O_762,N_24908,N_24970);
or UO_763 (O_763,N_24899,N_24952);
or UO_764 (O_764,N_24922,N_24869);
nor UO_765 (O_765,N_24848,N_24839);
nor UO_766 (O_766,N_24879,N_24822);
xor UO_767 (O_767,N_24995,N_24946);
or UO_768 (O_768,N_24868,N_24828);
nor UO_769 (O_769,N_24980,N_24961);
nor UO_770 (O_770,N_24835,N_24919);
and UO_771 (O_771,N_24919,N_24831);
nand UO_772 (O_772,N_24886,N_24851);
xnor UO_773 (O_773,N_24859,N_24843);
or UO_774 (O_774,N_24958,N_24968);
xor UO_775 (O_775,N_24824,N_24865);
and UO_776 (O_776,N_24823,N_24962);
nor UO_777 (O_777,N_24823,N_24919);
and UO_778 (O_778,N_24949,N_24988);
xnor UO_779 (O_779,N_24885,N_24958);
nor UO_780 (O_780,N_24906,N_24984);
xor UO_781 (O_781,N_24865,N_24962);
or UO_782 (O_782,N_24948,N_24831);
xnor UO_783 (O_783,N_24936,N_24843);
nand UO_784 (O_784,N_24901,N_24916);
nand UO_785 (O_785,N_24905,N_24945);
nand UO_786 (O_786,N_24908,N_24824);
and UO_787 (O_787,N_24842,N_24882);
nor UO_788 (O_788,N_24882,N_24932);
nand UO_789 (O_789,N_24807,N_24940);
nor UO_790 (O_790,N_24888,N_24811);
nor UO_791 (O_791,N_24809,N_24822);
or UO_792 (O_792,N_24963,N_24977);
and UO_793 (O_793,N_24821,N_24857);
xnor UO_794 (O_794,N_24874,N_24851);
and UO_795 (O_795,N_24953,N_24871);
and UO_796 (O_796,N_24911,N_24897);
nand UO_797 (O_797,N_24834,N_24901);
nor UO_798 (O_798,N_24950,N_24890);
nor UO_799 (O_799,N_24883,N_24977);
xor UO_800 (O_800,N_24999,N_24908);
nand UO_801 (O_801,N_24820,N_24889);
xor UO_802 (O_802,N_24909,N_24806);
or UO_803 (O_803,N_24935,N_24997);
nor UO_804 (O_804,N_24954,N_24911);
nand UO_805 (O_805,N_24957,N_24890);
or UO_806 (O_806,N_24882,N_24956);
and UO_807 (O_807,N_24928,N_24945);
or UO_808 (O_808,N_24868,N_24831);
nor UO_809 (O_809,N_24966,N_24985);
nor UO_810 (O_810,N_24937,N_24960);
nand UO_811 (O_811,N_24929,N_24879);
nor UO_812 (O_812,N_24920,N_24902);
nor UO_813 (O_813,N_24998,N_24852);
xnor UO_814 (O_814,N_24933,N_24884);
nor UO_815 (O_815,N_24800,N_24922);
nand UO_816 (O_816,N_24854,N_24805);
and UO_817 (O_817,N_24998,N_24841);
nor UO_818 (O_818,N_24972,N_24933);
and UO_819 (O_819,N_24924,N_24933);
and UO_820 (O_820,N_24896,N_24869);
and UO_821 (O_821,N_24990,N_24934);
or UO_822 (O_822,N_24917,N_24974);
or UO_823 (O_823,N_24950,N_24802);
or UO_824 (O_824,N_24937,N_24824);
or UO_825 (O_825,N_24830,N_24942);
xnor UO_826 (O_826,N_24844,N_24970);
xor UO_827 (O_827,N_24960,N_24802);
nand UO_828 (O_828,N_24807,N_24840);
xnor UO_829 (O_829,N_24941,N_24875);
and UO_830 (O_830,N_24920,N_24986);
xnor UO_831 (O_831,N_24804,N_24867);
nand UO_832 (O_832,N_24889,N_24901);
and UO_833 (O_833,N_24890,N_24964);
nor UO_834 (O_834,N_24881,N_24824);
xnor UO_835 (O_835,N_24875,N_24969);
or UO_836 (O_836,N_24971,N_24827);
and UO_837 (O_837,N_24878,N_24923);
nand UO_838 (O_838,N_24893,N_24940);
nand UO_839 (O_839,N_24857,N_24925);
xor UO_840 (O_840,N_24929,N_24919);
nand UO_841 (O_841,N_24960,N_24835);
and UO_842 (O_842,N_24915,N_24866);
or UO_843 (O_843,N_24928,N_24963);
nand UO_844 (O_844,N_24904,N_24853);
or UO_845 (O_845,N_24994,N_24953);
or UO_846 (O_846,N_24910,N_24923);
nor UO_847 (O_847,N_24973,N_24906);
and UO_848 (O_848,N_24824,N_24955);
xnor UO_849 (O_849,N_24951,N_24950);
nand UO_850 (O_850,N_24934,N_24899);
nand UO_851 (O_851,N_24907,N_24851);
nor UO_852 (O_852,N_24979,N_24925);
nand UO_853 (O_853,N_24839,N_24904);
and UO_854 (O_854,N_24967,N_24983);
and UO_855 (O_855,N_24917,N_24800);
nor UO_856 (O_856,N_24974,N_24870);
xnor UO_857 (O_857,N_24832,N_24993);
xor UO_858 (O_858,N_24998,N_24862);
xor UO_859 (O_859,N_24910,N_24911);
xnor UO_860 (O_860,N_24978,N_24954);
and UO_861 (O_861,N_24809,N_24856);
or UO_862 (O_862,N_24943,N_24891);
xnor UO_863 (O_863,N_24820,N_24973);
and UO_864 (O_864,N_24933,N_24850);
and UO_865 (O_865,N_24852,N_24891);
or UO_866 (O_866,N_24925,N_24835);
or UO_867 (O_867,N_24995,N_24972);
xor UO_868 (O_868,N_24952,N_24859);
xor UO_869 (O_869,N_24881,N_24847);
or UO_870 (O_870,N_24962,N_24956);
nor UO_871 (O_871,N_24877,N_24800);
and UO_872 (O_872,N_24991,N_24908);
or UO_873 (O_873,N_24856,N_24929);
and UO_874 (O_874,N_24973,N_24920);
nand UO_875 (O_875,N_24865,N_24971);
or UO_876 (O_876,N_24939,N_24863);
xnor UO_877 (O_877,N_24856,N_24877);
nor UO_878 (O_878,N_24993,N_24871);
nor UO_879 (O_879,N_24916,N_24908);
and UO_880 (O_880,N_24837,N_24818);
nor UO_881 (O_881,N_24931,N_24974);
nand UO_882 (O_882,N_24931,N_24900);
xor UO_883 (O_883,N_24907,N_24896);
nand UO_884 (O_884,N_24925,N_24854);
nand UO_885 (O_885,N_24817,N_24898);
and UO_886 (O_886,N_24904,N_24921);
nand UO_887 (O_887,N_24925,N_24986);
nand UO_888 (O_888,N_24998,N_24964);
nor UO_889 (O_889,N_24919,N_24909);
and UO_890 (O_890,N_24847,N_24916);
and UO_891 (O_891,N_24863,N_24973);
and UO_892 (O_892,N_24832,N_24815);
nand UO_893 (O_893,N_24886,N_24836);
and UO_894 (O_894,N_24877,N_24802);
nand UO_895 (O_895,N_24996,N_24999);
and UO_896 (O_896,N_24952,N_24886);
and UO_897 (O_897,N_24978,N_24868);
nor UO_898 (O_898,N_24914,N_24885);
xnor UO_899 (O_899,N_24802,N_24976);
or UO_900 (O_900,N_24868,N_24847);
nor UO_901 (O_901,N_24843,N_24978);
nor UO_902 (O_902,N_24923,N_24920);
and UO_903 (O_903,N_24879,N_24809);
nor UO_904 (O_904,N_24996,N_24869);
or UO_905 (O_905,N_24879,N_24984);
and UO_906 (O_906,N_24965,N_24864);
xnor UO_907 (O_907,N_24901,N_24964);
or UO_908 (O_908,N_24812,N_24841);
nand UO_909 (O_909,N_24837,N_24844);
nor UO_910 (O_910,N_24956,N_24800);
or UO_911 (O_911,N_24838,N_24979);
or UO_912 (O_912,N_24929,N_24872);
and UO_913 (O_913,N_24972,N_24839);
nand UO_914 (O_914,N_24825,N_24999);
nand UO_915 (O_915,N_24962,N_24983);
and UO_916 (O_916,N_24994,N_24812);
xnor UO_917 (O_917,N_24975,N_24966);
or UO_918 (O_918,N_24962,N_24927);
or UO_919 (O_919,N_24993,N_24973);
nor UO_920 (O_920,N_24911,N_24859);
nand UO_921 (O_921,N_24982,N_24831);
nor UO_922 (O_922,N_24922,N_24969);
xnor UO_923 (O_923,N_24970,N_24845);
xnor UO_924 (O_924,N_24943,N_24962);
and UO_925 (O_925,N_24938,N_24834);
and UO_926 (O_926,N_24814,N_24909);
nor UO_927 (O_927,N_24959,N_24981);
xnor UO_928 (O_928,N_24986,N_24917);
nor UO_929 (O_929,N_24850,N_24846);
or UO_930 (O_930,N_24836,N_24857);
nand UO_931 (O_931,N_24849,N_24919);
xnor UO_932 (O_932,N_24858,N_24983);
or UO_933 (O_933,N_24862,N_24852);
nand UO_934 (O_934,N_24823,N_24936);
nand UO_935 (O_935,N_24892,N_24870);
nand UO_936 (O_936,N_24992,N_24933);
nor UO_937 (O_937,N_24973,N_24843);
nor UO_938 (O_938,N_24900,N_24850);
nand UO_939 (O_939,N_24864,N_24938);
and UO_940 (O_940,N_24999,N_24879);
nor UO_941 (O_941,N_24863,N_24961);
or UO_942 (O_942,N_24970,N_24934);
nand UO_943 (O_943,N_24939,N_24839);
or UO_944 (O_944,N_24859,N_24928);
or UO_945 (O_945,N_24847,N_24903);
or UO_946 (O_946,N_24993,N_24885);
nor UO_947 (O_947,N_24951,N_24842);
or UO_948 (O_948,N_24946,N_24837);
nor UO_949 (O_949,N_24975,N_24878);
nor UO_950 (O_950,N_24873,N_24964);
nor UO_951 (O_951,N_24879,N_24953);
xnor UO_952 (O_952,N_24824,N_24879);
nor UO_953 (O_953,N_24919,N_24949);
xor UO_954 (O_954,N_24990,N_24915);
or UO_955 (O_955,N_24907,N_24878);
nand UO_956 (O_956,N_24888,N_24878);
or UO_957 (O_957,N_24950,N_24895);
nor UO_958 (O_958,N_24925,N_24927);
or UO_959 (O_959,N_24909,N_24956);
or UO_960 (O_960,N_24914,N_24964);
or UO_961 (O_961,N_24916,N_24802);
nor UO_962 (O_962,N_24946,N_24914);
nand UO_963 (O_963,N_24990,N_24945);
nand UO_964 (O_964,N_24907,N_24830);
nor UO_965 (O_965,N_24968,N_24980);
and UO_966 (O_966,N_24900,N_24854);
or UO_967 (O_967,N_24998,N_24982);
and UO_968 (O_968,N_24803,N_24924);
xnor UO_969 (O_969,N_24905,N_24800);
nand UO_970 (O_970,N_24902,N_24857);
nor UO_971 (O_971,N_24906,N_24888);
nor UO_972 (O_972,N_24820,N_24873);
nor UO_973 (O_973,N_24850,N_24984);
and UO_974 (O_974,N_24966,N_24928);
nand UO_975 (O_975,N_24817,N_24813);
nor UO_976 (O_976,N_24868,N_24817);
nor UO_977 (O_977,N_24825,N_24897);
or UO_978 (O_978,N_24973,N_24979);
and UO_979 (O_979,N_24945,N_24880);
or UO_980 (O_980,N_24810,N_24974);
and UO_981 (O_981,N_24831,N_24872);
or UO_982 (O_982,N_24918,N_24964);
nor UO_983 (O_983,N_24911,N_24880);
and UO_984 (O_984,N_24879,N_24819);
nand UO_985 (O_985,N_24888,N_24917);
or UO_986 (O_986,N_24962,N_24944);
nor UO_987 (O_987,N_24837,N_24815);
nor UO_988 (O_988,N_24923,N_24946);
nand UO_989 (O_989,N_24886,N_24978);
xnor UO_990 (O_990,N_24859,N_24844);
or UO_991 (O_991,N_24836,N_24873);
or UO_992 (O_992,N_24995,N_24817);
xnor UO_993 (O_993,N_24885,N_24849);
or UO_994 (O_994,N_24844,N_24903);
nand UO_995 (O_995,N_24967,N_24921);
nand UO_996 (O_996,N_24804,N_24901);
xnor UO_997 (O_997,N_24810,N_24864);
and UO_998 (O_998,N_24808,N_24844);
or UO_999 (O_999,N_24918,N_24841);
nand UO_1000 (O_1000,N_24925,N_24875);
xnor UO_1001 (O_1001,N_24928,N_24911);
nor UO_1002 (O_1002,N_24946,N_24917);
nor UO_1003 (O_1003,N_24895,N_24966);
xor UO_1004 (O_1004,N_24969,N_24907);
nand UO_1005 (O_1005,N_24861,N_24858);
and UO_1006 (O_1006,N_24845,N_24868);
nor UO_1007 (O_1007,N_24927,N_24865);
and UO_1008 (O_1008,N_24948,N_24886);
xnor UO_1009 (O_1009,N_24843,N_24840);
and UO_1010 (O_1010,N_24946,N_24910);
and UO_1011 (O_1011,N_24913,N_24917);
xor UO_1012 (O_1012,N_24853,N_24848);
or UO_1013 (O_1013,N_24894,N_24865);
nor UO_1014 (O_1014,N_24893,N_24963);
nand UO_1015 (O_1015,N_24866,N_24825);
and UO_1016 (O_1016,N_24834,N_24836);
nor UO_1017 (O_1017,N_24853,N_24883);
nand UO_1018 (O_1018,N_24927,N_24874);
or UO_1019 (O_1019,N_24873,N_24850);
nand UO_1020 (O_1020,N_24870,N_24955);
or UO_1021 (O_1021,N_24877,N_24964);
or UO_1022 (O_1022,N_24976,N_24808);
xor UO_1023 (O_1023,N_24965,N_24910);
nor UO_1024 (O_1024,N_24808,N_24817);
nand UO_1025 (O_1025,N_24985,N_24988);
or UO_1026 (O_1026,N_24804,N_24817);
or UO_1027 (O_1027,N_24824,N_24856);
nor UO_1028 (O_1028,N_24856,N_24844);
and UO_1029 (O_1029,N_24987,N_24887);
or UO_1030 (O_1030,N_24820,N_24957);
nand UO_1031 (O_1031,N_24998,N_24818);
nor UO_1032 (O_1032,N_24986,N_24910);
xor UO_1033 (O_1033,N_24957,N_24938);
or UO_1034 (O_1034,N_24898,N_24929);
and UO_1035 (O_1035,N_24843,N_24950);
nor UO_1036 (O_1036,N_24908,N_24847);
nor UO_1037 (O_1037,N_24951,N_24835);
nand UO_1038 (O_1038,N_24861,N_24811);
nor UO_1039 (O_1039,N_24911,N_24940);
nand UO_1040 (O_1040,N_24852,N_24990);
xor UO_1041 (O_1041,N_24961,N_24912);
or UO_1042 (O_1042,N_24909,N_24810);
and UO_1043 (O_1043,N_24832,N_24886);
nor UO_1044 (O_1044,N_24996,N_24980);
xor UO_1045 (O_1045,N_24963,N_24905);
or UO_1046 (O_1046,N_24939,N_24898);
or UO_1047 (O_1047,N_24981,N_24924);
and UO_1048 (O_1048,N_24835,N_24820);
xnor UO_1049 (O_1049,N_24838,N_24974);
nand UO_1050 (O_1050,N_24842,N_24972);
nand UO_1051 (O_1051,N_24893,N_24802);
and UO_1052 (O_1052,N_24986,N_24902);
and UO_1053 (O_1053,N_24913,N_24858);
nor UO_1054 (O_1054,N_24810,N_24975);
nor UO_1055 (O_1055,N_24838,N_24956);
xor UO_1056 (O_1056,N_24972,N_24960);
nor UO_1057 (O_1057,N_24902,N_24854);
xor UO_1058 (O_1058,N_24940,N_24847);
nand UO_1059 (O_1059,N_24853,N_24943);
xnor UO_1060 (O_1060,N_24882,N_24921);
xnor UO_1061 (O_1061,N_24936,N_24973);
or UO_1062 (O_1062,N_24850,N_24871);
xor UO_1063 (O_1063,N_24809,N_24881);
and UO_1064 (O_1064,N_24920,N_24869);
xor UO_1065 (O_1065,N_24830,N_24922);
or UO_1066 (O_1066,N_24805,N_24850);
and UO_1067 (O_1067,N_24988,N_24905);
nand UO_1068 (O_1068,N_24846,N_24993);
nor UO_1069 (O_1069,N_24980,N_24921);
nand UO_1070 (O_1070,N_24959,N_24923);
and UO_1071 (O_1071,N_24954,N_24986);
nor UO_1072 (O_1072,N_24804,N_24825);
nor UO_1073 (O_1073,N_24845,N_24882);
xor UO_1074 (O_1074,N_24857,N_24987);
and UO_1075 (O_1075,N_24981,N_24955);
nand UO_1076 (O_1076,N_24876,N_24845);
nand UO_1077 (O_1077,N_24979,N_24870);
and UO_1078 (O_1078,N_24811,N_24830);
or UO_1079 (O_1079,N_24983,N_24980);
xnor UO_1080 (O_1080,N_24981,N_24971);
nand UO_1081 (O_1081,N_24801,N_24825);
or UO_1082 (O_1082,N_24989,N_24890);
xnor UO_1083 (O_1083,N_24856,N_24901);
xor UO_1084 (O_1084,N_24875,N_24948);
nand UO_1085 (O_1085,N_24824,N_24901);
or UO_1086 (O_1086,N_24914,N_24977);
xor UO_1087 (O_1087,N_24941,N_24919);
nor UO_1088 (O_1088,N_24926,N_24914);
nand UO_1089 (O_1089,N_24935,N_24981);
nor UO_1090 (O_1090,N_24902,N_24932);
and UO_1091 (O_1091,N_24854,N_24984);
nand UO_1092 (O_1092,N_24803,N_24928);
nor UO_1093 (O_1093,N_24810,N_24942);
xnor UO_1094 (O_1094,N_24936,N_24909);
xor UO_1095 (O_1095,N_24907,N_24856);
nand UO_1096 (O_1096,N_24930,N_24800);
nand UO_1097 (O_1097,N_24822,N_24982);
xor UO_1098 (O_1098,N_24961,N_24901);
xnor UO_1099 (O_1099,N_24817,N_24874);
nor UO_1100 (O_1100,N_24819,N_24994);
nand UO_1101 (O_1101,N_24959,N_24807);
or UO_1102 (O_1102,N_24846,N_24927);
xor UO_1103 (O_1103,N_24844,N_24895);
nand UO_1104 (O_1104,N_24891,N_24952);
nand UO_1105 (O_1105,N_24974,N_24963);
nor UO_1106 (O_1106,N_24828,N_24886);
and UO_1107 (O_1107,N_24966,N_24958);
and UO_1108 (O_1108,N_24866,N_24823);
and UO_1109 (O_1109,N_24969,N_24934);
and UO_1110 (O_1110,N_24852,N_24968);
nor UO_1111 (O_1111,N_24960,N_24913);
or UO_1112 (O_1112,N_24954,N_24992);
xnor UO_1113 (O_1113,N_24991,N_24914);
nand UO_1114 (O_1114,N_24865,N_24879);
nand UO_1115 (O_1115,N_24908,N_24815);
nand UO_1116 (O_1116,N_24971,N_24876);
or UO_1117 (O_1117,N_24969,N_24911);
xor UO_1118 (O_1118,N_24891,N_24885);
xnor UO_1119 (O_1119,N_24892,N_24951);
or UO_1120 (O_1120,N_24823,N_24863);
nor UO_1121 (O_1121,N_24864,N_24951);
and UO_1122 (O_1122,N_24824,N_24828);
xor UO_1123 (O_1123,N_24973,N_24893);
or UO_1124 (O_1124,N_24859,N_24998);
xnor UO_1125 (O_1125,N_24972,N_24958);
nor UO_1126 (O_1126,N_24919,N_24853);
xnor UO_1127 (O_1127,N_24984,N_24962);
and UO_1128 (O_1128,N_24992,N_24871);
or UO_1129 (O_1129,N_24853,N_24935);
or UO_1130 (O_1130,N_24833,N_24961);
xor UO_1131 (O_1131,N_24988,N_24806);
and UO_1132 (O_1132,N_24852,N_24933);
nand UO_1133 (O_1133,N_24848,N_24833);
nor UO_1134 (O_1134,N_24893,N_24843);
nor UO_1135 (O_1135,N_24824,N_24914);
or UO_1136 (O_1136,N_24926,N_24912);
xor UO_1137 (O_1137,N_24998,N_24924);
or UO_1138 (O_1138,N_24871,N_24965);
or UO_1139 (O_1139,N_24868,N_24995);
or UO_1140 (O_1140,N_24920,N_24988);
or UO_1141 (O_1141,N_24860,N_24828);
or UO_1142 (O_1142,N_24918,N_24803);
nor UO_1143 (O_1143,N_24819,N_24943);
nand UO_1144 (O_1144,N_24897,N_24809);
or UO_1145 (O_1145,N_24964,N_24919);
and UO_1146 (O_1146,N_24939,N_24882);
xnor UO_1147 (O_1147,N_24975,N_24834);
xnor UO_1148 (O_1148,N_24800,N_24979);
xor UO_1149 (O_1149,N_24913,N_24972);
nand UO_1150 (O_1150,N_24967,N_24846);
and UO_1151 (O_1151,N_24904,N_24899);
nand UO_1152 (O_1152,N_24836,N_24918);
or UO_1153 (O_1153,N_24871,N_24853);
nor UO_1154 (O_1154,N_24820,N_24829);
nor UO_1155 (O_1155,N_24827,N_24968);
nor UO_1156 (O_1156,N_24837,N_24969);
and UO_1157 (O_1157,N_24868,N_24909);
and UO_1158 (O_1158,N_24953,N_24987);
xnor UO_1159 (O_1159,N_24819,N_24835);
xnor UO_1160 (O_1160,N_24856,N_24918);
and UO_1161 (O_1161,N_24881,N_24936);
or UO_1162 (O_1162,N_24958,N_24830);
xnor UO_1163 (O_1163,N_24940,N_24853);
and UO_1164 (O_1164,N_24907,N_24956);
or UO_1165 (O_1165,N_24889,N_24819);
and UO_1166 (O_1166,N_24818,N_24812);
nand UO_1167 (O_1167,N_24967,N_24929);
nor UO_1168 (O_1168,N_24837,N_24853);
nor UO_1169 (O_1169,N_24991,N_24805);
nand UO_1170 (O_1170,N_24835,N_24866);
nand UO_1171 (O_1171,N_24973,N_24914);
nand UO_1172 (O_1172,N_24879,N_24886);
nor UO_1173 (O_1173,N_24995,N_24967);
nor UO_1174 (O_1174,N_24852,N_24985);
and UO_1175 (O_1175,N_24881,N_24918);
nand UO_1176 (O_1176,N_24993,N_24917);
nand UO_1177 (O_1177,N_24800,N_24882);
xor UO_1178 (O_1178,N_24970,N_24862);
and UO_1179 (O_1179,N_24885,N_24853);
or UO_1180 (O_1180,N_24853,N_24991);
nor UO_1181 (O_1181,N_24855,N_24888);
or UO_1182 (O_1182,N_24871,N_24951);
and UO_1183 (O_1183,N_24803,N_24828);
xor UO_1184 (O_1184,N_24889,N_24848);
or UO_1185 (O_1185,N_24831,N_24828);
xor UO_1186 (O_1186,N_24901,N_24809);
or UO_1187 (O_1187,N_24810,N_24995);
xnor UO_1188 (O_1188,N_24852,N_24807);
xnor UO_1189 (O_1189,N_24918,N_24898);
nor UO_1190 (O_1190,N_24881,N_24925);
xor UO_1191 (O_1191,N_24810,N_24970);
and UO_1192 (O_1192,N_24812,N_24832);
and UO_1193 (O_1193,N_24842,N_24865);
or UO_1194 (O_1194,N_24961,N_24864);
and UO_1195 (O_1195,N_24842,N_24867);
nand UO_1196 (O_1196,N_24989,N_24940);
nand UO_1197 (O_1197,N_24830,N_24889);
nand UO_1198 (O_1198,N_24898,N_24807);
nor UO_1199 (O_1199,N_24920,N_24955);
nor UO_1200 (O_1200,N_24803,N_24948);
xor UO_1201 (O_1201,N_24850,N_24976);
nand UO_1202 (O_1202,N_24830,N_24989);
nand UO_1203 (O_1203,N_24975,N_24968);
xor UO_1204 (O_1204,N_24885,N_24952);
nor UO_1205 (O_1205,N_24972,N_24923);
xnor UO_1206 (O_1206,N_24988,N_24939);
or UO_1207 (O_1207,N_24807,N_24969);
nor UO_1208 (O_1208,N_24950,N_24989);
or UO_1209 (O_1209,N_24810,N_24981);
nor UO_1210 (O_1210,N_24901,N_24807);
nor UO_1211 (O_1211,N_24902,N_24866);
nand UO_1212 (O_1212,N_24940,N_24908);
nand UO_1213 (O_1213,N_24959,N_24911);
nor UO_1214 (O_1214,N_24870,N_24810);
nand UO_1215 (O_1215,N_24995,N_24848);
nand UO_1216 (O_1216,N_24979,N_24885);
and UO_1217 (O_1217,N_24962,N_24841);
nand UO_1218 (O_1218,N_24943,N_24944);
nand UO_1219 (O_1219,N_24805,N_24820);
nand UO_1220 (O_1220,N_24841,N_24803);
and UO_1221 (O_1221,N_24842,N_24830);
or UO_1222 (O_1222,N_24884,N_24975);
and UO_1223 (O_1223,N_24880,N_24852);
xnor UO_1224 (O_1224,N_24853,N_24840);
and UO_1225 (O_1225,N_24908,N_24830);
or UO_1226 (O_1226,N_24922,N_24999);
xnor UO_1227 (O_1227,N_24804,N_24991);
nand UO_1228 (O_1228,N_24860,N_24975);
nand UO_1229 (O_1229,N_24918,N_24858);
and UO_1230 (O_1230,N_24916,N_24885);
nand UO_1231 (O_1231,N_24899,N_24861);
or UO_1232 (O_1232,N_24976,N_24951);
or UO_1233 (O_1233,N_24810,N_24972);
and UO_1234 (O_1234,N_24996,N_24873);
nor UO_1235 (O_1235,N_24808,N_24811);
and UO_1236 (O_1236,N_24897,N_24964);
and UO_1237 (O_1237,N_24949,N_24983);
or UO_1238 (O_1238,N_24837,N_24948);
and UO_1239 (O_1239,N_24983,N_24942);
nand UO_1240 (O_1240,N_24816,N_24989);
or UO_1241 (O_1241,N_24940,N_24883);
xnor UO_1242 (O_1242,N_24822,N_24959);
nor UO_1243 (O_1243,N_24915,N_24928);
and UO_1244 (O_1244,N_24845,N_24825);
xor UO_1245 (O_1245,N_24929,N_24930);
or UO_1246 (O_1246,N_24998,N_24842);
and UO_1247 (O_1247,N_24836,N_24972);
or UO_1248 (O_1248,N_24902,N_24910);
nand UO_1249 (O_1249,N_24822,N_24804);
nand UO_1250 (O_1250,N_24877,N_24897);
and UO_1251 (O_1251,N_24856,N_24994);
xor UO_1252 (O_1252,N_24932,N_24872);
nor UO_1253 (O_1253,N_24947,N_24859);
xnor UO_1254 (O_1254,N_24811,N_24919);
or UO_1255 (O_1255,N_24855,N_24989);
xor UO_1256 (O_1256,N_24903,N_24962);
and UO_1257 (O_1257,N_24977,N_24946);
and UO_1258 (O_1258,N_24904,N_24859);
and UO_1259 (O_1259,N_24818,N_24951);
or UO_1260 (O_1260,N_24988,N_24864);
xnor UO_1261 (O_1261,N_24992,N_24930);
nand UO_1262 (O_1262,N_24906,N_24889);
xor UO_1263 (O_1263,N_24832,N_24897);
nor UO_1264 (O_1264,N_24969,N_24831);
nor UO_1265 (O_1265,N_24808,N_24908);
nor UO_1266 (O_1266,N_24958,N_24809);
or UO_1267 (O_1267,N_24833,N_24992);
xor UO_1268 (O_1268,N_24976,N_24920);
nor UO_1269 (O_1269,N_24844,N_24989);
nor UO_1270 (O_1270,N_24942,N_24850);
nor UO_1271 (O_1271,N_24808,N_24878);
nor UO_1272 (O_1272,N_24825,N_24950);
and UO_1273 (O_1273,N_24815,N_24909);
and UO_1274 (O_1274,N_24949,N_24800);
xnor UO_1275 (O_1275,N_24810,N_24912);
or UO_1276 (O_1276,N_24869,N_24901);
nor UO_1277 (O_1277,N_24862,N_24973);
nand UO_1278 (O_1278,N_24992,N_24997);
nor UO_1279 (O_1279,N_24884,N_24888);
or UO_1280 (O_1280,N_24859,N_24847);
xnor UO_1281 (O_1281,N_24998,N_24984);
or UO_1282 (O_1282,N_24872,N_24916);
and UO_1283 (O_1283,N_24898,N_24852);
nand UO_1284 (O_1284,N_24947,N_24895);
xnor UO_1285 (O_1285,N_24849,N_24869);
xor UO_1286 (O_1286,N_24893,N_24807);
nand UO_1287 (O_1287,N_24935,N_24817);
nor UO_1288 (O_1288,N_24822,N_24817);
or UO_1289 (O_1289,N_24806,N_24801);
or UO_1290 (O_1290,N_24853,N_24952);
nor UO_1291 (O_1291,N_24889,N_24980);
and UO_1292 (O_1292,N_24850,N_24808);
nand UO_1293 (O_1293,N_24940,N_24877);
nand UO_1294 (O_1294,N_24984,N_24943);
xnor UO_1295 (O_1295,N_24890,N_24999);
and UO_1296 (O_1296,N_24867,N_24931);
nor UO_1297 (O_1297,N_24985,N_24891);
nor UO_1298 (O_1298,N_24971,N_24835);
or UO_1299 (O_1299,N_24958,N_24893);
nor UO_1300 (O_1300,N_24801,N_24903);
and UO_1301 (O_1301,N_24947,N_24897);
or UO_1302 (O_1302,N_24966,N_24969);
and UO_1303 (O_1303,N_24884,N_24988);
nand UO_1304 (O_1304,N_24825,N_24925);
nand UO_1305 (O_1305,N_24996,N_24845);
xnor UO_1306 (O_1306,N_24833,N_24917);
xnor UO_1307 (O_1307,N_24917,N_24999);
nand UO_1308 (O_1308,N_24903,N_24957);
xor UO_1309 (O_1309,N_24931,N_24807);
nand UO_1310 (O_1310,N_24921,N_24859);
and UO_1311 (O_1311,N_24986,N_24901);
or UO_1312 (O_1312,N_24921,N_24818);
xnor UO_1313 (O_1313,N_24811,N_24812);
or UO_1314 (O_1314,N_24883,N_24915);
nand UO_1315 (O_1315,N_24842,N_24928);
xor UO_1316 (O_1316,N_24952,N_24822);
nor UO_1317 (O_1317,N_24873,N_24898);
and UO_1318 (O_1318,N_24832,N_24861);
or UO_1319 (O_1319,N_24943,N_24916);
nor UO_1320 (O_1320,N_24938,N_24868);
xnor UO_1321 (O_1321,N_24940,N_24856);
and UO_1322 (O_1322,N_24957,N_24959);
nand UO_1323 (O_1323,N_24901,N_24990);
or UO_1324 (O_1324,N_24853,N_24977);
and UO_1325 (O_1325,N_24986,N_24903);
nor UO_1326 (O_1326,N_24819,N_24823);
and UO_1327 (O_1327,N_24817,N_24805);
nor UO_1328 (O_1328,N_24879,N_24915);
or UO_1329 (O_1329,N_24930,N_24981);
and UO_1330 (O_1330,N_24966,N_24933);
nand UO_1331 (O_1331,N_24869,N_24981);
xor UO_1332 (O_1332,N_24950,N_24815);
and UO_1333 (O_1333,N_24839,N_24865);
xnor UO_1334 (O_1334,N_24872,N_24927);
nor UO_1335 (O_1335,N_24942,N_24833);
nor UO_1336 (O_1336,N_24955,N_24872);
nand UO_1337 (O_1337,N_24891,N_24944);
xnor UO_1338 (O_1338,N_24881,N_24942);
nand UO_1339 (O_1339,N_24962,N_24854);
or UO_1340 (O_1340,N_24883,N_24982);
nand UO_1341 (O_1341,N_24861,N_24872);
xnor UO_1342 (O_1342,N_24813,N_24800);
xnor UO_1343 (O_1343,N_24986,N_24996);
nor UO_1344 (O_1344,N_24922,N_24827);
xor UO_1345 (O_1345,N_24898,N_24855);
nand UO_1346 (O_1346,N_24949,N_24965);
and UO_1347 (O_1347,N_24982,N_24995);
nor UO_1348 (O_1348,N_24801,N_24868);
or UO_1349 (O_1349,N_24848,N_24819);
and UO_1350 (O_1350,N_24912,N_24846);
and UO_1351 (O_1351,N_24851,N_24948);
or UO_1352 (O_1352,N_24933,N_24853);
and UO_1353 (O_1353,N_24915,N_24945);
or UO_1354 (O_1354,N_24860,N_24935);
nor UO_1355 (O_1355,N_24961,N_24992);
xor UO_1356 (O_1356,N_24922,N_24945);
nand UO_1357 (O_1357,N_24911,N_24943);
xor UO_1358 (O_1358,N_24949,N_24936);
nor UO_1359 (O_1359,N_24813,N_24945);
xnor UO_1360 (O_1360,N_24951,N_24927);
nor UO_1361 (O_1361,N_24958,N_24990);
or UO_1362 (O_1362,N_24955,N_24917);
xor UO_1363 (O_1363,N_24997,N_24970);
or UO_1364 (O_1364,N_24967,N_24884);
nand UO_1365 (O_1365,N_24972,N_24997);
and UO_1366 (O_1366,N_24920,N_24814);
or UO_1367 (O_1367,N_24989,N_24885);
nand UO_1368 (O_1368,N_24852,N_24958);
nand UO_1369 (O_1369,N_24854,N_24855);
and UO_1370 (O_1370,N_24875,N_24877);
xnor UO_1371 (O_1371,N_24933,N_24915);
or UO_1372 (O_1372,N_24975,N_24826);
xor UO_1373 (O_1373,N_24880,N_24902);
xor UO_1374 (O_1374,N_24887,N_24816);
and UO_1375 (O_1375,N_24804,N_24879);
and UO_1376 (O_1376,N_24982,N_24891);
or UO_1377 (O_1377,N_24821,N_24982);
xor UO_1378 (O_1378,N_24886,N_24878);
nand UO_1379 (O_1379,N_24956,N_24899);
xnor UO_1380 (O_1380,N_24891,N_24828);
xor UO_1381 (O_1381,N_24997,N_24934);
and UO_1382 (O_1382,N_24950,N_24851);
nand UO_1383 (O_1383,N_24903,N_24821);
or UO_1384 (O_1384,N_24839,N_24942);
xor UO_1385 (O_1385,N_24801,N_24837);
nor UO_1386 (O_1386,N_24814,N_24937);
xnor UO_1387 (O_1387,N_24815,N_24940);
xnor UO_1388 (O_1388,N_24834,N_24877);
nand UO_1389 (O_1389,N_24862,N_24856);
nor UO_1390 (O_1390,N_24869,N_24828);
xnor UO_1391 (O_1391,N_24923,N_24876);
or UO_1392 (O_1392,N_24801,N_24954);
or UO_1393 (O_1393,N_24833,N_24800);
and UO_1394 (O_1394,N_24924,N_24917);
nand UO_1395 (O_1395,N_24801,N_24846);
xor UO_1396 (O_1396,N_24923,N_24817);
and UO_1397 (O_1397,N_24850,N_24882);
nand UO_1398 (O_1398,N_24877,N_24805);
or UO_1399 (O_1399,N_24974,N_24978);
nand UO_1400 (O_1400,N_24842,N_24901);
or UO_1401 (O_1401,N_24926,N_24858);
or UO_1402 (O_1402,N_24829,N_24898);
or UO_1403 (O_1403,N_24958,N_24937);
or UO_1404 (O_1404,N_24829,N_24943);
nand UO_1405 (O_1405,N_24809,N_24877);
and UO_1406 (O_1406,N_24829,N_24870);
or UO_1407 (O_1407,N_24813,N_24832);
and UO_1408 (O_1408,N_24872,N_24804);
nor UO_1409 (O_1409,N_24862,N_24933);
nor UO_1410 (O_1410,N_24846,N_24854);
or UO_1411 (O_1411,N_24802,N_24959);
nor UO_1412 (O_1412,N_24889,N_24879);
or UO_1413 (O_1413,N_24916,N_24828);
xnor UO_1414 (O_1414,N_24911,N_24847);
xnor UO_1415 (O_1415,N_24973,N_24829);
nand UO_1416 (O_1416,N_24828,N_24813);
and UO_1417 (O_1417,N_24974,N_24843);
nor UO_1418 (O_1418,N_24971,N_24811);
xor UO_1419 (O_1419,N_24911,N_24874);
xnor UO_1420 (O_1420,N_24835,N_24908);
nor UO_1421 (O_1421,N_24861,N_24905);
nor UO_1422 (O_1422,N_24959,N_24872);
or UO_1423 (O_1423,N_24854,N_24994);
nor UO_1424 (O_1424,N_24857,N_24878);
or UO_1425 (O_1425,N_24907,N_24873);
xor UO_1426 (O_1426,N_24891,N_24879);
nand UO_1427 (O_1427,N_24874,N_24900);
or UO_1428 (O_1428,N_24895,N_24965);
nand UO_1429 (O_1429,N_24834,N_24808);
nor UO_1430 (O_1430,N_24832,N_24959);
or UO_1431 (O_1431,N_24916,N_24800);
xor UO_1432 (O_1432,N_24848,N_24818);
xnor UO_1433 (O_1433,N_24940,N_24839);
and UO_1434 (O_1434,N_24922,N_24946);
and UO_1435 (O_1435,N_24888,N_24899);
nand UO_1436 (O_1436,N_24832,N_24907);
nor UO_1437 (O_1437,N_24845,N_24864);
nor UO_1438 (O_1438,N_24966,N_24853);
nand UO_1439 (O_1439,N_24981,N_24992);
xor UO_1440 (O_1440,N_24917,N_24960);
nand UO_1441 (O_1441,N_24937,N_24976);
or UO_1442 (O_1442,N_24920,N_24867);
and UO_1443 (O_1443,N_24807,N_24834);
xor UO_1444 (O_1444,N_24851,N_24916);
or UO_1445 (O_1445,N_24949,N_24934);
xor UO_1446 (O_1446,N_24955,N_24821);
xor UO_1447 (O_1447,N_24853,N_24956);
nand UO_1448 (O_1448,N_24897,N_24841);
nor UO_1449 (O_1449,N_24947,N_24806);
nor UO_1450 (O_1450,N_24939,N_24974);
and UO_1451 (O_1451,N_24884,N_24987);
nor UO_1452 (O_1452,N_24933,N_24840);
xor UO_1453 (O_1453,N_24825,N_24957);
nand UO_1454 (O_1454,N_24871,N_24908);
nand UO_1455 (O_1455,N_24942,N_24961);
xor UO_1456 (O_1456,N_24968,N_24988);
nor UO_1457 (O_1457,N_24836,N_24956);
or UO_1458 (O_1458,N_24837,N_24893);
xor UO_1459 (O_1459,N_24907,N_24849);
and UO_1460 (O_1460,N_24865,N_24920);
nor UO_1461 (O_1461,N_24995,N_24912);
and UO_1462 (O_1462,N_24997,N_24939);
nand UO_1463 (O_1463,N_24981,N_24948);
and UO_1464 (O_1464,N_24950,N_24946);
and UO_1465 (O_1465,N_24949,N_24821);
or UO_1466 (O_1466,N_24885,N_24890);
xor UO_1467 (O_1467,N_24876,N_24841);
and UO_1468 (O_1468,N_24912,N_24975);
and UO_1469 (O_1469,N_24836,N_24822);
or UO_1470 (O_1470,N_24809,N_24838);
nor UO_1471 (O_1471,N_24909,N_24880);
xor UO_1472 (O_1472,N_24964,N_24905);
nor UO_1473 (O_1473,N_24899,N_24920);
and UO_1474 (O_1474,N_24934,N_24896);
or UO_1475 (O_1475,N_24966,N_24816);
xnor UO_1476 (O_1476,N_24864,N_24969);
and UO_1477 (O_1477,N_24991,N_24896);
nand UO_1478 (O_1478,N_24895,N_24875);
or UO_1479 (O_1479,N_24900,N_24866);
or UO_1480 (O_1480,N_24900,N_24890);
or UO_1481 (O_1481,N_24914,N_24818);
or UO_1482 (O_1482,N_24803,N_24871);
nor UO_1483 (O_1483,N_24964,N_24989);
xor UO_1484 (O_1484,N_24878,N_24838);
nor UO_1485 (O_1485,N_24974,N_24896);
nor UO_1486 (O_1486,N_24954,N_24828);
xor UO_1487 (O_1487,N_24818,N_24935);
nor UO_1488 (O_1488,N_24806,N_24847);
or UO_1489 (O_1489,N_24880,N_24975);
nor UO_1490 (O_1490,N_24999,N_24982);
or UO_1491 (O_1491,N_24834,N_24966);
and UO_1492 (O_1492,N_24953,N_24843);
or UO_1493 (O_1493,N_24820,N_24844);
nand UO_1494 (O_1494,N_24986,N_24990);
xnor UO_1495 (O_1495,N_24914,N_24966);
and UO_1496 (O_1496,N_24826,N_24876);
nor UO_1497 (O_1497,N_24978,N_24913);
nor UO_1498 (O_1498,N_24931,N_24883);
xnor UO_1499 (O_1499,N_24852,N_24863);
nand UO_1500 (O_1500,N_24998,N_24837);
nor UO_1501 (O_1501,N_24898,N_24890);
nor UO_1502 (O_1502,N_24933,N_24976);
nor UO_1503 (O_1503,N_24845,N_24946);
xor UO_1504 (O_1504,N_24924,N_24818);
or UO_1505 (O_1505,N_24927,N_24875);
nand UO_1506 (O_1506,N_24947,N_24832);
and UO_1507 (O_1507,N_24948,N_24977);
nor UO_1508 (O_1508,N_24802,N_24872);
or UO_1509 (O_1509,N_24982,N_24819);
and UO_1510 (O_1510,N_24863,N_24806);
and UO_1511 (O_1511,N_24956,N_24804);
and UO_1512 (O_1512,N_24968,N_24959);
nand UO_1513 (O_1513,N_24969,N_24984);
and UO_1514 (O_1514,N_24990,N_24833);
and UO_1515 (O_1515,N_24990,N_24936);
nor UO_1516 (O_1516,N_24856,N_24935);
and UO_1517 (O_1517,N_24975,N_24827);
and UO_1518 (O_1518,N_24923,N_24875);
nand UO_1519 (O_1519,N_24940,N_24944);
xnor UO_1520 (O_1520,N_24811,N_24828);
or UO_1521 (O_1521,N_24922,N_24935);
nand UO_1522 (O_1522,N_24924,N_24854);
or UO_1523 (O_1523,N_24903,N_24977);
xor UO_1524 (O_1524,N_24879,N_24979);
or UO_1525 (O_1525,N_24835,N_24903);
and UO_1526 (O_1526,N_24984,N_24898);
and UO_1527 (O_1527,N_24997,N_24892);
and UO_1528 (O_1528,N_24811,N_24914);
nor UO_1529 (O_1529,N_24889,N_24803);
nor UO_1530 (O_1530,N_24957,N_24884);
nor UO_1531 (O_1531,N_24825,N_24930);
and UO_1532 (O_1532,N_24827,N_24983);
xnor UO_1533 (O_1533,N_24912,N_24958);
or UO_1534 (O_1534,N_24919,N_24885);
xor UO_1535 (O_1535,N_24876,N_24880);
and UO_1536 (O_1536,N_24809,N_24935);
xor UO_1537 (O_1537,N_24988,N_24858);
and UO_1538 (O_1538,N_24869,N_24935);
or UO_1539 (O_1539,N_24981,N_24865);
or UO_1540 (O_1540,N_24952,N_24962);
and UO_1541 (O_1541,N_24912,N_24842);
xnor UO_1542 (O_1542,N_24885,N_24804);
or UO_1543 (O_1543,N_24803,N_24938);
and UO_1544 (O_1544,N_24905,N_24990);
xor UO_1545 (O_1545,N_24977,N_24890);
or UO_1546 (O_1546,N_24954,N_24884);
xnor UO_1547 (O_1547,N_24862,N_24950);
nand UO_1548 (O_1548,N_24827,N_24896);
or UO_1549 (O_1549,N_24813,N_24899);
xor UO_1550 (O_1550,N_24951,N_24969);
and UO_1551 (O_1551,N_24802,N_24913);
xnor UO_1552 (O_1552,N_24906,N_24810);
xnor UO_1553 (O_1553,N_24814,N_24856);
and UO_1554 (O_1554,N_24838,N_24830);
or UO_1555 (O_1555,N_24952,N_24939);
or UO_1556 (O_1556,N_24879,N_24992);
nand UO_1557 (O_1557,N_24893,N_24993);
or UO_1558 (O_1558,N_24825,N_24823);
or UO_1559 (O_1559,N_24859,N_24815);
or UO_1560 (O_1560,N_24957,N_24958);
or UO_1561 (O_1561,N_24831,N_24871);
or UO_1562 (O_1562,N_24953,N_24828);
nor UO_1563 (O_1563,N_24836,N_24867);
nor UO_1564 (O_1564,N_24937,N_24944);
xnor UO_1565 (O_1565,N_24942,N_24979);
or UO_1566 (O_1566,N_24897,N_24868);
nand UO_1567 (O_1567,N_24802,N_24919);
nor UO_1568 (O_1568,N_24829,N_24811);
nand UO_1569 (O_1569,N_24981,N_24912);
nor UO_1570 (O_1570,N_24941,N_24948);
nand UO_1571 (O_1571,N_24801,N_24871);
xnor UO_1572 (O_1572,N_24963,N_24904);
xnor UO_1573 (O_1573,N_24826,N_24999);
nand UO_1574 (O_1574,N_24878,N_24951);
and UO_1575 (O_1575,N_24896,N_24834);
nand UO_1576 (O_1576,N_24862,N_24964);
and UO_1577 (O_1577,N_24988,N_24959);
nor UO_1578 (O_1578,N_24967,N_24845);
nor UO_1579 (O_1579,N_24873,N_24897);
xor UO_1580 (O_1580,N_24934,N_24892);
or UO_1581 (O_1581,N_24852,N_24865);
xor UO_1582 (O_1582,N_24912,N_24892);
or UO_1583 (O_1583,N_24977,N_24975);
nand UO_1584 (O_1584,N_24944,N_24982);
nor UO_1585 (O_1585,N_24895,N_24986);
nand UO_1586 (O_1586,N_24972,N_24878);
and UO_1587 (O_1587,N_24913,N_24945);
nand UO_1588 (O_1588,N_24863,N_24881);
or UO_1589 (O_1589,N_24879,N_24864);
xnor UO_1590 (O_1590,N_24803,N_24857);
and UO_1591 (O_1591,N_24944,N_24973);
nand UO_1592 (O_1592,N_24987,N_24913);
nand UO_1593 (O_1593,N_24834,N_24837);
xor UO_1594 (O_1594,N_24973,N_24922);
and UO_1595 (O_1595,N_24898,N_24992);
nor UO_1596 (O_1596,N_24816,N_24860);
and UO_1597 (O_1597,N_24874,N_24837);
xor UO_1598 (O_1598,N_24955,N_24951);
nand UO_1599 (O_1599,N_24876,N_24897);
and UO_1600 (O_1600,N_24824,N_24810);
xor UO_1601 (O_1601,N_24929,N_24804);
and UO_1602 (O_1602,N_24953,N_24860);
xnor UO_1603 (O_1603,N_24819,N_24924);
xnor UO_1604 (O_1604,N_24990,N_24967);
xnor UO_1605 (O_1605,N_24980,N_24907);
xor UO_1606 (O_1606,N_24899,N_24817);
nand UO_1607 (O_1607,N_24872,N_24821);
nand UO_1608 (O_1608,N_24992,N_24867);
xnor UO_1609 (O_1609,N_24872,N_24890);
or UO_1610 (O_1610,N_24850,N_24963);
nor UO_1611 (O_1611,N_24999,N_24919);
xnor UO_1612 (O_1612,N_24921,N_24987);
xor UO_1613 (O_1613,N_24902,N_24842);
nor UO_1614 (O_1614,N_24925,N_24932);
nand UO_1615 (O_1615,N_24973,N_24960);
nor UO_1616 (O_1616,N_24943,N_24832);
and UO_1617 (O_1617,N_24817,N_24939);
and UO_1618 (O_1618,N_24945,N_24818);
or UO_1619 (O_1619,N_24889,N_24983);
and UO_1620 (O_1620,N_24884,N_24892);
xnor UO_1621 (O_1621,N_24986,N_24973);
or UO_1622 (O_1622,N_24837,N_24829);
or UO_1623 (O_1623,N_24969,N_24802);
nor UO_1624 (O_1624,N_24934,N_24974);
xnor UO_1625 (O_1625,N_24807,N_24987);
and UO_1626 (O_1626,N_24996,N_24807);
nor UO_1627 (O_1627,N_24809,N_24943);
nand UO_1628 (O_1628,N_24947,N_24949);
nand UO_1629 (O_1629,N_24872,N_24914);
xnor UO_1630 (O_1630,N_24961,N_24995);
xnor UO_1631 (O_1631,N_24951,N_24928);
nor UO_1632 (O_1632,N_24834,N_24895);
or UO_1633 (O_1633,N_24881,N_24976);
nor UO_1634 (O_1634,N_24929,N_24812);
nand UO_1635 (O_1635,N_24962,N_24904);
or UO_1636 (O_1636,N_24834,N_24883);
and UO_1637 (O_1637,N_24828,N_24871);
nor UO_1638 (O_1638,N_24953,N_24861);
and UO_1639 (O_1639,N_24959,N_24809);
nand UO_1640 (O_1640,N_24937,N_24945);
nand UO_1641 (O_1641,N_24831,N_24959);
nor UO_1642 (O_1642,N_24878,N_24846);
nand UO_1643 (O_1643,N_24991,N_24867);
xnor UO_1644 (O_1644,N_24851,N_24901);
nor UO_1645 (O_1645,N_24987,N_24985);
nand UO_1646 (O_1646,N_24904,N_24860);
or UO_1647 (O_1647,N_24960,N_24889);
or UO_1648 (O_1648,N_24939,N_24991);
xnor UO_1649 (O_1649,N_24823,N_24882);
or UO_1650 (O_1650,N_24837,N_24847);
xor UO_1651 (O_1651,N_24882,N_24912);
and UO_1652 (O_1652,N_24951,N_24844);
and UO_1653 (O_1653,N_24859,N_24887);
xor UO_1654 (O_1654,N_24982,N_24962);
xor UO_1655 (O_1655,N_24970,N_24938);
and UO_1656 (O_1656,N_24964,N_24912);
nor UO_1657 (O_1657,N_24907,N_24923);
nor UO_1658 (O_1658,N_24811,N_24983);
xnor UO_1659 (O_1659,N_24958,N_24817);
nand UO_1660 (O_1660,N_24924,N_24913);
or UO_1661 (O_1661,N_24837,N_24836);
nand UO_1662 (O_1662,N_24934,N_24853);
and UO_1663 (O_1663,N_24880,N_24815);
xor UO_1664 (O_1664,N_24951,N_24968);
xnor UO_1665 (O_1665,N_24978,N_24977);
nor UO_1666 (O_1666,N_24921,N_24893);
xor UO_1667 (O_1667,N_24869,N_24895);
or UO_1668 (O_1668,N_24887,N_24835);
nand UO_1669 (O_1669,N_24876,N_24819);
xor UO_1670 (O_1670,N_24939,N_24919);
nand UO_1671 (O_1671,N_24851,N_24975);
nand UO_1672 (O_1672,N_24987,N_24951);
nand UO_1673 (O_1673,N_24818,N_24887);
xor UO_1674 (O_1674,N_24917,N_24806);
xnor UO_1675 (O_1675,N_24877,N_24868);
nand UO_1676 (O_1676,N_24811,N_24856);
nand UO_1677 (O_1677,N_24997,N_24960);
xor UO_1678 (O_1678,N_24923,N_24860);
nor UO_1679 (O_1679,N_24974,N_24808);
nor UO_1680 (O_1680,N_24847,N_24938);
or UO_1681 (O_1681,N_24974,N_24830);
nand UO_1682 (O_1682,N_24810,N_24858);
xor UO_1683 (O_1683,N_24856,N_24850);
and UO_1684 (O_1684,N_24992,N_24950);
xor UO_1685 (O_1685,N_24990,N_24954);
xnor UO_1686 (O_1686,N_24860,N_24827);
xor UO_1687 (O_1687,N_24926,N_24884);
nor UO_1688 (O_1688,N_24886,N_24936);
xor UO_1689 (O_1689,N_24862,N_24940);
xor UO_1690 (O_1690,N_24921,N_24841);
or UO_1691 (O_1691,N_24897,N_24916);
and UO_1692 (O_1692,N_24926,N_24849);
nand UO_1693 (O_1693,N_24931,N_24831);
nor UO_1694 (O_1694,N_24961,N_24880);
and UO_1695 (O_1695,N_24983,N_24930);
nand UO_1696 (O_1696,N_24970,N_24896);
nand UO_1697 (O_1697,N_24912,N_24901);
nor UO_1698 (O_1698,N_24867,N_24872);
or UO_1699 (O_1699,N_24923,N_24877);
nor UO_1700 (O_1700,N_24907,N_24986);
or UO_1701 (O_1701,N_24992,N_24902);
or UO_1702 (O_1702,N_24824,N_24931);
nand UO_1703 (O_1703,N_24899,N_24883);
or UO_1704 (O_1704,N_24897,N_24891);
xor UO_1705 (O_1705,N_24939,N_24881);
nor UO_1706 (O_1706,N_24845,N_24952);
nor UO_1707 (O_1707,N_24937,N_24867);
nor UO_1708 (O_1708,N_24935,N_24910);
or UO_1709 (O_1709,N_24877,N_24931);
or UO_1710 (O_1710,N_24836,N_24999);
or UO_1711 (O_1711,N_24810,N_24862);
or UO_1712 (O_1712,N_24804,N_24931);
nand UO_1713 (O_1713,N_24823,N_24906);
xnor UO_1714 (O_1714,N_24960,N_24932);
xor UO_1715 (O_1715,N_24929,N_24912);
and UO_1716 (O_1716,N_24834,N_24944);
xnor UO_1717 (O_1717,N_24837,N_24934);
nor UO_1718 (O_1718,N_24834,N_24939);
nand UO_1719 (O_1719,N_24882,N_24890);
nor UO_1720 (O_1720,N_24837,N_24848);
and UO_1721 (O_1721,N_24831,N_24980);
nand UO_1722 (O_1722,N_24802,N_24812);
nand UO_1723 (O_1723,N_24945,N_24859);
nor UO_1724 (O_1724,N_24981,N_24947);
or UO_1725 (O_1725,N_24860,N_24911);
nand UO_1726 (O_1726,N_24852,N_24962);
nand UO_1727 (O_1727,N_24951,N_24989);
and UO_1728 (O_1728,N_24805,N_24938);
or UO_1729 (O_1729,N_24936,N_24805);
xnor UO_1730 (O_1730,N_24936,N_24913);
xor UO_1731 (O_1731,N_24923,N_24961);
or UO_1732 (O_1732,N_24970,N_24890);
nor UO_1733 (O_1733,N_24843,N_24980);
or UO_1734 (O_1734,N_24871,N_24822);
and UO_1735 (O_1735,N_24925,N_24892);
nand UO_1736 (O_1736,N_24818,N_24961);
nor UO_1737 (O_1737,N_24985,N_24817);
nor UO_1738 (O_1738,N_24855,N_24923);
nand UO_1739 (O_1739,N_24920,N_24866);
xnor UO_1740 (O_1740,N_24833,N_24981);
or UO_1741 (O_1741,N_24875,N_24973);
nor UO_1742 (O_1742,N_24824,N_24919);
or UO_1743 (O_1743,N_24851,N_24846);
xor UO_1744 (O_1744,N_24838,N_24988);
and UO_1745 (O_1745,N_24815,N_24885);
or UO_1746 (O_1746,N_24992,N_24966);
nand UO_1747 (O_1747,N_24906,N_24971);
nand UO_1748 (O_1748,N_24899,N_24830);
nor UO_1749 (O_1749,N_24889,N_24941);
or UO_1750 (O_1750,N_24968,N_24906);
xor UO_1751 (O_1751,N_24983,N_24909);
nand UO_1752 (O_1752,N_24887,N_24819);
or UO_1753 (O_1753,N_24992,N_24999);
xnor UO_1754 (O_1754,N_24840,N_24934);
or UO_1755 (O_1755,N_24881,N_24894);
or UO_1756 (O_1756,N_24919,N_24968);
nand UO_1757 (O_1757,N_24860,N_24819);
nor UO_1758 (O_1758,N_24831,N_24882);
and UO_1759 (O_1759,N_24808,N_24993);
or UO_1760 (O_1760,N_24909,N_24951);
or UO_1761 (O_1761,N_24883,N_24823);
nor UO_1762 (O_1762,N_24975,N_24865);
or UO_1763 (O_1763,N_24924,N_24839);
xor UO_1764 (O_1764,N_24989,N_24959);
nand UO_1765 (O_1765,N_24967,N_24819);
or UO_1766 (O_1766,N_24835,N_24852);
or UO_1767 (O_1767,N_24931,N_24976);
and UO_1768 (O_1768,N_24822,N_24920);
nor UO_1769 (O_1769,N_24986,N_24824);
xor UO_1770 (O_1770,N_24849,N_24991);
or UO_1771 (O_1771,N_24810,N_24919);
or UO_1772 (O_1772,N_24970,N_24880);
nor UO_1773 (O_1773,N_24856,N_24998);
or UO_1774 (O_1774,N_24827,N_24863);
or UO_1775 (O_1775,N_24886,N_24863);
xnor UO_1776 (O_1776,N_24961,N_24983);
nand UO_1777 (O_1777,N_24990,N_24977);
xnor UO_1778 (O_1778,N_24823,N_24846);
and UO_1779 (O_1779,N_24865,N_24988);
nand UO_1780 (O_1780,N_24948,N_24949);
nand UO_1781 (O_1781,N_24828,N_24984);
and UO_1782 (O_1782,N_24893,N_24920);
and UO_1783 (O_1783,N_24827,N_24889);
or UO_1784 (O_1784,N_24921,N_24846);
and UO_1785 (O_1785,N_24811,N_24878);
and UO_1786 (O_1786,N_24853,N_24859);
or UO_1787 (O_1787,N_24949,N_24953);
or UO_1788 (O_1788,N_24930,N_24976);
or UO_1789 (O_1789,N_24987,N_24957);
nor UO_1790 (O_1790,N_24894,N_24982);
and UO_1791 (O_1791,N_24861,N_24865);
nand UO_1792 (O_1792,N_24980,N_24872);
nor UO_1793 (O_1793,N_24972,N_24849);
nor UO_1794 (O_1794,N_24860,N_24843);
nand UO_1795 (O_1795,N_24882,N_24875);
nand UO_1796 (O_1796,N_24981,N_24958);
nand UO_1797 (O_1797,N_24900,N_24882);
nand UO_1798 (O_1798,N_24934,N_24947);
or UO_1799 (O_1799,N_24829,N_24885);
nor UO_1800 (O_1800,N_24859,N_24941);
or UO_1801 (O_1801,N_24804,N_24888);
or UO_1802 (O_1802,N_24835,N_24816);
nand UO_1803 (O_1803,N_24932,N_24949);
and UO_1804 (O_1804,N_24861,N_24814);
and UO_1805 (O_1805,N_24955,N_24866);
and UO_1806 (O_1806,N_24882,N_24980);
and UO_1807 (O_1807,N_24836,N_24992);
and UO_1808 (O_1808,N_24849,N_24925);
nor UO_1809 (O_1809,N_24845,N_24843);
or UO_1810 (O_1810,N_24935,N_24904);
or UO_1811 (O_1811,N_24895,N_24940);
or UO_1812 (O_1812,N_24847,N_24833);
nor UO_1813 (O_1813,N_24964,N_24902);
xor UO_1814 (O_1814,N_24867,N_24963);
nor UO_1815 (O_1815,N_24994,N_24987);
xor UO_1816 (O_1816,N_24859,N_24971);
nand UO_1817 (O_1817,N_24858,N_24960);
and UO_1818 (O_1818,N_24893,N_24972);
nor UO_1819 (O_1819,N_24878,N_24904);
nor UO_1820 (O_1820,N_24819,N_24988);
xor UO_1821 (O_1821,N_24907,N_24964);
and UO_1822 (O_1822,N_24913,N_24821);
or UO_1823 (O_1823,N_24965,N_24958);
or UO_1824 (O_1824,N_24883,N_24987);
nor UO_1825 (O_1825,N_24843,N_24802);
nand UO_1826 (O_1826,N_24916,N_24892);
and UO_1827 (O_1827,N_24958,N_24992);
and UO_1828 (O_1828,N_24897,N_24969);
or UO_1829 (O_1829,N_24865,N_24984);
and UO_1830 (O_1830,N_24818,N_24976);
or UO_1831 (O_1831,N_24950,N_24800);
nand UO_1832 (O_1832,N_24922,N_24835);
or UO_1833 (O_1833,N_24916,N_24984);
nor UO_1834 (O_1834,N_24848,N_24994);
nor UO_1835 (O_1835,N_24820,N_24899);
nor UO_1836 (O_1836,N_24942,N_24800);
nand UO_1837 (O_1837,N_24995,N_24866);
or UO_1838 (O_1838,N_24997,N_24984);
nand UO_1839 (O_1839,N_24893,N_24828);
or UO_1840 (O_1840,N_24820,N_24859);
xor UO_1841 (O_1841,N_24968,N_24816);
or UO_1842 (O_1842,N_24852,N_24931);
xor UO_1843 (O_1843,N_24813,N_24891);
and UO_1844 (O_1844,N_24972,N_24983);
nor UO_1845 (O_1845,N_24869,N_24958);
and UO_1846 (O_1846,N_24932,N_24952);
or UO_1847 (O_1847,N_24945,N_24888);
or UO_1848 (O_1848,N_24999,N_24986);
nand UO_1849 (O_1849,N_24887,N_24844);
and UO_1850 (O_1850,N_24839,N_24920);
or UO_1851 (O_1851,N_24809,N_24875);
or UO_1852 (O_1852,N_24861,N_24856);
nor UO_1853 (O_1853,N_24958,N_24950);
and UO_1854 (O_1854,N_24845,N_24957);
and UO_1855 (O_1855,N_24934,N_24882);
and UO_1856 (O_1856,N_24974,N_24865);
nand UO_1857 (O_1857,N_24981,N_24832);
xor UO_1858 (O_1858,N_24870,N_24958);
nor UO_1859 (O_1859,N_24872,N_24893);
nand UO_1860 (O_1860,N_24862,N_24913);
and UO_1861 (O_1861,N_24842,N_24917);
nor UO_1862 (O_1862,N_24971,N_24964);
and UO_1863 (O_1863,N_24874,N_24898);
and UO_1864 (O_1864,N_24958,N_24839);
and UO_1865 (O_1865,N_24813,N_24924);
or UO_1866 (O_1866,N_24928,N_24900);
nor UO_1867 (O_1867,N_24814,N_24921);
nand UO_1868 (O_1868,N_24972,N_24876);
xor UO_1869 (O_1869,N_24947,N_24876);
xnor UO_1870 (O_1870,N_24952,N_24807);
xnor UO_1871 (O_1871,N_24967,N_24820);
and UO_1872 (O_1872,N_24805,N_24984);
or UO_1873 (O_1873,N_24939,N_24831);
and UO_1874 (O_1874,N_24876,N_24807);
and UO_1875 (O_1875,N_24978,N_24837);
nor UO_1876 (O_1876,N_24928,N_24977);
nor UO_1877 (O_1877,N_24846,N_24825);
nand UO_1878 (O_1878,N_24817,N_24904);
nand UO_1879 (O_1879,N_24879,N_24853);
or UO_1880 (O_1880,N_24879,N_24878);
and UO_1881 (O_1881,N_24849,N_24995);
or UO_1882 (O_1882,N_24871,N_24864);
nand UO_1883 (O_1883,N_24949,N_24939);
xnor UO_1884 (O_1884,N_24927,N_24800);
xor UO_1885 (O_1885,N_24924,N_24849);
nand UO_1886 (O_1886,N_24946,N_24986);
and UO_1887 (O_1887,N_24927,N_24860);
nor UO_1888 (O_1888,N_24846,N_24963);
or UO_1889 (O_1889,N_24938,N_24996);
and UO_1890 (O_1890,N_24867,N_24887);
and UO_1891 (O_1891,N_24926,N_24960);
nand UO_1892 (O_1892,N_24946,N_24821);
and UO_1893 (O_1893,N_24941,N_24839);
xor UO_1894 (O_1894,N_24800,N_24887);
nor UO_1895 (O_1895,N_24824,N_24891);
xnor UO_1896 (O_1896,N_24850,N_24989);
or UO_1897 (O_1897,N_24968,N_24800);
and UO_1898 (O_1898,N_24866,N_24881);
or UO_1899 (O_1899,N_24939,N_24856);
and UO_1900 (O_1900,N_24843,N_24852);
or UO_1901 (O_1901,N_24821,N_24850);
or UO_1902 (O_1902,N_24928,N_24858);
and UO_1903 (O_1903,N_24904,N_24874);
nor UO_1904 (O_1904,N_24845,N_24872);
and UO_1905 (O_1905,N_24960,N_24923);
xnor UO_1906 (O_1906,N_24847,N_24948);
xor UO_1907 (O_1907,N_24805,N_24826);
xnor UO_1908 (O_1908,N_24818,N_24988);
and UO_1909 (O_1909,N_24918,N_24921);
nor UO_1910 (O_1910,N_24812,N_24806);
nor UO_1911 (O_1911,N_24998,N_24945);
or UO_1912 (O_1912,N_24894,N_24946);
or UO_1913 (O_1913,N_24893,N_24869);
xor UO_1914 (O_1914,N_24939,N_24942);
and UO_1915 (O_1915,N_24934,N_24945);
xor UO_1916 (O_1916,N_24839,N_24816);
xor UO_1917 (O_1917,N_24974,N_24854);
nor UO_1918 (O_1918,N_24960,N_24873);
nor UO_1919 (O_1919,N_24922,N_24994);
or UO_1920 (O_1920,N_24882,N_24852);
xnor UO_1921 (O_1921,N_24907,N_24965);
nor UO_1922 (O_1922,N_24826,N_24913);
and UO_1923 (O_1923,N_24844,N_24988);
and UO_1924 (O_1924,N_24893,N_24925);
xnor UO_1925 (O_1925,N_24878,N_24989);
nand UO_1926 (O_1926,N_24806,N_24901);
nand UO_1927 (O_1927,N_24832,N_24983);
or UO_1928 (O_1928,N_24943,N_24860);
xor UO_1929 (O_1929,N_24909,N_24972);
nor UO_1930 (O_1930,N_24950,N_24900);
or UO_1931 (O_1931,N_24814,N_24885);
or UO_1932 (O_1932,N_24837,N_24850);
nand UO_1933 (O_1933,N_24976,N_24845);
and UO_1934 (O_1934,N_24893,N_24930);
nor UO_1935 (O_1935,N_24873,N_24965);
or UO_1936 (O_1936,N_24954,N_24904);
and UO_1937 (O_1937,N_24832,N_24899);
and UO_1938 (O_1938,N_24834,N_24949);
or UO_1939 (O_1939,N_24974,N_24883);
or UO_1940 (O_1940,N_24892,N_24896);
and UO_1941 (O_1941,N_24954,N_24803);
and UO_1942 (O_1942,N_24851,N_24895);
and UO_1943 (O_1943,N_24946,N_24991);
or UO_1944 (O_1944,N_24876,N_24954);
and UO_1945 (O_1945,N_24813,N_24949);
xor UO_1946 (O_1946,N_24994,N_24945);
and UO_1947 (O_1947,N_24985,N_24983);
and UO_1948 (O_1948,N_24976,N_24806);
xor UO_1949 (O_1949,N_24864,N_24913);
or UO_1950 (O_1950,N_24962,N_24836);
nor UO_1951 (O_1951,N_24897,N_24834);
and UO_1952 (O_1952,N_24871,N_24902);
and UO_1953 (O_1953,N_24977,N_24828);
xnor UO_1954 (O_1954,N_24900,N_24945);
nor UO_1955 (O_1955,N_24896,N_24881);
and UO_1956 (O_1956,N_24934,N_24832);
and UO_1957 (O_1957,N_24839,N_24814);
nor UO_1958 (O_1958,N_24865,N_24805);
xor UO_1959 (O_1959,N_24946,N_24997);
and UO_1960 (O_1960,N_24835,N_24803);
or UO_1961 (O_1961,N_24976,N_24856);
nand UO_1962 (O_1962,N_24953,N_24948);
nand UO_1963 (O_1963,N_24957,N_24832);
or UO_1964 (O_1964,N_24831,N_24834);
xor UO_1965 (O_1965,N_24984,N_24806);
nand UO_1966 (O_1966,N_24855,N_24960);
nor UO_1967 (O_1967,N_24926,N_24906);
nor UO_1968 (O_1968,N_24924,N_24928);
or UO_1969 (O_1969,N_24976,N_24978);
and UO_1970 (O_1970,N_24840,N_24875);
and UO_1971 (O_1971,N_24898,N_24830);
nand UO_1972 (O_1972,N_24990,N_24978);
or UO_1973 (O_1973,N_24869,N_24802);
nor UO_1974 (O_1974,N_24868,N_24887);
or UO_1975 (O_1975,N_24986,N_24957);
or UO_1976 (O_1976,N_24941,N_24986);
nand UO_1977 (O_1977,N_24895,N_24939);
xnor UO_1978 (O_1978,N_24913,N_24886);
xor UO_1979 (O_1979,N_24918,N_24975);
or UO_1980 (O_1980,N_24851,N_24871);
and UO_1981 (O_1981,N_24865,N_24851);
xor UO_1982 (O_1982,N_24949,N_24941);
nor UO_1983 (O_1983,N_24990,N_24973);
nor UO_1984 (O_1984,N_24888,N_24997);
nand UO_1985 (O_1985,N_24968,N_24803);
nand UO_1986 (O_1986,N_24994,N_24802);
nor UO_1987 (O_1987,N_24944,N_24889);
xor UO_1988 (O_1988,N_24925,N_24938);
nand UO_1989 (O_1989,N_24875,N_24986);
nor UO_1990 (O_1990,N_24927,N_24965);
xnor UO_1991 (O_1991,N_24999,N_24838);
nand UO_1992 (O_1992,N_24847,N_24981);
and UO_1993 (O_1993,N_24968,N_24877);
and UO_1994 (O_1994,N_24867,N_24933);
and UO_1995 (O_1995,N_24909,N_24941);
xor UO_1996 (O_1996,N_24837,N_24990);
and UO_1997 (O_1997,N_24895,N_24853);
and UO_1998 (O_1998,N_24855,N_24881);
nand UO_1999 (O_1999,N_24910,N_24815);
nor UO_2000 (O_2000,N_24967,N_24808);
xnor UO_2001 (O_2001,N_24962,N_24965);
nand UO_2002 (O_2002,N_24955,N_24907);
or UO_2003 (O_2003,N_24854,N_24987);
xor UO_2004 (O_2004,N_24963,N_24809);
or UO_2005 (O_2005,N_24961,N_24840);
or UO_2006 (O_2006,N_24996,N_24947);
nand UO_2007 (O_2007,N_24919,N_24978);
nor UO_2008 (O_2008,N_24850,N_24987);
xnor UO_2009 (O_2009,N_24907,N_24970);
nor UO_2010 (O_2010,N_24828,N_24825);
or UO_2011 (O_2011,N_24824,N_24900);
nand UO_2012 (O_2012,N_24895,N_24856);
or UO_2013 (O_2013,N_24983,N_24870);
or UO_2014 (O_2014,N_24945,N_24946);
and UO_2015 (O_2015,N_24814,N_24846);
xnor UO_2016 (O_2016,N_24875,N_24887);
nor UO_2017 (O_2017,N_24843,N_24819);
or UO_2018 (O_2018,N_24848,N_24968);
or UO_2019 (O_2019,N_24965,N_24829);
nand UO_2020 (O_2020,N_24940,N_24894);
and UO_2021 (O_2021,N_24861,N_24977);
and UO_2022 (O_2022,N_24929,N_24936);
nor UO_2023 (O_2023,N_24979,N_24825);
nor UO_2024 (O_2024,N_24915,N_24953);
or UO_2025 (O_2025,N_24931,N_24984);
nor UO_2026 (O_2026,N_24952,N_24820);
xor UO_2027 (O_2027,N_24876,N_24935);
nor UO_2028 (O_2028,N_24936,N_24898);
xnor UO_2029 (O_2029,N_24843,N_24897);
nand UO_2030 (O_2030,N_24952,N_24970);
nand UO_2031 (O_2031,N_24853,N_24882);
nand UO_2032 (O_2032,N_24861,N_24873);
nor UO_2033 (O_2033,N_24842,N_24911);
nand UO_2034 (O_2034,N_24874,N_24827);
or UO_2035 (O_2035,N_24991,N_24905);
nor UO_2036 (O_2036,N_24932,N_24980);
nand UO_2037 (O_2037,N_24990,N_24839);
or UO_2038 (O_2038,N_24986,N_24927);
nand UO_2039 (O_2039,N_24968,N_24841);
xor UO_2040 (O_2040,N_24876,N_24951);
or UO_2041 (O_2041,N_24949,N_24833);
xor UO_2042 (O_2042,N_24883,N_24841);
or UO_2043 (O_2043,N_24967,N_24930);
and UO_2044 (O_2044,N_24899,N_24822);
xnor UO_2045 (O_2045,N_24984,N_24877);
nand UO_2046 (O_2046,N_24836,N_24884);
nor UO_2047 (O_2047,N_24845,N_24921);
nand UO_2048 (O_2048,N_24997,N_24811);
xnor UO_2049 (O_2049,N_24886,N_24859);
and UO_2050 (O_2050,N_24903,N_24945);
or UO_2051 (O_2051,N_24895,N_24961);
or UO_2052 (O_2052,N_24929,N_24950);
or UO_2053 (O_2053,N_24994,N_24949);
and UO_2054 (O_2054,N_24911,N_24932);
xor UO_2055 (O_2055,N_24886,N_24961);
nor UO_2056 (O_2056,N_24850,N_24838);
nand UO_2057 (O_2057,N_24993,N_24924);
xnor UO_2058 (O_2058,N_24951,N_24935);
nand UO_2059 (O_2059,N_24874,N_24905);
and UO_2060 (O_2060,N_24828,N_24930);
nand UO_2061 (O_2061,N_24841,N_24810);
xnor UO_2062 (O_2062,N_24802,N_24814);
nand UO_2063 (O_2063,N_24992,N_24901);
nand UO_2064 (O_2064,N_24820,N_24988);
or UO_2065 (O_2065,N_24833,N_24940);
nand UO_2066 (O_2066,N_24934,N_24890);
and UO_2067 (O_2067,N_24822,N_24949);
nand UO_2068 (O_2068,N_24843,N_24836);
and UO_2069 (O_2069,N_24909,N_24840);
and UO_2070 (O_2070,N_24889,N_24831);
nand UO_2071 (O_2071,N_24992,N_24824);
xnor UO_2072 (O_2072,N_24945,N_24800);
nand UO_2073 (O_2073,N_24990,N_24924);
nor UO_2074 (O_2074,N_24907,N_24863);
xor UO_2075 (O_2075,N_24965,N_24933);
and UO_2076 (O_2076,N_24930,N_24829);
nor UO_2077 (O_2077,N_24892,N_24837);
nand UO_2078 (O_2078,N_24922,N_24874);
xnor UO_2079 (O_2079,N_24930,N_24918);
nand UO_2080 (O_2080,N_24929,N_24937);
and UO_2081 (O_2081,N_24956,N_24840);
or UO_2082 (O_2082,N_24973,N_24933);
nand UO_2083 (O_2083,N_24971,N_24987);
nand UO_2084 (O_2084,N_24897,N_24980);
nand UO_2085 (O_2085,N_24832,N_24894);
xnor UO_2086 (O_2086,N_24943,N_24925);
nor UO_2087 (O_2087,N_24877,N_24845);
nor UO_2088 (O_2088,N_24834,N_24817);
nand UO_2089 (O_2089,N_24876,N_24800);
xnor UO_2090 (O_2090,N_24916,N_24835);
and UO_2091 (O_2091,N_24965,N_24862);
nor UO_2092 (O_2092,N_24902,N_24944);
and UO_2093 (O_2093,N_24996,N_24976);
and UO_2094 (O_2094,N_24941,N_24933);
and UO_2095 (O_2095,N_24826,N_24987);
or UO_2096 (O_2096,N_24988,N_24970);
nor UO_2097 (O_2097,N_24833,N_24873);
xor UO_2098 (O_2098,N_24820,N_24905);
or UO_2099 (O_2099,N_24884,N_24953);
nand UO_2100 (O_2100,N_24901,N_24899);
xnor UO_2101 (O_2101,N_24938,N_24948);
or UO_2102 (O_2102,N_24937,N_24917);
xor UO_2103 (O_2103,N_24981,N_24841);
nand UO_2104 (O_2104,N_24887,N_24855);
or UO_2105 (O_2105,N_24867,N_24893);
nand UO_2106 (O_2106,N_24878,N_24804);
or UO_2107 (O_2107,N_24805,N_24882);
and UO_2108 (O_2108,N_24975,N_24994);
nor UO_2109 (O_2109,N_24852,N_24987);
xnor UO_2110 (O_2110,N_24992,N_24916);
nor UO_2111 (O_2111,N_24981,N_24926);
or UO_2112 (O_2112,N_24836,N_24826);
or UO_2113 (O_2113,N_24808,N_24929);
nand UO_2114 (O_2114,N_24991,N_24952);
xor UO_2115 (O_2115,N_24845,N_24818);
xnor UO_2116 (O_2116,N_24878,N_24906);
nor UO_2117 (O_2117,N_24947,N_24880);
and UO_2118 (O_2118,N_24937,N_24983);
nor UO_2119 (O_2119,N_24992,N_24971);
nor UO_2120 (O_2120,N_24874,N_24862);
xnor UO_2121 (O_2121,N_24992,N_24839);
nor UO_2122 (O_2122,N_24830,N_24887);
nand UO_2123 (O_2123,N_24857,N_24893);
nand UO_2124 (O_2124,N_24906,N_24990);
nand UO_2125 (O_2125,N_24949,N_24979);
and UO_2126 (O_2126,N_24886,N_24937);
and UO_2127 (O_2127,N_24868,N_24958);
and UO_2128 (O_2128,N_24850,N_24804);
and UO_2129 (O_2129,N_24897,N_24856);
nand UO_2130 (O_2130,N_24942,N_24875);
nand UO_2131 (O_2131,N_24964,N_24852);
or UO_2132 (O_2132,N_24821,N_24984);
xor UO_2133 (O_2133,N_24859,N_24837);
or UO_2134 (O_2134,N_24878,N_24977);
xnor UO_2135 (O_2135,N_24829,N_24948);
and UO_2136 (O_2136,N_24842,N_24913);
nand UO_2137 (O_2137,N_24951,N_24982);
nor UO_2138 (O_2138,N_24823,N_24966);
nand UO_2139 (O_2139,N_24827,N_24872);
nand UO_2140 (O_2140,N_24988,N_24892);
nand UO_2141 (O_2141,N_24931,N_24963);
nor UO_2142 (O_2142,N_24973,N_24807);
nand UO_2143 (O_2143,N_24997,N_24809);
or UO_2144 (O_2144,N_24907,N_24871);
nor UO_2145 (O_2145,N_24896,N_24937);
or UO_2146 (O_2146,N_24859,N_24870);
and UO_2147 (O_2147,N_24838,N_24872);
nor UO_2148 (O_2148,N_24877,N_24938);
nor UO_2149 (O_2149,N_24978,N_24956);
or UO_2150 (O_2150,N_24882,N_24898);
and UO_2151 (O_2151,N_24817,N_24932);
nor UO_2152 (O_2152,N_24848,N_24938);
nor UO_2153 (O_2153,N_24883,N_24958);
xnor UO_2154 (O_2154,N_24802,N_24921);
or UO_2155 (O_2155,N_24821,N_24885);
nand UO_2156 (O_2156,N_24955,N_24895);
nand UO_2157 (O_2157,N_24919,N_24857);
nor UO_2158 (O_2158,N_24907,N_24909);
xor UO_2159 (O_2159,N_24926,N_24982);
nor UO_2160 (O_2160,N_24986,N_24856);
or UO_2161 (O_2161,N_24914,N_24899);
xor UO_2162 (O_2162,N_24814,N_24901);
nor UO_2163 (O_2163,N_24802,N_24894);
nand UO_2164 (O_2164,N_24879,N_24935);
or UO_2165 (O_2165,N_24876,N_24998);
or UO_2166 (O_2166,N_24886,N_24962);
or UO_2167 (O_2167,N_24922,N_24811);
or UO_2168 (O_2168,N_24953,N_24943);
or UO_2169 (O_2169,N_24872,N_24967);
xnor UO_2170 (O_2170,N_24878,N_24805);
nor UO_2171 (O_2171,N_24962,N_24800);
nand UO_2172 (O_2172,N_24802,N_24972);
xor UO_2173 (O_2173,N_24883,N_24838);
nor UO_2174 (O_2174,N_24877,N_24882);
and UO_2175 (O_2175,N_24810,N_24888);
nand UO_2176 (O_2176,N_24898,N_24914);
nand UO_2177 (O_2177,N_24959,N_24929);
xor UO_2178 (O_2178,N_24876,N_24961);
or UO_2179 (O_2179,N_24879,N_24994);
nor UO_2180 (O_2180,N_24814,N_24822);
and UO_2181 (O_2181,N_24808,N_24950);
xnor UO_2182 (O_2182,N_24896,N_24854);
or UO_2183 (O_2183,N_24813,N_24975);
and UO_2184 (O_2184,N_24922,N_24898);
nor UO_2185 (O_2185,N_24849,N_24946);
and UO_2186 (O_2186,N_24872,N_24986);
or UO_2187 (O_2187,N_24833,N_24812);
and UO_2188 (O_2188,N_24937,N_24835);
or UO_2189 (O_2189,N_24882,N_24927);
nor UO_2190 (O_2190,N_24981,N_24945);
xnor UO_2191 (O_2191,N_24822,N_24906);
nor UO_2192 (O_2192,N_24928,N_24893);
xor UO_2193 (O_2193,N_24825,N_24863);
nor UO_2194 (O_2194,N_24873,N_24917);
xnor UO_2195 (O_2195,N_24814,N_24999);
or UO_2196 (O_2196,N_24936,N_24801);
nand UO_2197 (O_2197,N_24923,N_24980);
xnor UO_2198 (O_2198,N_24801,N_24874);
nand UO_2199 (O_2199,N_24907,N_24882);
and UO_2200 (O_2200,N_24875,N_24893);
and UO_2201 (O_2201,N_24855,N_24832);
or UO_2202 (O_2202,N_24960,N_24966);
xor UO_2203 (O_2203,N_24839,N_24893);
nand UO_2204 (O_2204,N_24991,N_24825);
xor UO_2205 (O_2205,N_24824,N_24964);
nand UO_2206 (O_2206,N_24838,N_24856);
or UO_2207 (O_2207,N_24936,N_24972);
nand UO_2208 (O_2208,N_24900,N_24986);
or UO_2209 (O_2209,N_24912,N_24831);
or UO_2210 (O_2210,N_24908,N_24993);
nor UO_2211 (O_2211,N_24997,N_24846);
nor UO_2212 (O_2212,N_24844,N_24943);
xnor UO_2213 (O_2213,N_24853,N_24974);
xor UO_2214 (O_2214,N_24985,N_24938);
and UO_2215 (O_2215,N_24928,N_24873);
nor UO_2216 (O_2216,N_24982,N_24955);
nand UO_2217 (O_2217,N_24903,N_24933);
or UO_2218 (O_2218,N_24807,N_24941);
and UO_2219 (O_2219,N_24958,N_24820);
nor UO_2220 (O_2220,N_24888,N_24969);
nor UO_2221 (O_2221,N_24958,N_24933);
nor UO_2222 (O_2222,N_24969,N_24904);
or UO_2223 (O_2223,N_24918,N_24886);
or UO_2224 (O_2224,N_24918,N_24901);
nor UO_2225 (O_2225,N_24954,N_24833);
nor UO_2226 (O_2226,N_24961,N_24867);
nand UO_2227 (O_2227,N_24826,N_24849);
xor UO_2228 (O_2228,N_24952,N_24943);
xnor UO_2229 (O_2229,N_24933,N_24849);
nor UO_2230 (O_2230,N_24887,N_24902);
xnor UO_2231 (O_2231,N_24931,N_24828);
xor UO_2232 (O_2232,N_24845,N_24896);
or UO_2233 (O_2233,N_24837,N_24885);
nor UO_2234 (O_2234,N_24874,N_24943);
or UO_2235 (O_2235,N_24874,N_24893);
nand UO_2236 (O_2236,N_24904,N_24824);
or UO_2237 (O_2237,N_24806,N_24831);
or UO_2238 (O_2238,N_24886,N_24988);
and UO_2239 (O_2239,N_24851,N_24845);
or UO_2240 (O_2240,N_24855,N_24800);
and UO_2241 (O_2241,N_24977,N_24885);
nor UO_2242 (O_2242,N_24825,N_24840);
and UO_2243 (O_2243,N_24946,N_24828);
nor UO_2244 (O_2244,N_24899,N_24908);
nand UO_2245 (O_2245,N_24974,N_24952);
xor UO_2246 (O_2246,N_24821,N_24988);
or UO_2247 (O_2247,N_24905,N_24803);
nand UO_2248 (O_2248,N_24897,N_24803);
nor UO_2249 (O_2249,N_24903,N_24875);
nand UO_2250 (O_2250,N_24908,N_24851);
nand UO_2251 (O_2251,N_24835,N_24905);
and UO_2252 (O_2252,N_24800,N_24802);
and UO_2253 (O_2253,N_24942,N_24809);
nor UO_2254 (O_2254,N_24946,N_24956);
nand UO_2255 (O_2255,N_24950,N_24986);
nand UO_2256 (O_2256,N_24996,N_24943);
and UO_2257 (O_2257,N_24894,N_24942);
or UO_2258 (O_2258,N_24846,N_24863);
and UO_2259 (O_2259,N_24913,N_24853);
and UO_2260 (O_2260,N_24811,N_24900);
and UO_2261 (O_2261,N_24970,N_24874);
nand UO_2262 (O_2262,N_24989,N_24881);
xor UO_2263 (O_2263,N_24989,N_24915);
xnor UO_2264 (O_2264,N_24856,N_24878);
and UO_2265 (O_2265,N_24969,N_24999);
and UO_2266 (O_2266,N_24902,N_24849);
xnor UO_2267 (O_2267,N_24916,N_24813);
xor UO_2268 (O_2268,N_24981,N_24808);
nand UO_2269 (O_2269,N_24928,N_24836);
and UO_2270 (O_2270,N_24852,N_24969);
xnor UO_2271 (O_2271,N_24875,N_24904);
nor UO_2272 (O_2272,N_24825,N_24872);
nor UO_2273 (O_2273,N_24901,N_24928);
and UO_2274 (O_2274,N_24930,N_24936);
and UO_2275 (O_2275,N_24942,N_24832);
xnor UO_2276 (O_2276,N_24973,N_24927);
xnor UO_2277 (O_2277,N_24899,N_24816);
and UO_2278 (O_2278,N_24893,N_24922);
xnor UO_2279 (O_2279,N_24955,N_24921);
and UO_2280 (O_2280,N_24957,N_24869);
nand UO_2281 (O_2281,N_24853,N_24979);
or UO_2282 (O_2282,N_24996,N_24806);
nand UO_2283 (O_2283,N_24945,N_24980);
or UO_2284 (O_2284,N_24866,N_24977);
or UO_2285 (O_2285,N_24971,N_24878);
and UO_2286 (O_2286,N_24941,N_24962);
xnor UO_2287 (O_2287,N_24957,N_24859);
xor UO_2288 (O_2288,N_24828,N_24989);
nand UO_2289 (O_2289,N_24933,N_24865);
and UO_2290 (O_2290,N_24907,N_24886);
xnor UO_2291 (O_2291,N_24904,N_24882);
nor UO_2292 (O_2292,N_24910,N_24889);
xnor UO_2293 (O_2293,N_24900,N_24878);
nor UO_2294 (O_2294,N_24979,N_24857);
xnor UO_2295 (O_2295,N_24922,N_24826);
and UO_2296 (O_2296,N_24856,N_24993);
nor UO_2297 (O_2297,N_24834,N_24882);
nor UO_2298 (O_2298,N_24882,N_24917);
and UO_2299 (O_2299,N_24958,N_24962);
nor UO_2300 (O_2300,N_24987,N_24949);
or UO_2301 (O_2301,N_24818,N_24954);
nand UO_2302 (O_2302,N_24977,N_24981);
nand UO_2303 (O_2303,N_24869,N_24805);
xor UO_2304 (O_2304,N_24987,N_24972);
nand UO_2305 (O_2305,N_24859,N_24875);
nor UO_2306 (O_2306,N_24894,N_24830);
or UO_2307 (O_2307,N_24848,N_24945);
xor UO_2308 (O_2308,N_24812,N_24941);
nor UO_2309 (O_2309,N_24815,N_24853);
and UO_2310 (O_2310,N_24810,N_24847);
nand UO_2311 (O_2311,N_24882,N_24808);
xnor UO_2312 (O_2312,N_24899,N_24880);
or UO_2313 (O_2313,N_24848,N_24871);
and UO_2314 (O_2314,N_24821,N_24855);
or UO_2315 (O_2315,N_24830,N_24890);
xnor UO_2316 (O_2316,N_24939,N_24854);
nand UO_2317 (O_2317,N_24904,N_24958);
xnor UO_2318 (O_2318,N_24995,N_24965);
and UO_2319 (O_2319,N_24841,N_24958);
and UO_2320 (O_2320,N_24902,N_24829);
xor UO_2321 (O_2321,N_24985,N_24857);
and UO_2322 (O_2322,N_24942,N_24815);
nor UO_2323 (O_2323,N_24911,N_24901);
nand UO_2324 (O_2324,N_24857,N_24957);
and UO_2325 (O_2325,N_24912,N_24817);
xor UO_2326 (O_2326,N_24964,N_24868);
nor UO_2327 (O_2327,N_24908,N_24868);
nand UO_2328 (O_2328,N_24826,N_24895);
nor UO_2329 (O_2329,N_24804,N_24839);
xnor UO_2330 (O_2330,N_24946,N_24912);
nor UO_2331 (O_2331,N_24956,N_24950);
xor UO_2332 (O_2332,N_24970,N_24914);
xnor UO_2333 (O_2333,N_24840,N_24929);
and UO_2334 (O_2334,N_24893,N_24952);
nand UO_2335 (O_2335,N_24885,N_24934);
xnor UO_2336 (O_2336,N_24813,N_24888);
and UO_2337 (O_2337,N_24811,N_24968);
or UO_2338 (O_2338,N_24833,N_24881);
xor UO_2339 (O_2339,N_24890,N_24902);
and UO_2340 (O_2340,N_24907,N_24819);
nor UO_2341 (O_2341,N_24919,N_24884);
nand UO_2342 (O_2342,N_24819,N_24829);
nand UO_2343 (O_2343,N_24828,N_24973);
and UO_2344 (O_2344,N_24827,N_24935);
and UO_2345 (O_2345,N_24952,N_24810);
nor UO_2346 (O_2346,N_24802,N_24957);
nor UO_2347 (O_2347,N_24886,N_24814);
xor UO_2348 (O_2348,N_24825,N_24834);
or UO_2349 (O_2349,N_24853,N_24827);
or UO_2350 (O_2350,N_24800,N_24849);
and UO_2351 (O_2351,N_24918,N_24878);
nor UO_2352 (O_2352,N_24969,N_24986);
nand UO_2353 (O_2353,N_24884,N_24997);
and UO_2354 (O_2354,N_24962,N_24918);
xor UO_2355 (O_2355,N_24987,N_24814);
or UO_2356 (O_2356,N_24865,N_24860);
nor UO_2357 (O_2357,N_24814,N_24813);
nor UO_2358 (O_2358,N_24881,N_24992);
xnor UO_2359 (O_2359,N_24844,N_24912);
xnor UO_2360 (O_2360,N_24887,N_24974);
or UO_2361 (O_2361,N_24974,N_24918);
or UO_2362 (O_2362,N_24954,N_24817);
nor UO_2363 (O_2363,N_24894,N_24967);
xor UO_2364 (O_2364,N_24951,N_24933);
and UO_2365 (O_2365,N_24921,N_24924);
xor UO_2366 (O_2366,N_24828,N_24970);
or UO_2367 (O_2367,N_24945,N_24831);
nor UO_2368 (O_2368,N_24964,N_24973);
and UO_2369 (O_2369,N_24962,N_24988);
and UO_2370 (O_2370,N_24993,N_24878);
nand UO_2371 (O_2371,N_24968,N_24813);
and UO_2372 (O_2372,N_24859,N_24938);
or UO_2373 (O_2373,N_24990,N_24922);
and UO_2374 (O_2374,N_24925,N_24987);
nand UO_2375 (O_2375,N_24907,N_24902);
nand UO_2376 (O_2376,N_24872,N_24975);
nand UO_2377 (O_2377,N_24906,N_24989);
and UO_2378 (O_2378,N_24914,N_24955);
nor UO_2379 (O_2379,N_24907,N_24833);
nor UO_2380 (O_2380,N_24816,N_24936);
nand UO_2381 (O_2381,N_24864,N_24868);
or UO_2382 (O_2382,N_24922,N_24956);
and UO_2383 (O_2383,N_24865,N_24900);
nor UO_2384 (O_2384,N_24807,N_24880);
nand UO_2385 (O_2385,N_24836,N_24896);
or UO_2386 (O_2386,N_24821,N_24958);
xor UO_2387 (O_2387,N_24862,N_24835);
and UO_2388 (O_2388,N_24930,N_24885);
and UO_2389 (O_2389,N_24981,N_24957);
nand UO_2390 (O_2390,N_24890,N_24966);
nor UO_2391 (O_2391,N_24981,N_24978);
and UO_2392 (O_2392,N_24893,N_24841);
nand UO_2393 (O_2393,N_24804,N_24851);
nand UO_2394 (O_2394,N_24887,N_24918);
nand UO_2395 (O_2395,N_24928,N_24917);
xor UO_2396 (O_2396,N_24824,N_24897);
nor UO_2397 (O_2397,N_24849,N_24892);
nand UO_2398 (O_2398,N_24913,N_24827);
nand UO_2399 (O_2399,N_24804,N_24895);
and UO_2400 (O_2400,N_24887,N_24989);
and UO_2401 (O_2401,N_24869,N_24865);
nand UO_2402 (O_2402,N_24965,N_24852);
nor UO_2403 (O_2403,N_24901,N_24857);
xor UO_2404 (O_2404,N_24996,N_24824);
nand UO_2405 (O_2405,N_24921,N_24899);
nand UO_2406 (O_2406,N_24835,N_24942);
and UO_2407 (O_2407,N_24997,N_24963);
and UO_2408 (O_2408,N_24967,N_24881);
or UO_2409 (O_2409,N_24984,N_24986);
xor UO_2410 (O_2410,N_24949,N_24884);
nor UO_2411 (O_2411,N_24886,N_24822);
and UO_2412 (O_2412,N_24813,N_24939);
nor UO_2413 (O_2413,N_24924,N_24937);
and UO_2414 (O_2414,N_24847,N_24995);
and UO_2415 (O_2415,N_24937,N_24827);
nor UO_2416 (O_2416,N_24919,N_24969);
nand UO_2417 (O_2417,N_24830,N_24981);
nor UO_2418 (O_2418,N_24964,N_24955);
or UO_2419 (O_2419,N_24892,N_24813);
or UO_2420 (O_2420,N_24936,N_24905);
or UO_2421 (O_2421,N_24935,N_24871);
nor UO_2422 (O_2422,N_24873,N_24831);
xor UO_2423 (O_2423,N_24817,N_24819);
or UO_2424 (O_2424,N_24866,N_24886);
and UO_2425 (O_2425,N_24944,N_24848);
nor UO_2426 (O_2426,N_24972,N_24931);
xor UO_2427 (O_2427,N_24825,N_24992);
xnor UO_2428 (O_2428,N_24986,N_24943);
nor UO_2429 (O_2429,N_24930,N_24858);
and UO_2430 (O_2430,N_24898,N_24891);
nor UO_2431 (O_2431,N_24865,N_24864);
and UO_2432 (O_2432,N_24902,N_24845);
nand UO_2433 (O_2433,N_24907,N_24827);
xor UO_2434 (O_2434,N_24990,N_24927);
and UO_2435 (O_2435,N_24837,N_24814);
and UO_2436 (O_2436,N_24848,N_24988);
or UO_2437 (O_2437,N_24956,N_24806);
or UO_2438 (O_2438,N_24985,N_24935);
nor UO_2439 (O_2439,N_24932,N_24828);
nand UO_2440 (O_2440,N_24808,N_24856);
xor UO_2441 (O_2441,N_24858,N_24947);
nor UO_2442 (O_2442,N_24963,N_24857);
or UO_2443 (O_2443,N_24914,N_24903);
nand UO_2444 (O_2444,N_24966,N_24864);
and UO_2445 (O_2445,N_24922,N_24807);
nand UO_2446 (O_2446,N_24898,N_24977);
xnor UO_2447 (O_2447,N_24958,N_24864);
xnor UO_2448 (O_2448,N_24918,N_24808);
or UO_2449 (O_2449,N_24867,N_24901);
nor UO_2450 (O_2450,N_24931,N_24843);
nor UO_2451 (O_2451,N_24897,N_24975);
xnor UO_2452 (O_2452,N_24909,N_24901);
and UO_2453 (O_2453,N_24923,N_24887);
or UO_2454 (O_2454,N_24858,N_24900);
nor UO_2455 (O_2455,N_24816,N_24850);
nor UO_2456 (O_2456,N_24894,N_24976);
nand UO_2457 (O_2457,N_24985,N_24934);
and UO_2458 (O_2458,N_24851,N_24967);
or UO_2459 (O_2459,N_24831,N_24985);
nor UO_2460 (O_2460,N_24812,N_24922);
xnor UO_2461 (O_2461,N_24910,N_24953);
xnor UO_2462 (O_2462,N_24961,N_24855);
xnor UO_2463 (O_2463,N_24989,N_24873);
nand UO_2464 (O_2464,N_24809,N_24857);
nor UO_2465 (O_2465,N_24949,N_24986);
xor UO_2466 (O_2466,N_24946,N_24882);
nor UO_2467 (O_2467,N_24821,N_24936);
or UO_2468 (O_2468,N_24952,N_24866);
or UO_2469 (O_2469,N_24918,N_24900);
and UO_2470 (O_2470,N_24861,N_24885);
nor UO_2471 (O_2471,N_24957,N_24988);
or UO_2472 (O_2472,N_24976,N_24895);
and UO_2473 (O_2473,N_24986,N_24961);
nand UO_2474 (O_2474,N_24960,N_24847);
nand UO_2475 (O_2475,N_24976,N_24884);
or UO_2476 (O_2476,N_24809,N_24878);
or UO_2477 (O_2477,N_24994,N_24804);
or UO_2478 (O_2478,N_24853,N_24972);
or UO_2479 (O_2479,N_24804,N_24856);
and UO_2480 (O_2480,N_24950,N_24879);
and UO_2481 (O_2481,N_24812,N_24906);
or UO_2482 (O_2482,N_24817,N_24981);
or UO_2483 (O_2483,N_24841,N_24967);
xor UO_2484 (O_2484,N_24887,N_24968);
nor UO_2485 (O_2485,N_24871,N_24829);
xnor UO_2486 (O_2486,N_24967,N_24957);
nand UO_2487 (O_2487,N_24899,N_24951);
and UO_2488 (O_2488,N_24824,N_24875);
nor UO_2489 (O_2489,N_24802,N_24876);
and UO_2490 (O_2490,N_24947,N_24927);
xor UO_2491 (O_2491,N_24992,N_24979);
or UO_2492 (O_2492,N_24974,N_24851);
nand UO_2493 (O_2493,N_24981,N_24839);
or UO_2494 (O_2494,N_24975,N_24825);
or UO_2495 (O_2495,N_24864,N_24892);
and UO_2496 (O_2496,N_24943,N_24931);
nor UO_2497 (O_2497,N_24974,N_24989);
or UO_2498 (O_2498,N_24973,N_24937);
xor UO_2499 (O_2499,N_24878,N_24908);
xor UO_2500 (O_2500,N_24817,N_24905);
nand UO_2501 (O_2501,N_24868,N_24943);
nand UO_2502 (O_2502,N_24835,N_24931);
nor UO_2503 (O_2503,N_24870,N_24987);
nand UO_2504 (O_2504,N_24923,N_24895);
or UO_2505 (O_2505,N_24861,N_24995);
nor UO_2506 (O_2506,N_24920,N_24802);
nand UO_2507 (O_2507,N_24873,N_24998);
nand UO_2508 (O_2508,N_24932,N_24977);
or UO_2509 (O_2509,N_24967,N_24861);
xnor UO_2510 (O_2510,N_24874,N_24822);
xor UO_2511 (O_2511,N_24924,N_24922);
nand UO_2512 (O_2512,N_24868,N_24882);
nor UO_2513 (O_2513,N_24923,N_24811);
and UO_2514 (O_2514,N_24889,N_24801);
xnor UO_2515 (O_2515,N_24904,N_24938);
nor UO_2516 (O_2516,N_24871,N_24823);
nor UO_2517 (O_2517,N_24822,N_24905);
nor UO_2518 (O_2518,N_24906,N_24979);
or UO_2519 (O_2519,N_24912,N_24978);
or UO_2520 (O_2520,N_24932,N_24971);
xnor UO_2521 (O_2521,N_24855,N_24840);
or UO_2522 (O_2522,N_24957,N_24826);
xnor UO_2523 (O_2523,N_24843,N_24979);
and UO_2524 (O_2524,N_24801,N_24917);
nand UO_2525 (O_2525,N_24891,N_24908);
nor UO_2526 (O_2526,N_24999,N_24918);
nand UO_2527 (O_2527,N_24931,N_24947);
or UO_2528 (O_2528,N_24856,N_24960);
and UO_2529 (O_2529,N_24812,N_24886);
and UO_2530 (O_2530,N_24889,N_24854);
nand UO_2531 (O_2531,N_24885,N_24970);
nand UO_2532 (O_2532,N_24864,N_24973);
and UO_2533 (O_2533,N_24953,N_24921);
nor UO_2534 (O_2534,N_24826,N_24990);
or UO_2535 (O_2535,N_24967,N_24913);
nor UO_2536 (O_2536,N_24965,N_24832);
and UO_2537 (O_2537,N_24808,N_24812);
nor UO_2538 (O_2538,N_24838,N_24828);
or UO_2539 (O_2539,N_24891,N_24992);
or UO_2540 (O_2540,N_24870,N_24991);
nor UO_2541 (O_2541,N_24831,N_24910);
nor UO_2542 (O_2542,N_24982,N_24960);
nor UO_2543 (O_2543,N_24829,N_24862);
and UO_2544 (O_2544,N_24894,N_24965);
xnor UO_2545 (O_2545,N_24988,N_24916);
xor UO_2546 (O_2546,N_24918,N_24961);
and UO_2547 (O_2547,N_24901,N_24954);
xnor UO_2548 (O_2548,N_24925,N_24937);
nor UO_2549 (O_2549,N_24950,N_24964);
xor UO_2550 (O_2550,N_24926,N_24886);
nand UO_2551 (O_2551,N_24858,N_24946);
and UO_2552 (O_2552,N_24843,N_24896);
or UO_2553 (O_2553,N_24988,N_24934);
or UO_2554 (O_2554,N_24960,N_24974);
or UO_2555 (O_2555,N_24900,N_24868);
or UO_2556 (O_2556,N_24861,N_24910);
xnor UO_2557 (O_2557,N_24806,N_24867);
or UO_2558 (O_2558,N_24934,N_24839);
and UO_2559 (O_2559,N_24986,N_24810);
nor UO_2560 (O_2560,N_24907,N_24930);
nor UO_2561 (O_2561,N_24990,N_24858);
or UO_2562 (O_2562,N_24983,N_24802);
or UO_2563 (O_2563,N_24801,N_24827);
and UO_2564 (O_2564,N_24896,N_24821);
xor UO_2565 (O_2565,N_24886,N_24860);
nand UO_2566 (O_2566,N_24848,N_24908);
xor UO_2567 (O_2567,N_24989,N_24908);
xnor UO_2568 (O_2568,N_24927,N_24994);
nor UO_2569 (O_2569,N_24880,N_24926);
nand UO_2570 (O_2570,N_24962,N_24942);
xor UO_2571 (O_2571,N_24805,N_24895);
and UO_2572 (O_2572,N_24883,N_24816);
nand UO_2573 (O_2573,N_24840,N_24952);
xnor UO_2574 (O_2574,N_24903,N_24990);
nand UO_2575 (O_2575,N_24842,N_24989);
and UO_2576 (O_2576,N_24875,N_24851);
and UO_2577 (O_2577,N_24808,N_24896);
nand UO_2578 (O_2578,N_24958,N_24805);
and UO_2579 (O_2579,N_24917,N_24859);
xnor UO_2580 (O_2580,N_24844,N_24973);
nor UO_2581 (O_2581,N_24809,N_24950);
and UO_2582 (O_2582,N_24964,N_24863);
and UO_2583 (O_2583,N_24876,N_24866);
and UO_2584 (O_2584,N_24999,N_24830);
and UO_2585 (O_2585,N_24807,N_24801);
or UO_2586 (O_2586,N_24925,N_24993);
and UO_2587 (O_2587,N_24804,N_24818);
and UO_2588 (O_2588,N_24849,N_24899);
or UO_2589 (O_2589,N_24902,N_24952);
xor UO_2590 (O_2590,N_24889,N_24998);
nor UO_2591 (O_2591,N_24852,N_24939);
or UO_2592 (O_2592,N_24881,N_24873);
nor UO_2593 (O_2593,N_24940,N_24969);
and UO_2594 (O_2594,N_24987,N_24928);
or UO_2595 (O_2595,N_24926,N_24989);
nor UO_2596 (O_2596,N_24872,N_24887);
and UO_2597 (O_2597,N_24886,N_24985);
and UO_2598 (O_2598,N_24960,N_24914);
nor UO_2599 (O_2599,N_24816,N_24949);
and UO_2600 (O_2600,N_24906,N_24847);
nor UO_2601 (O_2601,N_24855,N_24951);
nor UO_2602 (O_2602,N_24814,N_24952);
and UO_2603 (O_2603,N_24916,N_24989);
xor UO_2604 (O_2604,N_24876,N_24840);
xor UO_2605 (O_2605,N_24955,N_24978);
nand UO_2606 (O_2606,N_24913,N_24856);
nor UO_2607 (O_2607,N_24988,N_24853);
xnor UO_2608 (O_2608,N_24813,N_24974);
and UO_2609 (O_2609,N_24823,N_24852);
or UO_2610 (O_2610,N_24922,N_24957);
nor UO_2611 (O_2611,N_24818,N_24925);
or UO_2612 (O_2612,N_24989,N_24847);
xnor UO_2613 (O_2613,N_24961,N_24914);
or UO_2614 (O_2614,N_24834,N_24879);
nand UO_2615 (O_2615,N_24818,N_24944);
and UO_2616 (O_2616,N_24941,N_24899);
or UO_2617 (O_2617,N_24943,N_24989);
or UO_2618 (O_2618,N_24846,N_24813);
and UO_2619 (O_2619,N_24890,N_24936);
or UO_2620 (O_2620,N_24866,N_24953);
xnor UO_2621 (O_2621,N_24801,N_24910);
nand UO_2622 (O_2622,N_24854,N_24848);
or UO_2623 (O_2623,N_24861,N_24943);
nand UO_2624 (O_2624,N_24831,N_24975);
nand UO_2625 (O_2625,N_24942,N_24997);
and UO_2626 (O_2626,N_24910,N_24825);
nor UO_2627 (O_2627,N_24825,N_24907);
or UO_2628 (O_2628,N_24993,N_24868);
xor UO_2629 (O_2629,N_24981,N_24956);
and UO_2630 (O_2630,N_24926,N_24951);
or UO_2631 (O_2631,N_24972,N_24975);
and UO_2632 (O_2632,N_24943,N_24827);
nand UO_2633 (O_2633,N_24919,N_24943);
nor UO_2634 (O_2634,N_24912,N_24845);
nor UO_2635 (O_2635,N_24809,N_24895);
nor UO_2636 (O_2636,N_24827,N_24982);
and UO_2637 (O_2637,N_24892,N_24941);
nand UO_2638 (O_2638,N_24875,N_24823);
and UO_2639 (O_2639,N_24800,N_24977);
xor UO_2640 (O_2640,N_24942,N_24843);
nor UO_2641 (O_2641,N_24990,N_24961);
and UO_2642 (O_2642,N_24833,N_24953);
and UO_2643 (O_2643,N_24997,N_24987);
nor UO_2644 (O_2644,N_24888,N_24865);
xnor UO_2645 (O_2645,N_24906,N_24838);
xnor UO_2646 (O_2646,N_24934,N_24858);
nor UO_2647 (O_2647,N_24860,N_24895);
or UO_2648 (O_2648,N_24860,N_24933);
nand UO_2649 (O_2649,N_24806,N_24861);
xor UO_2650 (O_2650,N_24910,N_24836);
nor UO_2651 (O_2651,N_24974,N_24823);
and UO_2652 (O_2652,N_24988,N_24929);
nor UO_2653 (O_2653,N_24869,N_24933);
nor UO_2654 (O_2654,N_24863,N_24870);
nor UO_2655 (O_2655,N_24897,N_24908);
nand UO_2656 (O_2656,N_24804,N_24864);
nand UO_2657 (O_2657,N_24862,N_24981);
nand UO_2658 (O_2658,N_24835,N_24802);
nand UO_2659 (O_2659,N_24998,N_24833);
and UO_2660 (O_2660,N_24940,N_24907);
and UO_2661 (O_2661,N_24987,N_24872);
nor UO_2662 (O_2662,N_24824,N_24993);
nor UO_2663 (O_2663,N_24910,N_24907);
nand UO_2664 (O_2664,N_24895,N_24803);
xor UO_2665 (O_2665,N_24841,N_24987);
and UO_2666 (O_2666,N_24861,N_24826);
or UO_2667 (O_2667,N_24869,N_24881);
or UO_2668 (O_2668,N_24939,N_24855);
or UO_2669 (O_2669,N_24840,N_24820);
nand UO_2670 (O_2670,N_24939,N_24888);
or UO_2671 (O_2671,N_24874,N_24976);
nor UO_2672 (O_2672,N_24975,N_24911);
or UO_2673 (O_2673,N_24815,N_24804);
nor UO_2674 (O_2674,N_24869,N_24824);
or UO_2675 (O_2675,N_24967,N_24869);
nand UO_2676 (O_2676,N_24962,N_24890);
xor UO_2677 (O_2677,N_24983,N_24852);
or UO_2678 (O_2678,N_24814,N_24812);
xnor UO_2679 (O_2679,N_24958,N_24858);
nand UO_2680 (O_2680,N_24831,N_24804);
or UO_2681 (O_2681,N_24996,N_24907);
and UO_2682 (O_2682,N_24812,N_24953);
or UO_2683 (O_2683,N_24954,N_24870);
nand UO_2684 (O_2684,N_24878,N_24999);
and UO_2685 (O_2685,N_24829,N_24844);
and UO_2686 (O_2686,N_24852,N_24948);
or UO_2687 (O_2687,N_24954,N_24984);
and UO_2688 (O_2688,N_24895,N_24828);
xor UO_2689 (O_2689,N_24970,N_24854);
nor UO_2690 (O_2690,N_24908,N_24983);
xor UO_2691 (O_2691,N_24910,N_24800);
nor UO_2692 (O_2692,N_24801,N_24820);
nor UO_2693 (O_2693,N_24978,N_24904);
xor UO_2694 (O_2694,N_24920,N_24927);
and UO_2695 (O_2695,N_24881,N_24877);
or UO_2696 (O_2696,N_24979,N_24970);
nand UO_2697 (O_2697,N_24810,N_24978);
nand UO_2698 (O_2698,N_24960,N_24897);
and UO_2699 (O_2699,N_24812,N_24835);
and UO_2700 (O_2700,N_24907,N_24917);
nor UO_2701 (O_2701,N_24890,N_24847);
nand UO_2702 (O_2702,N_24813,N_24964);
xnor UO_2703 (O_2703,N_24872,N_24888);
nand UO_2704 (O_2704,N_24990,N_24955);
and UO_2705 (O_2705,N_24947,N_24830);
xnor UO_2706 (O_2706,N_24814,N_24804);
xnor UO_2707 (O_2707,N_24828,N_24964);
xor UO_2708 (O_2708,N_24834,N_24909);
or UO_2709 (O_2709,N_24883,N_24969);
and UO_2710 (O_2710,N_24815,N_24842);
nand UO_2711 (O_2711,N_24901,N_24843);
xor UO_2712 (O_2712,N_24886,N_24837);
nand UO_2713 (O_2713,N_24906,N_24912);
xor UO_2714 (O_2714,N_24881,N_24984);
nor UO_2715 (O_2715,N_24818,N_24983);
and UO_2716 (O_2716,N_24988,N_24837);
or UO_2717 (O_2717,N_24810,N_24857);
nor UO_2718 (O_2718,N_24931,N_24988);
nand UO_2719 (O_2719,N_24872,N_24996);
nand UO_2720 (O_2720,N_24982,N_24816);
and UO_2721 (O_2721,N_24938,N_24965);
nand UO_2722 (O_2722,N_24889,N_24874);
nor UO_2723 (O_2723,N_24931,N_24840);
or UO_2724 (O_2724,N_24858,N_24908);
or UO_2725 (O_2725,N_24948,N_24975);
and UO_2726 (O_2726,N_24808,N_24861);
xor UO_2727 (O_2727,N_24854,N_24895);
nand UO_2728 (O_2728,N_24838,N_24888);
nor UO_2729 (O_2729,N_24865,N_24908);
xor UO_2730 (O_2730,N_24837,N_24846);
or UO_2731 (O_2731,N_24965,N_24954);
and UO_2732 (O_2732,N_24844,N_24980);
or UO_2733 (O_2733,N_24925,N_24846);
nand UO_2734 (O_2734,N_24911,N_24807);
nand UO_2735 (O_2735,N_24989,N_24836);
or UO_2736 (O_2736,N_24893,N_24890);
and UO_2737 (O_2737,N_24951,N_24834);
nand UO_2738 (O_2738,N_24916,N_24939);
nor UO_2739 (O_2739,N_24916,N_24931);
nand UO_2740 (O_2740,N_24838,N_24926);
nor UO_2741 (O_2741,N_24861,N_24884);
nand UO_2742 (O_2742,N_24976,N_24830);
or UO_2743 (O_2743,N_24946,N_24907);
xnor UO_2744 (O_2744,N_24811,N_24819);
xnor UO_2745 (O_2745,N_24834,N_24849);
and UO_2746 (O_2746,N_24935,N_24917);
xnor UO_2747 (O_2747,N_24949,N_24940);
xor UO_2748 (O_2748,N_24844,N_24853);
nor UO_2749 (O_2749,N_24847,N_24992);
xnor UO_2750 (O_2750,N_24945,N_24923);
and UO_2751 (O_2751,N_24872,N_24988);
xor UO_2752 (O_2752,N_24817,N_24962);
and UO_2753 (O_2753,N_24978,N_24802);
xor UO_2754 (O_2754,N_24867,N_24968);
and UO_2755 (O_2755,N_24938,N_24923);
or UO_2756 (O_2756,N_24957,N_24912);
nor UO_2757 (O_2757,N_24808,N_24889);
or UO_2758 (O_2758,N_24939,N_24905);
and UO_2759 (O_2759,N_24969,N_24810);
or UO_2760 (O_2760,N_24930,N_24902);
and UO_2761 (O_2761,N_24835,N_24809);
or UO_2762 (O_2762,N_24903,N_24887);
xor UO_2763 (O_2763,N_24806,N_24845);
and UO_2764 (O_2764,N_24848,N_24867);
and UO_2765 (O_2765,N_24915,N_24811);
nor UO_2766 (O_2766,N_24948,N_24912);
nand UO_2767 (O_2767,N_24954,N_24987);
or UO_2768 (O_2768,N_24936,N_24960);
nor UO_2769 (O_2769,N_24849,N_24985);
xor UO_2770 (O_2770,N_24829,N_24863);
xnor UO_2771 (O_2771,N_24966,N_24894);
and UO_2772 (O_2772,N_24937,N_24878);
nor UO_2773 (O_2773,N_24948,N_24811);
nand UO_2774 (O_2774,N_24863,N_24949);
nor UO_2775 (O_2775,N_24869,N_24841);
nor UO_2776 (O_2776,N_24890,N_24991);
nor UO_2777 (O_2777,N_24899,N_24805);
nor UO_2778 (O_2778,N_24938,N_24831);
nor UO_2779 (O_2779,N_24871,N_24874);
and UO_2780 (O_2780,N_24950,N_24898);
and UO_2781 (O_2781,N_24896,N_24806);
or UO_2782 (O_2782,N_24804,N_24917);
nand UO_2783 (O_2783,N_24990,N_24929);
nand UO_2784 (O_2784,N_24880,N_24960);
nand UO_2785 (O_2785,N_24840,N_24995);
and UO_2786 (O_2786,N_24888,N_24850);
nand UO_2787 (O_2787,N_24956,N_24851);
nor UO_2788 (O_2788,N_24907,N_24903);
and UO_2789 (O_2789,N_24806,N_24833);
xnor UO_2790 (O_2790,N_24894,N_24806);
nand UO_2791 (O_2791,N_24859,N_24996);
and UO_2792 (O_2792,N_24934,N_24940);
nand UO_2793 (O_2793,N_24933,N_24811);
xnor UO_2794 (O_2794,N_24931,N_24860);
nor UO_2795 (O_2795,N_24995,N_24942);
xnor UO_2796 (O_2796,N_24824,N_24982);
and UO_2797 (O_2797,N_24931,N_24977);
and UO_2798 (O_2798,N_24943,N_24859);
xnor UO_2799 (O_2799,N_24920,N_24845);
or UO_2800 (O_2800,N_24816,N_24819);
nand UO_2801 (O_2801,N_24867,N_24846);
and UO_2802 (O_2802,N_24921,N_24801);
nor UO_2803 (O_2803,N_24995,N_24842);
and UO_2804 (O_2804,N_24909,N_24985);
and UO_2805 (O_2805,N_24805,N_24822);
nand UO_2806 (O_2806,N_24854,N_24878);
nor UO_2807 (O_2807,N_24857,N_24802);
nor UO_2808 (O_2808,N_24953,N_24917);
nand UO_2809 (O_2809,N_24882,N_24981);
nand UO_2810 (O_2810,N_24810,N_24825);
nor UO_2811 (O_2811,N_24810,N_24891);
and UO_2812 (O_2812,N_24930,N_24939);
xor UO_2813 (O_2813,N_24959,N_24893);
nor UO_2814 (O_2814,N_24959,N_24868);
and UO_2815 (O_2815,N_24854,N_24814);
or UO_2816 (O_2816,N_24969,N_24980);
xnor UO_2817 (O_2817,N_24806,N_24885);
or UO_2818 (O_2818,N_24813,N_24921);
or UO_2819 (O_2819,N_24897,N_24934);
nor UO_2820 (O_2820,N_24881,N_24978);
or UO_2821 (O_2821,N_24904,N_24854);
nor UO_2822 (O_2822,N_24809,N_24854);
nand UO_2823 (O_2823,N_24878,N_24802);
or UO_2824 (O_2824,N_24836,N_24977);
nor UO_2825 (O_2825,N_24810,N_24811);
and UO_2826 (O_2826,N_24921,N_24844);
nand UO_2827 (O_2827,N_24800,N_24834);
xnor UO_2828 (O_2828,N_24902,N_24840);
xnor UO_2829 (O_2829,N_24931,N_24819);
nand UO_2830 (O_2830,N_24950,N_24876);
or UO_2831 (O_2831,N_24903,N_24908);
nor UO_2832 (O_2832,N_24943,N_24949);
and UO_2833 (O_2833,N_24970,N_24992);
nor UO_2834 (O_2834,N_24895,N_24896);
xnor UO_2835 (O_2835,N_24939,N_24943);
xnor UO_2836 (O_2836,N_24936,N_24964);
nor UO_2837 (O_2837,N_24970,N_24878);
nor UO_2838 (O_2838,N_24885,N_24825);
xnor UO_2839 (O_2839,N_24958,N_24913);
and UO_2840 (O_2840,N_24802,N_24968);
nand UO_2841 (O_2841,N_24894,N_24916);
nand UO_2842 (O_2842,N_24963,N_24914);
or UO_2843 (O_2843,N_24938,N_24954);
and UO_2844 (O_2844,N_24936,N_24926);
nand UO_2845 (O_2845,N_24865,N_24821);
xnor UO_2846 (O_2846,N_24832,N_24950);
and UO_2847 (O_2847,N_24843,N_24955);
xor UO_2848 (O_2848,N_24827,N_24929);
nor UO_2849 (O_2849,N_24918,N_24826);
xor UO_2850 (O_2850,N_24854,N_24914);
and UO_2851 (O_2851,N_24940,N_24880);
or UO_2852 (O_2852,N_24829,N_24961);
or UO_2853 (O_2853,N_24983,N_24807);
and UO_2854 (O_2854,N_24918,N_24948);
nand UO_2855 (O_2855,N_24828,N_24833);
and UO_2856 (O_2856,N_24879,N_24835);
or UO_2857 (O_2857,N_24947,N_24816);
xor UO_2858 (O_2858,N_24904,N_24883);
or UO_2859 (O_2859,N_24850,N_24802);
xnor UO_2860 (O_2860,N_24870,N_24847);
nand UO_2861 (O_2861,N_24903,N_24941);
xnor UO_2862 (O_2862,N_24942,N_24884);
and UO_2863 (O_2863,N_24993,N_24946);
xnor UO_2864 (O_2864,N_24809,N_24821);
or UO_2865 (O_2865,N_24886,N_24855);
and UO_2866 (O_2866,N_24947,N_24874);
nor UO_2867 (O_2867,N_24860,N_24966);
and UO_2868 (O_2868,N_24856,N_24999);
nand UO_2869 (O_2869,N_24922,N_24963);
xor UO_2870 (O_2870,N_24951,N_24814);
nand UO_2871 (O_2871,N_24927,N_24998);
nand UO_2872 (O_2872,N_24973,N_24858);
nand UO_2873 (O_2873,N_24907,N_24837);
and UO_2874 (O_2874,N_24828,N_24849);
and UO_2875 (O_2875,N_24827,N_24833);
nand UO_2876 (O_2876,N_24872,N_24990);
and UO_2877 (O_2877,N_24824,N_24883);
or UO_2878 (O_2878,N_24980,N_24938);
xor UO_2879 (O_2879,N_24966,N_24803);
and UO_2880 (O_2880,N_24977,N_24904);
nand UO_2881 (O_2881,N_24804,N_24843);
nand UO_2882 (O_2882,N_24840,N_24893);
nand UO_2883 (O_2883,N_24879,N_24806);
nand UO_2884 (O_2884,N_24819,N_24977);
nand UO_2885 (O_2885,N_24991,N_24801);
nand UO_2886 (O_2886,N_24958,N_24944);
nand UO_2887 (O_2887,N_24992,N_24980);
nor UO_2888 (O_2888,N_24969,N_24952);
xor UO_2889 (O_2889,N_24984,N_24927);
and UO_2890 (O_2890,N_24945,N_24950);
and UO_2891 (O_2891,N_24984,N_24848);
nand UO_2892 (O_2892,N_24804,N_24812);
or UO_2893 (O_2893,N_24919,N_24808);
nor UO_2894 (O_2894,N_24984,N_24843);
xor UO_2895 (O_2895,N_24919,N_24904);
nor UO_2896 (O_2896,N_24963,N_24882);
nor UO_2897 (O_2897,N_24840,N_24839);
nand UO_2898 (O_2898,N_24838,N_24812);
nand UO_2899 (O_2899,N_24890,N_24846);
nand UO_2900 (O_2900,N_24983,N_24844);
or UO_2901 (O_2901,N_24970,N_24835);
xnor UO_2902 (O_2902,N_24892,N_24851);
or UO_2903 (O_2903,N_24812,N_24961);
and UO_2904 (O_2904,N_24897,N_24807);
xor UO_2905 (O_2905,N_24806,N_24844);
nand UO_2906 (O_2906,N_24970,N_24913);
nor UO_2907 (O_2907,N_24831,N_24845);
and UO_2908 (O_2908,N_24807,N_24925);
or UO_2909 (O_2909,N_24903,N_24916);
xnor UO_2910 (O_2910,N_24892,N_24928);
or UO_2911 (O_2911,N_24985,N_24882);
xnor UO_2912 (O_2912,N_24906,N_24804);
and UO_2913 (O_2913,N_24920,N_24800);
nor UO_2914 (O_2914,N_24927,N_24818);
or UO_2915 (O_2915,N_24804,N_24862);
and UO_2916 (O_2916,N_24940,N_24919);
nand UO_2917 (O_2917,N_24903,N_24926);
xnor UO_2918 (O_2918,N_24930,N_24998);
or UO_2919 (O_2919,N_24803,N_24911);
and UO_2920 (O_2920,N_24856,N_24866);
nor UO_2921 (O_2921,N_24943,N_24892);
or UO_2922 (O_2922,N_24975,N_24818);
xor UO_2923 (O_2923,N_24951,N_24921);
or UO_2924 (O_2924,N_24949,N_24887);
xnor UO_2925 (O_2925,N_24956,N_24913);
xor UO_2926 (O_2926,N_24934,N_24820);
or UO_2927 (O_2927,N_24815,N_24886);
xor UO_2928 (O_2928,N_24829,N_24857);
and UO_2929 (O_2929,N_24967,N_24801);
nor UO_2930 (O_2930,N_24970,N_24817);
and UO_2931 (O_2931,N_24812,N_24815);
nor UO_2932 (O_2932,N_24991,N_24969);
xnor UO_2933 (O_2933,N_24931,N_24961);
xnor UO_2934 (O_2934,N_24813,N_24823);
or UO_2935 (O_2935,N_24847,N_24800);
and UO_2936 (O_2936,N_24935,N_24948);
nand UO_2937 (O_2937,N_24895,N_24920);
nand UO_2938 (O_2938,N_24867,N_24844);
and UO_2939 (O_2939,N_24826,N_24933);
and UO_2940 (O_2940,N_24979,N_24934);
and UO_2941 (O_2941,N_24869,N_24995);
nand UO_2942 (O_2942,N_24931,N_24882);
and UO_2943 (O_2943,N_24933,N_24814);
xnor UO_2944 (O_2944,N_24943,N_24922);
and UO_2945 (O_2945,N_24824,N_24888);
or UO_2946 (O_2946,N_24993,N_24820);
or UO_2947 (O_2947,N_24964,N_24872);
or UO_2948 (O_2948,N_24844,N_24933);
and UO_2949 (O_2949,N_24805,N_24902);
nand UO_2950 (O_2950,N_24939,N_24840);
or UO_2951 (O_2951,N_24825,N_24814);
xnor UO_2952 (O_2952,N_24918,N_24888);
nand UO_2953 (O_2953,N_24916,N_24926);
nand UO_2954 (O_2954,N_24984,N_24908);
nand UO_2955 (O_2955,N_24847,N_24943);
nand UO_2956 (O_2956,N_24832,N_24863);
or UO_2957 (O_2957,N_24830,N_24882);
or UO_2958 (O_2958,N_24920,N_24880);
nand UO_2959 (O_2959,N_24980,N_24875);
or UO_2960 (O_2960,N_24877,N_24915);
xor UO_2961 (O_2961,N_24911,N_24937);
nor UO_2962 (O_2962,N_24851,N_24877);
nor UO_2963 (O_2963,N_24859,N_24964);
nand UO_2964 (O_2964,N_24963,N_24926);
and UO_2965 (O_2965,N_24823,N_24984);
and UO_2966 (O_2966,N_24863,N_24854);
nand UO_2967 (O_2967,N_24891,N_24820);
nor UO_2968 (O_2968,N_24896,N_24801);
or UO_2969 (O_2969,N_24925,N_24948);
nor UO_2970 (O_2970,N_24883,N_24937);
and UO_2971 (O_2971,N_24836,N_24924);
nand UO_2972 (O_2972,N_24858,N_24844);
xnor UO_2973 (O_2973,N_24850,N_24945);
nand UO_2974 (O_2974,N_24825,N_24830);
nand UO_2975 (O_2975,N_24931,N_24919);
nand UO_2976 (O_2976,N_24852,N_24830);
or UO_2977 (O_2977,N_24920,N_24811);
xnor UO_2978 (O_2978,N_24970,N_24864);
or UO_2979 (O_2979,N_24970,N_24941);
nor UO_2980 (O_2980,N_24990,N_24907);
nand UO_2981 (O_2981,N_24806,N_24946);
or UO_2982 (O_2982,N_24943,N_24908);
or UO_2983 (O_2983,N_24980,N_24859);
nor UO_2984 (O_2984,N_24829,N_24908);
or UO_2985 (O_2985,N_24849,N_24805);
nor UO_2986 (O_2986,N_24833,N_24844);
and UO_2987 (O_2987,N_24853,N_24845);
or UO_2988 (O_2988,N_24839,N_24952);
nand UO_2989 (O_2989,N_24930,N_24975);
nand UO_2990 (O_2990,N_24883,N_24890);
nand UO_2991 (O_2991,N_24888,N_24812);
nand UO_2992 (O_2992,N_24936,N_24996);
nor UO_2993 (O_2993,N_24959,N_24961);
or UO_2994 (O_2994,N_24950,N_24829);
or UO_2995 (O_2995,N_24814,N_24902);
and UO_2996 (O_2996,N_24983,N_24853);
and UO_2997 (O_2997,N_24963,N_24814);
xor UO_2998 (O_2998,N_24931,N_24832);
and UO_2999 (O_2999,N_24928,N_24943);
endmodule