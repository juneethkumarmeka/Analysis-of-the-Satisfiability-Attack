module basic_750_5000_1000_5_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_33,In_512);
xnor U1 (N_1,In_17,In_349);
nor U2 (N_2,In_115,In_620);
nand U3 (N_3,In_709,In_538);
or U4 (N_4,In_467,In_505);
and U5 (N_5,In_70,In_734);
and U6 (N_6,In_180,In_317);
or U7 (N_7,In_314,In_188);
nand U8 (N_8,In_657,In_112);
or U9 (N_9,In_143,In_627);
or U10 (N_10,In_700,In_743);
nand U11 (N_11,In_660,In_581);
and U12 (N_12,In_378,In_334);
or U13 (N_13,In_219,In_706);
and U14 (N_14,In_47,In_663);
nand U15 (N_15,In_533,In_511);
or U16 (N_16,In_38,In_123);
or U17 (N_17,In_636,In_465);
and U18 (N_18,In_719,In_4);
nand U19 (N_19,In_152,In_52);
nand U20 (N_20,In_128,In_56);
xnor U21 (N_21,In_428,In_655);
nor U22 (N_22,In_102,In_237);
and U23 (N_23,In_583,In_500);
and U24 (N_24,In_479,In_483);
and U25 (N_25,In_28,In_517);
nand U26 (N_26,In_269,In_76);
nor U27 (N_27,In_560,In_726);
nand U28 (N_28,In_279,In_599);
or U29 (N_29,In_498,In_430);
and U30 (N_30,In_255,In_258);
and U31 (N_31,In_194,In_11);
or U32 (N_32,In_699,In_578);
and U33 (N_33,In_118,In_189);
nand U34 (N_34,In_714,In_679);
nor U35 (N_35,In_166,In_526);
nor U36 (N_36,In_216,In_354);
nand U37 (N_37,In_649,In_594);
nor U38 (N_38,In_631,In_531);
or U39 (N_39,In_360,In_674);
and U40 (N_40,In_515,In_420);
and U41 (N_41,In_294,In_292);
and U42 (N_42,In_329,In_617);
and U43 (N_43,In_528,In_43);
and U44 (N_44,In_235,In_400);
nor U45 (N_45,In_254,In_411);
nand U46 (N_46,In_697,In_319);
or U47 (N_47,In_730,In_615);
and U48 (N_48,In_724,In_576);
nand U49 (N_49,In_275,In_481);
nand U50 (N_50,In_105,In_701);
nor U51 (N_51,In_86,In_382);
nand U52 (N_52,In_160,In_335);
nor U53 (N_53,In_151,In_705);
nor U54 (N_54,In_73,In_363);
and U55 (N_55,In_453,In_278);
and U56 (N_56,In_2,In_504);
and U57 (N_57,In_584,In_713);
nand U58 (N_58,In_622,In_519);
or U59 (N_59,In_720,In_646);
nand U60 (N_60,In_311,In_285);
or U61 (N_61,In_321,In_192);
nor U62 (N_62,In_508,In_67);
nand U63 (N_63,In_568,In_213);
nand U64 (N_64,In_5,In_690);
or U65 (N_65,In_342,In_482);
and U66 (N_66,In_643,In_195);
and U67 (N_67,In_49,In_405);
or U68 (N_68,In_745,In_600);
nor U69 (N_69,In_164,In_604);
and U70 (N_70,In_221,In_381);
and U71 (N_71,In_79,In_345);
nor U72 (N_72,In_582,In_635);
and U73 (N_73,In_553,In_191);
and U74 (N_74,In_293,In_145);
nor U75 (N_75,In_474,In_383);
and U76 (N_76,In_549,In_18);
and U77 (N_77,In_638,In_364);
or U78 (N_78,In_336,In_348);
nand U79 (N_79,In_394,In_630);
or U80 (N_80,In_676,In_178);
nor U81 (N_81,In_562,In_44);
xor U82 (N_82,In_530,In_670);
and U83 (N_83,In_327,In_135);
nor U84 (N_84,In_499,In_429);
and U85 (N_85,In_406,In_108);
or U86 (N_86,In_666,In_288);
xor U87 (N_87,In_518,In_410);
and U88 (N_88,In_675,In_95);
nand U89 (N_89,In_212,In_637);
nand U90 (N_90,In_211,In_395);
nor U91 (N_91,In_522,In_148);
nand U92 (N_92,In_544,In_190);
nor U93 (N_93,In_287,In_346);
nor U94 (N_94,In_35,In_40);
xor U95 (N_95,In_99,In_592);
and U96 (N_96,In_274,In_477);
nand U97 (N_97,In_248,In_7);
xnor U98 (N_98,In_650,In_427);
nor U99 (N_99,In_263,In_238);
or U100 (N_100,In_422,In_401);
or U101 (N_101,In_132,In_542);
nor U102 (N_102,In_10,In_157);
xnor U103 (N_103,In_352,In_142);
or U104 (N_104,In_116,In_8);
and U105 (N_105,In_181,In_298);
xnor U106 (N_106,In_149,In_739);
and U107 (N_107,In_454,In_446);
and U108 (N_108,In_535,In_527);
nand U109 (N_109,In_236,In_659);
xnor U110 (N_110,In_579,In_305);
nand U111 (N_111,In_672,In_645);
nor U112 (N_112,In_272,In_585);
and U113 (N_113,In_391,In_165);
xor U114 (N_114,In_552,In_629);
nand U115 (N_115,In_75,In_486);
and U116 (N_116,In_299,In_94);
nor U117 (N_117,In_71,In_385);
nand U118 (N_118,In_639,In_53);
and U119 (N_119,In_452,In_667);
and U120 (N_120,In_710,In_728);
and U121 (N_121,In_738,In_618);
or U122 (N_122,In_525,In_545);
nor U123 (N_123,In_81,In_440);
xor U124 (N_124,In_114,In_359);
and U125 (N_125,In_137,In_344);
or U126 (N_126,In_356,In_580);
nand U127 (N_127,In_613,In_662);
nand U128 (N_128,In_177,In_156);
nor U129 (N_129,In_315,In_561);
and U130 (N_130,In_507,In_96);
nor U131 (N_131,In_362,In_223);
and U132 (N_132,In_612,In_436);
and U133 (N_133,In_426,In_1);
xor U134 (N_134,In_24,In_320);
nand U135 (N_135,In_403,In_412);
or U136 (N_136,In_459,In_494);
and U137 (N_137,In_413,In_677);
nand U138 (N_138,In_606,In_204);
nor U139 (N_139,In_379,In_265);
nor U140 (N_140,In_341,In_225);
and U141 (N_141,In_6,In_313);
and U142 (N_142,In_742,In_451);
or U143 (N_143,In_110,In_228);
or U144 (N_144,In_551,In_302);
xnor U145 (N_145,In_685,In_103);
or U146 (N_146,In_716,In_122);
or U147 (N_147,In_707,In_26);
nand U148 (N_148,In_303,In_371);
xor U149 (N_149,In_273,In_744);
nor U150 (N_150,In_21,In_611);
or U151 (N_151,In_597,In_497);
nand U152 (N_152,In_113,In_524);
and U153 (N_153,In_441,In_433);
nor U154 (N_154,In_169,In_227);
and U155 (N_155,In_370,In_106);
nand U156 (N_156,In_57,In_537);
nand U157 (N_157,In_698,In_457);
or U158 (N_158,In_632,In_139);
or U159 (N_159,In_176,In_610);
or U160 (N_160,In_397,In_90);
and U161 (N_161,In_554,In_608);
xnor U162 (N_162,In_708,In_340);
nand U163 (N_163,In_61,In_434);
and U164 (N_164,In_201,In_493);
nand U165 (N_165,In_571,In_572);
or U166 (N_166,In_30,In_239);
and U167 (N_167,In_418,In_172);
xor U168 (N_168,In_136,In_324);
or U169 (N_169,In_215,In_277);
or U170 (N_170,In_27,In_141);
or U171 (N_171,In_727,In_111);
and U172 (N_172,In_575,In_731);
or U173 (N_173,In_475,In_357);
or U174 (N_174,In_485,In_337);
and U175 (N_175,In_127,In_19);
nand U176 (N_176,In_644,In_722);
xnor U177 (N_177,In_207,In_331);
or U178 (N_178,In_693,In_58);
xnor U179 (N_179,In_361,In_39);
nor U180 (N_180,In_529,In_69);
nor U181 (N_181,In_267,In_619);
nor U182 (N_182,In_489,In_55);
nand U183 (N_183,In_316,In_651);
or U184 (N_184,In_398,In_387);
nand U185 (N_185,In_621,In_392);
nor U186 (N_186,In_668,In_588);
nor U187 (N_187,In_161,In_669);
xnor U188 (N_188,In_741,In_573);
or U189 (N_189,In_29,In_251);
nor U190 (N_190,In_87,In_557);
nor U191 (N_191,In_182,In_488);
or U192 (N_192,In_423,In_230);
nor U193 (N_193,In_642,In_664);
xnor U194 (N_194,In_513,In_22);
nor U195 (N_195,In_460,In_435);
nand U196 (N_196,In_32,In_246);
nor U197 (N_197,In_439,In_147);
or U198 (N_198,In_472,In_536);
or U199 (N_199,In_46,In_193);
and U200 (N_200,In_15,In_31);
nor U201 (N_201,In_14,In_384);
nand U202 (N_202,In_23,In_280);
nor U203 (N_203,In_591,In_541);
nand U204 (N_204,In_308,In_289);
nand U205 (N_205,In_445,In_129);
or U206 (N_206,In_13,In_569);
or U207 (N_207,In_749,In_623);
nor U208 (N_208,In_737,In_520);
or U209 (N_209,In_678,In_48);
or U210 (N_210,In_186,In_417);
nor U211 (N_211,In_175,In_478);
xnor U212 (N_212,In_249,In_242);
and U213 (N_213,In_307,In_634);
and U214 (N_214,In_539,In_640);
or U215 (N_215,In_358,In_574);
nand U216 (N_216,In_159,In_495);
xor U217 (N_217,In_244,In_268);
or U218 (N_218,In_146,In_54);
xor U219 (N_219,In_449,In_656);
nor U220 (N_220,In_301,In_692);
nor U221 (N_221,In_256,In_390);
nand U222 (N_222,In_375,In_466);
and U223 (N_223,In_470,In_206);
or U224 (N_224,In_347,In_514);
and U225 (N_225,In_155,In_284);
and U226 (N_226,In_264,In_154);
xnor U227 (N_227,In_88,In_310);
nand U228 (N_228,In_605,In_684);
or U229 (N_229,In_628,In_100);
nand U230 (N_230,In_715,In_282);
and U231 (N_231,In_616,In_408);
xnor U232 (N_232,In_665,In_92);
nand U233 (N_233,In_131,In_78);
and U234 (N_234,In_197,In_72);
nor U235 (N_235,In_218,In_484);
or U236 (N_236,In_210,In_222);
and U237 (N_237,In_566,In_424);
nand U238 (N_238,In_295,In_480);
nand U239 (N_239,In_546,In_245);
nand U240 (N_240,In_442,In_174);
xor U241 (N_241,In_603,In_686);
xor U242 (N_242,In_373,In_85);
nand U243 (N_243,In_704,In_202);
or U244 (N_244,In_702,In_648);
nand U245 (N_245,In_502,In_60);
nor U246 (N_246,In_25,In_89);
nor U247 (N_247,In_388,In_104);
nor U248 (N_248,In_107,In_240);
nand U249 (N_249,In_409,In_333);
or U250 (N_250,In_77,In_609);
nor U251 (N_251,In_570,In_641);
nand U252 (N_252,In_501,In_593);
and U253 (N_253,In_718,In_404);
nand U254 (N_254,In_377,In_595);
nand U255 (N_255,In_183,In_200);
xnor U256 (N_256,In_421,In_270);
nor U257 (N_257,In_456,In_214);
or U258 (N_258,In_602,In_332);
or U259 (N_259,In_63,In_703);
nor U260 (N_260,In_45,In_589);
or U261 (N_261,In_283,In_695);
nand U262 (N_262,In_721,In_746);
or U263 (N_263,In_126,In_80);
xor U264 (N_264,In_260,In_0);
nand U265 (N_265,In_323,In_16);
nand U266 (N_266,In_652,In_443);
nand U267 (N_267,In_607,In_736);
or U268 (N_268,In_556,In_476);
nand U269 (N_269,In_134,In_209);
or U270 (N_270,In_59,In_687);
and U271 (N_271,In_170,In_414);
or U272 (N_272,In_252,In_97);
nor U273 (N_273,In_243,In_747);
nand U274 (N_274,In_372,In_98);
nor U275 (N_275,In_34,In_688);
nand U276 (N_276,In_124,In_50);
or U277 (N_277,In_487,In_91);
and U278 (N_278,In_425,In_300);
nand U279 (N_279,In_444,In_516);
xnor U280 (N_280,In_732,In_671);
and U281 (N_281,In_694,In_220);
nor U282 (N_282,In_625,In_735);
nor U283 (N_283,In_343,In_399);
or U284 (N_284,In_555,In_179);
and U285 (N_285,In_121,In_168);
nor U286 (N_286,In_119,In_355);
nor U287 (N_287,In_455,In_226);
xor U288 (N_288,In_437,In_419);
nor U289 (N_289,In_550,In_534);
nor U290 (N_290,In_503,In_130);
nand U291 (N_291,In_725,In_458);
xor U292 (N_292,In_9,In_723);
nor U293 (N_293,In_339,In_491);
or U294 (N_294,In_402,In_184);
nor U295 (N_295,In_509,In_185);
and U296 (N_296,In_140,In_450);
and U297 (N_297,In_586,In_448);
xor U298 (N_298,In_328,In_281);
nand U299 (N_299,In_748,In_740);
nor U300 (N_300,In_462,In_37);
nand U301 (N_301,In_432,In_125);
or U302 (N_302,In_564,In_682);
or U303 (N_303,In_567,In_691);
nor U304 (N_304,In_661,In_120);
and U305 (N_305,In_3,In_187);
nor U306 (N_306,In_492,In_559);
nor U307 (N_307,In_173,In_366);
or U308 (N_308,In_681,In_389);
nor U309 (N_309,In_309,In_144);
nor U310 (N_310,In_490,In_93);
nand U311 (N_311,In_647,In_523);
xor U312 (N_312,In_368,In_224);
nor U313 (N_313,In_367,In_653);
xnor U314 (N_314,In_250,In_601);
or U315 (N_315,In_262,In_374);
and U316 (N_316,In_416,In_696);
xor U317 (N_317,In_547,In_683);
or U318 (N_318,In_376,In_614);
and U319 (N_319,In_205,In_306);
and U320 (N_320,In_163,In_286);
nor U321 (N_321,In_259,In_633);
nand U322 (N_322,In_150,In_624);
nor U323 (N_323,In_654,In_68);
nor U324 (N_324,In_318,In_158);
or U325 (N_325,In_521,In_469);
nor U326 (N_326,In_74,In_330);
nor U327 (N_327,In_468,In_117);
and U328 (N_328,In_271,In_565);
nand U329 (N_329,In_717,In_711);
nand U330 (N_330,In_138,In_338);
nor U331 (N_331,In_84,In_233);
or U332 (N_332,In_447,In_234);
nor U333 (N_333,In_596,In_217);
nor U334 (N_334,In_101,In_461);
and U335 (N_335,In_208,In_229);
nand U336 (N_336,In_203,In_673);
nor U337 (N_337,In_82,In_350);
nand U338 (N_338,In_198,In_253);
nand U339 (N_339,In_153,In_353);
nand U340 (N_340,In_506,In_62);
nor U341 (N_341,In_471,In_199);
nand U342 (N_342,In_162,In_312);
nand U343 (N_343,In_473,In_247);
and U344 (N_344,In_386,In_510);
nor U345 (N_345,In_65,In_689);
or U346 (N_346,In_304,In_563);
or U347 (N_347,In_407,In_351);
nand U348 (N_348,In_257,In_626);
nor U349 (N_349,In_540,In_41);
and U350 (N_350,In_396,In_109);
nor U351 (N_351,In_658,In_133);
nor U352 (N_352,In_496,In_543);
nor U353 (N_353,In_438,In_266);
nor U354 (N_354,In_297,In_590);
nor U355 (N_355,In_290,In_276);
and U356 (N_356,In_431,In_171);
and U357 (N_357,In_729,In_291);
xor U358 (N_358,In_532,In_393);
xnor U359 (N_359,In_261,In_558);
or U360 (N_360,In_36,In_66);
and U361 (N_361,In_463,In_42);
xor U362 (N_362,In_598,In_733);
and U363 (N_363,In_326,In_83);
nor U364 (N_364,In_296,In_712);
or U365 (N_365,In_577,In_680);
and U366 (N_366,In_587,In_167);
nor U367 (N_367,In_196,In_241);
or U368 (N_368,In_322,In_415);
nor U369 (N_369,In_12,In_20);
nor U370 (N_370,In_232,In_325);
xor U371 (N_371,In_365,In_369);
nand U372 (N_372,In_380,In_231);
xnor U373 (N_373,In_51,In_548);
and U374 (N_374,In_64,In_464);
or U375 (N_375,In_434,In_690);
nand U376 (N_376,In_505,In_422);
and U377 (N_377,In_116,In_61);
or U378 (N_378,In_465,In_628);
nor U379 (N_379,In_614,In_281);
nand U380 (N_380,In_477,In_247);
nor U381 (N_381,In_204,In_565);
nand U382 (N_382,In_479,In_368);
and U383 (N_383,In_544,In_608);
or U384 (N_384,In_130,In_381);
or U385 (N_385,In_486,In_544);
xnor U386 (N_386,In_501,In_591);
or U387 (N_387,In_104,In_684);
and U388 (N_388,In_336,In_573);
nor U389 (N_389,In_384,In_193);
and U390 (N_390,In_32,In_83);
and U391 (N_391,In_516,In_512);
nand U392 (N_392,In_417,In_212);
and U393 (N_393,In_296,In_710);
nand U394 (N_394,In_178,In_632);
or U395 (N_395,In_388,In_73);
or U396 (N_396,In_382,In_77);
and U397 (N_397,In_264,In_540);
and U398 (N_398,In_671,In_455);
and U399 (N_399,In_624,In_300);
nand U400 (N_400,In_104,In_616);
nor U401 (N_401,In_513,In_492);
nor U402 (N_402,In_454,In_210);
xor U403 (N_403,In_380,In_275);
and U404 (N_404,In_518,In_644);
nor U405 (N_405,In_136,In_720);
nor U406 (N_406,In_619,In_563);
nor U407 (N_407,In_76,In_5);
and U408 (N_408,In_51,In_464);
nor U409 (N_409,In_744,In_60);
and U410 (N_410,In_725,In_397);
or U411 (N_411,In_275,In_161);
or U412 (N_412,In_421,In_658);
nand U413 (N_413,In_434,In_335);
nor U414 (N_414,In_208,In_273);
nand U415 (N_415,In_477,In_691);
nor U416 (N_416,In_632,In_291);
nor U417 (N_417,In_355,In_542);
or U418 (N_418,In_444,In_437);
or U419 (N_419,In_162,In_369);
nand U420 (N_420,In_405,In_684);
nor U421 (N_421,In_304,In_148);
nand U422 (N_422,In_230,In_35);
nor U423 (N_423,In_283,In_408);
or U424 (N_424,In_549,In_411);
nand U425 (N_425,In_522,In_84);
nor U426 (N_426,In_500,In_378);
and U427 (N_427,In_73,In_234);
or U428 (N_428,In_673,In_400);
nor U429 (N_429,In_399,In_735);
nor U430 (N_430,In_635,In_462);
and U431 (N_431,In_672,In_77);
or U432 (N_432,In_528,In_710);
nor U433 (N_433,In_411,In_293);
and U434 (N_434,In_274,In_659);
and U435 (N_435,In_734,In_2);
nor U436 (N_436,In_64,In_380);
nand U437 (N_437,In_612,In_247);
nor U438 (N_438,In_466,In_209);
nand U439 (N_439,In_199,In_314);
nand U440 (N_440,In_228,In_80);
or U441 (N_441,In_15,In_392);
nand U442 (N_442,In_53,In_20);
nand U443 (N_443,In_161,In_425);
nor U444 (N_444,In_598,In_692);
nand U445 (N_445,In_332,In_489);
xor U446 (N_446,In_361,In_669);
or U447 (N_447,In_89,In_37);
nand U448 (N_448,In_404,In_505);
nand U449 (N_449,In_605,In_202);
xor U450 (N_450,In_236,In_610);
or U451 (N_451,In_143,In_52);
or U452 (N_452,In_156,In_325);
and U453 (N_453,In_347,In_548);
nor U454 (N_454,In_533,In_448);
nand U455 (N_455,In_570,In_393);
xnor U456 (N_456,In_344,In_99);
and U457 (N_457,In_120,In_652);
nand U458 (N_458,In_451,In_14);
nor U459 (N_459,In_506,In_354);
or U460 (N_460,In_700,In_315);
or U461 (N_461,In_449,In_362);
nor U462 (N_462,In_23,In_183);
nor U463 (N_463,In_348,In_411);
and U464 (N_464,In_323,In_195);
xor U465 (N_465,In_173,In_343);
nand U466 (N_466,In_394,In_725);
nor U467 (N_467,In_222,In_625);
nor U468 (N_468,In_699,In_372);
xnor U469 (N_469,In_82,In_253);
nor U470 (N_470,In_396,In_337);
nand U471 (N_471,In_112,In_340);
nand U472 (N_472,In_439,In_31);
nor U473 (N_473,In_396,In_214);
nand U474 (N_474,In_273,In_17);
nor U475 (N_475,In_24,In_349);
or U476 (N_476,In_719,In_476);
nand U477 (N_477,In_347,In_521);
and U478 (N_478,In_90,In_254);
and U479 (N_479,In_713,In_741);
and U480 (N_480,In_238,In_23);
and U481 (N_481,In_123,In_154);
nand U482 (N_482,In_574,In_334);
or U483 (N_483,In_109,In_355);
nand U484 (N_484,In_196,In_438);
or U485 (N_485,In_139,In_616);
or U486 (N_486,In_513,In_132);
and U487 (N_487,In_281,In_726);
xor U488 (N_488,In_515,In_17);
xor U489 (N_489,In_492,In_226);
or U490 (N_490,In_174,In_479);
nor U491 (N_491,In_2,In_253);
or U492 (N_492,In_585,In_492);
nor U493 (N_493,In_315,In_81);
nor U494 (N_494,In_746,In_549);
nand U495 (N_495,In_38,In_681);
nand U496 (N_496,In_291,In_491);
or U497 (N_497,In_43,In_236);
and U498 (N_498,In_282,In_157);
and U499 (N_499,In_307,In_428);
or U500 (N_500,In_465,In_561);
nand U501 (N_501,In_105,In_365);
and U502 (N_502,In_415,In_673);
nand U503 (N_503,In_598,In_110);
nor U504 (N_504,In_286,In_588);
xor U505 (N_505,In_606,In_217);
or U506 (N_506,In_187,In_724);
nand U507 (N_507,In_76,In_492);
and U508 (N_508,In_620,In_657);
nor U509 (N_509,In_586,In_723);
and U510 (N_510,In_387,In_600);
and U511 (N_511,In_87,In_649);
nor U512 (N_512,In_740,In_29);
nand U513 (N_513,In_638,In_174);
nand U514 (N_514,In_64,In_113);
nand U515 (N_515,In_29,In_7);
xor U516 (N_516,In_372,In_486);
and U517 (N_517,In_639,In_551);
and U518 (N_518,In_705,In_139);
and U519 (N_519,In_345,In_360);
xnor U520 (N_520,In_16,In_190);
and U521 (N_521,In_179,In_682);
or U522 (N_522,In_675,In_361);
nand U523 (N_523,In_384,In_23);
and U524 (N_524,In_291,In_23);
or U525 (N_525,In_48,In_271);
nor U526 (N_526,In_650,In_572);
and U527 (N_527,In_432,In_255);
nand U528 (N_528,In_461,In_98);
and U529 (N_529,In_72,In_647);
nor U530 (N_530,In_724,In_206);
nand U531 (N_531,In_660,In_222);
and U532 (N_532,In_557,In_0);
nand U533 (N_533,In_303,In_32);
nand U534 (N_534,In_339,In_632);
and U535 (N_535,In_30,In_349);
or U536 (N_536,In_259,In_64);
nor U537 (N_537,In_87,In_456);
nor U538 (N_538,In_475,In_252);
or U539 (N_539,In_362,In_580);
and U540 (N_540,In_267,In_249);
nor U541 (N_541,In_519,In_639);
and U542 (N_542,In_20,In_36);
and U543 (N_543,In_672,In_163);
nand U544 (N_544,In_170,In_556);
or U545 (N_545,In_223,In_680);
nand U546 (N_546,In_300,In_110);
nand U547 (N_547,In_17,In_31);
xor U548 (N_548,In_241,In_585);
nand U549 (N_549,In_743,In_441);
nand U550 (N_550,In_655,In_468);
or U551 (N_551,In_437,In_251);
nor U552 (N_552,In_647,In_236);
nand U553 (N_553,In_20,In_481);
nand U554 (N_554,In_723,In_23);
and U555 (N_555,In_623,In_615);
and U556 (N_556,In_638,In_501);
nand U557 (N_557,In_172,In_440);
and U558 (N_558,In_403,In_342);
nor U559 (N_559,In_326,In_629);
and U560 (N_560,In_747,In_198);
nand U561 (N_561,In_226,In_354);
nor U562 (N_562,In_220,In_594);
or U563 (N_563,In_251,In_676);
or U564 (N_564,In_42,In_322);
xnor U565 (N_565,In_493,In_645);
nand U566 (N_566,In_258,In_501);
or U567 (N_567,In_742,In_672);
and U568 (N_568,In_136,In_5);
and U569 (N_569,In_586,In_259);
or U570 (N_570,In_197,In_591);
nand U571 (N_571,In_697,In_379);
or U572 (N_572,In_527,In_653);
nor U573 (N_573,In_627,In_226);
nand U574 (N_574,In_263,In_413);
nor U575 (N_575,In_99,In_470);
nand U576 (N_576,In_120,In_617);
and U577 (N_577,In_85,In_42);
and U578 (N_578,In_248,In_149);
xor U579 (N_579,In_678,In_394);
and U580 (N_580,In_39,In_30);
xnor U581 (N_581,In_544,In_26);
nor U582 (N_582,In_389,In_517);
nand U583 (N_583,In_106,In_609);
nand U584 (N_584,In_420,In_423);
or U585 (N_585,In_478,In_309);
and U586 (N_586,In_283,In_199);
nor U587 (N_587,In_695,In_330);
nand U588 (N_588,In_488,In_651);
and U589 (N_589,In_18,In_288);
xnor U590 (N_590,In_51,In_373);
xnor U591 (N_591,In_117,In_273);
nand U592 (N_592,In_577,In_447);
or U593 (N_593,In_610,In_66);
nor U594 (N_594,In_733,In_640);
nor U595 (N_595,In_325,In_294);
and U596 (N_596,In_58,In_636);
and U597 (N_597,In_343,In_415);
nor U598 (N_598,In_448,In_428);
nand U599 (N_599,In_591,In_200);
nand U600 (N_600,In_126,In_521);
and U601 (N_601,In_311,In_312);
nand U602 (N_602,In_679,In_555);
or U603 (N_603,In_711,In_521);
or U604 (N_604,In_638,In_460);
or U605 (N_605,In_277,In_30);
and U606 (N_606,In_374,In_740);
and U607 (N_607,In_632,In_738);
and U608 (N_608,In_720,In_450);
and U609 (N_609,In_728,In_738);
nor U610 (N_610,In_545,In_329);
nand U611 (N_611,In_688,In_124);
or U612 (N_612,In_690,In_47);
nand U613 (N_613,In_356,In_211);
nor U614 (N_614,In_411,In_553);
nor U615 (N_615,In_454,In_148);
or U616 (N_616,In_397,In_137);
nor U617 (N_617,In_239,In_522);
xor U618 (N_618,In_76,In_284);
or U619 (N_619,In_53,In_549);
nand U620 (N_620,In_394,In_646);
nand U621 (N_621,In_642,In_101);
and U622 (N_622,In_602,In_408);
nor U623 (N_623,In_192,In_95);
nor U624 (N_624,In_88,In_747);
or U625 (N_625,In_690,In_400);
and U626 (N_626,In_441,In_364);
or U627 (N_627,In_272,In_237);
nand U628 (N_628,In_214,In_350);
or U629 (N_629,In_22,In_131);
and U630 (N_630,In_436,In_382);
nor U631 (N_631,In_158,In_387);
nand U632 (N_632,In_105,In_632);
nor U633 (N_633,In_218,In_742);
nand U634 (N_634,In_6,In_487);
and U635 (N_635,In_43,In_661);
nand U636 (N_636,In_319,In_77);
and U637 (N_637,In_517,In_233);
or U638 (N_638,In_590,In_732);
or U639 (N_639,In_620,In_33);
nor U640 (N_640,In_330,In_420);
nand U641 (N_641,In_394,In_346);
or U642 (N_642,In_114,In_132);
nor U643 (N_643,In_52,In_479);
nor U644 (N_644,In_598,In_153);
and U645 (N_645,In_436,In_670);
and U646 (N_646,In_688,In_48);
nor U647 (N_647,In_482,In_530);
and U648 (N_648,In_708,In_237);
and U649 (N_649,In_720,In_449);
or U650 (N_650,In_460,In_360);
or U651 (N_651,In_437,In_712);
or U652 (N_652,In_400,In_397);
or U653 (N_653,In_471,In_366);
nor U654 (N_654,In_245,In_699);
nand U655 (N_655,In_344,In_287);
or U656 (N_656,In_84,In_588);
nor U657 (N_657,In_375,In_663);
and U658 (N_658,In_108,In_156);
nand U659 (N_659,In_69,In_423);
nand U660 (N_660,In_451,In_664);
and U661 (N_661,In_16,In_304);
nand U662 (N_662,In_85,In_222);
nor U663 (N_663,In_328,In_491);
nand U664 (N_664,In_219,In_205);
or U665 (N_665,In_554,In_319);
nor U666 (N_666,In_95,In_540);
or U667 (N_667,In_368,In_713);
nor U668 (N_668,In_521,In_713);
or U669 (N_669,In_265,In_351);
and U670 (N_670,In_138,In_449);
and U671 (N_671,In_172,In_193);
nor U672 (N_672,In_171,In_653);
nor U673 (N_673,In_532,In_705);
xor U674 (N_674,In_312,In_264);
nor U675 (N_675,In_575,In_190);
or U676 (N_676,In_556,In_372);
or U677 (N_677,In_226,In_186);
or U678 (N_678,In_98,In_690);
and U679 (N_679,In_21,In_251);
xor U680 (N_680,In_722,In_287);
nor U681 (N_681,In_615,In_739);
nand U682 (N_682,In_154,In_107);
nand U683 (N_683,In_424,In_592);
nor U684 (N_684,In_715,In_177);
nand U685 (N_685,In_694,In_412);
or U686 (N_686,In_260,In_579);
or U687 (N_687,In_253,In_737);
nor U688 (N_688,In_586,In_237);
or U689 (N_689,In_648,In_584);
or U690 (N_690,In_693,In_241);
and U691 (N_691,In_735,In_192);
nand U692 (N_692,In_553,In_175);
and U693 (N_693,In_517,In_423);
nor U694 (N_694,In_721,In_189);
or U695 (N_695,In_587,In_90);
nor U696 (N_696,In_430,In_628);
nand U697 (N_697,In_485,In_66);
or U698 (N_698,In_112,In_633);
nand U699 (N_699,In_27,In_29);
nor U700 (N_700,In_606,In_682);
xnor U701 (N_701,In_291,In_667);
nand U702 (N_702,In_258,In_35);
nor U703 (N_703,In_75,In_251);
and U704 (N_704,In_132,In_320);
nor U705 (N_705,In_413,In_198);
and U706 (N_706,In_433,In_673);
xor U707 (N_707,In_519,In_596);
and U708 (N_708,In_512,In_181);
xnor U709 (N_709,In_268,In_482);
nand U710 (N_710,In_190,In_271);
and U711 (N_711,In_271,In_60);
nor U712 (N_712,In_548,In_74);
nand U713 (N_713,In_638,In_59);
and U714 (N_714,In_524,In_396);
nor U715 (N_715,In_293,In_34);
and U716 (N_716,In_183,In_110);
and U717 (N_717,In_580,In_651);
xnor U718 (N_718,In_120,In_418);
nand U719 (N_719,In_443,In_205);
or U720 (N_720,In_154,In_658);
nor U721 (N_721,In_588,In_407);
or U722 (N_722,In_534,In_479);
nor U723 (N_723,In_293,In_15);
nor U724 (N_724,In_635,In_90);
and U725 (N_725,In_498,In_743);
and U726 (N_726,In_421,In_2);
nand U727 (N_727,In_299,In_682);
or U728 (N_728,In_712,In_86);
or U729 (N_729,In_326,In_571);
xor U730 (N_730,In_250,In_194);
or U731 (N_731,In_155,In_551);
and U732 (N_732,In_552,In_275);
xnor U733 (N_733,In_529,In_430);
nor U734 (N_734,In_47,In_98);
and U735 (N_735,In_535,In_730);
xnor U736 (N_736,In_339,In_478);
or U737 (N_737,In_515,In_368);
nor U738 (N_738,In_303,In_596);
xor U739 (N_739,In_710,In_698);
nor U740 (N_740,In_259,In_504);
nor U741 (N_741,In_278,In_479);
and U742 (N_742,In_223,In_22);
or U743 (N_743,In_70,In_225);
and U744 (N_744,In_498,In_258);
nor U745 (N_745,In_708,In_262);
nor U746 (N_746,In_646,In_247);
nand U747 (N_747,In_234,In_486);
xor U748 (N_748,In_703,In_79);
or U749 (N_749,In_507,In_440);
nand U750 (N_750,In_172,In_146);
nand U751 (N_751,In_591,In_128);
nand U752 (N_752,In_215,In_406);
and U753 (N_753,In_41,In_584);
nor U754 (N_754,In_472,In_513);
xor U755 (N_755,In_604,In_60);
xor U756 (N_756,In_85,In_401);
and U757 (N_757,In_105,In_164);
and U758 (N_758,In_190,In_492);
nand U759 (N_759,In_580,In_435);
or U760 (N_760,In_481,In_570);
nand U761 (N_761,In_157,In_306);
nor U762 (N_762,In_733,In_340);
nand U763 (N_763,In_126,In_594);
or U764 (N_764,In_672,In_652);
or U765 (N_765,In_598,In_534);
nand U766 (N_766,In_370,In_403);
nor U767 (N_767,In_335,In_166);
nand U768 (N_768,In_312,In_383);
and U769 (N_769,In_572,In_539);
nand U770 (N_770,In_501,In_618);
nor U771 (N_771,In_306,In_317);
nor U772 (N_772,In_402,In_713);
nand U773 (N_773,In_257,In_589);
nand U774 (N_774,In_654,In_299);
or U775 (N_775,In_603,In_241);
nor U776 (N_776,In_155,In_294);
xnor U777 (N_777,In_635,In_205);
xnor U778 (N_778,In_447,In_362);
and U779 (N_779,In_180,In_233);
and U780 (N_780,In_214,In_199);
or U781 (N_781,In_273,In_582);
or U782 (N_782,In_341,In_327);
or U783 (N_783,In_243,In_56);
or U784 (N_784,In_82,In_216);
and U785 (N_785,In_177,In_674);
and U786 (N_786,In_137,In_18);
or U787 (N_787,In_594,In_294);
and U788 (N_788,In_440,In_117);
nor U789 (N_789,In_45,In_378);
nor U790 (N_790,In_637,In_260);
and U791 (N_791,In_413,In_565);
and U792 (N_792,In_120,In_614);
nor U793 (N_793,In_488,In_372);
nor U794 (N_794,In_103,In_47);
nor U795 (N_795,In_271,In_53);
nand U796 (N_796,In_530,In_214);
and U797 (N_797,In_597,In_61);
and U798 (N_798,In_126,In_568);
and U799 (N_799,In_489,In_187);
nor U800 (N_800,In_505,In_11);
and U801 (N_801,In_136,In_634);
and U802 (N_802,In_489,In_230);
nand U803 (N_803,In_72,In_437);
and U804 (N_804,In_380,In_183);
xnor U805 (N_805,In_63,In_402);
nor U806 (N_806,In_36,In_420);
nand U807 (N_807,In_213,In_623);
xor U808 (N_808,In_561,In_413);
and U809 (N_809,In_554,In_547);
nor U810 (N_810,In_603,In_555);
nand U811 (N_811,In_679,In_117);
xnor U812 (N_812,In_494,In_323);
and U813 (N_813,In_131,In_303);
nand U814 (N_814,In_708,In_166);
nand U815 (N_815,In_642,In_256);
or U816 (N_816,In_696,In_357);
nor U817 (N_817,In_396,In_403);
nor U818 (N_818,In_311,In_711);
or U819 (N_819,In_292,In_266);
nand U820 (N_820,In_71,In_118);
and U821 (N_821,In_391,In_659);
nand U822 (N_822,In_342,In_373);
and U823 (N_823,In_74,In_607);
nand U824 (N_824,In_718,In_18);
nor U825 (N_825,In_191,In_205);
xnor U826 (N_826,In_665,In_636);
or U827 (N_827,In_404,In_152);
nand U828 (N_828,In_309,In_374);
nand U829 (N_829,In_214,In_358);
or U830 (N_830,In_62,In_345);
nor U831 (N_831,In_353,In_390);
and U832 (N_832,In_218,In_640);
nor U833 (N_833,In_281,In_745);
or U834 (N_834,In_543,In_577);
nor U835 (N_835,In_630,In_716);
nand U836 (N_836,In_31,In_392);
or U837 (N_837,In_177,In_262);
and U838 (N_838,In_535,In_713);
and U839 (N_839,In_161,In_744);
and U840 (N_840,In_619,In_213);
nor U841 (N_841,In_337,In_451);
nor U842 (N_842,In_514,In_177);
xnor U843 (N_843,In_683,In_127);
nand U844 (N_844,In_441,In_279);
nand U845 (N_845,In_283,In_551);
nor U846 (N_846,In_248,In_258);
or U847 (N_847,In_189,In_381);
and U848 (N_848,In_706,In_491);
and U849 (N_849,In_204,In_691);
or U850 (N_850,In_706,In_552);
or U851 (N_851,In_385,In_451);
xor U852 (N_852,In_66,In_666);
or U853 (N_853,In_698,In_51);
xnor U854 (N_854,In_629,In_626);
or U855 (N_855,In_533,In_699);
nor U856 (N_856,In_481,In_528);
nand U857 (N_857,In_130,In_319);
or U858 (N_858,In_409,In_706);
xor U859 (N_859,In_631,In_621);
nand U860 (N_860,In_452,In_511);
and U861 (N_861,In_111,In_518);
nand U862 (N_862,In_470,In_605);
nor U863 (N_863,In_677,In_373);
and U864 (N_864,In_19,In_524);
or U865 (N_865,In_396,In_746);
or U866 (N_866,In_46,In_161);
nor U867 (N_867,In_382,In_611);
nand U868 (N_868,In_15,In_524);
or U869 (N_869,In_270,In_317);
nor U870 (N_870,In_683,In_174);
nor U871 (N_871,In_210,In_624);
nand U872 (N_872,In_394,In_187);
nand U873 (N_873,In_46,In_97);
nor U874 (N_874,In_544,In_457);
nor U875 (N_875,In_513,In_158);
and U876 (N_876,In_404,In_160);
or U877 (N_877,In_538,In_503);
and U878 (N_878,In_566,In_723);
nor U879 (N_879,In_402,In_223);
nand U880 (N_880,In_426,In_447);
or U881 (N_881,In_257,In_31);
nand U882 (N_882,In_91,In_575);
nand U883 (N_883,In_647,In_16);
nand U884 (N_884,In_664,In_26);
and U885 (N_885,In_674,In_446);
nor U886 (N_886,In_105,In_600);
and U887 (N_887,In_559,In_474);
nand U888 (N_888,In_597,In_332);
nor U889 (N_889,In_718,In_197);
xor U890 (N_890,In_546,In_378);
nand U891 (N_891,In_590,In_231);
nand U892 (N_892,In_475,In_317);
nand U893 (N_893,In_66,In_213);
xor U894 (N_894,In_406,In_620);
nand U895 (N_895,In_514,In_135);
and U896 (N_896,In_581,In_693);
nor U897 (N_897,In_202,In_170);
and U898 (N_898,In_216,In_289);
xor U899 (N_899,In_602,In_393);
nand U900 (N_900,In_609,In_514);
nand U901 (N_901,In_253,In_566);
nor U902 (N_902,In_625,In_20);
nor U903 (N_903,In_607,In_575);
nor U904 (N_904,In_100,In_90);
nor U905 (N_905,In_319,In_210);
and U906 (N_906,In_397,In_232);
xor U907 (N_907,In_564,In_436);
nor U908 (N_908,In_269,In_522);
and U909 (N_909,In_89,In_638);
nand U910 (N_910,In_651,In_177);
nor U911 (N_911,In_509,In_491);
and U912 (N_912,In_519,In_142);
nand U913 (N_913,In_105,In_78);
or U914 (N_914,In_404,In_745);
nor U915 (N_915,In_732,In_578);
or U916 (N_916,In_524,In_711);
nand U917 (N_917,In_722,In_468);
and U918 (N_918,In_408,In_653);
xor U919 (N_919,In_738,In_283);
and U920 (N_920,In_646,In_342);
and U921 (N_921,In_511,In_682);
xnor U922 (N_922,In_742,In_375);
nor U923 (N_923,In_571,In_212);
nor U924 (N_924,In_662,In_180);
nor U925 (N_925,In_205,In_197);
xnor U926 (N_926,In_62,In_358);
or U927 (N_927,In_599,In_413);
nand U928 (N_928,In_292,In_319);
or U929 (N_929,In_640,In_288);
xnor U930 (N_930,In_625,In_706);
nand U931 (N_931,In_209,In_470);
nor U932 (N_932,In_655,In_431);
or U933 (N_933,In_251,In_17);
nor U934 (N_934,In_584,In_121);
nand U935 (N_935,In_609,In_331);
nor U936 (N_936,In_111,In_249);
or U937 (N_937,In_448,In_192);
or U938 (N_938,In_551,In_53);
xnor U939 (N_939,In_460,In_554);
or U940 (N_940,In_205,In_254);
nor U941 (N_941,In_115,In_594);
nor U942 (N_942,In_78,In_529);
and U943 (N_943,In_190,In_498);
xor U944 (N_944,In_354,In_475);
nor U945 (N_945,In_413,In_325);
nand U946 (N_946,In_176,In_734);
nor U947 (N_947,In_425,In_401);
or U948 (N_948,In_549,In_404);
xor U949 (N_949,In_525,In_544);
nor U950 (N_950,In_603,In_180);
or U951 (N_951,In_158,In_704);
and U952 (N_952,In_176,In_458);
xnor U953 (N_953,In_671,In_58);
or U954 (N_954,In_548,In_563);
xor U955 (N_955,In_666,In_620);
or U956 (N_956,In_568,In_30);
nand U957 (N_957,In_150,In_52);
or U958 (N_958,In_308,In_56);
nand U959 (N_959,In_326,In_546);
and U960 (N_960,In_669,In_431);
nor U961 (N_961,In_601,In_48);
nor U962 (N_962,In_130,In_703);
and U963 (N_963,In_747,In_586);
nor U964 (N_964,In_283,In_214);
and U965 (N_965,In_668,In_503);
nand U966 (N_966,In_430,In_133);
nor U967 (N_967,In_292,In_379);
nor U968 (N_968,In_332,In_278);
or U969 (N_969,In_148,In_333);
and U970 (N_970,In_514,In_491);
or U971 (N_971,In_634,In_686);
nand U972 (N_972,In_138,In_109);
and U973 (N_973,In_642,In_538);
nand U974 (N_974,In_717,In_364);
or U975 (N_975,In_527,In_645);
nor U976 (N_976,In_749,In_251);
nor U977 (N_977,In_425,In_60);
nand U978 (N_978,In_631,In_574);
or U979 (N_979,In_445,In_575);
or U980 (N_980,In_330,In_749);
or U981 (N_981,In_570,In_150);
nand U982 (N_982,In_115,In_333);
nand U983 (N_983,In_551,In_474);
nand U984 (N_984,In_170,In_18);
xnor U985 (N_985,In_543,In_719);
nand U986 (N_986,In_427,In_217);
nor U987 (N_987,In_173,In_719);
nor U988 (N_988,In_361,In_140);
and U989 (N_989,In_88,In_366);
and U990 (N_990,In_684,In_588);
and U991 (N_991,In_740,In_438);
or U992 (N_992,In_568,In_375);
xor U993 (N_993,In_528,In_24);
xor U994 (N_994,In_560,In_170);
or U995 (N_995,In_442,In_492);
nand U996 (N_996,In_664,In_497);
or U997 (N_997,In_105,In_426);
and U998 (N_998,In_518,In_376);
nand U999 (N_999,In_454,In_449);
nand U1000 (N_1000,N_890,N_284);
or U1001 (N_1001,N_838,N_738);
nor U1002 (N_1002,N_474,N_742);
nor U1003 (N_1003,N_987,N_143);
xnor U1004 (N_1004,N_723,N_264);
and U1005 (N_1005,N_487,N_872);
or U1006 (N_1006,N_33,N_856);
nand U1007 (N_1007,N_857,N_840);
nor U1008 (N_1008,N_712,N_548);
nor U1009 (N_1009,N_137,N_417);
or U1010 (N_1010,N_708,N_959);
nand U1011 (N_1011,N_256,N_821);
nand U1012 (N_1012,N_610,N_300);
xor U1013 (N_1013,N_608,N_989);
and U1014 (N_1014,N_414,N_392);
and U1015 (N_1015,N_914,N_584);
nor U1016 (N_1016,N_615,N_134);
or U1017 (N_1017,N_818,N_289);
nor U1018 (N_1018,N_244,N_568);
or U1019 (N_1019,N_450,N_728);
and U1020 (N_1020,N_697,N_198);
nor U1021 (N_1021,N_954,N_36);
and U1022 (N_1022,N_75,N_32);
nor U1023 (N_1023,N_910,N_80);
nor U1024 (N_1024,N_777,N_11);
or U1025 (N_1025,N_12,N_241);
or U1026 (N_1026,N_808,N_389);
or U1027 (N_1027,N_508,N_687);
and U1028 (N_1028,N_3,N_805);
nor U1029 (N_1029,N_62,N_762);
nand U1030 (N_1030,N_159,N_442);
nand U1031 (N_1031,N_893,N_119);
and U1032 (N_1032,N_197,N_138);
or U1033 (N_1033,N_550,N_169);
nor U1034 (N_1034,N_529,N_700);
and U1035 (N_1035,N_649,N_533);
or U1036 (N_1036,N_149,N_839);
nand U1037 (N_1037,N_382,N_116);
xor U1038 (N_1038,N_443,N_727);
and U1039 (N_1039,N_625,N_621);
and U1040 (N_1040,N_20,N_305);
nand U1041 (N_1041,N_176,N_929);
nand U1042 (N_1042,N_426,N_221);
and U1043 (N_1043,N_204,N_501);
nand U1044 (N_1044,N_146,N_322);
and U1045 (N_1045,N_254,N_222);
or U1046 (N_1046,N_431,N_235);
or U1047 (N_1047,N_633,N_819);
and U1048 (N_1048,N_829,N_704);
nor U1049 (N_1049,N_866,N_694);
nand U1050 (N_1050,N_884,N_199);
nand U1051 (N_1051,N_814,N_25);
or U1052 (N_1052,N_765,N_581);
or U1053 (N_1053,N_91,N_558);
nor U1054 (N_1054,N_683,N_577);
nand U1055 (N_1055,N_680,N_478);
xnor U1056 (N_1056,N_984,N_962);
and U1057 (N_1057,N_679,N_709);
nor U1058 (N_1058,N_988,N_183);
and U1059 (N_1059,N_76,N_698);
nor U1060 (N_1060,N_368,N_733);
nand U1061 (N_1061,N_78,N_418);
and U1062 (N_1062,N_869,N_547);
or U1063 (N_1063,N_736,N_441);
and U1064 (N_1064,N_835,N_609);
nor U1065 (N_1065,N_29,N_187);
and U1066 (N_1066,N_74,N_15);
nand U1067 (N_1067,N_308,N_271);
and U1068 (N_1068,N_390,N_117);
or U1069 (N_1069,N_461,N_191);
nor U1070 (N_1070,N_695,N_190);
and U1071 (N_1071,N_947,N_641);
or U1072 (N_1072,N_261,N_68);
or U1073 (N_1073,N_598,N_297);
nand U1074 (N_1074,N_94,N_302);
nor U1075 (N_1075,N_239,N_26);
or U1076 (N_1076,N_454,N_265);
nor U1077 (N_1077,N_259,N_445);
nand U1078 (N_1078,N_152,N_941);
nand U1079 (N_1079,N_404,N_333);
nor U1080 (N_1080,N_579,N_425);
nor U1081 (N_1081,N_65,N_429);
or U1082 (N_1082,N_787,N_446);
or U1083 (N_1083,N_544,N_525);
nand U1084 (N_1084,N_854,N_52);
nor U1085 (N_1085,N_699,N_258);
xnor U1086 (N_1086,N_904,N_714);
and U1087 (N_1087,N_58,N_435);
or U1088 (N_1088,N_275,N_479);
nor U1089 (N_1089,N_635,N_810);
and U1090 (N_1090,N_539,N_689);
nand U1091 (N_1091,N_459,N_121);
nor U1092 (N_1092,N_434,N_346);
or U1093 (N_1093,N_396,N_337);
or U1094 (N_1094,N_964,N_717);
or U1095 (N_1095,N_937,N_280);
xor U1096 (N_1096,N_654,N_780);
nor U1097 (N_1097,N_413,N_705);
or U1098 (N_1098,N_86,N_453);
or U1099 (N_1099,N_427,N_245);
nand U1100 (N_1100,N_512,N_739);
nand U1101 (N_1101,N_16,N_597);
and U1102 (N_1102,N_201,N_31);
or U1103 (N_1103,N_132,N_220);
xor U1104 (N_1104,N_386,N_309);
nor U1105 (N_1105,N_402,N_619);
nor U1106 (N_1106,N_89,N_341);
or U1107 (N_1107,N_406,N_400);
or U1108 (N_1108,N_384,N_125);
or U1109 (N_1109,N_129,N_273);
or U1110 (N_1110,N_724,N_836);
nor U1111 (N_1111,N_150,N_526);
nor U1112 (N_1112,N_685,N_706);
nor U1113 (N_1113,N_69,N_817);
nor U1114 (N_1114,N_573,N_42);
xor U1115 (N_1115,N_812,N_411);
and U1116 (N_1116,N_976,N_800);
and U1117 (N_1117,N_55,N_54);
nor U1118 (N_1118,N_905,N_969);
nor U1119 (N_1119,N_462,N_440);
nand U1120 (N_1120,N_967,N_175);
nor U1121 (N_1121,N_591,N_416);
or U1122 (N_1122,N_766,N_846);
or U1123 (N_1123,N_472,N_668);
and U1124 (N_1124,N_898,N_553);
nor U1125 (N_1125,N_921,N_98);
or U1126 (N_1126,N_575,N_243);
or U1127 (N_1127,N_673,N_971);
or U1128 (N_1128,N_761,N_184);
and U1129 (N_1129,N_877,N_595);
xor U1130 (N_1130,N_136,N_521);
nor U1131 (N_1131,N_776,N_523);
nand U1132 (N_1132,N_934,N_624);
or U1133 (N_1133,N_848,N_276);
xor U1134 (N_1134,N_630,N_38);
or U1135 (N_1135,N_855,N_45);
nand U1136 (N_1136,N_593,N_952);
nor U1137 (N_1137,N_93,N_931);
nor U1138 (N_1138,N_87,N_725);
and U1139 (N_1139,N_233,N_614);
nor U1140 (N_1140,N_513,N_607);
or U1141 (N_1141,N_586,N_2);
or U1142 (N_1142,N_639,N_692);
nand U1143 (N_1143,N_299,N_540);
or U1144 (N_1144,N_291,N_141);
nand U1145 (N_1145,N_102,N_27);
nand U1146 (N_1146,N_415,N_943);
nor U1147 (N_1147,N_385,N_737);
nand U1148 (N_1148,N_155,N_251);
nor U1149 (N_1149,N_966,N_110);
or U1150 (N_1150,N_930,N_887);
nor U1151 (N_1151,N_773,N_70);
xnor U1152 (N_1152,N_329,N_659);
nor U1153 (N_1153,N_843,N_899);
xor U1154 (N_1154,N_578,N_332);
or U1155 (N_1155,N_397,N_349);
nand U1156 (N_1156,N_262,N_174);
nand U1157 (N_1157,N_552,N_466);
nand U1158 (N_1158,N_73,N_358);
or U1159 (N_1159,N_327,N_561);
nor U1160 (N_1160,N_514,N_809);
nor U1161 (N_1161,N_935,N_892);
and U1162 (N_1162,N_306,N_528);
and U1163 (N_1163,N_486,N_993);
nand U1164 (N_1164,N_430,N_263);
or U1165 (N_1165,N_361,N_63);
or U1166 (N_1166,N_860,N_193);
nor U1167 (N_1167,N_122,N_179);
xor U1168 (N_1168,N_342,N_285);
nor U1169 (N_1169,N_380,N_99);
and U1170 (N_1170,N_824,N_6);
nand U1171 (N_1171,N_747,N_331);
or U1172 (N_1172,N_876,N_139);
nand U1173 (N_1173,N_806,N_288);
nand U1174 (N_1174,N_912,N_144);
nor U1175 (N_1175,N_407,N_433);
nand U1176 (N_1176,N_170,N_950);
xnor U1177 (N_1177,N_489,N_363);
or U1178 (N_1178,N_370,N_785);
xnor U1179 (N_1179,N_881,N_662);
nand U1180 (N_1180,N_750,N_744);
nand U1181 (N_1181,N_173,N_658);
nor U1182 (N_1182,N_627,N_815);
and U1183 (N_1183,N_596,N_644);
or U1184 (N_1184,N_565,N_335);
xnor U1185 (N_1185,N_447,N_768);
nand U1186 (N_1186,N_795,N_973);
and U1187 (N_1187,N_353,N_827);
nand U1188 (N_1188,N_22,N_622);
nand U1189 (N_1189,N_350,N_557);
nor U1190 (N_1190,N_778,N_663);
and U1191 (N_1191,N_786,N_998);
nor U1192 (N_1192,N_517,N_480);
xor U1193 (N_1193,N_8,N_985);
and U1194 (N_1194,N_151,N_383);
nand U1195 (N_1195,N_974,N_913);
nand U1196 (N_1196,N_799,N_393);
xnor U1197 (N_1197,N_760,N_781);
and U1198 (N_1198,N_295,N_538);
xnor U1199 (N_1199,N_497,N_95);
nor U1200 (N_1200,N_247,N_779);
nor U1201 (N_1201,N_774,N_516);
nor U1202 (N_1202,N_448,N_325);
nand U1203 (N_1203,N_981,N_732);
nor U1204 (N_1204,N_311,N_468);
and U1205 (N_1205,N_645,N_378);
and U1206 (N_1206,N_19,N_688);
nand U1207 (N_1207,N_163,N_522);
nand U1208 (N_1208,N_825,N_455);
nor U1209 (N_1209,N_807,N_938);
or U1210 (N_1210,N_784,N_324);
nand U1211 (N_1211,N_272,N_405);
nand U1212 (N_1212,N_602,N_372);
and U1213 (N_1213,N_131,N_842);
nand U1214 (N_1214,N_908,N_589);
or U1215 (N_1215,N_334,N_643);
nor U1216 (N_1216,N_990,N_371);
nand U1217 (N_1217,N_255,N_657);
or U1218 (N_1218,N_59,N_588);
and U1219 (N_1219,N_373,N_828);
nor U1220 (N_1220,N_932,N_339);
nand U1221 (N_1221,N_248,N_127);
nor U1222 (N_1222,N_457,N_381);
nor U1223 (N_1223,N_72,N_225);
xnor U1224 (N_1224,N_494,N_105);
or U1225 (N_1225,N_185,N_865);
nand U1226 (N_1226,N_319,N_572);
or U1227 (N_1227,N_231,N_287);
nand U1228 (N_1228,N_519,N_475);
nor U1229 (N_1229,N_328,N_214);
nand U1230 (N_1230,N_50,N_603);
and U1231 (N_1231,N_347,N_878);
and U1232 (N_1232,N_118,N_524);
nor U1233 (N_1233,N_57,N_182);
or U1234 (N_1234,N_5,N_868);
or U1235 (N_1235,N_7,N_377);
nor U1236 (N_1236,N_71,N_536);
or U1237 (N_1237,N_296,N_492);
nor U1238 (N_1238,N_640,N_563);
nor U1239 (N_1239,N_888,N_758);
and U1240 (N_1240,N_219,N_104);
nand U1241 (N_1241,N_154,N_240);
or U1242 (N_1242,N_298,N_85);
or U1243 (N_1243,N_13,N_730);
or U1244 (N_1244,N_391,N_318);
or U1245 (N_1245,N_902,N_918);
or U1246 (N_1246,N_437,N_796);
nor U1247 (N_1247,N_92,N_953);
and U1248 (N_1248,N_604,N_782);
nor U1249 (N_1249,N_142,N_180);
nor U1250 (N_1250,N_21,N_830);
xor U1251 (N_1251,N_879,N_18);
or U1252 (N_1252,N_543,N_678);
or U1253 (N_1253,N_194,N_629);
nor U1254 (N_1254,N_177,N_849);
and U1255 (N_1255,N_844,N_249);
nand U1256 (N_1256,N_148,N_826);
nand U1257 (N_1257,N_560,N_230);
nand U1258 (N_1258,N_106,N_977);
nand U1259 (N_1259,N_882,N_994);
or U1260 (N_1260,N_650,N_126);
nand U1261 (N_1261,N_567,N_253);
and U1262 (N_1262,N_471,N_853);
and U1263 (N_1263,N_651,N_115);
nor U1264 (N_1264,N_906,N_34);
nor U1265 (N_1265,N_23,N_798);
and U1266 (N_1266,N_636,N_701);
xnor U1267 (N_1267,N_502,N_229);
nand U1268 (N_1268,N_49,N_965);
xnor U1269 (N_1269,N_606,N_601);
or U1270 (N_1270,N_554,N_611);
nand U1271 (N_1271,N_939,N_83);
or U1272 (N_1272,N_963,N_123);
xor U1273 (N_1273,N_703,N_542);
nand U1274 (N_1274,N_851,N_304);
nand U1275 (N_1275,N_234,N_556);
and U1276 (N_1276,N_820,N_160);
nor U1277 (N_1277,N_566,N_250);
or U1278 (N_1278,N_203,N_637);
or U1279 (N_1279,N_338,N_504);
or U1280 (N_1280,N_590,N_436);
and U1281 (N_1281,N_911,N_356);
and U1282 (N_1282,N_51,N_549);
or U1283 (N_1283,N_569,N_767);
nand U1284 (N_1284,N_999,N_321);
and U1285 (N_1285,N_483,N_834);
or U1286 (N_1286,N_511,N_195);
xor U1287 (N_1287,N_942,N_669);
and U1288 (N_1288,N_653,N_46);
and U1289 (N_1289,N_422,N_545);
nor U1290 (N_1290,N_460,N_344);
nor U1291 (N_1291,N_359,N_770);
nor U1292 (N_1292,N_726,N_37);
xnor U1293 (N_1293,N_541,N_367);
xor U1294 (N_1294,N_690,N_617);
or U1295 (N_1295,N_790,N_801);
nor U1296 (N_1296,N_14,N_895);
nand U1297 (N_1297,N_355,N_398);
nand U1298 (N_1298,N_0,N_507);
nand U1299 (N_1299,N_43,N_237);
nand U1300 (N_1300,N_438,N_804);
or U1301 (N_1301,N_84,N_900);
nand U1302 (N_1302,N_583,N_232);
nand U1303 (N_1303,N_940,N_210);
and U1304 (N_1304,N_164,N_919);
nor U1305 (N_1305,N_216,N_978);
and U1306 (N_1306,N_850,N_419);
nand U1307 (N_1307,N_682,N_211);
nand U1308 (N_1308,N_242,N_917);
nor U1309 (N_1309,N_61,N_108);
and U1310 (N_1310,N_996,N_864);
nor U1311 (N_1311,N_403,N_326);
nor U1312 (N_1312,N_307,N_354);
and U1313 (N_1313,N_920,N_56);
nand U1314 (N_1314,N_503,N_626);
or U1315 (N_1315,N_722,N_30);
nand U1316 (N_1316,N_671,N_469);
nand U1317 (N_1317,N_420,N_520);
and U1318 (N_1318,N_213,N_493);
nand U1319 (N_1319,N_281,N_364);
nand U1320 (N_1320,N_867,N_186);
nand U1321 (N_1321,N_379,N_496);
nand U1322 (N_1322,N_217,N_861);
or U1323 (N_1323,N_746,N_456);
nor U1324 (N_1324,N_257,N_476);
nor U1325 (N_1325,N_238,N_120);
and U1326 (N_1326,N_582,N_870);
xnor U1327 (N_1327,N_499,N_376);
and U1328 (N_1328,N_67,N_880);
nor U1329 (N_1329,N_515,N_236);
or U1330 (N_1330,N_79,N_916);
nand U1331 (N_1331,N_477,N_290);
nor U1332 (N_1332,N_44,N_293);
or U1333 (N_1333,N_791,N_113);
nor U1334 (N_1334,N_847,N_948);
and U1335 (N_1335,N_312,N_410);
nand U1336 (N_1336,N_665,N_39);
nor U1337 (N_1337,N_759,N_388);
nor U1338 (N_1338,N_252,N_599);
and U1339 (N_1339,N_64,N_666);
and U1340 (N_1340,N_485,N_114);
nor U1341 (N_1341,N_467,N_686);
or U1342 (N_1342,N_684,N_632);
or U1343 (N_1343,N_421,N_945);
or U1344 (N_1344,N_794,N_670);
and U1345 (N_1345,N_693,N_133);
or U1346 (N_1346,N_412,N_831);
nand U1347 (N_1347,N_638,N_320);
nand U1348 (N_1348,N_505,N_729);
or U1349 (N_1349,N_423,N_681);
nand U1350 (N_1350,N_28,N_564);
or U1351 (N_1351,N_161,N_753);
and U1352 (N_1352,N_147,N_955);
nand U1353 (N_1353,N_47,N_162);
nor U1354 (N_1354,N_209,N_982);
xor U1355 (N_1355,N_153,N_696);
nor U1356 (N_1356,N_17,N_444);
nand U1357 (N_1357,N_343,N_616);
and U1358 (N_1358,N_53,N_4);
or U1359 (N_1359,N_178,N_628);
nor U1360 (N_1360,N_283,N_465);
nand U1361 (N_1361,N_317,N_270);
nor U1362 (N_1362,N_10,N_224);
and U1363 (N_1363,N_562,N_387);
nor U1364 (N_1364,N_896,N_927);
nand U1365 (N_1365,N_769,N_764);
xor U1366 (N_1366,N_731,N_600);
or U1367 (N_1367,N_823,N_316);
and U1368 (N_1368,N_451,N_227);
or U1369 (N_1369,N_605,N_648);
or U1370 (N_1370,N_623,N_357);
nor U1371 (N_1371,N_674,N_340);
or U1372 (N_1372,N_789,N_960);
nor U1373 (N_1373,N_631,N_510);
nor U1374 (N_1374,N_463,N_756);
or U1375 (N_1375,N_949,N_661);
xor U1376 (N_1376,N_352,N_702);
xnor U1377 (N_1377,N_852,N_375);
or U1378 (N_1378,N_351,N_715);
and U1379 (N_1379,N_832,N_1);
or U1380 (N_1380,N_837,N_792);
nand U1381 (N_1381,N_266,N_995);
or U1382 (N_1382,N_646,N_748);
nor U1383 (N_1383,N_202,N_741);
or U1384 (N_1384,N_535,N_972);
nand U1385 (N_1385,N_957,N_909);
or U1386 (N_1386,N_675,N_813);
nand U1387 (N_1387,N_278,N_189);
nor U1388 (N_1388,N_439,N_156);
nand U1389 (N_1389,N_532,N_571);
and U1390 (N_1390,N_793,N_537);
nor U1391 (N_1391,N_260,N_188);
nor U1392 (N_1392,N_207,N_167);
nor U1393 (N_1393,N_713,N_664);
nand U1394 (N_1394,N_845,N_192);
nand U1395 (N_1395,N_101,N_897);
or U1396 (N_1396,N_200,N_576);
xor U1397 (N_1397,N_409,N_212);
or U1398 (N_1398,N_886,N_481);
or U1399 (N_1399,N_775,N_656);
nand U1400 (N_1400,N_301,N_171);
and U1401 (N_1401,N_48,N_907);
and U1402 (N_1402,N_464,N_274);
nor U1403 (N_1403,N_369,N_587);
and U1404 (N_1404,N_992,N_710);
and U1405 (N_1405,N_797,N_961);
xor U1406 (N_1406,N_482,N_286);
and U1407 (N_1407,N_915,N_734);
or U1408 (N_1408,N_652,N_933);
xnor U1409 (N_1409,N_612,N_223);
nand U1410 (N_1410,N_721,N_506);
and U1411 (N_1411,N_925,N_802);
nand U1412 (N_1412,N_208,N_124);
and U1413 (N_1413,N_226,N_822);
nor U1414 (N_1414,N_894,N_130);
or U1415 (N_1415,N_858,N_763);
or U1416 (N_1416,N_530,N_719);
or U1417 (N_1417,N_432,N_313);
or U1418 (N_1418,N_975,N_720);
or U1419 (N_1419,N_707,N_757);
nand U1420 (N_1420,N_755,N_128);
and U1421 (N_1421,N_647,N_345);
or U1422 (N_1422,N_24,N_883);
nand U1423 (N_1423,N_958,N_196);
and U1424 (N_1424,N_570,N_394);
nand U1425 (N_1425,N_559,N_488);
and U1426 (N_1426,N_360,N_749);
xnor U1427 (N_1427,N_135,N_165);
and U1428 (N_1428,N_277,N_655);
or U1429 (N_1429,N_9,N_97);
nor U1430 (N_1430,N_551,N_452);
and U1431 (N_1431,N_336,N_60);
and U1432 (N_1432,N_555,N_449);
or U1433 (N_1433,N_470,N_677);
nand U1434 (N_1434,N_923,N_109);
nor U1435 (N_1435,N_862,N_592);
nand U1436 (N_1436,N_613,N_527);
or U1437 (N_1437,N_314,N_743);
xor U1438 (N_1438,N_330,N_811);
and U1439 (N_1439,N_100,N_783);
xor U1440 (N_1440,N_711,N_158);
nand U1441 (N_1441,N_282,N_107);
nand U1442 (N_1442,N_246,N_228);
and U1443 (N_1443,N_803,N_735);
or U1444 (N_1444,N_424,N_484);
nand U1445 (N_1445,N_90,N_218);
nand U1446 (N_1446,N_205,N_279);
nor U1447 (N_1447,N_303,N_983);
nand U1448 (N_1448,N_594,N_103);
and U1449 (N_1449,N_676,N_716);
or U1450 (N_1450,N_642,N_81);
nand U1451 (N_1451,N_691,N_745);
nand U1452 (N_1452,N_401,N_672);
and U1453 (N_1453,N_901,N_574);
and U1454 (N_1454,N_365,N_491);
nand U1455 (N_1455,N_458,N_951);
nand U1456 (N_1456,N_970,N_922);
and U1457 (N_1457,N_956,N_979);
nand U1458 (N_1458,N_399,N_618);
or U1459 (N_1459,N_772,N_986);
nand U1460 (N_1460,N_788,N_428);
nand U1461 (N_1461,N_751,N_172);
and U1462 (N_1462,N_871,N_112);
xnor U1463 (N_1463,N_924,N_473);
and U1464 (N_1464,N_408,N_859);
nand U1465 (N_1465,N_968,N_885);
nor U1466 (N_1466,N_891,N_267);
xor U1467 (N_1467,N_348,N_740);
nand U1468 (N_1468,N_874,N_667);
and U1469 (N_1469,N_928,N_889);
nand U1470 (N_1470,N_531,N_585);
and U1471 (N_1471,N_315,N_546);
or U1472 (N_1472,N_518,N_269);
or U1473 (N_1473,N_718,N_395);
or U1474 (N_1474,N_991,N_534);
or U1475 (N_1475,N_754,N_268);
nor U1476 (N_1476,N_873,N_980);
or U1477 (N_1477,N_77,N_168);
and U1478 (N_1478,N_944,N_157);
and U1479 (N_1479,N_35,N_96);
nand U1480 (N_1480,N_215,N_111);
nor U1481 (N_1481,N_660,N_294);
or U1482 (N_1482,N_997,N_875);
nand U1483 (N_1483,N_362,N_366);
nand U1484 (N_1484,N_374,N_310);
or U1485 (N_1485,N_292,N_946);
and U1486 (N_1486,N_580,N_771);
and U1487 (N_1487,N_145,N_926);
nand U1488 (N_1488,N_500,N_509);
xor U1489 (N_1489,N_88,N_936);
and U1490 (N_1490,N_833,N_140);
or U1491 (N_1491,N_498,N_863);
nand U1492 (N_1492,N_66,N_495);
nor U1493 (N_1493,N_41,N_323);
nor U1494 (N_1494,N_181,N_490);
nand U1495 (N_1495,N_206,N_816);
or U1496 (N_1496,N_841,N_634);
and U1497 (N_1497,N_40,N_82);
or U1498 (N_1498,N_166,N_620);
and U1499 (N_1499,N_903,N_752);
nor U1500 (N_1500,N_718,N_541);
nor U1501 (N_1501,N_706,N_827);
nand U1502 (N_1502,N_277,N_754);
and U1503 (N_1503,N_428,N_366);
xor U1504 (N_1504,N_728,N_202);
nand U1505 (N_1505,N_167,N_768);
nor U1506 (N_1506,N_463,N_354);
nor U1507 (N_1507,N_176,N_876);
or U1508 (N_1508,N_832,N_272);
nand U1509 (N_1509,N_375,N_403);
nor U1510 (N_1510,N_244,N_774);
nand U1511 (N_1511,N_329,N_364);
nand U1512 (N_1512,N_181,N_872);
and U1513 (N_1513,N_993,N_505);
nor U1514 (N_1514,N_96,N_250);
or U1515 (N_1515,N_560,N_110);
or U1516 (N_1516,N_247,N_713);
nor U1517 (N_1517,N_282,N_376);
nor U1518 (N_1518,N_920,N_162);
or U1519 (N_1519,N_477,N_128);
nand U1520 (N_1520,N_694,N_356);
or U1521 (N_1521,N_878,N_876);
or U1522 (N_1522,N_187,N_276);
nand U1523 (N_1523,N_10,N_853);
nand U1524 (N_1524,N_395,N_694);
nor U1525 (N_1525,N_586,N_842);
and U1526 (N_1526,N_10,N_530);
nand U1527 (N_1527,N_388,N_866);
and U1528 (N_1528,N_996,N_80);
and U1529 (N_1529,N_589,N_616);
or U1530 (N_1530,N_941,N_548);
or U1531 (N_1531,N_520,N_745);
nand U1532 (N_1532,N_554,N_8);
nor U1533 (N_1533,N_762,N_54);
and U1534 (N_1534,N_967,N_439);
xor U1535 (N_1535,N_457,N_539);
nand U1536 (N_1536,N_793,N_388);
nand U1537 (N_1537,N_842,N_535);
nor U1538 (N_1538,N_397,N_482);
or U1539 (N_1539,N_381,N_123);
or U1540 (N_1540,N_137,N_117);
nor U1541 (N_1541,N_341,N_109);
nand U1542 (N_1542,N_888,N_869);
and U1543 (N_1543,N_397,N_892);
and U1544 (N_1544,N_512,N_188);
nand U1545 (N_1545,N_134,N_67);
nand U1546 (N_1546,N_282,N_865);
and U1547 (N_1547,N_359,N_158);
xor U1548 (N_1548,N_839,N_144);
nand U1549 (N_1549,N_877,N_335);
nor U1550 (N_1550,N_544,N_595);
xor U1551 (N_1551,N_216,N_454);
and U1552 (N_1552,N_535,N_159);
or U1553 (N_1553,N_78,N_728);
nor U1554 (N_1554,N_11,N_121);
nor U1555 (N_1555,N_824,N_24);
nand U1556 (N_1556,N_991,N_591);
and U1557 (N_1557,N_632,N_813);
and U1558 (N_1558,N_673,N_792);
nand U1559 (N_1559,N_963,N_954);
and U1560 (N_1560,N_332,N_722);
or U1561 (N_1561,N_614,N_751);
or U1562 (N_1562,N_814,N_988);
or U1563 (N_1563,N_134,N_239);
nor U1564 (N_1564,N_785,N_206);
nand U1565 (N_1565,N_361,N_185);
and U1566 (N_1566,N_309,N_398);
nor U1567 (N_1567,N_314,N_938);
and U1568 (N_1568,N_334,N_590);
xor U1569 (N_1569,N_610,N_844);
and U1570 (N_1570,N_121,N_817);
nand U1571 (N_1571,N_554,N_602);
nor U1572 (N_1572,N_588,N_365);
and U1573 (N_1573,N_965,N_544);
nand U1574 (N_1574,N_551,N_109);
nor U1575 (N_1575,N_606,N_942);
nand U1576 (N_1576,N_993,N_417);
and U1577 (N_1577,N_72,N_821);
or U1578 (N_1578,N_546,N_515);
nor U1579 (N_1579,N_963,N_472);
nand U1580 (N_1580,N_428,N_445);
and U1581 (N_1581,N_595,N_362);
and U1582 (N_1582,N_307,N_528);
nor U1583 (N_1583,N_519,N_893);
nand U1584 (N_1584,N_178,N_318);
and U1585 (N_1585,N_143,N_540);
and U1586 (N_1586,N_194,N_30);
nand U1587 (N_1587,N_339,N_1);
nand U1588 (N_1588,N_173,N_541);
nand U1589 (N_1589,N_237,N_904);
nor U1590 (N_1590,N_214,N_460);
nand U1591 (N_1591,N_556,N_927);
and U1592 (N_1592,N_398,N_273);
and U1593 (N_1593,N_613,N_292);
or U1594 (N_1594,N_722,N_919);
nor U1595 (N_1595,N_116,N_655);
nor U1596 (N_1596,N_182,N_526);
and U1597 (N_1597,N_885,N_931);
nand U1598 (N_1598,N_106,N_47);
xnor U1599 (N_1599,N_442,N_131);
or U1600 (N_1600,N_889,N_931);
and U1601 (N_1601,N_500,N_66);
or U1602 (N_1602,N_716,N_989);
or U1603 (N_1603,N_967,N_45);
nor U1604 (N_1604,N_814,N_192);
and U1605 (N_1605,N_877,N_873);
and U1606 (N_1606,N_195,N_752);
or U1607 (N_1607,N_942,N_37);
nor U1608 (N_1608,N_962,N_143);
or U1609 (N_1609,N_121,N_19);
and U1610 (N_1610,N_111,N_820);
nor U1611 (N_1611,N_190,N_155);
or U1612 (N_1612,N_133,N_268);
and U1613 (N_1613,N_822,N_418);
nand U1614 (N_1614,N_397,N_775);
nor U1615 (N_1615,N_756,N_33);
or U1616 (N_1616,N_5,N_620);
nand U1617 (N_1617,N_935,N_890);
nand U1618 (N_1618,N_936,N_115);
nor U1619 (N_1619,N_720,N_617);
or U1620 (N_1620,N_677,N_526);
nand U1621 (N_1621,N_121,N_366);
nand U1622 (N_1622,N_822,N_934);
nor U1623 (N_1623,N_670,N_140);
or U1624 (N_1624,N_238,N_142);
nand U1625 (N_1625,N_811,N_374);
nand U1626 (N_1626,N_444,N_38);
xor U1627 (N_1627,N_401,N_366);
or U1628 (N_1628,N_264,N_223);
nor U1629 (N_1629,N_205,N_412);
or U1630 (N_1630,N_428,N_588);
nand U1631 (N_1631,N_647,N_884);
xnor U1632 (N_1632,N_787,N_171);
xnor U1633 (N_1633,N_727,N_429);
nand U1634 (N_1634,N_141,N_791);
nand U1635 (N_1635,N_797,N_218);
or U1636 (N_1636,N_8,N_908);
and U1637 (N_1637,N_37,N_941);
nor U1638 (N_1638,N_281,N_171);
or U1639 (N_1639,N_600,N_126);
nand U1640 (N_1640,N_632,N_132);
or U1641 (N_1641,N_17,N_1);
nor U1642 (N_1642,N_326,N_58);
nand U1643 (N_1643,N_19,N_543);
and U1644 (N_1644,N_770,N_55);
or U1645 (N_1645,N_40,N_619);
nor U1646 (N_1646,N_596,N_386);
nand U1647 (N_1647,N_597,N_245);
and U1648 (N_1648,N_274,N_426);
and U1649 (N_1649,N_313,N_848);
and U1650 (N_1650,N_904,N_657);
or U1651 (N_1651,N_298,N_917);
nor U1652 (N_1652,N_908,N_23);
and U1653 (N_1653,N_733,N_267);
or U1654 (N_1654,N_616,N_764);
and U1655 (N_1655,N_508,N_71);
or U1656 (N_1656,N_953,N_114);
nor U1657 (N_1657,N_313,N_991);
or U1658 (N_1658,N_39,N_459);
or U1659 (N_1659,N_778,N_465);
or U1660 (N_1660,N_609,N_103);
nor U1661 (N_1661,N_211,N_355);
xor U1662 (N_1662,N_675,N_644);
nand U1663 (N_1663,N_959,N_354);
nand U1664 (N_1664,N_491,N_413);
nor U1665 (N_1665,N_851,N_817);
or U1666 (N_1666,N_495,N_471);
or U1667 (N_1667,N_88,N_616);
nand U1668 (N_1668,N_127,N_29);
and U1669 (N_1669,N_169,N_519);
nand U1670 (N_1670,N_689,N_878);
and U1671 (N_1671,N_136,N_612);
or U1672 (N_1672,N_996,N_320);
and U1673 (N_1673,N_744,N_596);
or U1674 (N_1674,N_878,N_546);
nand U1675 (N_1675,N_505,N_70);
and U1676 (N_1676,N_304,N_723);
nand U1677 (N_1677,N_582,N_88);
or U1678 (N_1678,N_69,N_291);
nand U1679 (N_1679,N_869,N_930);
xor U1680 (N_1680,N_56,N_655);
nand U1681 (N_1681,N_557,N_121);
or U1682 (N_1682,N_586,N_476);
and U1683 (N_1683,N_481,N_806);
nor U1684 (N_1684,N_25,N_621);
nor U1685 (N_1685,N_2,N_493);
nand U1686 (N_1686,N_688,N_916);
and U1687 (N_1687,N_377,N_651);
nand U1688 (N_1688,N_784,N_304);
or U1689 (N_1689,N_792,N_947);
nand U1690 (N_1690,N_983,N_896);
or U1691 (N_1691,N_717,N_774);
nand U1692 (N_1692,N_667,N_737);
xnor U1693 (N_1693,N_156,N_647);
nor U1694 (N_1694,N_328,N_888);
nand U1695 (N_1695,N_803,N_833);
xor U1696 (N_1696,N_411,N_593);
and U1697 (N_1697,N_384,N_113);
xor U1698 (N_1698,N_533,N_145);
nand U1699 (N_1699,N_906,N_11);
or U1700 (N_1700,N_928,N_344);
nand U1701 (N_1701,N_851,N_268);
or U1702 (N_1702,N_760,N_835);
and U1703 (N_1703,N_754,N_718);
xor U1704 (N_1704,N_677,N_489);
nor U1705 (N_1705,N_901,N_634);
nand U1706 (N_1706,N_272,N_751);
nand U1707 (N_1707,N_309,N_511);
or U1708 (N_1708,N_449,N_732);
and U1709 (N_1709,N_391,N_45);
and U1710 (N_1710,N_390,N_70);
nand U1711 (N_1711,N_942,N_254);
nor U1712 (N_1712,N_630,N_331);
nor U1713 (N_1713,N_275,N_435);
nand U1714 (N_1714,N_851,N_923);
or U1715 (N_1715,N_588,N_809);
and U1716 (N_1716,N_628,N_711);
nor U1717 (N_1717,N_846,N_209);
and U1718 (N_1718,N_849,N_287);
nor U1719 (N_1719,N_220,N_848);
nand U1720 (N_1720,N_791,N_454);
and U1721 (N_1721,N_337,N_826);
and U1722 (N_1722,N_917,N_479);
nor U1723 (N_1723,N_409,N_620);
and U1724 (N_1724,N_733,N_10);
and U1725 (N_1725,N_982,N_108);
nand U1726 (N_1726,N_744,N_688);
nor U1727 (N_1727,N_765,N_583);
nor U1728 (N_1728,N_30,N_985);
nand U1729 (N_1729,N_192,N_614);
xor U1730 (N_1730,N_645,N_296);
nor U1731 (N_1731,N_348,N_388);
or U1732 (N_1732,N_40,N_452);
nor U1733 (N_1733,N_942,N_453);
nand U1734 (N_1734,N_700,N_818);
nor U1735 (N_1735,N_111,N_633);
nand U1736 (N_1736,N_897,N_955);
nand U1737 (N_1737,N_779,N_558);
nor U1738 (N_1738,N_179,N_327);
nand U1739 (N_1739,N_90,N_640);
or U1740 (N_1740,N_637,N_244);
nor U1741 (N_1741,N_254,N_777);
nor U1742 (N_1742,N_49,N_118);
and U1743 (N_1743,N_685,N_627);
or U1744 (N_1744,N_355,N_525);
nor U1745 (N_1745,N_909,N_685);
and U1746 (N_1746,N_31,N_728);
nand U1747 (N_1747,N_999,N_612);
and U1748 (N_1748,N_879,N_960);
nand U1749 (N_1749,N_126,N_880);
and U1750 (N_1750,N_786,N_238);
nor U1751 (N_1751,N_786,N_66);
nand U1752 (N_1752,N_142,N_263);
nand U1753 (N_1753,N_398,N_90);
nand U1754 (N_1754,N_992,N_484);
nor U1755 (N_1755,N_90,N_459);
and U1756 (N_1756,N_435,N_62);
or U1757 (N_1757,N_800,N_447);
nand U1758 (N_1758,N_292,N_730);
and U1759 (N_1759,N_422,N_204);
nor U1760 (N_1760,N_263,N_23);
and U1761 (N_1761,N_774,N_743);
or U1762 (N_1762,N_486,N_393);
or U1763 (N_1763,N_179,N_333);
xnor U1764 (N_1764,N_274,N_44);
nor U1765 (N_1765,N_373,N_921);
nor U1766 (N_1766,N_26,N_820);
nor U1767 (N_1767,N_267,N_846);
or U1768 (N_1768,N_332,N_642);
nor U1769 (N_1769,N_642,N_763);
or U1770 (N_1770,N_824,N_891);
nor U1771 (N_1771,N_107,N_748);
nor U1772 (N_1772,N_700,N_916);
nand U1773 (N_1773,N_656,N_763);
and U1774 (N_1774,N_229,N_475);
xnor U1775 (N_1775,N_113,N_808);
nor U1776 (N_1776,N_504,N_227);
or U1777 (N_1777,N_16,N_940);
xor U1778 (N_1778,N_115,N_672);
or U1779 (N_1779,N_758,N_434);
or U1780 (N_1780,N_475,N_878);
and U1781 (N_1781,N_544,N_68);
or U1782 (N_1782,N_352,N_343);
nor U1783 (N_1783,N_369,N_674);
nand U1784 (N_1784,N_463,N_424);
xnor U1785 (N_1785,N_491,N_56);
and U1786 (N_1786,N_715,N_558);
nor U1787 (N_1787,N_894,N_851);
nor U1788 (N_1788,N_386,N_57);
and U1789 (N_1789,N_150,N_343);
and U1790 (N_1790,N_748,N_531);
nand U1791 (N_1791,N_404,N_875);
or U1792 (N_1792,N_783,N_422);
and U1793 (N_1793,N_285,N_113);
and U1794 (N_1794,N_412,N_116);
or U1795 (N_1795,N_46,N_932);
nand U1796 (N_1796,N_815,N_937);
or U1797 (N_1797,N_498,N_578);
and U1798 (N_1798,N_897,N_439);
nand U1799 (N_1799,N_994,N_354);
nor U1800 (N_1800,N_190,N_370);
nor U1801 (N_1801,N_157,N_391);
nor U1802 (N_1802,N_962,N_373);
or U1803 (N_1803,N_520,N_409);
nand U1804 (N_1804,N_344,N_12);
nand U1805 (N_1805,N_975,N_498);
or U1806 (N_1806,N_69,N_463);
or U1807 (N_1807,N_913,N_322);
nor U1808 (N_1808,N_107,N_874);
or U1809 (N_1809,N_731,N_302);
nor U1810 (N_1810,N_195,N_737);
and U1811 (N_1811,N_275,N_457);
or U1812 (N_1812,N_691,N_165);
or U1813 (N_1813,N_920,N_164);
nor U1814 (N_1814,N_844,N_43);
nand U1815 (N_1815,N_486,N_813);
nor U1816 (N_1816,N_198,N_537);
or U1817 (N_1817,N_848,N_30);
nand U1818 (N_1818,N_195,N_441);
and U1819 (N_1819,N_759,N_438);
nor U1820 (N_1820,N_860,N_18);
nand U1821 (N_1821,N_373,N_212);
nand U1822 (N_1822,N_430,N_942);
nor U1823 (N_1823,N_73,N_123);
and U1824 (N_1824,N_445,N_973);
nor U1825 (N_1825,N_695,N_649);
or U1826 (N_1826,N_545,N_388);
nand U1827 (N_1827,N_463,N_681);
nor U1828 (N_1828,N_73,N_685);
xor U1829 (N_1829,N_682,N_997);
nand U1830 (N_1830,N_817,N_605);
or U1831 (N_1831,N_399,N_831);
nand U1832 (N_1832,N_531,N_490);
xnor U1833 (N_1833,N_356,N_178);
xnor U1834 (N_1834,N_647,N_302);
nand U1835 (N_1835,N_220,N_145);
nor U1836 (N_1836,N_172,N_6);
and U1837 (N_1837,N_548,N_757);
and U1838 (N_1838,N_147,N_7);
or U1839 (N_1839,N_492,N_44);
nor U1840 (N_1840,N_794,N_772);
or U1841 (N_1841,N_203,N_854);
xnor U1842 (N_1842,N_101,N_147);
nor U1843 (N_1843,N_126,N_601);
or U1844 (N_1844,N_212,N_710);
nand U1845 (N_1845,N_406,N_107);
xnor U1846 (N_1846,N_175,N_826);
nor U1847 (N_1847,N_722,N_955);
and U1848 (N_1848,N_88,N_19);
nor U1849 (N_1849,N_142,N_541);
or U1850 (N_1850,N_411,N_927);
nor U1851 (N_1851,N_434,N_238);
and U1852 (N_1852,N_597,N_731);
or U1853 (N_1853,N_306,N_118);
or U1854 (N_1854,N_633,N_621);
and U1855 (N_1855,N_287,N_197);
nand U1856 (N_1856,N_849,N_604);
or U1857 (N_1857,N_504,N_332);
xor U1858 (N_1858,N_87,N_840);
xnor U1859 (N_1859,N_949,N_160);
nor U1860 (N_1860,N_18,N_116);
nor U1861 (N_1861,N_987,N_360);
or U1862 (N_1862,N_457,N_935);
nand U1863 (N_1863,N_266,N_414);
or U1864 (N_1864,N_49,N_613);
nand U1865 (N_1865,N_612,N_865);
xnor U1866 (N_1866,N_31,N_42);
and U1867 (N_1867,N_769,N_579);
xor U1868 (N_1868,N_581,N_333);
or U1869 (N_1869,N_289,N_424);
and U1870 (N_1870,N_619,N_820);
xnor U1871 (N_1871,N_234,N_217);
nand U1872 (N_1872,N_232,N_370);
and U1873 (N_1873,N_114,N_576);
or U1874 (N_1874,N_245,N_635);
nor U1875 (N_1875,N_51,N_435);
or U1876 (N_1876,N_298,N_51);
nand U1877 (N_1877,N_837,N_876);
nor U1878 (N_1878,N_469,N_256);
or U1879 (N_1879,N_389,N_339);
nand U1880 (N_1880,N_43,N_341);
nand U1881 (N_1881,N_78,N_680);
and U1882 (N_1882,N_791,N_703);
nand U1883 (N_1883,N_493,N_918);
nor U1884 (N_1884,N_812,N_825);
nor U1885 (N_1885,N_774,N_586);
nand U1886 (N_1886,N_624,N_567);
and U1887 (N_1887,N_315,N_586);
or U1888 (N_1888,N_59,N_5);
and U1889 (N_1889,N_418,N_371);
or U1890 (N_1890,N_231,N_572);
and U1891 (N_1891,N_871,N_520);
and U1892 (N_1892,N_554,N_513);
nand U1893 (N_1893,N_568,N_462);
nor U1894 (N_1894,N_469,N_810);
nand U1895 (N_1895,N_444,N_133);
nand U1896 (N_1896,N_581,N_907);
nand U1897 (N_1897,N_624,N_799);
nor U1898 (N_1898,N_199,N_90);
nand U1899 (N_1899,N_446,N_480);
and U1900 (N_1900,N_890,N_743);
nand U1901 (N_1901,N_211,N_328);
nand U1902 (N_1902,N_549,N_849);
nand U1903 (N_1903,N_537,N_554);
nor U1904 (N_1904,N_71,N_929);
nand U1905 (N_1905,N_950,N_550);
nor U1906 (N_1906,N_582,N_363);
xnor U1907 (N_1907,N_424,N_864);
nand U1908 (N_1908,N_273,N_162);
or U1909 (N_1909,N_211,N_615);
nor U1910 (N_1910,N_321,N_440);
nor U1911 (N_1911,N_126,N_842);
and U1912 (N_1912,N_671,N_679);
and U1913 (N_1913,N_620,N_573);
and U1914 (N_1914,N_287,N_420);
or U1915 (N_1915,N_705,N_70);
or U1916 (N_1916,N_696,N_437);
nand U1917 (N_1917,N_283,N_228);
nor U1918 (N_1918,N_99,N_402);
nand U1919 (N_1919,N_753,N_578);
and U1920 (N_1920,N_875,N_175);
and U1921 (N_1921,N_668,N_64);
nor U1922 (N_1922,N_276,N_721);
and U1923 (N_1923,N_696,N_211);
xor U1924 (N_1924,N_786,N_939);
and U1925 (N_1925,N_627,N_347);
or U1926 (N_1926,N_843,N_853);
or U1927 (N_1927,N_292,N_158);
or U1928 (N_1928,N_332,N_820);
nand U1929 (N_1929,N_76,N_778);
and U1930 (N_1930,N_189,N_816);
and U1931 (N_1931,N_595,N_775);
nand U1932 (N_1932,N_811,N_324);
nand U1933 (N_1933,N_119,N_135);
nor U1934 (N_1934,N_940,N_728);
nor U1935 (N_1935,N_449,N_45);
nand U1936 (N_1936,N_583,N_324);
nor U1937 (N_1937,N_509,N_318);
or U1938 (N_1938,N_675,N_270);
nand U1939 (N_1939,N_973,N_155);
xnor U1940 (N_1940,N_146,N_269);
and U1941 (N_1941,N_765,N_988);
xnor U1942 (N_1942,N_731,N_180);
nor U1943 (N_1943,N_663,N_572);
nand U1944 (N_1944,N_796,N_685);
nand U1945 (N_1945,N_364,N_901);
or U1946 (N_1946,N_449,N_452);
or U1947 (N_1947,N_235,N_323);
nor U1948 (N_1948,N_89,N_632);
and U1949 (N_1949,N_27,N_664);
xnor U1950 (N_1950,N_750,N_582);
xor U1951 (N_1951,N_599,N_36);
and U1952 (N_1952,N_330,N_215);
nor U1953 (N_1953,N_199,N_327);
and U1954 (N_1954,N_840,N_707);
nor U1955 (N_1955,N_244,N_756);
or U1956 (N_1956,N_346,N_632);
nand U1957 (N_1957,N_553,N_965);
xor U1958 (N_1958,N_59,N_764);
nand U1959 (N_1959,N_810,N_38);
xor U1960 (N_1960,N_146,N_119);
nand U1961 (N_1961,N_686,N_650);
nor U1962 (N_1962,N_928,N_273);
nand U1963 (N_1963,N_725,N_727);
nor U1964 (N_1964,N_690,N_113);
nor U1965 (N_1965,N_121,N_442);
nand U1966 (N_1966,N_437,N_964);
and U1967 (N_1967,N_236,N_617);
nand U1968 (N_1968,N_956,N_657);
nor U1969 (N_1969,N_438,N_424);
nand U1970 (N_1970,N_416,N_425);
and U1971 (N_1971,N_271,N_937);
nand U1972 (N_1972,N_849,N_819);
or U1973 (N_1973,N_732,N_213);
nand U1974 (N_1974,N_364,N_148);
or U1975 (N_1975,N_42,N_934);
nand U1976 (N_1976,N_39,N_685);
nand U1977 (N_1977,N_603,N_387);
or U1978 (N_1978,N_234,N_589);
or U1979 (N_1979,N_162,N_658);
nor U1980 (N_1980,N_352,N_250);
and U1981 (N_1981,N_103,N_894);
nand U1982 (N_1982,N_736,N_170);
or U1983 (N_1983,N_95,N_569);
and U1984 (N_1984,N_127,N_189);
nand U1985 (N_1985,N_785,N_883);
nor U1986 (N_1986,N_115,N_488);
nor U1987 (N_1987,N_456,N_770);
and U1988 (N_1988,N_398,N_839);
nand U1989 (N_1989,N_317,N_472);
nor U1990 (N_1990,N_505,N_214);
nor U1991 (N_1991,N_645,N_951);
nor U1992 (N_1992,N_144,N_572);
xnor U1993 (N_1993,N_918,N_975);
nor U1994 (N_1994,N_398,N_761);
xor U1995 (N_1995,N_135,N_686);
or U1996 (N_1996,N_389,N_63);
nand U1997 (N_1997,N_514,N_611);
and U1998 (N_1998,N_333,N_689);
and U1999 (N_1999,N_137,N_354);
nor U2000 (N_2000,N_1990,N_1957);
and U2001 (N_2001,N_1815,N_1065);
and U2002 (N_2002,N_1518,N_1090);
xnor U2003 (N_2003,N_1036,N_1249);
or U2004 (N_2004,N_1513,N_1810);
nand U2005 (N_2005,N_1212,N_1565);
or U2006 (N_2006,N_1052,N_1145);
nand U2007 (N_2007,N_1690,N_1181);
nor U2008 (N_2008,N_1646,N_1244);
nor U2009 (N_2009,N_1847,N_1750);
or U2010 (N_2010,N_1542,N_1410);
xnor U2011 (N_2011,N_1562,N_1377);
and U2012 (N_2012,N_1226,N_1074);
or U2013 (N_2013,N_1595,N_1762);
or U2014 (N_2014,N_1722,N_1723);
and U2015 (N_2015,N_1480,N_1239);
and U2016 (N_2016,N_1128,N_1834);
or U2017 (N_2017,N_1407,N_1799);
and U2018 (N_2018,N_1923,N_1812);
or U2019 (N_2019,N_1972,N_1311);
or U2020 (N_2020,N_1567,N_1152);
nor U2021 (N_2021,N_1912,N_1117);
nand U2022 (N_2022,N_1461,N_1832);
and U2023 (N_2023,N_1136,N_1375);
and U2024 (N_2024,N_1008,N_1376);
nor U2025 (N_2025,N_1089,N_1132);
nand U2026 (N_2026,N_1666,N_1974);
and U2027 (N_2027,N_1028,N_1302);
nor U2028 (N_2028,N_1395,N_1357);
xnor U2029 (N_2029,N_1669,N_1007);
or U2030 (N_2030,N_1107,N_1267);
nand U2031 (N_2031,N_1875,N_1932);
nand U2032 (N_2032,N_1412,N_1018);
and U2033 (N_2033,N_1822,N_1185);
xor U2034 (N_2034,N_1908,N_1930);
or U2035 (N_2035,N_1858,N_1933);
and U2036 (N_2036,N_1103,N_1829);
xor U2037 (N_2037,N_1577,N_1728);
or U2038 (N_2038,N_1886,N_1654);
or U2039 (N_2039,N_1396,N_1462);
and U2040 (N_2040,N_1205,N_1176);
or U2041 (N_2041,N_1866,N_1721);
nor U2042 (N_2042,N_1326,N_1110);
nand U2043 (N_2043,N_1439,N_1167);
nand U2044 (N_2044,N_1287,N_1266);
nor U2045 (N_2045,N_1759,N_1689);
nand U2046 (N_2046,N_1257,N_1673);
nor U2047 (N_2047,N_1884,N_1082);
or U2048 (N_2048,N_1989,N_1623);
nand U2049 (N_2049,N_1401,N_1503);
and U2050 (N_2050,N_1992,N_1231);
nor U2051 (N_2051,N_1220,N_1964);
and U2052 (N_2052,N_1645,N_1647);
nand U2053 (N_2053,N_1434,N_1484);
or U2054 (N_2054,N_1072,N_1246);
nor U2055 (N_2055,N_1897,N_1020);
or U2056 (N_2056,N_1352,N_1800);
or U2057 (N_2057,N_1383,N_1892);
nand U2058 (N_2058,N_1667,N_1155);
nand U2059 (N_2059,N_1003,N_1741);
nand U2060 (N_2060,N_1600,N_1200);
and U2061 (N_2061,N_1280,N_1675);
nand U2062 (N_2062,N_1787,N_1877);
and U2063 (N_2063,N_1902,N_1499);
and U2064 (N_2064,N_1941,N_1724);
and U2065 (N_2065,N_1609,N_1825);
xnor U2066 (N_2066,N_1315,N_1517);
or U2067 (N_2067,N_1732,N_1096);
or U2068 (N_2068,N_1910,N_1823);
nor U2069 (N_2069,N_1298,N_1471);
nor U2070 (N_2070,N_1795,N_1828);
or U2071 (N_2071,N_1129,N_1234);
nand U2072 (N_2072,N_1275,N_1947);
or U2073 (N_2073,N_1424,N_1995);
nand U2074 (N_2074,N_1663,N_1585);
or U2075 (N_2075,N_1093,N_1535);
nor U2076 (N_2076,N_1279,N_1092);
and U2077 (N_2077,N_1235,N_1073);
and U2078 (N_2078,N_1804,N_1778);
or U2079 (N_2079,N_1415,N_1843);
nor U2080 (N_2080,N_1077,N_1579);
nor U2081 (N_2081,N_1105,N_1729);
nand U2082 (N_2082,N_1274,N_1839);
xor U2083 (N_2083,N_1840,N_1699);
or U2084 (N_2084,N_1447,N_1848);
and U2085 (N_2085,N_1608,N_1534);
nand U2086 (N_2086,N_1460,N_1855);
nand U2087 (N_2087,N_1801,N_1824);
nor U2088 (N_2088,N_1004,N_1539);
nand U2089 (N_2089,N_1134,N_1939);
nor U2090 (N_2090,N_1632,N_1940);
or U2091 (N_2091,N_1363,N_1219);
nor U2092 (N_2092,N_1678,N_1861);
and U2093 (N_2093,N_1948,N_1969);
nand U2094 (N_2094,N_1813,N_1224);
nor U2095 (N_2095,N_1726,N_1162);
nand U2096 (N_2096,N_1159,N_1251);
and U2097 (N_2097,N_1803,N_1068);
nor U2098 (N_2098,N_1730,N_1924);
xor U2099 (N_2099,N_1954,N_1710);
and U2100 (N_2100,N_1657,N_1709);
nor U2101 (N_2101,N_1037,N_1355);
or U2102 (N_2102,N_1367,N_1474);
and U2103 (N_2103,N_1700,N_1818);
nand U2104 (N_2104,N_1138,N_1867);
or U2105 (N_2105,N_1399,N_1528);
nand U2106 (N_2106,N_1414,N_1889);
and U2107 (N_2107,N_1350,N_1264);
or U2108 (N_2108,N_1859,N_1745);
and U2109 (N_2109,N_1289,N_1540);
nor U2110 (N_2110,N_1056,N_1488);
or U2111 (N_2111,N_1035,N_1466);
and U2112 (N_2112,N_1064,N_1846);
nand U2113 (N_2113,N_1365,N_1602);
and U2114 (N_2114,N_1620,N_1334);
nand U2115 (N_2115,N_1760,N_1015);
or U2116 (N_2116,N_1017,N_1895);
xor U2117 (N_2117,N_1921,N_1561);
nor U2118 (N_2118,N_1121,N_1172);
and U2119 (N_2119,N_1069,N_1960);
nand U2120 (N_2120,N_1254,N_1446);
or U2121 (N_2121,N_1448,N_1512);
and U2122 (N_2122,N_1899,N_1309);
nand U2123 (N_2123,N_1477,N_1458);
nor U2124 (N_2124,N_1599,N_1907);
and U2125 (N_2125,N_1354,N_1175);
nor U2126 (N_2126,N_1321,N_1160);
and U2127 (N_2127,N_1597,N_1000);
nor U2128 (N_2128,N_1042,N_1099);
nand U2129 (N_2129,N_1358,N_1331);
or U2130 (N_2130,N_1656,N_1850);
or U2131 (N_2131,N_1413,N_1238);
nor U2132 (N_2132,N_1631,N_1630);
xnor U2133 (N_2133,N_1978,N_1353);
and U2134 (N_2134,N_1956,N_1157);
and U2135 (N_2135,N_1273,N_1717);
nor U2136 (N_2136,N_1455,N_1479);
xor U2137 (N_2137,N_1767,N_1796);
and U2138 (N_2138,N_1691,N_1366);
and U2139 (N_2139,N_1572,N_1204);
or U2140 (N_2140,N_1190,N_1133);
or U2141 (N_2141,N_1423,N_1523);
nand U2142 (N_2142,N_1165,N_1874);
or U2143 (N_2143,N_1113,N_1443);
nor U2144 (N_2144,N_1592,N_1229);
xor U2145 (N_2145,N_1747,N_1849);
and U2146 (N_2146,N_1676,N_1719);
nor U2147 (N_2147,N_1641,N_1494);
xnor U2148 (N_2148,N_1573,N_1958);
and U2149 (N_2149,N_1078,N_1684);
and U2150 (N_2150,N_1432,N_1148);
or U2151 (N_2151,N_1782,N_1705);
or U2152 (N_2152,N_1170,N_1883);
and U2153 (N_2153,N_1463,N_1307);
or U2154 (N_2154,N_1487,N_1870);
and U2155 (N_2155,N_1614,N_1559);
and U2156 (N_2156,N_1217,N_1481);
and U2157 (N_2157,N_1711,N_1335);
or U2158 (N_2158,N_1519,N_1739);
or U2159 (N_2159,N_1928,N_1900);
and U2160 (N_2160,N_1380,N_1293);
and U2161 (N_2161,N_1420,N_1061);
and U2162 (N_2162,N_1215,N_1290);
nor U2163 (N_2163,N_1637,N_1112);
xor U2164 (N_2164,N_1524,N_1119);
or U2165 (N_2165,N_1755,N_1306);
or U2166 (N_2166,N_1046,N_1416);
nand U2167 (N_2167,N_1374,N_1173);
and U2168 (N_2168,N_1533,N_1256);
xnor U2169 (N_2169,N_1680,N_1442);
or U2170 (N_2170,N_1342,N_1965);
nand U2171 (N_2171,N_1905,N_1744);
xor U2172 (N_2172,N_1490,N_1913);
or U2173 (N_2173,N_1979,N_1329);
nor U2174 (N_2174,N_1652,N_1685);
nor U2175 (N_2175,N_1023,N_1580);
and U2176 (N_2176,N_1070,N_1033);
nor U2177 (N_2177,N_1550,N_1716);
nor U2178 (N_2178,N_1362,N_1146);
nor U2179 (N_2179,N_1793,N_1005);
nor U2180 (N_2180,N_1594,N_1486);
or U2181 (N_2181,N_1139,N_1402);
and U2182 (N_2182,N_1440,N_1987);
nor U2183 (N_2183,N_1582,N_1098);
or U2184 (N_2184,N_1704,N_1878);
nor U2185 (N_2185,N_1553,N_1318);
or U2186 (N_2186,N_1201,N_1944);
nor U2187 (N_2187,N_1817,N_1384);
and U2188 (N_2188,N_1497,N_1196);
nand U2189 (N_2189,N_1919,N_1010);
or U2190 (N_2190,N_1598,N_1214);
nor U2191 (N_2191,N_1109,N_1976);
nor U2192 (N_2192,N_1322,N_1578);
xor U2193 (N_2193,N_1001,N_1154);
or U2194 (N_2194,N_1814,N_1775);
or U2195 (N_2195,N_1453,N_1225);
nand U2196 (N_2196,N_1498,N_1435);
or U2197 (N_2197,N_1457,N_1785);
and U2198 (N_2198,N_1016,N_1029);
xor U2199 (N_2199,N_1714,N_1391);
or U2200 (N_2200,N_1809,N_1830);
nor U2201 (N_2201,N_1537,N_1909);
or U2202 (N_2202,N_1625,N_1918);
and U2203 (N_2203,N_1199,N_1421);
nor U2204 (N_2204,N_1805,N_1655);
nor U2205 (N_2205,N_1863,N_1299);
nor U2206 (N_2206,N_1104,N_1769);
and U2207 (N_2207,N_1731,N_1981);
or U2208 (N_2208,N_1544,N_1125);
nand U2209 (N_2209,N_1991,N_1097);
and U2210 (N_2210,N_1048,N_1406);
nand U2211 (N_2211,N_1764,N_1885);
nand U2212 (N_2212,N_1515,N_1386);
or U2213 (N_2213,N_1341,N_1917);
nor U2214 (N_2214,N_1945,N_1083);
nor U2215 (N_2215,N_1915,N_1161);
nor U2216 (N_2216,N_1473,N_1313);
nor U2217 (N_2217,N_1323,N_1633);
or U2218 (N_2218,N_1737,N_1236);
and U2219 (N_2219,N_1169,N_1095);
nand U2220 (N_2220,N_1664,N_1937);
nor U2221 (N_2221,N_1692,N_1901);
nor U2222 (N_2222,N_1779,N_1891);
or U2223 (N_2223,N_1683,N_1182);
nand U2224 (N_2224,N_1429,N_1661);
nand U2225 (N_2225,N_1998,N_1888);
nand U2226 (N_2226,N_1411,N_1790);
and U2227 (N_2227,N_1557,N_1021);
nor U2228 (N_2228,N_1943,N_1610);
nand U2229 (N_2229,N_1950,N_1483);
or U2230 (N_2230,N_1327,N_1147);
and U2231 (N_2231,N_1062,N_1043);
nor U2232 (N_2232,N_1911,N_1314);
nor U2233 (N_2233,N_1624,N_1142);
xnor U2234 (N_2234,N_1961,N_1752);
or U2235 (N_2235,N_1725,N_1606);
and U2236 (N_2236,N_1938,N_1963);
nand U2237 (N_2237,N_1994,N_1348);
xnor U2238 (N_2238,N_1143,N_1328);
nor U2239 (N_2239,N_1949,N_1507);
and U2240 (N_2240,N_1916,N_1765);
nand U2241 (N_2241,N_1833,N_1130);
nor U2242 (N_2242,N_1845,N_1852);
nand U2243 (N_2243,N_1842,N_1511);
nor U2244 (N_2244,N_1316,N_1558);
and U2245 (N_2245,N_1389,N_1295);
nor U2246 (N_2246,N_1748,N_1456);
and U2247 (N_2247,N_1002,N_1491);
xnor U2248 (N_2248,N_1955,N_1403);
nor U2249 (N_2249,N_1977,N_1291);
and U2250 (N_2250,N_1393,N_1914);
or U2251 (N_2251,N_1640,N_1548);
and U2252 (N_2252,N_1184,N_1698);
and U2253 (N_2253,N_1872,N_1135);
and U2254 (N_2254,N_1297,N_1011);
or U2255 (N_2255,N_1826,N_1896);
and U2256 (N_2256,N_1191,N_1492);
or U2257 (N_2257,N_1634,N_1243);
xnor U2258 (N_2258,N_1265,N_1574);
or U2259 (N_2259,N_1712,N_1970);
and U2260 (N_2260,N_1400,N_1233);
xor U2261 (N_2261,N_1319,N_1255);
nor U2262 (N_2262,N_1687,N_1301);
nand U2263 (N_2263,N_1733,N_1985);
and U2264 (N_2264,N_1869,N_1772);
nor U2265 (N_2265,N_1694,N_1276);
or U2266 (N_2266,N_1252,N_1838);
xnor U2267 (N_2267,N_1195,N_1756);
nor U2268 (N_2268,N_1841,N_1807);
xnor U2269 (N_2269,N_1080,N_1213);
xor U2270 (N_2270,N_1962,N_1405);
and U2271 (N_2271,N_1368,N_1619);
nor U2272 (N_2272,N_1397,N_1754);
and U2273 (N_2273,N_1178,N_1856);
nor U2274 (N_2274,N_1272,N_1164);
nor U2275 (N_2275,N_1269,N_1102);
nand U2276 (N_2276,N_1464,N_1379);
nand U2277 (N_2277,N_1681,N_1115);
and U2278 (N_2278,N_1171,N_1973);
xnor U2279 (N_2279,N_1552,N_1753);
nand U2280 (N_2280,N_1340,N_1952);
and U2281 (N_2281,N_1211,N_1288);
or U2282 (N_2282,N_1166,N_1783);
nor U2283 (N_2283,N_1345,N_1094);
or U2284 (N_2284,N_1108,N_1975);
or U2285 (N_2285,N_1882,N_1871);
nor U2286 (N_2286,N_1931,N_1612);
or U2287 (N_2287,N_1708,N_1425);
nor U2288 (N_2288,N_1873,N_1419);
nand U2289 (N_2289,N_1385,N_1569);
and U2290 (N_2290,N_1639,N_1715);
nor U2291 (N_2291,N_1501,N_1674);
nand U2292 (N_2292,N_1551,N_1727);
or U2293 (N_2293,N_1862,N_1476);
nand U2294 (N_2294,N_1151,N_1247);
nor U2295 (N_2295,N_1027,N_1971);
or U2296 (N_2296,N_1045,N_1696);
nand U2297 (N_2297,N_1038,N_1118);
xor U2298 (N_2298,N_1720,N_1898);
and U2299 (N_2299,N_1131,N_1041);
and U2300 (N_2300,N_1012,N_1966);
nor U2301 (N_2301,N_1428,N_1270);
nand U2302 (N_2302,N_1780,N_1359);
and U2303 (N_2303,N_1054,N_1194);
nor U2304 (N_2304,N_1051,N_1317);
and U2305 (N_2305,N_1050,N_1679);
and U2306 (N_2306,N_1344,N_1438);
or U2307 (N_2307,N_1347,N_1242);
or U2308 (N_2308,N_1268,N_1177);
nor U2309 (N_2309,N_1549,N_1183);
nor U2310 (N_2310,N_1677,N_1114);
and U2311 (N_2311,N_1806,N_1587);
and U2312 (N_2312,N_1980,N_1493);
or U2313 (N_2313,N_1394,N_1541);
xnor U2314 (N_2314,N_1308,N_1203);
and U2315 (N_2315,N_1066,N_1635);
nand U2316 (N_2316,N_1390,N_1786);
nor U2317 (N_2317,N_1221,N_1116);
nand U2318 (N_2318,N_1703,N_1351);
and U2319 (N_2319,N_1450,N_1188);
or U2320 (N_2320,N_1120,N_1819);
nand U2321 (N_2321,N_1568,N_1665);
nor U2322 (N_2322,N_1749,N_1929);
nand U2323 (N_2323,N_1469,N_1189);
nand U2324 (N_2324,N_1736,N_1281);
nand U2325 (N_2325,N_1589,N_1470);
and U2326 (N_2326,N_1526,N_1075);
and U2327 (N_2327,N_1153,N_1361);
or U2328 (N_2328,N_1248,N_1485);
and U2329 (N_2329,N_1508,N_1601);
xor U2330 (N_2330,N_1454,N_1427);
and U2331 (N_2331,N_1868,N_1777);
nand U2332 (N_2332,N_1701,N_1851);
and U2333 (N_2333,N_1022,N_1658);
nand U2334 (N_2334,N_1570,N_1381);
nor U2335 (N_2335,N_1791,N_1997);
nand U2336 (N_2336,N_1100,N_1478);
or U2337 (N_2337,N_1312,N_1071);
nand U2338 (N_2338,N_1032,N_1360);
and U2339 (N_2339,N_1536,N_1014);
nor U2340 (N_2340,N_1336,N_1996);
nor U2341 (N_2341,N_1343,N_1659);
nand U2342 (N_2342,N_1079,N_1398);
nand U2343 (N_2343,N_1575,N_1983);
nand U2344 (N_2344,N_1325,N_1529);
nor U2345 (N_2345,N_1583,N_1934);
nand U2346 (N_2346,N_1686,N_1670);
nand U2347 (N_2347,N_1009,N_1628);
nand U2348 (N_2348,N_1253,N_1743);
and U2349 (N_2349,N_1788,N_1993);
and U2350 (N_2350,N_1422,N_1451);
nand U2351 (N_2351,N_1449,N_1174);
or U2352 (N_2352,N_1141,N_1651);
or U2353 (N_2353,N_1636,N_1206);
nor U2354 (N_2354,N_1887,N_1209);
nor U2355 (N_2355,N_1649,N_1798);
nor U2356 (N_2356,N_1864,N_1564);
or U2357 (N_2357,N_1546,N_1495);
nor U2358 (N_2358,N_1218,N_1693);
nor U2359 (N_2359,N_1827,N_1586);
xnor U2360 (N_2360,N_1999,N_1025);
or U2361 (N_2361,N_1444,N_1835);
and U2362 (N_2362,N_1101,N_1417);
or U2363 (N_2363,N_1617,N_1522);
and U2364 (N_2364,N_1613,N_1713);
or U2365 (N_2365,N_1738,N_1590);
xor U2366 (N_2366,N_1063,N_1802);
or U2367 (N_2367,N_1426,N_1857);
or U2368 (N_2368,N_1773,N_1500);
and U2369 (N_2369,N_1509,N_1240);
and U2370 (N_2370,N_1452,N_1660);
nand U2371 (N_2371,N_1571,N_1387);
nor U2372 (N_2372,N_1740,N_1404);
nand U2373 (N_2373,N_1521,N_1925);
or U2374 (N_2374,N_1137,N_1808);
nand U2375 (N_2375,N_1149,N_1250);
or U2376 (N_2376,N_1186,N_1418);
nor U2377 (N_2377,N_1208,N_1935);
xnor U2378 (N_2378,N_1927,N_1262);
and U2379 (N_2379,N_1538,N_1922);
nand U2380 (N_2380,N_1192,N_1735);
and U2381 (N_2381,N_1688,N_1904);
or U2382 (N_2382,N_1627,N_1520);
nor U2383 (N_2383,N_1763,N_1081);
or U2384 (N_2384,N_1761,N_1084);
and U2385 (N_2385,N_1742,N_1860);
and U2386 (N_2386,N_1126,N_1707);
or U2387 (N_2387,N_1324,N_1230);
and U2388 (N_2388,N_1758,N_1622);
nor U2389 (N_2389,N_1320,N_1953);
nand U2390 (N_2390,N_1668,N_1545);
nand U2391 (N_2391,N_1525,N_1163);
and U2392 (N_2392,N_1346,N_1445);
and U2393 (N_2393,N_1168,N_1333);
or U2394 (N_2394,N_1278,N_1890);
nor U2395 (N_2395,N_1431,N_1926);
and U2396 (N_2396,N_1468,N_1106);
nand U2397 (N_2397,N_1467,N_1283);
nor U2398 (N_2398,N_1127,N_1088);
and U2399 (N_2399,N_1560,N_1370);
or U2400 (N_2400,N_1197,N_1356);
or U2401 (N_2401,N_1332,N_1202);
and U2402 (N_2402,N_1844,N_1210);
and U2403 (N_2403,N_1502,N_1430);
or U2404 (N_2404,N_1123,N_1330);
and U2405 (N_2405,N_1702,N_1496);
nor U2406 (N_2406,N_1055,N_1034);
or U2407 (N_2407,N_1364,N_1751);
nand U2408 (N_2408,N_1300,N_1768);
nand U2409 (N_2409,N_1019,N_1441);
or U2410 (N_2410,N_1604,N_1338);
nand U2411 (N_2411,N_1903,N_1388);
and U2412 (N_2412,N_1682,N_1555);
nand U2413 (N_2413,N_1662,N_1530);
nor U2414 (N_2414,N_1124,N_1816);
nand U2415 (N_2415,N_1285,N_1626);
nand U2416 (N_2416,N_1556,N_1643);
or U2417 (N_2417,N_1472,N_1820);
or U2418 (N_2418,N_1642,N_1672);
or U2419 (N_2419,N_1607,N_1227);
or U2420 (N_2420,N_1091,N_1067);
and U2421 (N_2421,N_1294,N_1505);
nand U2422 (N_2422,N_1876,N_1554);
and U2423 (N_2423,N_1865,N_1766);
xor U2424 (N_2424,N_1946,N_1282);
and U2425 (N_2425,N_1076,N_1349);
nand U2426 (N_2426,N_1611,N_1409);
xor U2427 (N_2427,N_1504,N_1581);
or U2428 (N_2428,N_1303,N_1638);
nand U2429 (N_2429,N_1261,N_1831);
xnor U2430 (N_2430,N_1771,N_1369);
nor U2431 (N_2431,N_1158,N_1543);
nand U2432 (N_2432,N_1514,N_1144);
and U2433 (N_2433,N_1087,N_1263);
nor U2434 (N_2434,N_1789,N_1982);
xnor U2435 (N_2435,N_1770,N_1854);
nor U2436 (N_2436,N_1193,N_1207);
nor U2437 (N_2437,N_1223,N_1988);
nand U2438 (N_2438,N_1967,N_1697);
nand U2439 (N_2439,N_1706,N_1436);
nand U2440 (N_2440,N_1811,N_1006);
nand U2441 (N_2441,N_1968,N_1237);
or U2442 (N_2442,N_1942,N_1746);
nand U2443 (N_2443,N_1792,N_1629);
and U2444 (N_2444,N_1615,N_1920);
and U2445 (N_2445,N_1049,N_1618);
or U2446 (N_2446,N_1337,N_1228);
nand U2447 (N_2447,N_1527,N_1584);
nor U2448 (N_2448,N_1296,N_1437);
nor U2449 (N_2449,N_1596,N_1057);
nand U2450 (N_2450,N_1603,N_1563);
or U2451 (N_2451,N_1371,N_1986);
or U2452 (N_2452,N_1111,N_1259);
or U2453 (N_2453,N_1122,N_1881);
nand U2454 (N_2454,N_1030,N_1757);
nor U2455 (N_2455,N_1392,N_1459);
nor U2456 (N_2456,N_1836,N_1059);
nor U2457 (N_2457,N_1284,N_1531);
and U2458 (N_2458,N_1286,N_1382);
nand U2459 (N_2459,N_1644,N_1893);
and U2460 (N_2460,N_1516,N_1216);
nand U2461 (N_2461,N_1794,N_1140);
and U2462 (N_2462,N_1653,N_1489);
or U2463 (N_2463,N_1879,N_1040);
xor U2464 (N_2464,N_1053,N_1566);
nor U2465 (N_2465,N_1482,N_1013);
or U2466 (N_2466,N_1305,N_1837);
nor U2467 (N_2467,N_1510,N_1245);
and U2468 (N_2468,N_1150,N_1047);
nor U2469 (N_2469,N_1547,N_1532);
and U2470 (N_2470,N_1718,N_1086);
or U2471 (N_2471,N_1621,N_1776);
or U2472 (N_2472,N_1588,N_1058);
and U2473 (N_2473,N_1085,N_1821);
or U2474 (N_2474,N_1734,N_1372);
or U2475 (N_2475,N_1906,N_1180);
or U2476 (N_2476,N_1465,N_1187);
xor U2477 (N_2477,N_1339,N_1222);
xor U2478 (N_2478,N_1671,N_1576);
and U2479 (N_2479,N_1277,N_1039);
xnor U2480 (N_2480,N_1593,N_1241);
or U2481 (N_2481,N_1894,N_1271);
nand U2482 (N_2482,N_1198,N_1784);
or U2483 (N_2483,N_1260,N_1310);
and U2484 (N_2484,N_1024,N_1648);
nor U2485 (N_2485,N_1951,N_1304);
and U2486 (N_2486,N_1774,N_1650);
nand U2487 (N_2487,N_1616,N_1475);
nor U2488 (N_2488,N_1060,N_1258);
or U2489 (N_2489,N_1695,N_1373);
nand U2490 (N_2490,N_1292,N_1506);
nor U2491 (N_2491,N_1031,N_1781);
xnor U2492 (N_2492,N_1044,N_1959);
xor U2493 (N_2493,N_1605,N_1179);
and U2494 (N_2494,N_1232,N_1026);
and U2495 (N_2495,N_1591,N_1408);
nand U2496 (N_2496,N_1936,N_1880);
xnor U2497 (N_2497,N_1433,N_1797);
nand U2498 (N_2498,N_1984,N_1156);
xor U2499 (N_2499,N_1853,N_1378);
nor U2500 (N_2500,N_1075,N_1194);
nand U2501 (N_2501,N_1155,N_1301);
nand U2502 (N_2502,N_1501,N_1897);
and U2503 (N_2503,N_1885,N_1994);
and U2504 (N_2504,N_1064,N_1987);
and U2505 (N_2505,N_1151,N_1505);
xor U2506 (N_2506,N_1006,N_1628);
and U2507 (N_2507,N_1046,N_1668);
or U2508 (N_2508,N_1842,N_1736);
or U2509 (N_2509,N_1948,N_1816);
nor U2510 (N_2510,N_1713,N_1592);
and U2511 (N_2511,N_1165,N_1986);
nor U2512 (N_2512,N_1881,N_1723);
or U2513 (N_2513,N_1387,N_1843);
nor U2514 (N_2514,N_1534,N_1276);
or U2515 (N_2515,N_1154,N_1036);
and U2516 (N_2516,N_1367,N_1767);
xor U2517 (N_2517,N_1682,N_1756);
nand U2518 (N_2518,N_1436,N_1232);
nand U2519 (N_2519,N_1284,N_1306);
or U2520 (N_2520,N_1847,N_1587);
nor U2521 (N_2521,N_1251,N_1347);
or U2522 (N_2522,N_1691,N_1618);
and U2523 (N_2523,N_1657,N_1205);
and U2524 (N_2524,N_1946,N_1286);
xor U2525 (N_2525,N_1058,N_1918);
nor U2526 (N_2526,N_1200,N_1284);
nor U2527 (N_2527,N_1226,N_1734);
and U2528 (N_2528,N_1218,N_1875);
nor U2529 (N_2529,N_1900,N_1005);
or U2530 (N_2530,N_1802,N_1053);
and U2531 (N_2531,N_1306,N_1365);
nand U2532 (N_2532,N_1349,N_1964);
nand U2533 (N_2533,N_1362,N_1101);
nand U2534 (N_2534,N_1941,N_1784);
nand U2535 (N_2535,N_1926,N_1590);
xor U2536 (N_2536,N_1036,N_1044);
nand U2537 (N_2537,N_1450,N_1086);
or U2538 (N_2538,N_1311,N_1570);
nor U2539 (N_2539,N_1568,N_1150);
nor U2540 (N_2540,N_1260,N_1822);
and U2541 (N_2541,N_1385,N_1298);
nand U2542 (N_2542,N_1515,N_1323);
or U2543 (N_2543,N_1621,N_1661);
and U2544 (N_2544,N_1221,N_1584);
nand U2545 (N_2545,N_1708,N_1582);
nand U2546 (N_2546,N_1744,N_1227);
nand U2547 (N_2547,N_1274,N_1766);
nand U2548 (N_2548,N_1533,N_1277);
xor U2549 (N_2549,N_1526,N_1062);
or U2550 (N_2550,N_1368,N_1110);
xnor U2551 (N_2551,N_1109,N_1231);
or U2552 (N_2552,N_1689,N_1139);
nand U2553 (N_2553,N_1412,N_1269);
or U2554 (N_2554,N_1320,N_1846);
or U2555 (N_2555,N_1468,N_1560);
xor U2556 (N_2556,N_1237,N_1226);
nand U2557 (N_2557,N_1757,N_1006);
nand U2558 (N_2558,N_1635,N_1460);
nor U2559 (N_2559,N_1918,N_1144);
and U2560 (N_2560,N_1363,N_1722);
nor U2561 (N_2561,N_1722,N_1136);
xnor U2562 (N_2562,N_1126,N_1387);
nand U2563 (N_2563,N_1770,N_1785);
and U2564 (N_2564,N_1593,N_1660);
and U2565 (N_2565,N_1512,N_1210);
nor U2566 (N_2566,N_1266,N_1045);
nor U2567 (N_2567,N_1479,N_1751);
and U2568 (N_2568,N_1454,N_1913);
nand U2569 (N_2569,N_1944,N_1185);
xnor U2570 (N_2570,N_1595,N_1063);
or U2571 (N_2571,N_1888,N_1446);
or U2572 (N_2572,N_1899,N_1747);
and U2573 (N_2573,N_1612,N_1444);
and U2574 (N_2574,N_1570,N_1691);
or U2575 (N_2575,N_1572,N_1407);
and U2576 (N_2576,N_1598,N_1792);
and U2577 (N_2577,N_1772,N_1561);
or U2578 (N_2578,N_1786,N_1336);
nand U2579 (N_2579,N_1532,N_1100);
and U2580 (N_2580,N_1604,N_1605);
nor U2581 (N_2581,N_1518,N_1805);
nor U2582 (N_2582,N_1744,N_1841);
nand U2583 (N_2583,N_1789,N_1405);
or U2584 (N_2584,N_1722,N_1862);
or U2585 (N_2585,N_1802,N_1632);
nor U2586 (N_2586,N_1228,N_1836);
xor U2587 (N_2587,N_1541,N_1793);
and U2588 (N_2588,N_1444,N_1474);
nor U2589 (N_2589,N_1360,N_1605);
or U2590 (N_2590,N_1824,N_1598);
nand U2591 (N_2591,N_1049,N_1986);
nor U2592 (N_2592,N_1048,N_1280);
nand U2593 (N_2593,N_1929,N_1094);
nor U2594 (N_2594,N_1964,N_1235);
xor U2595 (N_2595,N_1802,N_1044);
or U2596 (N_2596,N_1260,N_1709);
nand U2597 (N_2597,N_1796,N_1159);
or U2598 (N_2598,N_1612,N_1329);
or U2599 (N_2599,N_1918,N_1231);
xnor U2600 (N_2600,N_1450,N_1630);
xor U2601 (N_2601,N_1335,N_1070);
or U2602 (N_2602,N_1122,N_1094);
or U2603 (N_2603,N_1622,N_1319);
nor U2604 (N_2604,N_1191,N_1445);
nor U2605 (N_2605,N_1896,N_1192);
xnor U2606 (N_2606,N_1702,N_1194);
or U2607 (N_2607,N_1431,N_1140);
nand U2608 (N_2608,N_1475,N_1703);
or U2609 (N_2609,N_1072,N_1109);
nand U2610 (N_2610,N_1198,N_1116);
nor U2611 (N_2611,N_1866,N_1753);
nor U2612 (N_2612,N_1859,N_1311);
nand U2613 (N_2613,N_1834,N_1480);
xor U2614 (N_2614,N_1344,N_1610);
nand U2615 (N_2615,N_1823,N_1507);
nand U2616 (N_2616,N_1035,N_1899);
nand U2617 (N_2617,N_1276,N_1549);
and U2618 (N_2618,N_1403,N_1208);
or U2619 (N_2619,N_1313,N_1773);
or U2620 (N_2620,N_1720,N_1355);
nor U2621 (N_2621,N_1801,N_1283);
nand U2622 (N_2622,N_1292,N_1744);
nor U2623 (N_2623,N_1289,N_1811);
or U2624 (N_2624,N_1260,N_1607);
xnor U2625 (N_2625,N_1864,N_1678);
or U2626 (N_2626,N_1610,N_1011);
nand U2627 (N_2627,N_1251,N_1521);
xnor U2628 (N_2628,N_1947,N_1727);
nor U2629 (N_2629,N_1611,N_1947);
or U2630 (N_2630,N_1524,N_1084);
or U2631 (N_2631,N_1471,N_1431);
nand U2632 (N_2632,N_1358,N_1102);
and U2633 (N_2633,N_1108,N_1949);
nand U2634 (N_2634,N_1796,N_1898);
nor U2635 (N_2635,N_1128,N_1417);
or U2636 (N_2636,N_1584,N_1028);
nand U2637 (N_2637,N_1672,N_1741);
and U2638 (N_2638,N_1947,N_1062);
or U2639 (N_2639,N_1868,N_1565);
or U2640 (N_2640,N_1635,N_1647);
or U2641 (N_2641,N_1257,N_1193);
nand U2642 (N_2642,N_1314,N_1235);
and U2643 (N_2643,N_1876,N_1592);
or U2644 (N_2644,N_1218,N_1142);
or U2645 (N_2645,N_1717,N_1812);
and U2646 (N_2646,N_1681,N_1882);
nor U2647 (N_2647,N_1032,N_1422);
and U2648 (N_2648,N_1818,N_1922);
or U2649 (N_2649,N_1131,N_1804);
or U2650 (N_2650,N_1312,N_1126);
nand U2651 (N_2651,N_1606,N_1659);
or U2652 (N_2652,N_1469,N_1243);
nor U2653 (N_2653,N_1805,N_1997);
or U2654 (N_2654,N_1284,N_1891);
or U2655 (N_2655,N_1202,N_1705);
nor U2656 (N_2656,N_1388,N_1976);
nand U2657 (N_2657,N_1110,N_1484);
or U2658 (N_2658,N_1567,N_1068);
nand U2659 (N_2659,N_1916,N_1098);
and U2660 (N_2660,N_1376,N_1231);
or U2661 (N_2661,N_1459,N_1237);
xor U2662 (N_2662,N_1592,N_1514);
nor U2663 (N_2663,N_1685,N_1838);
or U2664 (N_2664,N_1537,N_1902);
nand U2665 (N_2665,N_1969,N_1650);
xnor U2666 (N_2666,N_1295,N_1650);
and U2667 (N_2667,N_1926,N_1875);
and U2668 (N_2668,N_1273,N_1955);
nor U2669 (N_2669,N_1539,N_1890);
or U2670 (N_2670,N_1266,N_1809);
nand U2671 (N_2671,N_1129,N_1735);
and U2672 (N_2672,N_1607,N_1997);
nor U2673 (N_2673,N_1773,N_1130);
nand U2674 (N_2674,N_1266,N_1651);
nand U2675 (N_2675,N_1078,N_1823);
or U2676 (N_2676,N_1390,N_1703);
or U2677 (N_2677,N_1493,N_1791);
nand U2678 (N_2678,N_1592,N_1712);
nor U2679 (N_2679,N_1626,N_1853);
xor U2680 (N_2680,N_1312,N_1891);
nor U2681 (N_2681,N_1866,N_1357);
nor U2682 (N_2682,N_1872,N_1159);
xor U2683 (N_2683,N_1546,N_1151);
nor U2684 (N_2684,N_1049,N_1885);
nor U2685 (N_2685,N_1581,N_1351);
and U2686 (N_2686,N_1415,N_1340);
or U2687 (N_2687,N_1040,N_1845);
nand U2688 (N_2688,N_1379,N_1767);
nand U2689 (N_2689,N_1381,N_1520);
or U2690 (N_2690,N_1114,N_1521);
nand U2691 (N_2691,N_1181,N_1139);
nand U2692 (N_2692,N_1886,N_1123);
nor U2693 (N_2693,N_1352,N_1839);
nand U2694 (N_2694,N_1692,N_1705);
or U2695 (N_2695,N_1000,N_1474);
or U2696 (N_2696,N_1721,N_1682);
or U2697 (N_2697,N_1882,N_1450);
and U2698 (N_2698,N_1048,N_1928);
and U2699 (N_2699,N_1743,N_1778);
nor U2700 (N_2700,N_1776,N_1682);
and U2701 (N_2701,N_1241,N_1106);
nor U2702 (N_2702,N_1960,N_1420);
and U2703 (N_2703,N_1792,N_1860);
or U2704 (N_2704,N_1081,N_1750);
nor U2705 (N_2705,N_1076,N_1212);
xor U2706 (N_2706,N_1557,N_1299);
xor U2707 (N_2707,N_1013,N_1526);
or U2708 (N_2708,N_1620,N_1096);
or U2709 (N_2709,N_1066,N_1878);
nor U2710 (N_2710,N_1518,N_1663);
and U2711 (N_2711,N_1742,N_1536);
nor U2712 (N_2712,N_1286,N_1490);
nand U2713 (N_2713,N_1343,N_1216);
nand U2714 (N_2714,N_1659,N_1764);
nor U2715 (N_2715,N_1533,N_1500);
or U2716 (N_2716,N_1791,N_1544);
nand U2717 (N_2717,N_1834,N_1192);
nor U2718 (N_2718,N_1438,N_1067);
nor U2719 (N_2719,N_1774,N_1160);
nor U2720 (N_2720,N_1672,N_1278);
nor U2721 (N_2721,N_1422,N_1328);
and U2722 (N_2722,N_1916,N_1320);
and U2723 (N_2723,N_1399,N_1040);
xor U2724 (N_2724,N_1346,N_1436);
and U2725 (N_2725,N_1610,N_1005);
or U2726 (N_2726,N_1202,N_1902);
nor U2727 (N_2727,N_1718,N_1474);
xnor U2728 (N_2728,N_1347,N_1122);
or U2729 (N_2729,N_1022,N_1643);
xnor U2730 (N_2730,N_1621,N_1772);
xnor U2731 (N_2731,N_1938,N_1664);
xnor U2732 (N_2732,N_1915,N_1382);
and U2733 (N_2733,N_1894,N_1807);
and U2734 (N_2734,N_1914,N_1879);
nor U2735 (N_2735,N_1883,N_1030);
nand U2736 (N_2736,N_1889,N_1296);
nand U2737 (N_2737,N_1122,N_1717);
nor U2738 (N_2738,N_1459,N_1585);
nor U2739 (N_2739,N_1730,N_1932);
xor U2740 (N_2740,N_1620,N_1952);
or U2741 (N_2741,N_1936,N_1310);
or U2742 (N_2742,N_1265,N_1807);
nand U2743 (N_2743,N_1544,N_1998);
nor U2744 (N_2744,N_1877,N_1991);
nor U2745 (N_2745,N_1437,N_1648);
nor U2746 (N_2746,N_1747,N_1210);
or U2747 (N_2747,N_1628,N_1107);
nor U2748 (N_2748,N_1183,N_1468);
nand U2749 (N_2749,N_1147,N_1331);
nand U2750 (N_2750,N_1279,N_1490);
and U2751 (N_2751,N_1045,N_1378);
nand U2752 (N_2752,N_1551,N_1334);
and U2753 (N_2753,N_1147,N_1269);
xor U2754 (N_2754,N_1896,N_1359);
nor U2755 (N_2755,N_1471,N_1537);
and U2756 (N_2756,N_1161,N_1789);
nand U2757 (N_2757,N_1581,N_1400);
nor U2758 (N_2758,N_1714,N_1918);
nor U2759 (N_2759,N_1996,N_1245);
or U2760 (N_2760,N_1883,N_1499);
or U2761 (N_2761,N_1993,N_1184);
nand U2762 (N_2762,N_1843,N_1587);
nor U2763 (N_2763,N_1298,N_1421);
and U2764 (N_2764,N_1374,N_1737);
nor U2765 (N_2765,N_1304,N_1893);
nor U2766 (N_2766,N_1355,N_1710);
and U2767 (N_2767,N_1110,N_1482);
nor U2768 (N_2768,N_1204,N_1881);
nor U2769 (N_2769,N_1123,N_1536);
nand U2770 (N_2770,N_1095,N_1552);
nor U2771 (N_2771,N_1029,N_1749);
or U2772 (N_2772,N_1831,N_1778);
nor U2773 (N_2773,N_1917,N_1156);
nand U2774 (N_2774,N_1740,N_1664);
nand U2775 (N_2775,N_1283,N_1721);
nor U2776 (N_2776,N_1452,N_1369);
and U2777 (N_2777,N_1564,N_1341);
nor U2778 (N_2778,N_1322,N_1171);
nor U2779 (N_2779,N_1733,N_1347);
or U2780 (N_2780,N_1401,N_1407);
nor U2781 (N_2781,N_1629,N_1994);
xnor U2782 (N_2782,N_1504,N_1526);
nand U2783 (N_2783,N_1056,N_1831);
xnor U2784 (N_2784,N_1793,N_1869);
xnor U2785 (N_2785,N_1610,N_1277);
nor U2786 (N_2786,N_1180,N_1237);
nor U2787 (N_2787,N_1750,N_1289);
nor U2788 (N_2788,N_1916,N_1602);
and U2789 (N_2789,N_1908,N_1266);
nand U2790 (N_2790,N_1557,N_1730);
or U2791 (N_2791,N_1444,N_1459);
nor U2792 (N_2792,N_1136,N_1926);
and U2793 (N_2793,N_1433,N_1690);
nand U2794 (N_2794,N_1804,N_1596);
and U2795 (N_2795,N_1469,N_1819);
nand U2796 (N_2796,N_1497,N_1365);
or U2797 (N_2797,N_1243,N_1948);
or U2798 (N_2798,N_1065,N_1284);
nor U2799 (N_2799,N_1755,N_1049);
xor U2800 (N_2800,N_1898,N_1979);
and U2801 (N_2801,N_1055,N_1951);
nand U2802 (N_2802,N_1717,N_1907);
or U2803 (N_2803,N_1966,N_1330);
nor U2804 (N_2804,N_1867,N_1210);
and U2805 (N_2805,N_1651,N_1579);
nand U2806 (N_2806,N_1032,N_1632);
nand U2807 (N_2807,N_1277,N_1171);
or U2808 (N_2808,N_1232,N_1726);
and U2809 (N_2809,N_1020,N_1880);
or U2810 (N_2810,N_1709,N_1063);
and U2811 (N_2811,N_1781,N_1043);
and U2812 (N_2812,N_1603,N_1809);
and U2813 (N_2813,N_1480,N_1172);
or U2814 (N_2814,N_1497,N_1951);
nor U2815 (N_2815,N_1271,N_1172);
nand U2816 (N_2816,N_1632,N_1698);
and U2817 (N_2817,N_1427,N_1519);
and U2818 (N_2818,N_1648,N_1030);
nand U2819 (N_2819,N_1828,N_1166);
nor U2820 (N_2820,N_1443,N_1463);
or U2821 (N_2821,N_1098,N_1049);
nand U2822 (N_2822,N_1983,N_1989);
nand U2823 (N_2823,N_1823,N_1057);
xnor U2824 (N_2824,N_1250,N_1630);
nand U2825 (N_2825,N_1146,N_1909);
nor U2826 (N_2826,N_1148,N_1064);
nor U2827 (N_2827,N_1616,N_1443);
and U2828 (N_2828,N_1410,N_1061);
or U2829 (N_2829,N_1121,N_1833);
or U2830 (N_2830,N_1608,N_1882);
nor U2831 (N_2831,N_1161,N_1625);
and U2832 (N_2832,N_1686,N_1653);
and U2833 (N_2833,N_1581,N_1393);
nor U2834 (N_2834,N_1168,N_1697);
nor U2835 (N_2835,N_1290,N_1128);
or U2836 (N_2836,N_1230,N_1714);
or U2837 (N_2837,N_1301,N_1782);
or U2838 (N_2838,N_1168,N_1755);
or U2839 (N_2839,N_1278,N_1995);
nor U2840 (N_2840,N_1111,N_1808);
xnor U2841 (N_2841,N_1760,N_1383);
nand U2842 (N_2842,N_1132,N_1487);
xnor U2843 (N_2843,N_1325,N_1124);
or U2844 (N_2844,N_1566,N_1932);
xnor U2845 (N_2845,N_1324,N_1539);
and U2846 (N_2846,N_1340,N_1349);
nor U2847 (N_2847,N_1225,N_1585);
and U2848 (N_2848,N_1886,N_1013);
or U2849 (N_2849,N_1219,N_1201);
nor U2850 (N_2850,N_1151,N_1842);
nand U2851 (N_2851,N_1831,N_1341);
or U2852 (N_2852,N_1468,N_1485);
and U2853 (N_2853,N_1045,N_1589);
and U2854 (N_2854,N_1895,N_1947);
nor U2855 (N_2855,N_1375,N_1754);
and U2856 (N_2856,N_1995,N_1848);
nor U2857 (N_2857,N_1620,N_1453);
and U2858 (N_2858,N_1420,N_1247);
nand U2859 (N_2859,N_1903,N_1673);
and U2860 (N_2860,N_1549,N_1026);
xnor U2861 (N_2861,N_1076,N_1279);
or U2862 (N_2862,N_1550,N_1208);
or U2863 (N_2863,N_1004,N_1886);
xnor U2864 (N_2864,N_1852,N_1866);
nand U2865 (N_2865,N_1442,N_1967);
nor U2866 (N_2866,N_1436,N_1210);
or U2867 (N_2867,N_1438,N_1398);
and U2868 (N_2868,N_1094,N_1865);
nor U2869 (N_2869,N_1503,N_1682);
nand U2870 (N_2870,N_1931,N_1364);
and U2871 (N_2871,N_1691,N_1300);
nand U2872 (N_2872,N_1227,N_1219);
nand U2873 (N_2873,N_1527,N_1989);
nor U2874 (N_2874,N_1062,N_1517);
and U2875 (N_2875,N_1156,N_1778);
or U2876 (N_2876,N_1988,N_1806);
and U2877 (N_2877,N_1525,N_1393);
nand U2878 (N_2878,N_1413,N_1451);
nor U2879 (N_2879,N_1283,N_1501);
nand U2880 (N_2880,N_1916,N_1810);
and U2881 (N_2881,N_1873,N_1855);
and U2882 (N_2882,N_1922,N_1486);
xor U2883 (N_2883,N_1888,N_1939);
or U2884 (N_2884,N_1696,N_1919);
and U2885 (N_2885,N_1434,N_1371);
and U2886 (N_2886,N_1839,N_1967);
nand U2887 (N_2887,N_1803,N_1308);
nor U2888 (N_2888,N_1195,N_1118);
nand U2889 (N_2889,N_1918,N_1945);
nand U2890 (N_2890,N_1565,N_1788);
or U2891 (N_2891,N_1195,N_1789);
nand U2892 (N_2892,N_1450,N_1354);
and U2893 (N_2893,N_1244,N_1842);
or U2894 (N_2894,N_1395,N_1525);
nor U2895 (N_2895,N_1189,N_1833);
nor U2896 (N_2896,N_1856,N_1926);
or U2897 (N_2897,N_1928,N_1130);
nor U2898 (N_2898,N_1948,N_1331);
and U2899 (N_2899,N_1732,N_1391);
or U2900 (N_2900,N_1811,N_1510);
or U2901 (N_2901,N_1742,N_1355);
nand U2902 (N_2902,N_1323,N_1102);
and U2903 (N_2903,N_1664,N_1033);
and U2904 (N_2904,N_1409,N_1056);
and U2905 (N_2905,N_1506,N_1681);
nor U2906 (N_2906,N_1047,N_1911);
nand U2907 (N_2907,N_1690,N_1948);
nor U2908 (N_2908,N_1590,N_1918);
xor U2909 (N_2909,N_1708,N_1687);
xnor U2910 (N_2910,N_1162,N_1096);
or U2911 (N_2911,N_1211,N_1063);
nor U2912 (N_2912,N_1154,N_1897);
and U2913 (N_2913,N_1695,N_1372);
and U2914 (N_2914,N_1756,N_1257);
and U2915 (N_2915,N_1697,N_1654);
nand U2916 (N_2916,N_1120,N_1797);
nor U2917 (N_2917,N_1275,N_1360);
nor U2918 (N_2918,N_1335,N_1805);
nand U2919 (N_2919,N_1811,N_1017);
nor U2920 (N_2920,N_1076,N_1245);
nor U2921 (N_2921,N_1203,N_1291);
and U2922 (N_2922,N_1174,N_1572);
nand U2923 (N_2923,N_1314,N_1480);
nand U2924 (N_2924,N_1784,N_1195);
xnor U2925 (N_2925,N_1559,N_1426);
and U2926 (N_2926,N_1578,N_1591);
and U2927 (N_2927,N_1852,N_1453);
xnor U2928 (N_2928,N_1275,N_1071);
and U2929 (N_2929,N_1592,N_1142);
or U2930 (N_2930,N_1455,N_1852);
and U2931 (N_2931,N_1926,N_1757);
or U2932 (N_2932,N_1656,N_1257);
or U2933 (N_2933,N_1510,N_1690);
nor U2934 (N_2934,N_1068,N_1100);
or U2935 (N_2935,N_1370,N_1530);
nand U2936 (N_2936,N_1063,N_1472);
xnor U2937 (N_2937,N_1598,N_1724);
and U2938 (N_2938,N_1655,N_1412);
xnor U2939 (N_2939,N_1162,N_1169);
and U2940 (N_2940,N_1908,N_1600);
nor U2941 (N_2941,N_1293,N_1624);
nor U2942 (N_2942,N_1429,N_1124);
or U2943 (N_2943,N_1100,N_1176);
nor U2944 (N_2944,N_1271,N_1534);
or U2945 (N_2945,N_1274,N_1623);
nand U2946 (N_2946,N_1140,N_1028);
or U2947 (N_2947,N_1041,N_1756);
and U2948 (N_2948,N_1560,N_1924);
and U2949 (N_2949,N_1291,N_1098);
nor U2950 (N_2950,N_1704,N_1543);
xnor U2951 (N_2951,N_1863,N_1383);
and U2952 (N_2952,N_1473,N_1753);
nand U2953 (N_2953,N_1056,N_1413);
nand U2954 (N_2954,N_1171,N_1693);
and U2955 (N_2955,N_1251,N_1666);
nor U2956 (N_2956,N_1395,N_1244);
and U2957 (N_2957,N_1677,N_1138);
xor U2958 (N_2958,N_1335,N_1721);
and U2959 (N_2959,N_1777,N_1152);
nor U2960 (N_2960,N_1482,N_1227);
and U2961 (N_2961,N_1925,N_1108);
and U2962 (N_2962,N_1383,N_1069);
or U2963 (N_2963,N_1739,N_1772);
nand U2964 (N_2964,N_1788,N_1370);
and U2965 (N_2965,N_1975,N_1369);
nor U2966 (N_2966,N_1692,N_1709);
or U2967 (N_2967,N_1070,N_1739);
nand U2968 (N_2968,N_1227,N_1821);
xnor U2969 (N_2969,N_1921,N_1324);
or U2970 (N_2970,N_1803,N_1822);
nor U2971 (N_2971,N_1071,N_1740);
and U2972 (N_2972,N_1728,N_1756);
or U2973 (N_2973,N_1860,N_1468);
and U2974 (N_2974,N_1361,N_1449);
nor U2975 (N_2975,N_1642,N_1086);
nor U2976 (N_2976,N_1898,N_1989);
and U2977 (N_2977,N_1193,N_1693);
nand U2978 (N_2978,N_1837,N_1906);
nor U2979 (N_2979,N_1190,N_1561);
or U2980 (N_2980,N_1669,N_1720);
and U2981 (N_2981,N_1422,N_1145);
nor U2982 (N_2982,N_1475,N_1301);
or U2983 (N_2983,N_1059,N_1189);
nand U2984 (N_2984,N_1375,N_1088);
nand U2985 (N_2985,N_1572,N_1256);
nor U2986 (N_2986,N_1300,N_1910);
nand U2987 (N_2987,N_1729,N_1069);
xor U2988 (N_2988,N_1723,N_1520);
nand U2989 (N_2989,N_1435,N_1820);
or U2990 (N_2990,N_1690,N_1172);
nand U2991 (N_2991,N_1682,N_1161);
nand U2992 (N_2992,N_1715,N_1220);
nor U2993 (N_2993,N_1041,N_1292);
nand U2994 (N_2994,N_1442,N_1644);
and U2995 (N_2995,N_1070,N_1536);
nand U2996 (N_2996,N_1770,N_1702);
or U2997 (N_2997,N_1877,N_1331);
nor U2998 (N_2998,N_1765,N_1523);
and U2999 (N_2999,N_1248,N_1155);
nor U3000 (N_3000,N_2318,N_2235);
or U3001 (N_3001,N_2268,N_2405);
or U3002 (N_3002,N_2526,N_2835);
xor U3003 (N_3003,N_2013,N_2919);
or U3004 (N_3004,N_2733,N_2173);
or U3005 (N_3005,N_2344,N_2059);
and U3006 (N_3006,N_2270,N_2399);
nor U3007 (N_3007,N_2219,N_2794);
and U3008 (N_3008,N_2109,N_2401);
xnor U3009 (N_3009,N_2834,N_2838);
and U3010 (N_3010,N_2700,N_2643);
or U3011 (N_3011,N_2293,N_2549);
nand U3012 (N_3012,N_2687,N_2648);
and U3013 (N_3013,N_2891,N_2029);
nor U3014 (N_3014,N_2617,N_2915);
xor U3015 (N_3015,N_2373,N_2618);
or U3016 (N_3016,N_2679,N_2443);
nand U3017 (N_3017,N_2407,N_2855);
and U3018 (N_3018,N_2005,N_2478);
and U3019 (N_3019,N_2299,N_2563);
or U3020 (N_3020,N_2079,N_2837);
nand U3021 (N_3021,N_2672,N_2368);
nor U3022 (N_3022,N_2767,N_2332);
and U3023 (N_3023,N_2028,N_2553);
or U3024 (N_3024,N_2611,N_2195);
or U3025 (N_3025,N_2513,N_2441);
and U3026 (N_3026,N_2681,N_2211);
nand U3027 (N_3027,N_2761,N_2004);
nand U3028 (N_3028,N_2626,N_2208);
nor U3029 (N_3029,N_2823,N_2938);
nand U3030 (N_3030,N_2587,N_2262);
and U3031 (N_3031,N_2985,N_2036);
or U3032 (N_3032,N_2912,N_2038);
and U3033 (N_3033,N_2755,N_2193);
and U3034 (N_3034,N_2062,N_2190);
nor U3035 (N_3035,N_2762,N_2381);
xor U3036 (N_3036,N_2135,N_2256);
or U3037 (N_3037,N_2530,N_2558);
and U3038 (N_3038,N_2123,N_2666);
and U3039 (N_3039,N_2593,N_2271);
or U3040 (N_3040,N_2683,N_2706);
or U3041 (N_3041,N_2205,N_2947);
and U3042 (N_3042,N_2063,N_2039);
nor U3043 (N_3043,N_2844,N_2157);
xor U3044 (N_3044,N_2186,N_2936);
and U3045 (N_3045,N_2247,N_2360);
and U3046 (N_3046,N_2065,N_2546);
or U3047 (N_3047,N_2636,N_2896);
nor U3048 (N_3048,N_2367,N_2759);
nor U3049 (N_3049,N_2199,N_2291);
and U3050 (N_3050,N_2612,N_2705);
nor U3051 (N_3051,N_2662,N_2459);
or U3052 (N_3052,N_2991,N_2045);
nor U3053 (N_3053,N_2719,N_2596);
and U3054 (N_3054,N_2818,N_2557);
xor U3055 (N_3055,N_2272,N_2006);
nor U3056 (N_3056,N_2020,N_2225);
or U3057 (N_3057,N_2415,N_2795);
nor U3058 (N_3058,N_2171,N_2031);
or U3059 (N_3059,N_2793,N_2099);
and U3060 (N_3060,N_2274,N_2337);
nand U3061 (N_3061,N_2507,N_2601);
nand U3062 (N_3062,N_2926,N_2144);
or U3063 (N_3063,N_2276,N_2866);
and U3064 (N_3064,N_2136,N_2046);
and U3065 (N_3065,N_2543,N_2469);
and U3066 (N_3066,N_2502,N_2750);
nand U3067 (N_3067,N_2942,N_2877);
nor U3068 (N_3068,N_2792,N_2480);
and U3069 (N_3069,N_2817,N_2691);
nand U3070 (N_3070,N_2956,N_2847);
and U3071 (N_3071,N_2773,N_2963);
or U3072 (N_3072,N_2581,N_2331);
and U3073 (N_3073,N_2395,N_2521);
nand U3074 (N_3074,N_2192,N_2467);
nand U3075 (N_3075,N_2808,N_2309);
and U3076 (N_3076,N_2995,N_2377);
and U3077 (N_3077,N_2231,N_2634);
nand U3078 (N_3078,N_2051,N_2204);
nand U3079 (N_3079,N_2210,N_2397);
nand U3080 (N_3080,N_2481,N_2885);
nand U3081 (N_3081,N_2196,N_2898);
nand U3082 (N_3082,N_2983,N_2206);
xor U3083 (N_3083,N_2506,N_2884);
nand U3084 (N_3084,N_2803,N_2172);
nand U3085 (N_3085,N_2385,N_2937);
or U3086 (N_3086,N_2166,N_2584);
nor U3087 (N_3087,N_2684,N_2154);
nor U3088 (N_3088,N_2765,N_2200);
nand U3089 (N_3089,N_2027,N_2899);
nand U3090 (N_3090,N_2236,N_2514);
nand U3091 (N_3091,N_2421,N_2954);
and U3092 (N_3092,N_2809,N_2856);
and U3093 (N_3093,N_2152,N_2722);
nor U3094 (N_3094,N_2378,N_2640);
nor U3095 (N_3095,N_2903,N_2893);
nor U3096 (N_3096,N_2629,N_2741);
nor U3097 (N_3097,N_2873,N_2649);
xnor U3098 (N_3098,N_2836,N_2772);
nand U3099 (N_3099,N_2253,N_2001);
or U3100 (N_3100,N_2708,N_2833);
nand U3101 (N_3101,N_2250,N_2440);
nand U3102 (N_3102,N_2339,N_2685);
and U3103 (N_3103,N_2758,N_2964);
or U3104 (N_3104,N_2140,N_2953);
and U3105 (N_3105,N_2310,N_2570);
nand U3106 (N_3106,N_2333,N_2313);
or U3107 (N_3107,N_2374,N_2744);
or U3108 (N_3108,N_2710,N_2734);
or U3109 (N_3109,N_2449,N_2701);
nor U3110 (N_3110,N_2163,N_2315);
nor U3111 (N_3111,N_2100,N_2160);
nand U3112 (N_3112,N_2107,N_2312);
nor U3113 (N_3113,N_2535,N_2479);
nor U3114 (N_3114,N_2106,N_2165);
nand U3115 (N_3115,N_2286,N_2141);
nand U3116 (N_3116,N_2533,N_2583);
nor U3117 (N_3117,N_2512,N_2913);
nor U3118 (N_3118,N_2879,N_2724);
nand U3119 (N_3119,N_2673,N_2789);
xnor U3120 (N_3120,N_2752,N_2158);
and U3121 (N_3121,N_2801,N_2391);
or U3122 (N_3122,N_2542,N_2962);
nor U3123 (N_3123,N_2328,N_2116);
nor U3124 (N_3124,N_2815,N_2070);
nor U3125 (N_3125,N_2861,N_2967);
or U3126 (N_3126,N_2414,N_2055);
nand U3127 (N_3127,N_2552,N_2468);
and U3128 (N_3128,N_2218,N_2184);
xor U3129 (N_3129,N_2126,N_2698);
nand U3130 (N_3130,N_2134,N_2806);
and U3131 (N_3131,N_2252,N_2343);
nor U3132 (N_3132,N_2580,N_2402);
and U3133 (N_3133,N_2457,N_2941);
or U3134 (N_3134,N_2900,N_2987);
and U3135 (N_3135,N_2153,N_2098);
and U3136 (N_3136,N_2411,N_2091);
nor U3137 (N_3137,N_2349,N_2233);
xor U3138 (N_3138,N_2798,N_2524);
nor U3139 (N_3139,N_2060,N_2639);
xor U3140 (N_3140,N_2745,N_2277);
nor U3141 (N_3141,N_2167,N_2709);
and U3142 (N_3142,N_2010,N_2357);
and U3143 (N_3143,N_2957,N_2671);
and U3144 (N_3144,N_2824,N_2830);
or U3145 (N_3145,N_2655,N_2554);
nor U3146 (N_3146,N_2538,N_2177);
nand U3147 (N_3147,N_2303,N_2927);
nor U3148 (N_3148,N_2675,N_2024);
nor U3149 (N_3149,N_2510,N_2279);
or U3150 (N_3150,N_2960,N_2347);
and U3151 (N_3151,N_2592,N_2696);
nand U3152 (N_3152,N_2260,N_2738);
or U3153 (N_3153,N_2689,N_2973);
and U3154 (N_3154,N_2609,N_2959);
nand U3155 (N_3155,N_2785,N_2370);
and U3156 (N_3156,N_2069,N_2658);
nor U3157 (N_3157,N_2298,N_2019);
or U3158 (N_3158,N_2693,N_2909);
nand U3159 (N_3159,N_2826,N_2409);
nor U3160 (N_3160,N_2198,N_2245);
nor U3161 (N_3161,N_2610,N_2930);
and U3162 (N_3162,N_2041,N_2472);
or U3163 (N_3163,N_2372,N_2654);
xnor U3164 (N_3164,N_2018,N_2283);
nand U3165 (N_3165,N_2131,N_2577);
and U3166 (N_3166,N_2676,N_2450);
nand U3167 (N_3167,N_2493,N_2661);
xnor U3168 (N_3168,N_2324,N_2904);
nand U3169 (N_3169,N_2138,N_2076);
nor U3170 (N_3170,N_2788,N_2735);
or U3171 (N_3171,N_2585,N_2846);
or U3172 (N_3172,N_2918,N_2489);
nand U3173 (N_3173,N_2682,N_2485);
nor U3174 (N_3174,N_2952,N_2820);
or U3175 (N_3175,N_2061,N_2223);
nand U3176 (N_3176,N_2525,N_2068);
nand U3177 (N_3177,N_2226,N_2294);
or U3178 (N_3178,N_2108,N_2518);
nor U3179 (N_3179,N_2338,N_2308);
or U3180 (N_3180,N_2089,N_2375);
or U3181 (N_3181,N_2032,N_2999);
nand U3182 (N_3182,N_2088,N_2764);
nor U3183 (N_3183,N_2790,N_2384);
nor U3184 (N_3184,N_2768,N_2541);
nand U3185 (N_3185,N_2906,N_2908);
nand U3186 (N_3186,N_2970,N_2497);
and U3187 (N_3187,N_2931,N_2151);
nor U3188 (N_3188,N_2561,N_2354);
and U3189 (N_3189,N_2121,N_2905);
or U3190 (N_3190,N_2828,N_2620);
and U3191 (N_3191,N_2008,N_2389);
or U3192 (N_3192,N_2113,N_2244);
and U3193 (N_3193,N_2117,N_2189);
or U3194 (N_3194,N_2376,N_2255);
nand U3195 (N_3195,N_2087,N_2132);
and U3196 (N_3196,N_2979,N_2142);
or U3197 (N_3197,N_2215,N_2130);
nand U3198 (N_3198,N_2437,N_2499);
and U3199 (N_3199,N_2394,N_2011);
or U3200 (N_3200,N_2660,N_2473);
nand U3201 (N_3201,N_2695,N_2417);
and U3202 (N_3202,N_2760,N_2320);
nor U3203 (N_3203,N_2984,N_2180);
nor U3204 (N_3204,N_2848,N_2564);
and U3205 (N_3205,N_2799,N_2605);
nand U3206 (N_3206,N_2924,N_2392);
nand U3207 (N_3207,N_2652,N_2319);
and U3208 (N_3208,N_2646,N_2476);
nor U3209 (N_3209,N_2273,N_2495);
and U3210 (N_3210,N_2653,N_2874);
nor U3211 (N_3211,N_2081,N_2150);
nand U3212 (N_3212,N_2348,N_2656);
nor U3213 (N_3213,N_2014,N_2015);
xnor U3214 (N_3214,N_2872,N_2509);
and U3215 (N_3215,N_2757,N_2878);
nand U3216 (N_3216,N_2842,N_2241);
or U3217 (N_3217,N_2560,N_2458);
xor U3218 (N_3218,N_2446,N_2914);
xnor U3219 (N_3219,N_2739,N_2935);
nor U3220 (N_3220,N_2187,N_2078);
nor U3221 (N_3221,N_2390,N_2017);
or U3222 (N_3222,N_2329,N_2582);
nand U3223 (N_3223,N_2539,N_2085);
nand U3224 (N_3224,N_2383,N_2220);
nor U3225 (N_3225,N_2197,N_2625);
and U3226 (N_3226,N_2148,N_2229);
or U3227 (N_3227,N_2571,N_2831);
and U3228 (N_3228,N_2246,N_2240);
xor U3229 (N_3229,N_2920,N_2556);
and U3230 (N_3230,N_2282,N_2254);
or U3231 (N_3231,N_2295,N_2025);
nor U3232 (N_3232,N_2145,N_2454);
nor U3233 (N_3233,N_2731,N_2183);
xnor U3234 (N_3234,N_2438,N_2517);
nand U3235 (N_3235,N_2222,N_2621);
nand U3236 (N_3236,N_2090,N_2104);
nand U3237 (N_3237,N_2551,N_2224);
or U3238 (N_3238,N_2988,N_2297);
nor U3239 (N_3239,N_2071,N_2317);
nor U3240 (N_3240,N_2659,N_2083);
or U3241 (N_3241,N_2398,N_2736);
nand U3242 (N_3242,N_2528,N_2420);
nor U3243 (N_3243,N_2769,N_2989);
nor U3244 (N_3244,N_2465,N_2112);
and U3245 (N_3245,N_2729,N_2712);
or U3246 (N_3246,N_2613,N_2436);
or U3247 (N_3247,N_2804,N_2287);
nand U3248 (N_3248,N_2737,N_2812);
and U3249 (N_3249,N_2619,N_2021);
or U3250 (N_3250,N_2054,N_2704);
nor U3251 (N_3251,N_2779,N_2118);
nand U3252 (N_3252,N_2248,N_2505);
or U3253 (N_3253,N_2249,N_2406);
nor U3254 (N_3254,N_2865,N_2470);
nand U3255 (N_3255,N_2500,N_2822);
nor U3256 (N_3256,N_2336,N_2690);
and U3257 (N_3257,N_2072,N_2651);
or U3258 (N_3258,N_2448,N_2486);
and U3259 (N_3259,N_2968,N_2547);
and U3260 (N_3260,N_2868,N_2670);
nand U3261 (N_3261,N_2600,N_2721);
nor U3262 (N_3262,N_2864,N_2545);
or U3263 (N_3263,N_2717,N_2867);
nor U3264 (N_3264,N_2889,N_2092);
or U3265 (N_3265,N_2771,N_2902);
and U3266 (N_3266,N_2049,N_2307);
and U3267 (N_3267,N_2544,N_2125);
or U3268 (N_3268,N_2124,N_2194);
xnor U3269 (N_3269,N_2699,N_2916);
or U3270 (N_3270,N_2413,N_2579);
and U3271 (N_3271,N_2396,N_2519);
nand U3272 (N_3272,N_2404,N_2713);
nor U3273 (N_3273,N_2678,N_2057);
nand U3274 (N_3274,N_2520,N_2073);
and U3275 (N_3275,N_2716,N_2992);
nand U3276 (N_3276,N_2943,N_2212);
nand U3277 (N_3277,N_2565,N_2674);
or U3278 (N_3278,N_2453,N_2201);
nor U3279 (N_3279,N_2400,N_2917);
or U3280 (N_3280,N_2251,N_2669);
nor U3281 (N_3281,N_2423,N_2426);
nand U3282 (N_3282,N_2503,N_2645);
or U3283 (N_3283,N_2977,N_2527);
and U3284 (N_3284,N_2482,N_2425);
and U3285 (N_3285,N_2529,N_2275);
and U3286 (N_3286,N_2657,N_2504);
and U3287 (N_3287,N_2037,N_2944);
nor U3288 (N_3288,N_2576,N_2326);
or U3289 (N_3289,N_2345,N_2149);
nor U3290 (N_3290,N_2366,N_2133);
nor U3291 (N_3291,N_2723,N_2778);
nand U3292 (N_3292,N_2362,N_2209);
and U3293 (N_3293,N_2747,N_2536);
nor U3294 (N_3294,N_2463,N_2179);
nand U3295 (N_3295,N_2464,N_2311);
nand U3296 (N_3296,N_2939,N_2958);
nand U3297 (N_3297,N_2776,N_2483);
and U3298 (N_3298,N_2568,N_2976);
and U3299 (N_3299,N_2614,N_2644);
and U3300 (N_3300,N_2883,N_2860);
and U3301 (N_3301,N_2093,N_2825);
or U3302 (N_3302,N_2791,N_2955);
nor U3303 (N_3303,N_2146,N_2050);
nor U3304 (N_3304,N_2047,N_2484);
nand U3305 (N_3305,N_2921,N_2002);
xor U3306 (N_3306,N_2466,N_2647);
nand U3307 (N_3307,N_2796,N_2129);
nor U3308 (N_3308,N_2871,N_2355);
nand U3309 (N_3309,N_2429,N_2269);
nand U3310 (N_3310,N_2603,N_2058);
and U3311 (N_3311,N_2292,N_2053);
xnor U3312 (N_3312,N_2170,N_2604);
nand U3313 (N_3313,N_2933,N_2756);
xor U3314 (N_3314,N_2892,N_2016);
nand U3315 (N_3315,N_2586,N_2819);
nand U3316 (N_3316,N_2314,N_2774);
nand U3317 (N_3317,N_2780,N_2574);
nand U3318 (N_3318,N_2534,N_2128);
and U3319 (N_3319,N_2492,N_2665);
and U3320 (N_3320,N_2439,N_2559);
xnor U3321 (N_3321,N_2487,N_2289);
or U3322 (N_3322,N_2531,N_2353);
or U3323 (N_3323,N_2412,N_2923);
nor U3324 (N_3324,N_2501,N_2259);
or U3325 (N_3325,N_2548,N_2278);
nor U3326 (N_3326,N_2843,N_2934);
nor U3327 (N_3327,N_2870,N_2203);
nand U3328 (N_3328,N_2410,N_2932);
and U3329 (N_3329,N_2816,N_2688);
or U3330 (N_3330,N_2718,N_2802);
or U3331 (N_3331,N_2114,N_2386);
and U3332 (N_3332,N_2418,N_2839);
nand U3333 (N_3333,N_2607,N_2147);
xnor U3334 (N_3334,N_2237,N_2875);
nand U3335 (N_3335,N_2230,N_2922);
nand U3336 (N_3336,N_2965,N_2052);
or U3337 (N_3337,N_2981,N_2630);
xnor U3338 (N_3338,N_2257,N_2234);
or U3339 (N_3339,N_2280,N_2886);
and U3340 (N_3340,N_2650,N_2990);
nor U3341 (N_3341,N_2101,N_2615);
nor U3342 (N_3342,N_2003,N_2035);
xor U3343 (N_3343,N_2267,N_2740);
and U3344 (N_3344,N_2832,N_2907);
nor U3345 (N_3345,N_2813,N_2416);
or U3346 (N_3346,N_2216,N_2007);
xnor U3347 (N_3347,N_2242,N_2228);
xor U3348 (N_3348,N_2895,N_2595);
or U3349 (N_3349,N_2388,N_2022);
nor U3350 (N_3350,N_2588,N_2598);
nor U3351 (N_3351,N_2911,N_2445);
and U3352 (N_3352,N_2746,N_2854);
and U3353 (N_3353,N_2232,N_2176);
and U3354 (N_3354,N_2940,N_2048);
and U3355 (N_3355,N_2522,N_2996);
and U3356 (N_3356,N_2261,N_2365);
or U3357 (N_3357,N_2703,N_2602);
or U3358 (N_3358,N_2350,N_2403);
and U3359 (N_3359,N_2361,N_2300);
or U3360 (N_3360,N_2488,N_2325);
or U3361 (N_3361,N_2508,N_2714);
and U3362 (N_3362,N_2633,N_2082);
and U3363 (N_3363,N_2097,N_2387);
nor U3364 (N_3364,N_2606,N_2890);
or U3365 (N_3365,N_2296,N_2238);
or U3366 (N_3366,N_2711,N_2221);
nand U3367 (N_3367,N_2102,N_2692);
or U3368 (N_3368,N_2663,N_2040);
nor U3369 (N_3369,N_2857,N_2686);
xor U3370 (N_3370,N_2498,N_2821);
nand U3371 (N_3371,N_2707,N_2239);
nand U3372 (N_3372,N_2202,N_2888);
nand U3373 (N_3373,N_2178,N_2335);
and U3374 (N_3374,N_2641,N_2869);
xor U3375 (N_3375,N_2858,N_2998);
nor U3376 (N_3376,N_2382,N_2105);
or U3377 (N_3377,N_2573,N_2523);
nand U3378 (N_3378,N_2110,N_2188);
and U3379 (N_3379,N_2444,N_2726);
and U3380 (N_3380,N_2594,N_2800);
nand U3381 (N_3381,N_2862,N_2422);
or U3382 (N_3382,N_2997,N_2243);
nor U3383 (N_3383,N_2447,N_2624);
xnor U3384 (N_3384,N_2622,N_2599);
or U3385 (N_3385,N_2972,N_2782);
nand U3386 (N_3386,N_2763,N_2080);
or U3387 (N_3387,N_2550,N_2213);
and U3388 (N_3388,N_2638,N_2748);
xor U3389 (N_3389,N_2590,N_2887);
nand U3390 (N_3390,N_2264,N_2702);
nor U3391 (N_3391,N_2316,N_2359);
xor U3392 (N_3392,N_2000,N_2496);
nand U3393 (N_3393,N_2342,N_2863);
or U3394 (N_3394,N_2288,N_2460);
and U3395 (N_3395,N_2428,N_2540);
nor U3396 (N_3396,N_2258,N_2949);
nor U3397 (N_3397,N_2728,N_2227);
nand U3398 (N_3398,N_2969,N_2012);
xnor U3399 (N_3399,N_2516,N_2044);
nor U3400 (N_3400,N_2845,N_2424);
and U3401 (N_3401,N_2978,N_2491);
xnor U3402 (N_3402,N_2191,N_2475);
nor U3403 (N_3403,N_2352,N_2302);
and U3404 (N_3404,N_2364,N_2589);
nand U3405 (N_3405,N_2948,N_2119);
or U3406 (N_3406,N_2009,N_2853);
or U3407 (N_3407,N_2026,N_2537);
and U3408 (N_3408,N_2749,N_2929);
nor U3409 (N_3409,N_2066,N_2694);
nor U3410 (N_3410,N_2980,N_2217);
nand U3411 (N_3411,N_2034,N_2074);
or U3412 (N_3412,N_2578,N_2301);
nor U3413 (N_3413,N_2419,N_2628);
nand U3414 (N_3414,N_2456,N_2322);
xor U3415 (N_3415,N_2371,N_2174);
nand U3416 (N_3416,N_2304,N_2966);
nor U3417 (N_3417,N_2851,N_2515);
or U3418 (N_3418,N_2994,N_2043);
nand U3419 (N_3419,N_2042,N_2623);
nor U3420 (N_3420,N_2430,N_2770);
nor U3421 (N_3421,N_2829,N_2814);
and U3422 (N_3422,N_2993,N_2122);
and U3423 (N_3423,N_2169,N_2901);
or U3424 (N_3424,N_2797,N_2265);
nand U3425 (N_3425,N_2910,N_2642);
xnor U3426 (N_3426,N_2408,N_2321);
nor U3427 (N_3427,N_2637,N_2358);
nor U3428 (N_3428,N_2777,N_2067);
nor U3429 (N_3429,N_2143,N_2766);
nor U3430 (N_3430,N_2435,N_2185);
nor U3431 (N_3431,N_2667,N_2876);
nor U3432 (N_3432,N_2668,N_2452);
and U3433 (N_3433,N_2427,N_2743);
or U3434 (N_3434,N_2442,N_2787);
nor U3435 (N_3435,N_2334,N_2103);
and U3436 (N_3436,N_2356,N_2168);
and U3437 (N_3437,N_2207,N_2285);
or U3438 (N_3438,N_2471,N_2164);
nor U3439 (N_3439,N_2086,N_2961);
nor U3440 (N_3440,N_2751,N_2075);
nor U3441 (N_3441,N_2730,N_2882);
xnor U3442 (N_3442,N_2971,N_2379);
nand U3443 (N_3443,N_2975,N_2290);
nand U3444 (N_3444,N_2462,N_2330);
or U3445 (N_3445,N_2635,N_2850);
and U3446 (N_3446,N_2680,N_2754);
and U3447 (N_3447,N_2175,N_2811);
nand U3448 (N_3448,N_2786,N_2742);
and U3449 (N_3449,N_2461,N_2030);
nand U3450 (N_3450,N_2162,N_2137);
nand U3451 (N_3451,N_2827,N_2572);
nand U3452 (N_3452,N_2715,N_2139);
nand U3453 (N_3453,N_2341,N_2511);
nor U3454 (N_3454,N_2182,N_2455);
and U3455 (N_3455,N_2120,N_2096);
or U3456 (N_3456,N_2982,N_2664);
and U3457 (N_3457,N_2897,N_2323);
nand U3458 (N_3458,N_2451,N_2608);
or U3459 (N_3459,N_2346,N_2783);
xnor U3460 (N_3460,N_2950,N_2266);
and U3461 (N_3461,N_2477,N_2095);
nor U3462 (N_3462,N_2064,N_2281);
and U3463 (N_3463,N_2807,N_2805);
nand U3464 (N_3464,N_2474,N_2566);
xnor U3465 (N_3465,N_2111,N_2894);
and U3466 (N_3466,N_2156,N_2161);
nor U3467 (N_3467,N_2363,N_2023);
nand U3468 (N_3468,N_2775,N_2155);
and U3469 (N_3469,N_2115,N_2627);
and U3470 (N_3470,N_2562,N_2084);
and U3471 (N_3471,N_2306,N_2431);
and U3472 (N_3472,N_2263,N_2434);
and U3473 (N_3473,N_2532,N_2946);
or U3474 (N_3474,N_2880,N_2725);
nand U3475 (N_3475,N_2951,N_2784);
or U3476 (N_3476,N_2631,N_2569);
nand U3477 (N_3477,N_2928,N_2351);
and U3478 (N_3478,N_2077,N_2327);
or U3479 (N_3479,N_2810,N_2986);
and U3480 (N_3480,N_2945,N_2974);
nor U3481 (N_3481,N_2033,N_2727);
and U3482 (N_3482,N_2567,N_2432);
or U3483 (N_3483,N_2616,N_2591);
xnor U3484 (N_3484,N_2433,N_2632);
nand U3485 (N_3485,N_2849,N_2881);
or U3486 (N_3486,N_2284,N_2340);
and U3487 (N_3487,N_2555,N_2859);
and U3488 (N_3488,N_2305,N_2597);
and U3489 (N_3489,N_2127,N_2575);
nor U3490 (N_3490,N_2380,N_2393);
or U3491 (N_3491,N_2494,N_2214);
or U3492 (N_3492,N_2490,N_2840);
nor U3493 (N_3493,N_2094,N_2841);
nand U3494 (N_3494,N_2781,N_2732);
and U3495 (N_3495,N_2056,N_2720);
nand U3496 (N_3496,N_2677,N_2852);
xor U3497 (N_3497,N_2697,N_2369);
nand U3498 (N_3498,N_2159,N_2181);
and U3499 (N_3499,N_2925,N_2753);
or U3500 (N_3500,N_2267,N_2036);
nor U3501 (N_3501,N_2886,N_2783);
and U3502 (N_3502,N_2106,N_2525);
nand U3503 (N_3503,N_2165,N_2412);
xor U3504 (N_3504,N_2918,N_2001);
or U3505 (N_3505,N_2057,N_2599);
and U3506 (N_3506,N_2010,N_2001);
and U3507 (N_3507,N_2241,N_2285);
nand U3508 (N_3508,N_2644,N_2162);
nor U3509 (N_3509,N_2742,N_2598);
or U3510 (N_3510,N_2676,N_2932);
and U3511 (N_3511,N_2154,N_2360);
nand U3512 (N_3512,N_2450,N_2521);
nand U3513 (N_3513,N_2495,N_2652);
nor U3514 (N_3514,N_2260,N_2120);
or U3515 (N_3515,N_2459,N_2002);
xnor U3516 (N_3516,N_2208,N_2232);
or U3517 (N_3517,N_2304,N_2700);
or U3518 (N_3518,N_2801,N_2732);
nand U3519 (N_3519,N_2101,N_2885);
xnor U3520 (N_3520,N_2610,N_2896);
nand U3521 (N_3521,N_2103,N_2862);
xnor U3522 (N_3522,N_2423,N_2193);
or U3523 (N_3523,N_2489,N_2140);
and U3524 (N_3524,N_2935,N_2823);
and U3525 (N_3525,N_2975,N_2343);
or U3526 (N_3526,N_2426,N_2608);
nand U3527 (N_3527,N_2089,N_2714);
nor U3528 (N_3528,N_2070,N_2332);
nand U3529 (N_3529,N_2148,N_2547);
or U3530 (N_3530,N_2455,N_2107);
nor U3531 (N_3531,N_2827,N_2845);
or U3532 (N_3532,N_2828,N_2139);
xnor U3533 (N_3533,N_2675,N_2268);
xor U3534 (N_3534,N_2954,N_2482);
or U3535 (N_3535,N_2633,N_2311);
xor U3536 (N_3536,N_2513,N_2733);
nor U3537 (N_3537,N_2652,N_2799);
nor U3538 (N_3538,N_2872,N_2966);
nor U3539 (N_3539,N_2335,N_2217);
or U3540 (N_3540,N_2373,N_2001);
nand U3541 (N_3541,N_2958,N_2743);
nand U3542 (N_3542,N_2230,N_2943);
xnor U3543 (N_3543,N_2861,N_2222);
nand U3544 (N_3544,N_2687,N_2012);
nor U3545 (N_3545,N_2453,N_2777);
nor U3546 (N_3546,N_2839,N_2876);
nand U3547 (N_3547,N_2265,N_2795);
xor U3548 (N_3548,N_2620,N_2771);
nand U3549 (N_3549,N_2256,N_2106);
nor U3550 (N_3550,N_2750,N_2964);
and U3551 (N_3551,N_2016,N_2947);
and U3552 (N_3552,N_2514,N_2534);
or U3553 (N_3553,N_2298,N_2395);
or U3554 (N_3554,N_2466,N_2239);
nor U3555 (N_3555,N_2213,N_2765);
or U3556 (N_3556,N_2837,N_2796);
or U3557 (N_3557,N_2353,N_2516);
and U3558 (N_3558,N_2437,N_2143);
nor U3559 (N_3559,N_2285,N_2399);
nor U3560 (N_3560,N_2465,N_2959);
nor U3561 (N_3561,N_2192,N_2766);
nand U3562 (N_3562,N_2985,N_2563);
nand U3563 (N_3563,N_2297,N_2593);
nand U3564 (N_3564,N_2303,N_2525);
nor U3565 (N_3565,N_2656,N_2502);
xnor U3566 (N_3566,N_2020,N_2053);
nor U3567 (N_3567,N_2587,N_2386);
nand U3568 (N_3568,N_2682,N_2814);
and U3569 (N_3569,N_2057,N_2768);
or U3570 (N_3570,N_2998,N_2267);
nor U3571 (N_3571,N_2822,N_2583);
nor U3572 (N_3572,N_2973,N_2353);
nand U3573 (N_3573,N_2622,N_2652);
and U3574 (N_3574,N_2889,N_2759);
and U3575 (N_3575,N_2525,N_2543);
xor U3576 (N_3576,N_2934,N_2689);
nor U3577 (N_3577,N_2231,N_2196);
nor U3578 (N_3578,N_2936,N_2716);
nand U3579 (N_3579,N_2524,N_2101);
and U3580 (N_3580,N_2283,N_2430);
xnor U3581 (N_3581,N_2287,N_2760);
nand U3582 (N_3582,N_2875,N_2094);
and U3583 (N_3583,N_2913,N_2418);
nand U3584 (N_3584,N_2694,N_2087);
or U3585 (N_3585,N_2065,N_2148);
or U3586 (N_3586,N_2113,N_2777);
nand U3587 (N_3587,N_2755,N_2044);
or U3588 (N_3588,N_2091,N_2121);
and U3589 (N_3589,N_2104,N_2083);
or U3590 (N_3590,N_2023,N_2514);
nand U3591 (N_3591,N_2020,N_2979);
and U3592 (N_3592,N_2291,N_2309);
nor U3593 (N_3593,N_2258,N_2927);
and U3594 (N_3594,N_2014,N_2299);
or U3595 (N_3595,N_2118,N_2512);
nand U3596 (N_3596,N_2410,N_2537);
nor U3597 (N_3597,N_2543,N_2850);
or U3598 (N_3598,N_2804,N_2087);
xnor U3599 (N_3599,N_2367,N_2575);
nor U3600 (N_3600,N_2661,N_2949);
nand U3601 (N_3601,N_2665,N_2977);
nand U3602 (N_3602,N_2481,N_2137);
nand U3603 (N_3603,N_2347,N_2962);
nand U3604 (N_3604,N_2037,N_2973);
nor U3605 (N_3605,N_2148,N_2131);
nor U3606 (N_3606,N_2331,N_2758);
and U3607 (N_3607,N_2110,N_2515);
nand U3608 (N_3608,N_2142,N_2597);
and U3609 (N_3609,N_2847,N_2708);
nand U3610 (N_3610,N_2521,N_2490);
and U3611 (N_3611,N_2422,N_2648);
or U3612 (N_3612,N_2382,N_2754);
and U3613 (N_3613,N_2051,N_2284);
xor U3614 (N_3614,N_2835,N_2047);
nand U3615 (N_3615,N_2490,N_2121);
nand U3616 (N_3616,N_2211,N_2720);
nand U3617 (N_3617,N_2683,N_2565);
nor U3618 (N_3618,N_2203,N_2003);
and U3619 (N_3619,N_2952,N_2948);
or U3620 (N_3620,N_2948,N_2522);
and U3621 (N_3621,N_2079,N_2959);
nand U3622 (N_3622,N_2403,N_2479);
or U3623 (N_3623,N_2520,N_2863);
nor U3624 (N_3624,N_2923,N_2549);
xnor U3625 (N_3625,N_2943,N_2726);
or U3626 (N_3626,N_2331,N_2536);
or U3627 (N_3627,N_2850,N_2706);
or U3628 (N_3628,N_2100,N_2731);
nor U3629 (N_3629,N_2382,N_2653);
nor U3630 (N_3630,N_2998,N_2017);
xnor U3631 (N_3631,N_2408,N_2704);
nand U3632 (N_3632,N_2242,N_2609);
nand U3633 (N_3633,N_2446,N_2013);
or U3634 (N_3634,N_2324,N_2191);
nand U3635 (N_3635,N_2045,N_2169);
and U3636 (N_3636,N_2888,N_2240);
and U3637 (N_3637,N_2319,N_2664);
or U3638 (N_3638,N_2119,N_2241);
or U3639 (N_3639,N_2730,N_2923);
nor U3640 (N_3640,N_2475,N_2701);
and U3641 (N_3641,N_2449,N_2729);
and U3642 (N_3642,N_2527,N_2815);
nor U3643 (N_3643,N_2726,N_2647);
or U3644 (N_3644,N_2995,N_2559);
xnor U3645 (N_3645,N_2738,N_2204);
xor U3646 (N_3646,N_2127,N_2825);
nor U3647 (N_3647,N_2015,N_2745);
nand U3648 (N_3648,N_2502,N_2031);
or U3649 (N_3649,N_2563,N_2913);
xnor U3650 (N_3650,N_2175,N_2087);
nand U3651 (N_3651,N_2597,N_2313);
nand U3652 (N_3652,N_2641,N_2940);
or U3653 (N_3653,N_2130,N_2207);
and U3654 (N_3654,N_2976,N_2695);
or U3655 (N_3655,N_2779,N_2570);
nor U3656 (N_3656,N_2482,N_2436);
and U3657 (N_3657,N_2419,N_2997);
nand U3658 (N_3658,N_2875,N_2886);
xnor U3659 (N_3659,N_2320,N_2801);
xnor U3660 (N_3660,N_2708,N_2921);
and U3661 (N_3661,N_2668,N_2152);
or U3662 (N_3662,N_2102,N_2449);
nand U3663 (N_3663,N_2869,N_2497);
xor U3664 (N_3664,N_2657,N_2107);
nor U3665 (N_3665,N_2203,N_2077);
or U3666 (N_3666,N_2587,N_2192);
and U3667 (N_3667,N_2469,N_2161);
nor U3668 (N_3668,N_2013,N_2663);
or U3669 (N_3669,N_2825,N_2461);
or U3670 (N_3670,N_2879,N_2365);
or U3671 (N_3671,N_2737,N_2576);
nand U3672 (N_3672,N_2897,N_2192);
and U3673 (N_3673,N_2145,N_2953);
xnor U3674 (N_3674,N_2891,N_2605);
or U3675 (N_3675,N_2035,N_2273);
or U3676 (N_3676,N_2775,N_2171);
xnor U3677 (N_3677,N_2307,N_2105);
nand U3678 (N_3678,N_2557,N_2463);
nor U3679 (N_3679,N_2581,N_2412);
and U3680 (N_3680,N_2128,N_2855);
or U3681 (N_3681,N_2722,N_2286);
and U3682 (N_3682,N_2184,N_2476);
and U3683 (N_3683,N_2719,N_2874);
or U3684 (N_3684,N_2977,N_2080);
nor U3685 (N_3685,N_2047,N_2697);
xnor U3686 (N_3686,N_2262,N_2667);
or U3687 (N_3687,N_2549,N_2487);
nand U3688 (N_3688,N_2291,N_2264);
nand U3689 (N_3689,N_2021,N_2047);
and U3690 (N_3690,N_2822,N_2716);
xnor U3691 (N_3691,N_2910,N_2817);
and U3692 (N_3692,N_2927,N_2513);
nand U3693 (N_3693,N_2517,N_2228);
or U3694 (N_3694,N_2353,N_2731);
or U3695 (N_3695,N_2841,N_2972);
nor U3696 (N_3696,N_2350,N_2683);
nand U3697 (N_3697,N_2096,N_2494);
or U3698 (N_3698,N_2585,N_2649);
nand U3699 (N_3699,N_2072,N_2212);
xnor U3700 (N_3700,N_2160,N_2485);
and U3701 (N_3701,N_2508,N_2270);
nand U3702 (N_3702,N_2021,N_2768);
and U3703 (N_3703,N_2422,N_2319);
and U3704 (N_3704,N_2149,N_2721);
xor U3705 (N_3705,N_2224,N_2777);
nand U3706 (N_3706,N_2923,N_2764);
or U3707 (N_3707,N_2617,N_2967);
nand U3708 (N_3708,N_2447,N_2313);
nor U3709 (N_3709,N_2445,N_2092);
and U3710 (N_3710,N_2863,N_2502);
nand U3711 (N_3711,N_2314,N_2969);
and U3712 (N_3712,N_2804,N_2604);
xnor U3713 (N_3713,N_2018,N_2193);
nand U3714 (N_3714,N_2601,N_2810);
nor U3715 (N_3715,N_2598,N_2185);
nor U3716 (N_3716,N_2257,N_2405);
nor U3717 (N_3717,N_2185,N_2750);
and U3718 (N_3718,N_2059,N_2218);
or U3719 (N_3719,N_2893,N_2475);
and U3720 (N_3720,N_2421,N_2713);
nand U3721 (N_3721,N_2810,N_2204);
nor U3722 (N_3722,N_2849,N_2328);
and U3723 (N_3723,N_2398,N_2486);
xnor U3724 (N_3724,N_2594,N_2795);
nor U3725 (N_3725,N_2937,N_2230);
and U3726 (N_3726,N_2514,N_2332);
nand U3727 (N_3727,N_2212,N_2153);
nor U3728 (N_3728,N_2320,N_2845);
and U3729 (N_3729,N_2871,N_2830);
nand U3730 (N_3730,N_2495,N_2615);
xor U3731 (N_3731,N_2689,N_2266);
and U3732 (N_3732,N_2427,N_2023);
nor U3733 (N_3733,N_2525,N_2474);
nor U3734 (N_3734,N_2938,N_2615);
nand U3735 (N_3735,N_2267,N_2890);
nand U3736 (N_3736,N_2105,N_2609);
nor U3737 (N_3737,N_2092,N_2935);
nor U3738 (N_3738,N_2588,N_2498);
nand U3739 (N_3739,N_2654,N_2637);
nand U3740 (N_3740,N_2974,N_2543);
nand U3741 (N_3741,N_2707,N_2182);
nor U3742 (N_3742,N_2828,N_2829);
xor U3743 (N_3743,N_2925,N_2018);
nor U3744 (N_3744,N_2238,N_2808);
and U3745 (N_3745,N_2514,N_2590);
nor U3746 (N_3746,N_2782,N_2519);
or U3747 (N_3747,N_2128,N_2331);
nor U3748 (N_3748,N_2901,N_2344);
xor U3749 (N_3749,N_2382,N_2717);
nor U3750 (N_3750,N_2386,N_2663);
nor U3751 (N_3751,N_2931,N_2348);
nand U3752 (N_3752,N_2739,N_2856);
and U3753 (N_3753,N_2750,N_2857);
and U3754 (N_3754,N_2849,N_2432);
xor U3755 (N_3755,N_2748,N_2974);
nor U3756 (N_3756,N_2664,N_2816);
and U3757 (N_3757,N_2261,N_2166);
and U3758 (N_3758,N_2912,N_2145);
nor U3759 (N_3759,N_2657,N_2065);
nand U3760 (N_3760,N_2863,N_2802);
nand U3761 (N_3761,N_2716,N_2072);
and U3762 (N_3762,N_2282,N_2955);
nand U3763 (N_3763,N_2306,N_2829);
nor U3764 (N_3764,N_2075,N_2470);
nand U3765 (N_3765,N_2432,N_2771);
or U3766 (N_3766,N_2754,N_2851);
nand U3767 (N_3767,N_2133,N_2498);
or U3768 (N_3768,N_2443,N_2113);
nand U3769 (N_3769,N_2703,N_2357);
nor U3770 (N_3770,N_2313,N_2031);
nor U3771 (N_3771,N_2759,N_2839);
nand U3772 (N_3772,N_2770,N_2922);
and U3773 (N_3773,N_2659,N_2195);
or U3774 (N_3774,N_2381,N_2729);
xor U3775 (N_3775,N_2021,N_2357);
or U3776 (N_3776,N_2829,N_2922);
nand U3777 (N_3777,N_2639,N_2597);
nor U3778 (N_3778,N_2287,N_2031);
or U3779 (N_3779,N_2102,N_2178);
or U3780 (N_3780,N_2098,N_2607);
nor U3781 (N_3781,N_2828,N_2459);
and U3782 (N_3782,N_2876,N_2850);
and U3783 (N_3783,N_2276,N_2634);
nand U3784 (N_3784,N_2192,N_2431);
xnor U3785 (N_3785,N_2197,N_2517);
nor U3786 (N_3786,N_2770,N_2283);
xor U3787 (N_3787,N_2780,N_2312);
nor U3788 (N_3788,N_2337,N_2159);
nor U3789 (N_3789,N_2915,N_2905);
or U3790 (N_3790,N_2363,N_2139);
xor U3791 (N_3791,N_2539,N_2577);
or U3792 (N_3792,N_2489,N_2226);
nand U3793 (N_3793,N_2544,N_2303);
xnor U3794 (N_3794,N_2678,N_2782);
nand U3795 (N_3795,N_2260,N_2431);
and U3796 (N_3796,N_2263,N_2791);
nor U3797 (N_3797,N_2497,N_2950);
or U3798 (N_3798,N_2379,N_2927);
and U3799 (N_3799,N_2541,N_2669);
xnor U3800 (N_3800,N_2531,N_2971);
nor U3801 (N_3801,N_2398,N_2315);
nor U3802 (N_3802,N_2093,N_2436);
or U3803 (N_3803,N_2053,N_2576);
nor U3804 (N_3804,N_2722,N_2982);
nor U3805 (N_3805,N_2392,N_2513);
or U3806 (N_3806,N_2503,N_2192);
or U3807 (N_3807,N_2005,N_2521);
or U3808 (N_3808,N_2125,N_2456);
and U3809 (N_3809,N_2809,N_2973);
nor U3810 (N_3810,N_2459,N_2676);
nor U3811 (N_3811,N_2507,N_2810);
nand U3812 (N_3812,N_2996,N_2102);
nand U3813 (N_3813,N_2023,N_2128);
xnor U3814 (N_3814,N_2824,N_2530);
and U3815 (N_3815,N_2871,N_2327);
and U3816 (N_3816,N_2970,N_2603);
nand U3817 (N_3817,N_2516,N_2077);
nor U3818 (N_3818,N_2261,N_2965);
nand U3819 (N_3819,N_2173,N_2863);
and U3820 (N_3820,N_2397,N_2544);
or U3821 (N_3821,N_2407,N_2754);
and U3822 (N_3822,N_2122,N_2897);
and U3823 (N_3823,N_2565,N_2573);
nor U3824 (N_3824,N_2535,N_2402);
xor U3825 (N_3825,N_2930,N_2762);
nand U3826 (N_3826,N_2083,N_2751);
or U3827 (N_3827,N_2418,N_2187);
nand U3828 (N_3828,N_2020,N_2446);
nor U3829 (N_3829,N_2299,N_2490);
and U3830 (N_3830,N_2823,N_2890);
nor U3831 (N_3831,N_2722,N_2701);
xnor U3832 (N_3832,N_2579,N_2522);
xor U3833 (N_3833,N_2619,N_2822);
or U3834 (N_3834,N_2134,N_2266);
nand U3835 (N_3835,N_2000,N_2656);
and U3836 (N_3836,N_2099,N_2528);
and U3837 (N_3837,N_2936,N_2650);
nand U3838 (N_3838,N_2279,N_2673);
or U3839 (N_3839,N_2136,N_2383);
nand U3840 (N_3840,N_2622,N_2026);
and U3841 (N_3841,N_2059,N_2419);
nor U3842 (N_3842,N_2807,N_2591);
or U3843 (N_3843,N_2739,N_2374);
or U3844 (N_3844,N_2876,N_2924);
and U3845 (N_3845,N_2151,N_2578);
or U3846 (N_3846,N_2740,N_2469);
nor U3847 (N_3847,N_2827,N_2025);
nand U3848 (N_3848,N_2400,N_2445);
and U3849 (N_3849,N_2316,N_2858);
or U3850 (N_3850,N_2084,N_2186);
nand U3851 (N_3851,N_2923,N_2146);
xnor U3852 (N_3852,N_2050,N_2699);
or U3853 (N_3853,N_2065,N_2681);
and U3854 (N_3854,N_2929,N_2932);
or U3855 (N_3855,N_2192,N_2539);
and U3856 (N_3856,N_2201,N_2864);
nand U3857 (N_3857,N_2221,N_2527);
and U3858 (N_3858,N_2968,N_2987);
and U3859 (N_3859,N_2080,N_2666);
nor U3860 (N_3860,N_2276,N_2397);
nor U3861 (N_3861,N_2373,N_2581);
xor U3862 (N_3862,N_2048,N_2594);
xnor U3863 (N_3863,N_2779,N_2073);
and U3864 (N_3864,N_2566,N_2282);
or U3865 (N_3865,N_2861,N_2242);
or U3866 (N_3866,N_2761,N_2445);
nor U3867 (N_3867,N_2136,N_2115);
nand U3868 (N_3868,N_2878,N_2597);
or U3869 (N_3869,N_2453,N_2830);
or U3870 (N_3870,N_2887,N_2048);
nand U3871 (N_3871,N_2072,N_2885);
or U3872 (N_3872,N_2321,N_2068);
nand U3873 (N_3873,N_2033,N_2621);
or U3874 (N_3874,N_2114,N_2128);
and U3875 (N_3875,N_2836,N_2159);
or U3876 (N_3876,N_2201,N_2649);
nand U3877 (N_3877,N_2767,N_2323);
or U3878 (N_3878,N_2292,N_2281);
or U3879 (N_3879,N_2690,N_2711);
xor U3880 (N_3880,N_2799,N_2987);
or U3881 (N_3881,N_2611,N_2567);
and U3882 (N_3882,N_2351,N_2404);
or U3883 (N_3883,N_2453,N_2310);
nand U3884 (N_3884,N_2145,N_2457);
nand U3885 (N_3885,N_2544,N_2914);
nand U3886 (N_3886,N_2305,N_2411);
or U3887 (N_3887,N_2687,N_2934);
nand U3888 (N_3888,N_2574,N_2178);
nor U3889 (N_3889,N_2290,N_2600);
or U3890 (N_3890,N_2598,N_2932);
nand U3891 (N_3891,N_2651,N_2573);
or U3892 (N_3892,N_2349,N_2635);
nor U3893 (N_3893,N_2860,N_2772);
nand U3894 (N_3894,N_2414,N_2145);
or U3895 (N_3895,N_2953,N_2344);
nand U3896 (N_3896,N_2370,N_2479);
nand U3897 (N_3897,N_2617,N_2279);
xnor U3898 (N_3898,N_2751,N_2328);
nand U3899 (N_3899,N_2975,N_2350);
nand U3900 (N_3900,N_2663,N_2828);
xor U3901 (N_3901,N_2697,N_2657);
nor U3902 (N_3902,N_2052,N_2685);
or U3903 (N_3903,N_2946,N_2344);
and U3904 (N_3904,N_2289,N_2461);
nand U3905 (N_3905,N_2385,N_2332);
xnor U3906 (N_3906,N_2372,N_2368);
nor U3907 (N_3907,N_2505,N_2279);
and U3908 (N_3908,N_2688,N_2457);
nor U3909 (N_3909,N_2500,N_2749);
and U3910 (N_3910,N_2815,N_2868);
and U3911 (N_3911,N_2531,N_2077);
and U3912 (N_3912,N_2153,N_2952);
or U3913 (N_3913,N_2943,N_2069);
and U3914 (N_3914,N_2850,N_2152);
nor U3915 (N_3915,N_2778,N_2904);
nand U3916 (N_3916,N_2724,N_2656);
nand U3917 (N_3917,N_2479,N_2660);
and U3918 (N_3918,N_2394,N_2998);
nand U3919 (N_3919,N_2716,N_2566);
xor U3920 (N_3920,N_2004,N_2484);
nand U3921 (N_3921,N_2892,N_2568);
nor U3922 (N_3922,N_2562,N_2060);
or U3923 (N_3923,N_2984,N_2350);
and U3924 (N_3924,N_2274,N_2858);
or U3925 (N_3925,N_2600,N_2160);
and U3926 (N_3926,N_2050,N_2127);
nor U3927 (N_3927,N_2112,N_2410);
and U3928 (N_3928,N_2995,N_2213);
nand U3929 (N_3929,N_2612,N_2445);
xnor U3930 (N_3930,N_2811,N_2374);
or U3931 (N_3931,N_2798,N_2964);
or U3932 (N_3932,N_2367,N_2334);
or U3933 (N_3933,N_2523,N_2582);
and U3934 (N_3934,N_2767,N_2787);
and U3935 (N_3935,N_2743,N_2970);
and U3936 (N_3936,N_2498,N_2251);
nand U3937 (N_3937,N_2009,N_2182);
nor U3938 (N_3938,N_2665,N_2042);
or U3939 (N_3939,N_2172,N_2794);
or U3940 (N_3940,N_2397,N_2054);
or U3941 (N_3941,N_2339,N_2436);
nor U3942 (N_3942,N_2827,N_2655);
and U3943 (N_3943,N_2540,N_2769);
or U3944 (N_3944,N_2888,N_2326);
nor U3945 (N_3945,N_2989,N_2839);
nor U3946 (N_3946,N_2677,N_2138);
nor U3947 (N_3947,N_2986,N_2252);
nand U3948 (N_3948,N_2843,N_2256);
nand U3949 (N_3949,N_2499,N_2605);
or U3950 (N_3950,N_2415,N_2625);
or U3951 (N_3951,N_2693,N_2993);
or U3952 (N_3952,N_2714,N_2532);
nor U3953 (N_3953,N_2328,N_2838);
xnor U3954 (N_3954,N_2717,N_2668);
and U3955 (N_3955,N_2114,N_2011);
and U3956 (N_3956,N_2689,N_2695);
or U3957 (N_3957,N_2650,N_2136);
or U3958 (N_3958,N_2346,N_2654);
and U3959 (N_3959,N_2802,N_2125);
and U3960 (N_3960,N_2170,N_2667);
nor U3961 (N_3961,N_2369,N_2211);
and U3962 (N_3962,N_2855,N_2283);
or U3963 (N_3963,N_2417,N_2963);
and U3964 (N_3964,N_2685,N_2675);
nor U3965 (N_3965,N_2057,N_2780);
or U3966 (N_3966,N_2724,N_2561);
nor U3967 (N_3967,N_2736,N_2930);
xor U3968 (N_3968,N_2208,N_2263);
and U3969 (N_3969,N_2321,N_2712);
and U3970 (N_3970,N_2033,N_2225);
nand U3971 (N_3971,N_2665,N_2065);
or U3972 (N_3972,N_2011,N_2273);
and U3973 (N_3973,N_2576,N_2137);
and U3974 (N_3974,N_2459,N_2610);
nand U3975 (N_3975,N_2420,N_2195);
nand U3976 (N_3976,N_2768,N_2604);
nand U3977 (N_3977,N_2612,N_2830);
nor U3978 (N_3978,N_2399,N_2133);
nor U3979 (N_3979,N_2127,N_2778);
nand U3980 (N_3980,N_2418,N_2386);
and U3981 (N_3981,N_2729,N_2866);
and U3982 (N_3982,N_2996,N_2712);
nand U3983 (N_3983,N_2553,N_2099);
or U3984 (N_3984,N_2280,N_2763);
nand U3985 (N_3985,N_2523,N_2983);
xnor U3986 (N_3986,N_2296,N_2040);
or U3987 (N_3987,N_2498,N_2414);
nor U3988 (N_3988,N_2454,N_2198);
and U3989 (N_3989,N_2512,N_2478);
or U3990 (N_3990,N_2086,N_2617);
nand U3991 (N_3991,N_2701,N_2597);
nor U3992 (N_3992,N_2499,N_2281);
or U3993 (N_3993,N_2987,N_2432);
and U3994 (N_3994,N_2220,N_2990);
and U3995 (N_3995,N_2737,N_2512);
xor U3996 (N_3996,N_2265,N_2608);
or U3997 (N_3997,N_2786,N_2518);
nand U3998 (N_3998,N_2614,N_2862);
and U3999 (N_3999,N_2210,N_2448);
nand U4000 (N_4000,N_3981,N_3342);
and U4001 (N_4001,N_3601,N_3063);
nor U4002 (N_4002,N_3686,N_3123);
or U4003 (N_4003,N_3191,N_3006);
nor U4004 (N_4004,N_3577,N_3495);
xnor U4005 (N_4005,N_3345,N_3631);
and U4006 (N_4006,N_3931,N_3125);
xor U4007 (N_4007,N_3825,N_3453);
and U4008 (N_4008,N_3782,N_3022);
and U4009 (N_4009,N_3179,N_3751);
nand U4010 (N_4010,N_3481,N_3851);
and U4011 (N_4011,N_3662,N_3441);
or U4012 (N_4012,N_3062,N_3479);
nand U4013 (N_4013,N_3461,N_3578);
nor U4014 (N_4014,N_3564,N_3717);
nand U4015 (N_4015,N_3771,N_3472);
or U4016 (N_4016,N_3701,N_3480);
nor U4017 (N_4017,N_3474,N_3672);
nor U4018 (N_4018,N_3285,N_3003);
nand U4019 (N_4019,N_3962,N_3895);
nor U4020 (N_4020,N_3834,N_3463);
nand U4021 (N_4021,N_3746,N_3506);
and U4022 (N_4022,N_3133,N_3198);
and U4023 (N_4023,N_3560,N_3685);
nor U4024 (N_4024,N_3024,N_3335);
nand U4025 (N_4025,N_3183,N_3148);
or U4026 (N_4026,N_3060,N_3162);
nand U4027 (N_4027,N_3720,N_3272);
nand U4028 (N_4028,N_3443,N_3009);
nor U4029 (N_4029,N_3399,N_3315);
and U4030 (N_4030,N_3450,N_3501);
nand U4031 (N_4031,N_3802,N_3901);
or U4032 (N_4032,N_3670,N_3846);
and U4033 (N_4033,N_3914,N_3558);
and U4034 (N_4034,N_3974,N_3423);
nor U4035 (N_4035,N_3530,N_3204);
nor U4036 (N_4036,N_3543,N_3805);
nor U4037 (N_4037,N_3169,N_3777);
or U4038 (N_4038,N_3677,N_3597);
and U4039 (N_4039,N_3076,N_3185);
or U4040 (N_4040,N_3697,N_3986);
nor U4041 (N_4041,N_3823,N_3683);
nor U4042 (N_4042,N_3862,N_3572);
nand U4043 (N_4043,N_3794,N_3235);
nand U4044 (N_4044,N_3816,N_3300);
or U4045 (N_4045,N_3039,N_3291);
and U4046 (N_4046,N_3769,N_3099);
nand U4047 (N_4047,N_3694,N_3987);
or U4048 (N_4048,N_3668,N_3080);
nor U4049 (N_4049,N_3562,N_3404);
and U4050 (N_4050,N_3579,N_3739);
nor U4051 (N_4051,N_3553,N_3407);
and U4052 (N_4052,N_3565,N_3468);
xor U4053 (N_4053,N_3596,N_3294);
and U4054 (N_4054,N_3083,N_3330);
xor U4055 (N_4055,N_3354,N_3103);
and U4056 (N_4056,N_3155,N_3585);
nand U4057 (N_4057,N_3071,N_3264);
nor U4058 (N_4058,N_3001,N_3841);
xnor U4059 (N_4059,N_3602,N_3245);
or U4060 (N_4060,N_3640,N_3035);
or U4061 (N_4061,N_3700,N_3610);
or U4062 (N_4062,N_3532,N_3112);
nor U4063 (N_4063,N_3554,N_3483);
xor U4064 (N_4064,N_3611,N_3533);
nand U4065 (N_4065,N_3184,N_3403);
or U4066 (N_4066,N_3867,N_3475);
nor U4067 (N_4067,N_3556,N_3695);
nor U4068 (N_4068,N_3084,N_3326);
nor U4069 (N_4069,N_3809,N_3959);
nor U4070 (N_4070,N_3352,N_3621);
nand U4071 (N_4071,N_3870,N_3837);
or U4072 (N_4072,N_3722,N_3815);
nand U4073 (N_4073,N_3958,N_3369);
nor U4074 (N_4074,N_3612,N_3160);
or U4075 (N_4075,N_3641,N_3220);
and U4076 (N_4076,N_3225,N_3535);
and U4077 (N_4077,N_3803,N_3885);
nand U4078 (N_4078,N_3027,N_3218);
nor U4079 (N_4079,N_3066,N_3905);
or U4080 (N_4080,N_3550,N_3969);
xnor U4081 (N_4081,N_3744,N_3977);
nor U4082 (N_4082,N_3241,N_3053);
xnor U4083 (N_4083,N_3889,N_3161);
or U4084 (N_4084,N_3199,N_3154);
nor U4085 (N_4085,N_3051,N_3521);
and U4086 (N_4086,N_3380,N_3435);
and U4087 (N_4087,N_3041,N_3627);
nor U4088 (N_4088,N_3747,N_3261);
nand U4089 (N_4089,N_3849,N_3568);
nor U4090 (N_4090,N_3709,N_3401);
and U4091 (N_4091,N_3473,N_3582);
xor U4092 (N_4092,N_3632,N_3364);
and U4093 (N_4093,N_3788,N_3279);
nand U4094 (N_4094,N_3793,N_3304);
or U4095 (N_4095,N_3433,N_3046);
nand U4096 (N_4096,N_3933,N_3016);
nand U4097 (N_4097,N_3363,N_3265);
or U4098 (N_4098,N_3386,N_3351);
and U4099 (N_4099,N_3190,N_3116);
xor U4100 (N_4100,N_3703,N_3504);
or U4101 (N_4101,N_3749,N_3766);
xor U4102 (N_4102,N_3015,N_3379);
nand U4103 (N_4103,N_3947,N_3079);
nand U4104 (N_4104,N_3661,N_3415);
and U4105 (N_4105,N_3107,N_3850);
nor U4106 (N_4106,N_3201,N_3678);
or U4107 (N_4107,N_3249,N_3238);
and U4108 (N_4108,N_3252,N_3708);
and U4109 (N_4109,N_3286,N_3312);
and U4110 (N_4110,N_3761,N_3874);
or U4111 (N_4111,N_3340,N_3247);
nor U4112 (N_4112,N_3037,N_3078);
and U4113 (N_4113,N_3875,N_3324);
and U4114 (N_4114,N_3406,N_3244);
nand U4115 (N_4115,N_3628,N_3956);
xnor U4116 (N_4116,N_3911,N_3593);
nor U4117 (N_4117,N_3555,N_3350);
and U4118 (N_4118,N_3365,N_3783);
xnor U4119 (N_4119,N_3492,N_3652);
or U4120 (N_4120,N_3548,N_3438);
xnor U4121 (N_4121,N_3892,N_3127);
and U4122 (N_4122,N_3036,N_3390);
or U4123 (N_4123,N_3411,N_3657);
or U4124 (N_4124,N_3493,N_3859);
nand U4125 (N_4125,N_3773,N_3471);
xor U4126 (N_4126,N_3392,N_3424);
or U4127 (N_4127,N_3636,N_3897);
nand U4128 (N_4128,N_3242,N_3417);
or U4129 (N_4129,N_3882,N_3835);
nand U4130 (N_4130,N_3707,N_3604);
or U4131 (N_4131,N_3362,N_3546);
nor U4132 (N_4132,N_3608,N_3687);
nand U4133 (N_4133,N_3868,N_3985);
nor U4134 (N_4134,N_3736,N_3638);
or U4135 (N_4135,N_3693,N_3821);
and U4136 (N_4136,N_3216,N_3332);
or U4137 (N_4137,N_3302,N_3781);
xnor U4138 (N_4138,N_3129,N_3826);
and U4139 (N_4139,N_3587,N_3305);
nand U4140 (N_4140,N_3861,N_3254);
nand U4141 (N_4141,N_3188,N_3716);
nand U4142 (N_4142,N_3538,N_3325);
nand U4143 (N_4143,N_3926,N_3192);
or U4144 (N_4144,N_3757,N_3624);
nand U4145 (N_4145,N_3671,N_3289);
or U4146 (N_4146,N_3232,N_3356);
and U4147 (N_4147,N_3923,N_3669);
nor U4148 (N_4148,N_3951,N_3055);
nand U4149 (N_4149,N_3786,N_3131);
and U4150 (N_4150,N_3371,N_3159);
nor U4151 (N_4151,N_3203,N_3303);
or U4152 (N_4152,N_3136,N_3113);
nand U4153 (N_4153,N_3385,N_3446);
and U4154 (N_4154,N_3246,N_3712);
nand U4155 (N_4155,N_3663,N_3007);
or U4156 (N_4156,N_3275,N_3347);
xor U4157 (N_4157,N_3607,N_3567);
nand U4158 (N_4158,N_3765,N_3944);
nand U4159 (N_4159,N_3266,N_3134);
nor U4160 (N_4160,N_3348,N_3137);
or U4161 (N_4161,N_3319,N_3282);
and U4162 (N_4162,N_3792,N_3171);
nand U4163 (N_4163,N_3298,N_3964);
nor U4164 (N_4164,N_3988,N_3732);
nor U4165 (N_4165,N_3963,N_3400);
or U4166 (N_4166,N_3519,N_3370);
or U4167 (N_4167,N_3509,N_3353);
and U4168 (N_4168,N_3308,N_3045);
xor U4169 (N_4169,N_3092,N_3307);
nand U4170 (N_4170,N_3421,N_3373);
xnor U4171 (N_4171,N_3320,N_3284);
nor U4172 (N_4172,N_3948,N_3108);
nor U4173 (N_4173,N_3212,N_3357);
nor U4174 (N_4174,N_3735,N_3605);
nand U4175 (N_4175,N_3237,N_3994);
or U4176 (N_4176,N_3594,N_3660);
xor U4177 (N_4177,N_3698,N_3295);
xor U4178 (N_4178,N_3946,N_3524);
and U4179 (N_4179,N_3102,N_3647);
and U4180 (N_4180,N_3917,N_3551);
nand U4181 (N_4181,N_3410,N_3454);
nor U4182 (N_4182,N_3448,N_3854);
and U4183 (N_4183,N_3710,N_3955);
and U4184 (N_4184,N_3592,N_3281);
and U4185 (N_4185,N_3419,N_3997);
nor U4186 (N_4186,N_3910,N_3081);
and U4187 (N_4187,N_3681,N_3827);
or U4188 (N_4188,N_3496,N_3017);
and U4189 (N_4189,N_3654,N_3459);
nor U4190 (N_4190,N_3590,N_3393);
nand U4191 (N_4191,N_3916,N_3609);
nor U4192 (N_4192,N_3919,N_3173);
xor U4193 (N_4193,N_3070,N_3737);
nor U4194 (N_4194,N_3230,N_3488);
nor U4195 (N_4195,N_3114,N_3341);
nor U4196 (N_4196,N_3526,N_3848);
or U4197 (N_4197,N_3240,N_3452);
or U4198 (N_4198,N_3011,N_3513);
nand U4199 (N_4199,N_3752,N_3855);
and U4200 (N_4200,N_3359,N_3429);
nand U4201 (N_4201,N_3738,N_3598);
or U4202 (N_4202,N_3925,N_3500);
or U4203 (N_4203,N_3844,N_3518);
and U4204 (N_4204,N_3048,N_3489);
and U4205 (N_4205,N_3288,N_3887);
nand U4206 (N_4206,N_3117,N_3121);
and U4207 (N_4207,N_3135,N_3536);
and U4208 (N_4208,N_3915,N_3293);
xnor U4209 (N_4209,N_3756,N_3360);
nor U4210 (N_4210,N_3091,N_3589);
nor U4211 (N_4211,N_3702,N_3516);
or U4212 (N_4212,N_3269,N_3845);
or U4213 (N_4213,N_3750,N_3615);
nor U4214 (N_4214,N_3881,N_3759);
or U4215 (N_4215,N_3434,N_3089);
and U4216 (N_4216,N_3329,N_3718);
nor U4217 (N_4217,N_3510,N_3943);
nand U4218 (N_4218,N_3623,N_3058);
nand U4219 (N_4219,N_3436,N_3745);
nor U4220 (N_4220,N_3234,N_3780);
nor U4221 (N_4221,N_3023,N_3648);
or U4222 (N_4222,N_3599,N_3912);
nand U4223 (N_4223,N_3402,N_3633);
nor U4224 (N_4224,N_3020,N_3896);
nand U4225 (N_4225,N_3142,N_3290);
xnor U4226 (N_4226,N_3233,N_3096);
and U4227 (N_4227,N_3065,N_3539);
or U4228 (N_4228,N_3511,N_3208);
nand U4229 (N_4229,N_3995,N_3832);
nor U4230 (N_4230,N_3748,N_3398);
or U4231 (N_4231,N_3965,N_3328);
and U4232 (N_4232,N_3343,N_3984);
nor U4233 (N_4233,N_3138,N_3649);
and U4234 (N_4234,N_3960,N_3658);
and U4235 (N_4235,N_3673,N_3166);
nand U4236 (N_4236,N_3014,N_3879);
nor U4237 (N_4237,N_3545,N_3991);
xor U4238 (N_4238,N_3779,N_3213);
or U4239 (N_4239,N_3177,N_3692);
nand U4240 (N_4240,N_3646,N_3833);
xnor U4241 (N_4241,N_3077,N_3067);
and U4242 (N_4242,N_3182,N_3175);
nand U4243 (N_4243,N_3082,N_3153);
and U4244 (N_4244,N_3442,N_3059);
or U4245 (N_4245,N_3257,N_3571);
or U4246 (N_4246,N_3529,N_3574);
nor U4247 (N_4247,N_3296,N_3032);
nand U4248 (N_4248,N_3278,N_3156);
xnor U4249 (N_4249,N_3405,N_3822);
xnor U4250 (N_4250,N_3789,N_3418);
and U4251 (N_4251,N_3219,N_3730);
and U4252 (N_4252,N_3666,N_3907);
and U4253 (N_4253,N_3097,N_3445);
nand U4254 (N_4254,N_3499,N_3795);
nor U4255 (N_4255,N_3828,N_3634);
or U4256 (N_4256,N_3346,N_3491);
and U4257 (N_4257,N_3618,N_3705);
xnor U4258 (N_4258,N_3796,N_3540);
nor U4259 (N_4259,N_3549,N_3000);
and U4260 (N_4260,N_3742,N_3439);
and U4261 (N_4261,N_3228,N_3455);
nand U4262 (N_4262,N_3484,N_3741);
or U4263 (N_4263,N_3952,N_3872);
nand U4264 (N_4264,N_3975,N_3763);
nand U4265 (N_4265,N_3149,N_3635);
nor U4266 (N_4266,N_3193,N_3819);
nor U4267 (N_4267,N_3922,N_3999);
nand U4268 (N_4268,N_3522,N_3258);
and U4269 (N_4269,N_3384,N_3679);
xnor U4270 (N_4270,N_3073,N_3903);
nor U4271 (N_4271,N_3561,N_3165);
nand U4272 (N_4272,N_3818,N_3432);
nand U4273 (N_4273,N_3557,N_3993);
nor U4274 (N_4274,N_3449,N_3010);
and U4275 (N_4275,N_3675,N_3918);
or U4276 (N_4276,N_3144,N_3021);
nor U4277 (N_4277,N_3909,N_3843);
and U4278 (N_4278,N_3847,N_3018);
or U4279 (N_4279,N_3791,N_3200);
nand U4280 (N_4280,N_3239,N_3387);
nand U4281 (N_4281,N_3194,N_3790);
nor U4282 (N_4282,N_3259,N_3236);
and U4283 (N_4283,N_3938,N_3170);
or U4284 (N_4284,N_3391,N_3978);
or U4285 (N_4285,N_3727,N_3580);
nor U4286 (N_4286,N_3031,N_3211);
or U4287 (N_4287,N_3711,N_3689);
nand U4288 (N_4288,N_3110,N_3665);
nor U4289 (N_4289,N_3316,N_3470);
nor U4290 (N_4290,N_3603,N_3101);
and U4291 (N_4291,N_3189,N_3214);
and U4292 (N_4292,N_3105,N_3936);
nand U4293 (N_4293,N_3824,N_3520);
nand U4294 (N_4294,N_3209,N_3318);
and U4295 (N_4295,N_3935,N_3715);
or U4296 (N_4296,N_3243,N_3957);
or U4297 (N_4297,N_3902,N_3575);
nand U4298 (N_4298,N_3327,N_3075);
xor U4299 (N_4299,N_3684,N_3622);
and U4300 (N_4300,N_3762,N_3880);
nor U4301 (N_4301,N_3842,N_3478);
nor U4302 (N_4302,N_3195,N_3667);
or U4303 (N_4303,N_3231,N_3613);
nor U4304 (N_4304,N_3940,N_3460);
nor U4305 (N_4305,N_3893,N_3966);
or U4306 (N_4306,N_3967,N_3772);
or U4307 (N_4307,N_3262,N_3462);
nor U4308 (N_4308,N_3857,N_3811);
nand U4309 (N_4309,N_3950,N_3040);
nand U4310 (N_4310,N_3871,N_3124);
and U4311 (N_4311,N_3397,N_3799);
or U4312 (N_4312,N_3458,N_3215);
nor U4313 (N_4313,N_3584,N_3486);
nor U4314 (N_4314,N_3682,N_3542);
nor U4315 (N_4315,N_3074,N_3038);
nand U4316 (N_4316,N_3726,N_3990);
xor U4317 (N_4317,N_3770,N_3147);
nor U4318 (N_4318,N_3992,N_3853);
xnor U4319 (N_4319,N_3674,N_3313);
or U4320 (N_4320,N_3619,N_3637);
nor U4321 (N_4321,N_3268,N_3900);
xnor U4322 (N_4322,N_3840,N_3644);
and U4323 (N_4323,N_3659,N_3425);
or U4324 (N_4324,N_3552,N_3664);
nor U4325 (N_4325,N_3476,N_3507);
or U4326 (N_4326,N_3733,N_3864);
nor U4327 (N_4327,N_3932,N_3734);
xor U4328 (N_4328,N_3143,N_3381);
nand U4329 (N_4329,N_3547,N_3466);
or U4330 (N_4330,N_3447,N_3140);
or U4331 (N_4331,N_3378,N_3383);
or U4332 (N_4332,N_3287,N_3388);
nand U4333 (N_4333,N_3515,N_3178);
or U4334 (N_4334,N_3115,N_3104);
or U4335 (N_4335,N_3030,N_3382);
and U4336 (N_4336,N_3093,N_3753);
or U4337 (N_4337,N_3299,N_3980);
nor U4338 (N_4338,N_3569,N_3427);
nor U4339 (N_4339,N_3202,N_3052);
nor U4340 (N_4340,N_3814,N_3050);
and U4341 (N_4341,N_3517,N_3339);
or U4342 (N_4342,N_3525,N_3422);
nand U4343 (N_4343,N_3998,N_3251);
and U4344 (N_4344,N_3883,N_3810);
nor U4345 (N_4345,N_3534,N_3187);
or U4346 (N_4346,N_3804,N_3323);
nor U4347 (N_4347,N_3801,N_3976);
or U4348 (N_4348,N_3586,N_3145);
nor U4349 (N_4349,N_3120,N_3537);
and U4350 (N_4350,N_3953,N_3205);
nor U4351 (N_4351,N_3004,N_3366);
nor U4352 (N_4352,N_3512,N_3273);
and U4353 (N_4353,N_3642,N_3152);
nor U4354 (N_4354,N_3563,N_3146);
or U4355 (N_4355,N_3111,N_3409);
nand U4356 (N_4356,N_3186,N_3614);
xnor U4357 (N_4357,N_3581,N_3729);
or U4358 (N_4358,N_3798,N_3248);
nor U4359 (N_4359,N_3349,N_3497);
or U4360 (N_4360,N_3724,N_3263);
nor U4361 (N_4361,N_3576,N_3355);
nand U4362 (N_4362,N_3157,N_3412);
nor U4363 (N_4363,N_3508,N_3921);
xor U4364 (N_4364,N_3150,N_3122);
nand U4365 (N_4365,N_3878,N_3069);
nor U4366 (N_4366,N_3856,N_3128);
nand U4367 (N_4367,N_3416,N_3968);
nor U4368 (N_4368,N_3767,N_3820);
or U4369 (N_4369,N_3168,N_3260);
and U4370 (N_4370,N_3222,N_3595);
nor U4371 (N_4371,N_3884,N_3297);
nand U4372 (N_4372,N_3095,N_3485);
nand U4373 (N_4373,N_3860,N_3514);
nand U4374 (N_4374,N_3172,N_3942);
and U4375 (N_4375,N_3930,N_3368);
or U4376 (N_4376,N_3088,N_3064);
or U4377 (N_4377,N_3056,N_3311);
nor U4378 (N_4378,N_3151,N_3954);
and U4379 (N_4379,N_3817,N_3072);
and U4380 (N_4380,N_3639,N_3087);
nor U4381 (N_4381,N_3440,N_3106);
and U4382 (N_4382,N_3784,N_3270);
nor U4383 (N_4383,N_3728,N_3797);
or U4384 (N_4384,N_3620,N_3743);
nand U4385 (N_4385,N_3713,N_3033);
and U4386 (N_4386,N_3283,N_3982);
or U4387 (N_4387,N_3026,N_3566);
nor U4388 (N_4388,N_3688,N_3929);
or U4389 (N_4389,N_3502,N_3334);
and U4390 (N_4390,N_3431,N_3731);
or U4391 (N_4391,N_3706,N_3367);
nor U4392 (N_4392,N_3787,N_3505);
nand U4393 (N_4393,N_3629,N_3886);
nand U4394 (N_4394,N_3467,N_3898);
or U4395 (N_4395,N_3464,N_3655);
and U4396 (N_4396,N_3650,N_3498);
nor U4397 (N_4397,N_3336,N_3869);
nor U4398 (N_4398,N_3894,N_3049);
and U4399 (N_4399,N_3544,N_3100);
and U4400 (N_4400,N_3180,N_3250);
and U4401 (N_4401,N_3028,N_3785);
and U4402 (N_4402,N_3126,N_3972);
and U4403 (N_4403,N_3426,N_3061);
nor U4404 (N_4404,N_3863,N_3754);
nand U4405 (N_4405,N_3600,N_3939);
nand U4406 (N_4406,N_3776,N_3457);
or U4407 (N_4407,N_3482,N_3331);
and U4408 (N_4408,N_3292,N_3904);
or U4409 (N_4409,N_3428,N_3344);
nor U4410 (N_4410,N_3420,N_3768);
nor U4411 (N_4411,N_3704,N_3255);
nor U4412 (N_4412,N_3691,N_3755);
or U4413 (N_4413,N_3043,N_3338);
and U4414 (N_4414,N_3276,N_3934);
nor U4415 (N_4415,N_3877,N_3888);
nor U4416 (N_4416,N_3927,N_3034);
nand U4417 (N_4417,N_3838,N_3174);
nand U4418 (N_4418,N_3314,N_3839);
or U4419 (N_4419,N_3807,N_3306);
nand U4420 (N_4420,N_3503,N_3164);
or U4421 (N_4421,N_3858,N_3337);
and U4422 (N_4422,N_3490,N_3760);
xor U4423 (N_4423,N_3696,N_3395);
nand U4424 (N_4424,N_3414,N_3451);
nand U4425 (N_4425,N_3961,N_3865);
nor U4426 (N_4426,N_3836,N_3158);
and U4427 (N_4427,N_3812,N_3197);
or U4428 (N_4428,N_3098,N_3224);
xnor U4429 (N_4429,N_3487,N_3394);
nand U4430 (N_4430,N_3430,N_3477);
nand U4431 (N_4431,N_3680,N_3651);
nand U4432 (N_4432,N_3937,N_3876);
xnor U4433 (N_4433,N_3196,N_3831);
nor U4434 (N_4434,N_3800,N_3778);
and U4435 (N_4435,N_3274,N_3676);
or U4436 (N_4436,N_3808,N_3042);
or U4437 (N_4437,N_3906,N_3899);
nand U4438 (N_4438,N_3389,N_3210);
or U4439 (N_4439,N_3139,N_3758);
and U4440 (N_4440,N_3090,N_3973);
nand U4441 (N_4441,N_3979,N_3583);
xnor U4442 (N_4442,N_3047,N_3253);
xor U4443 (N_4443,N_3333,N_3573);
or U4444 (N_4444,N_3372,N_3830);
and U4445 (N_4445,N_3813,N_3890);
nor U4446 (N_4446,N_3852,N_3223);
nor U4447 (N_4447,N_3068,N_3456);
nand U4448 (N_4448,N_3630,N_3920);
or U4449 (N_4449,N_3057,N_3690);
and U4450 (N_4450,N_3109,N_3271);
nor U4451 (N_4451,N_3626,N_3229);
xor U4452 (N_4452,N_3559,N_3181);
nand U4453 (N_4453,N_3764,N_3094);
or U4454 (N_4454,N_3656,N_3130);
nand U4455 (N_4455,N_3523,N_3012);
nor U4456 (N_4456,N_3374,N_3531);
and U4457 (N_4457,N_3321,N_3280);
nand U4458 (N_4458,N_3469,N_3141);
or U4459 (N_4459,N_3949,N_3358);
nand U4460 (N_4460,N_3008,N_3928);
nor U4461 (N_4461,N_3643,N_3829);
nand U4462 (N_4462,N_3444,N_3625);
or U4463 (N_4463,N_3019,N_3085);
and U4464 (N_4464,N_3616,N_3437);
nand U4465 (N_4465,N_3207,N_3044);
and U4466 (N_4466,N_3413,N_3873);
nor U4467 (N_4467,N_3163,N_3013);
nor U4468 (N_4468,N_3924,N_3617);
nor U4469 (N_4469,N_3408,N_3588);
or U4470 (N_4470,N_3971,N_3591);
and U4471 (N_4471,N_3309,N_3941);
and U4472 (N_4472,N_3653,N_3377);
nor U4473 (N_4473,N_3970,N_3221);
or U4474 (N_4474,N_3723,N_3317);
and U4475 (N_4475,N_3227,N_3029);
nand U4476 (N_4476,N_3527,N_3119);
nand U4477 (N_4477,N_3989,N_3913);
or U4478 (N_4478,N_3740,N_3996);
and U4479 (N_4479,N_3719,N_3774);
nand U4480 (N_4480,N_3375,N_3725);
and U4481 (N_4481,N_3310,N_3054);
xor U4482 (N_4482,N_3118,N_3301);
nand U4483 (N_4483,N_3217,N_3606);
or U4484 (N_4484,N_3721,N_3714);
or U4485 (N_4485,N_3866,N_3361);
nor U4486 (N_4486,N_3541,N_3206);
or U4487 (N_4487,N_3376,N_3396);
or U4488 (N_4488,N_3267,N_3005);
or U4489 (N_4489,N_3086,N_3806);
and U4490 (N_4490,N_3256,N_3167);
nor U4491 (N_4491,N_3983,N_3002);
or U4492 (N_4492,N_3322,N_3176);
or U4493 (N_4493,N_3528,N_3699);
and U4494 (N_4494,N_3775,N_3494);
nor U4495 (N_4495,N_3277,N_3226);
and U4496 (N_4496,N_3908,N_3891);
and U4497 (N_4497,N_3645,N_3465);
nand U4498 (N_4498,N_3132,N_3025);
nor U4499 (N_4499,N_3945,N_3570);
nor U4500 (N_4500,N_3926,N_3157);
nor U4501 (N_4501,N_3422,N_3806);
nor U4502 (N_4502,N_3166,N_3556);
or U4503 (N_4503,N_3123,N_3961);
and U4504 (N_4504,N_3068,N_3771);
nand U4505 (N_4505,N_3234,N_3444);
nand U4506 (N_4506,N_3639,N_3140);
nor U4507 (N_4507,N_3314,N_3552);
nand U4508 (N_4508,N_3967,N_3060);
or U4509 (N_4509,N_3760,N_3913);
and U4510 (N_4510,N_3798,N_3225);
nand U4511 (N_4511,N_3724,N_3693);
xnor U4512 (N_4512,N_3364,N_3970);
nand U4513 (N_4513,N_3512,N_3283);
and U4514 (N_4514,N_3380,N_3133);
nand U4515 (N_4515,N_3534,N_3065);
xnor U4516 (N_4516,N_3266,N_3780);
and U4517 (N_4517,N_3005,N_3071);
nand U4518 (N_4518,N_3562,N_3587);
or U4519 (N_4519,N_3038,N_3079);
nor U4520 (N_4520,N_3399,N_3035);
or U4521 (N_4521,N_3383,N_3987);
nor U4522 (N_4522,N_3042,N_3397);
nor U4523 (N_4523,N_3290,N_3577);
xnor U4524 (N_4524,N_3686,N_3318);
and U4525 (N_4525,N_3232,N_3724);
or U4526 (N_4526,N_3593,N_3077);
nor U4527 (N_4527,N_3729,N_3776);
and U4528 (N_4528,N_3251,N_3924);
nor U4529 (N_4529,N_3985,N_3791);
nor U4530 (N_4530,N_3820,N_3934);
or U4531 (N_4531,N_3308,N_3477);
nor U4532 (N_4532,N_3610,N_3348);
nand U4533 (N_4533,N_3900,N_3877);
nor U4534 (N_4534,N_3571,N_3298);
or U4535 (N_4535,N_3068,N_3081);
or U4536 (N_4536,N_3450,N_3835);
and U4537 (N_4537,N_3617,N_3763);
and U4538 (N_4538,N_3454,N_3664);
nand U4539 (N_4539,N_3857,N_3014);
nand U4540 (N_4540,N_3884,N_3544);
nand U4541 (N_4541,N_3768,N_3288);
nor U4542 (N_4542,N_3588,N_3724);
and U4543 (N_4543,N_3993,N_3829);
and U4544 (N_4544,N_3520,N_3409);
nand U4545 (N_4545,N_3746,N_3738);
or U4546 (N_4546,N_3953,N_3505);
nand U4547 (N_4547,N_3583,N_3190);
xor U4548 (N_4548,N_3063,N_3264);
nor U4549 (N_4549,N_3067,N_3650);
nand U4550 (N_4550,N_3669,N_3245);
nor U4551 (N_4551,N_3330,N_3656);
nand U4552 (N_4552,N_3680,N_3168);
and U4553 (N_4553,N_3443,N_3314);
nor U4554 (N_4554,N_3144,N_3935);
nand U4555 (N_4555,N_3474,N_3660);
nor U4556 (N_4556,N_3995,N_3622);
and U4557 (N_4557,N_3212,N_3978);
nor U4558 (N_4558,N_3643,N_3368);
nor U4559 (N_4559,N_3998,N_3558);
and U4560 (N_4560,N_3092,N_3865);
nand U4561 (N_4561,N_3437,N_3002);
and U4562 (N_4562,N_3935,N_3395);
nand U4563 (N_4563,N_3970,N_3579);
and U4564 (N_4564,N_3812,N_3941);
and U4565 (N_4565,N_3219,N_3009);
or U4566 (N_4566,N_3524,N_3208);
nor U4567 (N_4567,N_3947,N_3737);
xnor U4568 (N_4568,N_3592,N_3940);
and U4569 (N_4569,N_3847,N_3465);
nor U4570 (N_4570,N_3016,N_3614);
nand U4571 (N_4571,N_3785,N_3714);
and U4572 (N_4572,N_3879,N_3262);
or U4573 (N_4573,N_3663,N_3238);
and U4574 (N_4574,N_3275,N_3502);
nand U4575 (N_4575,N_3407,N_3286);
and U4576 (N_4576,N_3837,N_3474);
or U4577 (N_4577,N_3386,N_3043);
nor U4578 (N_4578,N_3677,N_3161);
or U4579 (N_4579,N_3730,N_3863);
or U4580 (N_4580,N_3339,N_3011);
xor U4581 (N_4581,N_3795,N_3887);
nor U4582 (N_4582,N_3118,N_3628);
nand U4583 (N_4583,N_3384,N_3280);
and U4584 (N_4584,N_3516,N_3449);
and U4585 (N_4585,N_3572,N_3668);
or U4586 (N_4586,N_3382,N_3410);
and U4587 (N_4587,N_3456,N_3944);
nand U4588 (N_4588,N_3560,N_3226);
or U4589 (N_4589,N_3350,N_3936);
nor U4590 (N_4590,N_3606,N_3048);
nand U4591 (N_4591,N_3866,N_3561);
nor U4592 (N_4592,N_3328,N_3239);
or U4593 (N_4593,N_3498,N_3569);
and U4594 (N_4594,N_3550,N_3143);
xnor U4595 (N_4595,N_3657,N_3416);
nor U4596 (N_4596,N_3583,N_3556);
or U4597 (N_4597,N_3304,N_3856);
and U4598 (N_4598,N_3075,N_3574);
nand U4599 (N_4599,N_3199,N_3197);
or U4600 (N_4600,N_3183,N_3669);
nor U4601 (N_4601,N_3864,N_3105);
nor U4602 (N_4602,N_3709,N_3241);
nand U4603 (N_4603,N_3647,N_3516);
and U4604 (N_4604,N_3577,N_3762);
nand U4605 (N_4605,N_3505,N_3269);
xor U4606 (N_4606,N_3599,N_3080);
nand U4607 (N_4607,N_3291,N_3792);
or U4608 (N_4608,N_3918,N_3765);
xor U4609 (N_4609,N_3524,N_3442);
nor U4610 (N_4610,N_3924,N_3114);
or U4611 (N_4611,N_3379,N_3409);
or U4612 (N_4612,N_3746,N_3235);
or U4613 (N_4613,N_3506,N_3021);
nand U4614 (N_4614,N_3614,N_3011);
xor U4615 (N_4615,N_3490,N_3409);
or U4616 (N_4616,N_3544,N_3776);
nand U4617 (N_4617,N_3344,N_3807);
nor U4618 (N_4618,N_3281,N_3173);
nor U4619 (N_4619,N_3830,N_3349);
or U4620 (N_4620,N_3120,N_3881);
nor U4621 (N_4621,N_3232,N_3999);
xor U4622 (N_4622,N_3782,N_3829);
and U4623 (N_4623,N_3114,N_3987);
nand U4624 (N_4624,N_3661,N_3856);
and U4625 (N_4625,N_3164,N_3391);
and U4626 (N_4626,N_3349,N_3745);
nor U4627 (N_4627,N_3820,N_3323);
nand U4628 (N_4628,N_3022,N_3158);
or U4629 (N_4629,N_3616,N_3536);
nand U4630 (N_4630,N_3511,N_3014);
xnor U4631 (N_4631,N_3699,N_3659);
or U4632 (N_4632,N_3819,N_3404);
or U4633 (N_4633,N_3915,N_3278);
nand U4634 (N_4634,N_3526,N_3378);
xnor U4635 (N_4635,N_3589,N_3680);
or U4636 (N_4636,N_3987,N_3986);
and U4637 (N_4637,N_3696,N_3536);
or U4638 (N_4638,N_3109,N_3537);
or U4639 (N_4639,N_3949,N_3505);
or U4640 (N_4640,N_3430,N_3313);
nor U4641 (N_4641,N_3848,N_3046);
nand U4642 (N_4642,N_3694,N_3129);
nor U4643 (N_4643,N_3385,N_3920);
nand U4644 (N_4644,N_3748,N_3820);
nor U4645 (N_4645,N_3620,N_3887);
nand U4646 (N_4646,N_3478,N_3339);
and U4647 (N_4647,N_3638,N_3011);
nor U4648 (N_4648,N_3758,N_3918);
and U4649 (N_4649,N_3303,N_3416);
nor U4650 (N_4650,N_3433,N_3713);
and U4651 (N_4651,N_3278,N_3367);
and U4652 (N_4652,N_3613,N_3756);
nor U4653 (N_4653,N_3137,N_3532);
or U4654 (N_4654,N_3683,N_3142);
and U4655 (N_4655,N_3140,N_3740);
and U4656 (N_4656,N_3788,N_3196);
nor U4657 (N_4657,N_3974,N_3320);
and U4658 (N_4658,N_3811,N_3222);
nand U4659 (N_4659,N_3005,N_3015);
or U4660 (N_4660,N_3893,N_3739);
or U4661 (N_4661,N_3614,N_3175);
nand U4662 (N_4662,N_3106,N_3625);
xor U4663 (N_4663,N_3192,N_3446);
nand U4664 (N_4664,N_3476,N_3497);
and U4665 (N_4665,N_3199,N_3736);
nor U4666 (N_4666,N_3108,N_3415);
nand U4667 (N_4667,N_3911,N_3007);
nor U4668 (N_4668,N_3514,N_3559);
or U4669 (N_4669,N_3363,N_3315);
and U4670 (N_4670,N_3061,N_3079);
nand U4671 (N_4671,N_3574,N_3943);
or U4672 (N_4672,N_3538,N_3165);
nor U4673 (N_4673,N_3662,N_3922);
nand U4674 (N_4674,N_3203,N_3847);
nand U4675 (N_4675,N_3036,N_3729);
nor U4676 (N_4676,N_3765,N_3468);
and U4677 (N_4677,N_3683,N_3374);
xor U4678 (N_4678,N_3968,N_3071);
nand U4679 (N_4679,N_3342,N_3039);
and U4680 (N_4680,N_3381,N_3150);
nor U4681 (N_4681,N_3032,N_3828);
or U4682 (N_4682,N_3330,N_3107);
nand U4683 (N_4683,N_3313,N_3298);
xor U4684 (N_4684,N_3485,N_3606);
and U4685 (N_4685,N_3493,N_3585);
or U4686 (N_4686,N_3338,N_3811);
nor U4687 (N_4687,N_3500,N_3980);
nor U4688 (N_4688,N_3074,N_3361);
or U4689 (N_4689,N_3555,N_3778);
nor U4690 (N_4690,N_3190,N_3267);
nor U4691 (N_4691,N_3497,N_3726);
or U4692 (N_4692,N_3664,N_3556);
or U4693 (N_4693,N_3768,N_3528);
and U4694 (N_4694,N_3819,N_3792);
nor U4695 (N_4695,N_3486,N_3313);
nor U4696 (N_4696,N_3240,N_3684);
or U4697 (N_4697,N_3609,N_3587);
xor U4698 (N_4698,N_3756,N_3092);
or U4699 (N_4699,N_3929,N_3266);
nand U4700 (N_4700,N_3278,N_3382);
nor U4701 (N_4701,N_3760,N_3700);
nand U4702 (N_4702,N_3558,N_3054);
nand U4703 (N_4703,N_3786,N_3839);
and U4704 (N_4704,N_3363,N_3644);
nand U4705 (N_4705,N_3152,N_3032);
or U4706 (N_4706,N_3342,N_3334);
or U4707 (N_4707,N_3914,N_3697);
nand U4708 (N_4708,N_3200,N_3782);
or U4709 (N_4709,N_3033,N_3702);
and U4710 (N_4710,N_3728,N_3322);
nand U4711 (N_4711,N_3966,N_3362);
nor U4712 (N_4712,N_3232,N_3530);
nor U4713 (N_4713,N_3157,N_3234);
and U4714 (N_4714,N_3853,N_3213);
nor U4715 (N_4715,N_3344,N_3094);
nand U4716 (N_4716,N_3539,N_3068);
nand U4717 (N_4717,N_3481,N_3856);
or U4718 (N_4718,N_3852,N_3777);
and U4719 (N_4719,N_3039,N_3769);
nand U4720 (N_4720,N_3309,N_3747);
nand U4721 (N_4721,N_3840,N_3009);
nor U4722 (N_4722,N_3289,N_3950);
xnor U4723 (N_4723,N_3130,N_3827);
xnor U4724 (N_4724,N_3812,N_3342);
or U4725 (N_4725,N_3065,N_3663);
nor U4726 (N_4726,N_3672,N_3693);
nor U4727 (N_4727,N_3263,N_3946);
xnor U4728 (N_4728,N_3558,N_3405);
and U4729 (N_4729,N_3710,N_3131);
or U4730 (N_4730,N_3830,N_3149);
nand U4731 (N_4731,N_3524,N_3102);
xnor U4732 (N_4732,N_3608,N_3101);
and U4733 (N_4733,N_3437,N_3447);
nor U4734 (N_4734,N_3317,N_3098);
nand U4735 (N_4735,N_3788,N_3546);
xnor U4736 (N_4736,N_3107,N_3193);
and U4737 (N_4737,N_3037,N_3116);
nand U4738 (N_4738,N_3606,N_3541);
or U4739 (N_4739,N_3387,N_3221);
nand U4740 (N_4740,N_3922,N_3359);
or U4741 (N_4741,N_3862,N_3500);
xnor U4742 (N_4742,N_3775,N_3211);
xnor U4743 (N_4743,N_3654,N_3830);
nand U4744 (N_4744,N_3210,N_3762);
or U4745 (N_4745,N_3029,N_3716);
and U4746 (N_4746,N_3598,N_3524);
nor U4747 (N_4747,N_3298,N_3255);
and U4748 (N_4748,N_3062,N_3783);
nor U4749 (N_4749,N_3059,N_3609);
nand U4750 (N_4750,N_3334,N_3958);
nand U4751 (N_4751,N_3764,N_3074);
and U4752 (N_4752,N_3584,N_3992);
or U4753 (N_4753,N_3114,N_3215);
and U4754 (N_4754,N_3112,N_3080);
nand U4755 (N_4755,N_3658,N_3536);
xnor U4756 (N_4756,N_3379,N_3081);
and U4757 (N_4757,N_3346,N_3388);
and U4758 (N_4758,N_3988,N_3641);
or U4759 (N_4759,N_3645,N_3803);
xnor U4760 (N_4760,N_3909,N_3305);
and U4761 (N_4761,N_3040,N_3617);
xnor U4762 (N_4762,N_3434,N_3588);
or U4763 (N_4763,N_3266,N_3578);
and U4764 (N_4764,N_3237,N_3604);
or U4765 (N_4765,N_3774,N_3769);
xor U4766 (N_4766,N_3653,N_3936);
xnor U4767 (N_4767,N_3192,N_3521);
or U4768 (N_4768,N_3649,N_3968);
xor U4769 (N_4769,N_3165,N_3218);
nand U4770 (N_4770,N_3779,N_3375);
and U4771 (N_4771,N_3322,N_3057);
nor U4772 (N_4772,N_3797,N_3323);
nand U4773 (N_4773,N_3432,N_3733);
or U4774 (N_4774,N_3592,N_3387);
or U4775 (N_4775,N_3271,N_3761);
or U4776 (N_4776,N_3311,N_3905);
nor U4777 (N_4777,N_3594,N_3087);
xor U4778 (N_4778,N_3209,N_3957);
nor U4779 (N_4779,N_3805,N_3388);
and U4780 (N_4780,N_3534,N_3760);
or U4781 (N_4781,N_3123,N_3434);
nor U4782 (N_4782,N_3319,N_3875);
and U4783 (N_4783,N_3841,N_3522);
or U4784 (N_4784,N_3822,N_3457);
or U4785 (N_4785,N_3209,N_3477);
and U4786 (N_4786,N_3802,N_3735);
and U4787 (N_4787,N_3759,N_3134);
or U4788 (N_4788,N_3118,N_3341);
nand U4789 (N_4789,N_3827,N_3039);
nor U4790 (N_4790,N_3144,N_3756);
nor U4791 (N_4791,N_3719,N_3377);
and U4792 (N_4792,N_3604,N_3243);
xor U4793 (N_4793,N_3799,N_3565);
nand U4794 (N_4794,N_3912,N_3375);
nor U4795 (N_4795,N_3711,N_3842);
nand U4796 (N_4796,N_3835,N_3348);
and U4797 (N_4797,N_3264,N_3232);
nor U4798 (N_4798,N_3440,N_3643);
nor U4799 (N_4799,N_3233,N_3760);
or U4800 (N_4800,N_3990,N_3295);
or U4801 (N_4801,N_3310,N_3844);
and U4802 (N_4802,N_3413,N_3593);
and U4803 (N_4803,N_3584,N_3398);
or U4804 (N_4804,N_3661,N_3867);
and U4805 (N_4805,N_3488,N_3757);
nand U4806 (N_4806,N_3517,N_3289);
nand U4807 (N_4807,N_3135,N_3202);
nand U4808 (N_4808,N_3307,N_3683);
or U4809 (N_4809,N_3732,N_3788);
and U4810 (N_4810,N_3129,N_3069);
nand U4811 (N_4811,N_3011,N_3348);
and U4812 (N_4812,N_3115,N_3872);
and U4813 (N_4813,N_3898,N_3442);
and U4814 (N_4814,N_3076,N_3949);
or U4815 (N_4815,N_3241,N_3344);
nor U4816 (N_4816,N_3144,N_3420);
xor U4817 (N_4817,N_3110,N_3374);
or U4818 (N_4818,N_3030,N_3254);
nand U4819 (N_4819,N_3642,N_3504);
nor U4820 (N_4820,N_3574,N_3427);
and U4821 (N_4821,N_3931,N_3925);
nor U4822 (N_4822,N_3875,N_3100);
or U4823 (N_4823,N_3027,N_3372);
or U4824 (N_4824,N_3519,N_3761);
or U4825 (N_4825,N_3722,N_3763);
nand U4826 (N_4826,N_3060,N_3144);
nand U4827 (N_4827,N_3894,N_3874);
nor U4828 (N_4828,N_3510,N_3972);
nor U4829 (N_4829,N_3581,N_3353);
or U4830 (N_4830,N_3661,N_3828);
nand U4831 (N_4831,N_3814,N_3318);
nor U4832 (N_4832,N_3196,N_3897);
xnor U4833 (N_4833,N_3315,N_3059);
nor U4834 (N_4834,N_3274,N_3531);
and U4835 (N_4835,N_3428,N_3490);
nand U4836 (N_4836,N_3041,N_3814);
xnor U4837 (N_4837,N_3788,N_3964);
and U4838 (N_4838,N_3650,N_3902);
and U4839 (N_4839,N_3925,N_3253);
xor U4840 (N_4840,N_3548,N_3665);
and U4841 (N_4841,N_3582,N_3998);
and U4842 (N_4842,N_3067,N_3782);
and U4843 (N_4843,N_3554,N_3339);
nand U4844 (N_4844,N_3397,N_3007);
nand U4845 (N_4845,N_3575,N_3088);
or U4846 (N_4846,N_3875,N_3697);
and U4847 (N_4847,N_3295,N_3574);
and U4848 (N_4848,N_3685,N_3102);
nor U4849 (N_4849,N_3825,N_3307);
nand U4850 (N_4850,N_3107,N_3489);
nor U4851 (N_4851,N_3128,N_3428);
nor U4852 (N_4852,N_3780,N_3269);
nand U4853 (N_4853,N_3469,N_3189);
nor U4854 (N_4854,N_3582,N_3155);
xor U4855 (N_4855,N_3063,N_3085);
nor U4856 (N_4856,N_3069,N_3463);
nand U4857 (N_4857,N_3584,N_3613);
or U4858 (N_4858,N_3534,N_3467);
nor U4859 (N_4859,N_3453,N_3345);
nand U4860 (N_4860,N_3927,N_3378);
nand U4861 (N_4861,N_3116,N_3315);
nor U4862 (N_4862,N_3481,N_3713);
xor U4863 (N_4863,N_3533,N_3463);
or U4864 (N_4864,N_3272,N_3360);
and U4865 (N_4865,N_3162,N_3967);
nand U4866 (N_4866,N_3683,N_3759);
or U4867 (N_4867,N_3032,N_3662);
nand U4868 (N_4868,N_3437,N_3974);
nand U4869 (N_4869,N_3898,N_3241);
nand U4870 (N_4870,N_3369,N_3729);
nor U4871 (N_4871,N_3446,N_3224);
nor U4872 (N_4872,N_3389,N_3423);
nor U4873 (N_4873,N_3428,N_3346);
and U4874 (N_4874,N_3153,N_3183);
or U4875 (N_4875,N_3589,N_3235);
nor U4876 (N_4876,N_3240,N_3416);
and U4877 (N_4877,N_3242,N_3957);
nand U4878 (N_4878,N_3234,N_3568);
nor U4879 (N_4879,N_3801,N_3075);
nand U4880 (N_4880,N_3470,N_3246);
and U4881 (N_4881,N_3131,N_3473);
nor U4882 (N_4882,N_3350,N_3434);
nor U4883 (N_4883,N_3167,N_3664);
or U4884 (N_4884,N_3304,N_3195);
nor U4885 (N_4885,N_3779,N_3801);
nand U4886 (N_4886,N_3721,N_3702);
nor U4887 (N_4887,N_3038,N_3504);
and U4888 (N_4888,N_3582,N_3291);
nand U4889 (N_4889,N_3521,N_3278);
and U4890 (N_4890,N_3040,N_3252);
nand U4891 (N_4891,N_3877,N_3875);
nand U4892 (N_4892,N_3494,N_3908);
nor U4893 (N_4893,N_3146,N_3603);
nand U4894 (N_4894,N_3854,N_3644);
nand U4895 (N_4895,N_3602,N_3994);
nand U4896 (N_4896,N_3324,N_3724);
xnor U4897 (N_4897,N_3558,N_3584);
and U4898 (N_4898,N_3806,N_3466);
xor U4899 (N_4899,N_3426,N_3055);
xnor U4900 (N_4900,N_3179,N_3541);
nand U4901 (N_4901,N_3274,N_3848);
and U4902 (N_4902,N_3654,N_3741);
and U4903 (N_4903,N_3270,N_3630);
xor U4904 (N_4904,N_3977,N_3403);
or U4905 (N_4905,N_3714,N_3923);
nand U4906 (N_4906,N_3739,N_3188);
nor U4907 (N_4907,N_3064,N_3354);
nand U4908 (N_4908,N_3832,N_3461);
or U4909 (N_4909,N_3333,N_3536);
nand U4910 (N_4910,N_3372,N_3152);
nand U4911 (N_4911,N_3403,N_3503);
nor U4912 (N_4912,N_3748,N_3728);
and U4913 (N_4913,N_3483,N_3512);
and U4914 (N_4914,N_3061,N_3776);
or U4915 (N_4915,N_3002,N_3780);
nand U4916 (N_4916,N_3293,N_3860);
nand U4917 (N_4917,N_3551,N_3847);
xnor U4918 (N_4918,N_3639,N_3358);
and U4919 (N_4919,N_3718,N_3440);
or U4920 (N_4920,N_3089,N_3748);
nor U4921 (N_4921,N_3198,N_3602);
and U4922 (N_4922,N_3589,N_3303);
and U4923 (N_4923,N_3789,N_3913);
nor U4924 (N_4924,N_3480,N_3912);
or U4925 (N_4925,N_3465,N_3783);
nor U4926 (N_4926,N_3281,N_3537);
and U4927 (N_4927,N_3357,N_3760);
nor U4928 (N_4928,N_3026,N_3794);
and U4929 (N_4929,N_3004,N_3671);
nand U4930 (N_4930,N_3543,N_3587);
or U4931 (N_4931,N_3061,N_3921);
and U4932 (N_4932,N_3923,N_3858);
and U4933 (N_4933,N_3767,N_3757);
or U4934 (N_4934,N_3242,N_3807);
nor U4935 (N_4935,N_3440,N_3414);
xnor U4936 (N_4936,N_3398,N_3516);
and U4937 (N_4937,N_3375,N_3829);
nor U4938 (N_4938,N_3638,N_3009);
nand U4939 (N_4939,N_3239,N_3438);
nor U4940 (N_4940,N_3275,N_3194);
or U4941 (N_4941,N_3262,N_3548);
nor U4942 (N_4942,N_3116,N_3615);
nand U4943 (N_4943,N_3568,N_3970);
xnor U4944 (N_4944,N_3649,N_3915);
nor U4945 (N_4945,N_3973,N_3592);
nor U4946 (N_4946,N_3972,N_3985);
or U4947 (N_4947,N_3471,N_3677);
or U4948 (N_4948,N_3422,N_3290);
and U4949 (N_4949,N_3177,N_3885);
and U4950 (N_4950,N_3084,N_3611);
and U4951 (N_4951,N_3173,N_3975);
or U4952 (N_4952,N_3266,N_3918);
and U4953 (N_4953,N_3616,N_3039);
xor U4954 (N_4954,N_3821,N_3196);
nor U4955 (N_4955,N_3469,N_3242);
or U4956 (N_4956,N_3334,N_3265);
nor U4957 (N_4957,N_3309,N_3359);
or U4958 (N_4958,N_3571,N_3348);
nor U4959 (N_4959,N_3469,N_3293);
nor U4960 (N_4960,N_3162,N_3581);
nand U4961 (N_4961,N_3117,N_3017);
or U4962 (N_4962,N_3716,N_3063);
xnor U4963 (N_4963,N_3520,N_3942);
or U4964 (N_4964,N_3524,N_3215);
nand U4965 (N_4965,N_3447,N_3810);
xnor U4966 (N_4966,N_3653,N_3381);
xnor U4967 (N_4967,N_3790,N_3650);
and U4968 (N_4968,N_3749,N_3560);
nor U4969 (N_4969,N_3315,N_3104);
nand U4970 (N_4970,N_3129,N_3598);
nand U4971 (N_4971,N_3837,N_3272);
and U4972 (N_4972,N_3579,N_3503);
or U4973 (N_4973,N_3851,N_3654);
xnor U4974 (N_4974,N_3579,N_3217);
xor U4975 (N_4975,N_3606,N_3688);
nand U4976 (N_4976,N_3276,N_3454);
and U4977 (N_4977,N_3660,N_3966);
nor U4978 (N_4978,N_3214,N_3709);
nand U4979 (N_4979,N_3624,N_3512);
nand U4980 (N_4980,N_3899,N_3669);
nand U4981 (N_4981,N_3552,N_3877);
and U4982 (N_4982,N_3267,N_3015);
nor U4983 (N_4983,N_3952,N_3462);
and U4984 (N_4984,N_3210,N_3045);
and U4985 (N_4985,N_3415,N_3444);
nor U4986 (N_4986,N_3487,N_3986);
nor U4987 (N_4987,N_3889,N_3071);
or U4988 (N_4988,N_3675,N_3920);
or U4989 (N_4989,N_3719,N_3841);
xor U4990 (N_4990,N_3549,N_3567);
nand U4991 (N_4991,N_3521,N_3018);
or U4992 (N_4992,N_3427,N_3587);
and U4993 (N_4993,N_3415,N_3122);
nor U4994 (N_4994,N_3712,N_3870);
and U4995 (N_4995,N_3715,N_3937);
nand U4996 (N_4996,N_3998,N_3290);
and U4997 (N_4997,N_3920,N_3881);
nor U4998 (N_4998,N_3887,N_3392);
or U4999 (N_4999,N_3267,N_3359);
xor UO_0 (O_0,N_4000,N_4185);
nand UO_1 (O_1,N_4855,N_4626);
or UO_2 (O_2,N_4090,N_4588);
and UO_3 (O_3,N_4919,N_4151);
nand UO_4 (O_4,N_4602,N_4788);
nand UO_5 (O_5,N_4763,N_4582);
nor UO_6 (O_6,N_4375,N_4775);
nor UO_7 (O_7,N_4664,N_4565);
nand UO_8 (O_8,N_4608,N_4340);
xnor UO_9 (O_9,N_4973,N_4689);
or UO_10 (O_10,N_4272,N_4121);
or UO_11 (O_11,N_4350,N_4743);
and UO_12 (O_12,N_4207,N_4378);
xnor UO_13 (O_13,N_4562,N_4753);
nand UO_14 (O_14,N_4130,N_4195);
or UO_15 (O_15,N_4591,N_4316);
nand UO_16 (O_16,N_4771,N_4766);
and UO_17 (O_17,N_4963,N_4639);
or UO_18 (O_18,N_4169,N_4699);
nand UO_19 (O_19,N_4358,N_4936);
or UO_20 (O_20,N_4509,N_4597);
nand UO_21 (O_21,N_4019,N_4967);
or UO_22 (O_22,N_4225,N_4533);
or UO_23 (O_23,N_4604,N_4240);
nor UO_24 (O_24,N_4387,N_4510);
and UO_25 (O_25,N_4152,N_4612);
nand UO_26 (O_26,N_4924,N_4023);
and UO_27 (O_27,N_4806,N_4999);
or UO_28 (O_28,N_4516,N_4268);
and UO_29 (O_29,N_4614,N_4912);
and UO_30 (O_30,N_4101,N_4552);
nor UO_31 (O_31,N_4459,N_4972);
or UO_32 (O_32,N_4096,N_4333);
nand UO_33 (O_33,N_4921,N_4535);
nand UO_34 (O_34,N_4424,N_4022);
and UO_35 (O_35,N_4851,N_4700);
and UO_36 (O_36,N_4188,N_4232);
and UO_37 (O_37,N_4498,N_4128);
or UO_38 (O_38,N_4482,N_4910);
nor UO_39 (O_39,N_4646,N_4768);
and UO_40 (O_40,N_4979,N_4944);
nand UO_41 (O_41,N_4359,N_4094);
or UO_42 (O_42,N_4795,N_4113);
nor UO_43 (O_43,N_4881,N_4901);
nor UO_44 (O_44,N_4647,N_4469);
nor UO_45 (O_45,N_4466,N_4114);
and UO_46 (O_46,N_4012,N_4236);
nor UO_47 (O_47,N_4968,N_4291);
and UO_48 (O_48,N_4808,N_4030);
xor UO_49 (O_49,N_4941,N_4220);
nand UO_50 (O_50,N_4460,N_4519);
and UO_51 (O_51,N_4837,N_4040);
nor UO_52 (O_52,N_4628,N_4401);
nand UO_53 (O_53,N_4418,N_4002);
or UO_54 (O_54,N_4122,N_4727);
or UO_55 (O_55,N_4391,N_4678);
and UO_56 (O_56,N_4497,N_4405);
and UO_57 (O_57,N_4539,N_4632);
nor UO_58 (O_58,N_4015,N_4731);
and UO_59 (O_59,N_4421,N_4398);
and UO_60 (O_60,N_4849,N_4112);
or UO_61 (O_61,N_4988,N_4288);
or UO_62 (O_62,N_4934,N_4408);
or UO_63 (O_63,N_4357,N_4875);
xnor UO_64 (O_64,N_4645,N_4013);
nor UO_65 (O_65,N_4158,N_4654);
and UO_66 (O_66,N_4903,N_4897);
or UO_67 (O_67,N_4736,N_4131);
or UO_68 (O_68,N_4715,N_4947);
and UO_69 (O_69,N_4043,N_4992);
nand UO_70 (O_70,N_4267,N_4545);
and UO_71 (O_71,N_4540,N_4735);
and UO_72 (O_72,N_4784,N_4813);
and UO_73 (O_73,N_4377,N_4550);
and UO_74 (O_74,N_4426,N_4842);
or UO_75 (O_75,N_4184,N_4099);
or UO_76 (O_76,N_4242,N_4135);
nand UO_77 (O_77,N_4410,N_4517);
and UO_78 (O_78,N_4790,N_4153);
or UO_79 (O_79,N_4933,N_4662);
or UO_80 (O_80,N_4106,N_4073);
or UO_81 (O_81,N_4390,N_4446);
nor UO_82 (O_82,N_4801,N_4658);
and UO_83 (O_83,N_4235,N_4494);
nand UO_84 (O_84,N_4009,N_4385);
and UO_85 (O_85,N_4816,N_4622);
or UO_86 (O_86,N_4861,N_4351);
nand UO_87 (O_87,N_4422,N_4760);
nand UO_88 (O_88,N_4204,N_4470);
nor UO_89 (O_89,N_4275,N_4896);
or UO_90 (O_90,N_4889,N_4172);
nand UO_91 (O_91,N_4990,N_4276);
nand UO_92 (O_92,N_4441,N_4835);
xnor UO_93 (O_93,N_4782,N_4071);
and UO_94 (O_94,N_4825,N_4860);
or UO_95 (O_95,N_4521,N_4064);
and UO_96 (O_96,N_4799,N_4066);
nand UO_97 (O_97,N_4303,N_4681);
or UO_98 (O_98,N_4491,N_4812);
xor UO_99 (O_99,N_4286,N_4167);
nand UO_100 (O_100,N_4804,N_4862);
or UO_101 (O_101,N_4037,N_4916);
or UO_102 (O_102,N_4674,N_4199);
and UO_103 (O_103,N_4794,N_4530);
and UO_104 (O_104,N_4697,N_4415);
nor UO_105 (O_105,N_4708,N_4124);
and UO_106 (O_106,N_4176,N_4007);
nand UO_107 (O_107,N_4512,N_4493);
nor UO_108 (O_108,N_4179,N_4698);
or UO_109 (O_109,N_4954,N_4585);
xor UO_110 (O_110,N_4214,N_4140);
and UO_111 (O_111,N_4939,N_4624);
or UO_112 (O_112,N_4311,N_4822);
or UO_113 (O_113,N_4156,N_4453);
or UO_114 (O_114,N_4706,N_4984);
or UO_115 (O_115,N_4998,N_4909);
and UO_116 (O_116,N_4435,N_4331);
nand UO_117 (O_117,N_4504,N_4050);
or UO_118 (O_118,N_4868,N_4117);
nand UO_119 (O_119,N_4738,N_4783);
xor UO_120 (O_120,N_4887,N_4219);
or UO_121 (O_121,N_4792,N_4922);
nand UO_122 (O_122,N_4252,N_4301);
or UO_123 (O_123,N_4427,N_4567);
nand UO_124 (O_124,N_4356,N_4273);
nor UO_125 (O_125,N_4171,N_4474);
and UO_126 (O_126,N_4492,N_4890);
nand UO_127 (O_127,N_4619,N_4338);
nand UO_128 (O_128,N_4430,N_4029);
nand UO_129 (O_129,N_4513,N_4383);
and UO_130 (O_130,N_4717,N_4611);
nor UO_131 (O_131,N_4758,N_4857);
or UO_132 (O_132,N_4661,N_4069);
nor UO_133 (O_133,N_4118,N_4249);
xor UO_134 (O_134,N_4160,N_4336);
nand UO_135 (O_135,N_4278,N_4823);
and UO_136 (O_136,N_4977,N_4584);
nand UO_137 (O_137,N_4650,N_4965);
xor UO_138 (O_138,N_4993,N_4821);
nor UO_139 (O_139,N_4770,N_4480);
nand UO_140 (O_140,N_4058,N_4168);
xnor UO_141 (O_141,N_4300,N_4399);
and UO_142 (O_142,N_4483,N_4100);
nor UO_143 (O_143,N_4814,N_4985);
and UO_144 (O_144,N_4044,N_4828);
xnor UO_145 (O_145,N_4244,N_4779);
nor UO_146 (O_146,N_4871,N_4014);
or UO_147 (O_147,N_4729,N_4579);
and UO_148 (O_148,N_4226,N_4655);
and UO_149 (O_149,N_4248,N_4210);
nand UO_150 (O_150,N_4544,N_4008);
nand UO_151 (O_151,N_4233,N_4320);
and UO_152 (O_152,N_4913,N_4221);
nand UO_153 (O_153,N_4891,N_4894);
or UO_154 (O_154,N_4949,N_4297);
or UO_155 (O_155,N_4149,N_4292);
xor UO_156 (O_156,N_4634,N_4379);
nor UO_157 (O_157,N_4344,N_4083);
or UO_158 (O_158,N_4730,N_4187);
nor UO_159 (O_159,N_4028,N_4082);
nor UO_160 (O_160,N_4127,N_4329);
nand UO_161 (O_161,N_4175,N_4917);
xor UO_162 (O_162,N_4580,N_4609);
nand UO_163 (O_163,N_4927,N_4734);
nand UO_164 (O_164,N_4852,N_4873);
xor UO_165 (O_165,N_4874,N_4695);
or UO_166 (O_166,N_4092,N_4606);
and UO_167 (O_167,N_4613,N_4648);
or UO_168 (O_168,N_4209,N_4380);
nor UO_169 (O_169,N_4104,N_4756);
or UO_170 (O_170,N_4136,N_4328);
or UO_171 (O_171,N_4367,N_4259);
nor UO_172 (O_172,N_4159,N_4772);
or UO_173 (O_173,N_4895,N_4991);
nor UO_174 (O_174,N_4507,N_4712);
and UO_175 (O_175,N_4419,N_4728);
nand UO_176 (O_176,N_4425,N_4062);
xor UO_177 (O_177,N_4462,N_4599);
and UO_178 (O_178,N_4803,N_4392);
xnor UO_179 (O_179,N_4886,N_4053);
nor UO_180 (O_180,N_4475,N_4583);
or UO_181 (O_181,N_4036,N_4141);
nand UO_182 (O_182,N_4631,N_4722);
xor UO_183 (O_183,N_4087,N_4039);
nand UO_184 (O_184,N_4797,N_4411);
and UO_185 (O_185,N_4557,N_4250);
nand UO_186 (O_186,N_4749,N_4701);
and UO_187 (O_187,N_4366,N_4508);
nor UO_188 (O_188,N_4072,N_4395);
and UO_189 (O_189,N_4637,N_4742);
or UO_190 (O_190,N_4145,N_4164);
and UO_191 (O_191,N_4590,N_4757);
nand UO_192 (O_192,N_4810,N_4070);
and UO_193 (O_193,N_4865,N_4528);
or UO_194 (O_194,N_4971,N_4067);
nand UO_195 (O_195,N_4417,N_4203);
and UO_196 (O_196,N_4080,N_4900);
or UO_197 (O_197,N_4433,N_4057);
xor UO_198 (O_198,N_4989,N_4705);
nand UO_199 (O_199,N_4047,N_4975);
nand UO_200 (O_200,N_4313,N_4107);
and UO_201 (O_201,N_4659,N_4386);
nand UO_202 (O_202,N_4274,N_4515);
nand UO_203 (O_203,N_4520,N_4490);
nor UO_204 (O_204,N_4110,N_4413);
nor UO_205 (O_205,N_4031,N_4093);
nor UO_206 (O_206,N_4183,N_4181);
xnor UO_207 (O_207,N_4231,N_4665);
xnor UO_208 (O_208,N_4255,N_4294);
nor UO_209 (O_209,N_4502,N_4981);
and UO_210 (O_210,N_4677,N_4572);
and UO_211 (O_211,N_4952,N_4819);
or UO_212 (O_212,N_4923,N_4234);
nand UO_213 (O_213,N_4098,N_4690);
and UO_214 (O_214,N_4287,N_4341);
nor UO_215 (O_215,N_4120,N_4123);
and UO_216 (O_216,N_4404,N_4832);
or UO_217 (O_217,N_4230,N_4443);
xnor UO_218 (O_218,N_4780,N_4452);
and UO_219 (O_219,N_4623,N_4636);
nand UO_220 (O_220,N_4551,N_4553);
xor UO_221 (O_221,N_4505,N_4721);
and UO_222 (O_222,N_4696,N_4056);
or UO_223 (O_223,N_4615,N_4154);
or UO_224 (O_224,N_4033,N_4996);
and UO_225 (O_225,N_4845,N_4467);
nand UO_226 (O_226,N_4461,N_4538);
and UO_227 (O_227,N_4724,N_4293);
nand UO_228 (O_228,N_4960,N_4027);
nand UO_229 (O_229,N_4620,N_4046);
nor UO_230 (O_230,N_4206,N_4005);
nand UO_231 (O_231,N_4077,N_4532);
nand UO_232 (O_232,N_4915,N_4270);
nor UO_233 (O_233,N_4683,N_4866);
nor UO_234 (O_234,N_4197,N_4431);
nor UO_235 (O_235,N_4885,N_4076);
and UO_236 (O_236,N_4192,N_4983);
nor UO_237 (O_237,N_4725,N_4966);
or UO_238 (O_238,N_4877,N_4353);
or UO_239 (O_239,N_4908,N_4327);
and UO_240 (O_240,N_4693,N_4003);
xnor UO_241 (O_241,N_4440,N_4878);
or UO_242 (O_242,N_4173,N_4126);
and UO_243 (O_243,N_4537,N_4299);
nor UO_244 (O_244,N_4254,N_4578);
or UO_245 (O_245,N_4097,N_4116);
and UO_246 (O_246,N_4266,N_4133);
or UO_247 (O_247,N_4381,N_4246);
or UO_248 (O_248,N_4525,N_4777);
and UO_249 (O_249,N_4481,N_4935);
nor UO_250 (O_250,N_4503,N_4263);
nor UO_251 (O_251,N_4305,N_4447);
nand UO_252 (O_252,N_4575,N_4224);
nand UO_253 (O_253,N_4931,N_4959);
xor UO_254 (O_254,N_4563,N_4476);
or UO_255 (O_255,N_4256,N_4884);
xnor UO_256 (O_256,N_4858,N_4409);
and UO_257 (O_257,N_4864,N_4957);
nor UO_258 (O_258,N_4764,N_4215);
nor UO_259 (O_259,N_4928,N_4325);
nor UO_260 (O_260,N_4995,N_4869);
xor UO_261 (O_261,N_4484,N_4834);
nor UO_262 (O_262,N_4307,N_4017);
and UO_263 (O_263,N_4618,N_4593);
nor UO_264 (O_264,N_4354,N_4719);
nand UO_265 (O_265,N_4004,N_4295);
or UO_266 (O_266,N_4940,N_4531);
and UO_267 (O_267,N_4867,N_4463);
or UO_268 (O_268,N_4376,N_4671);
or UO_269 (O_269,N_4312,N_4450);
or UO_270 (O_270,N_4704,N_4271);
and UO_271 (O_271,N_4045,N_4211);
or UO_272 (O_272,N_4198,N_4456);
nand UO_273 (O_273,N_4364,N_4337);
xor UO_274 (O_274,N_4111,N_4581);
nor UO_275 (O_275,N_4147,N_4946);
nor UO_276 (O_276,N_4938,N_4554);
nand UO_277 (O_277,N_4950,N_4601);
or UO_278 (O_278,N_4129,N_4257);
and UO_279 (O_279,N_4281,N_4429);
nand UO_280 (O_280,N_4514,N_4798);
and UO_281 (O_281,N_4302,N_4888);
nor UO_282 (O_282,N_4929,N_4744);
and UO_283 (O_283,N_4347,N_4943);
nand UO_284 (O_284,N_4279,N_4407);
nor UO_285 (O_285,N_4883,N_4846);
and UO_286 (O_286,N_4346,N_4564);
or UO_287 (O_287,N_4853,N_4899);
nand UO_288 (O_288,N_4872,N_4711);
nand UO_289 (O_289,N_4063,N_4652);
xor UO_290 (O_290,N_4826,N_4166);
xnor UO_291 (O_291,N_4177,N_4746);
nor UO_292 (O_292,N_4132,N_4091);
nor UO_293 (O_293,N_4412,N_4818);
xnor UO_294 (O_294,N_4710,N_4994);
nor UO_295 (O_295,N_4194,N_4548);
and UO_296 (O_296,N_4925,N_4560);
xor UO_297 (O_297,N_4605,N_4789);
nor UO_298 (O_298,N_4880,N_4032);
nor UO_299 (O_299,N_4633,N_4109);
nand UO_300 (O_300,N_4958,N_4389);
nand UO_301 (O_301,N_4892,N_4260);
nand UO_302 (O_302,N_4060,N_4685);
and UO_303 (O_303,N_4393,N_4640);
and UO_304 (O_304,N_4824,N_4360);
nand UO_305 (O_305,N_4059,N_4061);
nand UO_306 (O_306,N_4807,N_4522);
and UO_307 (O_307,N_4773,N_4987);
nand UO_308 (O_308,N_4449,N_4369);
nand UO_309 (O_309,N_4568,N_4144);
and UO_310 (O_310,N_4355,N_4682);
nor UO_311 (O_311,N_4397,N_4428);
and UO_312 (O_312,N_4241,N_4577);
xnor UO_313 (O_313,N_4629,N_4285);
or UO_314 (O_314,N_4054,N_4223);
or UO_315 (O_315,N_4870,N_4751);
or UO_316 (O_316,N_4339,N_4786);
and UO_317 (O_317,N_4836,N_4603);
nand UO_318 (O_318,N_4186,N_4833);
nand UO_319 (O_319,N_4669,N_4208);
nand UO_320 (O_320,N_4205,N_4394);
nor UO_321 (O_321,N_4815,N_4907);
or UO_322 (O_322,N_4472,N_4638);
xor UO_323 (O_323,N_4089,N_4086);
and UO_324 (O_324,N_4034,N_4666);
nand UO_325 (O_325,N_4660,N_4668);
or UO_326 (O_326,N_4400,N_4559);
nor UO_327 (O_327,N_4477,N_4523);
nand UO_328 (O_328,N_4103,N_4684);
xor UO_329 (O_329,N_4332,N_4318);
nor UO_330 (O_330,N_4956,N_4371);
nand UO_331 (O_331,N_4253,N_4511);
nand UO_332 (O_332,N_4189,N_4001);
and UO_333 (O_333,N_4905,N_4157);
nor UO_334 (O_334,N_4420,N_4163);
nor UO_335 (O_335,N_4536,N_4844);
nor UO_336 (O_336,N_4774,N_4304);
nor UO_337 (O_337,N_4641,N_4269);
nand UO_338 (O_338,N_4840,N_4841);
nor UO_339 (O_339,N_4762,N_4561);
and UO_340 (O_340,N_4951,N_4595);
nor UO_341 (O_341,N_4587,N_4384);
or UO_342 (O_342,N_4627,N_4778);
or UO_343 (O_343,N_4437,N_4296);
or UO_344 (O_344,N_4937,N_4079);
nand UO_345 (O_345,N_4343,N_4918);
and UO_346 (O_346,N_4914,N_4191);
or UO_347 (O_347,N_4306,N_4330);
and UO_348 (O_348,N_4196,N_4709);
or UO_349 (O_349,N_4458,N_4974);
nor UO_350 (O_350,N_4193,N_4718);
and UO_351 (O_351,N_4524,N_4997);
nor UO_352 (O_352,N_4362,N_4970);
nor UO_353 (O_353,N_4178,N_4969);
nand UO_354 (O_354,N_4882,N_4500);
or UO_355 (O_355,N_4911,N_4457);
and UO_356 (O_356,N_4809,N_4675);
and UO_357 (O_357,N_4839,N_4566);
or UO_358 (O_358,N_4703,N_4906);
nor UO_359 (O_359,N_4251,N_4055);
or UO_360 (O_360,N_4434,N_4657);
nor UO_361 (O_361,N_4679,N_4543);
nor UO_362 (O_362,N_4932,N_4863);
nor UO_363 (O_363,N_4594,N_4010);
or UO_364 (O_364,N_4573,N_4800);
and UO_365 (O_365,N_4085,N_4237);
nor UO_366 (O_366,N_4372,N_4656);
and UO_367 (O_367,N_4737,N_4289);
and UO_368 (O_368,N_4243,N_4326);
or UO_369 (O_369,N_4468,N_4961);
and UO_370 (O_370,N_4048,N_4964);
and UO_371 (O_371,N_4688,N_4438);
nor UO_372 (O_372,N_4478,N_4643);
and UO_373 (O_373,N_4796,N_4370);
nand UO_374 (O_374,N_4290,N_4649);
nor UO_375 (O_375,N_4487,N_4651);
nor UO_376 (O_376,N_4811,N_4451);
nand UO_377 (O_377,N_4432,N_4170);
and UO_378 (O_378,N_4108,N_4444);
nand UO_379 (O_379,N_4838,N_4694);
or UO_380 (O_380,N_4785,N_4038);
or UO_381 (O_381,N_4495,N_4119);
or UO_382 (O_382,N_4222,N_4319);
xnor UO_383 (O_383,N_4436,N_4228);
nand UO_384 (O_384,N_4202,N_4345);
xor UO_385 (O_385,N_4817,N_4042);
and UO_386 (O_386,N_4365,N_4388);
and UO_387 (O_387,N_4542,N_4464);
xor UO_388 (O_388,N_4569,N_4239);
nand UO_389 (O_389,N_4741,N_4716);
nor UO_390 (O_390,N_4315,N_4748);
nand UO_391 (O_391,N_4663,N_4283);
nand UO_392 (O_392,N_4556,N_4454);
nand UO_393 (O_393,N_4733,N_4879);
and UO_394 (O_394,N_4282,N_4948);
nor UO_395 (O_395,N_4499,N_4396);
or UO_396 (O_396,N_4732,N_4174);
or UO_397 (O_397,N_4547,N_4755);
and UO_398 (O_398,N_4115,N_4625);
or UO_399 (O_399,N_4361,N_4754);
nor UO_400 (O_400,N_4217,N_4363);
nor UO_401 (O_401,N_4025,N_4317);
nand UO_402 (O_402,N_4201,N_4750);
xnor UO_403 (O_403,N_4518,N_4150);
or UO_404 (O_404,N_4075,N_4382);
and UO_405 (O_405,N_4769,N_4955);
nand UO_406 (O_406,N_4739,N_4667);
or UO_407 (O_407,N_4713,N_4617);
and UO_408 (O_408,N_4616,N_4155);
nor UO_409 (O_409,N_4308,N_4549);
or UO_410 (O_410,N_4829,N_4827);
and UO_411 (O_411,N_4759,N_4501);
and UO_412 (O_412,N_4479,N_4526);
and UO_413 (O_413,N_4847,N_4767);
nor UO_414 (O_414,N_4607,N_4621);
or UO_415 (O_415,N_4335,N_4247);
nor UO_416 (O_416,N_4793,N_4238);
or UO_417 (O_417,N_4740,N_4374);
or UO_418 (O_418,N_4102,N_4323);
and UO_419 (O_419,N_4555,N_4488);
nand UO_420 (O_420,N_4850,N_4787);
or UO_421 (O_421,N_4496,N_4898);
or UO_422 (O_422,N_4541,N_4848);
nor UO_423 (O_423,N_4920,N_4084);
nor UO_424 (O_424,N_4720,N_4021);
nor UO_425 (O_425,N_4723,N_4714);
nand UO_426 (O_426,N_4200,N_4781);
or UO_427 (O_427,N_4527,N_4074);
and UO_428 (O_428,N_4471,N_4776);
nand UO_429 (O_429,N_4423,N_4105);
or UO_430 (O_430,N_4190,N_4342);
and UO_431 (O_431,N_4026,N_4635);
nor UO_432 (O_432,N_4416,N_4747);
and UO_433 (O_433,N_4644,N_4506);
nand UO_434 (O_434,N_4321,N_4180);
nand UO_435 (O_435,N_4653,N_4485);
nand UO_436 (O_436,N_4610,N_4258);
and UO_437 (O_437,N_4314,N_4065);
xnor UO_438 (O_438,N_4402,N_4686);
nand UO_439 (O_439,N_4672,N_4707);
and UO_440 (O_440,N_4489,N_4596);
nand UO_441 (O_441,N_4264,N_4265);
nor UO_442 (O_442,N_4902,N_4962);
xor UO_443 (O_443,N_4081,N_4843);
or UO_444 (O_444,N_4349,N_4529);
nand UO_445 (O_445,N_4820,N_4765);
and UO_446 (O_446,N_4041,N_4138);
nand UO_447 (O_447,N_4280,N_4830);
nor UO_448 (O_448,N_4162,N_4049);
nand UO_449 (O_449,N_4348,N_4142);
and UO_450 (O_450,N_4859,N_4245);
or UO_451 (O_451,N_4893,N_4805);
or UO_452 (O_452,N_4670,N_4448);
nand UO_453 (O_453,N_4791,N_4051);
and UO_454 (O_454,N_4035,N_4182);
and UO_455 (O_455,N_4558,N_4455);
and UO_456 (O_456,N_4831,N_4761);
nand UO_457 (O_457,N_4016,N_4006);
nor UO_458 (O_458,N_4691,N_4227);
nor UO_459 (O_459,N_4322,N_4352);
xor UO_460 (O_460,N_4692,N_4143);
or UO_461 (O_461,N_4020,N_4024);
nor UO_462 (O_462,N_4368,N_4702);
or UO_463 (O_463,N_4403,N_4953);
or UO_464 (O_464,N_4442,N_4473);
nand UO_465 (O_465,N_4574,N_4465);
nor UO_466 (O_466,N_4125,N_4078);
nand UO_467 (O_467,N_4570,N_4095);
or UO_468 (O_468,N_4600,N_4134);
nor UO_469 (O_469,N_4676,N_4687);
and UO_470 (O_470,N_4229,N_4088);
or UO_471 (O_471,N_4011,N_4976);
xor UO_472 (O_472,N_4146,N_4148);
or UO_473 (O_473,N_4598,N_4218);
and UO_474 (O_474,N_4298,N_4262);
and UO_475 (O_475,N_4592,N_4680);
nor UO_476 (O_476,N_4534,N_4576);
nand UO_477 (O_477,N_4726,N_4589);
and UO_478 (O_478,N_4439,N_4930);
nand UO_479 (O_479,N_4216,N_4261);
nor UO_480 (O_480,N_4310,N_4277);
nand UO_481 (O_481,N_4904,N_4052);
nand UO_482 (O_482,N_4068,N_4876);
xor UO_483 (O_483,N_4752,N_4982);
xnor UO_484 (O_484,N_4980,N_4942);
xnor UO_485 (O_485,N_4139,N_4926);
or UO_486 (O_486,N_4137,N_4630);
nor UO_487 (O_487,N_4642,N_4486);
or UO_488 (O_488,N_4673,N_4945);
nor UO_489 (O_489,N_4802,N_4546);
nand UO_490 (O_490,N_4165,N_4212);
or UO_491 (O_491,N_4213,N_4406);
nor UO_492 (O_492,N_4414,N_4586);
nor UO_493 (O_493,N_4978,N_4324);
and UO_494 (O_494,N_4854,N_4986);
nand UO_495 (O_495,N_4018,N_4445);
nand UO_496 (O_496,N_4856,N_4284);
nand UO_497 (O_497,N_4373,N_4334);
and UO_498 (O_498,N_4161,N_4309);
nor UO_499 (O_499,N_4745,N_4571);
and UO_500 (O_500,N_4395,N_4759);
or UO_501 (O_501,N_4588,N_4895);
and UO_502 (O_502,N_4119,N_4650);
and UO_503 (O_503,N_4677,N_4761);
nor UO_504 (O_504,N_4562,N_4920);
xor UO_505 (O_505,N_4894,N_4999);
and UO_506 (O_506,N_4061,N_4226);
nor UO_507 (O_507,N_4403,N_4871);
or UO_508 (O_508,N_4987,N_4356);
and UO_509 (O_509,N_4873,N_4213);
and UO_510 (O_510,N_4338,N_4925);
and UO_511 (O_511,N_4896,N_4384);
and UO_512 (O_512,N_4302,N_4329);
nand UO_513 (O_513,N_4765,N_4455);
and UO_514 (O_514,N_4079,N_4640);
and UO_515 (O_515,N_4763,N_4363);
and UO_516 (O_516,N_4201,N_4244);
or UO_517 (O_517,N_4222,N_4096);
or UO_518 (O_518,N_4938,N_4743);
or UO_519 (O_519,N_4212,N_4448);
or UO_520 (O_520,N_4189,N_4948);
and UO_521 (O_521,N_4570,N_4168);
nand UO_522 (O_522,N_4623,N_4714);
or UO_523 (O_523,N_4998,N_4442);
or UO_524 (O_524,N_4757,N_4198);
or UO_525 (O_525,N_4162,N_4167);
nor UO_526 (O_526,N_4577,N_4442);
nor UO_527 (O_527,N_4399,N_4019);
and UO_528 (O_528,N_4460,N_4525);
nand UO_529 (O_529,N_4162,N_4497);
or UO_530 (O_530,N_4987,N_4604);
nand UO_531 (O_531,N_4367,N_4699);
or UO_532 (O_532,N_4393,N_4036);
nor UO_533 (O_533,N_4971,N_4129);
or UO_534 (O_534,N_4858,N_4493);
or UO_535 (O_535,N_4212,N_4949);
or UO_536 (O_536,N_4507,N_4432);
nor UO_537 (O_537,N_4975,N_4708);
nor UO_538 (O_538,N_4124,N_4715);
nor UO_539 (O_539,N_4669,N_4515);
nand UO_540 (O_540,N_4070,N_4292);
nand UO_541 (O_541,N_4779,N_4055);
and UO_542 (O_542,N_4012,N_4061);
nand UO_543 (O_543,N_4769,N_4718);
nand UO_544 (O_544,N_4109,N_4801);
and UO_545 (O_545,N_4788,N_4553);
or UO_546 (O_546,N_4112,N_4205);
nor UO_547 (O_547,N_4673,N_4259);
and UO_548 (O_548,N_4699,N_4892);
nor UO_549 (O_549,N_4709,N_4687);
and UO_550 (O_550,N_4046,N_4393);
nor UO_551 (O_551,N_4783,N_4043);
or UO_552 (O_552,N_4486,N_4852);
nor UO_553 (O_553,N_4659,N_4445);
nor UO_554 (O_554,N_4579,N_4524);
and UO_555 (O_555,N_4791,N_4161);
nand UO_556 (O_556,N_4580,N_4081);
nor UO_557 (O_557,N_4078,N_4361);
nand UO_558 (O_558,N_4914,N_4096);
nand UO_559 (O_559,N_4001,N_4346);
nor UO_560 (O_560,N_4455,N_4758);
nor UO_561 (O_561,N_4652,N_4537);
and UO_562 (O_562,N_4637,N_4816);
nand UO_563 (O_563,N_4248,N_4821);
or UO_564 (O_564,N_4506,N_4637);
and UO_565 (O_565,N_4554,N_4861);
nand UO_566 (O_566,N_4899,N_4549);
xor UO_567 (O_567,N_4812,N_4389);
and UO_568 (O_568,N_4995,N_4000);
nor UO_569 (O_569,N_4240,N_4760);
nor UO_570 (O_570,N_4122,N_4914);
nand UO_571 (O_571,N_4633,N_4964);
and UO_572 (O_572,N_4201,N_4600);
xnor UO_573 (O_573,N_4814,N_4957);
nand UO_574 (O_574,N_4435,N_4910);
nand UO_575 (O_575,N_4464,N_4569);
nor UO_576 (O_576,N_4185,N_4601);
xnor UO_577 (O_577,N_4490,N_4760);
nand UO_578 (O_578,N_4904,N_4692);
nor UO_579 (O_579,N_4321,N_4213);
and UO_580 (O_580,N_4015,N_4170);
xor UO_581 (O_581,N_4494,N_4218);
nand UO_582 (O_582,N_4894,N_4403);
xor UO_583 (O_583,N_4484,N_4901);
nand UO_584 (O_584,N_4597,N_4900);
and UO_585 (O_585,N_4732,N_4475);
nand UO_586 (O_586,N_4113,N_4032);
nor UO_587 (O_587,N_4746,N_4173);
and UO_588 (O_588,N_4465,N_4595);
nor UO_589 (O_589,N_4190,N_4209);
and UO_590 (O_590,N_4222,N_4703);
and UO_591 (O_591,N_4614,N_4171);
or UO_592 (O_592,N_4384,N_4381);
and UO_593 (O_593,N_4941,N_4860);
nor UO_594 (O_594,N_4446,N_4409);
nor UO_595 (O_595,N_4310,N_4343);
nor UO_596 (O_596,N_4593,N_4867);
nor UO_597 (O_597,N_4003,N_4096);
nand UO_598 (O_598,N_4431,N_4488);
or UO_599 (O_599,N_4640,N_4785);
and UO_600 (O_600,N_4153,N_4551);
or UO_601 (O_601,N_4710,N_4808);
nand UO_602 (O_602,N_4979,N_4557);
nand UO_603 (O_603,N_4342,N_4267);
nand UO_604 (O_604,N_4532,N_4014);
nor UO_605 (O_605,N_4734,N_4269);
and UO_606 (O_606,N_4412,N_4017);
or UO_607 (O_607,N_4444,N_4709);
xnor UO_608 (O_608,N_4629,N_4617);
xor UO_609 (O_609,N_4867,N_4806);
and UO_610 (O_610,N_4936,N_4202);
nand UO_611 (O_611,N_4744,N_4317);
nor UO_612 (O_612,N_4031,N_4964);
and UO_613 (O_613,N_4500,N_4153);
nand UO_614 (O_614,N_4272,N_4915);
and UO_615 (O_615,N_4938,N_4233);
nor UO_616 (O_616,N_4429,N_4875);
and UO_617 (O_617,N_4784,N_4876);
xor UO_618 (O_618,N_4304,N_4767);
nand UO_619 (O_619,N_4184,N_4747);
nand UO_620 (O_620,N_4995,N_4531);
and UO_621 (O_621,N_4605,N_4877);
xor UO_622 (O_622,N_4735,N_4719);
and UO_623 (O_623,N_4244,N_4702);
or UO_624 (O_624,N_4350,N_4389);
or UO_625 (O_625,N_4589,N_4105);
and UO_626 (O_626,N_4895,N_4763);
nand UO_627 (O_627,N_4915,N_4379);
nand UO_628 (O_628,N_4659,N_4717);
nor UO_629 (O_629,N_4598,N_4640);
nor UO_630 (O_630,N_4812,N_4525);
nand UO_631 (O_631,N_4499,N_4098);
nor UO_632 (O_632,N_4915,N_4885);
or UO_633 (O_633,N_4468,N_4981);
and UO_634 (O_634,N_4112,N_4765);
and UO_635 (O_635,N_4193,N_4734);
or UO_636 (O_636,N_4212,N_4419);
nor UO_637 (O_637,N_4994,N_4190);
and UO_638 (O_638,N_4041,N_4174);
and UO_639 (O_639,N_4228,N_4498);
and UO_640 (O_640,N_4432,N_4370);
or UO_641 (O_641,N_4451,N_4833);
or UO_642 (O_642,N_4293,N_4102);
or UO_643 (O_643,N_4724,N_4230);
nor UO_644 (O_644,N_4915,N_4048);
and UO_645 (O_645,N_4075,N_4395);
nor UO_646 (O_646,N_4079,N_4926);
nor UO_647 (O_647,N_4352,N_4935);
nor UO_648 (O_648,N_4697,N_4719);
nor UO_649 (O_649,N_4938,N_4887);
xnor UO_650 (O_650,N_4623,N_4849);
nor UO_651 (O_651,N_4105,N_4645);
nor UO_652 (O_652,N_4507,N_4844);
xor UO_653 (O_653,N_4654,N_4632);
or UO_654 (O_654,N_4719,N_4431);
and UO_655 (O_655,N_4947,N_4089);
or UO_656 (O_656,N_4566,N_4961);
nand UO_657 (O_657,N_4779,N_4010);
nand UO_658 (O_658,N_4598,N_4309);
and UO_659 (O_659,N_4584,N_4931);
xnor UO_660 (O_660,N_4532,N_4701);
xor UO_661 (O_661,N_4581,N_4275);
xnor UO_662 (O_662,N_4248,N_4772);
xor UO_663 (O_663,N_4435,N_4574);
or UO_664 (O_664,N_4996,N_4052);
or UO_665 (O_665,N_4439,N_4028);
or UO_666 (O_666,N_4582,N_4564);
and UO_667 (O_667,N_4640,N_4344);
nand UO_668 (O_668,N_4498,N_4892);
and UO_669 (O_669,N_4303,N_4489);
nor UO_670 (O_670,N_4745,N_4875);
xnor UO_671 (O_671,N_4972,N_4319);
or UO_672 (O_672,N_4748,N_4226);
nand UO_673 (O_673,N_4692,N_4728);
or UO_674 (O_674,N_4961,N_4652);
and UO_675 (O_675,N_4957,N_4850);
xor UO_676 (O_676,N_4695,N_4456);
nand UO_677 (O_677,N_4258,N_4120);
and UO_678 (O_678,N_4232,N_4531);
xnor UO_679 (O_679,N_4491,N_4723);
nand UO_680 (O_680,N_4084,N_4794);
nand UO_681 (O_681,N_4299,N_4144);
nand UO_682 (O_682,N_4804,N_4385);
nor UO_683 (O_683,N_4448,N_4813);
nor UO_684 (O_684,N_4969,N_4718);
and UO_685 (O_685,N_4288,N_4244);
nand UO_686 (O_686,N_4484,N_4370);
or UO_687 (O_687,N_4119,N_4847);
or UO_688 (O_688,N_4442,N_4864);
or UO_689 (O_689,N_4082,N_4309);
nor UO_690 (O_690,N_4215,N_4181);
and UO_691 (O_691,N_4092,N_4951);
or UO_692 (O_692,N_4808,N_4884);
nand UO_693 (O_693,N_4562,N_4733);
or UO_694 (O_694,N_4403,N_4127);
nor UO_695 (O_695,N_4915,N_4847);
or UO_696 (O_696,N_4108,N_4521);
and UO_697 (O_697,N_4323,N_4201);
and UO_698 (O_698,N_4240,N_4666);
nor UO_699 (O_699,N_4962,N_4353);
nor UO_700 (O_700,N_4444,N_4488);
nor UO_701 (O_701,N_4681,N_4659);
xnor UO_702 (O_702,N_4229,N_4837);
or UO_703 (O_703,N_4568,N_4709);
or UO_704 (O_704,N_4408,N_4233);
and UO_705 (O_705,N_4070,N_4297);
or UO_706 (O_706,N_4177,N_4294);
or UO_707 (O_707,N_4816,N_4416);
nand UO_708 (O_708,N_4250,N_4394);
or UO_709 (O_709,N_4609,N_4810);
nor UO_710 (O_710,N_4943,N_4828);
nor UO_711 (O_711,N_4396,N_4738);
nand UO_712 (O_712,N_4664,N_4123);
nor UO_713 (O_713,N_4137,N_4754);
or UO_714 (O_714,N_4560,N_4501);
nor UO_715 (O_715,N_4435,N_4449);
and UO_716 (O_716,N_4391,N_4879);
and UO_717 (O_717,N_4458,N_4991);
nor UO_718 (O_718,N_4683,N_4122);
nor UO_719 (O_719,N_4521,N_4947);
nor UO_720 (O_720,N_4552,N_4873);
or UO_721 (O_721,N_4969,N_4705);
nand UO_722 (O_722,N_4717,N_4826);
xor UO_723 (O_723,N_4978,N_4721);
nand UO_724 (O_724,N_4528,N_4329);
nand UO_725 (O_725,N_4951,N_4361);
nor UO_726 (O_726,N_4679,N_4467);
and UO_727 (O_727,N_4241,N_4206);
or UO_728 (O_728,N_4672,N_4619);
and UO_729 (O_729,N_4665,N_4697);
xor UO_730 (O_730,N_4793,N_4353);
xnor UO_731 (O_731,N_4372,N_4776);
and UO_732 (O_732,N_4429,N_4631);
nor UO_733 (O_733,N_4149,N_4581);
or UO_734 (O_734,N_4892,N_4055);
xnor UO_735 (O_735,N_4274,N_4603);
and UO_736 (O_736,N_4245,N_4023);
and UO_737 (O_737,N_4234,N_4644);
and UO_738 (O_738,N_4010,N_4093);
or UO_739 (O_739,N_4660,N_4653);
or UO_740 (O_740,N_4065,N_4184);
or UO_741 (O_741,N_4916,N_4794);
and UO_742 (O_742,N_4424,N_4392);
nand UO_743 (O_743,N_4030,N_4803);
xor UO_744 (O_744,N_4064,N_4622);
and UO_745 (O_745,N_4720,N_4216);
and UO_746 (O_746,N_4045,N_4590);
nand UO_747 (O_747,N_4380,N_4302);
and UO_748 (O_748,N_4872,N_4873);
nand UO_749 (O_749,N_4757,N_4544);
nor UO_750 (O_750,N_4701,N_4590);
nand UO_751 (O_751,N_4414,N_4885);
nand UO_752 (O_752,N_4262,N_4736);
nor UO_753 (O_753,N_4853,N_4622);
nand UO_754 (O_754,N_4097,N_4648);
nand UO_755 (O_755,N_4677,N_4927);
and UO_756 (O_756,N_4539,N_4063);
and UO_757 (O_757,N_4020,N_4291);
and UO_758 (O_758,N_4472,N_4361);
or UO_759 (O_759,N_4915,N_4452);
or UO_760 (O_760,N_4146,N_4122);
nor UO_761 (O_761,N_4317,N_4197);
or UO_762 (O_762,N_4313,N_4813);
nand UO_763 (O_763,N_4117,N_4676);
or UO_764 (O_764,N_4810,N_4243);
nor UO_765 (O_765,N_4135,N_4478);
and UO_766 (O_766,N_4587,N_4830);
and UO_767 (O_767,N_4036,N_4215);
nor UO_768 (O_768,N_4318,N_4170);
nand UO_769 (O_769,N_4786,N_4381);
nor UO_770 (O_770,N_4016,N_4362);
nor UO_771 (O_771,N_4401,N_4721);
and UO_772 (O_772,N_4449,N_4077);
or UO_773 (O_773,N_4368,N_4853);
xnor UO_774 (O_774,N_4866,N_4429);
nor UO_775 (O_775,N_4611,N_4701);
nand UO_776 (O_776,N_4846,N_4265);
and UO_777 (O_777,N_4637,N_4930);
or UO_778 (O_778,N_4320,N_4053);
nor UO_779 (O_779,N_4855,N_4391);
nand UO_780 (O_780,N_4118,N_4562);
and UO_781 (O_781,N_4402,N_4114);
nor UO_782 (O_782,N_4847,N_4843);
nand UO_783 (O_783,N_4634,N_4943);
nand UO_784 (O_784,N_4332,N_4686);
nor UO_785 (O_785,N_4677,N_4097);
xor UO_786 (O_786,N_4830,N_4450);
or UO_787 (O_787,N_4940,N_4682);
nor UO_788 (O_788,N_4894,N_4760);
nor UO_789 (O_789,N_4439,N_4876);
nand UO_790 (O_790,N_4893,N_4912);
nand UO_791 (O_791,N_4235,N_4787);
or UO_792 (O_792,N_4882,N_4717);
xnor UO_793 (O_793,N_4294,N_4686);
and UO_794 (O_794,N_4626,N_4942);
or UO_795 (O_795,N_4908,N_4795);
or UO_796 (O_796,N_4138,N_4443);
and UO_797 (O_797,N_4424,N_4622);
and UO_798 (O_798,N_4800,N_4552);
or UO_799 (O_799,N_4967,N_4339);
and UO_800 (O_800,N_4167,N_4164);
or UO_801 (O_801,N_4909,N_4693);
nor UO_802 (O_802,N_4449,N_4148);
nor UO_803 (O_803,N_4073,N_4449);
nand UO_804 (O_804,N_4876,N_4176);
nor UO_805 (O_805,N_4181,N_4140);
nor UO_806 (O_806,N_4404,N_4073);
nor UO_807 (O_807,N_4112,N_4886);
and UO_808 (O_808,N_4350,N_4453);
and UO_809 (O_809,N_4930,N_4661);
and UO_810 (O_810,N_4228,N_4127);
nand UO_811 (O_811,N_4048,N_4255);
or UO_812 (O_812,N_4722,N_4270);
nand UO_813 (O_813,N_4265,N_4739);
or UO_814 (O_814,N_4377,N_4870);
nand UO_815 (O_815,N_4746,N_4335);
nand UO_816 (O_816,N_4029,N_4396);
and UO_817 (O_817,N_4675,N_4699);
nor UO_818 (O_818,N_4319,N_4470);
and UO_819 (O_819,N_4970,N_4469);
nor UO_820 (O_820,N_4111,N_4261);
nand UO_821 (O_821,N_4730,N_4997);
nand UO_822 (O_822,N_4091,N_4220);
nor UO_823 (O_823,N_4980,N_4197);
nor UO_824 (O_824,N_4431,N_4453);
nor UO_825 (O_825,N_4528,N_4273);
or UO_826 (O_826,N_4145,N_4562);
or UO_827 (O_827,N_4563,N_4633);
nor UO_828 (O_828,N_4678,N_4461);
nor UO_829 (O_829,N_4722,N_4811);
or UO_830 (O_830,N_4191,N_4184);
nor UO_831 (O_831,N_4011,N_4134);
nand UO_832 (O_832,N_4293,N_4313);
nand UO_833 (O_833,N_4163,N_4962);
or UO_834 (O_834,N_4960,N_4722);
and UO_835 (O_835,N_4396,N_4850);
or UO_836 (O_836,N_4401,N_4408);
nor UO_837 (O_837,N_4989,N_4547);
and UO_838 (O_838,N_4507,N_4978);
xnor UO_839 (O_839,N_4106,N_4395);
nor UO_840 (O_840,N_4423,N_4089);
and UO_841 (O_841,N_4964,N_4962);
or UO_842 (O_842,N_4419,N_4555);
xnor UO_843 (O_843,N_4671,N_4163);
nor UO_844 (O_844,N_4958,N_4945);
nor UO_845 (O_845,N_4299,N_4791);
or UO_846 (O_846,N_4665,N_4357);
nand UO_847 (O_847,N_4008,N_4196);
or UO_848 (O_848,N_4078,N_4055);
or UO_849 (O_849,N_4656,N_4985);
or UO_850 (O_850,N_4129,N_4791);
or UO_851 (O_851,N_4014,N_4293);
or UO_852 (O_852,N_4508,N_4455);
or UO_853 (O_853,N_4576,N_4690);
and UO_854 (O_854,N_4464,N_4113);
and UO_855 (O_855,N_4636,N_4832);
or UO_856 (O_856,N_4200,N_4151);
or UO_857 (O_857,N_4823,N_4694);
nor UO_858 (O_858,N_4379,N_4436);
xor UO_859 (O_859,N_4507,N_4527);
or UO_860 (O_860,N_4179,N_4623);
xor UO_861 (O_861,N_4718,N_4382);
and UO_862 (O_862,N_4393,N_4859);
and UO_863 (O_863,N_4844,N_4112);
or UO_864 (O_864,N_4924,N_4917);
xnor UO_865 (O_865,N_4912,N_4933);
nor UO_866 (O_866,N_4901,N_4146);
nand UO_867 (O_867,N_4748,N_4309);
and UO_868 (O_868,N_4006,N_4880);
and UO_869 (O_869,N_4617,N_4389);
nor UO_870 (O_870,N_4623,N_4071);
and UO_871 (O_871,N_4849,N_4240);
xnor UO_872 (O_872,N_4869,N_4164);
nand UO_873 (O_873,N_4054,N_4977);
nand UO_874 (O_874,N_4597,N_4572);
or UO_875 (O_875,N_4690,N_4404);
nor UO_876 (O_876,N_4374,N_4632);
nand UO_877 (O_877,N_4711,N_4158);
xor UO_878 (O_878,N_4444,N_4254);
or UO_879 (O_879,N_4512,N_4739);
nand UO_880 (O_880,N_4028,N_4106);
nor UO_881 (O_881,N_4086,N_4189);
and UO_882 (O_882,N_4272,N_4329);
and UO_883 (O_883,N_4240,N_4665);
or UO_884 (O_884,N_4504,N_4315);
xnor UO_885 (O_885,N_4376,N_4749);
nor UO_886 (O_886,N_4302,N_4273);
and UO_887 (O_887,N_4177,N_4015);
or UO_888 (O_888,N_4233,N_4587);
and UO_889 (O_889,N_4200,N_4597);
nand UO_890 (O_890,N_4105,N_4485);
nor UO_891 (O_891,N_4229,N_4581);
nand UO_892 (O_892,N_4965,N_4572);
xor UO_893 (O_893,N_4737,N_4700);
and UO_894 (O_894,N_4831,N_4474);
xor UO_895 (O_895,N_4019,N_4115);
and UO_896 (O_896,N_4133,N_4883);
nand UO_897 (O_897,N_4618,N_4067);
or UO_898 (O_898,N_4748,N_4069);
and UO_899 (O_899,N_4008,N_4241);
nor UO_900 (O_900,N_4151,N_4589);
or UO_901 (O_901,N_4624,N_4346);
nor UO_902 (O_902,N_4441,N_4701);
and UO_903 (O_903,N_4844,N_4624);
nor UO_904 (O_904,N_4908,N_4837);
nand UO_905 (O_905,N_4706,N_4508);
nand UO_906 (O_906,N_4132,N_4285);
and UO_907 (O_907,N_4434,N_4115);
or UO_908 (O_908,N_4436,N_4977);
or UO_909 (O_909,N_4102,N_4462);
nor UO_910 (O_910,N_4989,N_4636);
nand UO_911 (O_911,N_4375,N_4674);
nor UO_912 (O_912,N_4726,N_4300);
nand UO_913 (O_913,N_4103,N_4003);
nor UO_914 (O_914,N_4467,N_4219);
xor UO_915 (O_915,N_4707,N_4909);
nor UO_916 (O_916,N_4735,N_4770);
or UO_917 (O_917,N_4541,N_4218);
or UO_918 (O_918,N_4788,N_4192);
and UO_919 (O_919,N_4514,N_4245);
and UO_920 (O_920,N_4194,N_4340);
nand UO_921 (O_921,N_4676,N_4661);
nor UO_922 (O_922,N_4373,N_4196);
and UO_923 (O_923,N_4793,N_4489);
nand UO_924 (O_924,N_4343,N_4559);
nand UO_925 (O_925,N_4582,N_4291);
nor UO_926 (O_926,N_4405,N_4816);
nand UO_927 (O_927,N_4663,N_4800);
xor UO_928 (O_928,N_4310,N_4348);
nor UO_929 (O_929,N_4521,N_4265);
nor UO_930 (O_930,N_4735,N_4242);
or UO_931 (O_931,N_4745,N_4162);
nand UO_932 (O_932,N_4408,N_4333);
xnor UO_933 (O_933,N_4081,N_4002);
or UO_934 (O_934,N_4859,N_4416);
and UO_935 (O_935,N_4038,N_4012);
and UO_936 (O_936,N_4318,N_4866);
and UO_937 (O_937,N_4329,N_4095);
and UO_938 (O_938,N_4701,N_4040);
and UO_939 (O_939,N_4883,N_4209);
and UO_940 (O_940,N_4682,N_4767);
nor UO_941 (O_941,N_4086,N_4462);
xor UO_942 (O_942,N_4269,N_4319);
nand UO_943 (O_943,N_4972,N_4988);
or UO_944 (O_944,N_4366,N_4913);
nand UO_945 (O_945,N_4549,N_4389);
nor UO_946 (O_946,N_4960,N_4275);
nand UO_947 (O_947,N_4450,N_4716);
nor UO_948 (O_948,N_4975,N_4122);
nand UO_949 (O_949,N_4009,N_4158);
and UO_950 (O_950,N_4727,N_4387);
nor UO_951 (O_951,N_4905,N_4890);
or UO_952 (O_952,N_4797,N_4538);
nand UO_953 (O_953,N_4904,N_4640);
or UO_954 (O_954,N_4874,N_4689);
and UO_955 (O_955,N_4352,N_4096);
nor UO_956 (O_956,N_4982,N_4976);
xnor UO_957 (O_957,N_4164,N_4497);
and UO_958 (O_958,N_4156,N_4719);
or UO_959 (O_959,N_4373,N_4848);
nand UO_960 (O_960,N_4426,N_4330);
nand UO_961 (O_961,N_4779,N_4047);
and UO_962 (O_962,N_4152,N_4717);
or UO_963 (O_963,N_4959,N_4077);
nand UO_964 (O_964,N_4409,N_4299);
nor UO_965 (O_965,N_4589,N_4549);
or UO_966 (O_966,N_4881,N_4333);
and UO_967 (O_967,N_4317,N_4161);
and UO_968 (O_968,N_4430,N_4662);
xor UO_969 (O_969,N_4943,N_4378);
or UO_970 (O_970,N_4766,N_4910);
nand UO_971 (O_971,N_4871,N_4468);
nor UO_972 (O_972,N_4610,N_4781);
nand UO_973 (O_973,N_4995,N_4306);
and UO_974 (O_974,N_4505,N_4063);
and UO_975 (O_975,N_4905,N_4549);
nand UO_976 (O_976,N_4428,N_4074);
xor UO_977 (O_977,N_4925,N_4727);
or UO_978 (O_978,N_4380,N_4881);
or UO_979 (O_979,N_4908,N_4070);
nor UO_980 (O_980,N_4064,N_4868);
nor UO_981 (O_981,N_4999,N_4573);
nand UO_982 (O_982,N_4919,N_4814);
xnor UO_983 (O_983,N_4335,N_4206);
nor UO_984 (O_984,N_4850,N_4822);
and UO_985 (O_985,N_4236,N_4369);
and UO_986 (O_986,N_4008,N_4023);
nor UO_987 (O_987,N_4687,N_4324);
and UO_988 (O_988,N_4122,N_4283);
or UO_989 (O_989,N_4003,N_4924);
or UO_990 (O_990,N_4553,N_4350);
nor UO_991 (O_991,N_4870,N_4723);
nor UO_992 (O_992,N_4223,N_4418);
and UO_993 (O_993,N_4125,N_4233);
and UO_994 (O_994,N_4714,N_4961);
nor UO_995 (O_995,N_4457,N_4535);
or UO_996 (O_996,N_4070,N_4366);
nor UO_997 (O_997,N_4773,N_4717);
nor UO_998 (O_998,N_4075,N_4410);
or UO_999 (O_999,N_4738,N_4812);
endmodule