module basic_750_5000_1000_2_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2544,N_2545,N_2546,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2557,N_2560,N_2562,N_2563,N_2564,N_2565,N_2567,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2577,N_2578,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2604,N_2605,N_2606,N_2608,N_2609,N_2610,N_2612,N_2613,N_2614,N_2615,N_2617,N_2618,N_2620,N_2622,N_2623,N_2624,N_2625,N_2626,N_2628,N_2629,N_2630,N_2632,N_2633,N_2634,N_2635,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2647,N_2648,N_2649,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2661,N_2662,N_2663,N_2664,N_2666,N_2667,N_2669,N_2670,N_2671,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2682,N_2683,N_2684,N_2685,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2696,N_2697,N_2698,N_2699,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2719,N_2720,N_2721,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2733,N_2735,N_2736,N_2739,N_2740,N_2742,N_2743,N_2745,N_2746,N_2748,N_2749,N_2750,N_2751,N_2753,N_2755,N_2757,N_2758,N_2759,N_2760,N_2761,N_2763,N_2764,N_2766,N_2767,N_2768,N_2769,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2791,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2809,N_2810,N_2812,N_2813,N_2814,N_2815,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2834,N_2835,N_2836,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2858,N_2859,N_2860,N_2861,N_2862,N_2864,N_2865,N_2867,N_2868,N_2869,N_2871,N_2873,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2891,N_2892,N_2893,N_2896,N_2897,N_2899,N_2900,N_2901,N_2904,N_2905,N_2906,N_2907,N_2908,N_2910,N_2911,N_2912,N_2913,N_2915,N_2916,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2942,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2957,N_2959,N_2960,N_2961,N_2962,N_2964,N_2965,N_2966,N_2967,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2980,N_2982,N_2983,N_2984,N_2986,N_2987,N_2989,N_2990,N_2991,N_2993,N_2994,N_2995,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3006,N_3007,N_3009,N_3011,N_3012,N_3013,N_3014,N_3016,N_3018,N_3019,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3034,N_3036,N_3038,N_3039,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3097,N_3098,N_3099,N_3100,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3115,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3125,N_3126,N_3127,N_3128,N_3130,N_3131,N_3132,N_3133,N_3134,N_3136,N_3138,N_3140,N_3141,N_3142,N_3144,N_3145,N_3146,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3176,N_3177,N_3178,N_3180,N_3181,N_3182,N_3183,N_3185,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3206,N_3208,N_3209,N_3210,N_3212,N_3213,N_3214,N_3215,N_3216,N_3218,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3229,N_3230,N_3231,N_3232,N_3233,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3243,N_3245,N_3246,N_3247,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3273,N_3274,N_3275,N_3276,N_3277,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3325,N_3326,N_3327,N_3328,N_3329,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3357,N_3358,N_3362,N_3363,N_3364,N_3365,N_3366,N_3368,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3381,N_3384,N_3386,N_3387,N_3388,N_3389,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3409,N_3410,N_3411,N_3412,N_3414,N_3415,N_3416,N_3417,N_3419,N_3420,N_3421,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3434,N_3435,N_3436,N_3437,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3449,N_3450,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3459,N_3461,N_3462,N_3463,N_3466,N_3467,N_3468,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3481,N_3482,N_3483,N_3485,N_3487,N_3488,N_3490,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3511,N_3512,N_3514,N_3515,N_3517,N_3519,N_3520,N_3521,N_3523,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3532,N_3534,N_3535,N_3536,N_3537,N_3539,N_3540,N_3541,N_3543,N_3544,N_3546,N_3547,N_3548,N_3549,N_3551,N_3552,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3604,N_3605,N_3606,N_3610,N_3612,N_3613,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3623,N_3624,N_3625,N_3628,N_3629,N_3630,N_3632,N_3633,N_3634,N_3635,N_3636,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3664,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3674,N_3676,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3706,N_3707,N_3708,N_3709,N_3710,N_3712,N_3713,N_3714,N_3715,N_3717,N_3718,N_3719,N_3721,N_3722,N_3723,N_3724,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3734,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3752,N_3753,N_3754,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3768,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3783,N_3784,N_3785,N_3786,N_3788,N_3789,N_3791,N_3792,N_3793,N_3795,N_3797,N_3798,N_3801,N_3802,N_3804,N_3807,N_3808,N_3809,N_3810,N_3812,N_3813,N_3814,N_3816,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3829,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3841,N_3842,N_3844,N_3845,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3859,N_3861,N_3863,N_3864,N_3866,N_3867,N_3868,N_3870,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3892,N_3893,N_3894,N_3896,N_3897,N_3900,N_3903,N_3904,N_3907,N_3908,N_3909,N_3911,N_3912,N_3913,N_3914,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3926,N_3927,N_3928,N_3929,N_3930,N_3932,N_3933,N_3935,N_3936,N_3937,N_3938,N_3940,N_3941,N_3942,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3960,N_3962,N_3963,N_3964,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3977,N_3978,N_3979,N_3980,N_3983,N_3985,N_3987,N_3988,N_3990,N_3992,N_3993,N_3994,N_3995,N_3996,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4021,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4033,N_4034,N_4035,N_4036,N_4038,N_4039,N_4043,N_4045,N_4046,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4057,N_4058,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4068,N_4069,N_4070,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4084,N_4085,N_4087,N_4088,N_4089,N_4090,N_4091,N_4094,N_4095,N_4097,N_4098,N_4103,N_4104,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4113,N_4114,N_4117,N_4118,N_4120,N_4121,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4133,N_4134,N_4135,N_4136,N_4139,N_4140,N_4141,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4152,N_4153,N_4154,N_4156,N_4157,N_4158,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4167,N_4168,N_4169,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4183,N_4185,N_4186,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4196,N_4198,N_4199,N_4200,N_4202,N_4203,N_4205,N_4206,N_4207,N_4208,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4219,N_4221,N_4223,N_4224,N_4225,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4242,N_4244,N_4245,N_4246,N_4248,N_4249,N_4250,N_4251,N_4252,N_4254,N_4255,N_4256,N_4257,N_4258,N_4260,N_4261,N_4262,N_4263,N_4264,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4289,N_4291,N_4292,N_4294,N_4295,N_4296,N_4297,N_4299,N_4302,N_4304,N_4306,N_4309,N_4310,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4319,N_4321,N_4322,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4335,N_4336,N_4338,N_4339,N_4340,N_4341,N_4342,N_4344,N_4345,N_4346,N_4347,N_4348,N_4350,N_4351,N_4352,N_4354,N_4355,N_4356,N_4357,N_4358,N_4360,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4391,N_4392,N_4393,N_4394,N_4395,N_4397,N_4399,N_4401,N_4402,N_4405,N_4406,N_4407,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4459,N_4462,N_4463,N_4464,N_4466,N_4467,N_4468,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4481,N_4482,N_4483,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4527,N_4528,N_4529,N_4532,N_4533,N_4534,N_4535,N_4537,N_4538,N_4539,N_4540,N_4543,N_4544,N_4545,N_4546,N_4548,N_4549,N_4550,N_4551,N_4552,N_4554,N_4555,N_4556,N_4557,N_4558,N_4561,N_4562,N_4563,N_4565,N_4568,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4592,N_4593,N_4594,N_4595,N_4598,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4608,N_4609,N_4610,N_4611,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4634,N_4635,N_4636,N_4637,N_4640,N_4641,N_4642,N_4643,N_4645,N_4647,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4680,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4701,N_4702,N_4703,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4717,N_4719,N_4720,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4736,N_4737,N_4741,N_4742,N_4744,N_4746,N_4747,N_4748,N_4749,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4760,N_4761,N_4762,N_4763,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4777,N_4778,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4787,N_4788,N_4790,N_4791,N_4792,N_4793,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4809,N_4812,N_4813,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4823,N_4824,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4857,N_4859,N_4860,N_4862,N_4863,N_4865,N_4866,N_4868,N_4869,N_4870,N_4874,N_4875,N_4876,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4890,N_4891,N_4892,N_4894,N_4895,N_4896,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4907,N_4908,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4922,N_4924,N_4925,N_4927,N_4928,N_4929,N_4931,N_4933,N_4935,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4966,N_4967,N_4968,N_4970,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4990,N_4991,N_4992,N_4993,N_4994,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_683,In_572);
or U1 (N_1,In_33,In_580);
xnor U2 (N_2,In_309,In_460);
xor U3 (N_3,In_590,In_449);
nand U4 (N_4,In_584,In_414);
and U5 (N_5,In_600,In_227);
nand U6 (N_6,In_209,In_125);
or U7 (N_7,In_696,In_51);
nand U8 (N_8,In_338,In_684);
nor U9 (N_9,In_477,In_439);
and U10 (N_10,In_559,In_496);
xor U11 (N_11,In_435,In_129);
nand U12 (N_12,In_14,In_42);
nor U13 (N_13,In_10,In_647);
nand U14 (N_14,In_365,In_77);
nor U15 (N_15,In_485,In_26);
and U16 (N_16,In_398,In_339);
xor U17 (N_17,In_52,In_143);
and U18 (N_18,In_631,In_470);
or U19 (N_19,In_680,In_709);
nand U20 (N_20,In_259,In_434);
and U21 (N_21,In_220,In_640);
or U22 (N_22,In_617,In_746);
nor U23 (N_23,In_603,In_598);
nor U24 (N_24,In_351,In_69);
and U25 (N_25,In_423,In_728);
or U26 (N_26,In_330,In_94);
nand U27 (N_27,In_137,In_250);
nor U28 (N_28,In_587,In_501);
and U29 (N_29,In_233,In_614);
nor U30 (N_30,In_539,In_433);
xor U31 (N_31,In_370,In_86);
nand U32 (N_32,In_208,In_245);
and U33 (N_33,In_326,In_97);
and U34 (N_34,In_113,In_353);
nand U35 (N_35,In_57,In_312);
nor U36 (N_36,In_126,In_482);
nor U37 (N_37,In_384,In_716);
nand U38 (N_38,In_185,In_318);
nand U39 (N_39,In_672,In_576);
or U40 (N_40,In_413,In_355);
nand U41 (N_41,In_715,In_379);
or U42 (N_42,In_290,In_387);
or U43 (N_43,In_668,In_34);
xor U44 (N_44,In_275,In_521);
nand U45 (N_45,In_381,In_236);
and U46 (N_46,In_497,In_720);
and U47 (N_47,In_8,In_687);
nor U48 (N_48,In_217,In_76);
xor U49 (N_49,In_690,In_3);
xor U50 (N_50,In_335,In_622);
or U51 (N_51,In_131,In_360);
nor U52 (N_52,In_356,In_652);
nand U53 (N_53,In_404,In_239);
nor U54 (N_54,In_23,In_135);
nor U55 (N_55,In_21,In_729);
or U56 (N_56,In_29,In_20);
or U57 (N_57,In_128,In_701);
and U58 (N_58,In_577,In_402);
and U59 (N_59,In_134,In_643);
or U60 (N_60,In_509,In_327);
or U61 (N_61,In_679,In_124);
or U62 (N_62,In_105,In_218);
nand U63 (N_63,In_475,In_139);
and U64 (N_64,In_197,In_726);
or U65 (N_65,In_349,In_582);
nor U66 (N_66,In_513,In_568);
xnor U67 (N_67,In_85,In_297);
and U68 (N_68,In_249,In_558);
or U69 (N_69,In_575,In_657);
and U70 (N_70,In_455,In_594);
nor U71 (N_71,In_606,In_0);
nor U72 (N_72,In_548,In_141);
nor U73 (N_73,In_291,In_146);
and U74 (N_74,In_171,In_114);
and U75 (N_75,In_697,In_664);
nor U76 (N_76,In_397,In_224);
and U77 (N_77,In_240,In_495);
or U78 (N_78,In_39,In_302);
or U79 (N_79,In_13,In_260);
or U80 (N_80,In_706,In_656);
or U81 (N_81,In_90,In_537);
and U82 (N_82,In_295,In_120);
xor U83 (N_83,In_107,In_691);
or U84 (N_84,In_130,In_517);
nand U85 (N_85,In_655,In_713);
xor U86 (N_86,In_148,In_694);
or U87 (N_87,In_2,In_545);
or U88 (N_88,In_632,In_203);
or U89 (N_89,In_747,In_6);
or U90 (N_90,In_454,In_425);
nand U91 (N_91,In_740,In_328);
and U92 (N_92,In_358,In_98);
and U93 (N_93,In_563,In_415);
xnor U94 (N_94,In_686,In_95);
nor U95 (N_95,In_262,In_286);
nand U96 (N_96,In_314,In_391);
nand U97 (N_97,In_653,In_47);
and U98 (N_98,In_738,In_93);
xnor U99 (N_99,In_458,In_462);
or U100 (N_100,In_255,In_348);
and U101 (N_101,In_408,In_183);
and U102 (N_102,In_204,In_735);
xnor U103 (N_103,In_639,In_463);
and U104 (N_104,In_182,In_89);
and U105 (N_105,In_287,In_553);
or U106 (N_106,In_111,In_361);
or U107 (N_107,In_333,In_368);
and U108 (N_108,In_170,In_91);
and U109 (N_109,In_46,In_7);
nand U110 (N_110,In_303,In_396);
and U111 (N_111,In_426,In_292);
and U112 (N_112,In_212,In_147);
and U113 (N_113,In_494,In_607);
and U114 (N_114,In_734,In_608);
and U115 (N_115,In_564,In_25);
or U116 (N_116,In_591,In_18);
nand U117 (N_117,In_116,In_191);
and U118 (N_118,In_741,In_79);
nand U119 (N_119,In_108,In_123);
nand U120 (N_120,In_538,In_445);
xor U121 (N_121,In_403,In_298);
xor U122 (N_122,In_346,In_133);
and U123 (N_123,In_164,In_669);
nand U124 (N_124,In_595,In_12);
xnor U125 (N_125,In_241,In_343);
xor U126 (N_126,In_390,In_311);
nor U127 (N_127,In_596,In_48);
and U128 (N_128,In_407,In_82);
nor U129 (N_129,In_464,In_480);
nand U130 (N_130,In_552,In_288);
nand U131 (N_131,In_22,In_385);
nor U132 (N_132,In_196,In_556);
and U133 (N_133,In_99,In_161);
nor U134 (N_134,In_58,In_670);
and U135 (N_135,In_362,In_665);
or U136 (N_136,In_394,In_188);
or U137 (N_137,In_38,In_267);
nand U138 (N_138,In_447,In_533);
and U139 (N_139,In_499,In_375);
nor U140 (N_140,In_49,In_525);
or U141 (N_141,In_602,In_535);
and U142 (N_142,In_543,In_507);
or U143 (N_143,In_221,In_200);
and U144 (N_144,In_635,In_467);
nand U145 (N_145,In_616,In_673);
and U146 (N_146,In_417,In_276);
xnor U147 (N_147,In_44,In_341);
nor U148 (N_148,In_121,In_562);
nor U149 (N_149,In_392,In_40);
nor U150 (N_150,In_555,In_549);
and U151 (N_151,In_410,In_293);
xor U152 (N_152,In_702,In_367);
nand U153 (N_153,In_536,In_674);
xor U154 (N_154,In_307,In_363);
nor U155 (N_155,In_748,In_41);
nor U156 (N_156,In_393,In_416);
nor U157 (N_157,In_605,In_83);
and U158 (N_158,In_246,In_366);
and U159 (N_159,In_187,In_624);
nand U160 (N_160,In_714,In_479);
and U161 (N_161,In_345,In_725);
nor U162 (N_162,In_660,In_65);
nor U163 (N_163,In_154,In_322);
nand U164 (N_164,In_5,In_736);
xor U165 (N_165,In_461,In_332);
xor U166 (N_166,In_519,In_440);
nor U167 (N_167,In_510,In_55);
nor U168 (N_168,In_263,In_723);
nor U169 (N_169,In_283,In_560);
nor U170 (N_170,In_374,In_274);
nand U171 (N_171,In_109,In_618);
and U172 (N_172,In_15,In_305);
xor U173 (N_173,In_75,In_707);
nand U174 (N_174,In_427,In_437);
nand U175 (N_175,In_554,In_579);
and U176 (N_176,In_269,In_127);
nor U177 (N_177,In_68,In_167);
nor U178 (N_178,In_593,In_638);
and U179 (N_179,In_35,In_621);
and U180 (N_180,In_428,In_304);
nand U181 (N_181,In_251,In_421);
or U182 (N_182,In_484,In_371);
and U183 (N_183,In_72,In_406);
nor U184 (N_184,In_486,In_31);
xnor U185 (N_185,In_248,In_103);
or U186 (N_186,In_228,In_145);
or U187 (N_187,In_630,In_438);
nand U188 (N_188,In_611,In_60);
or U189 (N_189,In_92,In_277);
nor U190 (N_190,In_490,In_237);
xnor U191 (N_191,In_78,In_468);
or U192 (N_192,In_722,In_692);
nand U193 (N_193,In_500,In_420);
or U194 (N_194,In_573,In_229);
or U195 (N_195,In_289,In_336);
or U196 (N_196,In_599,In_636);
nor U197 (N_197,In_739,In_294);
and U198 (N_198,In_699,In_117);
or U199 (N_199,In_169,In_551);
nand U200 (N_200,In_529,In_411);
and U201 (N_201,In_742,In_62);
and U202 (N_202,In_613,In_192);
nor U203 (N_203,In_432,In_645);
and U204 (N_204,In_194,In_281);
or U205 (N_205,In_659,In_162);
nand U206 (N_206,In_676,In_493);
or U207 (N_207,In_321,In_210);
nand U208 (N_208,In_395,In_571);
nor U209 (N_209,In_610,In_745);
nor U210 (N_210,In_628,In_705);
or U211 (N_211,In_373,In_347);
or U212 (N_212,In_100,In_708);
and U213 (N_213,In_476,In_419);
or U214 (N_214,In_81,In_405);
xor U215 (N_215,In_544,In_733);
nand U216 (N_216,In_442,In_483);
or U217 (N_217,In_173,In_585);
or U218 (N_218,In_342,In_1);
nor U219 (N_219,In_534,In_527);
nor U220 (N_220,In_430,In_202);
and U221 (N_221,In_518,In_504);
and U222 (N_222,In_258,In_119);
nor U223 (N_223,In_743,In_542);
or U224 (N_224,In_324,In_214);
or U225 (N_225,In_418,In_567);
nand U226 (N_226,In_565,In_50);
nand U227 (N_227,In_609,In_446);
nor U228 (N_228,In_524,In_666);
nor U229 (N_229,In_727,In_400);
nand U230 (N_230,In_63,In_222);
nand U231 (N_231,In_43,In_383);
and U232 (N_232,In_531,In_234);
and U233 (N_233,In_732,In_369);
xor U234 (N_234,In_152,In_264);
xnor U235 (N_235,In_308,In_457);
and U236 (N_236,In_282,In_583);
and U237 (N_237,In_118,In_189);
or U238 (N_238,In_681,In_329);
and U239 (N_239,In_195,In_11);
nand U240 (N_240,In_487,In_731);
xor U241 (N_241,In_151,In_646);
or U242 (N_242,In_71,In_488);
nor U243 (N_243,In_516,In_604);
nor U244 (N_244,In_181,In_511);
xnor U245 (N_245,In_550,In_456);
nor U246 (N_246,In_528,In_651);
or U247 (N_247,In_546,In_633);
and U248 (N_248,In_174,In_478);
xor U249 (N_249,In_448,In_87);
nor U250 (N_250,In_597,In_515);
nor U251 (N_251,In_357,In_472);
xor U252 (N_252,In_378,In_177);
nand U253 (N_253,In_156,In_581);
xnor U254 (N_254,In_491,In_331);
and U255 (N_255,In_429,In_615);
or U256 (N_256,In_223,In_532);
nand U257 (N_257,In_466,In_216);
nand U258 (N_258,In_201,In_73);
and U259 (N_259,In_589,In_110);
and U260 (N_260,In_557,In_540);
or U261 (N_261,In_629,In_372);
and U262 (N_262,In_149,In_32);
nor U263 (N_263,In_522,In_678);
nor U264 (N_264,In_711,In_340);
nand U265 (N_265,In_16,In_64);
or U266 (N_266,In_213,In_252);
and U267 (N_267,In_285,In_588);
nand U268 (N_268,In_159,In_17);
and U269 (N_269,In_37,In_503);
and U270 (N_270,In_231,In_443);
nor U271 (N_271,In_319,In_310);
xor U272 (N_272,In_299,In_465);
or U273 (N_273,In_718,In_337);
and U274 (N_274,In_136,In_649);
or U275 (N_275,In_724,In_278);
xnor U276 (N_276,In_452,In_389);
nand U277 (N_277,In_586,In_693);
nor U278 (N_278,In_625,In_254);
xnor U279 (N_279,In_569,In_24);
or U280 (N_280,In_498,In_492);
or U281 (N_281,In_526,In_279);
and U282 (N_282,In_67,In_165);
or U283 (N_283,In_225,In_219);
and U284 (N_284,In_206,In_667);
nor U285 (N_285,In_45,In_422);
nor U286 (N_286,In_184,In_523);
or U287 (N_287,In_459,In_574);
nand U288 (N_288,In_424,In_721);
nand U289 (N_289,In_61,In_359);
nand U290 (N_290,In_637,In_520);
nand U291 (N_291,In_737,In_193);
nor U292 (N_292,In_730,In_481);
and U293 (N_293,In_541,In_243);
or U294 (N_294,In_257,In_566);
nor U295 (N_295,In_698,In_654);
nand U296 (N_296,In_626,In_489);
nand U297 (N_297,In_163,In_354);
and U298 (N_298,In_627,In_199);
and U299 (N_299,In_140,In_386);
or U300 (N_300,In_238,In_648);
nor U301 (N_301,In_112,In_634);
nand U302 (N_302,In_273,In_380);
and U303 (N_303,In_247,In_512);
nor U304 (N_304,In_689,In_473);
or U305 (N_305,In_334,In_168);
xor U306 (N_306,In_226,In_166);
nor U307 (N_307,In_695,In_106);
or U308 (N_308,In_271,In_54);
or U309 (N_309,In_102,In_436);
nor U310 (N_310,In_36,In_570);
and U311 (N_311,In_620,In_703);
xnor U312 (N_312,In_284,In_198);
or U313 (N_313,In_80,In_176);
nor U314 (N_314,In_104,In_677);
or U315 (N_315,In_320,In_235);
nand U316 (N_316,In_306,In_296);
or U317 (N_317,In_508,In_712);
or U318 (N_318,In_641,In_179);
or U319 (N_319,In_74,In_316);
and U320 (N_320,In_612,In_56);
and U321 (N_321,In_19,In_450);
nor U322 (N_322,In_230,In_138);
and U323 (N_323,In_253,In_658);
and U324 (N_324,In_661,In_242);
nand U325 (N_325,In_96,In_190);
nor U326 (N_326,In_301,In_453);
and U327 (N_327,In_592,In_685);
nand U328 (N_328,In_474,In_601);
nor U329 (N_329,In_261,In_272);
nor U330 (N_330,In_28,In_364);
nand U331 (N_331,In_300,In_142);
nor U332 (N_332,In_27,In_471);
or U333 (N_333,In_160,In_101);
xor U334 (N_334,In_401,In_642);
xor U335 (N_335,In_215,In_376);
or U336 (N_336,In_749,In_313);
nor U337 (N_337,In_409,In_717);
nand U338 (N_338,In_441,In_270);
and U339 (N_339,In_178,In_682);
nor U340 (N_340,In_382,In_155);
or U341 (N_341,In_315,In_623);
or U342 (N_342,In_266,In_172);
and U343 (N_343,In_505,In_325);
nor U344 (N_344,In_561,In_547);
nor U345 (N_345,In_744,In_710);
nor U346 (N_346,In_530,In_88);
or U347 (N_347,In_650,In_244);
nor U348 (N_348,In_444,In_344);
xnor U349 (N_349,In_70,In_4);
or U350 (N_350,In_469,In_506);
nand U351 (N_351,In_578,In_317);
nor U352 (N_352,In_502,In_431);
xnor U353 (N_353,In_700,In_186);
nor U354 (N_354,In_323,In_451);
nand U355 (N_355,In_388,In_719);
nor U356 (N_356,In_211,In_268);
xor U357 (N_357,In_671,In_30);
and U358 (N_358,In_377,In_232);
or U359 (N_359,In_207,In_644);
nor U360 (N_360,In_399,In_280);
nand U361 (N_361,In_175,In_514);
xor U362 (N_362,In_662,In_132);
xnor U363 (N_363,In_350,In_158);
xor U364 (N_364,In_9,In_59);
nand U365 (N_365,In_619,In_205);
xnor U366 (N_366,In_180,In_675);
nor U367 (N_367,In_150,In_53);
or U368 (N_368,In_688,In_115);
nand U369 (N_369,In_153,In_412);
and U370 (N_370,In_122,In_352);
nand U371 (N_371,In_265,In_66);
or U372 (N_372,In_256,In_84);
nor U373 (N_373,In_704,In_663);
and U374 (N_374,In_144,In_157);
nor U375 (N_375,In_99,In_529);
nor U376 (N_376,In_139,In_102);
nor U377 (N_377,In_622,In_244);
nand U378 (N_378,In_228,In_309);
or U379 (N_379,In_323,In_206);
or U380 (N_380,In_10,In_29);
or U381 (N_381,In_500,In_579);
xnor U382 (N_382,In_670,In_356);
nand U383 (N_383,In_2,In_128);
nor U384 (N_384,In_172,In_337);
or U385 (N_385,In_230,In_424);
nand U386 (N_386,In_77,In_252);
and U387 (N_387,In_598,In_480);
nand U388 (N_388,In_7,In_548);
nand U389 (N_389,In_256,In_107);
or U390 (N_390,In_622,In_711);
nand U391 (N_391,In_728,In_404);
nand U392 (N_392,In_271,In_85);
and U393 (N_393,In_707,In_502);
and U394 (N_394,In_512,In_203);
nor U395 (N_395,In_364,In_217);
nand U396 (N_396,In_254,In_578);
and U397 (N_397,In_561,In_258);
nand U398 (N_398,In_530,In_211);
and U399 (N_399,In_220,In_479);
nor U400 (N_400,In_347,In_731);
or U401 (N_401,In_68,In_116);
nand U402 (N_402,In_455,In_681);
or U403 (N_403,In_453,In_131);
nand U404 (N_404,In_223,In_309);
and U405 (N_405,In_488,In_100);
or U406 (N_406,In_56,In_432);
nor U407 (N_407,In_317,In_141);
and U408 (N_408,In_282,In_683);
and U409 (N_409,In_155,In_472);
nor U410 (N_410,In_64,In_467);
and U411 (N_411,In_222,In_513);
nand U412 (N_412,In_390,In_65);
nor U413 (N_413,In_305,In_713);
and U414 (N_414,In_176,In_402);
nand U415 (N_415,In_353,In_397);
nand U416 (N_416,In_148,In_358);
nand U417 (N_417,In_471,In_657);
or U418 (N_418,In_163,In_532);
nor U419 (N_419,In_537,In_259);
nand U420 (N_420,In_356,In_559);
and U421 (N_421,In_117,In_689);
nor U422 (N_422,In_595,In_279);
and U423 (N_423,In_276,In_510);
or U424 (N_424,In_290,In_331);
nand U425 (N_425,In_563,In_235);
nor U426 (N_426,In_394,In_292);
xor U427 (N_427,In_548,In_502);
and U428 (N_428,In_667,In_634);
and U429 (N_429,In_541,In_156);
nand U430 (N_430,In_553,In_329);
xor U431 (N_431,In_555,In_211);
nand U432 (N_432,In_168,In_478);
nand U433 (N_433,In_85,In_203);
nand U434 (N_434,In_279,In_6);
and U435 (N_435,In_272,In_195);
nand U436 (N_436,In_24,In_212);
nand U437 (N_437,In_203,In_12);
nand U438 (N_438,In_365,In_533);
nand U439 (N_439,In_437,In_647);
or U440 (N_440,In_122,In_362);
nor U441 (N_441,In_130,In_736);
nand U442 (N_442,In_419,In_87);
nand U443 (N_443,In_645,In_619);
xnor U444 (N_444,In_329,In_301);
xnor U445 (N_445,In_497,In_356);
or U446 (N_446,In_10,In_126);
nor U447 (N_447,In_428,In_404);
or U448 (N_448,In_310,In_444);
nor U449 (N_449,In_67,In_570);
and U450 (N_450,In_123,In_242);
nand U451 (N_451,In_86,In_318);
or U452 (N_452,In_495,In_636);
nand U453 (N_453,In_404,In_450);
nand U454 (N_454,In_538,In_673);
and U455 (N_455,In_538,In_340);
nor U456 (N_456,In_613,In_657);
or U457 (N_457,In_651,In_606);
nor U458 (N_458,In_64,In_280);
nand U459 (N_459,In_626,In_576);
xnor U460 (N_460,In_138,In_533);
nand U461 (N_461,In_60,In_100);
nor U462 (N_462,In_564,In_400);
and U463 (N_463,In_559,In_717);
nand U464 (N_464,In_386,In_86);
or U465 (N_465,In_348,In_645);
nand U466 (N_466,In_547,In_475);
nor U467 (N_467,In_684,In_309);
nor U468 (N_468,In_359,In_423);
nand U469 (N_469,In_533,In_372);
and U470 (N_470,In_456,In_38);
and U471 (N_471,In_160,In_23);
nand U472 (N_472,In_445,In_638);
or U473 (N_473,In_600,In_195);
nand U474 (N_474,In_524,In_292);
nand U475 (N_475,In_676,In_606);
nand U476 (N_476,In_304,In_29);
nor U477 (N_477,In_703,In_262);
or U478 (N_478,In_142,In_205);
or U479 (N_479,In_218,In_598);
nor U480 (N_480,In_297,In_80);
nand U481 (N_481,In_731,In_568);
nor U482 (N_482,In_280,In_329);
nor U483 (N_483,In_598,In_140);
and U484 (N_484,In_384,In_516);
nand U485 (N_485,In_600,In_303);
and U486 (N_486,In_728,In_242);
nor U487 (N_487,In_655,In_15);
and U488 (N_488,In_673,In_708);
nand U489 (N_489,In_693,In_701);
nand U490 (N_490,In_167,In_80);
nand U491 (N_491,In_10,In_101);
and U492 (N_492,In_209,In_97);
nor U493 (N_493,In_373,In_20);
and U494 (N_494,In_227,In_625);
and U495 (N_495,In_416,In_728);
nor U496 (N_496,In_589,In_46);
xor U497 (N_497,In_696,In_545);
and U498 (N_498,In_164,In_156);
and U499 (N_499,In_396,In_745);
nand U500 (N_500,In_221,In_228);
or U501 (N_501,In_31,In_341);
or U502 (N_502,In_404,In_245);
or U503 (N_503,In_479,In_52);
and U504 (N_504,In_295,In_567);
nor U505 (N_505,In_739,In_602);
nand U506 (N_506,In_370,In_87);
nand U507 (N_507,In_473,In_629);
or U508 (N_508,In_386,In_493);
nand U509 (N_509,In_82,In_483);
or U510 (N_510,In_721,In_194);
nand U511 (N_511,In_661,In_360);
nand U512 (N_512,In_143,In_596);
and U513 (N_513,In_361,In_428);
nand U514 (N_514,In_306,In_653);
or U515 (N_515,In_494,In_141);
and U516 (N_516,In_381,In_94);
or U517 (N_517,In_91,In_395);
or U518 (N_518,In_538,In_242);
and U519 (N_519,In_436,In_612);
nand U520 (N_520,In_542,In_38);
and U521 (N_521,In_441,In_554);
or U522 (N_522,In_295,In_373);
xnor U523 (N_523,In_351,In_37);
and U524 (N_524,In_610,In_363);
nor U525 (N_525,In_315,In_536);
and U526 (N_526,In_3,In_186);
and U527 (N_527,In_462,In_149);
and U528 (N_528,In_563,In_600);
xor U529 (N_529,In_737,In_96);
or U530 (N_530,In_390,In_264);
or U531 (N_531,In_412,In_296);
and U532 (N_532,In_324,In_294);
nand U533 (N_533,In_657,In_233);
xor U534 (N_534,In_672,In_348);
or U535 (N_535,In_230,In_538);
xnor U536 (N_536,In_409,In_577);
and U537 (N_537,In_682,In_365);
and U538 (N_538,In_586,In_142);
and U539 (N_539,In_167,In_745);
or U540 (N_540,In_651,In_81);
nor U541 (N_541,In_712,In_484);
or U542 (N_542,In_484,In_627);
nand U543 (N_543,In_69,In_98);
nand U544 (N_544,In_568,In_45);
and U545 (N_545,In_508,In_66);
and U546 (N_546,In_297,In_629);
and U547 (N_547,In_321,In_498);
nand U548 (N_548,In_390,In_491);
nor U549 (N_549,In_522,In_52);
nand U550 (N_550,In_378,In_24);
or U551 (N_551,In_650,In_415);
nor U552 (N_552,In_307,In_370);
and U553 (N_553,In_19,In_66);
nand U554 (N_554,In_153,In_53);
or U555 (N_555,In_644,In_465);
or U556 (N_556,In_23,In_269);
nand U557 (N_557,In_232,In_230);
nor U558 (N_558,In_555,In_646);
nand U559 (N_559,In_240,In_56);
nor U560 (N_560,In_129,In_183);
nand U561 (N_561,In_624,In_251);
nor U562 (N_562,In_278,In_127);
or U563 (N_563,In_207,In_360);
and U564 (N_564,In_190,In_340);
and U565 (N_565,In_257,In_49);
nor U566 (N_566,In_610,In_113);
nor U567 (N_567,In_618,In_429);
nor U568 (N_568,In_635,In_16);
and U569 (N_569,In_666,In_242);
xnor U570 (N_570,In_404,In_104);
nand U571 (N_571,In_390,In_629);
or U572 (N_572,In_43,In_630);
xor U573 (N_573,In_571,In_457);
nor U574 (N_574,In_534,In_92);
nand U575 (N_575,In_614,In_578);
nor U576 (N_576,In_526,In_287);
nand U577 (N_577,In_302,In_483);
and U578 (N_578,In_297,In_72);
nor U579 (N_579,In_274,In_331);
nor U580 (N_580,In_337,In_169);
xor U581 (N_581,In_515,In_314);
and U582 (N_582,In_363,In_577);
or U583 (N_583,In_310,In_505);
nand U584 (N_584,In_268,In_296);
nor U585 (N_585,In_89,In_146);
nand U586 (N_586,In_726,In_748);
or U587 (N_587,In_204,In_137);
or U588 (N_588,In_117,In_286);
nand U589 (N_589,In_47,In_716);
or U590 (N_590,In_407,In_106);
and U591 (N_591,In_522,In_628);
or U592 (N_592,In_231,In_437);
nor U593 (N_593,In_730,In_667);
xnor U594 (N_594,In_132,In_105);
and U595 (N_595,In_320,In_286);
and U596 (N_596,In_275,In_625);
xor U597 (N_597,In_134,In_651);
xor U598 (N_598,In_548,In_327);
nor U599 (N_599,In_396,In_554);
or U600 (N_600,In_373,In_348);
nor U601 (N_601,In_169,In_506);
nor U602 (N_602,In_22,In_669);
and U603 (N_603,In_359,In_497);
and U604 (N_604,In_313,In_296);
and U605 (N_605,In_548,In_540);
nand U606 (N_606,In_507,In_680);
or U607 (N_607,In_529,In_649);
nand U608 (N_608,In_560,In_87);
nor U609 (N_609,In_435,In_699);
and U610 (N_610,In_0,In_426);
or U611 (N_611,In_637,In_621);
or U612 (N_612,In_702,In_200);
nor U613 (N_613,In_707,In_527);
or U614 (N_614,In_232,In_87);
nand U615 (N_615,In_489,In_376);
xor U616 (N_616,In_645,In_389);
and U617 (N_617,In_468,In_16);
nor U618 (N_618,In_117,In_639);
xnor U619 (N_619,In_624,In_444);
and U620 (N_620,In_84,In_626);
nand U621 (N_621,In_711,In_743);
or U622 (N_622,In_63,In_699);
nor U623 (N_623,In_437,In_353);
or U624 (N_624,In_528,In_398);
or U625 (N_625,In_216,In_666);
nor U626 (N_626,In_138,In_423);
nor U627 (N_627,In_475,In_616);
and U628 (N_628,In_16,In_702);
xor U629 (N_629,In_266,In_487);
nor U630 (N_630,In_526,In_148);
xor U631 (N_631,In_383,In_388);
nor U632 (N_632,In_99,In_595);
nor U633 (N_633,In_375,In_339);
or U634 (N_634,In_614,In_476);
and U635 (N_635,In_290,In_7);
and U636 (N_636,In_438,In_689);
and U637 (N_637,In_744,In_607);
nor U638 (N_638,In_599,In_234);
nand U639 (N_639,In_526,In_199);
or U640 (N_640,In_147,In_279);
nor U641 (N_641,In_257,In_420);
or U642 (N_642,In_244,In_420);
nand U643 (N_643,In_364,In_581);
xor U644 (N_644,In_697,In_295);
nor U645 (N_645,In_647,In_673);
nor U646 (N_646,In_570,In_201);
or U647 (N_647,In_506,In_188);
and U648 (N_648,In_201,In_493);
nand U649 (N_649,In_201,In_342);
nand U650 (N_650,In_351,In_260);
nand U651 (N_651,In_178,In_475);
and U652 (N_652,In_414,In_15);
nor U653 (N_653,In_230,In_612);
or U654 (N_654,In_358,In_666);
nor U655 (N_655,In_295,In_606);
or U656 (N_656,In_716,In_311);
and U657 (N_657,In_490,In_588);
and U658 (N_658,In_624,In_332);
nand U659 (N_659,In_268,In_269);
nand U660 (N_660,In_620,In_126);
or U661 (N_661,In_644,In_604);
nor U662 (N_662,In_635,In_83);
nor U663 (N_663,In_232,In_556);
nand U664 (N_664,In_384,In_549);
nand U665 (N_665,In_73,In_80);
nor U666 (N_666,In_669,In_48);
or U667 (N_667,In_31,In_546);
nand U668 (N_668,In_221,In_446);
or U669 (N_669,In_591,In_119);
xor U670 (N_670,In_667,In_435);
or U671 (N_671,In_625,In_510);
and U672 (N_672,In_215,In_621);
nor U673 (N_673,In_270,In_484);
or U674 (N_674,In_375,In_735);
and U675 (N_675,In_474,In_217);
or U676 (N_676,In_519,In_46);
nor U677 (N_677,In_172,In_475);
nor U678 (N_678,In_607,In_649);
and U679 (N_679,In_154,In_599);
or U680 (N_680,In_733,In_678);
and U681 (N_681,In_741,In_450);
nor U682 (N_682,In_119,In_584);
nor U683 (N_683,In_127,In_528);
nand U684 (N_684,In_519,In_723);
and U685 (N_685,In_74,In_254);
nand U686 (N_686,In_430,In_431);
or U687 (N_687,In_59,In_12);
and U688 (N_688,In_310,In_238);
nand U689 (N_689,In_295,In_618);
nand U690 (N_690,In_491,In_2);
nand U691 (N_691,In_541,In_55);
nor U692 (N_692,In_601,In_48);
or U693 (N_693,In_41,In_137);
nand U694 (N_694,In_558,In_46);
nand U695 (N_695,In_719,In_430);
nand U696 (N_696,In_509,In_635);
and U697 (N_697,In_97,In_505);
and U698 (N_698,In_301,In_391);
nand U699 (N_699,In_75,In_39);
nand U700 (N_700,In_303,In_519);
and U701 (N_701,In_79,In_670);
nor U702 (N_702,In_444,In_734);
and U703 (N_703,In_730,In_405);
nor U704 (N_704,In_554,In_286);
and U705 (N_705,In_702,In_470);
nor U706 (N_706,In_141,In_501);
nor U707 (N_707,In_539,In_598);
or U708 (N_708,In_568,In_1);
nor U709 (N_709,In_164,In_703);
or U710 (N_710,In_684,In_40);
nor U711 (N_711,In_49,In_8);
nor U712 (N_712,In_352,In_637);
xor U713 (N_713,In_711,In_289);
and U714 (N_714,In_749,In_713);
nand U715 (N_715,In_279,In_227);
and U716 (N_716,In_244,In_186);
or U717 (N_717,In_636,In_282);
and U718 (N_718,In_178,In_553);
or U719 (N_719,In_648,In_348);
or U720 (N_720,In_400,In_470);
and U721 (N_721,In_516,In_296);
nor U722 (N_722,In_737,In_133);
nand U723 (N_723,In_198,In_105);
nand U724 (N_724,In_207,In_579);
nand U725 (N_725,In_493,In_437);
nor U726 (N_726,In_501,In_474);
and U727 (N_727,In_187,In_452);
and U728 (N_728,In_249,In_700);
nand U729 (N_729,In_494,In_591);
and U730 (N_730,In_584,In_357);
and U731 (N_731,In_37,In_431);
and U732 (N_732,In_579,In_402);
nand U733 (N_733,In_128,In_717);
nand U734 (N_734,In_99,In_670);
xor U735 (N_735,In_112,In_64);
nor U736 (N_736,In_91,In_601);
nor U737 (N_737,In_713,In_299);
or U738 (N_738,In_421,In_649);
and U739 (N_739,In_703,In_647);
or U740 (N_740,In_62,In_377);
nor U741 (N_741,In_674,In_646);
xor U742 (N_742,In_652,In_61);
and U743 (N_743,In_717,In_711);
or U744 (N_744,In_65,In_355);
nand U745 (N_745,In_319,In_438);
nand U746 (N_746,In_372,In_213);
or U747 (N_747,In_36,In_462);
and U748 (N_748,In_456,In_304);
or U749 (N_749,In_234,In_738);
or U750 (N_750,In_29,In_393);
xnor U751 (N_751,In_659,In_0);
and U752 (N_752,In_527,In_256);
or U753 (N_753,In_544,In_557);
nor U754 (N_754,In_612,In_704);
nand U755 (N_755,In_705,In_591);
xor U756 (N_756,In_208,In_241);
and U757 (N_757,In_508,In_596);
or U758 (N_758,In_621,In_359);
and U759 (N_759,In_696,In_337);
or U760 (N_760,In_368,In_628);
or U761 (N_761,In_199,In_163);
xnor U762 (N_762,In_313,In_456);
and U763 (N_763,In_749,In_21);
nand U764 (N_764,In_247,In_430);
or U765 (N_765,In_665,In_157);
or U766 (N_766,In_111,In_41);
nor U767 (N_767,In_665,In_545);
or U768 (N_768,In_733,In_288);
xnor U769 (N_769,In_15,In_419);
xnor U770 (N_770,In_26,In_432);
xor U771 (N_771,In_633,In_306);
or U772 (N_772,In_739,In_214);
xor U773 (N_773,In_692,In_31);
nor U774 (N_774,In_668,In_283);
or U775 (N_775,In_554,In_584);
or U776 (N_776,In_222,In_147);
xnor U777 (N_777,In_472,In_429);
and U778 (N_778,In_545,In_82);
nand U779 (N_779,In_366,In_449);
nor U780 (N_780,In_654,In_671);
nor U781 (N_781,In_48,In_104);
and U782 (N_782,In_313,In_596);
or U783 (N_783,In_144,In_529);
xnor U784 (N_784,In_503,In_471);
nor U785 (N_785,In_258,In_207);
or U786 (N_786,In_275,In_608);
and U787 (N_787,In_407,In_703);
nor U788 (N_788,In_200,In_239);
nor U789 (N_789,In_113,In_597);
nor U790 (N_790,In_335,In_365);
nand U791 (N_791,In_347,In_436);
nor U792 (N_792,In_602,In_654);
or U793 (N_793,In_256,In_157);
nor U794 (N_794,In_375,In_288);
nand U795 (N_795,In_179,In_419);
nand U796 (N_796,In_711,In_529);
nand U797 (N_797,In_362,In_569);
nand U798 (N_798,In_22,In_465);
or U799 (N_799,In_303,In_645);
or U800 (N_800,In_256,In_549);
xnor U801 (N_801,In_531,In_523);
or U802 (N_802,In_3,In_357);
xor U803 (N_803,In_375,In_380);
xnor U804 (N_804,In_341,In_732);
and U805 (N_805,In_34,In_633);
or U806 (N_806,In_323,In_468);
or U807 (N_807,In_539,In_248);
nand U808 (N_808,In_630,In_486);
or U809 (N_809,In_110,In_666);
and U810 (N_810,In_470,In_102);
nand U811 (N_811,In_681,In_476);
nor U812 (N_812,In_56,In_461);
and U813 (N_813,In_189,In_303);
or U814 (N_814,In_189,In_172);
or U815 (N_815,In_268,In_142);
nand U816 (N_816,In_622,In_421);
nor U817 (N_817,In_347,In_272);
and U818 (N_818,In_466,In_204);
nand U819 (N_819,In_447,In_266);
nand U820 (N_820,In_142,In_474);
nor U821 (N_821,In_660,In_509);
nand U822 (N_822,In_355,In_562);
nor U823 (N_823,In_100,In_531);
and U824 (N_824,In_632,In_680);
and U825 (N_825,In_435,In_438);
or U826 (N_826,In_472,In_299);
nor U827 (N_827,In_532,In_58);
or U828 (N_828,In_7,In_452);
nor U829 (N_829,In_344,In_713);
nand U830 (N_830,In_295,In_415);
nor U831 (N_831,In_592,In_167);
xor U832 (N_832,In_281,In_58);
or U833 (N_833,In_497,In_294);
and U834 (N_834,In_20,In_102);
or U835 (N_835,In_633,In_733);
and U836 (N_836,In_545,In_258);
nor U837 (N_837,In_198,In_397);
and U838 (N_838,In_175,In_323);
nand U839 (N_839,In_279,In_488);
nand U840 (N_840,In_510,In_545);
nand U841 (N_841,In_284,In_87);
and U842 (N_842,In_705,In_55);
and U843 (N_843,In_493,In_707);
or U844 (N_844,In_343,In_397);
or U845 (N_845,In_233,In_728);
and U846 (N_846,In_147,In_208);
nor U847 (N_847,In_28,In_185);
nor U848 (N_848,In_29,In_419);
or U849 (N_849,In_659,In_134);
and U850 (N_850,In_138,In_266);
nor U851 (N_851,In_108,In_333);
nor U852 (N_852,In_338,In_108);
nor U853 (N_853,In_396,In_483);
nand U854 (N_854,In_120,In_729);
nor U855 (N_855,In_25,In_526);
or U856 (N_856,In_319,In_427);
or U857 (N_857,In_7,In_110);
xnor U858 (N_858,In_48,In_68);
and U859 (N_859,In_52,In_95);
nand U860 (N_860,In_63,In_614);
and U861 (N_861,In_575,In_742);
nand U862 (N_862,In_459,In_348);
xor U863 (N_863,In_225,In_530);
nor U864 (N_864,In_609,In_628);
or U865 (N_865,In_163,In_601);
nor U866 (N_866,In_577,In_37);
or U867 (N_867,In_689,In_158);
or U868 (N_868,In_108,In_323);
or U869 (N_869,In_459,In_104);
nand U870 (N_870,In_25,In_680);
or U871 (N_871,In_748,In_462);
and U872 (N_872,In_184,In_623);
nor U873 (N_873,In_529,In_512);
nor U874 (N_874,In_68,In_633);
and U875 (N_875,In_12,In_211);
and U876 (N_876,In_330,In_54);
or U877 (N_877,In_315,In_537);
and U878 (N_878,In_129,In_474);
nor U879 (N_879,In_410,In_643);
nand U880 (N_880,In_670,In_135);
xor U881 (N_881,In_416,In_43);
nor U882 (N_882,In_312,In_481);
nand U883 (N_883,In_137,In_621);
and U884 (N_884,In_217,In_287);
or U885 (N_885,In_514,In_670);
or U886 (N_886,In_678,In_318);
nor U887 (N_887,In_263,In_277);
nor U888 (N_888,In_346,In_189);
nor U889 (N_889,In_129,In_108);
or U890 (N_890,In_578,In_50);
and U891 (N_891,In_357,In_18);
nor U892 (N_892,In_697,In_738);
and U893 (N_893,In_279,In_544);
nand U894 (N_894,In_322,In_614);
or U895 (N_895,In_581,In_543);
nand U896 (N_896,In_594,In_1);
xnor U897 (N_897,In_156,In_589);
nand U898 (N_898,In_397,In_379);
and U899 (N_899,In_438,In_132);
nand U900 (N_900,In_158,In_185);
and U901 (N_901,In_63,In_377);
and U902 (N_902,In_242,In_316);
xor U903 (N_903,In_618,In_495);
and U904 (N_904,In_507,In_285);
xor U905 (N_905,In_564,In_651);
xnor U906 (N_906,In_210,In_636);
and U907 (N_907,In_334,In_607);
nor U908 (N_908,In_495,In_739);
nor U909 (N_909,In_414,In_700);
nor U910 (N_910,In_365,In_338);
or U911 (N_911,In_563,In_173);
and U912 (N_912,In_477,In_175);
nor U913 (N_913,In_200,In_157);
and U914 (N_914,In_659,In_15);
and U915 (N_915,In_138,In_650);
nor U916 (N_916,In_465,In_396);
and U917 (N_917,In_66,In_15);
nand U918 (N_918,In_115,In_586);
and U919 (N_919,In_249,In_362);
or U920 (N_920,In_386,In_113);
nand U921 (N_921,In_441,In_140);
and U922 (N_922,In_643,In_361);
and U923 (N_923,In_47,In_439);
nand U924 (N_924,In_685,In_148);
or U925 (N_925,In_678,In_255);
xor U926 (N_926,In_433,In_409);
nor U927 (N_927,In_285,In_397);
or U928 (N_928,In_722,In_496);
nor U929 (N_929,In_724,In_49);
nand U930 (N_930,In_19,In_451);
nor U931 (N_931,In_605,In_492);
or U932 (N_932,In_250,In_53);
nor U933 (N_933,In_305,In_469);
and U934 (N_934,In_466,In_0);
and U935 (N_935,In_437,In_716);
or U936 (N_936,In_43,In_746);
and U937 (N_937,In_447,In_690);
nand U938 (N_938,In_551,In_695);
nand U939 (N_939,In_584,In_739);
and U940 (N_940,In_391,In_267);
or U941 (N_941,In_66,In_112);
nor U942 (N_942,In_481,In_377);
and U943 (N_943,In_669,In_297);
nor U944 (N_944,In_168,In_611);
nand U945 (N_945,In_542,In_511);
nor U946 (N_946,In_569,In_700);
and U947 (N_947,In_613,In_59);
nand U948 (N_948,In_717,In_48);
nor U949 (N_949,In_497,In_660);
nand U950 (N_950,In_661,In_518);
or U951 (N_951,In_284,In_749);
nor U952 (N_952,In_48,In_321);
or U953 (N_953,In_1,In_690);
or U954 (N_954,In_533,In_744);
and U955 (N_955,In_268,In_449);
nor U956 (N_956,In_604,In_450);
or U957 (N_957,In_695,In_584);
nor U958 (N_958,In_219,In_499);
and U959 (N_959,In_279,In_389);
nand U960 (N_960,In_40,In_212);
nor U961 (N_961,In_83,In_325);
nor U962 (N_962,In_0,In_435);
nand U963 (N_963,In_137,In_311);
or U964 (N_964,In_710,In_169);
nand U965 (N_965,In_94,In_507);
nor U966 (N_966,In_303,In_158);
xnor U967 (N_967,In_613,In_240);
nor U968 (N_968,In_40,In_209);
or U969 (N_969,In_45,In_697);
nor U970 (N_970,In_138,In_520);
and U971 (N_971,In_224,In_405);
or U972 (N_972,In_677,In_294);
or U973 (N_973,In_246,In_542);
nor U974 (N_974,In_325,In_741);
or U975 (N_975,In_57,In_164);
nor U976 (N_976,In_388,In_392);
nor U977 (N_977,In_730,In_652);
nand U978 (N_978,In_52,In_609);
xnor U979 (N_979,In_427,In_502);
nor U980 (N_980,In_109,In_176);
nor U981 (N_981,In_139,In_36);
and U982 (N_982,In_113,In_131);
nand U983 (N_983,In_211,In_736);
xnor U984 (N_984,In_518,In_517);
nor U985 (N_985,In_245,In_365);
nor U986 (N_986,In_565,In_101);
and U987 (N_987,In_4,In_2);
nor U988 (N_988,In_86,In_27);
and U989 (N_989,In_647,In_539);
nand U990 (N_990,In_383,In_316);
and U991 (N_991,In_305,In_43);
xor U992 (N_992,In_506,In_428);
xor U993 (N_993,In_262,In_33);
xor U994 (N_994,In_655,In_371);
and U995 (N_995,In_509,In_748);
or U996 (N_996,In_95,In_460);
or U997 (N_997,In_735,In_250);
and U998 (N_998,In_435,In_352);
nand U999 (N_999,In_377,In_565);
and U1000 (N_1000,In_735,In_38);
nor U1001 (N_1001,In_137,In_18);
and U1002 (N_1002,In_37,In_185);
and U1003 (N_1003,In_201,In_748);
nand U1004 (N_1004,In_30,In_589);
or U1005 (N_1005,In_420,In_134);
or U1006 (N_1006,In_426,In_721);
nor U1007 (N_1007,In_409,In_66);
or U1008 (N_1008,In_326,In_247);
or U1009 (N_1009,In_428,In_370);
or U1010 (N_1010,In_1,In_593);
nor U1011 (N_1011,In_139,In_438);
or U1012 (N_1012,In_509,In_109);
nor U1013 (N_1013,In_587,In_58);
nor U1014 (N_1014,In_616,In_440);
nand U1015 (N_1015,In_376,In_410);
nor U1016 (N_1016,In_307,In_679);
or U1017 (N_1017,In_340,In_368);
or U1018 (N_1018,In_72,In_224);
nor U1019 (N_1019,In_690,In_718);
and U1020 (N_1020,In_76,In_490);
or U1021 (N_1021,In_638,In_150);
xnor U1022 (N_1022,In_69,In_225);
xnor U1023 (N_1023,In_188,In_569);
nor U1024 (N_1024,In_654,In_526);
xor U1025 (N_1025,In_205,In_255);
and U1026 (N_1026,In_711,In_167);
nand U1027 (N_1027,In_121,In_510);
nand U1028 (N_1028,In_235,In_204);
or U1029 (N_1029,In_599,In_284);
nor U1030 (N_1030,In_448,In_296);
nor U1031 (N_1031,In_569,In_562);
and U1032 (N_1032,In_731,In_101);
nand U1033 (N_1033,In_453,In_729);
nor U1034 (N_1034,In_568,In_444);
and U1035 (N_1035,In_151,In_135);
and U1036 (N_1036,In_131,In_164);
nor U1037 (N_1037,In_299,In_336);
and U1038 (N_1038,In_628,In_741);
and U1039 (N_1039,In_745,In_516);
or U1040 (N_1040,In_688,In_12);
and U1041 (N_1041,In_253,In_558);
or U1042 (N_1042,In_358,In_701);
and U1043 (N_1043,In_54,In_425);
or U1044 (N_1044,In_684,In_458);
or U1045 (N_1045,In_662,In_479);
xnor U1046 (N_1046,In_19,In_447);
nand U1047 (N_1047,In_631,In_344);
and U1048 (N_1048,In_137,In_632);
xor U1049 (N_1049,In_632,In_453);
nand U1050 (N_1050,In_219,In_257);
nand U1051 (N_1051,In_55,In_481);
or U1052 (N_1052,In_227,In_746);
or U1053 (N_1053,In_654,In_384);
or U1054 (N_1054,In_114,In_255);
and U1055 (N_1055,In_745,In_663);
nor U1056 (N_1056,In_106,In_287);
nand U1057 (N_1057,In_486,In_712);
or U1058 (N_1058,In_388,In_293);
nor U1059 (N_1059,In_152,In_441);
nor U1060 (N_1060,In_554,In_173);
or U1061 (N_1061,In_633,In_253);
and U1062 (N_1062,In_201,In_175);
and U1063 (N_1063,In_249,In_597);
nor U1064 (N_1064,In_480,In_412);
and U1065 (N_1065,In_144,In_399);
and U1066 (N_1066,In_428,In_31);
nor U1067 (N_1067,In_561,In_117);
or U1068 (N_1068,In_289,In_200);
and U1069 (N_1069,In_100,In_560);
nand U1070 (N_1070,In_337,In_291);
xnor U1071 (N_1071,In_358,In_132);
xnor U1072 (N_1072,In_511,In_44);
nor U1073 (N_1073,In_480,In_262);
or U1074 (N_1074,In_700,In_236);
or U1075 (N_1075,In_224,In_469);
nor U1076 (N_1076,In_478,In_184);
or U1077 (N_1077,In_391,In_304);
nor U1078 (N_1078,In_49,In_337);
or U1079 (N_1079,In_337,In_498);
nor U1080 (N_1080,In_59,In_393);
xnor U1081 (N_1081,In_512,In_333);
nor U1082 (N_1082,In_329,In_72);
xor U1083 (N_1083,In_123,In_333);
nor U1084 (N_1084,In_121,In_329);
nor U1085 (N_1085,In_611,In_335);
nand U1086 (N_1086,In_160,In_616);
nand U1087 (N_1087,In_439,In_414);
nor U1088 (N_1088,In_695,In_355);
nor U1089 (N_1089,In_317,In_535);
and U1090 (N_1090,In_76,In_113);
nor U1091 (N_1091,In_733,In_645);
nor U1092 (N_1092,In_141,In_53);
and U1093 (N_1093,In_132,In_718);
and U1094 (N_1094,In_98,In_361);
and U1095 (N_1095,In_659,In_502);
nand U1096 (N_1096,In_202,In_263);
and U1097 (N_1097,In_126,In_259);
and U1098 (N_1098,In_692,In_122);
xnor U1099 (N_1099,In_41,In_411);
nor U1100 (N_1100,In_122,In_540);
nor U1101 (N_1101,In_89,In_283);
and U1102 (N_1102,In_177,In_550);
nor U1103 (N_1103,In_60,In_42);
xnor U1104 (N_1104,In_317,In_729);
nand U1105 (N_1105,In_308,In_618);
nand U1106 (N_1106,In_158,In_280);
nand U1107 (N_1107,In_684,In_575);
or U1108 (N_1108,In_725,In_610);
and U1109 (N_1109,In_469,In_666);
xnor U1110 (N_1110,In_153,In_109);
and U1111 (N_1111,In_91,In_90);
nand U1112 (N_1112,In_434,In_228);
or U1113 (N_1113,In_84,In_118);
or U1114 (N_1114,In_403,In_227);
or U1115 (N_1115,In_267,In_304);
or U1116 (N_1116,In_14,In_491);
or U1117 (N_1117,In_748,In_68);
nor U1118 (N_1118,In_42,In_740);
or U1119 (N_1119,In_38,In_694);
xnor U1120 (N_1120,In_359,In_24);
nand U1121 (N_1121,In_682,In_337);
or U1122 (N_1122,In_736,In_622);
or U1123 (N_1123,In_560,In_695);
nand U1124 (N_1124,In_292,In_24);
and U1125 (N_1125,In_155,In_322);
nor U1126 (N_1126,In_18,In_265);
xor U1127 (N_1127,In_399,In_230);
nor U1128 (N_1128,In_621,In_49);
and U1129 (N_1129,In_728,In_48);
and U1130 (N_1130,In_397,In_363);
or U1131 (N_1131,In_189,In_667);
or U1132 (N_1132,In_225,In_203);
nand U1133 (N_1133,In_398,In_609);
or U1134 (N_1134,In_721,In_31);
nor U1135 (N_1135,In_299,In_108);
or U1136 (N_1136,In_334,In_591);
nor U1137 (N_1137,In_431,In_61);
or U1138 (N_1138,In_108,In_260);
nand U1139 (N_1139,In_403,In_575);
or U1140 (N_1140,In_384,In_287);
and U1141 (N_1141,In_417,In_625);
nor U1142 (N_1142,In_414,In_357);
nor U1143 (N_1143,In_630,In_239);
nor U1144 (N_1144,In_20,In_460);
xor U1145 (N_1145,In_256,In_361);
nand U1146 (N_1146,In_259,In_511);
and U1147 (N_1147,In_157,In_646);
xnor U1148 (N_1148,In_556,In_249);
nand U1149 (N_1149,In_457,In_86);
xnor U1150 (N_1150,In_599,In_466);
and U1151 (N_1151,In_131,In_259);
xnor U1152 (N_1152,In_94,In_484);
and U1153 (N_1153,In_479,In_403);
and U1154 (N_1154,In_279,In_415);
nand U1155 (N_1155,In_137,In_534);
nor U1156 (N_1156,In_417,In_272);
and U1157 (N_1157,In_489,In_242);
or U1158 (N_1158,In_646,In_24);
and U1159 (N_1159,In_321,In_719);
nor U1160 (N_1160,In_504,In_544);
or U1161 (N_1161,In_313,In_544);
xor U1162 (N_1162,In_444,In_185);
nand U1163 (N_1163,In_224,In_178);
or U1164 (N_1164,In_448,In_187);
or U1165 (N_1165,In_293,In_513);
nand U1166 (N_1166,In_261,In_39);
nor U1167 (N_1167,In_669,In_737);
and U1168 (N_1168,In_132,In_198);
or U1169 (N_1169,In_503,In_338);
nand U1170 (N_1170,In_61,In_63);
and U1171 (N_1171,In_6,In_27);
nor U1172 (N_1172,In_270,In_747);
nand U1173 (N_1173,In_120,In_402);
nand U1174 (N_1174,In_83,In_227);
and U1175 (N_1175,In_694,In_402);
nand U1176 (N_1176,In_622,In_574);
or U1177 (N_1177,In_356,In_515);
nand U1178 (N_1178,In_302,In_682);
nand U1179 (N_1179,In_687,In_586);
nand U1180 (N_1180,In_245,In_96);
nand U1181 (N_1181,In_547,In_558);
nor U1182 (N_1182,In_728,In_461);
or U1183 (N_1183,In_88,In_697);
and U1184 (N_1184,In_40,In_360);
or U1185 (N_1185,In_86,In_738);
nor U1186 (N_1186,In_155,In_340);
and U1187 (N_1187,In_123,In_546);
nand U1188 (N_1188,In_495,In_253);
xnor U1189 (N_1189,In_284,In_271);
nand U1190 (N_1190,In_716,In_327);
or U1191 (N_1191,In_199,In_733);
nor U1192 (N_1192,In_611,In_664);
xor U1193 (N_1193,In_522,In_321);
and U1194 (N_1194,In_166,In_682);
xnor U1195 (N_1195,In_620,In_496);
and U1196 (N_1196,In_561,In_654);
nand U1197 (N_1197,In_280,In_572);
or U1198 (N_1198,In_603,In_439);
nor U1199 (N_1199,In_218,In_219);
nor U1200 (N_1200,In_632,In_445);
or U1201 (N_1201,In_266,In_570);
and U1202 (N_1202,In_215,In_395);
nand U1203 (N_1203,In_377,In_61);
or U1204 (N_1204,In_614,In_150);
nand U1205 (N_1205,In_105,In_713);
nor U1206 (N_1206,In_335,In_413);
nand U1207 (N_1207,In_142,In_451);
nor U1208 (N_1208,In_161,In_14);
or U1209 (N_1209,In_21,In_633);
and U1210 (N_1210,In_269,In_726);
nand U1211 (N_1211,In_329,In_538);
or U1212 (N_1212,In_368,In_539);
or U1213 (N_1213,In_362,In_262);
nand U1214 (N_1214,In_550,In_91);
and U1215 (N_1215,In_300,In_470);
and U1216 (N_1216,In_623,In_228);
nor U1217 (N_1217,In_259,In_159);
xor U1218 (N_1218,In_624,In_532);
nor U1219 (N_1219,In_691,In_174);
or U1220 (N_1220,In_315,In_567);
nand U1221 (N_1221,In_672,In_60);
and U1222 (N_1222,In_647,In_439);
nor U1223 (N_1223,In_374,In_541);
nor U1224 (N_1224,In_513,In_110);
or U1225 (N_1225,In_459,In_131);
nand U1226 (N_1226,In_701,In_418);
or U1227 (N_1227,In_375,In_178);
xor U1228 (N_1228,In_683,In_243);
nor U1229 (N_1229,In_62,In_743);
or U1230 (N_1230,In_112,In_726);
and U1231 (N_1231,In_509,In_280);
xnor U1232 (N_1232,In_701,In_455);
nand U1233 (N_1233,In_343,In_500);
and U1234 (N_1234,In_101,In_525);
or U1235 (N_1235,In_234,In_31);
nand U1236 (N_1236,In_368,In_639);
nor U1237 (N_1237,In_511,In_687);
nor U1238 (N_1238,In_737,In_642);
and U1239 (N_1239,In_144,In_689);
nand U1240 (N_1240,In_193,In_166);
nand U1241 (N_1241,In_54,In_216);
nand U1242 (N_1242,In_576,In_248);
or U1243 (N_1243,In_609,In_76);
or U1244 (N_1244,In_631,In_299);
nor U1245 (N_1245,In_444,In_29);
nor U1246 (N_1246,In_162,In_619);
or U1247 (N_1247,In_163,In_555);
nor U1248 (N_1248,In_482,In_100);
nor U1249 (N_1249,In_448,In_38);
and U1250 (N_1250,In_61,In_235);
nand U1251 (N_1251,In_222,In_172);
nor U1252 (N_1252,In_115,In_296);
nor U1253 (N_1253,In_513,In_739);
or U1254 (N_1254,In_265,In_263);
xor U1255 (N_1255,In_544,In_558);
xor U1256 (N_1256,In_713,In_453);
and U1257 (N_1257,In_510,In_269);
nand U1258 (N_1258,In_19,In_713);
xor U1259 (N_1259,In_547,In_285);
or U1260 (N_1260,In_281,In_113);
and U1261 (N_1261,In_307,In_447);
nor U1262 (N_1262,In_542,In_614);
and U1263 (N_1263,In_228,In_304);
xor U1264 (N_1264,In_266,In_50);
nor U1265 (N_1265,In_459,In_350);
and U1266 (N_1266,In_312,In_101);
or U1267 (N_1267,In_91,In_468);
or U1268 (N_1268,In_605,In_451);
nand U1269 (N_1269,In_339,In_259);
nor U1270 (N_1270,In_485,In_365);
and U1271 (N_1271,In_423,In_441);
or U1272 (N_1272,In_700,In_517);
nor U1273 (N_1273,In_668,In_42);
nand U1274 (N_1274,In_719,In_470);
nor U1275 (N_1275,In_639,In_148);
xor U1276 (N_1276,In_237,In_367);
nor U1277 (N_1277,In_310,In_59);
nor U1278 (N_1278,In_321,In_235);
nor U1279 (N_1279,In_209,In_364);
and U1280 (N_1280,In_387,In_288);
or U1281 (N_1281,In_300,In_149);
or U1282 (N_1282,In_0,In_45);
and U1283 (N_1283,In_16,In_487);
or U1284 (N_1284,In_229,In_503);
nor U1285 (N_1285,In_340,In_551);
or U1286 (N_1286,In_389,In_366);
nor U1287 (N_1287,In_113,In_107);
nand U1288 (N_1288,In_712,In_705);
nor U1289 (N_1289,In_659,In_573);
nand U1290 (N_1290,In_207,In_67);
and U1291 (N_1291,In_270,In_487);
or U1292 (N_1292,In_71,In_126);
and U1293 (N_1293,In_194,In_691);
or U1294 (N_1294,In_19,In_680);
nor U1295 (N_1295,In_167,In_133);
nor U1296 (N_1296,In_238,In_102);
and U1297 (N_1297,In_17,In_513);
and U1298 (N_1298,In_249,In_35);
and U1299 (N_1299,In_267,In_498);
or U1300 (N_1300,In_583,In_358);
nor U1301 (N_1301,In_658,In_386);
or U1302 (N_1302,In_129,In_281);
and U1303 (N_1303,In_159,In_539);
nand U1304 (N_1304,In_635,In_571);
nand U1305 (N_1305,In_286,In_35);
or U1306 (N_1306,In_657,In_193);
nor U1307 (N_1307,In_129,In_316);
nor U1308 (N_1308,In_368,In_532);
xnor U1309 (N_1309,In_619,In_599);
or U1310 (N_1310,In_664,In_372);
xor U1311 (N_1311,In_57,In_449);
nand U1312 (N_1312,In_142,In_702);
nand U1313 (N_1313,In_695,In_356);
nand U1314 (N_1314,In_465,In_602);
and U1315 (N_1315,In_233,In_449);
and U1316 (N_1316,In_492,In_584);
xor U1317 (N_1317,In_429,In_681);
and U1318 (N_1318,In_282,In_721);
or U1319 (N_1319,In_680,In_62);
nand U1320 (N_1320,In_672,In_570);
nor U1321 (N_1321,In_619,In_92);
nor U1322 (N_1322,In_745,In_698);
nor U1323 (N_1323,In_55,In_373);
nor U1324 (N_1324,In_540,In_90);
xnor U1325 (N_1325,In_278,In_728);
and U1326 (N_1326,In_369,In_363);
and U1327 (N_1327,In_577,In_277);
xor U1328 (N_1328,In_187,In_297);
and U1329 (N_1329,In_452,In_469);
and U1330 (N_1330,In_169,In_484);
xnor U1331 (N_1331,In_566,In_431);
and U1332 (N_1332,In_76,In_502);
nand U1333 (N_1333,In_550,In_34);
nand U1334 (N_1334,In_239,In_75);
or U1335 (N_1335,In_524,In_371);
or U1336 (N_1336,In_447,In_710);
and U1337 (N_1337,In_517,In_655);
or U1338 (N_1338,In_648,In_37);
nand U1339 (N_1339,In_146,In_163);
or U1340 (N_1340,In_496,In_184);
nand U1341 (N_1341,In_73,In_556);
or U1342 (N_1342,In_494,In_89);
nand U1343 (N_1343,In_716,In_137);
xnor U1344 (N_1344,In_193,In_284);
nor U1345 (N_1345,In_316,In_516);
nor U1346 (N_1346,In_471,In_573);
and U1347 (N_1347,In_235,In_720);
nand U1348 (N_1348,In_325,In_202);
xor U1349 (N_1349,In_740,In_275);
nor U1350 (N_1350,In_616,In_158);
and U1351 (N_1351,In_393,In_719);
or U1352 (N_1352,In_71,In_412);
xnor U1353 (N_1353,In_137,In_301);
and U1354 (N_1354,In_526,In_436);
or U1355 (N_1355,In_461,In_418);
nand U1356 (N_1356,In_317,In_431);
nor U1357 (N_1357,In_597,In_550);
nor U1358 (N_1358,In_494,In_720);
nand U1359 (N_1359,In_601,In_279);
nand U1360 (N_1360,In_503,In_482);
xor U1361 (N_1361,In_368,In_713);
nor U1362 (N_1362,In_197,In_578);
nor U1363 (N_1363,In_153,In_503);
xor U1364 (N_1364,In_491,In_564);
nor U1365 (N_1365,In_81,In_475);
and U1366 (N_1366,In_439,In_163);
and U1367 (N_1367,In_86,In_32);
and U1368 (N_1368,In_162,In_323);
or U1369 (N_1369,In_258,In_268);
nand U1370 (N_1370,In_363,In_55);
nand U1371 (N_1371,In_712,In_572);
nand U1372 (N_1372,In_629,In_577);
and U1373 (N_1373,In_463,In_460);
xor U1374 (N_1374,In_555,In_115);
or U1375 (N_1375,In_313,In_132);
and U1376 (N_1376,In_740,In_114);
and U1377 (N_1377,In_427,In_231);
xor U1378 (N_1378,In_707,In_647);
nand U1379 (N_1379,In_415,In_486);
nand U1380 (N_1380,In_409,In_390);
and U1381 (N_1381,In_48,In_649);
or U1382 (N_1382,In_435,In_119);
xor U1383 (N_1383,In_631,In_731);
xnor U1384 (N_1384,In_696,In_48);
or U1385 (N_1385,In_54,In_26);
xnor U1386 (N_1386,In_595,In_214);
xor U1387 (N_1387,In_689,In_354);
nand U1388 (N_1388,In_440,In_302);
nand U1389 (N_1389,In_255,In_591);
or U1390 (N_1390,In_416,In_341);
xnor U1391 (N_1391,In_172,In_97);
nor U1392 (N_1392,In_582,In_224);
or U1393 (N_1393,In_648,In_507);
nand U1394 (N_1394,In_326,In_447);
nor U1395 (N_1395,In_624,In_468);
nand U1396 (N_1396,In_382,In_337);
and U1397 (N_1397,In_644,In_139);
nor U1398 (N_1398,In_463,In_403);
xnor U1399 (N_1399,In_330,In_105);
nor U1400 (N_1400,In_167,In_550);
or U1401 (N_1401,In_121,In_674);
xor U1402 (N_1402,In_228,In_371);
nand U1403 (N_1403,In_709,In_213);
and U1404 (N_1404,In_670,In_104);
xor U1405 (N_1405,In_6,In_413);
nor U1406 (N_1406,In_80,In_587);
nor U1407 (N_1407,In_496,In_335);
or U1408 (N_1408,In_277,In_561);
and U1409 (N_1409,In_28,In_233);
nor U1410 (N_1410,In_143,In_709);
or U1411 (N_1411,In_161,In_630);
nor U1412 (N_1412,In_749,In_532);
nand U1413 (N_1413,In_262,In_129);
nor U1414 (N_1414,In_322,In_237);
nor U1415 (N_1415,In_503,In_622);
and U1416 (N_1416,In_445,In_120);
and U1417 (N_1417,In_511,In_2);
or U1418 (N_1418,In_125,In_331);
xnor U1419 (N_1419,In_252,In_510);
nand U1420 (N_1420,In_536,In_463);
and U1421 (N_1421,In_673,In_510);
and U1422 (N_1422,In_458,In_432);
or U1423 (N_1423,In_475,In_421);
xor U1424 (N_1424,In_513,In_256);
and U1425 (N_1425,In_679,In_359);
or U1426 (N_1426,In_262,In_546);
and U1427 (N_1427,In_177,In_298);
nor U1428 (N_1428,In_182,In_79);
or U1429 (N_1429,In_274,In_202);
or U1430 (N_1430,In_96,In_174);
and U1431 (N_1431,In_647,In_104);
xnor U1432 (N_1432,In_213,In_420);
and U1433 (N_1433,In_648,In_472);
or U1434 (N_1434,In_160,In_415);
nor U1435 (N_1435,In_248,In_747);
nor U1436 (N_1436,In_127,In_423);
or U1437 (N_1437,In_20,In_589);
and U1438 (N_1438,In_115,In_302);
and U1439 (N_1439,In_304,In_328);
nand U1440 (N_1440,In_506,In_111);
nand U1441 (N_1441,In_189,In_220);
nor U1442 (N_1442,In_584,In_89);
and U1443 (N_1443,In_526,In_711);
and U1444 (N_1444,In_714,In_616);
nand U1445 (N_1445,In_517,In_96);
or U1446 (N_1446,In_92,In_418);
nand U1447 (N_1447,In_136,In_427);
and U1448 (N_1448,In_387,In_416);
nor U1449 (N_1449,In_516,In_409);
or U1450 (N_1450,In_124,In_450);
or U1451 (N_1451,In_397,In_689);
and U1452 (N_1452,In_68,In_64);
nor U1453 (N_1453,In_653,In_85);
or U1454 (N_1454,In_53,In_567);
and U1455 (N_1455,In_422,In_127);
or U1456 (N_1456,In_52,In_9);
and U1457 (N_1457,In_364,In_489);
nor U1458 (N_1458,In_723,In_701);
nand U1459 (N_1459,In_727,In_187);
and U1460 (N_1460,In_563,In_528);
nor U1461 (N_1461,In_522,In_424);
nor U1462 (N_1462,In_638,In_487);
nand U1463 (N_1463,In_363,In_480);
nor U1464 (N_1464,In_177,In_416);
or U1465 (N_1465,In_164,In_555);
or U1466 (N_1466,In_638,In_513);
or U1467 (N_1467,In_15,In_683);
nand U1468 (N_1468,In_441,In_341);
or U1469 (N_1469,In_717,In_520);
nand U1470 (N_1470,In_641,In_243);
nor U1471 (N_1471,In_190,In_9);
or U1472 (N_1472,In_169,In_286);
nand U1473 (N_1473,In_579,In_656);
xnor U1474 (N_1474,In_548,In_71);
nor U1475 (N_1475,In_425,In_368);
and U1476 (N_1476,In_688,In_525);
or U1477 (N_1477,In_229,In_400);
or U1478 (N_1478,In_328,In_127);
or U1479 (N_1479,In_193,In_39);
and U1480 (N_1480,In_166,In_311);
nand U1481 (N_1481,In_544,In_612);
or U1482 (N_1482,In_356,In_40);
or U1483 (N_1483,In_524,In_150);
nand U1484 (N_1484,In_287,In_295);
and U1485 (N_1485,In_667,In_357);
and U1486 (N_1486,In_673,In_289);
or U1487 (N_1487,In_496,In_556);
and U1488 (N_1488,In_321,In_618);
nand U1489 (N_1489,In_201,In_388);
nand U1490 (N_1490,In_393,In_529);
nand U1491 (N_1491,In_384,In_302);
nand U1492 (N_1492,In_55,In_692);
nand U1493 (N_1493,In_98,In_137);
nor U1494 (N_1494,In_248,In_358);
or U1495 (N_1495,In_333,In_156);
nor U1496 (N_1496,In_202,In_642);
xnor U1497 (N_1497,In_421,In_341);
and U1498 (N_1498,In_386,In_298);
nor U1499 (N_1499,In_274,In_528);
or U1500 (N_1500,In_233,In_276);
and U1501 (N_1501,In_692,In_88);
and U1502 (N_1502,In_707,In_528);
nand U1503 (N_1503,In_487,In_123);
xnor U1504 (N_1504,In_539,In_156);
and U1505 (N_1505,In_635,In_488);
nor U1506 (N_1506,In_157,In_84);
and U1507 (N_1507,In_567,In_562);
xnor U1508 (N_1508,In_335,In_483);
nor U1509 (N_1509,In_206,In_356);
nand U1510 (N_1510,In_130,In_608);
nor U1511 (N_1511,In_258,In_630);
nor U1512 (N_1512,In_108,In_258);
and U1513 (N_1513,In_431,In_353);
nor U1514 (N_1514,In_380,In_521);
nor U1515 (N_1515,In_139,In_748);
or U1516 (N_1516,In_517,In_302);
xor U1517 (N_1517,In_486,In_450);
nand U1518 (N_1518,In_575,In_653);
nand U1519 (N_1519,In_336,In_727);
nand U1520 (N_1520,In_276,In_585);
and U1521 (N_1521,In_128,In_749);
xor U1522 (N_1522,In_531,In_290);
or U1523 (N_1523,In_129,In_682);
nor U1524 (N_1524,In_514,In_277);
nand U1525 (N_1525,In_259,In_674);
or U1526 (N_1526,In_514,In_165);
nand U1527 (N_1527,In_246,In_607);
nor U1528 (N_1528,In_72,In_331);
and U1529 (N_1529,In_521,In_495);
and U1530 (N_1530,In_707,In_396);
nor U1531 (N_1531,In_522,In_581);
nor U1532 (N_1532,In_465,In_608);
nor U1533 (N_1533,In_475,In_556);
or U1534 (N_1534,In_579,In_110);
and U1535 (N_1535,In_653,In_138);
and U1536 (N_1536,In_36,In_349);
nor U1537 (N_1537,In_53,In_188);
and U1538 (N_1538,In_320,In_450);
or U1539 (N_1539,In_596,In_140);
nor U1540 (N_1540,In_660,In_37);
nor U1541 (N_1541,In_350,In_216);
or U1542 (N_1542,In_534,In_697);
nor U1543 (N_1543,In_718,In_407);
nand U1544 (N_1544,In_472,In_394);
and U1545 (N_1545,In_92,In_497);
or U1546 (N_1546,In_225,In_492);
or U1547 (N_1547,In_271,In_277);
and U1548 (N_1548,In_409,In_146);
nor U1549 (N_1549,In_525,In_16);
or U1550 (N_1550,In_574,In_342);
nor U1551 (N_1551,In_101,In_251);
nand U1552 (N_1552,In_264,In_47);
nor U1553 (N_1553,In_482,In_388);
nor U1554 (N_1554,In_7,In_454);
nand U1555 (N_1555,In_561,In_184);
and U1556 (N_1556,In_180,In_748);
and U1557 (N_1557,In_242,In_198);
and U1558 (N_1558,In_104,In_217);
and U1559 (N_1559,In_251,In_198);
nor U1560 (N_1560,In_135,In_366);
nor U1561 (N_1561,In_339,In_129);
nand U1562 (N_1562,In_595,In_300);
and U1563 (N_1563,In_359,In_394);
or U1564 (N_1564,In_59,In_606);
xor U1565 (N_1565,In_19,In_685);
and U1566 (N_1566,In_421,In_232);
and U1567 (N_1567,In_303,In_46);
nand U1568 (N_1568,In_76,In_105);
xnor U1569 (N_1569,In_203,In_342);
nand U1570 (N_1570,In_19,In_89);
nand U1571 (N_1571,In_573,In_338);
xnor U1572 (N_1572,In_216,In_186);
nor U1573 (N_1573,In_228,In_67);
or U1574 (N_1574,In_679,In_666);
and U1575 (N_1575,In_9,In_372);
nand U1576 (N_1576,In_91,In_386);
nor U1577 (N_1577,In_162,In_14);
xor U1578 (N_1578,In_710,In_398);
or U1579 (N_1579,In_401,In_374);
and U1580 (N_1580,In_527,In_726);
xnor U1581 (N_1581,In_446,In_93);
xnor U1582 (N_1582,In_555,In_434);
nor U1583 (N_1583,In_88,In_362);
nand U1584 (N_1584,In_132,In_523);
and U1585 (N_1585,In_342,In_239);
nor U1586 (N_1586,In_685,In_744);
and U1587 (N_1587,In_717,In_535);
and U1588 (N_1588,In_178,In_351);
and U1589 (N_1589,In_605,In_524);
and U1590 (N_1590,In_112,In_48);
and U1591 (N_1591,In_691,In_182);
or U1592 (N_1592,In_684,In_80);
xor U1593 (N_1593,In_371,In_714);
or U1594 (N_1594,In_736,In_722);
or U1595 (N_1595,In_455,In_686);
and U1596 (N_1596,In_10,In_719);
and U1597 (N_1597,In_221,In_224);
nand U1598 (N_1598,In_293,In_564);
nor U1599 (N_1599,In_496,In_364);
nand U1600 (N_1600,In_310,In_467);
and U1601 (N_1601,In_454,In_616);
nand U1602 (N_1602,In_168,In_329);
xnor U1603 (N_1603,In_237,In_59);
or U1604 (N_1604,In_196,In_702);
and U1605 (N_1605,In_468,In_514);
or U1606 (N_1606,In_690,In_356);
or U1607 (N_1607,In_60,In_630);
or U1608 (N_1608,In_218,In_40);
or U1609 (N_1609,In_293,In_19);
nand U1610 (N_1610,In_209,In_281);
nand U1611 (N_1611,In_448,In_489);
nor U1612 (N_1612,In_382,In_673);
nor U1613 (N_1613,In_438,In_306);
or U1614 (N_1614,In_687,In_627);
or U1615 (N_1615,In_603,In_397);
or U1616 (N_1616,In_289,In_285);
nor U1617 (N_1617,In_16,In_24);
nor U1618 (N_1618,In_740,In_44);
or U1619 (N_1619,In_626,In_627);
xor U1620 (N_1620,In_619,In_742);
or U1621 (N_1621,In_78,In_230);
nand U1622 (N_1622,In_110,In_379);
or U1623 (N_1623,In_658,In_512);
and U1624 (N_1624,In_432,In_218);
nor U1625 (N_1625,In_34,In_718);
xor U1626 (N_1626,In_624,In_629);
and U1627 (N_1627,In_139,In_40);
nand U1628 (N_1628,In_451,In_496);
or U1629 (N_1629,In_646,In_729);
or U1630 (N_1630,In_258,In_177);
or U1631 (N_1631,In_348,In_424);
xnor U1632 (N_1632,In_457,In_381);
nand U1633 (N_1633,In_546,In_365);
and U1634 (N_1634,In_686,In_15);
nand U1635 (N_1635,In_115,In_437);
nand U1636 (N_1636,In_452,In_165);
nand U1637 (N_1637,In_137,In_248);
nor U1638 (N_1638,In_237,In_193);
and U1639 (N_1639,In_4,In_160);
and U1640 (N_1640,In_252,In_28);
and U1641 (N_1641,In_741,In_568);
and U1642 (N_1642,In_529,In_146);
or U1643 (N_1643,In_304,In_171);
and U1644 (N_1644,In_485,In_92);
and U1645 (N_1645,In_369,In_136);
nor U1646 (N_1646,In_267,In_734);
nand U1647 (N_1647,In_529,In_675);
and U1648 (N_1648,In_688,In_15);
nand U1649 (N_1649,In_41,In_535);
nand U1650 (N_1650,In_622,In_485);
and U1651 (N_1651,In_117,In_714);
and U1652 (N_1652,In_316,In_735);
or U1653 (N_1653,In_298,In_463);
nand U1654 (N_1654,In_693,In_146);
nor U1655 (N_1655,In_6,In_149);
nand U1656 (N_1656,In_314,In_75);
or U1657 (N_1657,In_380,In_149);
nand U1658 (N_1658,In_293,In_263);
nor U1659 (N_1659,In_371,In_190);
nor U1660 (N_1660,In_235,In_358);
and U1661 (N_1661,In_163,In_67);
or U1662 (N_1662,In_531,In_519);
or U1663 (N_1663,In_366,In_583);
or U1664 (N_1664,In_20,In_689);
nor U1665 (N_1665,In_489,In_65);
nor U1666 (N_1666,In_436,In_687);
or U1667 (N_1667,In_93,In_186);
nand U1668 (N_1668,In_615,In_688);
nand U1669 (N_1669,In_150,In_15);
xor U1670 (N_1670,In_234,In_430);
nor U1671 (N_1671,In_598,In_695);
nor U1672 (N_1672,In_208,In_51);
or U1673 (N_1673,In_259,In_379);
and U1674 (N_1674,In_635,In_272);
or U1675 (N_1675,In_522,In_616);
and U1676 (N_1676,In_147,In_334);
or U1677 (N_1677,In_697,In_743);
nand U1678 (N_1678,In_247,In_695);
xor U1679 (N_1679,In_19,In_309);
nor U1680 (N_1680,In_483,In_595);
nand U1681 (N_1681,In_581,In_253);
nand U1682 (N_1682,In_371,In_428);
and U1683 (N_1683,In_600,In_377);
and U1684 (N_1684,In_460,In_128);
nand U1685 (N_1685,In_169,In_725);
and U1686 (N_1686,In_671,In_263);
xnor U1687 (N_1687,In_125,In_27);
or U1688 (N_1688,In_445,In_547);
or U1689 (N_1689,In_47,In_591);
and U1690 (N_1690,In_1,In_299);
nand U1691 (N_1691,In_541,In_210);
nand U1692 (N_1692,In_613,In_578);
nand U1693 (N_1693,In_339,In_158);
and U1694 (N_1694,In_399,In_129);
nor U1695 (N_1695,In_721,In_457);
or U1696 (N_1696,In_498,In_677);
or U1697 (N_1697,In_367,In_740);
nor U1698 (N_1698,In_595,In_673);
or U1699 (N_1699,In_535,In_189);
nor U1700 (N_1700,In_725,In_708);
nor U1701 (N_1701,In_313,In_536);
xnor U1702 (N_1702,In_75,In_717);
and U1703 (N_1703,In_49,In_279);
nand U1704 (N_1704,In_368,In_427);
nor U1705 (N_1705,In_551,In_595);
and U1706 (N_1706,In_659,In_565);
nand U1707 (N_1707,In_338,In_166);
or U1708 (N_1708,In_81,In_233);
and U1709 (N_1709,In_286,In_570);
and U1710 (N_1710,In_166,In_537);
nor U1711 (N_1711,In_69,In_204);
nand U1712 (N_1712,In_117,In_95);
or U1713 (N_1713,In_308,In_154);
xnor U1714 (N_1714,In_577,In_473);
and U1715 (N_1715,In_447,In_559);
or U1716 (N_1716,In_63,In_166);
nor U1717 (N_1717,In_253,In_566);
or U1718 (N_1718,In_223,In_235);
and U1719 (N_1719,In_361,In_233);
or U1720 (N_1720,In_46,In_362);
xor U1721 (N_1721,In_403,In_160);
or U1722 (N_1722,In_28,In_543);
nor U1723 (N_1723,In_146,In_515);
or U1724 (N_1724,In_147,In_411);
nand U1725 (N_1725,In_466,In_478);
and U1726 (N_1726,In_372,In_450);
nand U1727 (N_1727,In_280,In_401);
nor U1728 (N_1728,In_330,In_498);
or U1729 (N_1729,In_683,In_59);
nand U1730 (N_1730,In_192,In_556);
nand U1731 (N_1731,In_405,In_96);
xnor U1732 (N_1732,In_178,In_577);
nand U1733 (N_1733,In_37,In_534);
and U1734 (N_1734,In_377,In_651);
nand U1735 (N_1735,In_538,In_593);
nand U1736 (N_1736,In_344,In_235);
and U1737 (N_1737,In_258,In_740);
or U1738 (N_1738,In_118,In_607);
or U1739 (N_1739,In_394,In_350);
and U1740 (N_1740,In_657,In_663);
nand U1741 (N_1741,In_592,In_608);
or U1742 (N_1742,In_11,In_389);
nand U1743 (N_1743,In_437,In_620);
nand U1744 (N_1744,In_596,In_220);
nand U1745 (N_1745,In_424,In_100);
nor U1746 (N_1746,In_132,In_375);
and U1747 (N_1747,In_94,In_46);
nor U1748 (N_1748,In_162,In_46);
xnor U1749 (N_1749,In_525,In_429);
or U1750 (N_1750,In_258,In_97);
xor U1751 (N_1751,In_137,In_730);
and U1752 (N_1752,In_22,In_600);
nand U1753 (N_1753,In_501,In_534);
and U1754 (N_1754,In_451,In_156);
nor U1755 (N_1755,In_727,In_546);
and U1756 (N_1756,In_691,In_487);
or U1757 (N_1757,In_253,In_618);
xnor U1758 (N_1758,In_75,In_196);
nor U1759 (N_1759,In_456,In_636);
nand U1760 (N_1760,In_458,In_183);
nor U1761 (N_1761,In_464,In_441);
nor U1762 (N_1762,In_235,In_132);
xnor U1763 (N_1763,In_731,In_163);
and U1764 (N_1764,In_52,In_109);
xor U1765 (N_1765,In_664,In_274);
and U1766 (N_1766,In_102,In_301);
and U1767 (N_1767,In_508,In_492);
or U1768 (N_1768,In_209,In_376);
or U1769 (N_1769,In_104,In_639);
nand U1770 (N_1770,In_364,In_122);
xor U1771 (N_1771,In_123,In_182);
nand U1772 (N_1772,In_432,In_646);
xnor U1773 (N_1773,In_379,In_558);
and U1774 (N_1774,In_154,In_166);
or U1775 (N_1775,In_316,In_362);
or U1776 (N_1776,In_45,In_73);
xnor U1777 (N_1777,In_646,In_404);
or U1778 (N_1778,In_339,In_559);
and U1779 (N_1779,In_222,In_553);
nor U1780 (N_1780,In_431,In_508);
or U1781 (N_1781,In_41,In_540);
nor U1782 (N_1782,In_526,In_362);
and U1783 (N_1783,In_357,In_524);
and U1784 (N_1784,In_397,In_366);
nor U1785 (N_1785,In_262,In_476);
or U1786 (N_1786,In_441,In_542);
and U1787 (N_1787,In_455,In_687);
or U1788 (N_1788,In_140,In_597);
or U1789 (N_1789,In_696,In_488);
nand U1790 (N_1790,In_409,In_169);
nand U1791 (N_1791,In_564,In_490);
and U1792 (N_1792,In_636,In_273);
nand U1793 (N_1793,In_304,In_243);
nand U1794 (N_1794,In_656,In_478);
or U1795 (N_1795,In_203,In_598);
nand U1796 (N_1796,In_133,In_522);
nor U1797 (N_1797,In_656,In_703);
and U1798 (N_1798,In_343,In_75);
nand U1799 (N_1799,In_152,In_64);
and U1800 (N_1800,In_736,In_497);
nor U1801 (N_1801,In_118,In_553);
and U1802 (N_1802,In_732,In_296);
and U1803 (N_1803,In_600,In_24);
xnor U1804 (N_1804,In_470,In_332);
xor U1805 (N_1805,In_672,In_355);
and U1806 (N_1806,In_708,In_297);
or U1807 (N_1807,In_105,In_548);
nand U1808 (N_1808,In_146,In_597);
nor U1809 (N_1809,In_340,In_561);
nand U1810 (N_1810,In_589,In_169);
xnor U1811 (N_1811,In_0,In_624);
nand U1812 (N_1812,In_77,In_623);
or U1813 (N_1813,In_543,In_673);
nor U1814 (N_1814,In_459,In_30);
and U1815 (N_1815,In_631,In_336);
or U1816 (N_1816,In_581,In_132);
or U1817 (N_1817,In_314,In_118);
or U1818 (N_1818,In_587,In_241);
nand U1819 (N_1819,In_55,In_648);
nand U1820 (N_1820,In_686,In_473);
nand U1821 (N_1821,In_328,In_44);
nand U1822 (N_1822,In_523,In_562);
or U1823 (N_1823,In_3,In_404);
nor U1824 (N_1824,In_15,In_657);
xnor U1825 (N_1825,In_212,In_63);
and U1826 (N_1826,In_161,In_294);
nor U1827 (N_1827,In_329,In_274);
nand U1828 (N_1828,In_12,In_676);
or U1829 (N_1829,In_406,In_61);
nand U1830 (N_1830,In_537,In_732);
nand U1831 (N_1831,In_343,In_626);
and U1832 (N_1832,In_628,In_289);
and U1833 (N_1833,In_720,In_589);
xnor U1834 (N_1834,In_144,In_413);
nor U1835 (N_1835,In_462,In_591);
and U1836 (N_1836,In_233,In_150);
and U1837 (N_1837,In_127,In_150);
and U1838 (N_1838,In_26,In_150);
or U1839 (N_1839,In_373,In_68);
xnor U1840 (N_1840,In_292,In_206);
nand U1841 (N_1841,In_594,In_535);
nand U1842 (N_1842,In_247,In_374);
nand U1843 (N_1843,In_603,In_599);
or U1844 (N_1844,In_349,In_273);
and U1845 (N_1845,In_4,In_551);
or U1846 (N_1846,In_47,In_458);
and U1847 (N_1847,In_69,In_295);
or U1848 (N_1848,In_318,In_445);
nand U1849 (N_1849,In_77,In_18);
nor U1850 (N_1850,In_590,In_150);
nor U1851 (N_1851,In_374,In_74);
or U1852 (N_1852,In_449,In_625);
and U1853 (N_1853,In_237,In_359);
nor U1854 (N_1854,In_559,In_327);
and U1855 (N_1855,In_585,In_2);
or U1856 (N_1856,In_547,In_570);
nor U1857 (N_1857,In_528,In_251);
nand U1858 (N_1858,In_675,In_34);
nand U1859 (N_1859,In_169,In_584);
nand U1860 (N_1860,In_250,In_90);
or U1861 (N_1861,In_630,In_461);
or U1862 (N_1862,In_656,In_690);
xnor U1863 (N_1863,In_542,In_699);
nand U1864 (N_1864,In_237,In_646);
and U1865 (N_1865,In_288,In_93);
or U1866 (N_1866,In_466,In_746);
nor U1867 (N_1867,In_20,In_59);
and U1868 (N_1868,In_235,In_198);
and U1869 (N_1869,In_95,In_418);
xnor U1870 (N_1870,In_42,In_100);
and U1871 (N_1871,In_666,In_369);
nand U1872 (N_1872,In_705,In_731);
nor U1873 (N_1873,In_267,In_326);
nor U1874 (N_1874,In_385,In_112);
nor U1875 (N_1875,In_386,In_745);
nand U1876 (N_1876,In_346,In_168);
or U1877 (N_1877,In_472,In_308);
and U1878 (N_1878,In_606,In_276);
nand U1879 (N_1879,In_219,In_21);
xor U1880 (N_1880,In_95,In_734);
or U1881 (N_1881,In_612,In_748);
nand U1882 (N_1882,In_171,In_258);
nand U1883 (N_1883,In_586,In_40);
or U1884 (N_1884,In_532,In_143);
nor U1885 (N_1885,In_433,In_698);
nand U1886 (N_1886,In_566,In_263);
or U1887 (N_1887,In_584,In_298);
nand U1888 (N_1888,In_61,In_569);
nand U1889 (N_1889,In_30,In_572);
nand U1890 (N_1890,In_307,In_552);
nand U1891 (N_1891,In_119,In_472);
and U1892 (N_1892,In_508,In_243);
nand U1893 (N_1893,In_275,In_426);
nand U1894 (N_1894,In_458,In_706);
nand U1895 (N_1895,In_168,In_731);
and U1896 (N_1896,In_450,In_340);
xor U1897 (N_1897,In_690,In_192);
nand U1898 (N_1898,In_641,In_648);
nand U1899 (N_1899,In_454,In_733);
and U1900 (N_1900,In_14,In_236);
or U1901 (N_1901,In_688,In_364);
or U1902 (N_1902,In_331,In_474);
nand U1903 (N_1903,In_29,In_369);
nand U1904 (N_1904,In_661,In_377);
nand U1905 (N_1905,In_491,In_650);
or U1906 (N_1906,In_425,In_687);
or U1907 (N_1907,In_273,In_550);
and U1908 (N_1908,In_426,In_693);
nor U1909 (N_1909,In_606,In_275);
nor U1910 (N_1910,In_101,In_237);
or U1911 (N_1911,In_287,In_655);
or U1912 (N_1912,In_625,In_596);
and U1913 (N_1913,In_304,In_721);
or U1914 (N_1914,In_123,In_541);
xor U1915 (N_1915,In_323,In_263);
xnor U1916 (N_1916,In_604,In_733);
nand U1917 (N_1917,In_398,In_411);
nand U1918 (N_1918,In_279,In_636);
and U1919 (N_1919,In_678,In_53);
and U1920 (N_1920,In_690,In_342);
nand U1921 (N_1921,In_145,In_372);
and U1922 (N_1922,In_240,In_531);
nor U1923 (N_1923,In_410,In_203);
and U1924 (N_1924,In_730,In_444);
nand U1925 (N_1925,In_291,In_96);
nand U1926 (N_1926,In_119,In_2);
nand U1927 (N_1927,In_148,In_163);
nor U1928 (N_1928,In_310,In_635);
or U1929 (N_1929,In_71,In_7);
xnor U1930 (N_1930,In_437,In_622);
or U1931 (N_1931,In_101,In_250);
or U1932 (N_1932,In_526,In_303);
nor U1933 (N_1933,In_146,In_350);
or U1934 (N_1934,In_695,In_68);
and U1935 (N_1935,In_571,In_637);
nor U1936 (N_1936,In_181,In_631);
or U1937 (N_1937,In_635,In_173);
or U1938 (N_1938,In_82,In_571);
and U1939 (N_1939,In_24,In_545);
xnor U1940 (N_1940,In_156,In_622);
nand U1941 (N_1941,In_26,In_317);
and U1942 (N_1942,In_744,In_474);
or U1943 (N_1943,In_196,In_233);
or U1944 (N_1944,In_659,In_476);
nor U1945 (N_1945,In_445,In_425);
or U1946 (N_1946,In_466,In_106);
nor U1947 (N_1947,In_667,In_125);
nor U1948 (N_1948,In_145,In_721);
nand U1949 (N_1949,In_642,In_408);
or U1950 (N_1950,In_423,In_305);
nand U1951 (N_1951,In_209,In_661);
nor U1952 (N_1952,In_218,In_318);
and U1953 (N_1953,In_254,In_518);
nand U1954 (N_1954,In_125,In_246);
nor U1955 (N_1955,In_685,In_568);
and U1956 (N_1956,In_570,In_157);
nand U1957 (N_1957,In_289,In_596);
or U1958 (N_1958,In_288,In_655);
nor U1959 (N_1959,In_735,In_25);
nand U1960 (N_1960,In_178,In_88);
and U1961 (N_1961,In_423,In_526);
nor U1962 (N_1962,In_286,In_692);
and U1963 (N_1963,In_499,In_340);
nor U1964 (N_1964,In_546,In_203);
and U1965 (N_1965,In_697,In_160);
and U1966 (N_1966,In_634,In_552);
nand U1967 (N_1967,In_144,In_279);
or U1968 (N_1968,In_551,In_113);
and U1969 (N_1969,In_603,In_566);
or U1970 (N_1970,In_302,In_149);
nand U1971 (N_1971,In_443,In_722);
nand U1972 (N_1972,In_105,In_351);
and U1973 (N_1973,In_363,In_333);
and U1974 (N_1974,In_536,In_182);
nand U1975 (N_1975,In_570,In_332);
xor U1976 (N_1976,In_307,In_220);
xor U1977 (N_1977,In_298,In_88);
nand U1978 (N_1978,In_345,In_39);
or U1979 (N_1979,In_219,In_521);
and U1980 (N_1980,In_233,In_518);
or U1981 (N_1981,In_425,In_168);
nor U1982 (N_1982,In_634,In_350);
xnor U1983 (N_1983,In_44,In_512);
and U1984 (N_1984,In_393,In_546);
or U1985 (N_1985,In_525,In_636);
nand U1986 (N_1986,In_486,In_507);
nand U1987 (N_1987,In_286,In_408);
nor U1988 (N_1988,In_616,In_424);
and U1989 (N_1989,In_737,In_731);
and U1990 (N_1990,In_313,In_377);
and U1991 (N_1991,In_458,In_290);
nand U1992 (N_1992,In_718,In_372);
and U1993 (N_1993,In_719,In_396);
nor U1994 (N_1994,In_260,In_137);
and U1995 (N_1995,In_401,In_551);
or U1996 (N_1996,In_571,In_225);
nor U1997 (N_1997,In_46,In_388);
nor U1998 (N_1998,In_513,In_246);
nor U1999 (N_1999,In_693,In_605);
or U2000 (N_2000,In_552,In_697);
and U2001 (N_2001,In_13,In_233);
nor U2002 (N_2002,In_687,In_283);
nor U2003 (N_2003,In_548,In_218);
and U2004 (N_2004,In_387,In_676);
and U2005 (N_2005,In_27,In_425);
and U2006 (N_2006,In_288,In_736);
and U2007 (N_2007,In_490,In_723);
or U2008 (N_2008,In_36,In_648);
xnor U2009 (N_2009,In_149,In_43);
and U2010 (N_2010,In_328,In_433);
or U2011 (N_2011,In_497,In_280);
nand U2012 (N_2012,In_390,In_720);
nor U2013 (N_2013,In_236,In_239);
or U2014 (N_2014,In_416,In_652);
xor U2015 (N_2015,In_572,In_582);
or U2016 (N_2016,In_672,In_216);
or U2017 (N_2017,In_140,In_738);
nand U2018 (N_2018,In_539,In_360);
or U2019 (N_2019,In_680,In_522);
nor U2020 (N_2020,In_421,In_319);
or U2021 (N_2021,In_35,In_138);
and U2022 (N_2022,In_676,In_116);
nor U2023 (N_2023,In_62,In_212);
or U2024 (N_2024,In_451,In_230);
xor U2025 (N_2025,In_739,In_550);
nor U2026 (N_2026,In_656,In_520);
xor U2027 (N_2027,In_445,In_504);
or U2028 (N_2028,In_261,In_316);
nand U2029 (N_2029,In_516,In_249);
nand U2030 (N_2030,In_383,In_724);
or U2031 (N_2031,In_266,In_730);
nor U2032 (N_2032,In_666,In_219);
xnor U2033 (N_2033,In_256,In_155);
nand U2034 (N_2034,In_141,In_225);
nor U2035 (N_2035,In_468,In_155);
nor U2036 (N_2036,In_472,In_695);
nand U2037 (N_2037,In_482,In_119);
or U2038 (N_2038,In_259,In_437);
xnor U2039 (N_2039,In_372,In_538);
and U2040 (N_2040,In_561,In_101);
nor U2041 (N_2041,In_579,In_526);
nand U2042 (N_2042,In_131,In_626);
xor U2043 (N_2043,In_450,In_46);
nor U2044 (N_2044,In_576,In_749);
or U2045 (N_2045,In_309,In_28);
xnor U2046 (N_2046,In_532,In_99);
and U2047 (N_2047,In_273,In_322);
or U2048 (N_2048,In_691,In_78);
and U2049 (N_2049,In_118,In_356);
nor U2050 (N_2050,In_16,In_422);
or U2051 (N_2051,In_477,In_617);
nor U2052 (N_2052,In_725,In_693);
and U2053 (N_2053,In_720,In_593);
nor U2054 (N_2054,In_239,In_449);
nand U2055 (N_2055,In_207,In_194);
or U2056 (N_2056,In_54,In_570);
or U2057 (N_2057,In_54,In_328);
nor U2058 (N_2058,In_41,In_187);
nor U2059 (N_2059,In_692,In_166);
and U2060 (N_2060,In_120,In_505);
nand U2061 (N_2061,In_743,In_484);
or U2062 (N_2062,In_331,In_506);
xnor U2063 (N_2063,In_13,In_385);
nand U2064 (N_2064,In_658,In_539);
or U2065 (N_2065,In_140,In_218);
and U2066 (N_2066,In_115,In_677);
nand U2067 (N_2067,In_179,In_238);
nand U2068 (N_2068,In_742,In_120);
nor U2069 (N_2069,In_528,In_49);
and U2070 (N_2070,In_598,In_396);
and U2071 (N_2071,In_603,In_219);
or U2072 (N_2072,In_58,In_257);
nand U2073 (N_2073,In_748,In_467);
nor U2074 (N_2074,In_455,In_464);
nor U2075 (N_2075,In_386,In_509);
nand U2076 (N_2076,In_178,In_75);
and U2077 (N_2077,In_634,In_310);
or U2078 (N_2078,In_491,In_307);
nand U2079 (N_2079,In_671,In_351);
nor U2080 (N_2080,In_120,In_97);
xnor U2081 (N_2081,In_431,In_501);
or U2082 (N_2082,In_191,In_150);
and U2083 (N_2083,In_623,In_449);
nand U2084 (N_2084,In_391,In_242);
xnor U2085 (N_2085,In_417,In_269);
and U2086 (N_2086,In_218,In_160);
or U2087 (N_2087,In_446,In_435);
nand U2088 (N_2088,In_688,In_708);
nand U2089 (N_2089,In_125,In_309);
nand U2090 (N_2090,In_605,In_93);
and U2091 (N_2091,In_345,In_598);
nor U2092 (N_2092,In_455,In_398);
or U2093 (N_2093,In_701,In_562);
or U2094 (N_2094,In_683,In_457);
nor U2095 (N_2095,In_25,In_419);
and U2096 (N_2096,In_323,In_493);
nor U2097 (N_2097,In_509,In_11);
or U2098 (N_2098,In_364,In_205);
or U2099 (N_2099,In_736,In_123);
and U2100 (N_2100,In_32,In_665);
nand U2101 (N_2101,In_180,In_681);
or U2102 (N_2102,In_334,In_28);
or U2103 (N_2103,In_59,In_156);
or U2104 (N_2104,In_444,In_280);
or U2105 (N_2105,In_379,In_8);
nor U2106 (N_2106,In_317,In_61);
nor U2107 (N_2107,In_1,In_456);
or U2108 (N_2108,In_385,In_307);
and U2109 (N_2109,In_95,In_130);
nand U2110 (N_2110,In_606,In_657);
nor U2111 (N_2111,In_479,In_377);
nor U2112 (N_2112,In_523,In_645);
nor U2113 (N_2113,In_456,In_17);
and U2114 (N_2114,In_384,In_295);
nor U2115 (N_2115,In_570,In_445);
or U2116 (N_2116,In_600,In_295);
nand U2117 (N_2117,In_674,In_565);
or U2118 (N_2118,In_243,In_559);
nor U2119 (N_2119,In_135,In_723);
or U2120 (N_2120,In_532,In_332);
nand U2121 (N_2121,In_381,In_287);
and U2122 (N_2122,In_730,In_249);
nor U2123 (N_2123,In_654,In_0);
or U2124 (N_2124,In_147,In_451);
nor U2125 (N_2125,In_617,In_432);
nand U2126 (N_2126,In_169,In_494);
or U2127 (N_2127,In_63,In_697);
nor U2128 (N_2128,In_347,In_346);
xor U2129 (N_2129,In_124,In_302);
nand U2130 (N_2130,In_226,In_592);
or U2131 (N_2131,In_71,In_175);
and U2132 (N_2132,In_137,In_543);
or U2133 (N_2133,In_358,In_500);
xor U2134 (N_2134,In_75,In_324);
xor U2135 (N_2135,In_323,In_577);
or U2136 (N_2136,In_739,In_660);
or U2137 (N_2137,In_326,In_680);
nor U2138 (N_2138,In_520,In_41);
or U2139 (N_2139,In_277,In_195);
and U2140 (N_2140,In_748,In_584);
or U2141 (N_2141,In_239,In_675);
and U2142 (N_2142,In_5,In_551);
or U2143 (N_2143,In_668,In_276);
or U2144 (N_2144,In_713,In_428);
or U2145 (N_2145,In_51,In_73);
or U2146 (N_2146,In_681,In_495);
or U2147 (N_2147,In_240,In_28);
nor U2148 (N_2148,In_315,In_28);
nand U2149 (N_2149,In_593,In_715);
nor U2150 (N_2150,In_347,In_226);
and U2151 (N_2151,In_495,In_527);
nand U2152 (N_2152,In_459,In_333);
and U2153 (N_2153,In_29,In_253);
nand U2154 (N_2154,In_377,In_182);
xor U2155 (N_2155,In_66,In_639);
and U2156 (N_2156,In_170,In_594);
nand U2157 (N_2157,In_630,In_221);
xor U2158 (N_2158,In_188,In_504);
or U2159 (N_2159,In_516,In_272);
and U2160 (N_2160,In_33,In_717);
and U2161 (N_2161,In_69,In_555);
nor U2162 (N_2162,In_625,In_569);
nand U2163 (N_2163,In_683,In_233);
and U2164 (N_2164,In_98,In_282);
and U2165 (N_2165,In_21,In_444);
and U2166 (N_2166,In_685,In_226);
nand U2167 (N_2167,In_565,In_496);
or U2168 (N_2168,In_518,In_544);
nor U2169 (N_2169,In_501,In_711);
xor U2170 (N_2170,In_724,In_114);
and U2171 (N_2171,In_314,In_376);
or U2172 (N_2172,In_565,In_164);
or U2173 (N_2173,In_351,In_385);
nor U2174 (N_2174,In_335,In_403);
and U2175 (N_2175,In_38,In_132);
and U2176 (N_2176,In_281,In_688);
or U2177 (N_2177,In_253,In_16);
nor U2178 (N_2178,In_296,In_662);
xnor U2179 (N_2179,In_29,In_343);
nor U2180 (N_2180,In_679,In_492);
and U2181 (N_2181,In_564,In_340);
and U2182 (N_2182,In_511,In_130);
nand U2183 (N_2183,In_445,In_64);
and U2184 (N_2184,In_118,In_280);
nor U2185 (N_2185,In_332,In_200);
nor U2186 (N_2186,In_41,In_492);
nor U2187 (N_2187,In_78,In_451);
and U2188 (N_2188,In_736,In_712);
xnor U2189 (N_2189,In_633,In_252);
nand U2190 (N_2190,In_433,In_488);
and U2191 (N_2191,In_333,In_340);
nor U2192 (N_2192,In_243,In_165);
and U2193 (N_2193,In_409,In_445);
or U2194 (N_2194,In_641,In_632);
xor U2195 (N_2195,In_307,In_170);
and U2196 (N_2196,In_626,In_117);
or U2197 (N_2197,In_579,In_644);
nor U2198 (N_2198,In_66,In_504);
and U2199 (N_2199,In_169,In_497);
or U2200 (N_2200,In_94,In_538);
or U2201 (N_2201,In_360,In_341);
nand U2202 (N_2202,In_369,In_51);
xor U2203 (N_2203,In_112,In_85);
nor U2204 (N_2204,In_84,In_215);
and U2205 (N_2205,In_43,In_360);
nand U2206 (N_2206,In_740,In_40);
nand U2207 (N_2207,In_101,In_422);
nand U2208 (N_2208,In_87,In_609);
and U2209 (N_2209,In_402,In_628);
nor U2210 (N_2210,In_9,In_689);
nor U2211 (N_2211,In_438,In_286);
nor U2212 (N_2212,In_550,In_142);
and U2213 (N_2213,In_11,In_154);
nand U2214 (N_2214,In_91,In_436);
nand U2215 (N_2215,In_97,In_511);
nor U2216 (N_2216,In_1,In_634);
nand U2217 (N_2217,In_172,In_397);
or U2218 (N_2218,In_232,In_647);
and U2219 (N_2219,In_273,In_744);
or U2220 (N_2220,In_434,In_455);
and U2221 (N_2221,In_175,In_254);
and U2222 (N_2222,In_562,In_187);
and U2223 (N_2223,In_247,In_483);
or U2224 (N_2224,In_614,In_261);
or U2225 (N_2225,In_104,In_534);
and U2226 (N_2226,In_454,In_470);
or U2227 (N_2227,In_576,In_278);
and U2228 (N_2228,In_598,In_526);
xnor U2229 (N_2229,In_112,In_479);
or U2230 (N_2230,In_326,In_528);
nand U2231 (N_2231,In_694,In_60);
and U2232 (N_2232,In_421,In_566);
or U2233 (N_2233,In_527,In_748);
and U2234 (N_2234,In_130,In_662);
and U2235 (N_2235,In_66,In_677);
nand U2236 (N_2236,In_72,In_347);
nor U2237 (N_2237,In_669,In_536);
or U2238 (N_2238,In_219,In_150);
nor U2239 (N_2239,In_702,In_350);
or U2240 (N_2240,In_687,In_405);
and U2241 (N_2241,In_404,In_146);
nand U2242 (N_2242,In_128,In_195);
nor U2243 (N_2243,In_716,In_591);
or U2244 (N_2244,In_711,In_85);
and U2245 (N_2245,In_585,In_567);
xor U2246 (N_2246,In_619,In_172);
xnor U2247 (N_2247,In_104,In_507);
nand U2248 (N_2248,In_361,In_158);
nor U2249 (N_2249,In_84,In_136);
or U2250 (N_2250,In_160,In_205);
and U2251 (N_2251,In_574,In_353);
nand U2252 (N_2252,In_184,In_94);
xnor U2253 (N_2253,In_223,In_607);
xnor U2254 (N_2254,In_313,In_251);
or U2255 (N_2255,In_694,In_28);
nand U2256 (N_2256,In_641,In_314);
or U2257 (N_2257,In_568,In_454);
nand U2258 (N_2258,In_575,In_192);
and U2259 (N_2259,In_237,In_172);
or U2260 (N_2260,In_57,In_736);
nor U2261 (N_2261,In_109,In_31);
and U2262 (N_2262,In_262,In_459);
nand U2263 (N_2263,In_161,In_225);
nand U2264 (N_2264,In_79,In_437);
or U2265 (N_2265,In_428,In_688);
and U2266 (N_2266,In_731,In_160);
xnor U2267 (N_2267,In_41,In_583);
nand U2268 (N_2268,In_161,In_4);
nand U2269 (N_2269,In_705,In_36);
or U2270 (N_2270,In_127,In_15);
nor U2271 (N_2271,In_337,In_746);
xnor U2272 (N_2272,In_739,In_113);
nor U2273 (N_2273,In_383,In_126);
and U2274 (N_2274,In_533,In_128);
nand U2275 (N_2275,In_7,In_229);
nand U2276 (N_2276,In_663,In_124);
or U2277 (N_2277,In_384,In_712);
nor U2278 (N_2278,In_378,In_109);
and U2279 (N_2279,In_474,In_551);
nor U2280 (N_2280,In_335,In_454);
nand U2281 (N_2281,In_352,In_342);
or U2282 (N_2282,In_663,In_746);
nand U2283 (N_2283,In_672,In_383);
nand U2284 (N_2284,In_188,In_646);
nand U2285 (N_2285,In_31,In_385);
nand U2286 (N_2286,In_100,In_441);
xnor U2287 (N_2287,In_380,In_383);
or U2288 (N_2288,In_446,In_186);
nor U2289 (N_2289,In_727,In_630);
nand U2290 (N_2290,In_469,In_574);
nor U2291 (N_2291,In_342,In_357);
or U2292 (N_2292,In_475,In_80);
or U2293 (N_2293,In_99,In_284);
and U2294 (N_2294,In_460,In_439);
and U2295 (N_2295,In_324,In_542);
and U2296 (N_2296,In_323,In_434);
nor U2297 (N_2297,In_243,In_621);
nor U2298 (N_2298,In_713,In_360);
or U2299 (N_2299,In_431,In_486);
or U2300 (N_2300,In_459,In_196);
or U2301 (N_2301,In_543,In_349);
or U2302 (N_2302,In_489,In_300);
and U2303 (N_2303,In_8,In_553);
nor U2304 (N_2304,In_430,In_140);
or U2305 (N_2305,In_46,In_479);
nand U2306 (N_2306,In_75,In_371);
nor U2307 (N_2307,In_120,In_368);
nor U2308 (N_2308,In_483,In_416);
and U2309 (N_2309,In_381,In_220);
or U2310 (N_2310,In_406,In_298);
nor U2311 (N_2311,In_485,In_386);
nand U2312 (N_2312,In_608,In_302);
nor U2313 (N_2313,In_110,In_40);
or U2314 (N_2314,In_218,In_429);
nand U2315 (N_2315,In_703,In_580);
nand U2316 (N_2316,In_90,In_272);
nor U2317 (N_2317,In_511,In_301);
or U2318 (N_2318,In_152,In_226);
and U2319 (N_2319,In_375,In_680);
xnor U2320 (N_2320,In_512,In_448);
or U2321 (N_2321,In_123,In_208);
xnor U2322 (N_2322,In_574,In_590);
nor U2323 (N_2323,In_285,In_343);
xor U2324 (N_2324,In_357,In_173);
and U2325 (N_2325,In_81,In_149);
and U2326 (N_2326,In_362,In_450);
nand U2327 (N_2327,In_126,In_251);
xor U2328 (N_2328,In_477,In_17);
or U2329 (N_2329,In_474,In_556);
nand U2330 (N_2330,In_53,In_627);
nor U2331 (N_2331,In_219,In_579);
or U2332 (N_2332,In_732,In_556);
and U2333 (N_2333,In_578,In_326);
xor U2334 (N_2334,In_484,In_398);
or U2335 (N_2335,In_451,In_453);
xnor U2336 (N_2336,In_130,In_520);
or U2337 (N_2337,In_643,In_220);
and U2338 (N_2338,In_107,In_645);
nor U2339 (N_2339,In_88,In_398);
and U2340 (N_2340,In_191,In_188);
and U2341 (N_2341,In_423,In_401);
nand U2342 (N_2342,In_64,In_309);
and U2343 (N_2343,In_261,In_286);
and U2344 (N_2344,In_230,In_642);
nor U2345 (N_2345,In_520,In_310);
and U2346 (N_2346,In_592,In_486);
nor U2347 (N_2347,In_115,In_716);
and U2348 (N_2348,In_269,In_622);
and U2349 (N_2349,In_610,In_426);
nand U2350 (N_2350,In_280,In_426);
or U2351 (N_2351,In_357,In_106);
or U2352 (N_2352,In_496,In_347);
xnor U2353 (N_2353,In_365,In_415);
nor U2354 (N_2354,In_639,In_430);
and U2355 (N_2355,In_745,In_410);
nand U2356 (N_2356,In_353,In_140);
or U2357 (N_2357,In_47,In_413);
nor U2358 (N_2358,In_424,In_133);
xor U2359 (N_2359,In_272,In_521);
and U2360 (N_2360,In_485,In_607);
xor U2361 (N_2361,In_714,In_527);
or U2362 (N_2362,In_530,In_146);
nor U2363 (N_2363,In_290,In_537);
nand U2364 (N_2364,In_7,In_352);
or U2365 (N_2365,In_466,In_299);
or U2366 (N_2366,In_356,In_97);
xnor U2367 (N_2367,In_495,In_130);
and U2368 (N_2368,In_231,In_661);
nor U2369 (N_2369,In_221,In_214);
nor U2370 (N_2370,In_12,In_308);
nor U2371 (N_2371,In_299,In_78);
or U2372 (N_2372,In_383,In_13);
xor U2373 (N_2373,In_360,In_542);
nor U2374 (N_2374,In_183,In_126);
and U2375 (N_2375,In_143,In_19);
or U2376 (N_2376,In_72,In_658);
xnor U2377 (N_2377,In_617,In_62);
and U2378 (N_2378,In_285,In_536);
nor U2379 (N_2379,In_203,In_381);
xor U2380 (N_2380,In_487,In_24);
nor U2381 (N_2381,In_203,In_143);
nor U2382 (N_2382,In_593,In_675);
xor U2383 (N_2383,In_160,In_703);
nand U2384 (N_2384,In_484,In_303);
nand U2385 (N_2385,In_653,In_142);
and U2386 (N_2386,In_171,In_550);
nand U2387 (N_2387,In_624,In_429);
nand U2388 (N_2388,In_411,In_351);
nor U2389 (N_2389,In_350,In_442);
xnor U2390 (N_2390,In_265,In_392);
or U2391 (N_2391,In_234,In_588);
nand U2392 (N_2392,In_172,In_81);
or U2393 (N_2393,In_109,In_538);
or U2394 (N_2394,In_354,In_511);
or U2395 (N_2395,In_254,In_618);
or U2396 (N_2396,In_730,In_426);
nor U2397 (N_2397,In_203,In_302);
and U2398 (N_2398,In_539,In_238);
or U2399 (N_2399,In_478,In_62);
nand U2400 (N_2400,In_342,In_205);
nor U2401 (N_2401,In_361,In_283);
or U2402 (N_2402,In_63,In_217);
xnor U2403 (N_2403,In_549,In_433);
or U2404 (N_2404,In_301,In_724);
and U2405 (N_2405,In_84,In_692);
nand U2406 (N_2406,In_599,In_36);
and U2407 (N_2407,In_314,In_125);
or U2408 (N_2408,In_655,In_589);
or U2409 (N_2409,In_405,In_703);
or U2410 (N_2410,In_459,In_359);
nor U2411 (N_2411,In_400,In_204);
or U2412 (N_2412,In_88,In_257);
and U2413 (N_2413,In_49,In_187);
or U2414 (N_2414,In_67,In_592);
or U2415 (N_2415,In_442,In_423);
nor U2416 (N_2416,In_255,In_39);
and U2417 (N_2417,In_296,In_617);
nand U2418 (N_2418,In_92,In_269);
nand U2419 (N_2419,In_535,In_104);
nand U2420 (N_2420,In_92,In_94);
and U2421 (N_2421,In_30,In_694);
nor U2422 (N_2422,In_265,In_415);
and U2423 (N_2423,In_647,In_138);
and U2424 (N_2424,In_46,In_293);
or U2425 (N_2425,In_694,In_639);
nand U2426 (N_2426,In_61,In_58);
nand U2427 (N_2427,In_185,In_310);
nand U2428 (N_2428,In_368,In_11);
or U2429 (N_2429,In_564,In_685);
nor U2430 (N_2430,In_430,In_425);
or U2431 (N_2431,In_302,In_274);
xnor U2432 (N_2432,In_488,In_245);
or U2433 (N_2433,In_439,In_381);
xor U2434 (N_2434,In_345,In_442);
nand U2435 (N_2435,In_142,In_8);
nand U2436 (N_2436,In_619,In_656);
or U2437 (N_2437,In_214,In_690);
nand U2438 (N_2438,In_380,In_262);
and U2439 (N_2439,In_374,In_325);
nor U2440 (N_2440,In_735,In_329);
and U2441 (N_2441,In_79,In_153);
nand U2442 (N_2442,In_3,In_9);
nand U2443 (N_2443,In_396,In_427);
and U2444 (N_2444,In_28,In_192);
nor U2445 (N_2445,In_655,In_620);
or U2446 (N_2446,In_619,In_99);
or U2447 (N_2447,In_447,In_616);
xor U2448 (N_2448,In_482,In_165);
nor U2449 (N_2449,In_703,In_531);
and U2450 (N_2450,In_392,In_617);
or U2451 (N_2451,In_165,In_240);
or U2452 (N_2452,In_324,In_566);
xnor U2453 (N_2453,In_315,In_732);
and U2454 (N_2454,In_608,In_203);
xor U2455 (N_2455,In_614,In_538);
and U2456 (N_2456,In_177,In_395);
nor U2457 (N_2457,In_479,In_666);
and U2458 (N_2458,In_313,In_546);
and U2459 (N_2459,In_740,In_728);
or U2460 (N_2460,In_147,In_644);
xnor U2461 (N_2461,In_133,In_74);
or U2462 (N_2462,In_139,In_744);
nand U2463 (N_2463,In_494,In_120);
or U2464 (N_2464,In_196,In_235);
nand U2465 (N_2465,In_351,In_610);
xnor U2466 (N_2466,In_427,In_312);
and U2467 (N_2467,In_69,In_542);
or U2468 (N_2468,In_503,In_668);
and U2469 (N_2469,In_702,In_716);
nor U2470 (N_2470,In_418,In_581);
or U2471 (N_2471,In_428,In_597);
nand U2472 (N_2472,In_314,In_365);
nor U2473 (N_2473,In_72,In_201);
nand U2474 (N_2474,In_356,In_576);
nor U2475 (N_2475,In_121,In_253);
and U2476 (N_2476,In_326,In_600);
nand U2477 (N_2477,In_386,In_383);
nor U2478 (N_2478,In_416,In_282);
and U2479 (N_2479,In_364,In_492);
and U2480 (N_2480,In_102,In_649);
nor U2481 (N_2481,In_553,In_192);
xnor U2482 (N_2482,In_383,In_701);
or U2483 (N_2483,In_277,In_568);
or U2484 (N_2484,In_410,In_67);
nor U2485 (N_2485,In_109,In_589);
or U2486 (N_2486,In_173,In_433);
nor U2487 (N_2487,In_4,In_224);
and U2488 (N_2488,In_691,In_377);
nand U2489 (N_2489,In_186,In_643);
and U2490 (N_2490,In_144,In_737);
or U2491 (N_2491,In_348,In_420);
and U2492 (N_2492,In_575,In_395);
or U2493 (N_2493,In_720,In_695);
nand U2494 (N_2494,In_47,In_663);
nand U2495 (N_2495,In_581,In_252);
nand U2496 (N_2496,In_311,In_265);
nor U2497 (N_2497,In_649,In_121);
nand U2498 (N_2498,In_403,In_727);
nand U2499 (N_2499,In_615,In_462);
nand U2500 (N_2500,N_1247,N_1193);
and U2501 (N_2501,N_1645,N_1889);
and U2502 (N_2502,N_725,N_1757);
nor U2503 (N_2503,N_267,N_2491);
and U2504 (N_2504,N_2391,N_332);
or U2505 (N_2505,N_2123,N_620);
nand U2506 (N_2506,N_1235,N_1002);
xor U2507 (N_2507,N_236,N_1709);
nor U2508 (N_2508,N_2397,N_1163);
or U2509 (N_2509,N_1839,N_1483);
and U2510 (N_2510,N_2335,N_1212);
nand U2511 (N_2511,N_1040,N_1975);
or U2512 (N_2512,N_276,N_52);
or U2513 (N_2513,N_122,N_526);
xnor U2514 (N_2514,N_1632,N_1367);
and U2515 (N_2515,N_319,N_462);
nor U2516 (N_2516,N_694,N_1359);
nand U2517 (N_2517,N_1157,N_1722);
nor U2518 (N_2518,N_898,N_443);
or U2519 (N_2519,N_1250,N_514);
and U2520 (N_2520,N_958,N_869);
nand U2521 (N_2521,N_1023,N_616);
nor U2522 (N_2522,N_504,N_1737);
or U2523 (N_2523,N_1291,N_1276);
and U2524 (N_2524,N_2196,N_818);
nand U2525 (N_2525,N_1734,N_1039);
nor U2526 (N_2526,N_25,N_2294);
nor U2527 (N_2527,N_1617,N_2314);
and U2528 (N_2528,N_348,N_341);
or U2529 (N_2529,N_2330,N_2437);
xnor U2530 (N_2530,N_1350,N_1444);
xnor U2531 (N_2531,N_2119,N_1517);
nand U2532 (N_2532,N_160,N_2244);
nand U2533 (N_2533,N_2031,N_237);
xnor U2534 (N_2534,N_1431,N_248);
nor U2535 (N_2535,N_1977,N_290);
nor U2536 (N_2536,N_2304,N_496);
or U2537 (N_2537,N_2452,N_5);
and U2538 (N_2538,N_366,N_1510);
nor U2539 (N_2539,N_2435,N_82);
nor U2540 (N_2540,N_2190,N_2469);
and U2541 (N_2541,N_603,N_989);
and U2542 (N_2542,N_2212,N_1602);
and U2543 (N_2543,N_1500,N_796);
nor U2544 (N_2544,N_1861,N_136);
or U2545 (N_2545,N_217,N_476);
or U2546 (N_2546,N_1448,N_895);
nor U2547 (N_2547,N_2178,N_1735);
or U2548 (N_2548,N_2310,N_921);
and U2549 (N_2549,N_1999,N_437);
nand U2550 (N_2550,N_1112,N_394);
and U2551 (N_2551,N_790,N_1683);
or U2552 (N_2552,N_892,N_1376);
or U2553 (N_2553,N_836,N_2456);
xor U2554 (N_2554,N_37,N_1091);
and U2555 (N_2555,N_153,N_2414);
or U2556 (N_2556,N_2027,N_765);
or U2557 (N_2557,N_527,N_1195);
xor U2558 (N_2558,N_1534,N_256);
nand U2559 (N_2559,N_2166,N_517);
or U2560 (N_2560,N_841,N_2409);
nand U2561 (N_2561,N_2353,N_710);
nand U2562 (N_2562,N_1729,N_1689);
xnor U2563 (N_2563,N_2405,N_1566);
or U2564 (N_2564,N_465,N_2361);
xor U2565 (N_2565,N_251,N_975);
nor U2566 (N_2566,N_752,N_2352);
xnor U2567 (N_2567,N_2245,N_600);
or U2568 (N_2568,N_2417,N_936);
xor U2569 (N_2569,N_241,N_1362);
nor U2570 (N_2570,N_684,N_970);
nand U2571 (N_2571,N_1875,N_402);
nor U2572 (N_2572,N_1493,N_809);
or U2573 (N_2573,N_583,N_1322);
and U2574 (N_2574,N_1259,N_2217);
or U2575 (N_2575,N_408,N_1760);
xnor U2576 (N_2576,N_1469,N_1671);
nor U2577 (N_2577,N_2264,N_58);
or U2578 (N_2578,N_2458,N_967);
nand U2579 (N_2579,N_1341,N_1800);
nand U2580 (N_2580,N_424,N_1321);
nor U2581 (N_2581,N_372,N_282);
xor U2582 (N_2582,N_356,N_1255);
nor U2583 (N_2583,N_1430,N_2042);
and U2584 (N_2584,N_1173,N_633);
nand U2585 (N_2585,N_686,N_146);
and U2586 (N_2586,N_1306,N_878);
nor U2587 (N_2587,N_1697,N_473);
or U2588 (N_2588,N_296,N_1959);
nor U2589 (N_2589,N_1663,N_165);
xor U2590 (N_2590,N_157,N_1287);
and U2591 (N_2591,N_1971,N_831);
nand U2592 (N_2592,N_2315,N_1575);
or U2593 (N_2593,N_1010,N_2356);
or U2594 (N_2594,N_284,N_2149);
nand U2595 (N_2595,N_250,N_821);
or U2596 (N_2596,N_1207,N_2343);
nand U2597 (N_2597,N_784,N_1458);
nand U2598 (N_2598,N_877,N_1042);
and U2599 (N_2599,N_938,N_553);
nand U2600 (N_2600,N_763,N_1873);
xnor U2601 (N_2601,N_750,N_935);
nor U2602 (N_2602,N_1147,N_1674);
xor U2603 (N_2603,N_1700,N_1135);
nor U2604 (N_2604,N_390,N_1642);
or U2605 (N_2605,N_1550,N_347);
or U2606 (N_2606,N_1050,N_1107);
nand U2607 (N_2607,N_1857,N_729);
or U2608 (N_2608,N_963,N_180);
or U2609 (N_2609,N_302,N_210);
and U2610 (N_2610,N_2246,N_2348);
or U2611 (N_2611,N_558,N_1423);
xor U2612 (N_2612,N_1634,N_2499);
or U2613 (N_2613,N_977,N_880);
and U2614 (N_2614,N_613,N_354);
and U2615 (N_2615,N_1723,N_2187);
nor U2616 (N_2616,N_1620,N_2043);
nor U2617 (N_2617,N_1636,N_2381);
nand U2618 (N_2618,N_1890,N_676);
or U2619 (N_2619,N_442,N_1878);
xnor U2620 (N_2620,N_2064,N_2215);
or U2621 (N_2621,N_1229,N_1044);
or U2622 (N_2622,N_1568,N_2101);
nand U2623 (N_2623,N_471,N_154);
nand U2624 (N_2624,N_283,N_1797);
nor U2625 (N_2625,N_1985,N_428);
nand U2626 (N_2626,N_1139,N_1599);
and U2627 (N_2627,N_2192,N_1481);
and U2628 (N_2628,N_814,N_1048);
nand U2629 (N_2629,N_619,N_1030);
and U2630 (N_2630,N_1887,N_1673);
and U2631 (N_2631,N_2168,N_682);
or U2632 (N_2632,N_1304,N_2366);
nor U2633 (N_2633,N_1810,N_2307);
nand U2634 (N_2634,N_358,N_1071);
or U2635 (N_2635,N_1931,N_2430);
or U2636 (N_2636,N_2250,N_315);
nand U2637 (N_2637,N_758,N_309);
nor U2638 (N_2638,N_2400,N_2270);
nor U2639 (N_2639,N_946,N_994);
or U2640 (N_2640,N_1144,N_1724);
nor U2641 (N_2641,N_1109,N_1606);
nand U2642 (N_2642,N_1137,N_1505);
or U2643 (N_2643,N_2211,N_1428);
nand U2644 (N_2644,N_1068,N_1134);
nand U2645 (N_2645,N_2200,N_1942);
and U2646 (N_2646,N_274,N_598);
nand U2647 (N_2647,N_1463,N_2005);
or U2648 (N_2648,N_1923,N_324);
or U2649 (N_2649,N_835,N_1509);
or U2650 (N_2650,N_1616,N_990);
nor U2651 (N_2651,N_2312,N_593);
xor U2652 (N_2652,N_1961,N_2401);
xnor U2653 (N_2653,N_571,N_1201);
nor U2654 (N_2654,N_463,N_1949);
and U2655 (N_2655,N_1074,N_965);
and U2656 (N_2656,N_2127,N_1987);
and U2657 (N_2657,N_2240,N_2354);
or U2658 (N_2658,N_1818,N_1282);
nor U2659 (N_2659,N_1929,N_12);
or U2660 (N_2660,N_137,N_705);
nor U2661 (N_2661,N_65,N_645);
or U2662 (N_2662,N_475,N_1824);
xnor U2663 (N_2663,N_1482,N_1946);
xnor U2664 (N_2664,N_901,N_2418);
nand U2665 (N_2665,N_1263,N_131);
and U2666 (N_2666,N_61,N_303);
and U2667 (N_2667,N_1548,N_1556);
and U2668 (N_2668,N_359,N_177);
and U2669 (N_2669,N_1006,N_1274);
nor U2670 (N_2670,N_66,N_149);
and U2671 (N_2671,N_1358,N_2332);
and U2672 (N_2672,N_1669,N_1773);
nand U2673 (N_2673,N_1821,N_461);
xor U2674 (N_2674,N_653,N_1440);
nor U2675 (N_2675,N_1624,N_40);
and U2676 (N_2676,N_2477,N_993);
nand U2677 (N_2677,N_2019,N_1392);
nor U2678 (N_2678,N_2362,N_278);
nand U2679 (N_2679,N_1069,N_2451);
nor U2680 (N_2680,N_574,N_1292);
and U2681 (N_2681,N_14,N_357);
nand U2682 (N_2682,N_49,N_1400);
nor U2683 (N_2683,N_824,N_1202);
or U2684 (N_2684,N_1925,N_1132);
nor U2685 (N_2685,N_124,N_71);
nor U2686 (N_2686,N_484,N_1111);
nand U2687 (N_2687,N_851,N_1191);
nand U2688 (N_2688,N_361,N_451);
nand U2689 (N_2689,N_996,N_2253);
and U2690 (N_2690,N_1795,N_327);
nor U2691 (N_2691,N_807,N_2220);
and U2692 (N_2692,N_2184,N_905);
or U2693 (N_2693,N_1621,N_503);
nand U2694 (N_2694,N_1143,N_2219);
or U2695 (N_2695,N_596,N_1300);
or U2696 (N_2696,N_1403,N_27);
or U2697 (N_2697,N_2191,N_737);
xnor U2698 (N_2698,N_1216,N_445);
and U2699 (N_2699,N_2047,N_486);
nor U2700 (N_2700,N_1982,N_1515);
or U2701 (N_2701,N_709,N_797);
and U2702 (N_2702,N_1348,N_515);
nor U2703 (N_2703,N_1591,N_1768);
nor U2704 (N_2704,N_135,N_1311);
nand U2705 (N_2705,N_1177,N_1969);
and U2706 (N_2706,N_1011,N_1037);
nand U2707 (N_2707,N_1547,N_1651);
nor U2708 (N_2708,N_401,N_1678);
nand U2709 (N_2709,N_1973,N_95);
and U2710 (N_2710,N_1034,N_2285);
or U2711 (N_2711,N_29,N_971);
nand U2712 (N_2712,N_1421,N_1145);
nor U2713 (N_2713,N_1559,N_379);
nor U2714 (N_2714,N_2498,N_539);
or U2715 (N_2715,N_1989,N_1117);
nor U2716 (N_2716,N_239,N_167);
nor U2717 (N_2717,N_2105,N_706);
or U2718 (N_2718,N_1631,N_1708);
and U2719 (N_2719,N_1283,N_806);
nand U2720 (N_2720,N_209,N_1166);
nand U2721 (N_2721,N_531,N_1995);
nand U2722 (N_2722,N_1933,N_1625);
and U2723 (N_2723,N_845,N_1904);
nor U2724 (N_2724,N_2468,N_223);
nor U2725 (N_2725,N_978,N_572);
nor U2726 (N_2726,N_2109,N_2111);
nand U2727 (N_2727,N_2302,N_426);
nor U2728 (N_2728,N_139,N_2049);
nor U2729 (N_2729,N_2298,N_1213);
or U2730 (N_2730,N_1736,N_1628);
nor U2731 (N_2731,N_1600,N_678);
and U2732 (N_2732,N_490,N_2459);
xor U2733 (N_2733,N_279,N_1604);
or U2734 (N_2734,N_2273,N_1520);
nand U2735 (N_2735,N_955,N_1864);
or U2736 (N_2736,N_1523,N_2035);
and U2737 (N_2737,N_1664,N_874);
and U2738 (N_2738,N_1707,N_2053);
nand U2739 (N_2739,N_744,N_182);
nand U2740 (N_2740,N_2470,N_1767);
and U2741 (N_2741,N_128,N_76);
or U2742 (N_2742,N_2207,N_2216);
xor U2743 (N_2743,N_453,N_2331);
nor U2744 (N_2744,N_533,N_1021);
nand U2745 (N_2745,N_232,N_838);
or U2746 (N_2746,N_852,N_2350);
nand U2747 (N_2747,N_138,N_2296);
and U2748 (N_2748,N_998,N_110);
nand U2749 (N_2749,N_1009,N_780);
nand U2750 (N_2750,N_1884,N_2388);
or U2751 (N_2751,N_871,N_675);
nor U2752 (N_2752,N_2083,N_1415);
or U2753 (N_2753,N_1314,N_464);
nand U2754 (N_2754,N_280,N_1964);
nor U2755 (N_2755,N_1972,N_524);
nor U2756 (N_2756,N_1504,N_1590);
and U2757 (N_2757,N_948,N_311);
nand U2758 (N_2758,N_1552,N_470);
nor U2759 (N_2759,N_2463,N_1294);
or U2760 (N_2760,N_1781,N_479);
or U2761 (N_2761,N_2293,N_529);
nand U2762 (N_2762,N_497,N_1332);
or U2763 (N_2763,N_1028,N_1271);
and U2764 (N_2764,N_1115,N_800);
nor U2765 (N_2765,N_339,N_1511);
nand U2766 (N_2766,N_36,N_582);
nand U2767 (N_2767,N_1200,N_1344);
nand U2768 (N_2768,N_1186,N_1179);
or U2769 (N_2769,N_2393,N_519);
nand U2770 (N_2770,N_2428,N_509);
nand U2771 (N_2771,N_2420,N_407);
nand U2772 (N_2772,N_2128,N_1257);
xnor U2773 (N_2773,N_655,N_646);
or U2774 (N_2774,N_828,N_1546);
nor U2775 (N_2775,N_293,N_1033);
and U2776 (N_2776,N_2102,N_244);
nor U2777 (N_2777,N_493,N_170);
or U2778 (N_2778,N_1756,N_634);
or U2779 (N_2779,N_1553,N_2136);
or U2780 (N_2780,N_411,N_1496);
nor U2781 (N_2781,N_1096,N_1439);
or U2782 (N_2782,N_1525,N_1528);
xor U2783 (N_2783,N_939,N_2374);
nand U2784 (N_2784,N_1780,N_132);
nor U2785 (N_2785,N_1089,N_1990);
nand U2786 (N_2786,N_732,N_887);
or U2787 (N_2787,N_2094,N_59);
or U2788 (N_2788,N_2457,N_301);
and U2789 (N_2789,N_155,N_2382);
nor U2790 (N_2790,N_2324,N_1876);
and U2791 (N_2791,N_1805,N_1075);
xor U2792 (N_2792,N_631,N_832);
and U2793 (N_2793,N_2440,N_2096);
nor U2794 (N_2794,N_1097,N_703);
and U2795 (N_2795,N_579,N_2475);
xnor U2796 (N_2796,N_1038,N_2436);
and U2797 (N_2797,N_164,N_1164);
xor U2798 (N_2798,N_875,N_1160);
or U2799 (N_2799,N_789,N_1082);
nand U2800 (N_2800,N_1437,N_2465);
nand U2801 (N_2801,N_950,N_1668);
nor U2802 (N_2802,N_1073,N_1491);
and U2803 (N_2803,N_333,N_1377);
and U2804 (N_2804,N_140,N_1336);
nand U2805 (N_2805,N_39,N_1753);
and U2806 (N_2806,N_367,N_2239);
or U2807 (N_2807,N_18,N_1791);
or U2808 (N_2808,N_1870,N_2197);
and U2809 (N_2809,N_446,N_542);
nor U2810 (N_2810,N_968,N_226);
nand U2811 (N_2811,N_1175,N_2089);
nand U2812 (N_2812,N_208,N_1739);
and U2813 (N_2813,N_528,N_748);
nor U2814 (N_2814,N_1380,N_1586);
and U2815 (N_2815,N_113,N_1869);
nand U2816 (N_2816,N_213,N_1908);
xor U2817 (N_2817,N_107,N_2347);
nor U2818 (N_2818,N_458,N_2448);
and U2819 (N_2819,N_1065,N_1831);
and U2820 (N_2820,N_425,N_100);
nor U2821 (N_2821,N_1842,N_985);
nand U2822 (N_2822,N_2446,N_1225);
nor U2823 (N_2823,N_768,N_242);
xor U2824 (N_2824,N_867,N_696);
nor U2825 (N_2825,N_1574,N_2365);
nor U2826 (N_2826,N_670,N_1778);
or U2827 (N_2827,N_667,N_1360);
xor U2828 (N_2828,N_355,N_441);
and U2829 (N_2829,N_1582,N_1003);
nor U2830 (N_2830,N_536,N_545);
nor U2831 (N_2831,N_2025,N_925);
and U2832 (N_2832,N_816,N_547);
nand U2833 (N_2833,N_1310,N_1531);
xor U2834 (N_2834,N_11,N_611);
nand U2835 (N_2835,N_1474,N_2221);
or U2836 (N_2836,N_2328,N_48);
and U2837 (N_2837,N_1860,N_983);
nand U2838 (N_2838,N_103,N_1436);
and U2839 (N_2839,N_823,N_1124);
and U2840 (N_2840,N_2235,N_1819);
xor U2841 (N_2841,N_1613,N_2069);
nand U2842 (N_2842,N_230,N_84);
nand U2843 (N_2843,N_692,N_1420);
nor U2844 (N_2844,N_1542,N_1701);
xor U2845 (N_2845,N_33,N_1637);
or U2846 (N_2846,N_1058,N_2070);
nand U2847 (N_2847,N_1747,N_1254);
or U2848 (N_2848,N_883,N_2295);
nor U2849 (N_2849,N_1140,N_726);
nand U2850 (N_2850,N_999,N_1623);
and U2851 (N_2851,N_488,N_1168);
or U2852 (N_2852,N_799,N_972);
nand U2853 (N_2853,N_1951,N_2208);
or U2854 (N_2854,N_343,N_2017);
nand U2855 (N_2855,N_1779,N_1221);
nor U2856 (N_2856,N_747,N_8);
xor U2857 (N_2857,N_1885,N_1236);
nand U2858 (N_2858,N_1273,N_576);
and U2859 (N_2859,N_1909,N_2081);
and U2860 (N_2860,N_1279,N_934);
xnor U2861 (N_2861,N_1830,N_1297);
or U2862 (N_2862,N_651,N_1543);
nor U2863 (N_2863,N_200,N_1749);
xor U2864 (N_2864,N_1921,N_2455);
and U2865 (N_2865,N_1782,N_2287);
and U2866 (N_2866,N_487,N_1906);
or U2867 (N_2867,N_1101,N_204);
nand U2868 (N_2868,N_491,N_53);
or U2869 (N_2869,N_417,N_2317);
or U2870 (N_2870,N_1149,N_2021);
or U2871 (N_2871,N_1583,N_1086);
nor U2872 (N_2872,N_2039,N_2008);
and U2873 (N_2873,N_447,N_262);
or U2874 (N_2874,N_1650,N_2198);
and U2875 (N_2875,N_1947,N_1763);
and U2876 (N_2876,N_1385,N_1640);
nand U2877 (N_2877,N_1497,N_2474);
nand U2878 (N_2878,N_219,N_981);
nand U2879 (N_2879,N_1138,N_67);
or U2880 (N_2880,N_1105,N_1232);
nand U2881 (N_2881,N_2398,N_1245);
or U2882 (N_2882,N_2185,N_1347);
or U2883 (N_2883,N_1968,N_489);
nor U2884 (N_2884,N_2218,N_1893);
and U2885 (N_2885,N_728,N_1281);
or U2886 (N_2886,N_1692,N_843);
and U2887 (N_2887,N_227,N_736);
nor U2888 (N_2888,N_2370,N_1465);
or U2889 (N_2889,N_454,N_1217);
and U2890 (N_2890,N_1537,N_1793);
or U2891 (N_2891,N_422,N_1324);
and U2892 (N_2892,N_556,N_1573);
nor U2893 (N_2893,N_1788,N_1379);
nor U2894 (N_2894,N_917,N_387);
nand U2895 (N_2895,N_1644,N_2238);
nand U2896 (N_2896,N_2243,N_1859);
xnor U2897 (N_2897,N_1478,N_1224);
nor U2898 (N_2898,N_117,N_270);
and U2899 (N_2899,N_434,N_2279);
nor U2900 (N_2900,N_2404,N_2416);
nor U2901 (N_2901,N_199,N_586);
nand U2902 (N_2902,N_21,N_1691);
and U2903 (N_2903,N_716,N_142);
nand U2904 (N_2904,N_2041,N_2341);
and U2905 (N_2905,N_1187,N_245);
and U2906 (N_2906,N_2093,N_1316);
nor U2907 (N_2907,N_1529,N_320);
nor U2908 (N_2908,N_1102,N_2326);
nand U2909 (N_2909,N_2303,N_2449);
nor U2910 (N_2910,N_2223,N_1936);
nor U2911 (N_2911,N_1384,N_2308);
and U2912 (N_2912,N_307,N_1506);
nor U2913 (N_2913,N_2020,N_1832);
nor U2914 (N_2914,N_988,N_2406);
nand U2915 (N_2915,N_1203,N_664);
and U2916 (N_2916,N_672,N_630);
nand U2917 (N_2917,N_1284,N_432);
nand U2918 (N_2918,N_592,N_2189);
nor U2919 (N_2919,N_1532,N_1442);
nand U2920 (N_2920,N_1325,N_444);
and U2921 (N_2921,N_391,N_1146);
and U2922 (N_2922,N_1967,N_563);
and U2923 (N_2923,N_1792,N_535);
nor U2924 (N_2924,N_1471,N_467);
and U2925 (N_2925,N_1333,N_2385);
nor U2926 (N_2926,N_468,N_2396);
nor U2927 (N_2927,N_888,N_933);
and U2928 (N_2928,N_70,N_2473);
and U2929 (N_2929,N_652,N_2268);
and U2930 (N_2930,N_2007,N_2234);
nor U2931 (N_2931,N_15,N_783);
or U2932 (N_2932,N_2126,N_492);
or U2933 (N_2933,N_2090,N_1576);
and U2934 (N_2934,N_19,N_1577);
nor U2935 (N_2935,N_1190,N_863);
and U2936 (N_2936,N_2497,N_1455);
and U2937 (N_2937,N_181,N_1764);
and U2938 (N_2938,N_1988,N_252);
nor U2939 (N_2939,N_30,N_1226);
nand U2940 (N_2940,N_949,N_295);
xnor U2941 (N_2941,N_1813,N_1560);
and U2942 (N_2942,N_187,N_330);
nand U2943 (N_2943,N_2305,N_2426);
nor U2944 (N_2944,N_205,N_261);
and U2945 (N_2945,N_2082,N_1120);
nand U2946 (N_2946,N_42,N_50);
and U2947 (N_2947,N_1991,N_1425);
nand U2948 (N_2948,N_1419,N_2232);
nor U2949 (N_2949,N_2058,N_953);
nor U2950 (N_2950,N_26,N_338);
or U2951 (N_2951,N_191,N_88);
xnor U2952 (N_2952,N_44,N_510);
and U2953 (N_2953,N_1001,N_2);
nand U2954 (N_2954,N_1501,N_1682);
and U2955 (N_2955,N_1502,N_868);
nor U2956 (N_2956,N_1252,N_1189);
and U2957 (N_2957,N_924,N_2125);
and U2958 (N_2958,N_2159,N_1858);
and U2959 (N_2959,N_2351,N_760);
nor U2960 (N_2960,N_1312,N_1794);
nand U2961 (N_2961,N_679,N_448);
nor U2962 (N_2962,N_4,N_578);
nand U2963 (N_2963,N_844,N_109);
nand U2964 (N_2964,N_656,N_2357);
nand U2965 (N_2965,N_2236,N_349);
or U2966 (N_2966,N_201,N_2065);
xnor U2967 (N_2967,N_636,N_1705);
and U2968 (N_2968,N_1565,N_63);
or U2969 (N_2969,N_286,N_1610);
nor U2970 (N_2970,N_847,N_2258);
nor U2971 (N_2971,N_1919,N_2161);
nand U2972 (N_2972,N_595,N_2063);
nand U2973 (N_2973,N_2467,N_1178);
nand U2974 (N_2974,N_300,N_1127);
and U2975 (N_2975,N_1389,N_198);
nand U2976 (N_2976,N_966,N_2155);
or U2977 (N_2977,N_1054,N_2051);
and U2978 (N_2978,N_427,N_954);
nand U2979 (N_2979,N_741,N_2297);
xor U2980 (N_2980,N_474,N_920);
nand U2981 (N_2981,N_308,N_1833);
or U2982 (N_2982,N_1470,N_1646);
nand U2983 (N_2983,N_1918,N_660);
nor U2984 (N_2984,N_1007,N_234);
or U2985 (N_2985,N_1728,N_557);
or U2986 (N_2986,N_1184,N_178);
nor U2987 (N_2987,N_739,N_229);
and U2988 (N_2988,N_2227,N_2073);
and U2989 (N_2989,N_1787,N_842);
or U2990 (N_2990,N_152,N_1301);
and U2991 (N_2991,N_1593,N_1046);
and U2992 (N_2992,N_1796,N_973);
nand U2993 (N_2993,N_1966,N_325);
nor U2994 (N_2994,N_1192,N_1204);
xor U2995 (N_2995,N_2000,N_206);
or U2996 (N_2996,N_2484,N_1323);
and U2997 (N_2997,N_855,N_116);
xnor U2998 (N_2998,N_854,N_485);
and U2999 (N_2999,N_2148,N_1476);
and U3000 (N_3000,N_452,N_1826);
nor U3001 (N_3001,N_2301,N_1446);
nand U3002 (N_3002,N_1328,N_346);
nor U3003 (N_3003,N_1445,N_2443);
and U3004 (N_3004,N_1142,N_1983);
and U3005 (N_3005,N_1834,N_1903);
and U3006 (N_3006,N_1712,N_544);
or U3007 (N_3007,N_943,N_2309);
nand U3008 (N_3008,N_647,N_755);
xnor U3009 (N_3009,N_176,N_1895);
or U3010 (N_3010,N_1853,N_1840);
nand U3011 (N_3011,N_1103,N_894);
nor U3012 (N_3012,N_2466,N_1512);
nand U3013 (N_3013,N_1720,N_1361);
xor U3014 (N_3014,N_2118,N_431);
nand U3015 (N_3015,N_795,N_2012);
nand U3016 (N_3016,N_1238,N_907);
or U3017 (N_3017,N_857,N_1167);
or U3018 (N_3018,N_397,N_1812);
nand U3019 (N_3019,N_727,N_360);
xnor U3020 (N_3020,N_909,N_2299);
nand U3021 (N_3021,N_2068,N_1267);
xor U3022 (N_3022,N_873,N_1104);
and U3023 (N_3023,N_913,N_1902);
nor U3024 (N_3024,N_141,N_865);
and U3025 (N_3025,N_126,N_1490);
and U3026 (N_3026,N_669,N_1121);
nand U3027 (N_3027,N_1937,N_1412);
nand U3028 (N_3028,N_258,N_203);
nand U3029 (N_3029,N_984,N_2222);
nand U3030 (N_3030,N_1752,N_1924);
nand U3031 (N_3031,N_914,N_1657);
nand U3032 (N_3032,N_1486,N_1473);
xnor U3033 (N_3033,N_565,N_2403);
nor U3034 (N_3034,N_876,N_46);
nand U3035 (N_3035,N_2263,N_1612);
or U3036 (N_3036,N_1798,N_2138);
or U3037 (N_3037,N_1253,N_1246);
xor U3038 (N_3038,N_1286,N_51);
nor U3039 (N_3039,N_189,N_612);
and U3040 (N_3040,N_2066,N_1088);
and U3041 (N_3041,N_254,N_1148);
xnor U3042 (N_3042,N_1618,N_987);
nand U3043 (N_3043,N_1670,N_1677);
and U3044 (N_3044,N_1713,N_1943);
and U3045 (N_3045,N_1879,N_35);
or U3046 (N_3046,N_626,N_899);
nor U3047 (N_3047,N_610,N_101);
or U3048 (N_3048,N_457,N_478);
nand U3049 (N_3049,N_345,N_1686);
nor U3050 (N_3050,N_403,N_2176);
and U3051 (N_3051,N_766,N_2368);
and U3052 (N_3052,N_1993,N_1154);
nor U3053 (N_3053,N_2276,N_911);
or U3054 (N_3054,N_2432,N_607);
nand U3055 (N_3055,N_174,N_221);
nand U3056 (N_3056,N_2407,N_381);
nor U3057 (N_3057,N_1461,N_1538);
or U3058 (N_3058,N_2337,N_1733);
nand U3059 (N_3059,N_92,N_1427);
nand U3060 (N_3060,N_54,N_1974);
and U3061 (N_3061,N_2251,N_575);
nand U3062 (N_3062,N_414,N_1656);
nor U3063 (N_3063,N_846,N_773);
xor U3064 (N_3064,N_738,N_3);
xnor U3065 (N_3065,N_1413,N_1174);
nor U3066 (N_3066,N_644,N_317);
nor U3067 (N_3067,N_1725,N_439);
or U3068 (N_3068,N_549,N_2050);
nor U3069 (N_3069,N_2267,N_1241);
and U3070 (N_3070,N_522,N_1675);
nor U3071 (N_3071,N_469,N_1130);
and U3072 (N_3072,N_1280,N_1366);
nand U3073 (N_3073,N_175,N_396);
and U3074 (N_3074,N_292,N_306);
nand U3075 (N_3075,N_756,N_1339);
and U3076 (N_3076,N_1424,N_1016);
nand U3077 (N_3077,N_811,N_163);
and U3078 (N_3078,N_577,N_774);
nand U3079 (N_3079,N_1372,N_884);
xor U3080 (N_3080,N_287,N_2271);
nand U3081 (N_3081,N_1319,N_148);
nor U3082 (N_3082,N_147,N_207);
or U3083 (N_3083,N_1406,N_605);
xor U3084 (N_3084,N_1004,N_121);
and U3085 (N_3085,N_1365,N_585);
or U3086 (N_3086,N_561,N_1000);
nand U3087 (N_3087,N_1375,N_1183);
nor U3088 (N_3088,N_997,N_1508);
and U3089 (N_3089,N_2322,N_1536);
nand U3090 (N_3090,N_416,N_2255);
xor U3091 (N_3091,N_1335,N_433);
nor U3092 (N_3092,N_781,N_373);
nor U3093 (N_3093,N_1741,N_1136);
nand U3094 (N_3094,N_1854,N_1799);
xor U3095 (N_3095,N_2037,N_624);
nand U3096 (N_3096,N_1293,N_507);
or U3097 (N_3097,N_1309,N_704);
or U3098 (N_3098,N_225,N_291);
nand U3099 (N_3099,N_2071,N_456);
or U3100 (N_3100,N_2163,N_1589);
or U3101 (N_3101,N_231,N_1378);
nor U3102 (N_3102,N_1169,N_1243);
xnor U3103 (N_3103,N_801,N_6);
and U3104 (N_3104,N_459,N_689);
nor U3105 (N_3105,N_782,N_926);
xnor U3106 (N_3106,N_1417,N_1611);
xor U3107 (N_3107,N_570,N_707);
or U3108 (N_3108,N_757,N_532);
and U3109 (N_3109,N_1188,N_1888);
nand U3110 (N_3110,N_930,N_1185);
nor U3111 (N_3111,N_685,N_1970);
nor U3112 (N_3112,N_212,N_961);
nand U3113 (N_3113,N_665,N_2329);
or U3114 (N_3114,N_614,N_893);
and U3115 (N_3115,N_243,N_2278);
or U3116 (N_3116,N_108,N_388);
nor U3117 (N_3117,N_1545,N_974);
nand U3118 (N_3118,N_1209,N_538);
and U3119 (N_3119,N_1789,N_2334);
nor U3120 (N_3120,N_185,N_249);
and U3121 (N_3121,N_627,N_28);
or U3122 (N_3122,N_992,N_277);
or U3123 (N_3123,N_742,N_1116);
or U3124 (N_3124,N_420,N_253);
or U3125 (N_3125,N_9,N_719);
or U3126 (N_3126,N_1036,N_1897);
xor U3127 (N_3127,N_1381,N_778);
and U3128 (N_3128,N_681,N_481);
and U3129 (N_3129,N_1499,N_1714);
or U3130 (N_3130,N_1345,N_1064);
nand U3131 (N_3131,N_1595,N_870);
xor U3132 (N_3132,N_2316,N_621);
or U3133 (N_3133,N_385,N_743);
nand U3134 (N_3134,N_430,N_1549);
nor U3135 (N_3135,N_1695,N_197);
or U3136 (N_3136,N_1219,N_617);
and U3137 (N_3137,N_353,N_932);
nand U3138 (N_3138,N_1814,N_2338);
nand U3139 (N_3139,N_1648,N_2321);
xnor U3140 (N_3140,N_910,N_1329);
nor U3141 (N_3141,N_1070,N_2112);
and U3142 (N_3142,N_321,N_915);
xnor U3143 (N_3143,N_677,N_127);
xor U3144 (N_3144,N_1416,N_1062);
or U3145 (N_3145,N_1945,N_2355);
and U3146 (N_3146,N_419,N_2170);
and U3147 (N_3147,N_1696,N_2306);
or U3148 (N_3148,N_1052,N_1161);
nor U3149 (N_3149,N_2461,N_602);
and U3150 (N_3150,N_2233,N_2392);
nor U3151 (N_3151,N_498,N_2427);
or U3152 (N_3152,N_1601,N_329);
xnor U3153 (N_3153,N_1353,N_775);
and U3154 (N_3154,N_1938,N_2194);
xnor U3155 (N_3155,N_2045,N_2346);
xnor U3156 (N_3156,N_588,N_2029);
xnor U3157 (N_3157,N_2364,N_2318);
nor U3158 (N_3158,N_1268,N_1603);
and U3159 (N_3159,N_1514,N_415);
and U3160 (N_3160,N_2460,N_2445);
or U3161 (N_3161,N_1521,N_322);
or U3162 (N_3162,N_1180,N_1487);
nor U3163 (N_3163,N_2036,N_1382);
and U3164 (N_3164,N_785,N_654);
and U3165 (N_3165,N_951,N_1661);
nor U3166 (N_3166,N_1868,N_2345);
nor U3167 (N_3167,N_2288,N_2380);
and U3168 (N_3168,N_1031,N_1998);
nor U3169 (N_3169,N_581,N_2015);
xor U3170 (N_3170,N_1053,N_2462);
nor U3171 (N_3171,N_1084,N_1704);
nand U3172 (N_3172,N_722,N_1125);
nand U3173 (N_3173,N_849,N_1208);
xor U3174 (N_3174,N_2103,N_2412);
nand U3175 (N_3175,N_1410,N_1);
nor U3176 (N_3176,N_2454,N_786);
xnor U3177 (N_3177,N_1554,N_2464);
nand U3178 (N_3178,N_247,N_1266);
and U3179 (N_3179,N_1026,N_2213);
and U3180 (N_3180,N_2092,N_1398);
nand U3181 (N_3181,N_440,N_1197);
nor U3182 (N_3182,N_663,N_1214);
nor U3183 (N_3183,N_941,N_1608);
nor U3184 (N_3184,N_1066,N_1562);
nand U3185 (N_3185,N_798,N_516);
nand U3186 (N_3186,N_123,N_2095);
xor U3187 (N_3187,N_370,N_2203);
nand U3188 (N_3188,N_1228,N_323);
nand U3189 (N_3189,N_721,N_506);
nor U3190 (N_3190,N_833,N_1666);
and U3191 (N_3191,N_2001,N_1719);
nand U3192 (N_3192,N_1939,N_885);
and U3193 (N_3193,N_1662,N_1941);
nand U3194 (N_3194,N_731,N_43);
xnor U3195 (N_3195,N_1485,N_72);
and U3196 (N_3196,N_2485,N_2395);
xor U3197 (N_3197,N_272,N_2205);
nor U3198 (N_3198,N_850,N_1716);
or U3199 (N_3199,N_701,N_1811);
nand U3200 (N_3200,N_1922,N_566);
and U3201 (N_3201,N_1049,N_1960);
xnor U3202 (N_3202,N_642,N_68);
xnor U3203 (N_3203,N_2077,N_1457);
or U3204 (N_3204,N_1630,N_1761);
xnor U3205 (N_3205,N_2280,N_688);
nand U3206 (N_3206,N_1804,N_1772);
and U3207 (N_3207,N_1220,N_991);
nand U3208 (N_3208,N_450,N_819);
nor U3209 (N_3209,N_1702,N_714);
and U3210 (N_3210,N_380,N_1688);
nand U3211 (N_3211,N_2183,N_2319);
or U3212 (N_3212,N_1363,N_1181);
xor U3213 (N_3213,N_1845,N_1495);
nand U3214 (N_3214,N_255,N_1330);
nand U3215 (N_3215,N_1592,N_1014);
and U3216 (N_3216,N_328,N_1892);
nand U3217 (N_3217,N_74,N_957);
nand U3218 (N_3218,N_1564,N_2453);
nand U3219 (N_3219,N_2106,N_184);
nor U3220 (N_3220,N_1467,N_518);
nor U3221 (N_3221,N_183,N_1249);
or U3222 (N_3222,N_2179,N_1997);
and U3223 (N_3223,N_1684,N_1710);
or U3224 (N_3224,N_1045,N_604);
nand U3225 (N_3225,N_1882,N_1438);
nand U3226 (N_3226,N_2145,N_1647);
and U3227 (N_3227,N_134,N_2137);
xnor U3228 (N_3228,N_161,N_1342);
nand U3229 (N_3229,N_2116,N_171);
nand U3230 (N_3230,N_1449,N_2057);
and U3231 (N_3231,N_530,N_1762);
nand U3232 (N_3232,N_1660,N_2157);
and U3233 (N_3233,N_1354,N_1817);
or U3234 (N_3234,N_928,N_406);
or U3235 (N_3235,N_299,N_2104);
and U3236 (N_3236,N_1081,N_216);
or U3237 (N_3237,N_2067,N_143);
and U3238 (N_3238,N_2230,N_2379);
or U3239 (N_3239,N_1726,N_1822);
and U3240 (N_3240,N_931,N_2016);
nand U3241 (N_3241,N_382,N_2442);
nand U3242 (N_3242,N_1388,N_2496);
or U3243 (N_3243,N_2254,N_754);
or U3244 (N_3244,N_2098,N_673);
and U3245 (N_3245,N_872,N_708);
or U3246 (N_3246,N_1915,N_1222);
and U3247 (N_3247,N_720,N_342);
or U3248 (N_3248,N_1288,N_2146);
nor U3249 (N_3249,N_1432,N_1561);
nor U3250 (N_3250,N_1072,N_375);
or U3251 (N_3251,N_1391,N_1296);
or U3252 (N_3252,N_525,N_513);
nor U3253 (N_3253,N_787,N_2281);
nor U3254 (N_3254,N_228,N_2413);
nor U3255 (N_3255,N_1441,N_2275);
and U3256 (N_3256,N_158,N_211);
nand U3257 (N_3257,N_829,N_853);
and U3258 (N_3258,N_297,N_2450);
and U3259 (N_3259,N_1313,N_224);
or U3260 (N_3260,N_1150,N_2014);
nand U3261 (N_3261,N_1141,N_86);
or U3262 (N_3262,N_1022,N_554);
or U3263 (N_3263,N_511,N_1730);
nor U3264 (N_3264,N_374,N_1622);
or U3265 (N_3265,N_1914,N_1343);
nor U3266 (N_3266,N_1317,N_2231);
or U3267 (N_3267,N_1544,N_1881);
or U3268 (N_3268,N_2143,N_1489);
xor U3269 (N_3269,N_1371,N_540);
or U3270 (N_3270,N_2438,N_825);
and U3271 (N_3271,N_861,N_1963);
nor U3272 (N_3272,N_1758,N_2124);
xor U3273 (N_3273,N_55,N_1866);
or U3274 (N_3274,N_2131,N_1746);
nand U3275 (N_3275,N_75,N_2113);
or U3276 (N_3276,N_2072,N_1877);
or U3277 (N_3277,N_1886,N_622);
nor U3278 (N_3278,N_908,N_32);
nor U3279 (N_3279,N_1242,N_1308);
and U3280 (N_3280,N_1654,N_104);
xor U3281 (N_3281,N_1952,N_1118);
and U3282 (N_3282,N_2099,N_734);
xnor U3283 (N_3283,N_2429,N_589);
and U3284 (N_3284,N_1626,N_2044);
nor U3285 (N_3285,N_87,N_2431);
or U3286 (N_3286,N_268,N_813);
xnor U3287 (N_3287,N_62,N_1459);
nor U3288 (N_3288,N_2171,N_2195);
nand U3289 (N_3289,N_1803,N_1315);
nand U3290 (N_3290,N_429,N_1837);
nor U3291 (N_3291,N_2199,N_1076);
or U3292 (N_3292,N_1850,N_218);
or U3293 (N_3293,N_815,N_1480);
nand U3294 (N_3294,N_2415,N_1667);
nand U3295 (N_3295,N_2023,N_423);
nor U3296 (N_3296,N_2153,N_1260);
nand U3297 (N_3297,N_384,N_1836);
nand U3298 (N_3298,N_2291,N_753);
nand U3299 (N_3299,N_2369,N_2482);
or U3300 (N_3300,N_1211,N_1194);
nor U3301 (N_3301,N_702,N_1862);
or U3302 (N_3302,N_1976,N_890);
xor U3303 (N_3303,N_505,N_2165);
and U3304 (N_3304,N_1641,N_1019);
nand U3305 (N_3305,N_2056,N_1090);
nor U3306 (N_3306,N_436,N_41);
and U3307 (N_3307,N_1863,N_1479);
or U3308 (N_3308,N_976,N_699);
nand U3309 (N_3309,N_2274,N_156);
xnor U3310 (N_3310,N_1777,N_2402);
nand U3311 (N_3311,N_2087,N_820);
or U3312 (N_3312,N_1614,N_657);
or U3313 (N_3313,N_1408,N_2488);
xor U3314 (N_3314,N_1205,N_1290);
or U3315 (N_3315,N_2247,N_826);
nand U3316 (N_3316,N_2490,N_1754);
nand U3317 (N_3317,N_1182,N_378);
nand U3318 (N_3318,N_2193,N_1093);
and U3319 (N_3319,N_632,N_314);
nand U3320 (N_3320,N_371,N_1901);
nand U3321 (N_3321,N_392,N_2156);
or U3322 (N_3322,N_580,N_923);
nor U3323 (N_3323,N_1958,N_922);
and U3324 (N_3324,N_2494,N_1551);
and U3325 (N_3325,N_591,N_1123);
and U3326 (N_3326,N_376,N_2479);
and U3327 (N_3327,N_1114,N_623);
nand U3328 (N_3328,N_304,N_2085);
xnor U3329 (N_3329,N_1774,N_717);
or U3330 (N_3330,N_1852,N_2373);
and U3331 (N_3331,N_1240,N_168);
nor U3332 (N_3332,N_1607,N_1672);
and U3333 (N_3333,N_2486,N_2372);
xnor U3334 (N_3334,N_648,N_2172);
nand U3335 (N_3335,N_1386,N_2371);
or U3336 (N_3336,N_2206,N_713);
and U3337 (N_3337,N_460,N_125);
or U3338 (N_3338,N_2311,N_776);
or U3339 (N_3339,N_1172,N_1357);
and U3340 (N_3340,N_1916,N_1061);
nand U3341 (N_3341,N_1694,N_1928);
or U3342 (N_3342,N_745,N_1447);
nor U3343 (N_3343,N_1051,N_1609);
and U3344 (N_3344,N_629,N_1555);
nor U3345 (N_3345,N_1872,N_2377);
nor U3346 (N_3346,N_2376,N_1098);
nor U3347 (N_3347,N_1270,N_1492);
nor U3348 (N_3348,N_2260,N_960);
nand U3349 (N_3349,N_661,N_1571);
nor U3350 (N_3350,N_190,N_2272);
xor U3351 (N_3351,N_2349,N_1206);
and U3352 (N_3352,N_2204,N_649);
nor U3353 (N_3353,N_1771,N_1638);
and U3354 (N_3354,N_597,N_1524);
and U3355 (N_3355,N_2493,N_618);
and U3356 (N_3356,N_34,N_2340);
nand U3357 (N_3357,N_404,N_1113);
nor U3358 (N_3358,N_1526,N_1092);
and U3359 (N_3359,N_1823,N_2300);
nand U3360 (N_3360,N_2142,N_1953);
and U3361 (N_3361,N_1917,N_275);
nand U3362 (N_3362,N_2492,N_1405);
xnor U3363 (N_3363,N_834,N_1176);
nor U3364 (N_3364,N_409,N_1151);
nor U3365 (N_3365,N_1383,N_947);
nand U3366 (N_3366,N_779,N_969);
nand U3367 (N_3367,N_1078,N_1462);
nor U3368 (N_3368,N_919,N_730);
nand U3369 (N_3369,N_1334,N_466);
nor U3370 (N_3370,N_2167,N_1851);
nor U3371 (N_3371,N_537,N_1825);
nand U3372 (N_3372,N_1785,N_1699);
and U3373 (N_3373,N_285,N_1802);
nor U3374 (N_3374,N_1374,N_839);
nand U3375 (N_3375,N_1426,N_1056);
nand U3376 (N_3376,N_1128,N_723);
nor U3377 (N_3377,N_1627,N_1856);
nor U3378 (N_3378,N_2261,N_1466);
nor U3379 (N_3379,N_1784,N_2202);
nor U3380 (N_3380,N_886,N_1373);
nand U3381 (N_3381,N_1979,N_2018);
nand U3382 (N_3382,N_691,N_2130);
or U3383 (N_3383,N_1816,N_1750);
nor U3384 (N_3384,N_1579,N_1956);
nor U3385 (N_3385,N_2241,N_2214);
nor U3386 (N_3386,N_383,N_1755);
and U3387 (N_3387,N_1477,N_2100);
and U3388 (N_3388,N_770,N_365);
nand U3389 (N_3389,N_635,N_2358);
and U3390 (N_3390,N_1429,N_1865);
nand U3391 (N_3391,N_194,N_1331);
and U3392 (N_3392,N_2325,N_73);
nor U3393 (N_3393,N_2252,N_2080);
nor U3394 (N_3394,N_1507,N_1659);
nor U3395 (N_3395,N_902,N_1156);
nor U3396 (N_3396,N_83,N_1233);
nor U3397 (N_3397,N_1563,N_482);
nor U3398 (N_3398,N_940,N_2210);
nor U3399 (N_3399,N_337,N_316);
nor U3400 (N_3400,N_979,N_1844);
or U3401 (N_3401,N_2292,N_864);
and U3402 (N_3402,N_2336,N_413);
and U3403 (N_3403,N_114,N_2425);
nor U3404 (N_3404,N_263,N_1698);
nand U3405 (N_3405,N_455,N_13);
nor U3406 (N_3406,N_1393,N_2344);
nand U3407 (N_3407,N_2160,N_2004);
or U3408 (N_3408,N_1025,N_2290);
or U3409 (N_3409,N_233,N_1783);
xnor U3410 (N_3410,N_331,N_318);
nor U3411 (N_3411,N_2224,N_2481);
or U3412 (N_3412,N_687,N_2433);
and U3413 (N_3413,N_944,N_637);
and U3414 (N_3414,N_336,N_1443);
or U3415 (N_3415,N_400,N_188);
nor U3416 (N_3416,N_1717,N_85);
or U3417 (N_3417,N_1927,N_144);
and U3418 (N_3418,N_1655,N_659);
nand U3419 (N_3419,N_1978,N_896);
or U3420 (N_3420,N_541,N_1635);
or U3421 (N_3421,N_1808,N_1248);
or U3422 (N_3422,N_1981,N_897);
nor U3423 (N_3423,N_313,N_840);
nand U3424 (N_3424,N_1687,N_1770);
nand U3425 (N_3425,N_929,N_47);
xor U3426 (N_3426,N_1395,N_2447);
and U3427 (N_3427,N_118,N_1569);
nand U3428 (N_3428,N_289,N_94);
and U3429 (N_3429,N_352,N_1633);
xnor U3430 (N_3430,N_1855,N_788);
xor U3431 (N_3431,N_2339,N_1318);
nand U3432 (N_3432,N_2320,N_2002);
nor U3433 (N_3433,N_2262,N_643);
nor U3434 (N_3434,N_764,N_312);
or U3435 (N_3435,N_344,N_1665);
and U3436 (N_3436,N_2444,N_1996);
xor U3437 (N_3437,N_1539,N_1843);
and U3438 (N_3438,N_1012,N_298);
xnor U3439 (N_3439,N_150,N_1801);
nor U3440 (N_3440,N_2419,N_368);
nand U3441 (N_3441,N_2237,N_671);
nand U3442 (N_3442,N_1404,N_179);
or U3443 (N_3443,N_1452,N_1434);
nor U3444 (N_3444,N_1435,N_1896);
and U3445 (N_3445,N_641,N_2040);
and U3446 (N_3446,N_771,N_2164);
nor U3447 (N_3447,N_2162,N_2487);
and U3448 (N_3448,N_1460,N_2286);
and U3449 (N_3449,N_2383,N_1298);
and U3450 (N_3450,N_130,N_942);
xnor U3451 (N_3451,N_1397,N_562);
nor U3452 (N_3452,N_2209,N_1402);
or U3453 (N_3453,N_2180,N_1957);
xor U3454 (N_3454,N_350,N_2013);
nor U3455 (N_3455,N_1751,N_435);
nor U3456 (N_3456,N_520,N_1944);
or U3457 (N_3457,N_1759,N_856);
or U3458 (N_3458,N_1883,N_2151);
or U3459 (N_3459,N_2107,N_1880);
or U3460 (N_3460,N_1433,N_882);
nor U3461 (N_3461,N_494,N_2150);
nor U3462 (N_3462,N_2097,N_215);
or U3463 (N_3463,N_1100,N_1899);
or U3464 (N_3464,N_1024,N_1980);
or U3465 (N_3465,N_2483,N_1251);
nand U3466 (N_3466,N_2256,N_1454);
or U3467 (N_3467,N_1676,N_650);
or U3468 (N_3468,N_1059,N_22);
nor U3469 (N_3469,N_1110,N_569);
or U3470 (N_3470,N_1401,N_1171);
and U3471 (N_3471,N_962,N_1170);
nor U3472 (N_3472,N_1498,N_761);
nor U3473 (N_3473,N_523,N_1199);
nor U3474 (N_3474,N_751,N_2062);
xor U3475 (N_3475,N_1234,N_794);
or U3476 (N_3476,N_2144,N_405);
or U3477 (N_3477,N_1680,N_2181);
and U3478 (N_3478,N_1018,N_680);
nand U3479 (N_3479,N_69,N_438);
nand U3480 (N_3480,N_808,N_2471);
and U3481 (N_3481,N_1223,N_2249);
and U3482 (N_3482,N_96,N_495);
nand U3483 (N_3483,N_1658,N_759);
nand U3484 (N_3484,N_1302,N_1721);
and U3485 (N_3485,N_1387,N_559);
xor U3486 (N_3486,N_1265,N_534);
and U3487 (N_3487,N_1264,N_1278);
and U3488 (N_3488,N_1275,N_508);
and U3489 (N_3489,N_399,N_551);
nor U3490 (N_3490,N_1584,N_1060);
nand U3491 (N_3491,N_334,N_715);
nor U3492 (N_3492,N_2439,N_1422);
nand U3493 (N_3493,N_1775,N_38);
nor U3494 (N_3494,N_1894,N_2055);
and U3495 (N_3495,N_625,N_115);
and U3496 (N_3496,N_1962,N_1129);
and U3497 (N_3497,N_837,N_1027);
nor U3498 (N_3498,N_1598,N_2386);
xor U3499 (N_3499,N_1153,N_1594);
and U3500 (N_3500,N_693,N_1955);
and U3501 (N_3501,N_449,N_1083);
xnor U3502 (N_3502,N_2359,N_472);
and U3503 (N_3503,N_266,N_1828);
nor U3504 (N_3504,N_386,N_418);
or U3505 (N_3505,N_986,N_2075);
nand U3506 (N_3506,N_1094,N_1418);
xnor U3507 (N_3507,N_326,N_2411);
nor U3508 (N_3508,N_735,N_1122);
or U3509 (N_3509,N_501,N_80);
nor U3510 (N_3510,N_590,N_567);
or U3511 (N_3511,N_2389,N_1126);
nand U3512 (N_3512,N_830,N_2277);
or U3513 (N_3513,N_858,N_1585);
or U3514 (N_3514,N_2378,N_1835);
nor U3515 (N_3515,N_24,N_1106);
and U3516 (N_3516,N_1732,N_1653);
nand U3517 (N_3517,N_568,N_1352);
nand U3518 (N_3518,N_1087,N_79);
nand U3519 (N_3519,N_1847,N_791);
nand U3520 (N_3520,N_1272,N_1597);
or U3521 (N_3521,N_2188,N_904);
nand U3522 (N_3522,N_1017,N_1776);
nor U3523 (N_3523,N_1472,N_410);
or U3524 (N_3524,N_1706,N_269);
nand U3525 (N_3525,N_1769,N_1475);
xor U3526 (N_3526,N_1748,N_548);
and U3527 (N_3527,N_1320,N_246);
and U3528 (N_3528,N_129,N_10);
and U3529 (N_3529,N_259,N_477);
and U3530 (N_3530,N_2408,N_2424);
and U3531 (N_3531,N_1685,N_1580);
or U3532 (N_3532,N_1718,N_288);
nor U3533 (N_3533,N_1766,N_640);
or U3534 (N_3534,N_89,N_2088);
nor U3535 (N_3535,N_1269,N_628);
nor U3536 (N_3536,N_31,N_220);
or U3537 (N_3537,N_1742,N_1557);
and U3538 (N_3538,N_1738,N_2169);
xor U3539 (N_3539,N_60,N_609);
xnor U3540 (N_3540,N_1727,N_1541);
or U3541 (N_3541,N_2154,N_1305);
and U3542 (N_3542,N_1390,N_2114);
nand U3543 (N_3543,N_1119,N_1043);
nand U3544 (N_3544,N_1639,N_2003);
and U3545 (N_3545,N_0,N_964);
nor U3546 (N_3546,N_1572,N_1848);
nor U3547 (N_3547,N_1681,N_1994);
nor U3548 (N_3548,N_1152,N_1596);
xor U3549 (N_3549,N_690,N_2434);
nand U3550 (N_3550,N_638,N_111);
nor U3551 (N_3551,N_1930,N_2489);
nand U3552 (N_3552,N_1108,N_2054);
or U3553 (N_3553,N_195,N_193);
or U3554 (N_3554,N_1519,N_2242);
and U3555 (N_3555,N_2079,N_2259);
or U3556 (N_3556,N_1231,N_2225);
or U3557 (N_3557,N_1920,N_2129);
nor U3558 (N_3558,N_1407,N_906);
or U3559 (N_3559,N_273,N_2158);
nor U3560 (N_3560,N_1159,N_658);
nor U3561 (N_3561,N_1277,N_395);
nor U3562 (N_3562,N_802,N_1629);
and U3563 (N_3563,N_1456,N_2289);
nor U3564 (N_3564,N_1468,N_1790);
and U3565 (N_3565,N_1740,N_64);
or U3566 (N_3566,N_1518,N_1605);
nand U3567 (N_3567,N_2313,N_2323);
nand U3568 (N_3568,N_550,N_2480);
nand U3569 (N_3569,N_599,N_421);
and U3570 (N_3570,N_1907,N_2139);
nor U3571 (N_3571,N_45,N_1965);
nand U3572 (N_3572,N_340,N_1484);
or U3573 (N_3573,N_1394,N_2011);
nor U3574 (N_3574,N_1815,N_952);
or U3575 (N_3575,N_1950,N_2423);
nor U3576 (N_3576,N_196,N_1745);
and U3577 (N_3577,N_1743,N_1261);
or U3578 (N_3578,N_2046,N_2120);
xor U3579 (N_3579,N_700,N_186);
xnor U3580 (N_3580,N_2327,N_822);
or U3581 (N_3581,N_240,N_698);
xnor U3582 (N_3582,N_1198,N_310);
or U3583 (N_3583,N_1239,N_1041);
xnor U3584 (N_3584,N_1898,N_398);
or U3585 (N_3585,N_151,N_521);
and U3586 (N_3586,N_1258,N_172);
or U3587 (N_3587,N_862,N_393);
nor U3588 (N_3588,N_543,N_2186);
xor U3589 (N_3589,N_767,N_78);
xnor U3590 (N_3590,N_369,N_1047);
nand U3591 (N_3591,N_587,N_1516);
nand U3592 (N_3592,N_606,N_483);
or U3593 (N_3593,N_1744,N_2034);
xnor U3594 (N_3594,N_1162,N_1703);
or U3595 (N_3595,N_1368,N_1295);
nor U3596 (N_3596,N_762,N_97);
or U3597 (N_3597,N_560,N_1230);
and U3598 (N_3598,N_1326,N_2283);
or U3599 (N_3599,N_2363,N_192);
nor U3600 (N_3600,N_20,N_2282);
or U3601 (N_3601,N_2059,N_1364);
nand U3602 (N_3602,N_945,N_552);
or U3603 (N_3603,N_1165,N_1196);
or U3604 (N_3604,N_106,N_1008);
nand U3605 (N_3605,N_859,N_1020);
or U3606 (N_3606,N_2140,N_1926);
nor U3607 (N_3607,N_305,N_1338);
nand U3608 (N_3608,N_1414,N_959);
nand U3609 (N_3609,N_1690,N_1992);
nand U3610 (N_3610,N_927,N_1067);
nor U3611 (N_3611,N_594,N_1340);
nand U3612 (N_3612,N_912,N_666);
or U3613 (N_3613,N_900,N_512);
and U3614 (N_3614,N_2086,N_335);
or U3615 (N_3615,N_982,N_1450);
or U3616 (N_3616,N_2422,N_56);
and U3617 (N_3617,N_120,N_2078);
nor U3618 (N_3618,N_1581,N_777);
nand U3619 (N_3619,N_697,N_81);
or U3620 (N_3620,N_1503,N_1133);
and U3621 (N_3621,N_2030,N_1934);
nor U3622 (N_3622,N_99,N_281);
and U3623 (N_3623,N_803,N_2269);
and U3624 (N_3624,N_1619,N_1711);
or U3625 (N_3625,N_1210,N_2390);
nor U3626 (N_3626,N_1307,N_2033);
or U3627 (N_3627,N_2024,N_351);
nand U3628 (N_3628,N_1913,N_98);
and U3629 (N_3629,N_1057,N_2228);
nor U3630 (N_3630,N_1355,N_1488);
nor U3631 (N_3631,N_1615,N_1765);
and U3632 (N_3632,N_1984,N_2032);
nor U3633 (N_3633,N_2173,N_1570);
and U3634 (N_3634,N_2061,N_805);
nand U3635 (N_3635,N_17,N_879);
or U3636 (N_3636,N_2052,N_2076);
nand U3637 (N_3637,N_2333,N_2121);
or U3638 (N_3638,N_1299,N_1567);
or U3639 (N_3639,N_2478,N_119);
and U3640 (N_3640,N_1285,N_792);
or U3641 (N_3641,N_7,N_1535);
nor U3642 (N_3642,N_102,N_2265);
or U3643 (N_3643,N_1588,N_1095);
nand U3644 (N_3644,N_793,N_1643);
nand U3645 (N_3645,N_173,N_2141);
nor U3646 (N_3646,N_1289,N_1451);
nand U3647 (N_3647,N_1131,N_2174);
xor U3648 (N_3648,N_1809,N_2132);
and U3649 (N_3649,N_2133,N_2122);
nand U3650 (N_3650,N_500,N_2266);
and U3651 (N_3651,N_1079,N_1369);
nand U3652 (N_3652,N_2152,N_889);
xnor U3653 (N_3653,N_1453,N_937);
and U3654 (N_3654,N_1786,N_1954);
and U3655 (N_3655,N_2110,N_980);
nand U3656 (N_3656,N_1227,N_674);
nor U3657 (N_3657,N_93,N_1715);
and U3658 (N_3658,N_389,N_1911);
nor U3659 (N_3659,N_1015,N_601);
nor U3660 (N_3660,N_1349,N_2229);
and U3661 (N_3661,N_1158,N_2182);
or U3662 (N_3662,N_2410,N_712);
and U3663 (N_3663,N_1935,N_2147);
and U3664 (N_3664,N_956,N_1829);
nand U3665 (N_3665,N_2421,N_1867);
nor U3666 (N_3666,N_555,N_1237);
or U3667 (N_3667,N_2108,N_1827);
and U3668 (N_3668,N_1932,N_2360);
nor U3669 (N_3669,N_2476,N_1013);
nand U3670 (N_3670,N_1346,N_265);
nor U3671 (N_3671,N_2399,N_1846);
or U3672 (N_3672,N_918,N_1910);
and U3673 (N_3673,N_1005,N_2006);
nand U3674 (N_3674,N_2074,N_891);
nand U3675 (N_3675,N_90,N_412);
and U3676 (N_3676,N_812,N_718);
or U3677 (N_3677,N_2026,N_377);
nand U3678 (N_3678,N_1370,N_202);
and U3679 (N_3679,N_740,N_1912);
nor U3680 (N_3680,N_608,N_238);
nor U3681 (N_3681,N_1849,N_2038);
or U3682 (N_3682,N_1337,N_1032);
nor U3683 (N_3683,N_2394,N_1807);
and U3684 (N_3684,N_1244,N_2472);
nand U3685 (N_3685,N_1527,N_2342);
and U3686 (N_3686,N_810,N_1820);
or U3687 (N_3687,N_2135,N_724);
or U3688 (N_3688,N_264,N_364);
nor U3689 (N_3689,N_1085,N_746);
or U3690 (N_3690,N_23,N_860);
or U3691 (N_3691,N_769,N_1540);
or U3692 (N_3692,N_1155,N_1399);
nor U3693 (N_3693,N_1679,N_2367);
or U3694 (N_3694,N_1077,N_260);
or U3695 (N_3695,N_2495,N_166);
and U3696 (N_3696,N_2028,N_1558);
nor U3697 (N_3697,N_2091,N_2284);
and U3698 (N_3698,N_1649,N_1948);
nand U3699 (N_3699,N_1652,N_214);
and U3700 (N_3700,N_16,N_639);
and U3701 (N_3701,N_1513,N_1731);
nor U3702 (N_3702,N_749,N_145);
nand U3703 (N_3703,N_1351,N_480);
and U3704 (N_3704,N_2201,N_903);
nand U3705 (N_3705,N_916,N_733);
xor U3706 (N_3706,N_1871,N_573);
or U3707 (N_3707,N_1035,N_1356);
or U3708 (N_3708,N_1986,N_827);
nor U3709 (N_3709,N_1409,N_881);
and U3710 (N_3710,N_1411,N_1303);
or U3711 (N_3711,N_502,N_546);
nor U3712 (N_3712,N_105,N_294);
or U3713 (N_3713,N_2022,N_133);
nand U3714 (N_3714,N_2387,N_2084);
nand U3715 (N_3715,N_2117,N_1578);
nor U3716 (N_3716,N_1494,N_615);
nor U3717 (N_3717,N_1841,N_817);
nor U3718 (N_3718,N_2177,N_711);
nor U3719 (N_3719,N_1396,N_362);
or U3720 (N_3720,N_1806,N_159);
and U3721 (N_3721,N_584,N_257);
or U3722 (N_3722,N_1262,N_77);
or U3723 (N_3723,N_1530,N_995);
or U3724 (N_3724,N_1838,N_564);
and U3725 (N_3725,N_2248,N_2441);
nand U3726 (N_3726,N_1029,N_91);
nor U3727 (N_3727,N_866,N_499);
nand U3728 (N_3728,N_2257,N_848);
or U3729 (N_3729,N_2048,N_1218);
nand U3730 (N_3730,N_2060,N_235);
or U3731 (N_3731,N_1080,N_112);
nand U3732 (N_3732,N_57,N_2009);
nand U3733 (N_3733,N_363,N_1256);
nand U3734 (N_3734,N_2010,N_1874);
nand U3735 (N_3735,N_804,N_1891);
nand U3736 (N_3736,N_772,N_1099);
or U3737 (N_3737,N_1587,N_683);
or U3738 (N_3738,N_2175,N_1905);
nor U3739 (N_3739,N_1464,N_1055);
nor U3740 (N_3740,N_1215,N_1327);
nand U3741 (N_3741,N_668,N_162);
nor U3742 (N_3742,N_1533,N_169);
and U3743 (N_3743,N_695,N_1063);
or U3744 (N_3744,N_2134,N_1940);
nand U3745 (N_3745,N_1522,N_2375);
and U3746 (N_3746,N_1693,N_2384);
nor U3747 (N_3747,N_662,N_2226);
or U3748 (N_3748,N_271,N_222);
or U3749 (N_3749,N_1900,N_2115);
nand U3750 (N_3750,N_49,N_22);
or U3751 (N_3751,N_1155,N_349);
nor U3752 (N_3752,N_181,N_1516);
nor U3753 (N_3753,N_523,N_2092);
xor U3754 (N_3754,N_2031,N_174);
and U3755 (N_3755,N_1900,N_589);
xnor U3756 (N_3756,N_472,N_1832);
nand U3757 (N_3757,N_863,N_1105);
or U3758 (N_3758,N_2002,N_1740);
or U3759 (N_3759,N_827,N_1327);
or U3760 (N_3760,N_1949,N_637);
and U3761 (N_3761,N_1177,N_864);
nand U3762 (N_3762,N_1448,N_2272);
and U3763 (N_3763,N_1195,N_1478);
or U3764 (N_3764,N_281,N_1306);
or U3765 (N_3765,N_2301,N_605);
nor U3766 (N_3766,N_2475,N_342);
xor U3767 (N_3767,N_1112,N_824);
nor U3768 (N_3768,N_513,N_2333);
nor U3769 (N_3769,N_887,N_460);
nand U3770 (N_3770,N_776,N_1344);
nor U3771 (N_3771,N_1118,N_1154);
and U3772 (N_3772,N_535,N_1029);
and U3773 (N_3773,N_754,N_872);
nor U3774 (N_3774,N_1052,N_2358);
nand U3775 (N_3775,N_1800,N_472);
or U3776 (N_3776,N_2470,N_515);
nor U3777 (N_3777,N_1574,N_1817);
or U3778 (N_3778,N_2145,N_1204);
nor U3779 (N_3779,N_328,N_138);
nor U3780 (N_3780,N_14,N_936);
nor U3781 (N_3781,N_464,N_2239);
or U3782 (N_3782,N_2078,N_2194);
and U3783 (N_3783,N_1669,N_888);
nor U3784 (N_3784,N_36,N_1436);
or U3785 (N_3785,N_1033,N_1180);
nand U3786 (N_3786,N_768,N_1646);
nor U3787 (N_3787,N_240,N_323);
or U3788 (N_3788,N_1850,N_1101);
and U3789 (N_3789,N_2206,N_1450);
or U3790 (N_3790,N_1594,N_2307);
nor U3791 (N_3791,N_146,N_1282);
nor U3792 (N_3792,N_1595,N_1203);
and U3793 (N_3793,N_1311,N_557);
nor U3794 (N_3794,N_1664,N_180);
xnor U3795 (N_3795,N_1263,N_840);
or U3796 (N_3796,N_1297,N_1050);
nor U3797 (N_3797,N_1952,N_1209);
and U3798 (N_3798,N_2110,N_2335);
or U3799 (N_3799,N_292,N_1349);
and U3800 (N_3800,N_943,N_824);
or U3801 (N_3801,N_1307,N_937);
and U3802 (N_3802,N_1846,N_192);
xnor U3803 (N_3803,N_477,N_995);
nor U3804 (N_3804,N_538,N_699);
nor U3805 (N_3805,N_1995,N_1116);
nor U3806 (N_3806,N_20,N_2034);
nor U3807 (N_3807,N_1604,N_341);
nor U3808 (N_3808,N_2288,N_1002);
nand U3809 (N_3809,N_1465,N_1943);
and U3810 (N_3810,N_1762,N_2451);
xnor U3811 (N_3811,N_967,N_1487);
and U3812 (N_3812,N_1080,N_1446);
or U3813 (N_3813,N_1106,N_1424);
nor U3814 (N_3814,N_60,N_601);
or U3815 (N_3815,N_1050,N_2144);
nand U3816 (N_3816,N_1485,N_323);
nor U3817 (N_3817,N_1754,N_810);
xnor U3818 (N_3818,N_1267,N_123);
nand U3819 (N_3819,N_2156,N_1825);
xor U3820 (N_3820,N_2298,N_612);
and U3821 (N_3821,N_2411,N_152);
nand U3822 (N_3822,N_2074,N_2218);
nor U3823 (N_3823,N_816,N_1887);
nand U3824 (N_3824,N_129,N_1938);
nor U3825 (N_3825,N_673,N_2258);
and U3826 (N_3826,N_164,N_544);
or U3827 (N_3827,N_2065,N_509);
and U3828 (N_3828,N_2187,N_1614);
or U3829 (N_3829,N_473,N_102);
nand U3830 (N_3830,N_1242,N_1073);
and U3831 (N_3831,N_988,N_674);
nor U3832 (N_3832,N_1621,N_2265);
nand U3833 (N_3833,N_2063,N_1890);
or U3834 (N_3834,N_2174,N_682);
xor U3835 (N_3835,N_1586,N_944);
nor U3836 (N_3836,N_765,N_669);
nor U3837 (N_3837,N_1163,N_1629);
nor U3838 (N_3838,N_2243,N_2382);
and U3839 (N_3839,N_2261,N_393);
or U3840 (N_3840,N_1433,N_440);
and U3841 (N_3841,N_431,N_2180);
nand U3842 (N_3842,N_190,N_84);
xnor U3843 (N_3843,N_2074,N_606);
or U3844 (N_3844,N_2236,N_1559);
xnor U3845 (N_3845,N_1253,N_1922);
and U3846 (N_3846,N_2115,N_2128);
nor U3847 (N_3847,N_982,N_1254);
nand U3848 (N_3848,N_142,N_1305);
and U3849 (N_3849,N_1576,N_1456);
or U3850 (N_3850,N_851,N_768);
nand U3851 (N_3851,N_2071,N_2230);
and U3852 (N_3852,N_286,N_1333);
or U3853 (N_3853,N_1086,N_2171);
and U3854 (N_3854,N_1393,N_331);
nor U3855 (N_3855,N_695,N_143);
xor U3856 (N_3856,N_1692,N_23);
nand U3857 (N_3857,N_1515,N_1883);
and U3858 (N_3858,N_1705,N_1929);
and U3859 (N_3859,N_980,N_1254);
or U3860 (N_3860,N_1218,N_1760);
nor U3861 (N_3861,N_1534,N_1170);
and U3862 (N_3862,N_1345,N_2228);
nand U3863 (N_3863,N_405,N_1486);
nand U3864 (N_3864,N_1074,N_2328);
and U3865 (N_3865,N_228,N_2147);
and U3866 (N_3866,N_1475,N_1513);
nand U3867 (N_3867,N_1384,N_2194);
nor U3868 (N_3868,N_309,N_2121);
nand U3869 (N_3869,N_1024,N_1210);
and U3870 (N_3870,N_1249,N_1011);
or U3871 (N_3871,N_26,N_1432);
nor U3872 (N_3872,N_386,N_1804);
nand U3873 (N_3873,N_196,N_1785);
and U3874 (N_3874,N_1911,N_716);
and U3875 (N_3875,N_200,N_72);
and U3876 (N_3876,N_1466,N_1268);
or U3877 (N_3877,N_1833,N_2143);
nand U3878 (N_3878,N_1976,N_526);
xor U3879 (N_3879,N_2139,N_1097);
or U3880 (N_3880,N_984,N_1481);
nor U3881 (N_3881,N_1260,N_1174);
nand U3882 (N_3882,N_1536,N_1256);
nor U3883 (N_3883,N_1976,N_1708);
nand U3884 (N_3884,N_1420,N_2241);
and U3885 (N_3885,N_1675,N_1054);
xor U3886 (N_3886,N_642,N_1879);
xor U3887 (N_3887,N_1476,N_60);
nand U3888 (N_3888,N_2196,N_44);
nand U3889 (N_3889,N_1566,N_2404);
or U3890 (N_3890,N_1880,N_2139);
xor U3891 (N_3891,N_2187,N_1916);
and U3892 (N_3892,N_844,N_1689);
and U3893 (N_3893,N_2380,N_2111);
nor U3894 (N_3894,N_2030,N_1598);
xor U3895 (N_3895,N_800,N_2494);
or U3896 (N_3896,N_1368,N_2100);
nand U3897 (N_3897,N_2146,N_1172);
and U3898 (N_3898,N_537,N_1216);
nand U3899 (N_3899,N_299,N_2091);
and U3900 (N_3900,N_2266,N_1347);
nand U3901 (N_3901,N_382,N_1569);
and U3902 (N_3902,N_746,N_576);
nor U3903 (N_3903,N_171,N_1036);
nand U3904 (N_3904,N_1691,N_1866);
nand U3905 (N_3905,N_677,N_953);
nor U3906 (N_3906,N_1403,N_1182);
nor U3907 (N_3907,N_95,N_191);
and U3908 (N_3908,N_1706,N_589);
or U3909 (N_3909,N_434,N_146);
xor U3910 (N_3910,N_523,N_1010);
and U3911 (N_3911,N_822,N_1353);
or U3912 (N_3912,N_134,N_1587);
or U3913 (N_3913,N_36,N_70);
and U3914 (N_3914,N_1867,N_578);
and U3915 (N_3915,N_2215,N_17);
and U3916 (N_3916,N_619,N_711);
nor U3917 (N_3917,N_1265,N_1271);
and U3918 (N_3918,N_67,N_569);
xnor U3919 (N_3919,N_207,N_1354);
nor U3920 (N_3920,N_851,N_1199);
nand U3921 (N_3921,N_487,N_4);
nor U3922 (N_3922,N_981,N_1886);
and U3923 (N_3923,N_616,N_542);
xor U3924 (N_3924,N_2049,N_113);
or U3925 (N_3925,N_2231,N_21);
nor U3926 (N_3926,N_890,N_2111);
or U3927 (N_3927,N_1303,N_2249);
nand U3928 (N_3928,N_626,N_586);
xor U3929 (N_3929,N_1086,N_378);
xnor U3930 (N_3930,N_2289,N_2194);
and U3931 (N_3931,N_639,N_2252);
or U3932 (N_3932,N_1800,N_1564);
nor U3933 (N_3933,N_2076,N_2494);
and U3934 (N_3934,N_953,N_583);
or U3935 (N_3935,N_179,N_1051);
nor U3936 (N_3936,N_293,N_1163);
nand U3937 (N_3937,N_1879,N_27);
nor U3938 (N_3938,N_1701,N_1615);
and U3939 (N_3939,N_1899,N_1246);
or U3940 (N_3940,N_136,N_1895);
nor U3941 (N_3941,N_136,N_1605);
or U3942 (N_3942,N_2007,N_1837);
and U3943 (N_3943,N_55,N_586);
nor U3944 (N_3944,N_597,N_491);
or U3945 (N_3945,N_1550,N_1579);
and U3946 (N_3946,N_1690,N_1321);
and U3947 (N_3947,N_131,N_2467);
or U3948 (N_3948,N_465,N_1167);
and U3949 (N_3949,N_2321,N_2426);
nand U3950 (N_3950,N_577,N_908);
and U3951 (N_3951,N_1876,N_1625);
and U3952 (N_3952,N_2342,N_1311);
nand U3953 (N_3953,N_1603,N_2083);
nand U3954 (N_3954,N_1041,N_946);
nor U3955 (N_3955,N_236,N_938);
or U3956 (N_3956,N_2491,N_375);
nand U3957 (N_3957,N_2390,N_259);
and U3958 (N_3958,N_1157,N_369);
xor U3959 (N_3959,N_1930,N_929);
and U3960 (N_3960,N_1988,N_1642);
xor U3961 (N_3961,N_1304,N_554);
or U3962 (N_3962,N_1979,N_1691);
nand U3963 (N_3963,N_1801,N_2049);
and U3964 (N_3964,N_2226,N_679);
or U3965 (N_3965,N_304,N_19);
or U3966 (N_3966,N_2380,N_42);
nand U3967 (N_3967,N_1291,N_1678);
and U3968 (N_3968,N_1516,N_991);
or U3969 (N_3969,N_1451,N_674);
nor U3970 (N_3970,N_1118,N_2220);
nand U3971 (N_3971,N_924,N_548);
nand U3972 (N_3972,N_928,N_1367);
nor U3973 (N_3973,N_1140,N_919);
nand U3974 (N_3974,N_443,N_834);
nor U3975 (N_3975,N_1811,N_620);
or U3976 (N_3976,N_2057,N_2371);
or U3977 (N_3977,N_659,N_52);
nor U3978 (N_3978,N_1732,N_355);
nor U3979 (N_3979,N_2376,N_2228);
nand U3980 (N_3980,N_2214,N_2002);
and U3981 (N_3981,N_1648,N_395);
and U3982 (N_3982,N_294,N_2300);
and U3983 (N_3983,N_1987,N_530);
xor U3984 (N_3984,N_365,N_698);
or U3985 (N_3985,N_937,N_2275);
or U3986 (N_3986,N_1246,N_745);
nor U3987 (N_3987,N_1470,N_1503);
and U3988 (N_3988,N_159,N_1829);
nor U3989 (N_3989,N_1304,N_249);
nand U3990 (N_3990,N_1349,N_1061);
xnor U3991 (N_3991,N_1901,N_1889);
and U3992 (N_3992,N_2020,N_626);
or U3993 (N_3993,N_2206,N_272);
nand U3994 (N_3994,N_1028,N_2250);
nand U3995 (N_3995,N_400,N_907);
and U3996 (N_3996,N_125,N_741);
xor U3997 (N_3997,N_2414,N_1568);
nor U3998 (N_3998,N_2316,N_1202);
xor U3999 (N_3999,N_118,N_272);
or U4000 (N_4000,N_832,N_1779);
and U4001 (N_4001,N_1060,N_1887);
nand U4002 (N_4002,N_2083,N_1890);
xor U4003 (N_4003,N_1960,N_1780);
or U4004 (N_4004,N_2372,N_65);
and U4005 (N_4005,N_1660,N_366);
nor U4006 (N_4006,N_73,N_2126);
or U4007 (N_4007,N_2312,N_71);
xor U4008 (N_4008,N_1470,N_2422);
or U4009 (N_4009,N_829,N_46);
or U4010 (N_4010,N_522,N_568);
nand U4011 (N_4011,N_466,N_619);
or U4012 (N_4012,N_2068,N_415);
and U4013 (N_4013,N_429,N_1198);
xnor U4014 (N_4014,N_1849,N_801);
xor U4015 (N_4015,N_567,N_2488);
or U4016 (N_4016,N_1204,N_311);
nor U4017 (N_4017,N_389,N_1263);
nand U4018 (N_4018,N_446,N_721);
and U4019 (N_4019,N_1222,N_890);
nand U4020 (N_4020,N_1571,N_568);
nor U4021 (N_4021,N_2423,N_473);
nor U4022 (N_4022,N_2084,N_1723);
nor U4023 (N_4023,N_1386,N_2152);
nand U4024 (N_4024,N_75,N_1354);
or U4025 (N_4025,N_2032,N_2361);
or U4026 (N_4026,N_1012,N_1768);
and U4027 (N_4027,N_1665,N_972);
nor U4028 (N_4028,N_343,N_2416);
nor U4029 (N_4029,N_263,N_328);
or U4030 (N_4030,N_264,N_701);
nor U4031 (N_4031,N_388,N_347);
or U4032 (N_4032,N_1696,N_1191);
nor U4033 (N_4033,N_980,N_1499);
nor U4034 (N_4034,N_1242,N_104);
or U4035 (N_4035,N_2230,N_1631);
and U4036 (N_4036,N_1741,N_183);
or U4037 (N_4037,N_759,N_1170);
or U4038 (N_4038,N_2115,N_749);
and U4039 (N_4039,N_325,N_1351);
xor U4040 (N_4040,N_1438,N_1875);
and U4041 (N_4041,N_1826,N_2417);
and U4042 (N_4042,N_1546,N_1260);
and U4043 (N_4043,N_2148,N_1480);
or U4044 (N_4044,N_636,N_2273);
and U4045 (N_4045,N_1112,N_1223);
nor U4046 (N_4046,N_244,N_730);
nand U4047 (N_4047,N_2028,N_1536);
nor U4048 (N_4048,N_0,N_2388);
nor U4049 (N_4049,N_1942,N_1245);
nand U4050 (N_4050,N_322,N_2263);
and U4051 (N_4051,N_314,N_1361);
nor U4052 (N_4052,N_1807,N_2149);
nand U4053 (N_4053,N_1577,N_1325);
nor U4054 (N_4054,N_292,N_1364);
nand U4055 (N_4055,N_1666,N_1677);
nand U4056 (N_4056,N_26,N_853);
nand U4057 (N_4057,N_1283,N_2150);
xor U4058 (N_4058,N_568,N_900);
and U4059 (N_4059,N_508,N_1323);
xnor U4060 (N_4060,N_86,N_1158);
and U4061 (N_4061,N_1230,N_1074);
and U4062 (N_4062,N_2387,N_2167);
and U4063 (N_4063,N_1490,N_2052);
and U4064 (N_4064,N_1818,N_961);
and U4065 (N_4065,N_756,N_1294);
xnor U4066 (N_4066,N_2054,N_1304);
or U4067 (N_4067,N_1224,N_305);
and U4068 (N_4068,N_908,N_1996);
and U4069 (N_4069,N_1734,N_509);
or U4070 (N_4070,N_937,N_1266);
nand U4071 (N_4071,N_1179,N_1341);
nor U4072 (N_4072,N_2428,N_1875);
or U4073 (N_4073,N_587,N_143);
or U4074 (N_4074,N_2499,N_311);
or U4075 (N_4075,N_538,N_259);
nor U4076 (N_4076,N_1511,N_2472);
nor U4077 (N_4077,N_1831,N_792);
and U4078 (N_4078,N_832,N_1084);
and U4079 (N_4079,N_565,N_2085);
nand U4080 (N_4080,N_1237,N_1355);
nor U4081 (N_4081,N_737,N_1639);
and U4082 (N_4082,N_1362,N_1755);
xnor U4083 (N_4083,N_989,N_1728);
nand U4084 (N_4084,N_2467,N_1190);
xnor U4085 (N_4085,N_1931,N_7);
nand U4086 (N_4086,N_955,N_377);
nor U4087 (N_4087,N_620,N_877);
nor U4088 (N_4088,N_246,N_1197);
nand U4089 (N_4089,N_453,N_449);
or U4090 (N_4090,N_2063,N_1408);
nor U4091 (N_4091,N_1994,N_1659);
nand U4092 (N_4092,N_1090,N_574);
or U4093 (N_4093,N_298,N_1487);
or U4094 (N_4094,N_1988,N_1972);
nor U4095 (N_4095,N_1018,N_1829);
and U4096 (N_4096,N_346,N_1712);
and U4097 (N_4097,N_1327,N_394);
and U4098 (N_4098,N_408,N_880);
nand U4099 (N_4099,N_788,N_513);
xor U4100 (N_4100,N_1468,N_2372);
and U4101 (N_4101,N_168,N_1129);
nor U4102 (N_4102,N_2151,N_222);
nor U4103 (N_4103,N_810,N_1609);
nand U4104 (N_4104,N_503,N_1116);
nor U4105 (N_4105,N_597,N_1556);
or U4106 (N_4106,N_499,N_668);
nand U4107 (N_4107,N_259,N_33);
or U4108 (N_4108,N_2353,N_2345);
nor U4109 (N_4109,N_516,N_469);
xor U4110 (N_4110,N_2427,N_1526);
or U4111 (N_4111,N_613,N_844);
nor U4112 (N_4112,N_1886,N_1477);
nor U4113 (N_4113,N_1653,N_166);
nor U4114 (N_4114,N_1983,N_1823);
xnor U4115 (N_4115,N_1729,N_1350);
nand U4116 (N_4116,N_735,N_1745);
or U4117 (N_4117,N_1230,N_699);
nand U4118 (N_4118,N_713,N_1147);
nor U4119 (N_4119,N_1917,N_1881);
or U4120 (N_4120,N_207,N_1073);
and U4121 (N_4121,N_821,N_1956);
nand U4122 (N_4122,N_150,N_1469);
xnor U4123 (N_4123,N_2135,N_1574);
nand U4124 (N_4124,N_1906,N_2253);
nand U4125 (N_4125,N_356,N_1169);
or U4126 (N_4126,N_1327,N_1279);
and U4127 (N_4127,N_1136,N_370);
or U4128 (N_4128,N_959,N_2395);
or U4129 (N_4129,N_866,N_941);
and U4130 (N_4130,N_954,N_1053);
or U4131 (N_4131,N_1384,N_485);
and U4132 (N_4132,N_1714,N_136);
nor U4133 (N_4133,N_1543,N_1862);
nor U4134 (N_4134,N_2428,N_832);
and U4135 (N_4135,N_1660,N_1790);
nor U4136 (N_4136,N_366,N_2330);
xnor U4137 (N_4137,N_1349,N_813);
xnor U4138 (N_4138,N_1960,N_636);
and U4139 (N_4139,N_1104,N_2107);
nand U4140 (N_4140,N_2013,N_1457);
and U4141 (N_4141,N_1924,N_619);
nor U4142 (N_4142,N_839,N_674);
nor U4143 (N_4143,N_870,N_738);
or U4144 (N_4144,N_2126,N_976);
nor U4145 (N_4145,N_2374,N_1757);
nand U4146 (N_4146,N_111,N_1332);
nand U4147 (N_4147,N_1999,N_173);
nor U4148 (N_4148,N_326,N_694);
nor U4149 (N_4149,N_446,N_1014);
nand U4150 (N_4150,N_508,N_600);
nor U4151 (N_4151,N_1161,N_2387);
xnor U4152 (N_4152,N_641,N_1469);
xor U4153 (N_4153,N_549,N_268);
nor U4154 (N_4154,N_440,N_996);
and U4155 (N_4155,N_855,N_246);
and U4156 (N_4156,N_510,N_858);
nor U4157 (N_4157,N_1685,N_1868);
and U4158 (N_4158,N_78,N_242);
xor U4159 (N_4159,N_630,N_1559);
and U4160 (N_4160,N_2447,N_1634);
nand U4161 (N_4161,N_1527,N_325);
or U4162 (N_4162,N_1391,N_1266);
nor U4163 (N_4163,N_295,N_235);
nand U4164 (N_4164,N_2041,N_256);
or U4165 (N_4165,N_534,N_1678);
and U4166 (N_4166,N_161,N_1355);
or U4167 (N_4167,N_1390,N_1089);
and U4168 (N_4168,N_293,N_1881);
nor U4169 (N_4169,N_478,N_2283);
or U4170 (N_4170,N_2418,N_1739);
nand U4171 (N_4171,N_885,N_619);
or U4172 (N_4172,N_1540,N_599);
nand U4173 (N_4173,N_1949,N_866);
nand U4174 (N_4174,N_636,N_317);
or U4175 (N_4175,N_125,N_114);
and U4176 (N_4176,N_675,N_2250);
xor U4177 (N_4177,N_825,N_1714);
nor U4178 (N_4178,N_1564,N_400);
nand U4179 (N_4179,N_2311,N_675);
or U4180 (N_4180,N_80,N_1571);
and U4181 (N_4181,N_2457,N_1084);
and U4182 (N_4182,N_1265,N_2189);
nand U4183 (N_4183,N_1514,N_629);
and U4184 (N_4184,N_2130,N_2367);
and U4185 (N_4185,N_307,N_1327);
nand U4186 (N_4186,N_691,N_1241);
nand U4187 (N_4187,N_1615,N_330);
or U4188 (N_4188,N_1335,N_1784);
or U4189 (N_4189,N_1508,N_503);
and U4190 (N_4190,N_1521,N_1134);
and U4191 (N_4191,N_1702,N_2207);
nand U4192 (N_4192,N_1495,N_2489);
or U4193 (N_4193,N_633,N_1104);
or U4194 (N_4194,N_1993,N_1839);
and U4195 (N_4195,N_608,N_1675);
nand U4196 (N_4196,N_2281,N_1673);
nor U4197 (N_4197,N_968,N_1485);
or U4198 (N_4198,N_906,N_387);
nor U4199 (N_4199,N_1652,N_2183);
nand U4200 (N_4200,N_26,N_1335);
nand U4201 (N_4201,N_1187,N_1113);
and U4202 (N_4202,N_230,N_1300);
and U4203 (N_4203,N_1869,N_1237);
or U4204 (N_4204,N_960,N_2262);
xnor U4205 (N_4205,N_568,N_204);
or U4206 (N_4206,N_2257,N_915);
and U4207 (N_4207,N_2163,N_2337);
and U4208 (N_4208,N_2076,N_344);
and U4209 (N_4209,N_832,N_690);
nor U4210 (N_4210,N_1252,N_536);
nor U4211 (N_4211,N_2020,N_981);
nor U4212 (N_4212,N_523,N_1761);
nor U4213 (N_4213,N_154,N_2372);
and U4214 (N_4214,N_2003,N_1600);
nand U4215 (N_4215,N_528,N_2223);
or U4216 (N_4216,N_1447,N_766);
and U4217 (N_4217,N_130,N_820);
and U4218 (N_4218,N_1521,N_1669);
nor U4219 (N_4219,N_1008,N_340);
nand U4220 (N_4220,N_2469,N_717);
nor U4221 (N_4221,N_2021,N_202);
nor U4222 (N_4222,N_436,N_2276);
xnor U4223 (N_4223,N_1869,N_208);
xnor U4224 (N_4224,N_2214,N_2398);
xor U4225 (N_4225,N_2198,N_948);
nand U4226 (N_4226,N_1907,N_1718);
or U4227 (N_4227,N_763,N_1934);
nand U4228 (N_4228,N_1529,N_1855);
nor U4229 (N_4229,N_1222,N_407);
nor U4230 (N_4230,N_1337,N_342);
or U4231 (N_4231,N_1956,N_1752);
and U4232 (N_4232,N_1351,N_327);
or U4233 (N_4233,N_1079,N_1651);
or U4234 (N_4234,N_410,N_51);
or U4235 (N_4235,N_2173,N_1473);
nand U4236 (N_4236,N_1135,N_326);
nor U4237 (N_4237,N_1429,N_2163);
and U4238 (N_4238,N_1765,N_1762);
nor U4239 (N_4239,N_2266,N_1152);
or U4240 (N_4240,N_1963,N_1438);
xor U4241 (N_4241,N_2309,N_940);
nand U4242 (N_4242,N_1904,N_1732);
xor U4243 (N_4243,N_1070,N_830);
and U4244 (N_4244,N_1275,N_65);
xnor U4245 (N_4245,N_806,N_575);
nand U4246 (N_4246,N_1688,N_2340);
or U4247 (N_4247,N_1211,N_1465);
or U4248 (N_4248,N_1177,N_113);
nor U4249 (N_4249,N_717,N_281);
and U4250 (N_4250,N_1225,N_230);
xnor U4251 (N_4251,N_315,N_970);
xor U4252 (N_4252,N_1806,N_1555);
or U4253 (N_4253,N_1410,N_491);
and U4254 (N_4254,N_1275,N_273);
xor U4255 (N_4255,N_2151,N_1387);
nor U4256 (N_4256,N_408,N_302);
nand U4257 (N_4257,N_949,N_1454);
nand U4258 (N_4258,N_1524,N_459);
xor U4259 (N_4259,N_23,N_423);
xor U4260 (N_4260,N_344,N_1729);
or U4261 (N_4261,N_2488,N_100);
nor U4262 (N_4262,N_871,N_461);
and U4263 (N_4263,N_1132,N_2);
and U4264 (N_4264,N_505,N_814);
and U4265 (N_4265,N_181,N_1560);
and U4266 (N_4266,N_220,N_2155);
nor U4267 (N_4267,N_600,N_1318);
nor U4268 (N_4268,N_151,N_2002);
or U4269 (N_4269,N_2450,N_516);
or U4270 (N_4270,N_1280,N_243);
nor U4271 (N_4271,N_1384,N_513);
and U4272 (N_4272,N_2311,N_1659);
nor U4273 (N_4273,N_1512,N_592);
nand U4274 (N_4274,N_1392,N_2139);
or U4275 (N_4275,N_2187,N_724);
and U4276 (N_4276,N_499,N_823);
nand U4277 (N_4277,N_2160,N_77);
nand U4278 (N_4278,N_911,N_1750);
or U4279 (N_4279,N_1408,N_1997);
xnor U4280 (N_4280,N_2040,N_2339);
nor U4281 (N_4281,N_566,N_2114);
and U4282 (N_4282,N_1765,N_2110);
nor U4283 (N_4283,N_414,N_34);
nor U4284 (N_4284,N_1658,N_2476);
and U4285 (N_4285,N_1922,N_1385);
nand U4286 (N_4286,N_1719,N_178);
and U4287 (N_4287,N_1607,N_2353);
or U4288 (N_4288,N_2083,N_933);
or U4289 (N_4289,N_2047,N_1984);
and U4290 (N_4290,N_254,N_255);
and U4291 (N_4291,N_1735,N_480);
xnor U4292 (N_4292,N_75,N_897);
and U4293 (N_4293,N_707,N_1675);
nor U4294 (N_4294,N_213,N_685);
and U4295 (N_4295,N_2156,N_805);
nor U4296 (N_4296,N_1937,N_1875);
xor U4297 (N_4297,N_1026,N_2066);
nand U4298 (N_4298,N_2155,N_309);
nor U4299 (N_4299,N_30,N_2373);
or U4300 (N_4300,N_476,N_263);
or U4301 (N_4301,N_1,N_1352);
nand U4302 (N_4302,N_207,N_321);
xnor U4303 (N_4303,N_113,N_1745);
or U4304 (N_4304,N_435,N_1341);
or U4305 (N_4305,N_1781,N_1441);
xnor U4306 (N_4306,N_2142,N_867);
nor U4307 (N_4307,N_2090,N_313);
or U4308 (N_4308,N_722,N_1328);
nor U4309 (N_4309,N_1783,N_1797);
and U4310 (N_4310,N_1608,N_633);
nor U4311 (N_4311,N_1310,N_1996);
nand U4312 (N_4312,N_2368,N_2212);
nor U4313 (N_4313,N_1763,N_1777);
nand U4314 (N_4314,N_871,N_630);
nor U4315 (N_4315,N_908,N_281);
nand U4316 (N_4316,N_765,N_2275);
and U4317 (N_4317,N_551,N_1270);
or U4318 (N_4318,N_1090,N_46);
nand U4319 (N_4319,N_1298,N_658);
nor U4320 (N_4320,N_2415,N_756);
and U4321 (N_4321,N_1977,N_1288);
and U4322 (N_4322,N_64,N_367);
and U4323 (N_4323,N_344,N_1447);
or U4324 (N_4324,N_674,N_1487);
or U4325 (N_4325,N_1178,N_2343);
or U4326 (N_4326,N_2135,N_1265);
and U4327 (N_4327,N_1476,N_1732);
xnor U4328 (N_4328,N_2233,N_1542);
and U4329 (N_4329,N_72,N_777);
nand U4330 (N_4330,N_1306,N_1854);
and U4331 (N_4331,N_868,N_1692);
nor U4332 (N_4332,N_1247,N_1657);
and U4333 (N_4333,N_3,N_1178);
nand U4334 (N_4334,N_1115,N_2141);
or U4335 (N_4335,N_393,N_457);
and U4336 (N_4336,N_773,N_2179);
and U4337 (N_4337,N_1987,N_1282);
nor U4338 (N_4338,N_2313,N_617);
or U4339 (N_4339,N_2333,N_2070);
nor U4340 (N_4340,N_968,N_1114);
nor U4341 (N_4341,N_688,N_2239);
nand U4342 (N_4342,N_1368,N_332);
nand U4343 (N_4343,N_1301,N_1287);
nand U4344 (N_4344,N_1053,N_1936);
nor U4345 (N_4345,N_1241,N_93);
xor U4346 (N_4346,N_928,N_633);
and U4347 (N_4347,N_1376,N_2171);
nor U4348 (N_4348,N_1696,N_1357);
or U4349 (N_4349,N_1119,N_2320);
nor U4350 (N_4350,N_1877,N_1074);
xnor U4351 (N_4351,N_1790,N_2042);
and U4352 (N_4352,N_1963,N_330);
nand U4353 (N_4353,N_1036,N_1851);
nand U4354 (N_4354,N_2370,N_39);
nor U4355 (N_4355,N_1170,N_561);
nor U4356 (N_4356,N_835,N_171);
xnor U4357 (N_4357,N_1658,N_1796);
nor U4358 (N_4358,N_1006,N_26);
xor U4359 (N_4359,N_708,N_1953);
or U4360 (N_4360,N_1743,N_945);
or U4361 (N_4361,N_1598,N_2337);
nor U4362 (N_4362,N_179,N_899);
nor U4363 (N_4363,N_457,N_339);
and U4364 (N_4364,N_976,N_850);
nor U4365 (N_4365,N_1879,N_28);
nor U4366 (N_4366,N_1978,N_2356);
nand U4367 (N_4367,N_1257,N_2227);
nand U4368 (N_4368,N_1640,N_2315);
and U4369 (N_4369,N_44,N_1864);
nor U4370 (N_4370,N_1896,N_794);
or U4371 (N_4371,N_1414,N_1656);
nand U4372 (N_4372,N_2060,N_1977);
nor U4373 (N_4373,N_1167,N_204);
nor U4374 (N_4374,N_709,N_2027);
nand U4375 (N_4375,N_19,N_1199);
nand U4376 (N_4376,N_2210,N_1684);
nand U4377 (N_4377,N_2339,N_1612);
nand U4378 (N_4378,N_1674,N_2213);
and U4379 (N_4379,N_1882,N_2381);
or U4380 (N_4380,N_1331,N_738);
and U4381 (N_4381,N_2459,N_2335);
nand U4382 (N_4382,N_1731,N_1225);
xnor U4383 (N_4383,N_2038,N_917);
and U4384 (N_4384,N_71,N_327);
xnor U4385 (N_4385,N_570,N_341);
nor U4386 (N_4386,N_2388,N_1652);
nand U4387 (N_4387,N_327,N_2212);
or U4388 (N_4388,N_576,N_646);
and U4389 (N_4389,N_1800,N_883);
xor U4390 (N_4390,N_233,N_927);
nor U4391 (N_4391,N_37,N_902);
nor U4392 (N_4392,N_988,N_926);
nand U4393 (N_4393,N_59,N_1423);
nand U4394 (N_4394,N_2334,N_1033);
nor U4395 (N_4395,N_2134,N_1722);
nand U4396 (N_4396,N_2325,N_1999);
nor U4397 (N_4397,N_1529,N_1624);
nand U4398 (N_4398,N_2021,N_1047);
nand U4399 (N_4399,N_1146,N_2088);
nand U4400 (N_4400,N_685,N_1517);
nand U4401 (N_4401,N_313,N_2468);
xnor U4402 (N_4402,N_2234,N_953);
nand U4403 (N_4403,N_1526,N_2423);
or U4404 (N_4404,N_1901,N_1486);
nand U4405 (N_4405,N_874,N_975);
or U4406 (N_4406,N_2410,N_1754);
xor U4407 (N_4407,N_2327,N_2177);
nand U4408 (N_4408,N_0,N_916);
or U4409 (N_4409,N_2026,N_2435);
and U4410 (N_4410,N_670,N_535);
nand U4411 (N_4411,N_726,N_339);
nand U4412 (N_4412,N_1998,N_2413);
nand U4413 (N_4413,N_675,N_850);
nand U4414 (N_4414,N_1335,N_640);
and U4415 (N_4415,N_2379,N_721);
and U4416 (N_4416,N_595,N_1325);
and U4417 (N_4417,N_1343,N_2243);
and U4418 (N_4418,N_1794,N_1287);
nor U4419 (N_4419,N_944,N_471);
nand U4420 (N_4420,N_618,N_1327);
or U4421 (N_4421,N_555,N_1031);
or U4422 (N_4422,N_413,N_1462);
or U4423 (N_4423,N_1569,N_1383);
nand U4424 (N_4424,N_970,N_1123);
nand U4425 (N_4425,N_1946,N_2292);
nor U4426 (N_4426,N_35,N_85);
nor U4427 (N_4427,N_334,N_1739);
and U4428 (N_4428,N_2495,N_356);
or U4429 (N_4429,N_2188,N_481);
and U4430 (N_4430,N_1560,N_688);
xor U4431 (N_4431,N_240,N_951);
nor U4432 (N_4432,N_1788,N_2066);
xor U4433 (N_4433,N_524,N_710);
nand U4434 (N_4434,N_2271,N_850);
and U4435 (N_4435,N_900,N_2051);
nor U4436 (N_4436,N_311,N_2118);
nand U4437 (N_4437,N_2267,N_719);
nand U4438 (N_4438,N_1857,N_1223);
and U4439 (N_4439,N_1458,N_320);
or U4440 (N_4440,N_2132,N_1987);
and U4441 (N_4441,N_658,N_303);
or U4442 (N_4442,N_745,N_1295);
and U4443 (N_4443,N_1628,N_509);
and U4444 (N_4444,N_2337,N_1045);
nand U4445 (N_4445,N_862,N_2299);
and U4446 (N_4446,N_584,N_1433);
and U4447 (N_4447,N_374,N_1388);
nand U4448 (N_4448,N_2446,N_1016);
nor U4449 (N_4449,N_1004,N_2259);
or U4450 (N_4450,N_1614,N_612);
and U4451 (N_4451,N_2063,N_805);
nand U4452 (N_4452,N_515,N_1870);
nor U4453 (N_4453,N_2024,N_860);
nand U4454 (N_4454,N_2043,N_981);
nor U4455 (N_4455,N_1808,N_312);
or U4456 (N_4456,N_798,N_2387);
nor U4457 (N_4457,N_1674,N_875);
nor U4458 (N_4458,N_1744,N_1456);
xnor U4459 (N_4459,N_1798,N_1575);
and U4460 (N_4460,N_1927,N_1626);
or U4461 (N_4461,N_596,N_2456);
nand U4462 (N_4462,N_1280,N_1075);
nand U4463 (N_4463,N_1301,N_8);
nand U4464 (N_4464,N_891,N_1064);
or U4465 (N_4465,N_119,N_2466);
nand U4466 (N_4466,N_1319,N_1779);
nor U4467 (N_4467,N_1198,N_2294);
nand U4468 (N_4468,N_2309,N_1455);
or U4469 (N_4469,N_1067,N_1230);
nand U4470 (N_4470,N_1841,N_1733);
nand U4471 (N_4471,N_1928,N_1005);
nor U4472 (N_4472,N_304,N_532);
or U4473 (N_4473,N_48,N_1663);
or U4474 (N_4474,N_1184,N_131);
nand U4475 (N_4475,N_355,N_1117);
nand U4476 (N_4476,N_815,N_1138);
or U4477 (N_4477,N_1088,N_438);
nand U4478 (N_4478,N_293,N_1936);
or U4479 (N_4479,N_1763,N_1734);
nand U4480 (N_4480,N_0,N_635);
or U4481 (N_4481,N_28,N_1616);
nor U4482 (N_4482,N_44,N_2470);
and U4483 (N_4483,N_2412,N_2192);
and U4484 (N_4484,N_1275,N_1418);
nand U4485 (N_4485,N_944,N_6);
and U4486 (N_4486,N_1993,N_654);
or U4487 (N_4487,N_898,N_1648);
and U4488 (N_4488,N_875,N_565);
nand U4489 (N_4489,N_1979,N_917);
or U4490 (N_4490,N_1496,N_849);
nor U4491 (N_4491,N_2014,N_232);
or U4492 (N_4492,N_1864,N_1775);
nor U4493 (N_4493,N_493,N_448);
and U4494 (N_4494,N_1375,N_1134);
or U4495 (N_4495,N_479,N_145);
nand U4496 (N_4496,N_604,N_760);
nor U4497 (N_4497,N_50,N_1509);
nand U4498 (N_4498,N_1030,N_1077);
or U4499 (N_4499,N_1769,N_1101);
nand U4500 (N_4500,N_908,N_1861);
and U4501 (N_4501,N_1238,N_835);
nand U4502 (N_4502,N_1445,N_1942);
nor U4503 (N_4503,N_317,N_884);
nor U4504 (N_4504,N_100,N_1102);
xnor U4505 (N_4505,N_20,N_3);
nor U4506 (N_4506,N_127,N_2115);
or U4507 (N_4507,N_610,N_820);
or U4508 (N_4508,N_427,N_1807);
nor U4509 (N_4509,N_205,N_560);
and U4510 (N_4510,N_2000,N_1890);
xor U4511 (N_4511,N_520,N_819);
nor U4512 (N_4512,N_486,N_947);
nand U4513 (N_4513,N_1261,N_271);
and U4514 (N_4514,N_2128,N_244);
nor U4515 (N_4515,N_1978,N_1898);
and U4516 (N_4516,N_598,N_1141);
xnor U4517 (N_4517,N_156,N_514);
nor U4518 (N_4518,N_1449,N_591);
nand U4519 (N_4519,N_28,N_1742);
and U4520 (N_4520,N_325,N_2461);
nor U4521 (N_4521,N_1031,N_218);
nand U4522 (N_4522,N_984,N_181);
nand U4523 (N_4523,N_1680,N_1608);
xor U4524 (N_4524,N_319,N_1462);
nand U4525 (N_4525,N_1731,N_1523);
or U4526 (N_4526,N_1066,N_93);
nand U4527 (N_4527,N_163,N_232);
and U4528 (N_4528,N_561,N_1798);
nor U4529 (N_4529,N_105,N_1023);
nor U4530 (N_4530,N_172,N_655);
nand U4531 (N_4531,N_1350,N_1296);
nor U4532 (N_4532,N_2079,N_1585);
and U4533 (N_4533,N_1579,N_1916);
or U4534 (N_4534,N_1163,N_236);
xnor U4535 (N_4535,N_636,N_1117);
xor U4536 (N_4536,N_1656,N_2281);
and U4537 (N_4537,N_315,N_142);
nor U4538 (N_4538,N_1687,N_2306);
or U4539 (N_4539,N_1605,N_2472);
or U4540 (N_4540,N_543,N_855);
and U4541 (N_4541,N_1233,N_193);
nor U4542 (N_4542,N_1214,N_1549);
nor U4543 (N_4543,N_600,N_1585);
nor U4544 (N_4544,N_2353,N_1494);
nand U4545 (N_4545,N_427,N_1333);
xor U4546 (N_4546,N_2359,N_1463);
nand U4547 (N_4547,N_2065,N_2244);
or U4548 (N_4548,N_1555,N_81);
or U4549 (N_4549,N_1621,N_59);
or U4550 (N_4550,N_1349,N_2347);
or U4551 (N_4551,N_2485,N_1396);
nor U4552 (N_4552,N_1071,N_496);
or U4553 (N_4553,N_1962,N_1261);
nand U4554 (N_4554,N_2134,N_503);
nor U4555 (N_4555,N_1791,N_2026);
nor U4556 (N_4556,N_745,N_2020);
nor U4557 (N_4557,N_1864,N_113);
nand U4558 (N_4558,N_2017,N_1900);
nand U4559 (N_4559,N_540,N_929);
nand U4560 (N_4560,N_985,N_2299);
nand U4561 (N_4561,N_1839,N_1291);
or U4562 (N_4562,N_234,N_1995);
nand U4563 (N_4563,N_1926,N_1715);
xor U4564 (N_4564,N_148,N_1472);
and U4565 (N_4565,N_1545,N_1379);
nor U4566 (N_4566,N_1057,N_465);
or U4567 (N_4567,N_33,N_1476);
or U4568 (N_4568,N_1803,N_137);
or U4569 (N_4569,N_1557,N_2451);
nor U4570 (N_4570,N_1258,N_1946);
and U4571 (N_4571,N_270,N_1133);
nor U4572 (N_4572,N_1212,N_1745);
nor U4573 (N_4573,N_462,N_2149);
xnor U4574 (N_4574,N_2259,N_2082);
and U4575 (N_4575,N_1998,N_220);
xnor U4576 (N_4576,N_2068,N_1701);
nand U4577 (N_4577,N_429,N_2415);
or U4578 (N_4578,N_1280,N_2265);
or U4579 (N_4579,N_2134,N_760);
nand U4580 (N_4580,N_857,N_480);
nand U4581 (N_4581,N_1715,N_333);
and U4582 (N_4582,N_317,N_1979);
nand U4583 (N_4583,N_2441,N_2149);
and U4584 (N_4584,N_85,N_1939);
or U4585 (N_4585,N_157,N_1045);
or U4586 (N_4586,N_397,N_2129);
and U4587 (N_4587,N_1106,N_1540);
or U4588 (N_4588,N_2249,N_507);
nand U4589 (N_4589,N_659,N_1709);
nand U4590 (N_4590,N_2202,N_2325);
or U4591 (N_4591,N_837,N_1642);
or U4592 (N_4592,N_195,N_1782);
or U4593 (N_4593,N_891,N_1022);
nor U4594 (N_4594,N_2184,N_846);
nand U4595 (N_4595,N_84,N_2035);
nand U4596 (N_4596,N_459,N_802);
xnor U4597 (N_4597,N_1371,N_692);
nand U4598 (N_4598,N_1050,N_1335);
or U4599 (N_4599,N_366,N_1061);
nand U4600 (N_4600,N_2088,N_805);
and U4601 (N_4601,N_1541,N_163);
nor U4602 (N_4602,N_2297,N_1134);
nor U4603 (N_4603,N_2102,N_962);
or U4604 (N_4604,N_2288,N_603);
nand U4605 (N_4605,N_464,N_970);
nand U4606 (N_4606,N_239,N_238);
or U4607 (N_4607,N_2288,N_1535);
nand U4608 (N_4608,N_1859,N_139);
nand U4609 (N_4609,N_1758,N_328);
xor U4610 (N_4610,N_1122,N_1964);
and U4611 (N_4611,N_1660,N_1320);
or U4612 (N_4612,N_1998,N_350);
or U4613 (N_4613,N_1862,N_760);
xnor U4614 (N_4614,N_279,N_788);
xor U4615 (N_4615,N_976,N_1231);
and U4616 (N_4616,N_449,N_961);
nand U4617 (N_4617,N_2480,N_1444);
or U4618 (N_4618,N_439,N_1961);
or U4619 (N_4619,N_571,N_1710);
nand U4620 (N_4620,N_198,N_1142);
nor U4621 (N_4621,N_545,N_1039);
nor U4622 (N_4622,N_2041,N_1296);
nor U4623 (N_4623,N_708,N_187);
nand U4624 (N_4624,N_24,N_1190);
or U4625 (N_4625,N_1402,N_1790);
xor U4626 (N_4626,N_1831,N_745);
nand U4627 (N_4627,N_301,N_1962);
or U4628 (N_4628,N_491,N_2320);
nor U4629 (N_4629,N_519,N_2436);
nor U4630 (N_4630,N_973,N_1232);
nand U4631 (N_4631,N_1397,N_368);
and U4632 (N_4632,N_1055,N_78);
and U4633 (N_4633,N_1298,N_1962);
or U4634 (N_4634,N_1507,N_1143);
nor U4635 (N_4635,N_524,N_1954);
or U4636 (N_4636,N_1219,N_1791);
and U4637 (N_4637,N_2265,N_803);
or U4638 (N_4638,N_1953,N_1351);
nor U4639 (N_4639,N_1172,N_22);
or U4640 (N_4640,N_217,N_628);
and U4641 (N_4641,N_420,N_739);
or U4642 (N_4642,N_1615,N_685);
and U4643 (N_4643,N_190,N_860);
or U4644 (N_4644,N_93,N_2373);
nor U4645 (N_4645,N_118,N_2223);
nand U4646 (N_4646,N_1396,N_1600);
nand U4647 (N_4647,N_1049,N_102);
or U4648 (N_4648,N_743,N_844);
and U4649 (N_4649,N_368,N_2460);
and U4650 (N_4650,N_1875,N_246);
xnor U4651 (N_4651,N_1891,N_1792);
or U4652 (N_4652,N_1199,N_2225);
nand U4653 (N_4653,N_554,N_2411);
and U4654 (N_4654,N_1611,N_2053);
and U4655 (N_4655,N_278,N_2069);
and U4656 (N_4656,N_87,N_1101);
nand U4657 (N_4657,N_411,N_1687);
or U4658 (N_4658,N_2191,N_1379);
nand U4659 (N_4659,N_1670,N_907);
nor U4660 (N_4660,N_244,N_584);
and U4661 (N_4661,N_2414,N_1302);
nor U4662 (N_4662,N_1719,N_643);
and U4663 (N_4663,N_352,N_124);
and U4664 (N_4664,N_2267,N_1971);
nand U4665 (N_4665,N_1364,N_1505);
or U4666 (N_4666,N_1608,N_149);
or U4667 (N_4667,N_186,N_567);
nor U4668 (N_4668,N_946,N_2311);
or U4669 (N_4669,N_1440,N_226);
nor U4670 (N_4670,N_2283,N_186);
nor U4671 (N_4671,N_359,N_542);
nor U4672 (N_4672,N_1681,N_667);
or U4673 (N_4673,N_2458,N_2003);
xor U4674 (N_4674,N_1410,N_2105);
nor U4675 (N_4675,N_1056,N_1316);
nand U4676 (N_4676,N_1423,N_1128);
nor U4677 (N_4677,N_514,N_142);
and U4678 (N_4678,N_1445,N_52);
or U4679 (N_4679,N_826,N_43);
nand U4680 (N_4680,N_2402,N_2394);
nand U4681 (N_4681,N_324,N_1824);
and U4682 (N_4682,N_1418,N_986);
or U4683 (N_4683,N_679,N_2430);
nand U4684 (N_4684,N_690,N_2332);
or U4685 (N_4685,N_68,N_1548);
and U4686 (N_4686,N_1245,N_186);
xnor U4687 (N_4687,N_297,N_1836);
nor U4688 (N_4688,N_886,N_2);
nor U4689 (N_4689,N_13,N_965);
nand U4690 (N_4690,N_2349,N_1975);
or U4691 (N_4691,N_2074,N_2100);
and U4692 (N_4692,N_680,N_302);
or U4693 (N_4693,N_1519,N_1342);
or U4694 (N_4694,N_1511,N_33);
nand U4695 (N_4695,N_1404,N_1357);
nand U4696 (N_4696,N_71,N_2424);
or U4697 (N_4697,N_2368,N_1757);
or U4698 (N_4698,N_1302,N_1713);
nand U4699 (N_4699,N_1100,N_246);
and U4700 (N_4700,N_1192,N_1786);
or U4701 (N_4701,N_1363,N_639);
and U4702 (N_4702,N_1402,N_362);
and U4703 (N_4703,N_1073,N_1798);
xnor U4704 (N_4704,N_657,N_26);
nand U4705 (N_4705,N_2337,N_591);
and U4706 (N_4706,N_1348,N_333);
nor U4707 (N_4707,N_1969,N_503);
or U4708 (N_4708,N_1134,N_1504);
or U4709 (N_4709,N_741,N_352);
nor U4710 (N_4710,N_265,N_496);
and U4711 (N_4711,N_878,N_1004);
nor U4712 (N_4712,N_113,N_383);
and U4713 (N_4713,N_1679,N_2293);
nor U4714 (N_4714,N_2050,N_812);
xor U4715 (N_4715,N_1209,N_2352);
nor U4716 (N_4716,N_2213,N_592);
nand U4717 (N_4717,N_1808,N_1936);
nand U4718 (N_4718,N_2192,N_1540);
and U4719 (N_4719,N_1491,N_112);
or U4720 (N_4720,N_824,N_668);
or U4721 (N_4721,N_2160,N_210);
nor U4722 (N_4722,N_1395,N_668);
xor U4723 (N_4723,N_1720,N_662);
and U4724 (N_4724,N_2029,N_2457);
nand U4725 (N_4725,N_2459,N_1022);
and U4726 (N_4726,N_344,N_469);
nor U4727 (N_4727,N_1999,N_303);
and U4728 (N_4728,N_279,N_809);
and U4729 (N_4729,N_226,N_456);
or U4730 (N_4730,N_2295,N_909);
and U4731 (N_4731,N_1,N_1398);
and U4732 (N_4732,N_1951,N_158);
nor U4733 (N_4733,N_1369,N_1763);
nand U4734 (N_4734,N_876,N_1001);
and U4735 (N_4735,N_1587,N_1028);
or U4736 (N_4736,N_32,N_1253);
nand U4737 (N_4737,N_1884,N_2253);
nor U4738 (N_4738,N_2400,N_883);
nand U4739 (N_4739,N_2006,N_1217);
and U4740 (N_4740,N_1867,N_1485);
xnor U4741 (N_4741,N_702,N_1457);
or U4742 (N_4742,N_2474,N_1946);
nand U4743 (N_4743,N_1021,N_950);
nand U4744 (N_4744,N_204,N_743);
nor U4745 (N_4745,N_271,N_1131);
or U4746 (N_4746,N_752,N_842);
nand U4747 (N_4747,N_330,N_2071);
nand U4748 (N_4748,N_66,N_2216);
nand U4749 (N_4749,N_97,N_1167);
nor U4750 (N_4750,N_2412,N_717);
nand U4751 (N_4751,N_1672,N_905);
or U4752 (N_4752,N_1397,N_1708);
nor U4753 (N_4753,N_1970,N_2196);
nand U4754 (N_4754,N_1323,N_279);
nand U4755 (N_4755,N_110,N_2019);
nand U4756 (N_4756,N_449,N_371);
nor U4757 (N_4757,N_1332,N_1148);
nand U4758 (N_4758,N_957,N_1533);
and U4759 (N_4759,N_1460,N_2460);
and U4760 (N_4760,N_2482,N_793);
xor U4761 (N_4761,N_1156,N_2265);
nand U4762 (N_4762,N_507,N_2436);
nor U4763 (N_4763,N_121,N_855);
and U4764 (N_4764,N_1007,N_801);
and U4765 (N_4765,N_2358,N_1344);
and U4766 (N_4766,N_2166,N_87);
nand U4767 (N_4767,N_217,N_2136);
nor U4768 (N_4768,N_2262,N_1240);
or U4769 (N_4769,N_1139,N_1424);
nor U4770 (N_4770,N_1781,N_1853);
or U4771 (N_4771,N_1104,N_1531);
nand U4772 (N_4772,N_592,N_554);
and U4773 (N_4773,N_2118,N_283);
nand U4774 (N_4774,N_803,N_468);
xor U4775 (N_4775,N_210,N_2060);
xnor U4776 (N_4776,N_620,N_1044);
and U4777 (N_4777,N_1248,N_1589);
or U4778 (N_4778,N_1983,N_1615);
and U4779 (N_4779,N_1443,N_839);
nand U4780 (N_4780,N_1216,N_2331);
and U4781 (N_4781,N_14,N_33);
or U4782 (N_4782,N_827,N_2310);
nand U4783 (N_4783,N_530,N_1890);
nor U4784 (N_4784,N_2468,N_614);
or U4785 (N_4785,N_1623,N_653);
and U4786 (N_4786,N_207,N_1961);
nand U4787 (N_4787,N_1055,N_2195);
or U4788 (N_4788,N_88,N_805);
nand U4789 (N_4789,N_715,N_2167);
xor U4790 (N_4790,N_296,N_713);
and U4791 (N_4791,N_1107,N_1248);
nand U4792 (N_4792,N_843,N_1026);
and U4793 (N_4793,N_1156,N_1867);
nor U4794 (N_4794,N_505,N_650);
or U4795 (N_4795,N_2014,N_2227);
nor U4796 (N_4796,N_360,N_1647);
and U4797 (N_4797,N_2137,N_326);
and U4798 (N_4798,N_2069,N_520);
xnor U4799 (N_4799,N_441,N_721);
and U4800 (N_4800,N_781,N_965);
and U4801 (N_4801,N_1293,N_2398);
and U4802 (N_4802,N_176,N_1578);
nor U4803 (N_4803,N_2228,N_752);
nand U4804 (N_4804,N_215,N_1108);
nor U4805 (N_4805,N_350,N_2189);
nand U4806 (N_4806,N_798,N_1454);
nor U4807 (N_4807,N_1799,N_1935);
nand U4808 (N_4808,N_191,N_990);
nand U4809 (N_4809,N_1243,N_465);
nor U4810 (N_4810,N_562,N_1190);
nor U4811 (N_4811,N_977,N_1081);
or U4812 (N_4812,N_365,N_421);
nor U4813 (N_4813,N_452,N_2004);
or U4814 (N_4814,N_26,N_2006);
nor U4815 (N_4815,N_1327,N_1680);
or U4816 (N_4816,N_373,N_270);
and U4817 (N_4817,N_1737,N_862);
nand U4818 (N_4818,N_1485,N_943);
nand U4819 (N_4819,N_1401,N_1478);
and U4820 (N_4820,N_1474,N_261);
or U4821 (N_4821,N_785,N_1419);
nor U4822 (N_4822,N_1021,N_2296);
nor U4823 (N_4823,N_232,N_1140);
nand U4824 (N_4824,N_1562,N_513);
nor U4825 (N_4825,N_1484,N_172);
nor U4826 (N_4826,N_2170,N_1919);
and U4827 (N_4827,N_1599,N_561);
or U4828 (N_4828,N_1518,N_1162);
nor U4829 (N_4829,N_1935,N_411);
nor U4830 (N_4830,N_1760,N_1080);
and U4831 (N_4831,N_2335,N_1565);
or U4832 (N_4832,N_1348,N_2018);
and U4833 (N_4833,N_930,N_1920);
nor U4834 (N_4834,N_1471,N_732);
nor U4835 (N_4835,N_2153,N_1852);
nand U4836 (N_4836,N_692,N_1057);
or U4837 (N_4837,N_535,N_19);
nand U4838 (N_4838,N_1637,N_137);
or U4839 (N_4839,N_1871,N_206);
nor U4840 (N_4840,N_2150,N_641);
nor U4841 (N_4841,N_2311,N_2192);
and U4842 (N_4842,N_1170,N_1679);
or U4843 (N_4843,N_1383,N_1680);
xor U4844 (N_4844,N_2466,N_1592);
nand U4845 (N_4845,N_907,N_2262);
nand U4846 (N_4846,N_1364,N_827);
nand U4847 (N_4847,N_1459,N_2495);
and U4848 (N_4848,N_393,N_2336);
nor U4849 (N_4849,N_785,N_394);
nor U4850 (N_4850,N_412,N_430);
and U4851 (N_4851,N_1648,N_918);
or U4852 (N_4852,N_985,N_630);
nor U4853 (N_4853,N_295,N_307);
and U4854 (N_4854,N_1794,N_2229);
or U4855 (N_4855,N_1322,N_2289);
or U4856 (N_4856,N_590,N_1697);
and U4857 (N_4857,N_1126,N_1831);
and U4858 (N_4858,N_1175,N_380);
nor U4859 (N_4859,N_988,N_278);
nor U4860 (N_4860,N_2259,N_141);
and U4861 (N_4861,N_2244,N_1421);
or U4862 (N_4862,N_2325,N_1157);
xor U4863 (N_4863,N_43,N_23);
and U4864 (N_4864,N_104,N_642);
or U4865 (N_4865,N_1965,N_917);
and U4866 (N_4866,N_1091,N_252);
and U4867 (N_4867,N_1892,N_519);
xor U4868 (N_4868,N_304,N_1847);
and U4869 (N_4869,N_1683,N_2318);
nor U4870 (N_4870,N_1763,N_2335);
or U4871 (N_4871,N_2029,N_1957);
nand U4872 (N_4872,N_1541,N_339);
or U4873 (N_4873,N_702,N_1310);
and U4874 (N_4874,N_2486,N_1485);
nand U4875 (N_4875,N_1284,N_516);
xor U4876 (N_4876,N_2489,N_1660);
and U4877 (N_4877,N_1832,N_2198);
nor U4878 (N_4878,N_1644,N_1032);
nand U4879 (N_4879,N_1382,N_710);
or U4880 (N_4880,N_1319,N_1726);
nand U4881 (N_4881,N_1677,N_553);
and U4882 (N_4882,N_1279,N_877);
nand U4883 (N_4883,N_2115,N_1251);
and U4884 (N_4884,N_1763,N_957);
and U4885 (N_4885,N_2071,N_874);
and U4886 (N_4886,N_1547,N_2181);
nand U4887 (N_4887,N_1958,N_160);
nor U4888 (N_4888,N_2347,N_33);
xnor U4889 (N_4889,N_952,N_963);
nor U4890 (N_4890,N_860,N_323);
or U4891 (N_4891,N_1542,N_2309);
and U4892 (N_4892,N_495,N_793);
nor U4893 (N_4893,N_2279,N_1744);
nand U4894 (N_4894,N_1075,N_1924);
xnor U4895 (N_4895,N_2152,N_2051);
and U4896 (N_4896,N_2209,N_407);
or U4897 (N_4897,N_688,N_2327);
nand U4898 (N_4898,N_1781,N_1956);
nand U4899 (N_4899,N_1104,N_1857);
and U4900 (N_4900,N_2128,N_1063);
nand U4901 (N_4901,N_1760,N_944);
or U4902 (N_4902,N_112,N_2216);
xor U4903 (N_4903,N_1971,N_708);
or U4904 (N_4904,N_1982,N_1994);
nand U4905 (N_4905,N_579,N_2013);
and U4906 (N_4906,N_407,N_606);
or U4907 (N_4907,N_239,N_539);
or U4908 (N_4908,N_636,N_30);
or U4909 (N_4909,N_100,N_353);
and U4910 (N_4910,N_1538,N_1984);
or U4911 (N_4911,N_2273,N_1934);
nor U4912 (N_4912,N_694,N_2091);
nor U4913 (N_4913,N_2010,N_2149);
or U4914 (N_4914,N_2356,N_1049);
or U4915 (N_4915,N_625,N_219);
nor U4916 (N_4916,N_298,N_1462);
nand U4917 (N_4917,N_2430,N_480);
and U4918 (N_4918,N_29,N_915);
nand U4919 (N_4919,N_2360,N_689);
nand U4920 (N_4920,N_2066,N_232);
or U4921 (N_4921,N_1191,N_598);
or U4922 (N_4922,N_1326,N_1155);
and U4923 (N_4923,N_1813,N_494);
xnor U4924 (N_4924,N_258,N_1508);
xnor U4925 (N_4925,N_1134,N_1428);
nor U4926 (N_4926,N_521,N_664);
nor U4927 (N_4927,N_13,N_1751);
or U4928 (N_4928,N_1709,N_189);
nor U4929 (N_4929,N_2309,N_748);
or U4930 (N_4930,N_2275,N_2351);
or U4931 (N_4931,N_2293,N_1584);
nand U4932 (N_4932,N_2456,N_2445);
nand U4933 (N_4933,N_1184,N_1358);
nand U4934 (N_4934,N_83,N_184);
and U4935 (N_4935,N_958,N_1800);
nand U4936 (N_4936,N_1763,N_916);
nor U4937 (N_4937,N_1234,N_369);
and U4938 (N_4938,N_604,N_478);
nand U4939 (N_4939,N_763,N_663);
or U4940 (N_4940,N_260,N_1291);
nor U4941 (N_4941,N_499,N_570);
or U4942 (N_4942,N_1401,N_830);
nor U4943 (N_4943,N_919,N_59);
or U4944 (N_4944,N_327,N_1718);
xnor U4945 (N_4945,N_873,N_147);
and U4946 (N_4946,N_548,N_2470);
nor U4947 (N_4947,N_2010,N_1135);
or U4948 (N_4948,N_1363,N_19);
and U4949 (N_4949,N_2202,N_1814);
or U4950 (N_4950,N_276,N_1287);
nor U4951 (N_4951,N_179,N_1120);
nor U4952 (N_4952,N_2081,N_422);
nor U4953 (N_4953,N_1104,N_673);
nor U4954 (N_4954,N_1412,N_666);
xor U4955 (N_4955,N_1218,N_937);
nand U4956 (N_4956,N_1265,N_2097);
xnor U4957 (N_4957,N_2194,N_1570);
nand U4958 (N_4958,N_1372,N_855);
xnor U4959 (N_4959,N_516,N_1785);
xnor U4960 (N_4960,N_939,N_1111);
or U4961 (N_4961,N_784,N_1288);
and U4962 (N_4962,N_1916,N_367);
nor U4963 (N_4963,N_2218,N_2113);
xnor U4964 (N_4964,N_661,N_762);
and U4965 (N_4965,N_910,N_1414);
or U4966 (N_4966,N_1733,N_2371);
nor U4967 (N_4967,N_414,N_808);
nor U4968 (N_4968,N_2018,N_998);
nand U4969 (N_4969,N_1954,N_2172);
nand U4970 (N_4970,N_1396,N_1892);
and U4971 (N_4971,N_1706,N_829);
or U4972 (N_4972,N_1943,N_1391);
nor U4973 (N_4973,N_1517,N_351);
nand U4974 (N_4974,N_2138,N_1129);
nor U4975 (N_4975,N_483,N_1422);
and U4976 (N_4976,N_9,N_1814);
and U4977 (N_4977,N_416,N_545);
or U4978 (N_4978,N_1571,N_2171);
and U4979 (N_4979,N_1247,N_740);
and U4980 (N_4980,N_712,N_1772);
or U4981 (N_4981,N_2418,N_1882);
or U4982 (N_4982,N_1666,N_1425);
or U4983 (N_4983,N_2420,N_1723);
or U4984 (N_4984,N_1988,N_1919);
xnor U4985 (N_4985,N_556,N_1439);
xor U4986 (N_4986,N_529,N_1347);
nand U4987 (N_4987,N_1379,N_196);
nor U4988 (N_4988,N_1278,N_2308);
or U4989 (N_4989,N_1763,N_1344);
and U4990 (N_4990,N_1912,N_2112);
nand U4991 (N_4991,N_1636,N_1715);
nor U4992 (N_4992,N_2193,N_2314);
or U4993 (N_4993,N_1796,N_1391);
or U4994 (N_4994,N_311,N_1737);
and U4995 (N_4995,N_1574,N_442);
and U4996 (N_4996,N_845,N_308);
nor U4997 (N_4997,N_2362,N_968);
or U4998 (N_4998,N_1920,N_1401);
and U4999 (N_4999,N_1735,N_514);
nor UO_0 (O_0,N_4868,N_4437);
or UO_1 (O_1,N_3078,N_4473);
nand UO_2 (O_2,N_3428,N_4016);
nor UO_3 (O_3,N_3907,N_4991);
and UO_4 (O_4,N_4207,N_3633);
and UO_5 (O_5,N_3876,N_4966);
or UO_6 (O_6,N_4836,N_2600);
and UO_7 (O_7,N_3746,N_4316);
nand UO_8 (O_8,N_3850,N_3768);
xnor UO_9 (O_9,N_4338,N_3506);
or UO_10 (O_10,N_4755,N_4322);
and UO_11 (O_11,N_4169,N_4335);
or UO_12 (O_12,N_2615,N_3708);
nor UO_13 (O_13,N_4089,N_4173);
nand UO_14 (O_14,N_3679,N_3851);
nor UO_15 (O_15,N_4313,N_2709);
or UO_16 (O_16,N_2776,N_4131);
and UO_17 (O_17,N_4387,N_2720);
or UO_18 (O_18,N_3619,N_4901);
or UO_19 (O_19,N_2832,N_3995);
nor UO_20 (O_20,N_4133,N_3493);
nor UO_21 (O_21,N_4161,N_3088);
and UO_22 (O_22,N_3178,N_3824);
nand UO_23 (O_23,N_2791,N_2959);
and UO_24 (O_24,N_2957,N_4332);
nand UO_25 (O_25,N_3914,N_3789);
xnor UO_26 (O_26,N_2514,N_3138);
nor UO_27 (O_27,N_2714,N_3969);
and UO_28 (O_28,N_3266,N_3339);
nor UO_29 (O_29,N_4350,N_3892);
or UO_30 (O_30,N_2795,N_4993);
and UO_31 (O_31,N_3930,N_3406);
nand UO_32 (O_32,N_4855,N_3321);
or UO_33 (O_33,N_3523,N_3718);
xnor UO_34 (O_34,N_4974,N_4256);
nor UO_35 (O_35,N_2763,N_3298);
xnor UO_36 (O_36,N_3095,N_4240);
or UO_37 (O_37,N_4429,N_2836);
nor UO_38 (O_38,N_3479,N_3029);
and UO_39 (O_39,N_4179,N_3181);
and UO_40 (O_40,N_3262,N_3141);
and UO_41 (O_41,N_3887,N_2751);
xor UO_42 (O_42,N_3113,N_3407);
nor UO_43 (O_43,N_3466,N_2858);
nand UO_44 (O_44,N_3000,N_4502);
nand UO_45 (O_45,N_3719,N_3588);
nor UO_46 (O_46,N_4467,N_3946);
and UO_47 (O_47,N_4760,N_3476);
or UO_48 (O_48,N_3102,N_3680);
xor UO_49 (O_49,N_3180,N_3239);
or UO_50 (O_50,N_3449,N_4233);
or UO_51 (O_51,N_2515,N_2851);
or UO_52 (O_52,N_4985,N_4996);
nor UO_53 (O_53,N_4057,N_4585);
or UO_54 (O_54,N_2519,N_3290);
and UO_55 (O_55,N_3791,N_2727);
or UO_56 (O_56,N_4630,N_3873);
nor UO_57 (O_57,N_3084,N_4523);
nand UO_58 (O_58,N_2511,N_3412);
nand UO_59 (O_59,N_3405,N_4378);
and UO_60 (O_60,N_4551,N_4653);
nor UO_61 (O_61,N_4587,N_2712);
nor UO_62 (O_62,N_3073,N_2575);
and UO_63 (O_63,N_3620,N_4894);
nor UO_64 (O_64,N_4845,N_4869);
xor UO_65 (O_65,N_3223,N_4438);
nand UO_66 (O_66,N_3852,N_4399);
nand UO_67 (O_67,N_2995,N_4266);
nor UO_68 (O_68,N_4556,N_2530);
or UO_69 (O_69,N_4430,N_3305);
and UO_70 (O_70,N_3338,N_2885);
nor UO_71 (O_71,N_3698,N_4675);
nor UO_72 (O_72,N_3859,N_4809);
nand UO_73 (O_73,N_4673,N_4522);
and UO_74 (O_74,N_4424,N_4106);
or UO_75 (O_75,N_3883,N_2861);
nor UO_76 (O_76,N_3597,N_4371);
nor UO_77 (O_77,N_4029,N_2550);
xnor UO_78 (O_78,N_3750,N_3365);
or UO_79 (O_79,N_3643,N_4053);
nor UO_80 (O_80,N_3958,N_4690);
nor UO_81 (O_81,N_4039,N_4406);
nand UO_82 (O_82,N_4643,N_3641);
nor UO_83 (O_83,N_3310,N_3133);
and UO_84 (O_84,N_3772,N_2860);
nor UO_85 (O_85,N_3042,N_3190);
nor UO_86 (O_86,N_4397,N_4317);
nor UO_87 (O_87,N_3404,N_2632);
nor UO_88 (O_88,N_3694,N_4705);
or UO_89 (O_89,N_4216,N_3528);
or UO_90 (O_90,N_2797,N_2730);
or UO_91 (O_91,N_4746,N_3215);
or UO_92 (O_92,N_4490,N_3236);
and UO_93 (O_93,N_4631,N_4944);
and UO_94 (O_94,N_4766,N_2900);
nand UO_95 (O_95,N_3870,N_2571);
and UO_96 (O_96,N_4476,N_4489);
or UO_97 (O_97,N_2926,N_4457);
or UO_98 (O_98,N_4129,N_2658);
nor UO_99 (O_99,N_3773,N_4446);
nand UO_100 (O_100,N_2748,N_3543);
or UO_101 (O_101,N_4104,N_3940);
nand UO_102 (O_102,N_4336,N_2934);
or UO_103 (O_103,N_3297,N_4533);
nand UO_104 (O_104,N_4685,N_2839);
and UO_105 (O_105,N_3311,N_2782);
nor UO_106 (O_106,N_4183,N_3714);
or UO_107 (O_107,N_3612,N_3544);
nand UO_108 (O_108,N_3625,N_3955);
and UO_109 (O_109,N_4752,N_3599);
nor UO_110 (O_110,N_3375,N_3259);
and UO_111 (O_111,N_2798,N_4958);
nand UO_112 (O_112,N_3507,N_4135);
nor UO_113 (O_113,N_2588,N_2696);
nor UO_114 (O_114,N_4539,N_4727);
and UO_115 (O_115,N_3739,N_3669);
and UO_116 (O_116,N_3896,N_3212);
or UO_117 (O_117,N_3706,N_4491);
xor UO_118 (O_118,N_2713,N_3950);
and UO_119 (O_119,N_4427,N_3168);
xnor UO_120 (O_120,N_2509,N_4455);
and UO_121 (O_121,N_2887,N_4887);
and UO_122 (O_122,N_3580,N_3659);
nor UO_123 (O_123,N_3396,N_4851);
nor UO_124 (O_124,N_3977,N_4051);
nand UO_125 (O_125,N_3674,N_2721);
nor UO_126 (O_126,N_4024,N_4941);
or UO_127 (O_127,N_3598,N_2950);
or UO_128 (O_128,N_3471,N_3713);
and UO_129 (O_129,N_4549,N_3462);
or UO_130 (O_130,N_3410,N_2523);
xnor UO_131 (O_131,N_4662,N_3877);
nand UO_132 (O_132,N_4413,N_4823);
nor UO_133 (O_133,N_2780,N_2645);
nand UO_134 (O_134,N_3971,N_4890);
and UO_135 (O_135,N_3926,N_3023);
nand UO_136 (O_136,N_3885,N_4817);
nand UO_137 (O_137,N_4262,N_3584);
nor UO_138 (O_138,N_3662,N_4695);
nand UO_139 (O_139,N_4986,N_3313);
and UO_140 (O_140,N_3842,N_3165);
xnor UO_141 (O_141,N_3710,N_2976);
nor UO_142 (O_142,N_3312,N_4834);
and UO_143 (O_143,N_3388,N_4791);
nor UO_144 (O_144,N_3485,N_4711);
nor UO_145 (O_145,N_4238,N_4733);
xor UO_146 (O_146,N_4006,N_3119);
nand UO_147 (O_147,N_4250,N_4698);
and UO_148 (O_148,N_4444,N_4544);
or UO_149 (O_149,N_4440,N_3214);
nand UO_150 (O_150,N_3837,N_3254);
nor UO_151 (O_151,N_2915,N_4616);
nor UO_152 (O_152,N_4883,N_3497);
and UO_153 (O_153,N_2503,N_3085);
nor UO_154 (O_154,N_4815,N_4911);
nor UO_155 (O_155,N_2967,N_2742);
nand UO_156 (O_156,N_2582,N_4758);
nand UO_157 (O_157,N_3723,N_2767);
nand UO_158 (O_158,N_4156,N_2913);
nor UO_159 (O_159,N_4793,N_3702);
and UO_160 (O_160,N_3070,N_3393);
nor UO_161 (O_161,N_4829,N_2775);
and UO_162 (O_162,N_3024,N_2538);
or UO_163 (O_163,N_2969,N_4190);
or UO_164 (O_164,N_2690,N_3468);
or UO_165 (O_165,N_4261,N_3126);
nor UO_166 (O_166,N_3947,N_3059);
xnor UO_167 (O_167,N_2716,N_3448);
xor UO_168 (O_168,N_3547,N_3350);
and UO_169 (O_169,N_3415,N_4712);
and UO_170 (O_170,N_3826,N_4011);
nor UO_171 (O_171,N_3848,N_4661);
nand UO_172 (O_172,N_4543,N_4124);
xor UO_173 (O_173,N_4557,N_3502);
or UO_174 (O_174,N_2638,N_3340);
xor UO_175 (O_175,N_2842,N_4421);
xnor UO_176 (O_176,N_4891,N_2924);
nor UO_177 (O_177,N_3792,N_4367);
nor UO_178 (O_178,N_4276,N_3777);
nand UO_179 (O_179,N_2796,N_3052);
xnor UO_180 (O_180,N_3954,N_3774);
nor UO_181 (O_181,N_3752,N_2512);
and UO_182 (O_182,N_3732,N_2689);
nand UO_183 (O_183,N_4975,N_4723);
and UO_184 (O_184,N_3890,N_2545);
or UO_185 (O_185,N_3736,N_3053);
and UO_186 (O_186,N_2951,N_2908);
and UO_187 (O_187,N_3093,N_4193);
nor UO_188 (O_188,N_4728,N_4434);
or UO_189 (O_189,N_2589,N_3246);
and UO_190 (O_190,N_4824,N_4748);
or UO_191 (O_191,N_2522,N_4152);
or UO_192 (O_192,N_3771,N_3280);
nor UO_193 (O_193,N_3342,N_3671);
nor UO_194 (O_194,N_4003,N_4045);
nand UO_195 (O_195,N_3120,N_2949);
nand UO_196 (O_196,N_4860,N_3764);
nand UO_197 (O_197,N_3900,N_3548);
or UO_198 (O_198,N_4200,N_2529);
and UO_199 (O_199,N_4763,N_3274);
and UO_200 (O_200,N_4120,N_4431);
nand UO_201 (O_201,N_4886,N_2554);
nand UO_202 (O_202,N_3307,N_4504);
and UO_203 (O_203,N_3423,N_4602);
or UO_204 (O_204,N_2527,N_2867);
and UO_205 (O_205,N_3668,N_3492);
nor UO_206 (O_206,N_4617,N_2906);
nand UO_207 (O_207,N_3443,N_4931);
nand UO_208 (O_208,N_4244,N_4352);
nor UO_209 (O_209,N_3916,N_2826);
nand UO_210 (O_210,N_4191,N_2986);
or UO_211 (O_211,N_4061,N_4475);
or UO_212 (O_212,N_3302,N_4570);
nor UO_213 (O_213,N_3648,N_2789);
or UO_214 (O_214,N_4203,N_2784);
and UO_215 (O_215,N_3068,N_4981);
nand UO_216 (O_216,N_3153,N_2733);
xor UO_217 (O_217,N_3435,N_4402);
and UO_218 (O_218,N_3802,N_3117);
nand UO_219 (O_219,N_3169,N_3928);
or UO_220 (O_220,N_4806,N_2962);
nor UO_221 (O_221,N_2807,N_3224);
and UO_222 (O_222,N_3967,N_2664);
and UO_223 (O_223,N_3391,N_3610);
nand UO_224 (O_224,N_3039,N_4162);
xnor UO_225 (O_225,N_2657,N_3952);
nand UO_226 (O_226,N_4485,N_2679);
nor UO_227 (O_227,N_3650,N_2777);
xnor UO_228 (O_228,N_4997,N_3596);
and UO_229 (O_229,N_2506,N_3701);
and UO_230 (O_230,N_2694,N_2786);
and UO_231 (O_231,N_3160,N_3992);
or UO_232 (O_232,N_3461,N_3681);
nand UO_233 (O_233,N_4885,N_2580);
or UO_234 (O_234,N_3623,N_4713);
and UO_235 (O_235,N_4672,N_3812);
and UO_236 (O_236,N_3457,N_4667);
or UO_237 (O_237,N_3099,N_4299);
and UO_238 (O_238,N_2546,N_4784);
and UO_239 (O_239,N_4268,N_2703);
or UO_240 (O_240,N_2945,N_4938);
xnor UO_241 (O_241,N_3208,N_4507);
and UO_242 (O_242,N_4325,N_3634);
or UO_243 (O_243,N_3226,N_4524);
and UO_244 (O_244,N_3047,N_4189);
nand UO_245 (O_245,N_3006,N_3519);
and UO_246 (O_246,N_4914,N_3062);
or UO_247 (O_247,N_2813,N_3477);
nor UO_248 (O_248,N_4506,N_4870);
or UO_249 (O_249,N_3478,N_2827);
nor UO_250 (O_250,N_4331,N_3177);
and UO_251 (O_251,N_3937,N_2876);
or UO_252 (O_252,N_4611,N_2810);
nand UO_253 (O_253,N_4050,N_3376);
or UO_254 (O_254,N_4664,N_4805);
xnor UO_255 (O_255,N_3373,N_4468);
nand UO_256 (O_256,N_4951,N_4984);
or UO_257 (O_257,N_2927,N_3722);
or UO_258 (O_258,N_3411,N_3503);
or UO_259 (O_259,N_4426,N_4908);
nand UO_260 (O_260,N_4807,N_4419);
nand UO_261 (O_261,N_2830,N_3766);
xor UO_262 (O_262,N_3285,N_4454);
xor UO_263 (O_263,N_4001,N_3216);
or UO_264 (O_264,N_3903,N_3514);
xnor UO_265 (O_265,N_4239,N_3293);
and UO_266 (O_266,N_4394,N_4565);
nor UO_267 (O_267,N_2693,N_3089);
nor UO_268 (O_268,N_3202,N_3558);
nand UO_269 (O_269,N_3326,N_4647);
nor UO_270 (O_270,N_3974,N_4952);
nand UO_271 (O_271,N_3018,N_2640);
nor UO_272 (O_272,N_3615,N_4841);
nor UO_273 (O_273,N_4732,N_2592);
or UO_274 (O_274,N_4609,N_3804);
nand UO_275 (O_275,N_3983,N_4798);
xor UO_276 (O_276,N_4967,N_2850);
or UO_277 (O_277,N_3225,N_4407);
nor UO_278 (O_278,N_2912,N_2656);
and UO_279 (O_279,N_3034,N_2923);
nand UO_280 (O_280,N_3164,N_2731);
and UO_281 (O_281,N_4111,N_3127);
and UO_282 (O_282,N_4982,N_3721);
nor UO_283 (O_283,N_4998,N_2975);
nand UO_284 (O_284,N_4368,N_4148);
xnor UO_285 (O_285,N_2920,N_2625);
or UO_286 (O_286,N_4655,N_4154);
nand UO_287 (O_287,N_4280,N_2997);
nor UO_288 (O_288,N_4820,N_4246);
or UO_289 (O_289,N_2991,N_3530);
and UO_290 (O_290,N_3409,N_4054);
xor UO_291 (O_291,N_4899,N_4821);
nand UO_292 (O_292,N_4272,N_4580);
xnor UO_293 (O_293,N_2977,N_3935);
or UO_294 (O_294,N_3585,N_3198);
or UO_295 (O_295,N_3499,N_4279);
or UO_296 (O_296,N_2740,N_3372);
nand UO_297 (O_297,N_4925,N_2766);
nand UO_298 (O_298,N_2812,N_3013);
nor UO_299 (O_299,N_3155,N_2551);
xor UO_300 (O_300,N_4634,N_4146);
and UO_301 (O_301,N_2916,N_3727);
and UO_302 (O_302,N_3617,N_4666);
xor UO_303 (O_303,N_3045,N_3689);
nor UO_304 (O_304,N_3056,N_3253);
and UO_305 (O_305,N_4094,N_4158);
and UO_306 (O_306,N_4962,N_4620);
nand UO_307 (O_307,N_3187,N_4002);
nor UO_308 (O_308,N_3816,N_4058);
nor UO_309 (O_309,N_3581,N_3031);
nand UO_310 (O_310,N_3193,N_3818);
nand UO_311 (O_311,N_2753,N_3071);
nand UO_312 (O_312,N_2953,N_2785);
xnor UO_313 (O_313,N_3835,N_4277);
and UO_314 (O_314,N_4144,N_4471);
or UO_315 (O_315,N_2570,N_3437);
xor UO_316 (O_316,N_3090,N_4835);
or UO_317 (O_317,N_4777,N_2960);
or UO_318 (O_318,N_4345,N_4703);
or UO_319 (O_319,N_3335,N_2573);
nor UO_320 (O_320,N_3505,N_3026);
or UO_321 (O_321,N_4498,N_3344);
or UO_322 (O_322,N_4314,N_4854);
or UO_323 (O_323,N_3081,N_4588);
nor UO_324 (O_324,N_4961,N_4346);
and UO_325 (O_325,N_4375,N_3866);
or UO_326 (O_326,N_4369,N_4330);
nand UO_327 (O_327,N_3158,N_2761);
nand UO_328 (O_328,N_2702,N_4903);
xnor UO_329 (O_329,N_4005,N_3316);
nand UO_330 (O_330,N_4761,N_2608);
and UO_331 (O_331,N_4360,N_4028);
nor UO_332 (O_332,N_3686,N_3025);
nand UO_333 (O_333,N_3798,N_2828);
or UO_334 (O_334,N_3844,N_4725);
nor UO_335 (O_335,N_4686,N_3072);
nand UO_336 (O_336,N_3389,N_3712);
or UO_337 (O_337,N_3807,N_3136);
nand UO_338 (O_338,N_3629,N_4852);
nand UO_339 (O_339,N_4692,N_4160);
xnor UO_340 (O_340,N_3352,N_3430);
xor UO_341 (O_341,N_3277,N_2935);
xor UO_342 (O_342,N_4186,N_3963);
nand UO_343 (O_343,N_4063,N_2889);
or UO_344 (O_344,N_4818,N_3346);
or UO_345 (O_345,N_2502,N_3209);
or UO_346 (O_346,N_3270,N_3703);
nand UO_347 (O_347,N_4859,N_4227);
nor UO_348 (O_348,N_3252,N_4321);
or UO_349 (O_349,N_3128,N_2877);
or UO_350 (O_350,N_3613,N_2966);
or UO_351 (O_351,N_4292,N_4788);
nor UO_352 (O_352,N_2574,N_3110);
xor UO_353 (O_353,N_4167,N_3016);
nand UO_354 (O_354,N_2806,N_2899);
nor UO_355 (O_355,N_2864,N_4720);
nor UO_356 (O_356,N_4928,N_4449);
xnor UO_357 (O_357,N_4983,N_3758);
and UO_358 (O_358,N_3783,N_3343);
nor UO_359 (O_359,N_4568,N_4949);
and UO_360 (O_360,N_3540,N_3003);
nor UO_361 (O_361,N_4714,N_3920);
xor UO_362 (O_362,N_4939,N_4826);
or UO_363 (O_363,N_3327,N_2528);
or UO_364 (O_364,N_2549,N_4649);
nand UO_365 (O_365,N_4278,N_3378);
or UO_366 (O_366,N_3427,N_3744);
xnor UO_367 (O_367,N_4584,N_2643);
nor UO_368 (O_368,N_3044,N_3590);
nand UO_369 (O_369,N_4354,N_4592);
nand UO_370 (O_370,N_2622,N_4796);
and UO_371 (O_371,N_2855,N_4790);
and UO_372 (O_372,N_2859,N_4125);
or UO_373 (O_373,N_2540,N_2888);
and UO_374 (O_374,N_3904,N_3606);
xor UO_375 (O_375,N_4948,N_2983);
nor UO_376 (O_376,N_4339,N_4283);
nand UO_377 (O_377,N_3303,N_4493);
xnor UO_378 (O_378,N_2717,N_2618);
and UO_379 (O_379,N_2524,N_2955);
and UO_380 (O_380,N_3429,N_4518);
or UO_381 (O_381,N_3861,N_4221);
xor UO_382 (O_382,N_2590,N_3104);
and UO_383 (O_383,N_3233,N_3549);
or UO_384 (O_384,N_3251,N_3639);
or UO_385 (O_385,N_4819,N_3436);
and UO_386 (O_386,N_3913,N_3973);
or UO_387 (O_387,N_2965,N_3576);
or UO_388 (O_388,N_4676,N_4882);
and UO_389 (O_389,N_4654,N_4517);
xor UO_390 (O_390,N_2704,N_3336);
nor UO_391 (O_391,N_4373,N_3616);
and UO_392 (O_392,N_3299,N_3834);
or UO_393 (O_393,N_4978,N_3172);
nand UO_394 (O_394,N_4563,N_3103);
nand UO_395 (O_395,N_2517,N_4285);
nand UO_396 (O_396,N_3425,N_3387);
nor UO_397 (O_397,N_3994,N_4211);
or UO_398 (O_398,N_4030,N_4065);
or UO_399 (O_399,N_4922,N_3809);
xor UO_400 (O_400,N_4802,N_3897);
nor UO_401 (O_401,N_4126,N_3354);
nor UO_402 (O_402,N_2773,N_3030);
xor UO_403 (O_403,N_3011,N_4496);
nor UO_404 (O_404,N_3148,N_3384);
xor UO_405 (O_405,N_3979,N_3027);
and UO_406 (O_406,N_4451,N_3864);
nand UO_407 (O_407,N_4060,N_3917);
xnor UO_408 (O_408,N_4857,N_3765);
nand UO_409 (O_409,N_2848,N_3453);
or UO_410 (O_410,N_4668,N_4513);
xnor UO_411 (O_411,N_3156,N_4503);
xnor UO_412 (O_412,N_2998,N_3551);
nor UO_413 (O_413,N_4249,N_4572);
nor UO_414 (O_414,N_2650,N_3715);
nand UO_415 (O_415,N_4202,N_4046);
or UO_416 (O_416,N_4935,N_4621);
nand UO_417 (O_417,N_3366,N_3194);
and UO_418 (O_418,N_4640,N_4940);
or UO_419 (O_419,N_2964,N_3586);
nand UO_420 (O_420,N_4532,N_3332);
nand UO_421 (O_421,N_3105,N_4707);
and UO_422 (O_422,N_3879,N_4281);
nor UO_423 (O_423,N_4619,N_4917);
or UO_424 (O_424,N_4194,N_2567);
nor UO_425 (O_425,N_4749,N_4391);
nand UO_426 (O_426,N_4736,N_3445);
nor UO_427 (O_427,N_4509,N_2662);
nand UO_428 (O_428,N_4593,N_3112);
nand UO_429 (O_429,N_4499,N_4579);
nand UO_430 (O_430,N_3434,N_4562);
or UO_431 (O_431,N_3788,N_2936);
nand UO_432 (O_432,N_3557,N_3894);
nor UO_433 (O_433,N_2683,N_4618);
or UO_434 (O_434,N_3289,N_4768);
and UO_435 (O_435,N_4370,N_4601);
nor UO_436 (O_436,N_3654,N_4987);
nor UO_437 (O_437,N_4874,N_2938);
or UO_438 (O_438,N_4838,N_3657);
and UO_439 (O_439,N_4880,N_2891);
nor UO_440 (O_440,N_2849,N_2521);
xnor UO_441 (O_441,N_3403,N_4514);
or UO_442 (O_442,N_4264,N_3454);
or UO_443 (O_443,N_2699,N_4577);
and UO_444 (O_444,N_2667,N_4849);
nor UO_445 (O_445,N_3481,N_2882);
nand UO_446 (O_446,N_2746,N_3605);
nand UO_447 (O_447,N_3508,N_2921);
or UO_448 (O_448,N_3709,N_4537);
or UO_449 (O_449,N_4048,N_3589);
and UO_450 (O_450,N_3587,N_4157);
nor UO_451 (O_451,N_2970,N_3111);
nand UO_452 (O_452,N_3521,N_3398);
nand UO_453 (O_453,N_2881,N_4107);
nor UO_454 (O_454,N_3057,N_4778);
nand UO_455 (O_455,N_4583,N_4687);
nor UO_456 (O_456,N_4595,N_3949);
or UO_457 (O_457,N_4535,N_3618);
nand UO_458 (O_458,N_3699,N_4143);
nand UO_459 (O_459,N_2628,N_2678);
and UO_460 (O_460,N_4358,N_4724);
and UO_461 (O_461,N_4865,N_3256);
and UO_462 (O_462,N_4347,N_4773);
and UO_463 (O_463,N_3728,N_2531);
or UO_464 (O_464,N_4409,N_4892);
nand UO_465 (O_465,N_3424,N_3683);
or UO_466 (O_466,N_2584,N_4478);
or UO_467 (O_467,N_2597,N_2805);
or UO_468 (O_468,N_2654,N_2647);
or UO_469 (O_469,N_4488,N_4401);
nor UO_470 (O_470,N_4355,N_4481);
and UO_471 (O_471,N_3700,N_4109);
nand UO_472 (O_472,N_2852,N_4635);
nor UO_473 (O_473,N_3797,N_4756);
or UO_474 (O_474,N_4574,N_4036);
nand UO_475 (O_475,N_2617,N_4780);
or UO_476 (O_476,N_3724,N_3296);
nand UO_477 (O_477,N_3532,N_3960);
or UO_478 (O_478,N_4230,N_3306);
xnor UO_479 (O_479,N_4964,N_3046);
or UO_480 (O_480,N_3761,N_3091);
nor UO_481 (O_481,N_4145,N_4453);
or UO_482 (O_482,N_3922,N_3658);
xnor UO_483 (O_483,N_4198,N_2542);
and UO_484 (O_484,N_3624,N_3573);
and UO_485 (O_485,N_4069,N_3621);
xor UO_486 (O_486,N_3731,N_4432);
nand UO_487 (O_487,N_3526,N_3123);
and UO_488 (O_488,N_3309,N_4295);
nor UO_489 (O_489,N_3474,N_3325);
nor UO_490 (O_490,N_4665,N_3707);
nor UO_491 (O_491,N_2516,N_4251);
or UO_492 (O_492,N_3315,N_4767);
nor UO_493 (O_493,N_3570,N_3951);
or UO_494 (O_494,N_4270,N_3183);
nor UO_495 (O_495,N_4670,N_3908);
or UO_496 (O_496,N_4830,N_2907);
and UO_497 (O_497,N_4573,N_4603);
nand UO_498 (O_498,N_2939,N_4552);
xor UO_499 (O_499,N_3222,N_4924);
nor UO_500 (O_500,N_4090,N_4581);
nand UO_501 (O_501,N_4388,N_3819);
nor UO_502 (O_502,N_3759,N_2904);
nor UO_503 (O_503,N_3363,N_4804);
nor UO_504 (O_504,N_4785,N_2666);
nand UO_505 (O_505,N_4717,N_2972);
and UO_506 (O_506,N_4237,N_3781);
nor UO_507 (O_507,N_4452,N_2728);
or UO_508 (O_508,N_3323,N_4605);
and UO_509 (O_509,N_2871,N_2685);
nand UO_510 (O_510,N_2982,N_2999);
nand UO_511 (O_511,N_4297,N_3260);
nand UO_512 (O_512,N_3919,N_4482);
nand UO_513 (O_513,N_3267,N_2541);
nor UO_514 (O_514,N_4702,N_3331);
xor UO_515 (O_515,N_2818,N_3821);
nand UO_516 (O_516,N_2801,N_2845);
or UO_517 (O_517,N_3051,N_3012);
nand UO_518 (O_518,N_3368,N_3693);
or UO_519 (O_519,N_3628,N_3911);
nand UO_520 (O_520,N_3394,N_4235);
nor UO_521 (O_521,N_4792,N_2557);
nand UO_522 (O_522,N_4121,N_2598);
nor UO_523 (O_523,N_4636,N_3320);
nand UO_524 (O_524,N_3083,N_4074);
nor UO_525 (O_525,N_4907,N_4715);
and UO_526 (O_526,N_3822,N_3785);
xnor UO_527 (O_527,N_4988,N_3058);
and UO_528 (O_528,N_3291,N_2612);
or UO_529 (O_529,N_3795,N_3483);
xnor UO_530 (O_530,N_3362,N_2989);
or UO_531 (O_531,N_2578,N_2781);
nand UO_532 (O_532,N_4863,N_3060);
or UO_533 (O_533,N_4615,N_4548);
or UO_534 (O_534,N_2510,N_3318);
nor UO_535 (O_535,N_4363,N_4178);
nor UO_536 (O_536,N_3292,N_2772);
nand UO_537 (O_537,N_4118,N_3636);
or UO_538 (O_538,N_3667,N_3632);
and UO_539 (O_539,N_4436,N_4520);
nor UO_540 (O_540,N_3998,N_4497);
or UO_541 (O_541,N_4055,N_2536);
or UO_542 (O_542,N_3978,N_2886);
or UO_543 (O_543,N_3355,N_4881);
xor UO_544 (O_544,N_3002,N_2707);
nand UO_545 (O_545,N_4015,N_3048);
and UO_546 (O_546,N_4366,N_3849);
or UO_547 (O_547,N_2583,N_3086);
and UO_548 (O_548,N_4267,N_4384);
nand UO_549 (O_549,N_4091,N_3317);
and UO_550 (O_550,N_4070,N_4433);
or UO_551 (O_551,N_2980,N_4274);
and UO_552 (O_552,N_4729,N_3504);
xnor UO_553 (O_553,N_2892,N_2873);
nor UO_554 (O_554,N_4742,N_4688);
and UO_555 (O_555,N_3880,N_4304);
or UO_556 (O_556,N_3061,N_2743);
nand UO_557 (O_557,N_4501,N_3097);
nor UO_558 (O_558,N_4787,N_2778);
nand UO_559 (O_559,N_3142,N_4624);
nor UO_560 (O_560,N_4177,N_2897);
or UO_561 (O_561,N_4683,N_3738);
nor UO_562 (O_562,N_2823,N_4710);
nand UO_563 (O_563,N_3972,N_3525);
or UO_564 (O_564,N_4208,N_4171);
xor UO_565 (O_565,N_2534,N_3152);
and UO_566 (O_566,N_3696,N_3855);
nand UO_567 (O_567,N_2726,N_4613);
nor UO_568 (O_568,N_2961,N_3279);
nor UO_569 (O_569,N_3121,N_3392);
nor UO_570 (O_570,N_2800,N_3450);
or UO_571 (O_571,N_4078,N_4782);
or UO_572 (O_572,N_4210,N_3829);
or UO_573 (O_573,N_2878,N_3975);
and UO_574 (O_574,N_2847,N_4632);
nand UO_575 (O_575,N_2553,N_3170);
and UO_576 (O_576,N_3936,N_3841);
or UO_577 (O_577,N_3122,N_3601);
and UO_578 (O_578,N_4734,N_2670);
nand UO_579 (O_579,N_3985,N_2526);
and UO_580 (O_580,N_4677,N_3402);
and UO_581 (O_581,N_4598,N_3494);
and UO_582 (O_582,N_3692,N_4900);
nor UO_583 (O_583,N_2620,N_3075);
nand UO_584 (O_584,N_3108,N_3498);
nand UO_585 (O_585,N_4417,N_3942);
nor UO_586 (O_586,N_4275,N_4164);
or UO_587 (O_587,N_3414,N_3562);
nand UO_588 (O_588,N_2841,N_4428);
nand UO_589 (O_589,N_3195,N_4709);
or UO_590 (O_590,N_2659,N_3263);
nand UO_591 (O_591,N_3022,N_2505);
nand UO_592 (O_592,N_4416,N_4487);
nor UO_593 (O_593,N_3163,N_3269);
or UO_594 (O_594,N_2535,N_4392);
xnor UO_595 (O_595,N_2682,N_3775);
nand UO_596 (O_596,N_3909,N_4088);
nand UO_597 (O_597,N_3087,N_4955);
nand UO_598 (O_598,N_3467,N_2862);
nor UO_599 (O_599,N_3371,N_4324);
nand UO_600 (O_600,N_4674,N_2639);
xor UO_601 (O_601,N_3990,N_2838);
nor UO_602 (O_602,N_3349,N_2809);
or UO_603 (O_603,N_3231,N_3552);
and UO_604 (O_604,N_3808,N_4594);
nor UO_605 (O_605,N_2518,N_4606);
nor UO_606 (O_606,N_3130,N_3534);
nand UO_607 (O_607,N_3283,N_2605);
and UO_608 (O_608,N_4977,N_2931);
xor UO_609 (O_609,N_3150,N_2946);
nor UO_610 (O_610,N_3074,N_3337);
nor UO_611 (O_611,N_4386,N_4495);
nor UO_612 (O_612,N_3591,N_3230);
xnor UO_613 (O_613,N_3753,N_3697);
nor UO_614 (O_614,N_4225,N_2613);
nor UO_615 (O_615,N_3386,N_3945);
or UO_616 (O_616,N_3778,N_4614);
or UO_617 (O_617,N_4916,N_3055);
and UO_618 (O_618,N_2856,N_4464);
xor UO_619 (O_619,N_2919,N_4085);
or UO_620 (O_620,N_3980,N_4172);
nand UO_621 (O_621,N_4521,N_4282);
or UO_622 (O_622,N_4878,N_4571);
nor UO_623 (O_623,N_2835,N_4212);
and UO_624 (O_624,N_2593,N_3541);
xnor UO_625 (O_625,N_4273,N_2865);
xor UO_626 (O_626,N_4128,N_3754);
nand UO_627 (O_627,N_2652,N_4098);
nand UO_628 (O_628,N_3268,N_2783);
or UO_629 (O_629,N_3536,N_4443);
nor UO_630 (O_630,N_3154,N_4258);
nand UO_631 (O_631,N_3441,N_4414);
xor UO_632 (O_632,N_4231,N_3054);
or UO_633 (O_633,N_4234,N_4669);
nand UO_634 (O_634,N_4694,N_3682);
or UO_635 (O_635,N_2520,N_3203);
nor UO_636 (O_636,N_3927,N_4372);
nand UO_637 (O_637,N_3893,N_4260);
nand UO_638 (O_638,N_3749,N_4744);
nand UO_639 (O_639,N_3288,N_3948);
nand UO_640 (O_640,N_3201,N_3833);
and UO_641 (O_641,N_3569,N_2829);
nor UO_642 (O_642,N_3092,N_4023);
and UO_643 (O_643,N_3872,N_4771);
or UO_644 (O_644,N_4365,N_4289);
and UO_645 (O_645,N_4021,N_2764);
or UO_646 (O_646,N_4229,N_2533);
or UO_647 (O_647,N_3455,N_2884);
nand UO_648 (O_648,N_3308,N_2684);
or UO_649 (O_649,N_3999,N_3473);
nor UO_650 (O_650,N_2586,N_3171);
or UO_651 (O_651,N_3238,N_4622);
nand UO_652 (O_652,N_2599,N_2952);
or UO_653 (O_653,N_4960,N_4130);
xor UO_654 (O_654,N_4168,N_3653);
nand UO_655 (O_655,N_2729,N_4393);
nand UO_656 (O_656,N_4302,N_4486);
or UO_657 (O_657,N_3801,N_4799);
or UO_658 (O_658,N_3257,N_3295);
nor UO_659 (O_659,N_3014,N_4979);
nand UO_660 (O_660,N_3432,N_4213);
or UO_661 (O_661,N_2674,N_2606);
and UO_662 (O_662,N_3912,N_3964);
nor UO_663 (O_663,N_3527,N_3395);
nand UO_664 (O_664,N_4842,N_4110);
nand UO_665 (O_665,N_3741,N_3577);
or UO_666 (O_666,N_3082,N_4862);
xnor UO_667 (O_667,N_4344,N_3762);
nor UO_668 (O_668,N_3080,N_4850);
nor UO_669 (O_669,N_4765,N_3814);
xnor UO_670 (O_670,N_4462,N_4762);
nor UO_671 (O_671,N_2653,N_4348);
xnor UO_672 (O_672,N_4362,N_2820);
or UO_673 (O_673,N_4546,N_3167);
xnor UO_674 (O_674,N_3115,N_4699);
xnor UO_675 (O_675,N_3825,N_4018);
or UO_676 (O_676,N_3770,N_4696);
or UO_677 (O_677,N_3374,N_4341);
nor UO_678 (O_678,N_4382,N_4312);
nor UO_679 (O_679,N_3300,N_4627);
nand UO_680 (O_680,N_2942,N_4127);
nor UO_681 (O_681,N_3459,N_3250);
and UO_682 (O_682,N_4943,N_4663);
xnor UO_683 (O_683,N_4590,N_2634);
and UO_684 (O_684,N_4309,N_4757);
or UO_685 (O_685,N_4236,N_4970);
nand UO_686 (O_686,N_3776,N_3444);
or UO_687 (O_687,N_4992,N_3592);
or UO_688 (O_688,N_3649,N_3511);
nand UO_689 (O_689,N_2648,N_3079);
nand UO_690 (O_690,N_4972,N_3007);
nor UO_691 (O_691,N_4254,N_4904);
nor UO_692 (O_692,N_4027,N_3490);
nand UO_693 (O_693,N_3192,N_4326);
nor UO_694 (O_694,N_3417,N_4340);
and UO_695 (O_695,N_2697,N_3575);
or UO_696 (O_696,N_4946,N_4329);
or UO_697 (O_697,N_2739,N_2623);
or UO_698 (O_698,N_4781,N_4108);
nor UO_699 (O_699,N_2954,N_3579);
xnor UO_700 (O_700,N_3756,N_4474);
nor UO_701 (O_701,N_4896,N_4064);
and UO_702 (O_702,N_2711,N_3475);
and UO_703 (O_703,N_3273,N_4448);
nand UO_704 (O_704,N_4252,N_2635);
or UO_705 (O_705,N_2819,N_3067);
nor UO_706 (O_706,N_3134,N_4113);
or UO_707 (O_707,N_2596,N_4722);
nor UO_708 (O_708,N_3938,N_3638);
or UO_709 (O_709,N_4066,N_4284);
or UO_710 (O_710,N_4123,N_4994);
nor UO_711 (O_711,N_4515,N_4528);
nand UO_712 (O_712,N_4035,N_3933);
nand UO_713 (O_713,N_4813,N_4052);
and UO_714 (O_714,N_2698,N_3546);
xnor UO_715 (O_715,N_4902,N_3348);
nor UO_716 (O_716,N_3247,N_3867);
nand UO_717 (O_717,N_3237,N_4999);
or UO_718 (O_718,N_3932,N_4450);
nand UO_719 (O_719,N_3341,N_2883);
and UO_720 (O_720,N_4192,N_2757);
nor UO_721 (O_721,N_3294,N_4351);
nor UO_722 (O_722,N_4816,N_3660);
nor UO_723 (O_723,N_2691,N_2537);
or UO_724 (O_724,N_4534,N_2624);
or UO_725 (O_725,N_3763,N_3255);
xor UO_726 (O_726,N_2799,N_2552);
and UO_727 (O_727,N_4719,N_4385);
or UO_728 (O_728,N_4651,N_3482);
nor UO_729 (O_729,N_2843,N_4383);
nor UO_730 (O_730,N_4554,N_3509);
or UO_731 (O_731,N_4512,N_3962);
and UO_732 (O_732,N_3678,N_3780);
nand UO_733 (O_733,N_3559,N_4848);
nand UO_734 (O_734,N_3691,N_3881);
or UO_735 (O_735,N_4356,N_4610);
nand UO_736 (O_736,N_4968,N_4652);
or UO_737 (O_737,N_3001,N_3281);
nor UO_738 (O_738,N_3561,N_2610);
nor UO_739 (O_739,N_2507,N_4139);
nor UO_740 (O_740,N_4242,N_4291);
or UO_741 (O_741,N_3282,N_3676);
or UO_742 (O_742,N_4418,N_3704);
or UO_743 (O_743,N_3539,N_2724);
nor UO_744 (O_744,N_2869,N_2513);
and UO_745 (O_745,N_3760,N_4753);
nor UO_746 (O_746,N_3651,N_4846);
xor UO_747 (O_747,N_2736,N_3578);
or UO_748 (O_748,N_3333,N_3440);
nor UO_749 (O_749,N_4844,N_3271);
nand UO_750 (O_750,N_3345,N_4073);
xor UO_751 (O_751,N_3240,N_2633);
or UO_752 (O_752,N_3672,N_2825);
nor UO_753 (O_753,N_3537,N_3426);
nor UO_754 (O_754,N_3495,N_4912);
xor UO_755 (O_755,N_3210,N_2539);
nor UO_756 (O_756,N_3555,N_4176);
and UO_757 (O_757,N_2508,N_4561);
nand UO_758 (O_758,N_3690,N_3243);
xnor UO_759 (O_759,N_2692,N_2671);
and UO_760 (O_760,N_2846,N_4980);
nor UO_761 (O_761,N_4420,N_3442);
nor UO_762 (O_762,N_4459,N_3032);
and UO_763 (O_763,N_3106,N_4206);
xor UO_764 (O_764,N_4327,N_3159);
or UO_765 (O_765,N_2644,N_2948);
xor UO_766 (O_766,N_3229,N_4650);
nor UO_767 (O_767,N_4084,N_4693);
or UO_768 (O_768,N_2708,N_4214);
and UO_769 (O_769,N_3245,N_4625);
or UO_770 (O_770,N_4828,N_3249);
and UO_771 (O_771,N_2868,N_3593);
nor UO_772 (O_772,N_3740,N_3695);
nand UO_773 (O_773,N_2978,N_4795);
nand UO_774 (O_774,N_3664,N_3151);
nand UO_775 (O_775,N_2500,N_2735);
xor UO_776 (O_776,N_4165,N_2973);
nand UO_777 (O_777,N_3748,N_4077);
and UO_778 (O_778,N_4477,N_2706);
nor UO_779 (O_779,N_2669,N_4701);
or UO_780 (O_780,N_4929,N_3640);
and UO_781 (O_781,N_4741,N_4228);
or UO_782 (O_782,N_4405,N_4447);
and UO_783 (O_783,N_3463,N_3100);
nand UO_784 (O_784,N_3512,N_2688);
nor UO_785 (O_785,N_4025,N_3647);
and UO_786 (O_786,N_4087,N_4578);
and UO_787 (O_787,N_4494,N_4257);
xnor UO_788 (O_788,N_3400,N_4410);
nor UO_789 (O_789,N_4017,N_2814);
xnor UO_790 (O_790,N_4589,N_3162);
nand UO_791 (O_791,N_3635,N_3517);
or UO_792 (O_792,N_3351,N_3554);
or UO_793 (O_793,N_3401,N_4076);
or UO_794 (O_794,N_3314,N_2905);
and UO_795 (O_795,N_3845,N_3218);
nor UO_796 (O_796,N_2929,N_4540);
or UO_797 (O_797,N_3941,N_3747);
nor UO_798 (O_798,N_4680,N_3131);
nor UO_799 (O_799,N_3145,N_3929);
nor UO_800 (O_800,N_3968,N_4287);
and UO_801 (O_801,N_4945,N_3370);
and UO_802 (O_802,N_3996,N_4315);
nor UO_803 (O_803,N_3779,N_2577);
xor UO_804 (O_804,N_3556,N_4174);
and UO_805 (O_805,N_4895,N_3381);
or UO_806 (O_806,N_2673,N_2760);
nand UO_807 (O_807,N_4657,N_3832);
nor UO_808 (O_808,N_2563,N_4905);
and UO_809 (O_809,N_4328,N_3050);
nor UO_810 (O_810,N_4918,N_2677);
or UO_811 (O_811,N_3076,N_4479);
and UO_812 (O_812,N_4223,N_3730);
or UO_813 (O_813,N_4963,N_4062);
xor UO_814 (O_814,N_4103,N_3729);
and UO_815 (O_815,N_3529,N_4950);
nor UO_816 (O_816,N_3399,N_2947);
or UO_817 (O_817,N_4959,N_3737);
nand UO_818 (O_818,N_4641,N_3149);
xor UO_819 (O_819,N_3421,N_4357);
xor UO_820 (O_820,N_4072,N_2788);
and UO_821 (O_821,N_4364,N_4068);
nand UO_822 (O_822,N_2771,N_4884);
or UO_823 (O_823,N_2663,N_3098);
nand UO_824 (O_824,N_4196,N_3094);
and UO_825 (O_825,N_2630,N_3921);
nand UO_826 (O_826,N_3066,N_3132);
or UO_827 (O_827,N_4456,N_3364);
nand UO_828 (O_828,N_2655,N_4879);
or UO_829 (O_829,N_2587,N_4840);
or UO_830 (O_830,N_3820,N_4575);
and UO_831 (O_831,N_2745,N_3456);
nand UO_832 (O_832,N_4608,N_4875);
nor UO_833 (O_833,N_3431,N_2821);
nor UO_834 (O_834,N_2564,N_3853);
nand UO_835 (O_835,N_4095,N_2723);
and UO_836 (O_836,N_3185,N_3287);
xnor UO_837 (O_837,N_3500,N_3028);
or UO_838 (O_838,N_3301,N_2585);
nor UO_839 (O_839,N_3358,N_4973);
nand UO_840 (O_840,N_3646,N_3357);
nand UO_841 (O_841,N_2626,N_3188);
nor UO_842 (O_842,N_3064,N_4141);
nand UO_843 (O_843,N_4628,N_2544);
nor UO_844 (O_844,N_3472,N_4898);
nor UO_845 (O_845,N_4175,N_2984);
nor UO_846 (O_846,N_3882,N_3199);
or UO_847 (O_847,N_4505,N_4954);
nand UO_848 (O_848,N_4545,N_3888);
nor UO_849 (O_849,N_3176,N_3191);
and UO_850 (O_850,N_2705,N_3196);
or UO_851 (O_851,N_2759,N_4395);
or UO_852 (O_852,N_3836,N_2824);
nand UO_853 (O_853,N_4827,N_3232);
or UO_854 (O_854,N_4492,N_4812);
nor UO_855 (O_855,N_2994,N_4296);
or UO_856 (O_856,N_4014,N_3161);
and UO_857 (O_857,N_4185,N_4747);
or UO_858 (O_858,N_3786,N_4269);
or UO_859 (O_859,N_4529,N_3757);
nand UO_860 (O_860,N_3987,N_3970);
nor UO_861 (O_861,N_2560,N_4038);
nor UO_862 (O_862,N_4215,N_3717);
nor UO_863 (O_863,N_4913,N_3377);
nor UO_864 (O_864,N_3884,N_2614);
xor UO_865 (O_865,N_3420,N_3810);
nand UO_866 (O_866,N_2768,N_4219);
nor UO_867 (O_867,N_4519,N_3036);
nor UO_868 (O_868,N_4310,N_3009);
or UO_869 (O_869,N_3043,N_3329);
or UO_870 (O_870,N_3107,N_4659);
or UO_871 (O_871,N_2933,N_2719);
nor UO_872 (O_872,N_4217,N_3334);
and UO_873 (O_873,N_2840,N_3823);
nand UO_874 (O_874,N_3670,N_2591);
xor UO_875 (O_875,N_4466,N_3684);
nor UO_876 (O_876,N_2930,N_4019);
nor UO_877 (O_877,N_3328,N_3745);
nand UO_878 (O_878,N_4012,N_4342);
nor UO_879 (O_879,N_4629,N_3063);
or UO_880 (O_880,N_3515,N_3953);
nand UO_881 (O_881,N_3157,N_3182);
or UO_882 (O_882,N_4319,N_3235);
nor UO_883 (O_883,N_2911,N_3416);
and UO_884 (O_884,N_3666,N_4199);
xor UO_885 (O_885,N_2993,N_2854);
or UO_886 (O_886,N_4731,N_4232);
or UO_887 (O_887,N_3889,N_3685);
nor UO_888 (O_888,N_3275,N_2822);
nand UO_889 (O_889,N_4245,N_4379);
or UO_890 (O_890,N_3258,N_2641);
nand UO_891 (O_891,N_4558,N_4538);
and UO_892 (O_892,N_4008,N_4645);
nand UO_893 (O_893,N_2569,N_4441);
and UO_894 (O_894,N_2725,N_2675);
nor UO_895 (O_895,N_4586,N_3419);
and UO_896 (O_896,N_2595,N_3594);
xor UO_897 (O_897,N_4114,N_4550);
xor UO_898 (O_898,N_3652,N_3261);
and UO_899 (O_899,N_3571,N_4374);
nor UO_900 (O_900,N_3886,N_4381);
nor UO_901 (O_901,N_2802,N_3956);
nor UO_902 (O_902,N_4516,N_4801);
nand UO_903 (O_903,N_3322,N_3353);
and UO_904 (O_904,N_3501,N_4853);
or UO_905 (O_905,N_2974,N_2940);
or UO_906 (O_906,N_4380,N_3874);
nor UO_907 (O_907,N_4658,N_2642);
or UO_908 (O_908,N_2971,N_3452);
and UO_909 (O_909,N_2649,N_2562);
or UO_910 (O_910,N_3019,N_4000);
and UO_911 (O_911,N_4294,N_3993);
or UO_912 (O_912,N_2937,N_4163);
xor UO_913 (O_913,N_4953,N_3918);
nor UO_914 (O_914,N_2715,N_3213);
nand UO_915 (O_915,N_4306,N_3397);
nand UO_916 (O_916,N_3447,N_3831);
nor UO_917 (O_917,N_3065,N_3189);
xnor UO_918 (O_918,N_3661,N_4255);
nand UO_919 (O_919,N_2774,N_2750);
nand UO_920 (O_920,N_3566,N_4915);
nor UO_921 (O_921,N_4445,N_3988);
and UO_922 (O_922,N_4876,N_3125);
and UO_923 (O_923,N_3875,N_4783);
xnor UO_924 (O_924,N_3630,N_4527);
nor UO_925 (O_925,N_4510,N_2555);
and UO_926 (O_926,N_2901,N_4754);
nand UO_927 (O_927,N_4205,N_4942);
and UO_928 (O_928,N_4009,N_4423);
and UO_929 (O_929,N_4976,N_3488);
and UO_930 (O_930,N_3863,N_4140);
and UO_931 (O_931,N_2893,N_4007);
or UO_932 (O_932,N_4837,N_3535);
and UO_933 (O_933,N_4730,N_3146);
nor UO_934 (O_934,N_4933,N_4990);
xnor UO_935 (O_935,N_4839,N_3600);
or UO_936 (O_936,N_2880,N_4947);
or UO_937 (O_937,N_3166,N_4706);
or UO_938 (O_938,N_3743,N_2581);
or UO_939 (O_939,N_4691,N_4097);
and UO_940 (O_940,N_4224,N_4637);
nand UO_941 (O_941,N_2803,N_3241);
and UO_942 (O_942,N_2749,N_4772);
nand UO_943 (O_943,N_4833,N_3734);
nor UO_944 (O_944,N_2853,N_3784);
or UO_945 (O_945,N_2896,N_3957);
and UO_946 (O_946,N_3204,N_2928);
or UO_947 (O_947,N_4726,N_3520);
or UO_948 (O_948,N_2879,N_3206);
or UO_949 (O_949,N_2572,N_2831);
or UO_950 (O_950,N_4684,N_3568);
nor UO_951 (O_951,N_4803,N_3140);
nand UO_952 (O_952,N_3487,N_4075);
nand UO_953 (O_953,N_3197,N_4271);
nor UO_954 (O_954,N_4136,N_3109);
nand UO_955 (O_955,N_2601,N_2769);
nand UO_956 (O_956,N_3604,N_3038);
and UO_957 (O_957,N_4800,N_4043);
or UO_958 (O_958,N_3868,N_4769);
and UO_959 (O_959,N_3602,N_3567);
or UO_960 (O_960,N_4843,N_3742);
xor UO_961 (O_961,N_4847,N_4737);
and UO_962 (O_962,N_2604,N_4576);
xor UO_963 (O_963,N_4472,N_3642);
and UO_964 (O_964,N_3118,N_4149);
nand UO_965 (O_965,N_3595,N_2787);
or UO_966 (O_966,N_4153,N_2548);
and UO_967 (O_967,N_3319,N_3284);
nor UO_968 (O_968,N_4463,N_4412);
nand UO_969 (O_969,N_2661,N_4642);
nand UO_970 (O_970,N_4415,N_4831);
nor UO_971 (O_971,N_3857,N_4263);
xor UO_972 (O_972,N_4656,N_4079);
xnor UO_973 (O_973,N_4927,N_3173);
and UO_974 (O_974,N_4049,N_4866);
xnor UO_975 (O_975,N_4010,N_3813);
nor UO_976 (O_976,N_4708,N_3144);
and UO_977 (O_977,N_4797,N_4770);
and UO_978 (O_978,N_2910,N_2629);
nand UO_979 (O_979,N_4411,N_2922);
xnor UO_980 (O_980,N_3793,N_3644);
nand UO_981 (O_981,N_4508,N_4604);
xor UO_982 (O_982,N_3276,N_4422);
xnor UO_983 (O_983,N_4483,N_2987);
or UO_984 (O_984,N_2637,N_3496);
xnor UO_985 (O_985,N_2817,N_3200);
or UO_986 (O_986,N_3227,N_3572);
or UO_987 (O_987,N_2834,N_2676);
and UO_988 (O_988,N_4439,N_2565);
xnor UO_989 (O_989,N_4026,N_4248);
xnor UO_990 (O_990,N_3021,N_3304);
xor UO_991 (O_991,N_2875,N_4033);
or UO_992 (O_992,N_2844,N_4919);
nand UO_993 (O_993,N_3854,N_2815);
or UO_994 (O_994,N_2804,N_2758);
or UO_995 (O_995,N_2602,N_2609);
nor UO_996 (O_996,N_4671,N_4555);
or UO_997 (O_997,N_3856,N_2755);
nor UO_998 (O_998,N_4117,N_4034);
and UO_999 (O_999,N_2990,N_4134);
endmodule