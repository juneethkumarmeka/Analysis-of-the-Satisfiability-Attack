module basic_500_3000_500_3_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_138,In_19);
and U1 (N_1,In_209,In_311);
xnor U2 (N_2,In_286,In_77);
and U3 (N_3,In_38,In_438);
xnor U4 (N_4,In_488,In_173);
or U5 (N_5,In_81,In_490);
and U6 (N_6,In_481,In_136);
xnor U7 (N_7,In_235,In_402);
nand U8 (N_8,In_79,In_171);
or U9 (N_9,In_52,In_53);
xnor U10 (N_10,In_320,In_266);
and U11 (N_11,In_116,In_483);
nand U12 (N_12,In_247,In_404);
nand U13 (N_13,In_225,In_400);
nand U14 (N_14,In_407,In_399);
and U15 (N_15,In_78,In_239);
nor U16 (N_16,In_122,In_299);
or U17 (N_17,In_195,In_434);
nand U18 (N_18,In_83,In_255);
or U19 (N_19,In_415,In_137);
xor U20 (N_20,In_289,In_62);
nor U21 (N_21,In_228,In_470);
and U22 (N_22,In_336,In_73);
and U23 (N_23,In_442,In_484);
or U24 (N_24,In_39,In_84);
nand U25 (N_25,In_242,In_460);
or U26 (N_26,In_129,In_319);
nor U27 (N_27,In_347,In_268);
or U28 (N_28,In_107,In_294);
nand U29 (N_29,In_212,In_193);
xnor U30 (N_30,In_218,In_448);
nor U31 (N_31,In_334,In_388);
and U32 (N_32,In_21,In_202);
nor U33 (N_33,In_271,In_42);
nor U34 (N_34,In_248,In_493);
or U35 (N_35,In_91,In_94);
or U36 (N_36,In_232,In_310);
nor U37 (N_37,In_439,In_31);
nor U38 (N_38,In_12,In_128);
nor U39 (N_39,In_132,In_449);
nand U40 (N_40,In_304,In_187);
and U41 (N_41,In_330,In_494);
and U42 (N_42,In_468,In_51);
xor U43 (N_43,In_204,In_170);
nand U44 (N_44,In_405,In_177);
nor U45 (N_45,In_121,In_223);
nand U46 (N_46,In_326,In_6);
or U47 (N_47,In_13,In_227);
or U48 (N_48,In_18,In_236);
nor U49 (N_49,In_179,In_420);
or U50 (N_50,In_348,In_131);
nor U51 (N_51,In_328,In_208);
nor U52 (N_52,In_335,In_469);
nand U53 (N_53,In_274,In_45);
nand U54 (N_54,In_422,In_443);
or U55 (N_55,In_251,In_48);
and U56 (N_56,In_215,In_359);
and U57 (N_57,In_314,In_30);
nand U58 (N_58,In_102,In_486);
nand U59 (N_59,In_67,In_34);
xnor U60 (N_60,In_72,In_161);
or U61 (N_61,In_124,In_267);
xnor U62 (N_62,In_292,In_57);
xnor U63 (N_63,In_188,In_40);
nor U64 (N_64,In_302,In_444);
nor U65 (N_65,In_146,In_385);
or U66 (N_66,In_387,In_303);
or U67 (N_67,In_35,In_164);
xnor U68 (N_68,In_190,In_279);
xor U69 (N_69,In_47,In_181);
and U70 (N_70,In_214,In_15);
nand U71 (N_71,In_126,In_368);
nor U72 (N_72,In_143,In_441);
or U73 (N_73,In_452,In_191);
nor U74 (N_74,In_224,In_440);
and U75 (N_75,In_307,In_245);
or U76 (N_76,In_284,In_298);
xnor U77 (N_77,In_380,In_36);
xor U78 (N_78,In_7,In_447);
or U79 (N_79,In_23,In_437);
and U80 (N_80,In_206,In_98);
nor U81 (N_81,In_60,In_489);
or U82 (N_82,In_345,In_382);
nand U83 (N_83,In_159,In_259);
xnor U84 (N_84,In_295,In_254);
nand U85 (N_85,In_133,In_360);
nor U86 (N_86,In_192,In_479);
nand U87 (N_87,In_65,In_55);
and U88 (N_88,In_166,In_419);
xor U89 (N_89,In_480,In_104);
nor U90 (N_90,In_197,In_211);
or U91 (N_91,In_134,In_340);
nand U92 (N_92,In_397,In_222);
nor U93 (N_93,In_27,In_401);
nand U94 (N_94,In_198,In_273);
and U95 (N_95,In_29,In_112);
nand U96 (N_96,In_463,In_33);
nand U97 (N_97,In_82,In_346);
or U98 (N_98,In_182,In_375);
nor U99 (N_99,In_100,In_99);
xor U100 (N_100,In_376,In_329);
and U101 (N_101,In_464,In_408);
nor U102 (N_102,In_264,In_312);
or U103 (N_103,In_277,In_50);
or U104 (N_104,In_260,In_466);
xnor U105 (N_105,In_8,In_66);
nor U106 (N_106,In_272,In_451);
xnor U107 (N_107,In_315,In_4);
nand U108 (N_108,In_213,In_325);
and U109 (N_109,In_243,In_395);
and U110 (N_110,In_357,In_123);
nand U111 (N_111,In_372,In_370);
nand U112 (N_112,In_231,In_280);
and U113 (N_113,In_109,In_432);
or U114 (N_114,In_85,In_467);
nor U115 (N_115,In_2,In_207);
nand U116 (N_116,In_369,In_64);
and U117 (N_117,In_416,In_409);
nand U118 (N_118,In_497,In_436);
or U119 (N_119,In_344,In_477);
and U120 (N_120,In_322,In_194);
or U121 (N_121,In_398,In_117);
xor U122 (N_122,In_257,In_285);
or U123 (N_123,In_461,In_165);
nor U124 (N_124,In_475,In_403);
nor U125 (N_125,In_374,In_185);
nand U126 (N_126,In_189,In_113);
nand U127 (N_127,In_278,In_324);
xnor U128 (N_128,In_371,In_427);
and U129 (N_129,In_183,In_144);
or U130 (N_130,In_366,In_421);
or U131 (N_131,In_41,In_269);
xnor U132 (N_132,In_96,In_390);
nor U133 (N_133,In_108,In_201);
nand U134 (N_134,In_430,In_332);
nand U135 (N_135,In_379,In_300);
nor U136 (N_136,In_384,In_450);
and U137 (N_137,In_97,In_22);
xnor U138 (N_138,In_262,In_381);
or U139 (N_139,In_17,In_354);
nand U140 (N_140,In_240,In_364);
and U141 (N_141,In_423,In_63);
nor U142 (N_142,In_59,In_200);
or U143 (N_143,In_323,In_418);
or U144 (N_144,In_9,In_281);
nor U145 (N_145,In_391,In_106);
nand U146 (N_146,In_20,In_424);
or U147 (N_147,In_317,In_141);
xnor U148 (N_148,In_76,In_458);
and U149 (N_149,In_496,In_69);
or U150 (N_150,In_275,In_352);
nand U151 (N_151,In_61,In_140);
nor U152 (N_152,In_338,In_435);
nor U153 (N_153,In_263,In_349);
nand U154 (N_154,In_162,In_238);
and U155 (N_155,In_25,In_168);
and U156 (N_156,In_495,In_355);
nor U157 (N_157,In_377,In_54);
or U158 (N_158,In_499,In_291);
or U159 (N_159,In_210,In_256);
nor U160 (N_160,In_158,In_417);
nor U161 (N_161,In_92,In_175);
or U162 (N_162,In_226,In_492);
nand U163 (N_163,In_205,In_341);
xnor U164 (N_164,In_428,In_49);
or U165 (N_165,In_396,In_101);
xor U166 (N_166,In_216,In_425);
or U167 (N_167,In_241,In_203);
nor U168 (N_168,In_220,In_176);
or U169 (N_169,In_44,In_414);
and U170 (N_170,In_130,In_118);
and U171 (N_171,In_270,In_174);
nor U172 (N_172,In_58,In_457);
nand U173 (N_173,In_482,In_71);
nor U174 (N_174,In_10,In_237);
nand U175 (N_175,In_337,In_393);
nor U176 (N_176,In_308,In_156);
and U177 (N_177,In_28,In_473);
nor U178 (N_178,In_343,In_86);
or U179 (N_179,In_485,In_43);
nand U180 (N_180,In_105,In_313);
nand U181 (N_181,In_253,In_155);
nor U182 (N_182,In_288,In_287);
and U183 (N_183,In_290,In_16);
or U184 (N_184,In_476,In_229);
or U185 (N_185,In_265,In_406);
or U186 (N_186,In_362,In_217);
or U187 (N_187,In_367,In_412);
nor U188 (N_188,In_306,In_180);
nand U189 (N_189,In_305,In_453);
nor U190 (N_190,In_454,In_321);
or U191 (N_191,In_353,In_37);
or U192 (N_192,In_465,In_250);
and U193 (N_193,In_445,In_14);
and U194 (N_194,In_246,In_361);
and U195 (N_195,In_178,In_373);
and U196 (N_196,In_87,In_145);
nor U197 (N_197,In_93,In_358);
xnor U198 (N_198,In_411,In_149);
nand U199 (N_199,In_433,In_498);
nand U200 (N_200,In_90,In_363);
nand U201 (N_201,In_462,In_301);
and U202 (N_202,In_413,In_426);
xor U203 (N_203,In_233,In_219);
or U204 (N_204,In_316,In_68);
and U205 (N_205,In_167,In_89);
and U206 (N_206,In_154,In_75);
or U207 (N_207,In_139,In_429);
or U208 (N_208,In_186,In_351);
nand U209 (N_209,In_160,In_386);
nand U210 (N_210,In_5,In_0);
nor U211 (N_211,In_276,In_157);
and U212 (N_212,In_318,In_148);
or U213 (N_213,In_56,In_70);
nor U214 (N_214,In_297,In_196);
or U215 (N_215,In_125,In_472);
nor U216 (N_216,In_249,In_169);
or U217 (N_217,In_103,In_95);
nand U218 (N_218,In_394,In_151);
nor U219 (N_219,In_356,In_410);
nor U220 (N_220,In_199,In_261);
or U221 (N_221,In_11,In_333);
nor U222 (N_222,In_150,In_392);
nor U223 (N_223,In_455,In_258);
and U224 (N_224,In_244,In_142);
nand U225 (N_225,In_350,In_456);
and U226 (N_226,In_365,In_46);
nor U227 (N_227,In_296,In_147);
nor U228 (N_228,In_110,In_293);
xor U229 (N_229,In_389,In_74);
or U230 (N_230,In_282,In_230);
and U231 (N_231,In_331,In_184);
or U232 (N_232,In_153,In_26);
or U233 (N_233,In_474,In_252);
and U234 (N_234,In_487,In_378);
or U235 (N_235,In_24,In_135);
or U236 (N_236,In_120,In_114);
nand U237 (N_237,In_446,In_172);
and U238 (N_238,In_339,In_127);
and U239 (N_239,In_431,In_115);
xor U240 (N_240,In_309,In_478);
or U241 (N_241,In_221,In_80);
nor U242 (N_242,In_3,In_471);
nor U243 (N_243,In_459,In_491);
xor U244 (N_244,In_32,In_342);
nand U245 (N_245,In_1,In_88);
nor U246 (N_246,In_152,In_111);
nor U247 (N_247,In_234,In_383);
nand U248 (N_248,In_119,In_163);
and U249 (N_249,In_283,In_327);
or U250 (N_250,In_233,In_216);
and U251 (N_251,In_416,In_57);
nand U252 (N_252,In_461,In_360);
nor U253 (N_253,In_454,In_406);
or U254 (N_254,In_361,In_62);
nand U255 (N_255,In_120,In_100);
nand U256 (N_256,In_84,In_243);
nor U257 (N_257,In_380,In_113);
or U258 (N_258,In_179,In_477);
nor U259 (N_259,In_219,In_143);
nand U260 (N_260,In_365,In_224);
or U261 (N_261,In_74,In_228);
and U262 (N_262,In_224,In_99);
nor U263 (N_263,In_348,In_35);
or U264 (N_264,In_465,In_427);
nand U265 (N_265,In_307,In_497);
and U266 (N_266,In_307,In_294);
and U267 (N_267,In_43,In_397);
and U268 (N_268,In_222,In_134);
nand U269 (N_269,In_478,In_433);
nand U270 (N_270,In_117,In_473);
nand U271 (N_271,In_189,In_172);
and U272 (N_272,In_295,In_401);
or U273 (N_273,In_288,In_337);
nor U274 (N_274,In_154,In_77);
nand U275 (N_275,In_412,In_142);
and U276 (N_276,In_172,In_109);
nor U277 (N_277,In_472,In_482);
nand U278 (N_278,In_126,In_8);
and U279 (N_279,In_299,In_399);
nor U280 (N_280,In_404,In_293);
or U281 (N_281,In_123,In_220);
nor U282 (N_282,In_30,In_29);
nand U283 (N_283,In_6,In_14);
or U284 (N_284,In_84,In_112);
or U285 (N_285,In_170,In_168);
and U286 (N_286,In_299,In_259);
and U287 (N_287,In_296,In_272);
or U288 (N_288,In_393,In_413);
or U289 (N_289,In_221,In_10);
or U290 (N_290,In_33,In_32);
nand U291 (N_291,In_458,In_385);
or U292 (N_292,In_304,In_165);
or U293 (N_293,In_55,In_275);
nor U294 (N_294,In_241,In_57);
nand U295 (N_295,In_141,In_168);
or U296 (N_296,In_375,In_50);
nor U297 (N_297,In_152,In_56);
or U298 (N_298,In_463,In_439);
or U299 (N_299,In_284,In_235);
nand U300 (N_300,In_205,In_90);
nor U301 (N_301,In_188,In_153);
nor U302 (N_302,In_251,In_270);
and U303 (N_303,In_426,In_243);
or U304 (N_304,In_489,In_496);
and U305 (N_305,In_190,In_469);
and U306 (N_306,In_430,In_225);
nand U307 (N_307,In_466,In_91);
nor U308 (N_308,In_475,In_220);
xnor U309 (N_309,In_278,In_249);
or U310 (N_310,In_191,In_356);
and U311 (N_311,In_442,In_16);
nand U312 (N_312,In_450,In_44);
nand U313 (N_313,In_124,In_185);
xor U314 (N_314,In_364,In_15);
nor U315 (N_315,In_118,In_412);
nand U316 (N_316,In_391,In_338);
or U317 (N_317,In_386,In_121);
or U318 (N_318,In_179,In_490);
or U319 (N_319,In_202,In_498);
nor U320 (N_320,In_190,In_71);
nand U321 (N_321,In_408,In_98);
nand U322 (N_322,In_201,In_198);
and U323 (N_323,In_341,In_315);
xnor U324 (N_324,In_425,In_358);
nand U325 (N_325,In_317,In_232);
nor U326 (N_326,In_158,In_290);
and U327 (N_327,In_208,In_477);
and U328 (N_328,In_158,In_234);
xnor U329 (N_329,In_273,In_463);
nor U330 (N_330,In_381,In_417);
nor U331 (N_331,In_352,In_237);
nor U332 (N_332,In_258,In_233);
nand U333 (N_333,In_346,In_418);
nor U334 (N_334,In_193,In_194);
nor U335 (N_335,In_268,In_424);
and U336 (N_336,In_121,In_132);
and U337 (N_337,In_279,In_344);
xnor U338 (N_338,In_298,In_494);
xor U339 (N_339,In_180,In_481);
or U340 (N_340,In_299,In_253);
or U341 (N_341,In_267,In_108);
and U342 (N_342,In_341,In_68);
xnor U343 (N_343,In_15,In_252);
nor U344 (N_344,In_391,In_262);
nor U345 (N_345,In_31,In_482);
and U346 (N_346,In_269,In_83);
or U347 (N_347,In_93,In_14);
and U348 (N_348,In_231,In_357);
and U349 (N_349,In_21,In_305);
nor U350 (N_350,In_454,In_438);
nor U351 (N_351,In_44,In_73);
nor U352 (N_352,In_164,In_145);
nand U353 (N_353,In_160,In_270);
xor U354 (N_354,In_279,In_75);
or U355 (N_355,In_116,In_136);
xor U356 (N_356,In_146,In_28);
nor U357 (N_357,In_336,In_27);
nor U358 (N_358,In_264,In_255);
nor U359 (N_359,In_73,In_260);
nor U360 (N_360,In_447,In_112);
nand U361 (N_361,In_112,In_120);
nand U362 (N_362,In_153,In_99);
or U363 (N_363,In_114,In_335);
nand U364 (N_364,In_306,In_375);
or U365 (N_365,In_119,In_446);
nor U366 (N_366,In_440,In_56);
nand U367 (N_367,In_69,In_113);
nor U368 (N_368,In_284,In_410);
and U369 (N_369,In_389,In_164);
and U370 (N_370,In_475,In_354);
and U371 (N_371,In_445,In_126);
nand U372 (N_372,In_90,In_369);
nand U373 (N_373,In_225,In_409);
and U374 (N_374,In_93,In_143);
nand U375 (N_375,In_308,In_470);
xor U376 (N_376,In_27,In_91);
nor U377 (N_377,In_419,In_37);
or U378 (N_378,In_16,In_94);
nand U379 (N_379,In_96,In_248);
or U380 (N_380,In_65,In_358);
and U381 (N_381,In_475,In_40);
nand U382 (N_382,In_407,In_166);
nor U383 (N_383,In_98,In_225);
or U384 (N_384,In_409,In_48);
or U385 (N_385,In_19,In_74);
and U386 (N_386,In_301,In_378);
nor U387 (N_387,In_451,In_104);
nor U388 (N_388,In_486,In_408);
xnor U389 (N_389,In_6,In_197);
or U390 (N_390,In_162,In_295);
nor U391 (N_391,In_219,In_231);
nand U392 (N_392,In_299,In_10);
nor U393 (N_393,In_248,In_289);
nor U394 (N_394,In_58,In_176);
nand U395 (N_395,In_253,In_319);
nand U396 (N_396,In_493,In_24);
nand U397 (N_397,In_258,In_428);
nand U398 (N_398,In_62,In_466);
or U399 (N_399,In_37,In_184);
nor U400 (N_400,In_325,In_17);
xnor U401 (N_401,In_404,In_407);
nand U402 (N_402,In_439,In_365);
and U403 (N_403,In_396,In_118);
or U404 (N_404,In_176,In_118);
or U405 (N_405,In_209,In_414);
or U406 (N_406,In_33,In_116);
nand U407 (N_407,In_96,In_169);
nand U408 (N_408,In_47,In_389);
nor U409 (N_409,In_288,In_208);
nand U410 (N_410,In_21,In_487);
or U411 (N_411,In_195,In_137);
and U412 (N_412,In_217,In_192);
nand U413 (N_413,In_206,In_23);
nand U414 (N_414,In_439,In_210);
and U415 (N_415,In_99,In_55);
nor U416 (N_416,In_395,In_443);
and U417 (N_417,In_403,In_81);
nor U418 (N_418,In_357,In_174);
xnor U419 (N_419,In_54,In_284);
nor U420 (N_420,In_352,In_243);
xnor U421 (N_421,In_474,In_202);
xor U422 (N_422,In_99,In_225);
and U423 (N_423,In_29,In_57);
nand U424 (N_424,In_157,In_291);
nor U425 (N_425,In_167,In_242);
xor U426 (N_426,In_104,In_83);
or U427 (N_427,In_384,In_442);
nor U428 (N_428,In_4,In_1);
and U429 (N_429,In_192,In_263);
or U430 (N_430,In_392,In_432);
or U431 (N_431,In_240,In_297);
nand U432 (N_432,In_40,In_397);
and U433 (N_433,In_108,In_493);
and U434 (N_434,In_299,In_410);
nor U435 (N_435,In_283,In_59);
nor U436 (N_436,In_98,In_450);
nor U437 (N_437,In_414,In_39);
or U438 (N_438,In_478,In_184);
or U439 (N_439,In_257,In_371);
xnor U440 (N_440,In_212,In_260);
or U441 (N_441,In_59,In_133);
xnor U442 (N_442,In_318,In_131);
or U443 (N_443,In_78,In_42);
nand U444 (N_444,In_4,In_104);
or U445 (N_445,In_438,In_97);
or U446 (N_446,In_65,In_247);
nor U447 (N_447,In_403,In_397);
and U448 (N_448,In_76,In_210);
nor U449 (N_449,In_112,In_385);
or U450 (N_450,In_271,In_388);
nor U451 (N_451,In_165,In_66);
nor U452 (N_452,In_206,In_335);
and U453 (N_453,In_221,In_139);
and U454 (N_454,In_428,In_365);
or U455 (N_455,In_403,In_479);
or U456 (N_456,In_125,In_261);
nor U457 (N_457,In_304,In_132);
nor U458 (N_458,In_423,In_278);
or U459 (N_459,In_325,In_5);
xnor U460 (N_460,In_123,In_410);
and U461 (N_461,In_454,In_220);
nand U462 (N_462,In_42,In_445);
and U463 (N_463,In_264,In_471);
nand U464 (N_464,In_397,In_256);
xnor U465 (N_465,In_282,In_234);
xor U466 (N_466,In_279,In_349);
nor U467 (N_467,In_194,In_445);
or U468 (N_468,In_205,In_0);
xnor U469 (N_469,In_348,In_219);
and U470 (N_470,In_68,In_52);
or U471 (N_471,In_235,In_305);
or U472 (N_472,In_484,In_490);
and U473 (N_473,In_481,In_445);
nand U474 (N_474,In_445,In_113);
or U475 (N_475,In_129,In_489);
and U476 (N_476,In_468,In_46);
and U477 (N_477,In_28,In_322);
nand U478 (N_478,In_32,In_44);
nand U479 (N_479,In_222,In_98);
or U480 (N_480,In_231,In_316);
nand U481 (N_481,In_267,In_235);
nor U482 (N_482,In_248,In_29);
nand U483 (N_483,In_325,In_244);
nand U484 (N_484,In_474,In_44);
nor U485 (N_485,In_261,In_471);
nor U486 (N_486,In_388,In_121);
nor U487 (N_487,In_199,In_243);
nand U488 (N_488,In_290,In_464);
and U489 (N_489,In_176,In_171);
and U490 (N_490,In_371,In_208);
nor U491 (N_491,In_388,In_482);
or U492 (N_492,In_17,In_168);
or U493 (N_493,In_181,In_128);
and U494 (N_494,In_45,In_41);
nor U495 (N_495,In_125,In_373);
nor U496 (N_496,In_96,In_361);
nand U497 (N_497,In_403,In_62);
and U498 (N_498,In_424,In_394);
nor U499 (N_499,In_213,In_319);
nand U500 (N_500,In_359,In_173);
and U501 (N_501,In_497,In_8);
or U502 (N_502,In_423,In_196);
nand U503 (N_503,In_334,In_417);
and U504 (N_504,In_475,In_305);
nor U505 (N_505,In_53,In_275);
and U506 (N_506,In_354,In_118);
and U507 (N_507,In_491,In_60);
or U508 (N_508,In_7,In_175);
nand U509 (N_509,In_249,In_443);
xnor U510 (N_510,In_103,In_371);
and U511 (N_511,In_353,In_141);
and U512 (N_512,In_411,In_194);
nand U513 (N_513,In_177,In_490);
nor U514 (N_514,In_352,In_340);
xnor U515 (N_515,In_42,In_182);
nand U516 (N_516,In_122,In_382);
nand U517 (N_517,In_188,In_17);
and U518 (N_518,In_236,In_381);
and U519 (N_519,In_370,In_380);
xor U520 (N_520,In_422,In_126);
or U521 (N_521,In_406,In_304);
or U522 (N_522,In_69,In_459);
and U523 (N_523,In_78,In_43);
nand U524 (N_524,In_249,In_388);
and U525 (N_525,In_160,In_395);
or U526 (N_526,In_125,In_84);
xor U527 (N_527,In_70,In_358);
or U528 (N_528,In_294,In_8);
and U529 (N_529,In_480,In_495);
or U530 (N_530,In_122,In_92);
xnor U531 (N_531,In_121,In_470);
xnor U532 (N_532,In_31,In_121);
nor U533 (N_533,In_129,In_76);
nor U534 (N_534,In_450,In_348);
or U535 (N_535,In_349,In_301);
nor U536 (N_536,In_276,In_260);
nor U537 (N_537,In_346,In_498);
or U538 (N_538,In_207,In_168);
and U539 (N_539,In_131,In_469);
nor U540 (N_540,In_222,In_226);
or U541 (N_541,In_75,In_165);
or U542 (N_542,In_483,In_417);
xnor U543 (N_543,In_219,In_180);
and U544 (N_544,In_34,In_398);
nor U545 (N_545,In_152,In_451);
nor U546 (N_546,In_322,In_17);
nor U547 (N_547,In_374,In_150);
and U548 (N_548,In_275,In_377);
nand U549 (N_549,In_135,In_462);
or U550 (N_550,In_290,In_353);
and U551 (N_551,In_157,In_433);
nor U552 (N_552,In_386,In_470);
xnor U553 (N_553,In_290,In_328);
nand U554 (N_554,In_287,In_264);
or U555 (N_555,In_295,In_4);
or U556 (N_556,In_20,In_201);
nor U557 (N_557,In_190,In_497);
or U558 (N_558,In_354,In_206);
nand U559 (N_559,In_184,In_13);
or U560 (N_560,In_447,In_139);
nand U561 (N_561,In_236,In_447);
nor U562 (N_562,In_227,In_314);
or U563 (N_563,In_140,In_121);
nand U564 (N_564,In_179,In_494);
nor U565 (N_565,In_265,In_358);
xnor U566 (N_566,In_401,In_192);
and U567 (N_567,In_165,In_351);
and U568 (N_568,In_74,In_36);
nand U569 (N_569,In_451,In_74);
and U570 (N_570,In_109,In_246);
or U571 (N_571,In_339,In_242);
nor U572 (N_572,In_164,In_88);
or U573 (N_573,In_215,In_387);
nand U574 (N_574,In_15,In_306);
and U575 (N_575,In_383,In_431);
xnor U576 (N_576,In_189,In_87);
and U577 (N_577,In_238,In_54);
nand U578 (N_578,In_16,In_392);
or U579 (N_579,In_328,In_262);
nor U580 (N_580,In_94,In_63);
nor U581 (N_581,In_207,In_493);
and U582 (N_582,In_168,In_428);
nand U583 (N_583,In_331,In_329);
and U584 (N_584,In_472,In_226);
and U585 (N_585,In_393,In_411);
nor U586 (N_586,In_102,In_258);
and U587 (N_587,In_447,In_151);
or U588 (N_588,In_27,In_394);
nand U589 (N_589,In_465,In_192);
or U590 (N_590,In_243,In_67);
nor U591 (N_591,In_450,In_449);
and U592 (N_592,In_50,In_469);
nor U593 (N_593,In_386,In_413);
nor U594 (N_594,In_149,In_369);
nor U595 (N_595,In_488,In_87);
nor U596 (N_596,In_192,In_415);
nand U597 (N_597,In_41,In_397);
or U598 (N_598,In_109,In_293);
and U599 (N_599,In_13,In_84);
nor U600 (N_600,In_398,In_106);
or U601 (N_601,In_143,In_154);
and U602 (N_602,In_261,In_359);
nand U603 (N_603,In_106,In_52);
and U604 (N_604,In_463,In_360);
nand U605 (N_605,In_391,In_172);
or U606 (N_606,In_391,In_145);
and U607 (N_607,In_319,In_54);
xnor U608 (N_608,In_83,In_442);
and U609 (N_609,In_35,In_349);
nand U610 (N_610,In_173,In_258);
nand U611 (N_611,In_181,In_130);
and U612 (N_612,In_232,In_133);
nor U613 (N_613,In_287,In_426);
or U614 (N_614,In_173,In_336);
or U615 (N_615,In_367,In_302);
or U616 (N_616,In_274,In_2);
and U617 (N_617,In_129,In_467);
nor U618 (N_618,In_244,In_464);
and U619 (N_619,In_307,In_304);
or U620 (N_620,In_489,In_486);
nor U621 (N_621,In_1,In_86);
nand U622 (N_622,In_333,In_318);
xnor U623 (N_623,In_496,In_196);
or U624 (N_624,In_362,In_206);
or U625 (N_625,In_217,In_170);
and U626 (N_626,In_310,In_182);
nand U627 (N_627,In_44,In_404);
or U628 (N_628,In_445,In_280);
nor U629 (N_629,In_317,In_113);
and U630 (N_630,In_290,In_285);
and U631 (N_631,In_53,In_451);
or U632 (N_632,In_359,In_35);
or U633 (N_633,In_239,In_67);
or U634 (N_634,In_316,In_249);
nand U635 (N_635,In_270,In_239);
or U636 (N_636,In_220,In_398);
xor U637 (N_637,In_394,In_106);
xor U638 (N_638,In_54,In_341);
xnor U639 (N_639,In_199,In_197);
nand U640 (N_640,In_146,In_350);
and U641 (N_641,In_212,In_37);
nor U642 (N_642,In_211,In_173);
and U643 (N_643,In_380,In_13);
nor U644 (N_644,In_332,In_54);
nand U645 (N_645,In_75,In_92);
or U646 (N_646,In_242,In_361);
or U647 (N_647,In_405,In_378);
nor U648 (N_648,In_26,In_375);
and U649 (N_649,In_14,In_86);
and U650 (N_650,In_108,In_347);
nor U651 (N_651,In_167,In_215);
or U652 (N_652,In_140,In_442);
and U653 (N_653,In_148,In_365);
and U654 (N_654,In_223,In_55);
xnor U655 (N_655,In_43,In_94);
or U656 (N_656,In_405,In_47);
or U657 (N_657,In_35,In_312);
nand U658 (N_658,In_206,In_443);
and U659 (N_659,In_28,In_228);
xor U660 (N_660,In_363,In_46);
nor U661 (N_661,In_95,In_406);
nand U662 (N_662,In_482,In_21);
nor U663 (N_663,In_259,In_412);
nor U664 (N_664,In_429,In_197);
nand U665 (N_665,In_234,In_217);
nand U666 (N_666,In_161,In_357);
xnor U667 (N_667,In_226,In_356);
nand U668 (N_668,In_312,In_58);
or U669 (N_669,In_250,In_11);
or U670 (N_670,In_146,In_270);
or U671 (N_671,In_349,In_68);
nand U672 (N_672,In_55,In_27);
nor U673 (N_673,In_483,In_160);
nor U674 (N_674,In_131,In_34);
nand U675 (N_675,In_475,In_259);
or U676 (N_676,In_106,In_419);
nor U677 (N_677,In_414,In_296);
nand U678 (N_678,In_419,In_468);
nor U679 (N_679,In_57,In_316);
and U680 (N_680,In_206,In_471);
nor U681 (N_681,In_32,In_293);
nor U682 (N_682,In_436,In_207);
nor U683 (N_683,In_329,In_127);
nor U684 (N_684,In_131,In_298);
xnor U685 (N_685,In_437,In_167);
and U686 (N_686,In_40,In_214);
nand U687 (N_687,In_241,In_373);
or U688 (N_688,In_325,In_264);
nor U689 (N_689,In_451,In_239);
nand U690 (N_690,In_77,In_39);
nand U691 (N_691,In_398,In_244);
and U692 (N_692,In_191,In_151);
and U693 (N_693,In_483,In_485);
and U694 (N_694,In_39,In_395);
nand U695 (N_695,In_247,In_151);
and U696 (N_696,In_313,In_206);
or U697 (N_697,In_24,In_123);
or U698 (N_698,In_414,In_186);
nand U699 (N_699,In_167,In_488);
and U700 (N_700,In_431,In_224);
or U701 (N_701,In_419,In_165);
or U702 (N_702,In_153,In_366);
and U703 (N_703,In_202,In_448);
nand U704 (N_704,In_76,In_331);
and U705 (N_705,In_287,In_476);
and U706 (N_706,In_68,In_198);
and U707 (N_707,In_408,In_102);
and U708 (N_708,In_195,In_401);
or U709 (N_709,In_8,In_474);
or U710 (N_710,In_254,In_274);
and U711 (N_711,In_400,In_1);
nor U712 (N_712,In_443,In_167);
nand U713 (N_713,In_163,In_144);
nand U714 (N_714,In_498,In_371);
nand U715 (N_715,In_488,In_199);
nand U716 (N_716,In_430,In_449);
and U717 (N_717,In_128,In_235);
nand U718 (N_718,In_227,In_396);
nor U719 (N_719,In_263,In_496);
nand U720 (N_720,In_176,In_385);
nor U721 (N_721,In_180,In_126);
nand U722 (N_722,In_491,In_57);
nor U723 (N_723,In_62,In_474);
nand U724 (N_724,In_227,In_66);
nand U725 (N_725,In_99,In_453);
nor U726 (N_726,In_76,In_422);
nor U727 (N_727,In_431,In_442);
or U728 (N_728,In_132,In_74);
or U729 (N_729,In_370,In_19);
nand U730 (N_730,In_87,In_164);
xnor U731 (N_731,In_474,In_357);
or U732 (N_732,In_299,In_151);
and U733 (N_733,In_129,In_397);
or U734 (N_734,In_375,In_115);
and U735 (N_735,In_98,In_257);
nand U736 (N_736,In_345,In_204);
or U737 (N_737,In_238,In_152);
nor U738 (N_738,In_39,In_455);
nand U739 (N_739,In_184,In_59);
or U740 (N_740,In_236,In_422);
and U741 (N_741,In_168,In_215);
nor U742 (N_742,In_329,In_357);
and U743 (N_743,In_495,In_492);
nor U744 (N_744,In_161,In_447);
nand U745 (N_745,In_215,In_143);
nor U746 (N_746,In_169,In_306);
nand U747 (N_747,In_303,In_136);
nor U748 (N_748,In_391,In_105);
or U749 (N_749,In_82,In_324);
or U750 (N_750,In_321,In_340);
or U751 (N_751,In_296,In_424);
nor U752 (N_752,In_493,In_70);
or U753 (N_753,In_247,In_234);
nand U754 (N_754,In_199,In_291);
or U755 (N_755,In_104,In_249);
and U756 (N_756,In_382,In_217);
and U757 (N_757,In_81,In_10);
nand U758 (N_758,In_110,In_371);
xor U759 (N_759,In_167,In_346);
or U760 (N_760,In_379,In_10);
nand U761 (N_761,In_494,In_342);
nand U762 (N_762,In_412,In_110);
and U763 (N_763,In_298,In_188);
nor U764 (N_764,In_28,In_419);
nand U765 (N_765,In_193,In_321);
nor U766 (N_766,In_475,In_323);
xor U767 (N_767,In_94,In_245);
nand U768 (N_768,In_466,In_49);
nor U769 (N_769,In_448,In_46);
and U770 (N_770,In_14,In_98);
and U771 (N_771,In_61,In_106);
or U772 (N_772,In_347,In_232);
nand U773 (N_773,In_353,In_28);
nor U774 (N_774,In_64,In_193);
nor U775 (N_775,In_35,In_3);
nand U776 (N_776,In_452,In_379);
nor U777 (N_777,In_484,In_55);
and U778 (N_778,In_433,In_36);
nand U779 (N_779,In_132,In_282);
nand U780 (N_780,In_442,In_353);
xor U781 (N_781,In_27,In_470);
xor U782 (N_782,In_65,In_334);
nand U783 (N_783,In_385,In_417);
nor U784 (N_784,In_290,In_26);
nand U785 (N_785,In_163,In_214);
xnor U786 (N_786,In_188,In_92);
and U787 (N_787,In_290,In_61);
nand U788 (N_788,In_377,In_14);
and U789 (N_789,In_377,In_254);
and U790 (N_790,In_214,In_75);
or U791 (N_791,In_230,In_260);
nand U792 (N_792,In_351,In_274);
or U793 (N_793,In_177,In_212);
nand U794 (N_794,In_250,In_0);
nor U795 (N_795,In_311,In_64);
nand U796 (N_796,In_13,In_476);
xnor U797 (N_797,In_334,In_391);
nand U798 (N_798,In_303,In_102);
xnor U799 (N_799,In_272,In_233);
nor U800 (N_800,In_264,In_132);
nor U801 (N_801,In_253,In_165);
nand U802 (N_802,In_250,In_322);
nor U803 (N_803,In_256,In_174);
nor U804 (N_804,In_9,In_19);
nand U805 (N_805,In_290,In_146);
nand U806 (N_806,In_200,In_319);
and U807 (N_807,In_446,In_377);
nor U808 (N_808,In_62,In_476);
nor U809 (N_809,In_170,In_487);
xnor U810 (N_810,In_209,In_112);
nor U811 (N_811,In_167,In_251);
nor U812 (N_812,In_37,In_205);
xnor U813 (N_813,In_160,In_377);
or U814 (N_814,In_168,In_82);
nand U815 (N_815,In_184,In_1);
and U816 (N_816,In_452,In_153);
and U817 (N_817,In_153,In_274);
or U818 (N_818,In_453,In_292);
and U819 (N_819,In_74,In_359);
or U820 (N_820,In_468,In_61);
nand U821 (N_821,In_435,In_402);
nand U822 (N_822,In_489,In_49);
and U823 (N_823,In_143,In_83);
xnor U824 (N_824,In_106,In_265);
xor U825 (N_825,In_36,In_10);
or U826 (N_826,In_214,In_367);
xnor U827 (N_827,In_180,In_203);
nor U828 (N_828,In_322,In_90);
or U829 (N_829,In_88,In_153);
or U830 (N_830,In_233,In_198);
or U831 (N_831,In_1,In_217);
and U832 (N_832,In_401,In_323);
and U833 (N_833,In_354,In_236);
nor U834 (N_834,In_94,In_498);
and U835 (N_835,In_10,In_5);
nand U836 (N_836,In_486,In_165);
or U837 (N_837,In_22,In_382);
or U838 (N_838,In_270,In_195);
nand U839 (N_839,In_425,In_428);
and U840 (N_840,In_45,In_320);
nand U841 (N_841,In_361,In_459);
and U842 (N_842,In_370,In_373);
nand U843 (N_843,In_299,In_478);
nor U844 (N_844,In_305,In_285);
and U845 (N_845,In_363,In_132);
and U846 (N_846,In_118,In_382);
nand U847 (N_847,In_379,In_199);
xnor U848 (N_848,In_268,In_198);
and U849 (N_849,In_244,In_212);
nor U850 (N_850,In_358,In_156);
nor U851 (N_851,In_340,In_164);
or U852 (N_852,In_144,In_373);
nand U853 (N_853,In_200,In_166);
or U854 (N_854,In_314,In_311);
nand U855 (N_855,In_207,In_157);
xor U856 (N_856,In_180,In_198);
nand U857 (N_857,In_261,In_5);
nor U858 (N_858,In_166,In_198);
or U859 (N_859,In_378,In_388);
nand U860 (N_860,In_385,In_57);
or U861 (N_861,In_420,In_437);
and U862 (N_862,In_93,In_192);
or U863 (N_863,In_295,In_411);
nand U864 (N_864,In_446,In_189);
and U865 (N_865,In_363,In_183);
or U866 (N_866,In_401,In_313);
or U867 (N_867,In_222,In_333);
and U868 (N_868,In_142,In_281);
nand U869 (N_869,In_64,In_0);
or U870 (N_870,In_173,In_203);
nand U871 (N_871,In_380,In_304);
or U872 (N_872,In_341,In_324);
and U873 (N_873,In_13,In_447);
nor U874 (N_874,In_113,In_471);
and U875 (N_875,In_398,In_237);
or U876 (N_876,In_11,In_99);
or U877 (N_877,In_0,In_318);
or U878 (N_878,In_421,In_239);
and U879 (N_879,In_27,In_254);
and U880 (N_880,In_437,In_52);
and U881 (N_881,In_10,In_202);
xnor U882 (N_882,In_297,In_365);
or U883 (N_883,In_384,In_328);
and U884 (N_884,In_73,In_189);
or U885 (N_885,In_203,In_198);
nor U886 (N_886,In_486,In_244);
and U887 (N_887,In_73,In_464);
and U888 (N_888,In_403,In_343);
xor U889 (N_889,In_91,In_54);
nor U890 (N_890,In_422,In_190);
and U891 (N_891,In_270,In_159);
nand U892 (N_892,In_434,In_78);
or U893 (N_893,In_109,In_480);
nand U894 (N_894,In_17,In_31);
and U895 (N_895,In_140,In_34);
or U896 (N_896,In_259,In_88);
or U897 (N_897,In_375,In_385);
and U898 (N_898,In_343,In_24);
nor U899 (N_899,In_437,In_67);
nand U900 (N_900,In_385,In_197);
nor U901 (N_901,In_148,In_404);
nand U902 (N_902,In_123,In_300);
nor U903 (N_903,In_287,In_149);
or U904 (N_904,In_195,In_330);
or U905 (N_905,In_267,In_35);
nor U906 (N_906,In_328,In_12);
and U907 (N_907,In_256,In_29);
and U908 (N_908,In_287,In_141);
nand U909 (N_909,In_337,In_95);
nand U910 (N_910,In_127,In_259);
nor U911 (N_911,In_213,In_146);
or U912 (N_912,In_187,In_268);
nand U913 (N_913,In_352,In_407);
xnor U914 (N_914,In_436,In_39);
xnor U915 (N_915,In_282,In_299);
nor U916 (N_916,In_182,In_327);
nor U917 (N_917,In_83,In_376);
xor U918 (N_918,In_372,In_21);
xor U919 (N_919,In_126,In_361);
nor U920 (N_920,In_471,In_482);
or U921 (N_921,In_167,In_382);
and U922 (N_922,In_52,In_300);
or U923 (N_923,In_486,In_50);
or U924 (N_924,In_99,In_232);
and U925 (N_925,In_440,In_383);
and U926 (N_926,In_137,In_369);
xnor U927 (N_927,In_460,In_383);
or U928 (N_928,In_237,In_156);
nor U929 (N_929,In_114,In_317);
nand U930 (N_930,In_233,In_387);
xor U931 (N_931,In_378,In_478);
or U932 (N_932,In_396,In_164);
or U933 (N_933,In_6,In_165);
nor U934 (N_934,In_8,In_464);
nor U935 (N_935,In_237,In_456);
and U936 (N_936,In_302,In_384);
or U937 (N_937,In_63,In_111);
xnor U938 (N_938,In_190,In_8);
nor U939 (N_939,In_28,In_470);
and U940 (N_940,In_11,In_284);
or U941 (N_941,In_411,In_492);
nand U942 (N_942,In_456,In_346);
and U943 (N_943,In_31,In_249);
nand U944 (N_944,In_395,In_154);
nor U945 (N_945,In_218,In_499);
xor U946 (N_946,In_417,In_327);
and U947 (N_947,In_212,In_158);
nand U948 (N_948,In_236,In_6);
xnor U949 (N_949,In_22,In_306);
or U950 (N_950,In_474,In_74);
or U951 (N_951,In_51,In_259);
nand U952 (N_952,In_409,In_305);
and U953 (N_953,In_29,In_499);
nor U954 (N_954,In_296,In_401);
xnor U955 (N_955,In_394,In_324);
nor U956 (N_956,In_438,In_330);
and U957 (N_957,In_258,In_228);
or U958 (N_958,In_466,In_120);
nand U959 (N_959,In_174,In_72);
and U960 (N_960,In_499,In_339);
xor U961 (N_961,In_28,In_384);
xor U962 (N_962,In_46,In_302);
or U963 (N_963,In_471,In_281);
or U964 (N_964,In_176,In_322);
and U965 (N_965,In_71,In_289);
or U966 (N_966,In_451,In_169);
or U967 (N_967,In_458,In_254);
nor U968 (N_968,In_337,In_346);
nand U969 (N_969,In_290,In_253);
or U970 (N_970,In_109,In_470);
nand U971 (N_971,In_371,In_276);
nand U972 (N_972,In_115,In_232);
or U973 (N_973,In_49,In_479);
nand U974 (N_974,In_403,In_171);
xor U975 (N_975,In_202,In_213);
nand U976 (N_976,In_303,In_351);
and U977 (N_977,In_441,In_439);
and U978 (N_978,In_418,In_260);
nor U979 (N_979,In_114,In_332);
or U980 (N_980,In_136,In_275);
nand U981 (N_981,In_4,In_106);
nand U982 (N_982,In_108,In_128);
nor U983 (N_983,In_490,In_157);
nor U984 (N_984,In_176,In_456);
and U985 (N_985,In_328,In_489);
nand U986 (N_986,In_56,In_256);
or U987 (N_987,In_54,In_49);
and U988 (N_988,In_174,In_350);
nor U989 (N_989,In_140,In_491);
or U990 (N_990,In_201,In_414);
xor U991 (N_991,In_322,In_432);
or U992 (N_992,In_200,In_70);
and U993 (N_993,In_168,In_263);
or U994 (N_994,In_314,In_59);
nor U995 (N_995,In_419,In_342);
and U996 (N_996,In_496,In_50);
and U997 (N_997,In_330,In_241);
and U998 (N_998,In_393,In_327);
nor U999 (N_999,In_36,In_429);
or U1000 (N_1000,N_222,N_914);
nor U1001 (N_1001,N_471,N_332);
or U1002 (N_1002,N_391,N_630);
or U1003 (N_1003,N_447,N_791);
xor U1004 (N_1004,N_955,N_572);
or U1005 (N_1005,N_740,N_498);
and U1006 (N_1006,N_592,N_629);
nor U1007 (N_1007,N_164,N_892);
nand U1008 (N_1008,N_602,N_472);
nand U1009 (N_1009,N_850,N_453);
nand U1010 (N_1010,N_198,N_81);
nor U1011 (N_1011,N_963,N_623);
nor U1012 (N_1012,N_474,N_321);
or U1013 (N_1013,N_751,N_839);
nor U1014 (N_1014,N_542,N_191);
nor U1015 (N_1015,N_460,N_253);
and U1016 (N_1016,N_678,N_399);
nor U1017 (N_1017,N_152,N_481);
and U1018 (N_1018,N_544,N_918);
nand U1019 (N_1019,N_965,N_350);
or U1020 (N_1020,N_113,N_41);
and U1021 (N_1021,N_288,N_652);
or U1022 (N_1022,N_414,N_229);
nand U1023 (N_1023,N_256,N_353);
and U1024 (N_1024,N_318,N_380);
or U1025 (N_1025,N_431,N_564);
nor U1026 (N_1026,N_181,N_452);
nor U1027 (N_1027,N_195,N_501);
and U1028 (N_1028,N_371,N_557);
nor U1029 (N_1029,N_618,N_190);
nor U1030 (N_1030,N_84,N_508);
nand U1031 (N_1031,N_593,N_323);
or U1032 (N_1032,N_856,N_283);
and U1033 (N_1033,N_880,N_891);
nand U1034 (N_1034,N_754,N_272);
nand U1035 (N_1035,N_582,N_274);
and U1036 (N_1036,N_598,N_275);
nor U1037 (N_1037,N_732,N_684);
nand U1038 (N_1038,N_107,N_70);
nor U1039 (N_1039,N_999,N_889);
nor U1040 (N_1040,N_178,N_349);
nor U1041 (N_1041,N_520,N_364);
nor U1042 (N_1042,N_951,N_549);
and U1043 (N_1043,N_369,N_642);
nand U1044 (N_1044,N_725,N_376);
xnor U1045 (N_1045,N_745,N_146);
nor U1046 (N_1046,N_182,N_527);
nand U1047 (N_1047,N_314,N_674);
nand U1048 (N_1048,N_217,N_424);
or U1049 (N_1049,N_798,N_329);
or U1050 (N_1050,N_579,N_224);
or U1051 (N_1051,N_241,N_931);
xnor U1052 (N_1052,N_915,N_874);
nor U1053 (N_1053,N_654,N_834);
nor U1054 (N_1054,N_586,N_752);
and U1055 (N_1055,N_422,N_112);
nand U1056 (N_1056,N_469,N_552);
xnor U1057 (N_1057,N_741,N_722);
or U1058 (N_1058,N_671,N_902);
or U1059 (N_1059,N_865,N_616);
or U1060 (N_1060,N_404,N_805);
nand U1061 (N_1061,N_971,N_800);
and U1062 (N_1062,N_55,N_277);
xnor U1063 (N_1063,N_120,N_123);
nand U1064 (N_1064,N_867,N_777);
xor U1065 (N_1065,N_773,N_137);
or U1066 (N_1066,N_615,N_637);
and U1067 (N_1067,N_263,N_382);
nand U1068 (N_1068,N_554,N_820);
and U1069 (N_1069,N_851,N_799);
or U1070 (N_1070,N_907,N_957);
or U1071 (N_1071,N_34,N_3);
nor U1072 (N_1072,N_410,N_646);
nor U1073 (N_1073,N_682,N_324);
nor U1074 (N_1074,N_973,N_655);
nand U1075 (N_1075,N_911,N_157);
nor U1076 (N_1076,N_220,N_534);
nor U1077 (N_1077,N_597,N_522);
xor U1078 (N_1078,N_609,N_286);
nand U1079 (N_1079,N_875,N_545);
nor U1080 (N_1080,N_644,N_90);
xor U1081 (N_1081,N_374,N_31);
nand U1082 (N_1082,N_988,N_306);
nand U1083 (N_1083,N_265,N_292);
or U1084 (N_1084,N_499,N_871);
and U1085 (N_1085,N_894,N_475);
and U1086 (N_1086,N_733,N_479);
and U1087 (N_1087,N_276,N_882);
nand U1088 (N_1088,N_864,N_86);
or U1089 (N_1089,N_994,N_67);
or U1090 (N_1090,N_862,N_964);
nor U1091 (N_1091,N_131,N_574);
nand U1092 (N_1092,N_816,N_702);
nor U1093 (N_1093,N_521,N_199);
nand U1094 (N_1094,N_138,N_419);
or U1095 (N_1095,N_956,N_437);
or U1096 (N_1096,N_402,N_885);
nand U1097 (N_1097,N_877,N_600);
and U1098 (N_1098,N_908,N_38);
nor U1099 (N_1099,N_692,N_640);
nand U1100 (N_1100,N_689,N_954);
or U1101 (N_1101,N_819,N_54);
and U1102 (N_1102,N_328,N_16);
nor U1103 (N_1103,N_480,N_768);
xor U1104 (N_1104,N_942,N_992);
xnor U1105 (N_1105,N_569,N_47);
or U1106 (N_1106,N_920,N_72);
xnor U1107 (N_1107,N_79,N_327);
or U1108 (N_1108,N_727,N_494);
nor U1109 (N_1109,N_632,N_270);
nand U1110 (N_1110,N_359,N_929);
nor U1111 (N_1111,N_581,N_518);
nor U1112 (N_1112,N_928,N_770);
and U1113 (N_1113,N_700,N_483);
or U1114 (N_1114,N_363,N_121);
xnor U1115 (N_1115,N_724,N_78);
nor U1116 (N_1116,N_168,N_715);
and U1117 (N_1117,N_662,N_886);
or U1118 (N_1118,N_192,N_30);
nor U1119 (N_1119,N_861,N_901);
or U1120 (N_1120,N_663,N_571);
nor U1121 (N_1121,N_633,N_857);
nand U1122 (N_1122,N_686,N_691);
nand U1123 (N_1123,N_560,N_831);
and U1124 (N_1124,N_604,N_977);
nand U1125 (N_1125,N_185,N_106);
nand U1126 (N_1126,N_218,N_507);
or U1127 (N_1127,N_559,N_526);
and U1128 (N_1128,N_311,N_599);
or U1129 (N_1129,N_243,N_665);
and U1130 (N_1130,N_114,N_340);
or U1131 (N_1131,N_242,N_337);
nor U1132 (N_1132,N_24,N_673);
and U1133 (N_1133,N_550,N_258);
nand U1134 (N_1134,N_840,N_523);
xor U1135 (N_1135,N_667,N_925);
nor U1136 (N_1136,N_32,N_688);
nand U1137 (N_1137,N_9,N_394);
and U1138 (N_1138,N_147,N_111);
and U1139 (N_1139,N_813,N_748);
or U1140 (N_1140,N_291,N_981);
nor U1141 (N_1141,N_228,N_470);
and U1142 (N_1142,N_653,N_10);
and U1143 (N_1143,N_279,N_505);
xnor U1144 (N_1144,N_130,N_492);
and U1145 (N_1145,N_860,N_325);
or U1146 (N_1146,N_305,N_177);
nor U1147 (N_1147,N_513,N_75);
and U1148 (N_1148,N_295,N_624);
or U1149 (N_1149,N_742,N_436);
nand U1150 (N_1150,N_514,N_893);
and U1151 (N_1151,N_246,N_695);
nand U1152 (N_1152,N_149,N_659);
nor U1153 (N_1153,N_440,N_836);
xnor U1154 (N_1154,N_393,N_685);
nor U1155 (N_1155,N_679,N_583);
nor U1156 (N_1156,N_83,N_225);
and U1157 (N_1157,N_917,N_390);
and U1158 (N_1158,N_968,N_676);
nor U1159 (N_1159,N_187,N_763);
or U1160 (N_1160,N_535,N_771);
nand U1161 (N_1161,N_236,N_338);
nor U1162 (N_1162,N_260,N_20);
nand U1163 (N_1163,N_196,N_797);
or U1164 (N_1164,N_783,N_859);
or U1165 (N_1165,N_669,N_807);
nand U1166 (N_1166,N_442,N_997);
or U1167 (N_1167,N_995,N_619);
and U1168 (N_1168,N_897,N_80);
or U1169 (N_1169,N_144,N_345);
or U1170 (N_1170,N_284,N_823);
nor U1171 (N_1171,N_815,N_405);
nor U1172 (N_1172,N_612,N_262);
nand U1173 (N_1173,N_814,N_308);
nor U1174 (N_1174,N_728,N_556);
xor U1175 (N_1175,N_720,N_884);
nand U1176 (N_1176,N_99,N_100);
and U1177 (N_1177,N_870,N_211);
nor U1178 (N_1178,N_53,N_497);
and U1179 (N_1179,N_959,N_140);
xnor U1180 (N_1180,N_767,N_822);
nor U1181 (N_1181,N_153,N_213);
nor U1182 (N_1182,N_517,N_301);
nor U1183 (N_1183,N_361,N_387);
nor U1184 (N_1184,N_268,N_764);
xnor U1185 (N_1185,N_351,N_575);
or U1186 (N_1186,N_916,N_869);
or U1187 (N_1187,N_945,N_628);
nand U1188 (N_1188,N_457,N_432);
and U1189 (N_1189,N_577,N_122);
nor U1190 (N_1190,N_761,N_296);
xor U1191 (N_1191,N_943,N_162);
and U1192 (N_1192,N_25,N_209);
nor U1193 (N_1193,N_386,N_919);
nand U1194 (N_1194,N_334,N_142);
and U1195 (N_1195,N_488,N_40);
or U1196 (N_1196,N_879,N_802);
nor U1197 (N_1197,N_753,N_610);
nand U1198 (N_1198,N_806,N_844);
nor U1199 (N_1199,N_37,N_743);
or U1200 (N_1200,N_546,N_650);
nor U1201 (N_1201,N_124,N_461);
nand U1202 (N_1202,N_565,N_289);
and U1203 (N_1203,N_530,N_750);
and U1204 (N_1204,N_48,N_626);
or U1205 (N_1205,N_8,N_22);
nor U1206 (N_1206,N_717,N_467);
nor U1207 (N_1207,N_948,N_677);
nand U1208 (N_1208,N_249,N_709);
nor U1209 (N_1209,N_409,N_317);
or U1210 (N_1210,N_825,N_881);
nor U1211 (N_1211,N_352,N_56);
nand U1212 (N_1212,N_448,N_976);
and U1213 (N_1213,N_921,N_952);
nor U1214 (N_1214,N_758,N_439);
or U1215 (N_1215,N_366,N_400);
nor U1216 (N_1216,N_937,N_412);
or U1217 (N_1217,N_341,N_990);
nand U1218 (N_1218,N_833,N_699);
or U1219 (N_1219,N_536,N_852);
or U1220 (N_1220,N_215,N_487);
and U1221 (N_1221,N_736,N_547);
nand U1222 (N_1222,N_233,N_322);
and U1223 (N_1223,N_312,N_6);
or U1224 (N_1224,N_372,N_622);
and U1225 (N_1225,N_335,N_273);
nor U1226 (N_1226,N_775,N_969);
nand U1227 (N_1227,N_485,N_941);
or U1228 (N_1228,N_239,N_45);
or U1229 (N_1229,N_74,N_656);
nor U1230 (N_1230,N_232,N_214);
or U1231 (N_1231,N_670,N_811);
or U1232 (N_1232,N_810,N_331);
nand U1233 (N_1233,N_502,N_596);
nor U1234 (N_1234,N_985,N_780);
and U1235 (N_1235,N_119,N_944);
or U1236 (N_1236,N_878,N_219);
or U1237 (N_1237,N_7,N_934);
and U1238 (N_1238,N_647,N_804);
nand U1239 (N_1239,N_978,N_202);
xor U1240 (N_1240,N_693,N_760);
nor U1241 (N_1241,N_384,N_365);
nand U1242 (N_1242,N_139,N_853);
and U1243 (N_1243,N_385,N_108);
nor U1244 (N_1244,N_420,N_61);
nor U1245 (N_1245,N_316,N_991);
nor U1246 (N_1246,N_343,N_562);
or U1247 (N_1247,N_890,N_675);
or U1248 (N_1248,N_357,N_208);
nand U1249 (N_1249,N_135,N_169);
nor U1250 (N_1250,N_872,N_533);
or U1251 (N_1251,N_666,N_660);
and U1252 (N_1252,N_772,N_484);
nand U1253 (N_1253,N_779,N_608);
nor U1254 (N_1254,N_982,N_319);
xnor U1255 (N_1255,N_972,N_762);
nand U1256 (N_1256,N_94,N_417);
xor U1257 (N_1257,N_326,N_636);
xnor U1258 (N_1258,N_787,N_854);
nor U1259 (N_1259,N_605,N_425);
nand U1260 (N_1260,N_873,N_735);
nand U1261 (N_1261,N_39,N_519);
nor U1262 (N_1262,N_290,N_996);
or U1263 (N_1263,N_620,N_809);
and U1264 (N_1264,N_903,N_817);
and U1265 (N_1265,N_355,N_221);
nand U1266 (N_1266,N_818,N_35);
nand U1267 (N_1267,N_132,N_93);
nor U1268 (N_1268,N_843,N_254);
or U1269 (N_1269,N_790,N_532);
nor U1270 (N_1270,N_749,N_466);
and U1271 (N_1271,N_658,N_287);
or U1272 (N_1272,N_540,N_993);
xor U1273 (N_1273,N_478,N_570);
nor U1274 (N_1274,N_173,N_826);
and U1275 (N_1275,N_418,N_52);
nor U1276 (N_1276,N_15,N_423);
or U1277 (N_1277,N_82,N_416);
and U1278 (N_1278,N_381,N_237);
nand U1279 (N_1279,N_12,N_63);
nand U1280 (N_1280,N_201,N_847);
nand U1281 (N_1281,N_774,N_989);
or U1282 (N_1282,N_176,N_2);
and U1283 (N_1283,N_701,N_59);
nand U1284 (N_1284,N_297,N_465);
or U1285 (N_1285,N_883,N_657);
xor U1286 (N_1286,N_697,N_960);
xor U1287 (N_1287,N_984,N_808);
xor U1288 (N_1288,N_525,N_607);
nor U1289 (N_1289,N_866,N_346);
or U1290 (N_1290,N_495,N_68);
xnor U1291 (N_1291,N_543,N_888);
nor U1292 (N_1292,N_179,N_784);
and U1293 (N_1293,N_643,N_603);
or U1294 (N_1294,N_348,N_585);
or U1295 (N_1295,N_486,N_189);
nand U1296 (N_1296,N_887,N_463);
or U1297 (N_1297,N_266,N_28);
and U1298 (N_1298,N_141,N_129);
nand U1299 (N_1299,N_298,N_974);
xnor U1300 (N_1300,N_240,N_5);
nor U1301 (N_1301,N_193,N_50);
and U1302 (N_1302,N_812,N_115);
nand U1303 (N_1303,N_489,N_967);
nor U1304 (N_1304,N_395,N_117);
nor U1305 (N_1305,N_60,N_573);
and U1306 (N_1306,N_389,N_595);
and U1307 (N_1307,N_46,N_958);
nand U1308 (N_1308,N_759,N_27);
or U1309 (N_1309,N_85,N_718);
or U1310 (N_1310,N_19,N_230);
or U1311 (N_1311,N_634,N_313);
xor U1312 (N_1312,N_49,N_975);
nand U1313 (N_1313,N_356,N_648);
nor U1314 (N_1314,N_726,N_795);
xor U1315 (N_1315,N_17,N_868);
and U1316 (N_1316,N_264,N_408);
xor U1317 (N_1317,N_576,N_428);
or U1318 (N_1318,N_77,N_373);
and U1319 (N_1319,N_69,N_370);
and U1320 (N_1320,N_294,N_962);
nor U1321 (N_1321,N_88,N_744);
xor U1322 (N_1322,N_101,N_938);
and U1323 (N_1323,N_635,N_704);
and U1324 (N_1324,N_829,N_785);
and U1325 (N_1325,N_690,N_250);
or U1326 (N_1326,N_302,N_11);
nor U1327 (N_1327,N_738,N_438);
xor U1328 (N_1328,N_427,N_589);
and U1329 (N_1329,N_392,N_133);
or U1330 (N_1330,N_776,N_21);
nor U1331 (N_1331,N_299,N_649);
nor U1332 (N_1332,N_450,N_231);
nand U1333 (N_1333,N_936,N_252);
and U1334 (N_1334,N_788,N_13);
or U1335 (N_1335,N_449,N_842);
xor U1336 (N_1336,N_568,N_567);
xor U1337 (N_1337,N_515,N_983);
xnor U1338 (N_1338,N_110,N_134);
xnor U1339 (N_1339,N_148,N_281);
nor U1340 (N_1340,N_234,N_280);
xnor U1341 (N_1341,N_163,N_42);
or U1342 (N_1342,N_824,N_269);
xor U1343 (N_1343,N_65,N_307);
or U1344 (N_1344,N_226,N_551);
nor U1345 (N_1345,N_606,N_707);
nand U1346 (N_1346,N_97,N_161);
nand U1347 (N_1347,N_832,N_126);
nor U1348 (N_1348,N_339,N_703);
and U1349 (N_1349,N_285,N_92);
nor U1350 (N_1350,N_212,N_443);
nand U1351 (N_1351,N_746,N_383);
nor U1352 (N_1352,N_613,N_933);
nand U1353 (N_1353,N_561,N_998);
or U1354 (N_1354,N_278,N_468);
nand U1355 (N_1355,N_109,N_203);
and U1356 (N_1356,N_358,N_939);
or U1357 (N_1357,N_714,N_651);
and U1358 (N_1358,N_713,N_698);
and U1359 (N_1359,N_104,N_792);
xor U1360 (N_1360,N_304,N_627);
or U1361 (N_1361,N_444,N_512);
and U1362 (N_1362,N_445,N_333);
xnor U1363 (N_1363,N_730,N_172);
nor U1364 (N_1364,N_858,N_433);
and U1365 (N_1365,N_838,N_464);
nand U1366 (N_1366,N_26,N_757);
nand U1367 (N_1367,N_159,N_946);
and U1368 (N_1368,N_504,N_765);
and U1369 (N_1369,N_524,N_789);
nor U1370 (N_1370,N_227,N_830);
nand U1371 (N_1371,N_491,N_127);
or U1372 (N_1372,N_1,N_206);
nor U1373 (N_1373,N_493,N_922);
nor U1374 (N_1374,N_828,N_267);
nor U1375 (N_1375,N_434,N_553);
nor U1376 (N_1376,N_455,N_731);
or U1377 (N_1377,N_406,N_155);
or U1378 (N_1378,N_128,N_330);
and U1379 (N_1379,N_71,N_261);
nand U1380 (N_1380,N_315,N_841);
nand U1381 (N_1381,N_247,N_446);
nand U1382 (N_1382,N_638,N_528);
nor U1383 (N_1383,N_377,N_706);
and U1384 (N_1384,N_103,N_245);
xnor U1385 (N_1385,N_477,N_490);
nor U1386 (N_1386,N_541,N_496);
nor U1387 (N_1387,N_906,N_723);
nor U1388 (N_1388,N_855,N_183);
nor U1389 (N_1389,N_300,N_205);
nor U1390 (N_1390,N_360,N_687);
nand U1391 (N_1391,N_905,N_578);
nor U1392 (N_1392,N_537,N_158);
and U1393 (N_1393,N_257,N_14);
or U1394 (N_1394,N_721,N_244);
or U1395 (N_1395,N_849,N_186);
or U1396 (N_1396,N_711,N_584);
nand U1397 (N_1397,N_899,N_398);
nor U1398 (N_1398,N_368,N_150);
nor U1399 (N_1399,N_451,N_621);
or U1400 (N_1400,N_781,N_166);
and U1401 (N_1401,N_803,N_712);
and U1402 (N_1402,N_342,N_238);
nand U1403 (N_1403,N_454,N_57);
xor U1404 (N_1404,N_716,N_835);
and U1405 (N_1405,N_910,N_441);
nor U1406 (N_1406,N_167,N_156);
or U1407 (N_1407,N_846,N_548);
or U1408 (N_1408,N_793,N_683);
nand U1409 (N_1409,N_476,N_309);
or U1410 (N_1410,N_89,N_43);
and U1411 (N_1411,N_429,N_953);
nor U1412 (N_1412,N_734,N_170);
and U1413 (N_1413,N_930,N_558);
or U1414 (N_1414,N_986,N_590);
xor U1415 (N_1415,N_909,N_375);
or U1416 (N_1416,N_29,N_200);
nand U1417 (N_1417,N_614,N_64);
or U1418 (N_1418,N_563,N_413);
nand U1419 (N_1419,N_566,N_303);
nand U1420 (N_1420,N_347,N_271);
nor U1421 (N_1421,N_210,N_435);
nand U1422 (N_1422,N_407,N_979);
or U1423 (N_1423,N_344,N_207);
and U1424 (N_1424,N_255,N_91);
nor U1425 (N_1425,N_511,N_970);
and U1426 (N_1426,N_645,N_354);
nor U1427 (N_1427,N_966,N_539);
nand U1428 (N_1428,N_672,N_459);
nand U1429 (N_1429,N_848,N_516);
and U1430 (N_1430,N_18,N_248);
nand U1431 (N_1431,N_949,N_950);
and U1432 (N_1432,N_204,N_194);
and U1433 (N_1433,N_932,N_591);
and U1434 (N_1434,N_786,N_118);
and U1435 (N_1435,N_611,N_506);
nor U1436 (N_1436,N_411,N_415);
nor U1437 (N_1437,N_136,N_62);
or U1438 (N_1438,N_473,N_367);
nand U1439 (N_1439,N_500,N_580);
nand U1440 (N_1440,N_151,N_503);
nand U1441 (N_1441,N_924,N_293);
xor U1442 (N_1442,N_73,N_729);
and U1443 (N_1443,N_125,N_36);
and U1444 (N_1444,N_895,N_766);
or U1445 (N_1445,N_947,N_96);
nand U1446 (N_1446,N_755,N_175);
or U1447 (N_1447,N_641,N_782);
and U1448 (N_1448,N_223,N_778);
and U1449 (N_1449,N_664,N_796);
nand U1450 (N_1450,N_320,N_961);
and U1451 (N_1451,N_509,N_631);
and U1452 (N_1452,N_251,N_756);
nor U1453 (N_1453,N_719,N_827);
nand U1454 (N_1454,N_336,N_681);
nand U1455 (N_1455,N_362,N_747);
nand U1456 (N_1456,N_594,N_876);
nor U1457 (N_1457,N_76,N_980);
nor U1458 (N_1458,N_379,N_143);
nand U1459 (N_1459,N_33,N_310);
nor U1460 (N_1460,N_4,N_388);
nor U1461 (N_1461,N_531,N_456);
or U1462 (N_1462,N_896,N_529);
and U1463 (N_1463,N_601,N_188);
and U1464 (N_1464,N_900,N_680);
or U1465 (N_1465,N_160,N_259);
nor U1466 (N_1466,N_462,N_180);
nor U1467 (N_1467,N_184,N_739);
or U1468 (N_1468,N_105,N_661);
nor U1469 (N_1469,N_116,N_987);
nand U1470 (N_1470,N_705,N_174);
nor U1471 (N_1471,N_801,N_913);
or U1472 (N_1472,N_694,N_396);
and U1473 (N_1473,N_397,N_87);
and U1474 (N_1474,N_912,N_23);
or U1475 (N_1475,N_66,N_458);
nor U1476 (N_1476,N_538,N_98);
nand U1477 (N_1477,N_165,N_837);
and U1478 (N_1478,N_625,N_421);
nand U1479 (N_1479,N_426,N_696);
nand U1480 (N_1480,N_145,N_668);
or U1481 (N_1481,N_794,N_401);
and U1482 (N_1482,N_940,N_588);
or U1483 (N_1483,N_935,N_51);
nor U1484 (N_1484,N_0,N_926);
nor U1485 (N_1485,N_510,N_708);
and U1486 (N_1486,N_95,N_154);
and U1487 (N_1487,N_737,N_197);
or U1488 (N_1488,N_430,N_403);
nor U1489 (N_1489,N_235,N_482);
nand U1490 (N_1490,N_845,N_587);
nand U1491 (N_1491,N_769,N_923);
nor U1492 (N_1492,N_639,N_898);
nor U1493 (N_1493,N_58,N_617);
nor U1494 (N_1494,N_378,N_171);
or U1495 (N_1495,N_216,N_102);
or U1496 (N_1496,N_821,N_555);
nor U1497 (N_1497,N_863,N_710);
xor U1498 (N_1498,N_927,N_904);
xor U1499 (N_1499,N_282,N_44);
nand U1500 (N_1500,N_399,N_395);
and U1501 (N_1501,N_885,N_757);
and U1502 (N_1502,N_519,N_114);
nor U1503 (N_1503,N_817,N_220);
nor U1504 (N_1504,N_370,N_360);
nand U1505 (N_1505,N_56,N_747);
and U1506 (N_1506,N_144,N_101);
and U1507 (N_1507,N_439,N_435);
nand U1508 (N_1508,N_407,N_246);
nand U1509 (N_1509,N_627,N_886);
nand U1510 (N_1510,N_77,N_154);
xnor U1511 (N_1511,N_238,N_584);
and U1512 (N_1512,N_604,N_606);
or U1513 (N_1513,N_845,N_465);
nand U1514 (N_1514,N_2,N_120);
xnor U1515 (N_1515,N_317,N_823);
or U1516 (N_1516,N_860,N_969);
or U1517 (N_1517,N_486,N_316);
nand U1518 (N_1518,N_635,N_435);
or U1519 (N_1519,N_998,N_388);
and U1520 (N_1520,N_688,N_124);
and U1521 (N_1521,N_61,N_566);
nor U1522 (N_1522,N_629,N_91);
or U1523 (N_1523,N_930,N_508);
nand U1524 (N_1524,N_205,N_937);
nor U1525 (N_1525,N_178,N_551);
or U1526 (N_1526,N_47,N_373);
nand U1527 (N_1527,N_299,N_257);
or U1528 (N_1528,N_648,N_521);
and U1529 (N_1529,N_785,N_176);
nor U1530 (N_1530,N_229,N_547);
or U1531 (N_1531,N_375,N_922);
xnor U1532 (N_1532,N_228,N_20);
nand U1533 (N_1533,N_955,N_57);
and U1534 (N_1534,N_242,N_254);
and U1535 (N_1535,N_235,N_542);
and U1536 (N_1536,N_410,N_957);
nand U1537 (N_1537,N_601,N_329);
nor U1538 (N_1538,N_503,N_397);
nand U1539 (N_1539,N_979,N_518);
xor U1540 (N_1540,N_543,N_708);
or U1541 (N_1541,N_441,N_886);
nand U1542 (N_1542,N_473,N_128);
nor U1543 (N_1543,N_542,N_390);
nand U1544 (N_1544,N_367,N_987);
nand U1545 (N_1545,N_264,N_54);
nor U1546 (N_1546,N_674,N_124);
nor U1547 (N_1547,N_960,N_250);
nand U1548 (N_1548,N_809,N_635);
nor U1549 (N_1549,N_642,N_257);
and U1550 (N_1550,N_709,N_378);
and U1551 (N_1551,N_416,N_203);
or U1552 (N_1552,N_455,N_879);
nor U1553 (N_1553,N_35,N_663);
and U1554 (N_1554,N_641,N_299);
and U1555 (N_1555,N_359,N_691);
nand U1556 (N_1556,N_348,N_826);
and U1557 (N_1557,N_428,N_970);
or U1558 (N_1558,N_566,N_794);
nor U1559 (N_1559,N_847,N_349);
or U1560 (N_1560,N_576,N_633);
and U1561 (N_1561,N_936,N_283);
or U1562 (N_1562,N_325,N_755);
or U1563 (N_1563,N_537,N_708);
or U1564 (N_1564,N_752,N_511);
nand U1565 (N_1565,N_517,N_452);
nand U1566 (N_1566,N_105,N_165);
and U1567 (N_1567,N_530,N_333);
or U1568 (N_1568,N_795,N_305);
or U1569 (N_1569,N_810,N_444);
nor U1570 (N_1570,N_105,N_705);
nand U1571 (N_1571,N_511,N_333);
and U1572 (N_1572,N_236,N_961);
and U1573 (N_1573,N_511,N_243);
or U1574 (N_1574,N_862,N_233);
and U1575 (N_1575,N_772,N_32);
or U1576 (N_1576,N_289,N_115);
and U1577 (N_1577,N_968,N_133);
or U1578 (N_1578,N_757,N_233);
nand U1579 (N_1579,N_803,N_871);
or U1580 (N_1580,N_396,N_644);
nor U1581 (N_1581,N_790,N_704);
or U1582 (N_1582,N_473,N_514);
nor U1583 (N_1583,N_313,N_802);
or U1584 (N_1584,N_162,N_688);
xor U1585 (N_1585,N_119,N_205);
nand U1586 (N_1586,N_803,N_119);
nor U1587 (N_1587,N_499,N_120);
or U1588 (N_1588,N_888,N_142);
or U1589 (N_1589,N_414,N_661);
and U1590 (N_1590,N_898,N_542);
or U1591 (N_1591,N_101,N_45);
xor U1592 (N_1592,N_118,N_604);
nand U1593 (N_1593,N_963,N_375);
and U1594 (N_1594,N_324,N_501);
or U1595 (N_1595,N_424,N_248);
xnor U1596 (N_1596,N_978,N_654);
or U1597 (N_1597,N_625,N_468);
and U1598 (N_1598,N_825,N_447);
nor U1599 (N_1599,N_28,N_265);
nor U1600 (N_1600,N_457,N_22);
nand U1601 (N_1601,N_549,N_904);
or U1602 (N_1602,N_367,N_999);
nand U1603 (N_1603,N_407,N_773);
and U1604 (N_1604,N_784,N_93);
or U1605 (N_1605,N_851,N_863);
nand U1606 (N_1606,N_507,N_528);
nand U1607 (N_1607,N_892,N_582);
or U1608 (N_1608,N_531,N_264);
nand U1609 (N_1609,N_656,N_826);
nor U1610 (N_1610,N_802,N_151);
and U1611 (N_1611,N_136,N_344);
and U1612 (N_1612,N_743,N_822);
or U1613 (N_1613,N_893,N_670);
nand U1614 (N_1614,N_543,N_227);
nand U1615 (N_1615,N_145,N_863);
and U1616 (N_1616,N_574,N_398);
or U1617 (N_1617,N_508,N_66);
nor U1618 (N_1618,N_96,N_174);
nand U1619 (N_1619,N_669,N_904);
xnor U1620 (N_1620,N_60,N_317);
nor U1621 (N_1621,N_205,N_191);
or U1622 (N_1622,N_51,N_62);
and U1623 (N_1623,N_789,N_664);
nor U1624 (N_1624,N_523,N_616);
or U1625 (N_1625,N_344,N_6);
or U1626 (N_1626,N_964,N_682);
nor U1627 (N_1627,N_892,N_796);
nand U1628 (N_1628,N_525,N_524);
and U1629 (N_1629,N_595,N_193);
or U1630 (N_1630,N_29,N_501);
or U1631 (N_1631,N_133,N_650);
xor U1632 (N_1632,N_876,N_535);
nand U1633 (N_1633,N_242,N_481);
nand U1634 (N_1634,N_982,N_221);
and U1635 (N_1635,N_487,N_532);
and U1636 (N_1636,N_299,N_31);
nor U1637 (N_1637,N_876,N_350);
or U1638 (N_1638,N_241,N_677);
nor U1639 (N_1639,N_378,N_411);
nand U1640 (N_1640,N_936,N_274);
nor U1641 (N_1641,N_699,N_931);
and U1642 (N_1642,N_107,N_643);
or U1643 (N_1643,N_577,N_528);
nand U1644 (N_1644,N_269,N_484);
nor U1645 (N_1645,N_416,N_295);
xnor U1646 (N_1646,N_755,N_352);
and U1647 (N_1647,N_873,N_290);
nor U1648 (N_1648,N_447,N_912);
and U1649 (N_1649,N_625,N_744);
nand U1650 (N_1650,N_476,N_203);
nor U1651 (N_1651,N_270,N_911);
nor U1652 (N_1652,N_955,N_765);
and U1653 (N_1653,N_730,N_510);
nor U1654 (N_1654,N_177,N_705);
nand U1655 (N_1655,N_126,N_744);
nand U1656 (N_1656,N_704,N_452);
nor U1657 (N_1657,N_874,N_392);
and U1658 (N_1658,N_74,N_125);
or U1659 (N_1659,N_683,N_412);
nand U1660 (N_1660,N_341,N_721);
and U1661 (N_1661,N_232,N_339);
nand U1662 (N_1662,N_805,N_472);
nand U1663 (N_1663,N_512,N_937);
and U1664 (N_1664,N_513,N_220);
nand U1665 (N_1665,N_353,N_161);
and U1666 (N_1666,N_903,N_850);
nand U1667 (N_1667,N_642,N_936);
nor U1668 (N_1668,N_245,N_868);
nor U1669 (N_1669,N_881,N_127);
nand U1670 (N_1670,N_581,N_37);
and U1671 (N_1671,N_519,N_966);
nand U1672 (N_1672,N_39,N_906);
and U1673 (N_1673,N_423,N_55);
nand U1674 (N_1674,N_514,N_973);
nand U1675 (N_1675,N_291,N_657);
and U1676 (N_1676,N_498,N_244);
or U1677 (N_1677,N_199,N_307);
or U1678 (N_1678,N_58,N_165);
or U1679 (N_1679,N_611,N_465);
nor U1680 (N_1680,N_380,N_65);
xor U1681 (N_1681,N_680,N_760);
nor U1682 (N_1682,N_376,N_667);
and U1683 (N_1683,N_836,N_377);
nor U1684 (N_1684,N_35,N_826);
and U1685 (N_1685,N_398,N_479);
nor U1686 (N_1686,N_679,N_379);
or U1687 (N_1687,N_729,N_513);
and U1688 (N_1688,N_97,N_632);
nand U1689 (N_1689,N_285,N_231);
xnor U1690 (N_1690,N_974,N_391);
and U1691 (N_1691,N_265,N_41);
nand U1692 (N_1692,N_397,N_432);
nor U1693 (N_1693,N_928,N_589);
nand U1694 (N_1694,N_578,N_649);
nand U1695 (N_1695,N_337,N_177);
or U1696 (N_1696,N_483,N_897);
nor U1697 (N_1697,N_558,N_578);
nor U1698 (N_1698,N_375,N_143);
nor U1699 (N_1699,N_611,N_669);
and U1700 (N_1700,N_622,N_632);
xor U1701 (N_1701,N_283,N_82);
or U1702 (N_1702,N_445,N_139);
nor U1703 (N_1703,N_906,N_333);
nor U1704 (N_1704,N_65,N_600);
nor U1705 (N_1705,N_551,N_550);
and U1706 (N_1706,N_699,N_636);
or U1707 (N_1707,N_764,N_211);
nor U1708 (N_1708,N_738,N_507);
or U1709 (N_1709,N_688,N_967);
nor U1710 (N_1710,N_535,N_776);
xnor U1711 (N_1711,N_173,N_758);
and U1712 (N_1712,N_97,N_54);
nor U1713 (N_1713,N_516,N_347);
and U1714 (N_1714,N_8,N_902);
nor U1715 (N_1715,N_802,N_791);
nand U1716 (N_1716,N_202,N_24);
nor U1717 (N_1717,N_213,N_752);
or U1718 (N_1718,N_154,N_829);
or U1719 (N_1719,N_835,N_221);
nand U1720 (N_1720,N_593,N_891);
xor U1721 (N_1721,N_664,N_208);
nand U1722 (N_1722,N_750,N_682);
nand U1723 (N_1723,N_580,N_268);
nand U1724 (N_1724,N_959,N_967);
nand U1725 (N_1725,N_854,N_24);
nand U1726 (N_1726,N_305,N_903);
or U1727 (N_1727,N_372,N_708);
nand U1728 (N_1728,N_72,N_627);
nand U1729 (N_1729,N_433,N_480);
or U1730 (N_1730,N_666,N_552);
or U1731 (N_1731,N_178,N_237);
nor U1732 (N_1732,N_923,N_349);
nand U1733 (N_1733,N_804,N_41);
nor U1734 (N_1734,N_981,N_694);
and U1735 (N_1735,N_42,N_829);
and U1736 (N_1736,N_716,N_391);
or U1737 (N_1737,N_291,N_841);
nand U1738 (N_1738,N_491,N_13);
or U1739 (N_1739,N_532,N_640);
or U1740 (N_1740,N_469,N_32);
nand U1741 (N_1741,N_195,N_904);
or U1742 (N_1742,N_374,N_461);
or U1743 (N_1743,N_248,N_73);
or U1744 (N_1744,N_993,N_229);
or U1745 (N_1745,N_80,N_305);
nand U1746 (N_1746,N_228,N_796);
nand U1747 (N_1747,N_567,N_957);
nor U1748 (N_1748,N_9,N_927);
and U1749 (N_1749,N_745,N_993);
nand U1750 (N_1750,N_613,N_85);
nor U1751 (N_1751,N_115,N_592);
nor U1752 (N_1752,N_724,N_443);
and U1753 (N_1753,N_540,N_201);
or U1754 (N_1754,N_768,N_156);
nand U1755 (N_1755,N_149,N_454);
nor U1756 (N_1756,N_849,N_711);
xor U1757 (N_1757,N_420,N_752);
or U1758 (N_1758,N_107,N_338);
and U1759 (N_1759,N_612,N_757);
nand U1760 (N_1760,N_313,N_837);
or U1761 (N_1761,N_993,N_330);
and U1762 (N_1762,N_331,N_784);
or U1763 (N_1763,N_87,N_135);
or U1764 (N_1764,N_279,N_373);
nand U1765 (N_1765,N_642,N_617);
nor U1766 (N_1766,N_655,N_315);
nand U1767 (N_1767,N_450,N_475);
or U1768 (N_1768,N_85,N_979);
xor U1769 (N_1769,N_523,N_206);
nor U1770 (N_1770,N_833,N_401);
nand U1771 (N_1771,N_876,N_671);
nor U1772 (N_1772,N_964,N_162);
nor U1773 (N_1773,N_272,N_123);
and U1774 (N_1774,N_662,N_605);
and U1775 (N_1775,N_384,N_687);
nor U1776 (N_1776,N_726,N_687);
nor U1777 (N_1777,N_128,N_57);
nand U1778 (N_1778,N_378,N_100);
nor U1779 (N_1779,N_567,N_417);
nor U1780 (N_1780,N_811,N_3);
nor U1781 (N_1781,N_2,N_290);
nand U1782 (N_1782,N_762,N_797);
or U1783 (N_1783,N_251,N_539);
nor U1784 (N_1784,N_960,N_902);
nand U1785 (N_1785,N_844,N_587);
or U1786 (N_1786,N_142,N_718);
and U1787 (N_1787,N_411,N_468);
nor U1788 (N_1788,N_179,N_154);
or U1789 (N_1789,N_817,N_843);
or U1790 (N_1790,N_821,N_232);
or U1791 (N_1791,N_424,N_584);
nor U1792 (N_1792,N_0,N_726);
nand U1793 (N_1793,N_392,N_149);
xnor U1794 (N_1794,N_297,N_647);
or U1795 (N_1795,N_993,N_695);
and U1796 (N_1796,N_490,N_853);
nor U1797 (N_1797,N_949,N_996);
or U1798 (N_1798,N_786,N_656);
xor U1799 (N_1799,N_39,N_778);
xor U1800 (N_1800,N_629,N_326);
xnor U1801 (N_1801,N_176,N_984);
and U1802 (N_1802,N_626,N_460);
and U1803 (N_1803,N_13,N_820);
or U1804 (N_1804,N_334,N_674);
or U1805 (N_1805,N_125,N_853);
or U1806 (N_1806,N_114,N_802);
nand U1807 (N_1807,N_894,N_687);
xor U1808 (N_1808,N_675,N_773);
and U1809 (N_1809,N_922,N_739);
xor U1810 (N_1810,N_489,N_829);
nand U1811 (N_1811,N_370,N_172);
nor U1812 (N_1812,N_80,N_84);
and U1813 (N_1813,N_977,N_523);
and U1814 (N_1814,N_623,N_220);
and U1815 (N_1815,N_441,N_401);
and U1816 (N_1816,N_728,N_536);
nand U1817 (N_1817,N_538,N_921);
and U1818 (N_1818,N_511,N_758);
or U1819 (N_1819,N_243,N_31);
nor U1820 (N_1820,N_408,N_853);
nor U1821 (N_1821,N_102,N_657);
or U1822 (N_1822,N_445,N_126);
xor U1823 (N_1823,N_649,N_125);
nand U1824 (N_1824,N_73,N_669);
nand U1825 (N_1825,N_866,N_412);
nand U1826 (N_1826,N_973,N_923);
and U1827 (N_1827,N_148,N_387);
nor U1828 (N_1828,N_476,N_229);
nor U1829 (N_1829,N_463,N_969);
or U1830 (N_1830,N_494,N_101);
and U1831 (N_1831,N_7,N_427);
or U1832 (N_1832,N_430,N_504);
xnor U1833 (N_1833,N_42,N_731);
or U1834 (N_1834,N_922,N_571);
and U1835 (N_1835,N_904,N_288);
and U1836 (N_1836,N_990,N_532);
and U1837 (N_1837,N_75,N_845);
and U1838 (N_1838,N_580,N_611);
and U1839 (N_1839,N_664,N_595);
nor U1840 (N_1840,N_45,N_751);
or U1841 (N_1841,N_796,N_566);
nor U1842 (N_1842,N_947,N_362);
xor U1843 (N_1843,N_514,N_305);
or U1844 (N_1844,N_73,N_13);
or U1845 (N_1845,N_816,N_883);
or U1846 (N_1846,N_659,N_433);
xor U1847 (N_1847,N_482,N_867);
nand U1848 (N_1848,N_79,N_15);
nor U1849 (N_1849,N_470,N_225);
nand U1850 (N_1850,N_907,N_84);
or U1851 (N_1851,N_202,N_940);
nor U1852 (N_1852,N_850,N_680);
nand U1853 (N_1853,N_447,N_936);
or U1854 (N_1854,N_396,N_218);
xnor U1855 (N_1855,N_278,N_690);
and U1856 (N_1856,N_279,N_932);
nor U1857 (N_1857,N_751,N_423);
nor U1858 (N_1858,N_191,N_684);
nand U1859 (N_1859,N_963,N_831);
nor U1860 (N_1860,N_924,N_229);
and U1861 (N_1861,N_422,N_442);
and U1862 (N_1862,N_899,N_30);
xnor U1863 (N_1863,N_957,N_152);
nand U1864 (N_1864,N_690,N_729);
or U1865 (N_1865,N_730,N_365);
xor U1866 (N_1866,N_179,N_876);
nor U1867 (N_1867,N_653,N_933);
nor U1868 (N_1868,N_778,N_568);
nor U1869 (N_1869,N_323,N_664);
nand U1870 (N_1870,N_55,N_43);
nor U1871 (N_1871,N_327,N_817);
and U1872 (N_1872,N_967,N_710);
nand U1873 (N_1873,N_112,N_773);
and U1874 (N_1874,N_929,N_875);
and U1875 (N_1875,N_470,N_125);
and U1876 (N_1876,N_401,N_745);
and U1877 (N_1877,N_89,N_300);
or U1878 (N_1878,N_348,N_686);
nand U1879 (N_1879,N_30,N_919);
or U1880 (N_1880,N_140,N_322);
nor U1881 (N_1881,N_718,N_842);
nand U1882 (N_1882,N_826,N_866);
nor U1883 (N_1883,N_160,N_366);
and U1884 (N_1884,N_32,N_432);
nand U1885 (N_1885,N_218,N_349);
nor U1886 (N_1886,N_695,N_529);
and U1887 (N_1887,N_16,N_628);
nand U1888 (N_1888,N_757,N_584);
nand U1889 (N_1889,N_217,N_590);
and U1890 (N_1890,N_455,N_495);
or U1891 (N_1891,N_958,N_813);
or U1892 (N_1892,N_245,N_918);
and U1893 (N_1893,N_313,N_248);
xnor U1894 (N_1894,N_522,N_882);
nand U1895 (N_1895,N_467,N_90);
nor U1896 (N_1896,N_329,N_788);
nor U1897 (N_1897,N_893,N_718);
nor U1898 (N_1898,N_343,N_789);
and U1899 (N_1899,N_443,N_881);
xnor U1900 (N_1900,N_209,N_686);
nor U1901 (N_1901,N_670,N_505);
nand U1902 (N_1902,N_532,N_679);
xnor U1903 (N_1903,N_893,N_965);
or U1904 (N_1904,N_252,N_645);
and U1905 (N_1905,N_585,N_96);
or U1906 (N_1906,N_871,N_684);
nand U1907 (N_1907,N_666,N_224);
or U1908 (N_1908,N_505,N_798);
xor U1909 (N_1909,N_474,N_773);
or U1910 (N_1910,N_134,N_31);
and U1911 (N_1911,N_557,N_230);
or U1912 (N_1912,N_180,N_978);
nor U1913 (N_1913,N_791,N_341);
and U1914 (N_1914,N_81,N_356);
nor U1915 (N_1915,N_34,N_68);
nand U1916 (N_1916,N_726,N_124);
nand U1917 (N_1917,N_45,N_414);
nor U1918 (N_1918,N_336,N_6);
nand U1919 (N_1919,N_640,N_865);
xnor U1920 (N_1920,N_109,N_932);
nand U1921 (N_1921,N_12,N_573);
nand U1922 (N_1922,N_664,N_820);
nor U1923 (N_1923,N_804,N_459);
nor U1924 (N_1924,N_562,N_709);
and U1925 (N_1925,N_31,N_1);
and U1926 (N_1926,N_234,N_992);
or U1927 (N_1927,N_737,N_438);
or U1928 (N_1928,N_286,N_751);
and U1929 (N_1929,N_366,N_131);
nor U1930 (N_1930,N_822,N_298);
nor U1931 (N_1931,N_261,N_724);
and U1932 (N_1932,N_8,N_605);
or U1933 (N_1933,N_119,N_302);
nand U1934 (N_1934,N_512,N_225);
and U1935 (N_1935,N_904,N_658);
and U1936 (N_1936,N_937,N_162);
or U1937 (N_1937,N_631,N_745);
nand U1938 (N_1938,N_668,N_998);
nor U1939 (N_1939,N_223,N_767);
or U1940 (N_1940,N_901,N_946);
and U1941 (N_1941,N_925,N_252);
xor U1942 (N_1942,N_297,N_26);
and U1943 (N_1943,N_390,N_960);
nand U1944 (N_1944,N_614,N_470);
xor U1945 (N_1945,N_546,N_175);
nand U1946 (N_1946,N_976,N_823);
and U1947 (N_1947,N_156,N_956);
nor U1948 (N_1948,N_454,N_965);
and U1949 (N_1949,N_429,N_210);
nand U1950 (N_1950,N_457,N_758);
nor U1951 (N_1951,N_634,N_131);
or U1952 (N_1952,N_646,N_1);
and U1953 (N_1953,N_730,N_228);
nand U1954 (N_1954,N_937,N_243);
nand U1955 (N_1955,N_44,N_562);
or U1956 (N_1956,N_995,N_484);
and U1957 (N_1957,N_919,N_994);
nor U1958 (N_1958,N_765,N_768);
or U1959 (N_1959,N_119,N_579);
xnor U1960 (N_1960,N_801,N_962);
xor U1961 (N_1961,N_979,N_625);
nor U1962 (N_1962,N_597,N_26);
nand U1963 (N_1963,N_327,N_632);
nor U1964 (N_1964,N_952,N_289);
or U1965 (N_1965,N_699,N_536);
nor U1966 (N_1966,N_705,N_513);
nor U1967 (N_1967,N_476,N_607);
nand U1968 (N_1968,N_569,N_581);
nand U1969 (N_1969,N_365,N_792);
and U1970 (N_1970,N_765,N_692);
and U1971 (N_1971,N_836,N_973);
nor U1972 (N_1972,N_693,N_317);
xor U1973 (N_1973,N_383,N_897);
and U1974 (N_1974,N_891,N_332);
nor U1975 (N_1975,N_917,N_731);
nand U1976 (N_1976,N_176,N_53);
nand U1977 (N_1977,N_618,N_347);
or U1978 (N_1978,N_556,N_136);
nor U1979 (N_1979,N_305,N_863);
or U1980 (N_1980,N_714,N_558);
and U1981 (N_1981,N_920,N_861);
nand U1982 (N_1982,N_632,N_427);
nor U1983 (N_1983,N_54,N_577);
xor U1984 (N_1984,N_903,N_869);
nand U1985 (N_1985,N_101,N_172);
nand U1986 (N_1986,N_538,N_681);
nand U1987 (N_1987,N_862,N_342);
xnor U1988 (N_1988,N_79,N_63);
or U1989 (N_1989,N_304,N_416);
and U1990 (N_1990,N_915,N_499);
nand U1991 (N_1991,N_281,N_309);
nand U1992 (N_1992,N_477,N_450);
xnor U1993 (N_1993,N_109,N_389);
and U1994 (N_1994,N_787,N_429);
nand U1995 (N_1995,N_793,N_633);
nand U1996 (N_1996,N_105,N_196);
nor U1997 (N_1997,N_772,N_748);
nor U1998 (N_1998,N_873,N_103);
nand U1999 (N_1999,N_73,N_245);
nand U2000 (N_2000,N_1947,N_1581);
nand U2001 (N_2001,N_1070,N_1973);
and U2002 (N_2002,N_1095,N_1414);
nand U2003 (N_2003,N_1406,N_1236);
nor U2004 (N_2004,N_1059,N_1339);
or U2005 (N_2005,N_1341,N_1412);
or U2006 (N_2006,N_1606,N_1665);
or U2007 (N_2007,N_1211,N_1092);
or U2008 (N_2008,N_1161,N_1175);
nand U2009 (N_2009,N_1895,N_1754);
and U2010 (N_2010,N_1894,N_1036);
or U2011 (N_2011,N_1787,N_1387);
nand U2012 (N_2012,N_1410,N_1584);
or U2013 (N_2013,N_1967,N_1859);
nand U2014 (N_2014,N_1363,N_1112);
or U2015 (N_2015,N_1110,N_1284);
or U2016 (N_2016,N_1248,N_1190);
nor U2017 (N_2017,N_1825,N_1186);
and U2018 (N_2018,N_1571,N_1328);
xnor U2019 (N_2019,N_1922,N_1409);
nor U2020 (N_2020,N_1702,N_1327);
nand U2021 (N_2021,N_1398,N_1537);
nor U2022 (N_2022,N_1631,N_1324);
and U2023 (N_2023,N_1645,N_1561);
nand U2024 (N_2024,N_1256,N_1336);
nor U2025 (N_2025,N_1290,N_1907);
and U2026 (N_2026,N_1260,N_1669);
nand U2027 (N_2027,N_1172,N_1831);
nand U2028 (N_2028,N_1629,N_1701);
nor U2029 (N_2029,N_1744,N_1055);
nand U2030 (N_2030,N_1488,N_1653);
or U2031 (N_2031,N_1782,N_1677);
or U2032 (N_2032,N_1026,N_1741);
nor U2033 (N_2033,N_1507,N_1963);
or U2034 (N_2034,N_1940,N_1345);
nor U2035 (N_2035,N_1297,N_1128);
nand U2036 (N_2036,N_1930,N_1289);
nor U2037 (N_2037,N_1021,N_1827);
nand U2038 (N_2038,N_1892,N_1288);
and U2039 (N_2039,N_1249,N_1252);
or U2040 (N_2040,N_1302,N_1797);
and U2041 (N_2041,N_1534,N_1514);
or U2042 (N_2042,N_1675,N_1313);
nand U2043 (N_2043,N_1893,N_1673);
or U2044 (N_2044,N_1857,N_1871);
xnor U2045 (N_2045,N_1109,N_1433);
xor U2046 (N_2046,N_1216,N_1725);
nor U2047 (N_2047,N_1119,N_1776);
and U2048 (N_2048,N_1380,N_1114);
and U2049 (N_2049,N_1937,N_1218);
xnor U2050 (N_2050,N_1411,N_1436);
or U2051 (N_2051,N_1033,N_1599);
or U2052 (N_2052,N_1564,N_1505);
nor U2053 (N_2053,N_1789,N_1971);
xor U2054 (N_2054,N_1699,N_1590);
nor U2055 (N_2055,N_1246,N_1272);
nand U2056 (N_2056,N_1586,N_1203);
nand U2057 (N_2057,N_1662,N_1781);
nand U2058 (N_2058,N_1157,N_1393);
or U2059 (N_2059,N_1113,N_1742);
nand U2060 (N_2060,N_1364,N_1147);
nor U2061 (N_2061,N_1220,N_1957);
nor U2062 (N_2062,N_1550,N_1862);
and U2063 (N_2063,N_1138,N_1126);
and U2064 (N_2064,N_1580,N_1987);
and U2065 (N_2065,N_1291,N_1108);
or U2066 (N_2066,N_1655,N_1259);
nor U2067 (N_2067,N_1262,N_1883);
nand U2068 (N_2068,N_1603,N_1080);
nor U2069 (N_2069,N_1887,N_1232);
and U2070 (N_2070,N_1545,N_1555);
or U2071 (N_2071,N_1698,N_1714);
or U2072 (N_2072,N_1576,N_1355);
nand U2073 (N_2073,N_1786,N_1484);
or U2074 (N_2074,N_1525,N_1356);
nand U2075 (N_2075,N_1891,N_1337);
and U2076 (N_2076,N_1391,N_1740);
or U2077 (N_2077,N_1899,N_1107);
nand U2078 (N_2078,N_1243,N_1239);
nor U2079 (N_2079,N_1913,N_1314);
nor U2080 (N_2080,N_1925,N_1150);
and U2081 (N_2081,N_1478,N_1533);
nor U2082 (N_2082,N_1148,N_1774);
and U2083 (N_2083,N_1997,N_1476);
and U2084 (N_2084,N_1097,N_1932);
nor U2085 (N_2085,N_1521,N_1501);
nand U2086 (N_2086,N_1156,N_1226);
nor U2087 (N_2087,N_1919,N_1060);
and U2088 (N_2088,N_1568,N_1622);
nand U2089 (N_2089,N_1096,N_1779);
and U2090 (N_2090,N_1106,N_1192);
and U2091 (N_2091,N_1303,N_1764);
nor U2092 (N_2092,N_1807,N_1610);
or U2093 (N_2093,N_1715,N_1441);
nand U2094 (N_2094,N_1196,N_1648);
and U2095 (N_2095,N_1105,N_1517);
and U2096 (N_2096,N_1258,N_1222);
nand U2097 (N_2097,N_1018,N_1408);
nand U2098 (N_2098,N_1277,N_1663);
nand U2099 (N_2099,N_1591,N_1049);
or U2100 (N_2100,N_1791,N_1560);
nor U2101 (N_2101,N_1473,N_1149);
nand U2102 (N_2102,N_1357,N_1605);
or U2103 (N_2103,N_1811,N_1856);
and U2104 (N_2104,N_1301,N_1998);
nand U2105 (N_2105,N_1170,N_1474);
nand U2106 (N_2106,N_1566,N_1162);
nand U2107 (N_2107,N_1888,N_1019);
nand U2108 (N_2108,N_1767,N_1295);
and U2109 (N_2109,N_1443,N_1445);
xnor U2110 (N_2110,N_1985,N_1898);
nand U2111 (N_2111,N_1952,N_1037);
nor U2112 (N_2112,N_1743,N_1270);
nand U2113 (N_2113,N_1536,N_1210);
nor U2114 (N_2114,N_1950,N_1159);
nand U2115 (N_2115,N_1184,N_1494);
nand U2116 (N_2116,N_1944,N_1510);
nor U2117 (N_2117,N_1678,N_1956);
nor U2118 (N_2118,N_1395,N_1373);
and U2119 (N_2119,N_1100,N_1469);
and U2120 (N_2120,N_1348,N_1145);
xor U2121 (N_2121,N_1233,N_1934);
nor U2122 (N_2122,N_1821,N_1200);
and U2123 (N_2123,N_1869,N_1617);
or U2124 (N_2124,N_1264,N_1959);
or U2125 (N_2125,N_1874,N_1072);
or U2126 (N_2126,N_1823,N_1083);
nor U2127 (N_2127,N_1578,N_1227);
nand U2128 (N_2128,N_1250,N_1317);
nand U2129 (N_2129,N_1735,N_1890);
and U2130 (N_2130,N_1692,N_1158);
nor U2131 (N_2131,N_1043,N_1378);
nor U2132 (N_2132,N_1838,N_1637);
and U2133 (N_2133,N_1736,N_1604);
or U2134 (N_2134,N_1416,N_1076);
nor U2135 (N_2135,N_1130,N_1608);
nor U2136 (N_2136,N_1589,N_1292);
nor U2137 (N_2137,N_1921,N_1583);
nor U2138 (N_2138,N_1795,N_1872);
nand U2139 (N_2139,N_1194,N_1727);
xor U2140 (N_2140,N_1513,N_1152);
or U2141 (N_2141,N_1897,N_1720);
and U2142 (N_2142,N_1929,N_1177);
nor U2143 (N_2143,N_1452,N_1480);
nand U2144 (N_2144,N_1592,N_1875);
nor U2145 (N_2145,N_1247,N_1667);
nand U2146 (N_2146,N_1319,N_1431);
nand U2147 (N_2147,N_1224,N_1722);
and U2148 (N_2148,N_1084,N_1668);
xor U2149 (N_2149,N_1496,N_1151);
nand U2150 (N_2150,N_1529,N_1091);
and U2151 (N_2151,N_1657,N_1309);
and U2152 (N_2152,N_1928,N_1418);
or U2153 (N_2153,N_1619,N_1207);
and U2154 (N_2154,N_1658,N_1293);
or U2155 (N_2155,N_1647,N_1738);
nor U2156 (N_2156,N_1274,N_1864);
or U2157 (N_2157,N_1772,N_1075);
or U2158 (N_2158,N_1552,N_1951);
or U2159 (N_2159,N_1818,N_1691);
nor U2160 (N_2160,N_1127,N_1174);
and U2161 (N_2161,N_1515,N_1674);
nor U2162 (N_2162,N_1731,N_1069);
or U2163 (N_2163,N_1164,N_1173);
nand U2164 (N_2164,N_1755,N_1547);
nand U2165 (N_2165,N_1168,N_1372);
or U2166 (N_2166,N_1090,N_1980);
or U2167 (N_2167,N_1300,N_1650);
xor U2168 (N_2168,N_1051,N_1509);
or U2169 (N_2169,N_1439,N_1326);
and U2170 (N_2170,N_1118,N_1009);
nor U2171 (N_2171,N_1392,N_1972);
and U2172 (N_2172,N_1073,N_1625);
and U2173 (N_2173,N_1935,N_1046);
and U2174 (N_2174,N_1464,N_1282);
or U2175 (N_2175,N_1349,N_1504);
nand U2176 (N_2176,N_1187,N_1188);
xor U2177 (N_2177,N_1633,N_1982);
nand U2178 (N_2178,N_1038,N_1557);
nand U2179 (N_2179,N_1041,N_1426);
and U2180 (N_2180,N_1362,N_1989);
and U2181 (N_2181,N_1384,N_1066);
nor U2182 (N_2182,N_1730,N_1749);
nor U2183 (N_2183,N_1679,N_1098);
and U2184 (N_2184,N_1966,N_1945);
or U2185 (N_2185,N_1153,N_1052);
nand U2186 (N_2186,N_1191,N_1732);
nand U2187 (N_2187,N_1056,N_1206);
nand U2188 (N_2188,N_1938,N_1129);
nand U2189 (N_2189,N_1866,N_1810);
nand U2190 (N_2190,N_1485,N_1962);
or U2191 (N_2191,N_1030,N_1794);
and U2192 (N_2192,N_1949,N_1830);
nor U2193 (N_2193,N_1569,N_1548);
and U2194 (N_2194,N_1718,N_1020);
nand U2195 (N_2195,N_1582,N_1961);
nand U2196 (N_2196,N_1636,N_1427);
nor U2197 (N_2197,N_1765,N_1242);
nand U2198 (N_2198,N_1429,N_1588);
or U2199 (N_2199,N_1401,N_1681);
or U2200 (N_2200,N_1824,N_1029);
and U2201 (N_2201,N_1487,N_1077);
nand U2202 (N_2202,N_1848,N_1993);
and U2203 (N_2203,N_1627,N_1438);
nand U2204 (N_2204,N_1390,N_1748);
nor U2205 (N_2205,N_1986,N_1179);
nand U2206 (N_2206,N_1121,N_1843);
nand U2207 (N_2207,N_1228,N_1757);
nand U2208 (N_2208,N_1027,N_1778);
nand U2209 (N_2209,N_1909,N_1538);
nand U2210 (N_2210,N_1523,N_1528);
nor U2211 (N_2211,N_1946,N_1616);
or U2212 (N_2212,N_1717,N_1331);
xor U2213 (N_2213,N_1155,N_1209);
nor U2214 (N_2214,N_1212,N_1139);
or U2215 (N_2215,N_1858,N_1388);
and U2216 (N_2216,N_1750,N_1450);
xor U2217 (N_2217,N_1775,N_1965);
and U2218 (N_2218,N_1885,N_1712);
nor U2219 (N_2219,N_1527,N_1976);
and U2220 (N_2220,N_1316,N_1422);
and U2221 (N_2221,N_1612,N_1465);
xnor U2222 (N_2222,N_1752,N_1086);
nor U2223 (N_2223,N_1470,N_1165);
or U2224 (N_2224,N_1048,N_1013);
or U2225 (N_2225,N_1031,N_1615);
xor U2226 (N_2226,N_1912,N_1461);
nor U2227 (N_2227,N_1405,N_1724);
nor U2228 (N_2228,N_1322,N_1889);
xnor U2229 (N_2229,N_1531,N_1710);
nor U2230 (N_2230,N_1978,N_1801);
xor U2231 (N_2231,N_1511,N_1558);
nand U2232 (N_2232,N_1201,N_1628);
or U2233 (N_2233,N_1497,N_1054);
and U2234 (N_2234,N_1995,N_1845);
nor U2235 (N_2235,N_1865,N_1773);
nand U2236 (N_2236,N_1884,N_1598);
nor U2237 (N_2237,N_1554,N_1133);
and U2238 (N_2238,N_1134,N_1948);
nor U2239 (N_2239,N_1245,N_1543);
nor U2240 (N_2240,N_1910,N_1841);
or U2241 (N_2241,N_1305,N_1325);
or U2242 (N_2242,N_1131,N_1984);
nor U2243 (N_2243,N_1917,N_1283);
and U2244 (N_2244,N_1280,N_1969);
or U2245 (N_2245,N_1546,N_1400);
nor U2246 (N_2246,N_1942,N_1861);
nor U2247 (N_2247,N_1342,N_1671);
nand U2248 (N_2248,N_1320,N_1522);
and U2249 (N_2249,N_1124,N_1215);
nor U2250 (N_2250,N_1563,N_1185);
or U2251 (N_2251,N_1205,N_1047);
or U2252 (N_2252,N_1904,N_1770);
nor U2253 (N_2253,N_1235,N_1813);
xnor U2254 (N_2254,N_1672,N_1955);
xor U2255 (N_2255,N_1758,N_1613);
or U2256 (N_2256,N_1491,N_1225);
nor U2257 (N_2257,N_1307,N_1784);
nor U2258 (N_2258,N_1687,N_1639);
and U2259 (N_2259,N_1111,N_1506);
nor U2260 (N_2260,N_1991,N_1901);
xnor U2261 (N_2261,N_1466,N_1382);
nand U2262 (N_2262,N_1936,N_1479);
nor U2263 (N_2263,N_1472,N_1449);
xnor U2264 (N_2264,N_1208,N_1846);
xnor U2265 (N_2265,N_1338,N_1979);
or U2266 (N_2266,N_1067,N_1352);
nand U2267 (N_2267,N_1454,N_1595);
or U2268 (N_2268,N_1611,N_1078);
and U2269 (N_2269,N_1646,N_1182);
or U2270 (N_2270,N_1815,N_1402);
and U2271 (N_2271,N_1844,N_1000);
and U2272 (N_2272,N_1540,N_1065);
nor U2273 (N_2273,N_1189,N_1435);
nor U2274 (N_2274,N_1163,N_1340);
and U2275 (N_2275,N_1882,N_1597);
nor U2276 (N_2276,N_1323,N_1970);
and U2277 (N_2277,N_1577,N_1694);
nand U2278 (N_2278,N_1876,N_1840);
and U2279 (N_2279,N_1267,N_1117);
and U2280 (N_2280,N_1101,N_1696);
or U2281 (N_2281,N_1217,N_1093);
or U2282 (N_2282,N_1202,N_1102);
nand U2283 (N_2283,N_1123,N_1853);
nor U2284 (N_2284,N_1640,N_1574);
nand U2285 (N_2285,N_1851,N_1624);
nor U2286 (N_2286,N_1837,N_1053);
nor U2287 (N_2287,N_1361,N_1500);
or U2288 (N_2288,N_1706,N_1819);
xor U2289 (N_2289,N_1759,N_1460);
or U2290 (N_2290,N_1330,N_1321);
or U2291 (N_2291,N_1508,N_1044);
xnor U2292 (N_2292,N_1828,N_1532);
or U2293 (N_2293,N_1146,N_1012);
xnor U2294 (N_2294,N_1171,N_1050);
nor U2295 (N_2295,N_1939,N_1136);
xor U2296 (N_2296,N_1286,N_1424);
nand U2297 (N_2297,N_1676,N_1644);
xor U2298 (N_2298,N_1142,N_1335);
and U2299 (N_2299,N_1562,N_1705);
nor U2300 (N_2300,N_1870,N_1607);
and U2301 (N_2301,N_1896,N_1032);
or U2302 (N_2302,N_1726,N_1016);
and U2303 (N_2303,N_1024,N_1253);
nand U2304 (N_2304,N_1343,N_1085);
nand U2305 (N_2305,N_1780,N_1255);
and U2306 (N_2306,N_1010,N_1834);
nand U2307 (N_2307,N_1544,N_1585);
nand U2308 (N_2308,N_1421,N_1854);
or U2309 (N_2309,N_1877,N_1251);
and U2310 (N_2310,N_1573,N_1299);
and U2311 (N_2311,N_1482,N_1737);
nor U2312 (N_2312,N_1733,N_1231);
or U2313 (N_2313,N_1370,N_1601);
or U2314 (N_2314,N_1502,N_1240);
and U2315 (N_2315,N_1087,N_1456);
xor U2316 (N_2316,N_1519,N_1761);
xor U2317 (N_2317,N_1279,N_1996);
nor U2318 (N_2318,N_1058,N_1924);
nand U2319 (N_2319,N_1968,N_1001);
nor U2320 (N_2320,N_1079,N_1809);
xor U2321 (N_2321,N_1351,N_1964);
nand U2322 (N_2322,N_1863,N_1788);
nor U2323 (N_2323,N_1596,N_1878);
nor U2324 (N_2324,N_1579,N_1835);
or U2325 (N_2325,N_1306,N_1448);
or U2326 (N_2326,N_1498,N_1799);
and U2327 (N_2327,N_1334,N_1195);
nand U2328 (N_2328,N_1183,N_1816);
nand U2329 (N_2329,N_1931,N_1539);
and U2330 (N_2330,N_1287,N_1354);
or U2331 (N_2331,N_1994,N_1587);
and U2332 (N_2332,N_1790,N_1695);
or U2333 (N_2333,N_1015,N_1425);
and U2334 (N_2334,N_1855,N_1007);
nand U2335 (N_2335,N_1365,N_1381);
nor U2336 (N_2336,N_1609,N_1689);
xnor U2337 (N_2337,N_1434,N_1632);
xnor U2338 (N_2338,N_1457,N_1081);
and U2339 (N_2339,N_1729,N_1120);
and U2340 (N_2340,N_1768,N_1011);
nand U2341 (N_2341,N_1804,N_1836);
nor U2342 (N_2342,N_1181,N_1359);
or U2343 (N_2343,N_1684,N_1908);
xor U2344 (N_2344,N_1620,N_1670);
nor U2345 (N_2345,N_1760,N_1035);
and U2346 (N_2346,N_1367,N_1927);
xnor U2347 (N_2347,N_1369,N_1103);
and U2348 (N_2348,N_1278,N_1920);
nand U2349 (N_2349,N_1413,N_1734);
or U2350 (N_2350,N_1376,N_1263);
nand U2351 (N_2351,N_1800,N_1600);
and U2352 (N_2352,N_1467,N_1902);
and U2353 (N_2353,N_1753,N_1180);
or U2354 (N_2354,N_1602,N_1666);
and U2355 (N_2355,N_1304,N_1423);
nor U2356 (N_2356,N_1333,N_1254);
nor U2357 (N_2357,N_1104,N_1281);
nand U2358 (N_2358,N_1643,N_1486);
and U2359 (N_2359,N_1771,N_1943);
nand U2360 (N_2360,N_1268,N_1005);
xnor U2361 (N_2361,N_1458,N_1808);
or U2362 (N_2362,N_1905,N_1347);
and U2363 (N_2363,N_1664,N_1137);
or U2364 (N_2364,N_1451,N_1792);
nor U2365 (N_2365,N_1914,N_1089);
and U2366 (N_2366,N_1198,N_1873);
nand U2367 (N_2367,N_1238,N_1783);
nand U2368 (N_2368,N_1432,N_1614);
and U2369 (N_2369,N_1704,N_1318);
and U2370 (N_2370,N_1453,N_1852);
and U2371 (N_2371,N_1366,N_1045);
and U2372 (N_2372,N_1237,N_1368);
nor U2373 (N_2373,N_1535,N_1298);
nor U2374 (N_2374,N_1829,N_1166);
nand U2375 (N_2375,N_1039,N_1082);
nor U2376 (N_2376,N_1623,N_1014);
and U2377 (N_2377,N_1886,N_1814);
nand U2378 (N_2378,N_1350,N_1805);
and U2379 (N_2379,N_1074,N_1798);
or U2380 (N_2380,N_1371,N_1812);
and U2381 (N_2381,N_1444,N_1746);
nand U2382 (N_2382,N_1040,N_1556);
and U2383 (N_2383,N_1656,N_1265);
and U2384 (N_2384,N_1983,N_1641);
or U2385 (N_2385,N_1132,N_1524);
or U2386 (N_2386,N_1002,N_1707);
nor U2387 (N_2387,N_1399,N_1826);
nor U2388 (N_2388,N_1918,N_1630);
nor U2389 (N_2389,N_1417,N_1833);
nand U2390 (N_2390,N_1709,N_1541);
nor U2391 (N_2391,N_1219,N_1273);
and U2392 (N_2392,N_1751,N_1385);
and U2393 (N_2393,N_1652,N_1419);
xnor U2394 (N_2394,N_1042,N_1868);
and U2395 (N_2395,N_1975,N_1880);
nand U2396 (N_2396,N_1638,N_1565);
xor U2397 (N_2397,N_1197,N_1716);
nor U2398 (N_2398,N_1064,N_1559);
or U2399 (N_2399,N_1926,N_1553);
xnor U2400 (N_2400,N_1777,N_1266);
and U2401 (N_2401,N_1839,N_1881);
nand U2402 (N_2402,N_1471,N_1257);
and U2403 (N_2403,N_1455,N_1404);
nand U2404 (N_2404,N_1981,N_1397);
nor U2405 (N_2405,N_1383,N_1358);
nor U2406 (N_2406,N_1437,N_1708);
or U2407 (N_2407,N_1923,N_1685);
or U2408 (N_2408,N_1477,N_1660);
or U2409 (N_2409,N_1017,N_1403);
xnor U2410 (N_2410,N_1008,N_1683);
xor U2411 (N_2411,N_1703,N_1430);
or U2412 (N_2412,N_1649,N_1475);
nand U2413 (N_2413,N_1329,N_1088);
nor U2414 (N_2414,N_1140,N_1221);
or U2415 (N_2415,N_1806,N_1642);
nor U2416 (N_2416,N_1719,N_1346);
nand U2417 (N_2417,N_1068,N_1567);
nor U2418 (N_2418,N_1493,N_1204);
and U2419 (N_2419,N_1115,N_1960);
nor U2420 (N_2420,N_1459,N_1551);
nor U2421 (N_2421,N_1481,N_1003);
or U2422 (N_2422,N_1276,N_1867);
nor U2423 (N_2423,N_1241,N_1374);
xnor U2424 (N_2424,N_1332,N_1739);
and U2425 (N_2425,N_1353,N_1802);
xor U2426 (N_2426,N_1769,N_1229);
nor U2427 (N_2427,N_1693,N_1499);
xor U2428 (N_2428,N_1025,N_1594);
xor U2429 (N_2429,N_1230,N_1713);
or U2430 (N_2430,N_1526,N_1682);
nand U2431 (N_2431,N_1879,N_1503);
nand U2432 (N_2432,N_1261,N_1094);
nor U2433 (N_2433,N_1160,N_1178);
nor U2434 (N_2434,N_1269,N_1141);
nand U2435 (N_2435,N_1661,N_1659);
and U2436 (N_2436,N_1394,N_1489);
xor U2437 (N_2437,N_1463,N_1958);
nand U2438 (N_2438,N_1062,N_1953);
and U2439 (N_2439,N_1822,N_1954);
or U2440 (N_2440,N_1933,N_1294);
and U2441 (N_2441,N_1199,N_1575);
and U2442 (N_2442,N_1762,N_1756);
nand U2443 (N_2443,N_1022,N_1244);
nor U2444 (N_2444,N_1721,N_1803);
xnor U2445 (N_2445,N_1296,N_1990);
or U2446 (N_2446,N_1974,N_1143);
and U2447 (N_2447,N_1135,N_1377);
xor U2448 (N_2448,N_1144,N_1462);
nand U2449 (N_2449,N_1728,N_1977);
nand U2450 (N_2450,N_1023,N_1379);
and U2451 (N_2451,N_1223,N_1442);
or U2452 (N_2452,N_1006,N_1389);
and U2453 (N_2453,N_1785,N_1651);
nor U2454 (N_2454,N_1315,N_1570);
or U2455 (N_2455,N_1483,N_1697);
nand U2456 (N_2456,N_1063,N_1654);
and U2457 (N_2457,N_1490,N_1999);
xnor U2458 (N_2458,N_1116,N_1832);
and U2459 (N_2459,N_1099,N_1793);
or U2460 (N_2460,N_1635,N_1700);
and U2461 (N_2461,N_1234,N_1723);
and U2462 (N_2462,N_1518,N_1688);
or U2463 (N_2463,N_1988,N_1407);
nor U2464 (N_2464,N_1344,N_1763);
nor U2465 (N_2465,N_1903,N_1214);
nor U2466 (N_2466,N_1167,N_1285);
and U2467 (N_2467,N_1028,N_1906);
and U2468 (N_2468,N_1428,N_1992);
nand U2469 (N_2469,N_1745,N_1193);
and U2470 (N_2470,N_1154,N_1271);
nand U2471 (N_2471,N_1446,N_1916);
xor U2472 (N_2472,N_1468,N_1593);
xnor U2473 (N_2473,N_1071,N_1440);
xor U2474 (N_2474,N_1542,N_1530);
nand U2475 (N_2475,N_1311,N_1911);
or U2476 (N_2476,N_1711,N_1213);
nand U2477 (N_2477,N_1420,N_1520);
and U2478 (N_2478,N_1447,N_1941);
nand U2479 (N_2479,N_1900,N_1850);
and U2480 (N_2480,N_1312,N_1061);
nor U2481 (N_2481,N_1626,N_1549);
and U2482 (N_2482,N_1747,N_1680);
nor U2483 (N_2483,N_1310,N_1176);
and U2484 (N_2484,N_1690,N_1396);
nand U2485 (N_2485,N_1275,N_1849);
or U2486 (N_2486,N_1057,N_1618);
nor U2487 (N_2487,N_1915,N_1860);
xnor U2488 (N_2488,N_1415,N_1634);
nor U2489 (N_2489,N_1796,N_1621);
or U2490 (N_2490,N_1004,N_1386);
and U2491 (N_2491,N_1842,N_1766);
or U2492 (N_2492,N_1817,N_1375);
xnor U2493 (N_2493,N_1820,N_1360);
or U2494 (N_2494,N_1512,N_1034);
and U2495 (N_2495,N_1308,N_1492);
and U2496 (N_2496,N_1686,N_1169);
or U2497 (N_2497,N_1495,N_1122);
or U2498 (N_2498,N_1847,N_1572);
and U2499 (N_2499,N_1125,N_1516);
and U2500 (N_2500,N_1920,N_1925);
nor U2501 (N_2501,N_1813,N_1897);
or U2502 (N_2502,N_1565,N_1106);
and U2503 (N_2503,N_1729,N_1111);
xor U2504 (N_2504,N_1859,N_1416);
or U2505 (N_2505,N_1561,N_1862);
xor U2506 (N_2506,N_1473,N_1194);
nor U2507 (N_2507,N_1270,N_1910);
or U2508 (N_2508,N_1017,N_1027);
and U2509 (N_2509,N_1071,N_1669);
or U2510 (N_2510,N_1278,N_1720);
nand U2511 (N_2511,N_1869,N_1427);
and U2512 (N_2512,N_1591,N_1155);
nand U2513 (N_2513,N_1709,N_1724);
nor U2514 (N_2514,N_1011,N_1850);
and U2515 (N_2515,N_1679,N_1584);
nand U2516 (N_2516,N_1892,N_1444);
nor U2517 (N_2517,N_1025,N_1576);
or U2518 (N_2518,N_1640,N_1223);
or U2519 (N_2519,N_1091,N_1756);
or U2520 (N_2520,N_1096,N_1184);
nor U2521 (N_2521,N_1429,N_1004);
or U2522 (N_2522,N_1673,N_1309);
nor U2523 (N_2523,N_1837,N_1277);
or U2524 (N_2524,N_1111,N_1542);
nand U2525 (N_2525,N_1438,N_1537);
nand U2526 (N_2526,N_1465,N_1169);
nor U2527 (N_2527,N_1072,N_1166);
or U2528 (N_2528,N_1019,N_1890);
xnor U2529 (N_2529,N_1359,N_1660);
and U2530 (N_2530,N_1897,N_1656);
or U2531 (N_2531,N_1068,N_1563);
and U2532 (N_2532,N_1005,N_1264);
nand U2533 (N_2533,N_1357,N_1689);
and U2534 (N_2534,N_1980,N_1874);
nand U2535 (N_2535,N_1582,N_1514);
nor U2536 (N_2536,N_1758,N_1386);
and U2537 (N_2537,N_1508,N_1243);
and U2538 (N_2538,N_1240,N_1816);
nor U2539 (N_2539,N_1994,N_1690);
nor U2540 (N_2540,N_1557,N_1512);
and U2541 (N_2541,N_1376,N_1794);
xor U2542 (N_2542,N_1599,N_1904);
nand U2543 (N_2543,N_1283,N_1896);
or U2544 (N_2544,N_1014,N_1543);
or U2545 (N_2545,N_1765,N_1169);
and U2546 (N_2546,N_1988,N_1447);
nand U2547 (N_2547,N_1499,N_1462);
or U2548 (N_2548,N_1137,N_1545);
or U2549 (N_2549,N_1200,N_1183);
nand U2550 (N_2550,N_1335,N_1464);
and U2551 (N_2551,N_1843,N_1936);
and U2552 (N_2552,N_1171,N_1026);
nor U2553 (N_2553,N_1595,N_1878);
nand U2554 (N_2554,N_1245,N_1423);
and U2555 (N_2555,N_1514,N_1522);
or U2556 (N_2556,N_1467,N_1436);
or U2557 (N_2557,N_1441,N_1725);
nor U2558 (N_2558,N_1314,N_1749);
or U2559 (N_2559,N_1491,N_1749);
nor U2560 (N_2560,N_1447,N_1107);
nor U2561 (N_2561,N_1949,N_1652);
or U2562 (N_2562,N_1669,N_1627);
xnor U2563 (N_2563,N_1656,N_1828);
nor U2564 (N_2564,N_1729,N_1639);
xor U2565 (N_2565,N_1827,N_1624);
or U2566 (N_2566,N_1653,N_1968);
nand U2567 (N_2567,N_1391,N_1303);
or U2568 (N_2568,N_1389,N_1573);
nand U2569 (N_2569,N_1967,N_1402);
or U2570 (N_2570,N_1604,N_1738);
xnor U2571 (N_2571,N_1999,N_1675);
nor U2572 (N_2572,N_1214,N_1216);
and U2573 (N_2573,N_1521,N_1787);
or U2574 (N_2574,N_1505,N_1129);
or U2575 (N_2575,N_1745,N_1314);
nand U2576 (N_2576,N_1104,N_1747);
or U2577 (N_2577,N_1475,N_1941);
nand U2578 (N_2578,N_1865,N_1874);
nor U2579 (N_2579,N_1559,N_1761);
and U2580 (N_2580,N_1630,N_1073);
or U2581 (N_2581,N_1948,N_1597);
or U2582 (N_2582,N_1207,N_1200);
nand U2583 (N_2583,N_1755,N_1109);
and U2584 (N_2584,N_1515,N_1173);
nor U2585 (N_2585,N_1358,N_1370);
xor U2586 (N_2586,N_1301,N_1921);
nand U2587 (N_2587,N_1257,N_1175);
or U2588 (N_2588,N_1684,N_1629);
nand U2589 (N_2589,N_1464,N_1050);
nand U2590 (N_2590,N_1161,N_1286);
nor U2591 (N_2591,N_1025,N_1511);
xnor U2592 (N_2592,N_1177,N_1780);
and U2593 (N_2593,N_1127,N_1037);
or U2594 (N_2594,N_1655,N_1665);
nand U2595 (N_2595,N_1889,N_1487);
nor U2596 (N_2596,N_1787,N_1241);
or U2597 (N_2597,N_1820,N_1851);
or U2598 (N_2598,N_1404,N_1437);
or U2599 (N_2599,N_1737,N_1525);
nand U2600 (N_2600,N_1406,N_1396);
and U2601 (N_2601,N_1453,N_1753);
and U2602 (N_2602,N_1173,N_1091);
and U2603 (N_2603,N_1659,N_1445);
nor U2604 (N_2604,N_1349,N_1109);
and U2605 (N_2605,N_1204,N_1746);
or U2606 (N_2606,N_1090,N_1802);
or U2607 (N_2607,N_1988,N_1877);
nor U2608 (N_2608,N_1361,N_1751);
nor U2609 (N_2609,N_1669,N_1292);
nor U2610 (N_2610,N_1613,N_1256);
nand U2611 (N_2611,N_1918,N_1085);
or U2612 (N_2612,N_1488,N_1179);
or U2613 (N_2613,N_1907,N_1703);
nor U2614 (N_2614,N_1475,N_1282);
nor U2615 (N_2615,N_1756,N_1189);
or U2616 (N_2616,N_1950,N_1522);
nand U2617 (N_2617,N_1530,N_1683);
nand U2618 (N_2618,N_1205,N_1038);
nor U2619 (N_2619,N_1294,N_1409);
nand U2620 (N_2620,N_1960,N_1796);
nor U2621 (N_2621,N_1259,N_1732);
nand U2622 (N_2622,N_1339,N_1898);
nand U2623 (N_2623,N_1701,N_1673);
or U2624 (N_2624,N_1890,N_1941);
and U2625 (N_2625,N_1775,N_1851);
xor U2626 (N_2626,N_1749,N_1354);
nor U2627 (N_2627,N_1050,N_1822);
nand U2628 (N_2628,N_1564,N_1805);
nor U2629 (N_2629,N_1747,N_1314);
and U2630 (N_2630,N_1137,N_1063);
or U2631 (N_2631,N_1598,N_1798);
nor U2632 (N_2632,N_1453,N_1794);
or U2633 (N_2633,N_1850,N_1932);
nand U2634 (N_2634,N_1242,N_1954);
nor U2635 (N_2635,N_1958,N_1661);
xnor U2636 (N_2636,N_1562,N_1786);
xnor U2637 (N_2637,N_1724,N_1296);
and U2638 (N_2638,N_1219,N_1342);
or U2639 (N_2639,N_1729,N_1275);
nor U2640 (N_2640,N_1545,N_1346);
nand U2641 (N_2641,N_1125,N_1068);
nand U2642 (N_2642,N_1872,N_1238);
and U2643 (N_2643,N_1443,N_1159);
nand U2644 (N_2644,N_1972,N_1749);
nand U2645 (N_2645,N_1156,N_1280);
nor U2646 (N_2646,N_1634,N_1566);
or U2647 (N_2647,N_1653,N_1606);
nor U2648 (N_2648,N_1950,N_1516);
nor U2649 (N_2649,N_1053,N_1912);
nand U2650 (N_2650,N_1103,N_1525);
xor U2651 (N_2651,N_1890,N_1610);
nand U2652 (N_2652,N_1432,N_1223);
nor U2653 (N_2653,N_1823,N_1181);
nand U2654 (N_2654,N_1053,N_1395);
nand U2655 (N_2655,N_1578,N_1257);
xnor U2656 (N_2656,N_1019,N_1512);
or U2657 (N_2657,N_1611,N_1652);
nor U2658 (N_2658,N_1923,N_1388);
and U2659 (N_2659,N_1660,N_1939);
and U2660 (N_2660,N_1158,N_1233);
xnor U2661 (N_2661,N_1265,N_1959);
or U2662 (N_2662,N_1848,N_1453);
nor U2663 (N_2663,N_1408,N_1758);
or U2664 (N_2664,N_1807,N_1736);
nand U2665 (N_2665,N_1785,N_1597);
and U2666 (N_2666,N_1096,N_1677);
or U2667 (N_2667,N_1817,N_1641);
xnor U2668 (N_2668,N_1582,N_1781);
nand U2669 (N_2669,N_1105,N_1825);
or U2670 (N_2670,N_1666,N_1636);
and U2671 (N_2671,N_1433,N_1924);
nor U2672 (N_2672,N_1416,N_1170);
and U2673 (N_2673,N_1584,N_1916);
xnor U2674 (N_2674,N_1496,N_1633);
or U2675 (N_2675,N_1004,N_1059);
nor U2676 (N_2676,N_1042,N_1939);
or U2677 (N_2677,N_1870,N_1932);
or U2678 (N_2678,N_1065,N_1507);
nand U2679 (N_2679,N_1507,N_1593);
or U2680 (N_2680,N_1800,N_1704);
nand U2681 (N_2681,N_1207,N_1457);
or U2682 (N_2682,N_1985,N_1703);
nand U2683 (N_2683,N_1675,N_1900);
and U2684 (N_2684,N_1603,N_1465);
and U2685 (N_2685,N_1349,N_1508);
or U2686 (N_2686,N_1816,N_1809);
or U2687 (N_2687,N_1417,N_1451);
nand U2688 (N_2688,N_1110,N_1627);
nor U2689 (N_2689,N_1061,N_1316);
or U2690 (N_2690,N_1167,N_1063);
nand U2691 (N_2691,N_1348,N_1717);
xnor U2692 (N_2692,N_1676,N_1893);
xor U2693 (N_2693,N_1130,N_1496);
or U2694 (N_2694,N_1056,N_1638);
nand U2695 (N_2695,N_1127,N_1753);
nand U2696 (N_2696,N_1012,N_1907);
and U2697 (N_2697,N_1301,N_1856);
xor U2698 (N_2698,N_1768,N_1076);
nor U2699 (N_2699,N_1851,N_1661);
nor U2700 (N_2700,N_1083,N_1057);
nor U2701 (N_2701,N_1694,N_1464);
nand U2702 (N_2702,N_1589,N_1619);
nand U2703 (N_2703,N_1079,N_1320);
nor U2704 (N_2704,N_1516,N_1999);
or U2705 (N_2705,N_1260,N_1067);
nor U2706 (N_2706,N_1485,N_1963);
or U2707 (N_2707,N_1650,N_1738);
nand U2708 (N_2708,N_1534,N_1159);
nand U2709 (N_2709,N_1136,N_1995);
or U2710 (N_2710,N_1042,N_1690);
or U2711 (N_2711,N_1066,N_1008);
or U2712 (N_2712,N_1624,N_1580);
xnor U2713 (N_2713,N_1763,N_1959);
or U2714 (N_2714,N_1761,N_1805);
nand U2715 (N_2715,N_1869,N_1817);
and U2716 (N_2716,N_1323,N_1179);
and U2717 (N_2717,N_1125,N_1815);
and U2718 (N_2718,N_1588,N_1166);
nand U2719 (N_2719,N_1108,N_1020);
nor U2720 (N_2720,N_1858,N_1619);
or U2721 (N_2721,N_1674,N_1486);
and U2722 (N_2722,N_1852,N_1774);
nand U2723 (N_2723,N_1831,N_1094);
and U2724 (N_2724,N_1995,N_1363);
nand U2725 (N_2725,N_1634,N_1365);
nand U2726 (N_2726,N_1617,N_1298);
or U2727 (N_2727,N_1762,N_1679);
or U2728 (N_2728,N_1989,N_1715);
or U2729 (N_2729,N_1212,N_1616);
nand U2730 (N_2730,N_1496,N_1978);
or U2731 (N_2731,N_1680,N_1052);
and U2732 (N_2732,N_1213,N_1183);
or U2733 (N_2733,N_1756,N_1864);
nand U2734 (N_2734,N_1015,N_1710);
nand U2735 (N_2735,N_1090,N_1621);
xor U2736 (N_2736,N_1003,N_1460);
and U2737 (N_2737,N_1915,N_1185);
or U2738 (N_2738,N_1829,N_1714);
nor U2739 (N_2739,N_1489,N_1705);
nor U2740 (N_2740,N_1756,N_1226);
or U2741 (N_2741,N_1030,N_1766);
nand U2742 (N_2742,N_1364,N_1551);
or U2743 (N_2743,N_1901,N_1849);
or U2744 (N_2744,N_1082,N_1317);
nor U2745 (N_2745,N_1421,N_1088);
nor U2746 (N_2746,N_1134,N_1429);
and U2747 (N_2747,N_1519,N_1532);
nor U2748 (N_2748,N_1220,N_1024);
nor U2749 (N_2749,N_1211,N_1207);
xor U2750 (N_2750,N_1723,N_1275);
and U2751 (N_2751,N_1935,N_1081);
and U2752 (N_2752,N_1484,N_1859);
and U2753 (N_2753,N_1758,N_1947);
nor U2754 (N_2754,N_1242,N_1760);
or U2755 (N_2755,N_1492,N_1784);
and U2756 (N_2756,N_1476,N_1507);
nand U2757 (N_2757,N_1550,N_1476);
nor U2758 (N_2758,N_1876,N_1682);
xnor U2759 (N_2759,N_1711,N_1535);
nand U2760 (N_2760,N_1787,N_1290);
nor U2761 (N_2761,N_1644,N_1055);
or U2762 (N_2762,N_1832,N_1239);
xnor U2763 (N_2763,N_1968,N_1037);
or U2764 (N_2764,N_1174,N_1547);
nor U2765 (N_2765,N_1765,N_1330);
nand U2766 (N_2766,N_1705,N_1023);
or U2767 (N_2767,N_1135,N_1151);
nor U2768 (N_2768,N_1087,N_1555);
and U2769 (N_2769,N_1018,N_1726);
or U2770 (N_2770,N_1958,N_1485);
or U2771 (N_2771,N_1944,N_1794);
xor U2772 (N_2772,N_1438,N_1481);
nor U2773 (N_2773,N_1600,N_1745);
or U2774 (N_2774,N_1815,N_1984);
and U2775 (N_2775,N_1054,N_1311);
and U2776 (N_2776,N_1155,N_1913);
nor U2777 (N_2777,N_1385,N_1739);
nand U2778 (N_2778,N_1363,N_1906);
and U2779 (N_2779,N_1026,N_1878);
and U2780 (N_2780,N_1044,N_1909);
nand U2781 (N_2781,N_1336,N_1016);
or U2782 (N_2782,N_1341,N_1120);
nand U2783 (N_2783,N_1300,N_1358);
nor U2784 (N_2784,N_1108,N_1366);
nor U2785 (N_2785,N_1153,N_1676);
nand U2786 (N_2786,N_1471,N_1519);
nand U2787 (N_2787,N_1844,N_1539);
nand U2788 (N_2788,N_1078,N_1936);
and U2789 (N_2789,N_1771,N_1127);
nor U2790 (N_2790,N_1241,N_1410);
and U2791 (N_2791,N_1151,N_1307);
and U2792 (N_2792,N_1405,N_1566);
and U2793 (N_2793,N_1144,N_1130);
nor U2794 (N_2794,N_1967,N_1963);
nor U2795 (N_2795,N_1989,N_1646);
xnor U2796 (N_2796,N_1777,N_1453);
or U2797 (N_2797,N_1697,N_1203);
xnor U2798 (N_2798,N_1913,N_1343);
or U2799 (N_2799,N_1218,N_1943);
nand U2800 (N_2800,N_1478,N_1838);
nand U2801 (N_2801,N_1206,N_1506);
nand U2802 (N_2802,N_1059,N_1944);
nor U2803 (N_2803,N_1589,N_1671);
nor U2804 (N_2804,N_1058,N_1097);
or U2805 (N_2805,N_1805,N_1006);
or U2806 (N_2806,N_1273,N_1466);
nand U2807 (N_2807,N_1675,N_1865);
or U2808 (N_2808,N_1345,N_1117);
or U2809 (N_2809,N_1922,N_1582);
or U2810 (N_2810,N_1771,N_1180);
nor U2811 (N_2811,N_1734,N_1688);
nand U2812 (N_2812,N_1703,N_1547);
nand U2813 (N_2813,N_1062,N_1747);
nand U2814 (N_2814,N_1483,N_1599);
or U2815 (N_2815,N_1097,N_1506);
nor U2816 (N_2816,N_1226,N_1267);
xor U2817 (N_2817,N_1941,N_1384);
nand U2818 (N_2818,N_1755,N_1146);
or U2819 (N_2819,N_1124,N_1238);
or U2820 (N_2820,N_1870,N_1175);
or U2821 (N_2821,N_1787,N_1160);
nand U2822 (N_2822,N_1479,N_1556);
nor U2823 (N_2823,N_1866,N_1079);
nand U2824 (N_2824,N_1140,N_1388);
or U2825 (N_2825,N_1139,N_1999);
nand U2826 (N_2826,N_1134,N_1463);
nand U2827 (N_2827,N_1267,N_1565);
nor U2828 (N_2828,N_1971,N_1524);
and U2829 (N_2829,N_1417,N_1616);
nand U2830 (N_2830,N_1424,N_1504);
or U2831 (N_2831,N_1360,N_1585);
nor U2832 (N_2832,N_1310,N_1683);
and U2833 (N_2833,N_1278,N_1153);
or U2834 (N_2834,N_1281,N_1942);
nand U2835 (N_2835,N_1087,N_1813);
nor U2836 (N_2836,N_1910,N_1282);
and U2837 (N_2837,N_1215,N_1366);
nand U2838 (N_2838,N_1949,N_1707);
and U2839 (N_2839,N_1516,N_1196);
or U2840 (N_2840,N_1587,N_1730);
and U2841 (N_2841,N_1746,N_1636);
or U2842 (N_2842,N_1151,N_1154);
or U2843 (N_2843,N_1098,N_1058);
and U2844 (N_2844,N_1233,N_1131);
nor U2845 (N_2845,N_1606,N_1357);
nor U2846 (N_2846,N_1728,N_1745);
and U2847 (N_2847,N_1347,N_1795);
and U2848 (N_2848,N_1657,N_1104);
nand U2849 (N_2849,N_1108,N_1992);
or U2850 (N_2850,N_1013,N_1814);
nor U2851 (N_2851,N_1661,N_1180);
and U2852 (N_2852,N_1144,N_1719);
or U2853 (N_2853,N_1736,N_1015);
nand U2854 (N_2854,N_1593,N_1735);
nand U2855 (N_2855,N_1120,N_1913);
or U2856 (N_2856,N_1488,N_1375);
nor U2857 (N_2857,N_1638,N_1305);
nand U2858 (N_2858,N_1713,N_1735);
nor U2859 (N_2859,N_1465,N_1788);
or U2860 (N_2860,N_1818,N_1281);
or U2861 (N_2861,N_1087,N_1495);
and U2862 (N_2862,N_1397,N_1756);
or U2863 (N_2863,N_1972,N_1411);
nor U2864 (N_2864,N_1169,N_1685);
nand U2865 (N_2865,N_1537,N_1945);
and U2866 (N_2866,N_1195,N_1596);
or U2867 (N_2867,N_1083,N_1228);
nor U2868 (N_2868,N_1493,N_1076);
nand U2869 (N_2869,N_1898,N_1515);
nand U2870 (N_2870,N_1722,N_1389);
and U2871 (N_2871,N_1178,N_1557);
and U2872 (N_2872,N_1951,N_1143);
or U2873 (N_2873,N_1122,N_1295);
and U2874 (N_2874,N_1725,N_1284);
or U2875 (N_2875,N_1790,N_1128);
nor U2876 (N_2876,N_1970,N_1801);
or U2877 (N_2877,N_1461,N_1712);
nor U2878 (N_2878,N_1869,N_1999);
or U2879 (N_2879,N_1762,N_1648);
nor U2880 (N_2880,N_1421,N_1342);
and U2881 (N_2881,N_1049,N_1195);
or U2882 (N_2882,N_1908,N_1300);
xor U2883 (N_2883,N_1527,N_1269);
and U2884 (N_2884,N_1035,N_1736);
and U2885 (N_2885,N_1439,N_1230);
or U2886 (N_2886,N_1679,N_1002);
nor U2887 (N_2887,N_1607,N_1159);
nor U2888 (N_2888,N_1025,N_1001);
or U2889 (N_2889,N_1581,N_1220);
nor U2890 (N_2890,N_1043,N_1006);
xor U2891 (N_2891,N_1096,N_1561);
and U2892 (N_2892,N_1519,N_1293);
and U2893 (N_2893,N_1228,N_1539);
nor U2894 (N_2894,N_1497,N_1592);
and U2895 (N_2895,N_1142,N_1211);
or U2896 (N_2896,N_1944,N_1961);
nand U2897 (N_2897,N_1170,N_1156);
nand U2898 (N_2898,N_1766,N_1492);
xor U2899 (N_2899,N_1833,N_1794);
or U2900 (N_2900,N_1656,N_1104);
nor U2901 (N_2901,N_1295,N_1681);
nor U2902 (N_2902,N_1765,N_1814);
xnor U2903 (N_2903,N_1237,N_1148);
nor U2904 (N_2904,N_1725,N_1374);
xor U2905 (N_2905,N_1566,N_1715);
and U2906 (N_2906,N_1750,N_1655);
nand U2907 (N_2907,N_1768,N_1206);
and U2908 (N_2908,N_1794,N_1688);
nand U2909 (N_2909,N_1151,N_1605);
and U2910 (N_2910,N_1902,N_1933);
and U2911 (N_2911,N_1371,N_1097);
nand U2912 (N_2912,N_1549,N_1685);
nand U2913 (N_2913,N_1602,N_1535);
nand U2914 (N_2914,N_1472,N_1360);
nor U2915 (N_2915,N_1376,N_1168);
nand U2916 (N_2916,N_1977,N_1600);
nand U2917 (N_2917,N_1224,N_1482);
and U2918 (N_2918,N_1198,N_1465);
nand U2919 (N_2919,N_1439,N_1151);
or U2920 (N_2920,N_1932,N_1756);
and U2921 (N_2921,N_1773,N_1828);
and U2922 (N_2922,N_1729,N_1973);
nor U2923 (N_2923,N_1663,N_1022);
nor U2924 (N_2924,N_1705,N_1336);
nor U2925 (N_2925,N_1963,N_1764);
nand U2926 (N_2926,N_1378,N_1805);
and U2927 (N_2927,N_1187,N_1875);
nor U2928 (N_2928,N_1149,N_1488);
or U2929 (N_2929,N_1439,N_1835);
or U2930 (N_2930,N_1015,N_1409);
nand U2931 (N_2931,N_1924,N_1106);
nor U2932 (N_2932,N_1833,N_1104);
nor U2933 (N_2933,N_1316,N_1853);
and U2934 (N_2934,N_1595,N_1056);
or U2935 (N_2935,N_1838,N_1651);
or U2936 (N_2936,N_1936,N_1981);
and U2937 (N_2937,N_1030,N_1797);
and U2938 (N_2938,N_1781,N_1123);
or U2939 (N_2939,N_1424,N_1213);
and U2940 (N_2940,N_1449,N_1981);
xor U2941 (N_2941,N_1509,N_1897);
nand U2942 (N_2942,N_1615,N_1045);
and U2943 (N_2943,N_1455,N_1521);
nand U2944 (N_2944,N_1217,N_1210);
nor U2945 (N_2945,N_1098,N_1523);
and U2946 (N_2946,N_1760,N_1248);
nor U2947 (N_2947,N_1958,N_1030);
nand U2948 (N_2948,N_1784,N_1601);
and U2949 (N_2949,N_1273,N_1138);
or U2950 (N_2950,N_1039,N_1808);
nor U2951 (N_2951,N_1586,N_1939);
or U2952 (N_2952,N_1240,N_1164);
nand U2953 (N_2953,N_1508,N_1222);
nand U2954 (N_2954,N_1737,N_1843);
and U2955 (N_2955,N_1553,N_1340);
and U2956 (N_2956,N_1178,N_1188);
and U2957 (N_2957,N_1777,N_1348);
nor U2958 (N_2958,N_1731,N_1608);
xor U2959 (N_2959,N_1044,N_1691);
or U2960 (N_2960,N_1764,N_1650);
and U2961 (N_2961,N_1699,N_1784);
xor U2962 (N_2962,N_1296,N_1192);
or U2963 (N_2963,N_1736,N_1611);
nor U2964 (N_2964,N_1151,N_1101);
nand U2965 (N_2965,N_1450,N_1998);
nor U2966 (N_2966,N_1840,N_1700);
or U2967 (N_2967,N_1545,N_1719);
xnor U2968 (N_2968,N_1961,N_1616);
xor U2969 (N_2969,N_1550,N_1186);
nand U2970 (N_2970,N_1622,N_1472);
xnor U2971 (N_2971,N_1251,N_1191);
nand U2972 (N_2972,N_1578,N_1605);
nor U2973 (N_2973,N_1751,N_1735);
nand U2974 (N_2974,N_1271,N_1020);
nand U2975 (N_2975,N_1459,N_1084);
or U2976 (N_2976,N_1634,N_1172);
nor U2977 (N_2977,N_1915,N_1703);
nor U2978 (N_2978,N_1345,N_1176);
and U2979 (N_2979,N_1673,N_1212);
nor U2980 (N_2980,N_1198,N_1277);
nor U2981 (N_2981,N_1466,N_1416);
or U2982 (N_2982,N_1324,N_1407);
nor U2983 (N_2983,N_1768,N_1367);
and U2984 (N_2984,N_1368,N_1534);
or U2985 (N_2985,N_1765,N_1894);
or U2986 (N_2986,N_1040,N_1404);
and U2987 (N_2987,N_1861,N_1853);
or U2988 (N_2988,N_1893,N_1540);
nand U2989 (N_2989,N_1278,N_1890);
or U2990 (N_2990,N_1984,N_1792);
nor U2991 (N_2991,N_1883,N_1829);
xnor U2992 (N_2992,N_1754,N_1138);
nor U2993 (N_2993,N_1898,N_1458);
and U2994 (N_2994,N_1752,N_1047);
or U2995 (N_2995,N_1798,N_1878);
nor U2996 (N_2996,N_1560,N_1474);
nor U2997 (N_2997,N_1444,N_1954);
nand U2998 (N_2998,N_1603,N_1919);
and U2999 (N_2999,N_1275,N_1327);
nor UO_0 (O_0,N_2053,N_2102);
and UO_1 (O_1,N_2842,N_2177);
and UO_2 (O_2,N_2270,N_2011);
nor UO_3 (O_3,N_2614,N_2736);
nor UO_4 (O_4,N_2310,N_2796);
nor UO_5 (O_5,N_2045,N_2859);
xor UO_6 (O_6,N_2056,N_2730);
and UO_7 (O_7,N_2823,N_2199);
nand UO_8 (O_8,N_2950,N_2575);
or UO_9 (O_9,N_2767,N_2111);
nand UO_10 (O_10,N_2794,N_2117);
or UO_11 (O_11,N_2927,N_2457);
nor UO_12 (O_12,N_2313,N_2151);
and UO_13 (O_13,N_2472,N_2863);
or UO_14 (O_14,N_2129,N_2670);
xnor UO_15 (O_15,N_2729,N_2816);
nor UO_16 (O_16,N_2822,N_2080);
xor UO_17 (O_17,N_2263,N_2790);
and UO_18 (O_18,N_2275,N_2027);
nor UO_19 (O_19,N_2081,N_2557);
and UO_20 (O_20,N_2001,N_2946);
and UO_21 (O_21,N_2008,N_2175);
nand UO_22 (O_22,N_2540,N_2188);
nor UO_23 (O_23,N_2029,N_2991);
nand UO_24 (O_24,N_2775,N_2022);
and UO_25 (O_25,N_2236,N_2641);
nand UO_26 (O_26,N_2414,N_2014);
nor UO_27 (O_27,N_2268,N_2259);
nand UO_28 (O_28,N_2776,N_2905);
and UO_29 (O_29,N_2615,N_2444);
and UO_30 (O_30,N_2307,N_2176);
and UO_31 (O_31,N_2826,N_2301);
nand UO_32 (O_32,N_2141,N_2123);
xnor UO_33 (O_33,N_2099,N_2560);
or UO_34 (O_34,N_2443,N_2198);
or UO_35 (O_35,N_2207,N_2544);
nor UO_36 (O_36,N_2972,N_2922);
nor UO_37 (O_37,N_2034,N_2913);
nand UO_38 (O_38,N_2007,N_2891);
nand UO_39 (O_39,N_2992,N_2574);
nand UO_40 (O_40,N_2719,N_2164);
nand UO_41 (O_41,N_2067,N_2205);
nor UO_42 (O_42,N_2391,N_2282);
or UO_43 (O_43,N_2356,N_2539);
xor UO_44 (O_44,N_2172,N_2203);
or UO_45 (O_45,N_2181,N_2358);
and UO_46 (O_46,N_2287,N_2785);
and UO_47 (O_47,N_2269,N_2572);
nor UO_48 (O_48,N_2653,N_2031);
and UO_49 (O_49,N_2168,N_2348);
nand UO_50 (O_50,N_2505,N_2622);
and UO_51 (O_51,N_2824,N_2144);
xor UO_52 (O_52,N_2097,N_2920);
nor UO_53 (O_53,N_2353,N_2724);
and UO_54 (O_54,N_2036,N_2570);
nor UO_55 (O_55,N_2299,N_2784);
and UO_56 (O_56,N_2229,N_2910);
nand UO_57 (O_57,N_2537,N_2284);
nand UO_58 (O_58,N_2618,N_2437);
or UO_59 (O_59,N_2947,N_2616);
or UO_60 (O_60,N_2213,N_2698);
nand UO_61 (O_61,N_2798,N_2037);
and UO_62 (O_62,N_2204,N_2899);
nor UO_63 (O_63,N_2739,N_2028);
or UO_64 (O_64,N_2835,N_2791);
nand UO_65 (O_65,N_2265,N_2377);
nor UO_66 (O_66,N_2302,N_2490);
nor UO_67 (O_67,N_2253,N_2825);
or UO_68 (O_68,N_2843,N_2743);
nor UO_69 (O_69,N_2128,N_2832);
nand UO_70 (O_70,N_2297,N_2059);
nor UO_71 (O_71,N_2362,N_2726);
nor UO_72 (O_72,N_2467,N_2535);
nor UO_73 (O_73,N_2054,N_2656);
nand UO_74 (O_74,N_2163,N_2644);
nor UO_75 (O_75,N_2751,N_2183);
nand UO_76 (O_76,N_2066,N_2600);
or UO_77 (O_77,N_2602,N_2519);
nor UO_78 (O_78,N_2318,N_2432);
xnor UO_79 (O_79,N_2161,N_2323);
xnor UO_80 (O_80,N_2897,N_2247);
nor UO_81 (O_81,N_2924,N_2710);
nor UO_82 (O_82,N_2235,N_2191);
or UO_83 (O_83,N_2871,N_2073);
and UO_84 (O_84,N_2065,N_2024);
xor UO_85 (O_85,N_2032,N_2898);
nand UO_86 (O_86,N_2674,N_2869);
or UO_87 (O_87,N_2981,N_2987);
nor UO_88 (O_88,N_2581,N_2304);
or UO_89 (O_89,N_2495,N_2217);
or UO_90 (O_90,N_2320,N_2885);
or UO_91 (O_91,N_2465,N_2846);
and UO_92 (O_92,N_2119,N_2760);
or UO_93 (O_93,N_2521,N_2441);
or UO_94 (O_94,N_2888,N_2608);
and UO_95 (O_95,N_2526,N_2691);
or UO_96 (O_96,N_2112,N_2699);
and UO_97 (O_97,N_2094,N_2901);
and UO_98 (O_98,N_2599,N_2558);
xor UO_99 (O_99,N_2973,N_2951);
and UO_100 (O_100,N_2245,N_2139);
and UO_101 (O_101,N_2484,N_2255);
and UO_102 (O_102,N_2440,N_2470);
nor UO_103 (O_103,N_2393,N_2604);
nand UO_104 (O_104,N_2435,N_2718);
nor UO_105 (O_105,N_2492,N_2254);
and UO_106 (O_106,N_2665,N_2930);
nand UO_107 (O_107,N_2769,N_2895);
nand UO_108 (O_108,N_2140,N_2873);
nor UO_109 (O_109,N_2912,N_2821);
and UO_110 (O_110,N_2087,N_2773);
and UO_111 (O_111,N_2564,N_2157);
nand UO_112 (O_112,N_2697,N_2208);
nor UO_113 (O_113,N_2116,N_2580);
xnor UO_114 (O_114,N_2293,N_2146);
nand UO_115 (O_115,N_2713,N_2419);
nand UO_116 (O_116,N_2830,N_2148);
and UO_117 (O_117,N_2850,N_2516);
or UO_118 (O_118,N_2635,N_2149);
xor UO_119 (O_119,N_2778,N_2279);
nor UO_120 (O_120,N_2807,N_2364);
or UO_121 (O_121,N_2145,N_2782);
nand UO_122 (O_122,N_2306,N_2433);
and UO_123 (O_123,N_2224,N_2324);
or UO_124 (O_124,N_2226,N_2219);
or UO_125 (O_125,N_2048,N_2035);
nand UO_126 (O_126,N_2372,N_2956);
and UO_127 (O_127,N_2496,N_2086);
nor UO_128 (O_128,N_2343,N_2668);
or UO_129 (O_129,N_2277,N_2789);
and UO_130 (O_130,N_2130,N_2940);
or UO_131 (O_131,N_2855,N_2637);
nand UO_132 (O_132,N_2013,N_2507);
and UO_133 (O_133,N_2969,N_2244);
nand UO_134 (O_134,N_2480,N_2765);
and UO_135 (O_135,N_2352,N_2742);
xor UO_136 (O_136,N_2017,N_2091);
or UO_137 (O_137,N_2122,N_2663);
or UO_138 (O_138,N_2043,N_2095);
nand UO_139 (O_139,N_2737,N_2988);
xnor UO_140 (O_140,N_2190,N_2395);
or UO_141 (O_141,N_2999,N_2209);
xnor UO_142 (O_142,N_2605,N_2997);
nand UO_143 (O_143,N_2196,N_2169);
nor UO_144 (O_144,N_2682,N_2120);
and UO_145 (O_145,N_2453,N_2162);
nand UO_146 (O_146,N_2904,N_2316);
or UO_147 (O_147,N_2068,N_2603);
xnor UO_148 (O_148,N_2945,N_2954);
nand UO_149 (O_149,N_2514,N_2482);
and UO_150 (O_150,N_2349,N_2555);
nor UO_151 (O_151,N_2382,N_2373);
and UO_152 (O_152,N_2648,N_2702);
or UO_153 (O_153,N_2587,N_2367);
or UO_154 (O_154,N_2407,N_2928);
nor UO_155 (O_155,N_2359,N_2016);
nand UO_156 (O_156,N_2877,N_2308);
or UO_157 (O_157,N_2588,N_2549);
or UO_158 (O_158,N_2523,N_2985);
and UO_159 (O_159,N_2462,N_2642);
nor UO_160 (O_160,N_2839,N_2401);
nor UO_161 (O_161,N_2517,N_2792);
or UO_162 (O_162,N_2103,N_2357);
or UO_163 (O_163,N_2077,N_2533);
and UO_164 (O_164,N_2361,N_2733);
nor UO_165 (O_165,N_2178,N_2452);
xnor UO_166 (O_166,N_2390,N_2478);
nor UO_167 (O_167,N_2929,N_2469);
and UO_168 (O_168,N_2611,N_2124);
nor UO_169 (O_169,N_2400,N_2942);
or UO_170 (O_170,N_2044,N_2098);
or UO_171 (O_171,N_2914,N_2315);
nor UO_172 (O_172,N_2326,N_2613);
or UO_173 (O_173,N_2610,N_2970);
nand UO_174 (O_174,N_2143,N_2110);
or UO_175 (O_175,N_2980,N_2703);
nor UO_176 (O_176,N_2062,N_2201);
nor UO_177 (O_177,N_2200,N_2650);
xor UO_178 (O_178,N_2689,N_2513);
nor UO_179 (O_179,N_2880,N_2690);
xor UO_180 (O_180,N_2319,N_2220);
nor UO_181 (O_181,N_2089,N_2757);
nand UO_182 (O_182,N_2696,N_2429);
or UO_183 (O_183,N_2550,N_2184);
nand UO_184 (O_184,N_2300,N_2448);
nor UO_185 (O_185,N_2844,N_2944);
nor UO_186 (O_186,N_2768,N_2640);
nand UO_187 (O_187,N_2777,N_2607);
nor UO_188 (O_188,N_2061,N_2397);
and UO_189 (O_189,N_2771,N_2589);
nand UO_190 (O_190,N_2154,N_2601);
nor UO_191 (O_191,N_2214,N_2179);
nand UO_192 (O_192,N_2399,N_2055);
or UO_193 (O_193,N_2683,N_2242);
nand UO_194 (O_194,N_2366,N_2687);
and UO_195 (O_195,N_2879,N_2903);
and UO_196 (O_196,N_2447,N_2957);
nor UO_197 (O_197,N_2829,N_2340);
and UO_198 (O_198,N_2747,N_2814);
nand UO_199 (O_199,N_2772,N_2576);
and UO_200 (O_200,N_2501,N_2396);
nand UO_201 (O_201,N_2314,N_2979);
nand UO_202 (O_202,N_2609,N_2886);
nand UO_203 (O_203,N_2221,N_2723);
xor UO_204 (O_204,N_2210,N_2959);
nand UO_205 (O_205,N_2369,N_2009);
or UO_206 (O_206,N_2446,N_2436);
and UO_207 (O_207,N_2185,N_2819);
nor UO_208 (O_208,N_2639,N_2153);
nand UO_209 (O_209,N_2673,N_2398);
and UO_210 (O_210,N_2454,N_2960);
nor UO_211 (O_211,N_2976,N_2865);
or UO_212 (O_212,N_2541,N_2530);
nand UO_213 (O_213,N_2620,N_2797);
nand UO_214 (O_214,N_2837,N_2451);
nor UO_215 (O_215,N_2460,N_2425);
or UO_216 (O_216,N_2974,N_2659);
nand UO_217 (O_217,N_2971,N_2392);
nor UO_218 (O_218,N_2799,N_2346);
nor UO_219 (O_219,N_2800,N_2071);
nor UO_220 (O_220,N_2223,N_2355);
nor UO_221 (O_221,N_2118,N_2759);
or UO_222 (O_222,N_2231,N_2677);
nor UO_223 (O_223,N_2894,N_2882);
nor UO_224 (O_224,N_2627,N_2458);
nand UO_225 (O_225,N_2333,N_2344);
and UO_226 (O_226,N_2965,N_2388);
and UO_227 (O_227,N_2786,N_2327);
and UO_228 (O_228,N_2935,N_2847);
nand UO_229 (O_229,N_2473,N_2336);
and UO_230 (O_230,N_2335,N_2745);
nand UO_231 (O_231,N_2593,N_2638);
or UO_232 (O_232,N_2193,N_2774);
or UO_233 (O_233,N_2006,N_2735);
nand UO_234 (O_234,N_2686,N_2820);
and UO_235 (O_235,N_2375,N_2815);
nor UO_236 (O_236,N_2722,N_2173);
or UO_237 (O_237,N_2552,N_2019);
and UO_238 (O_238,N_2961,N_2252);
or UO_239 (O_239,N_2290,N_2415);
and UO_240 (O_240,N_2136,N_2967);
and UO_241 (O_241,N_2548,N_2249);
nor UO_242 (O_242,N_2101,N_2626);
and UO_243 (O_243,N_2590,N_2261);
nand UO_244 (O_244,N_2752,N_2438);
xnor UO_245 (O_245,N_2288,N_2192);
nor UO_246 (O_246,N_2278,N_2949);
and UO_247 (O_247,N_2694,N_2975);
nand UO_248 (O_248,N_2840,N_2916);
nand UO_249 (O_249,N_2070,N_2695);
nand UO_250 (O_250,N_2408,N_2413);
and UO_251 (O_251,N_2106,N_2571);
nor UO_252 (O_252,N_2936,N_2990);
nand UO_253 (O_253,N_2456,N_2232);
and UO_254 (O_254,N_2039,N_2932);
nand UO_255 (O_255,N_2506,N_2060);
xor UO_256 (O_256,N_2250,N_2502);
nand UO_257 (O_257,N_2966,N_2554);
or UO_258 (O_258,N_2371,N_2836);
or UO_259 (O_259,N_2281,N_2854);
nand UO_260 (O_260,N_2679,N_2421);
and UO_261 (O_261,N_2442,N_2239);
nor UO_262 (O_262,N_2933,N_2058);
xor UO_263 (O_263,N_2165,N_2069);
nand UO_264 (O_264,N_2260,N_2360);
and UO_265 (O_265,N_2510,N_2906);
nor UO_266 (O_266,N_2422,N_2150);
nand UO_267 (O_267,N_2160,N_2631);
xor UO_268 (O_268,N_2728,N_2449);
nand UO_269 (O_269,N_2685,N_2700);
and UO_270 (O_270,N_2624,N_2115);
or UO_271 (O_271,N_2487,N_2410);
nor UO_272 (O_272,N_2135,N_2938);
or UO_273 (O_273,N_2579,N_2834);
or UO_274 (O_274,N_2475,N_2525);
nor UO_275 (O_275,N_2872,N_2108);
and UO_276 (O_276,N_2766,N_2701);
and UO_277 (O_277,N_2787,N_2114);
nand UO_278 (O_278,N_2127,N_2113);
nand UO_279 (O_279,N_2955,N_2021);
and UO_280 (O_280,N_2295,N_2707);
nand UO_281 (O_281,N_2584,N_2381);
xnor UO_282 (O_282,N_2547,N_2020);
xnor UO_283 (O_283,N_2345,N_2328);
nand UO_284 (O_284,N_2218,N_2948);
nor UO_285 (O_285,N_2902,N_2132);
nand UO_286 (O_286,N_2347,N_2100);
nand UO_287 (O_287,N_2134,N_2889);
xor UO_288 (O_288,N_2018,N_2234);
nor UO_289 (O_289,N_2420,N_2669);
nor UO_290 (O_290,N_2222,N_2937);
and UO_291 (O_291,N_2727,N_2380);
nand UO_292 (O_292,N_2817,N_2104);
and UO_293 (O_293,N_2636,N_2860);
or UO_294 (O_294,N_2900,N_2002);
and UO_295 (O_295,N_2802,N_2005);
or UO_296 (O_296,N_2658,N_2738);
nand UO_297 (O_297,N_2082,N_2803);
nor UO_298 (O_298,N_2655,N_2862);
and UO_299 (O_299,N_2121,N_2334);
or UO_300 (O_300,N_2908,N_2468);
and UO_301 (O_301,N_2418,N_2064);
nor UO_302 (O_302,N_2384,N_2717);
or UO_303 (O_303,N_2272,N_2493);
nand UO_304 (O_304,N_2878,N_2330);
and UO_305 (O_305,N_2994,N_2385);
nand UO_306 (O_306,N_2206,N_2654);
nand UO_307 (O_307,N_2194,N_2864);
nor UO_308 (O_308,N_2479,N_2676);
nor UO_309 (O_309,N_2688,N_2455);
or UO_310 (O_310,N_2856,N_2296);
xnor UO_311 (O_311,N_2088,N_2755);
nand UO_312 (O_312,N_2374,N_2074);
and UO_313 (O_313,N_2754,N_2015);
nor UO_314 (O_314,N_2405,N_2424);
and UO_315 (O_315,N_2305,N_2657);
or UO_316 (O_316,N_2241,N_2619);
and UO_317 (O_317,N_2746,N_2567);
and UO_318 (O_318,N_2569,N_2057);
and UO_319 (O_319,N_2716,N_2285);
or UO_320 (O_320,N_2998,N_2033);
and UO_321 (O_321,N_2753,N_2875);
nand UO_322 (O_322,N_2858,N_2133);
nor UO_323 (O_323,N_2725,N_2561);
nand UO_324 (O_324,N_2294,N_2881);
nor UO_325 (O_325,N_2818,N_2573);
and UO_326 (O_326,N_2508,N_2474);
nor UO_327 (O_327,N_2887,N_2721);
nor UO_328 (O_328,N_2923,N_2651);
and UO_329 (O_329,N_2926,N_2711);
nor UO_330 (O_330,N_2138,N_2159);
or UO_331 (O_331,N_2562,N_2617);
or UO_332 (O_332,N_2485,N_2341);
or UO_333 (O_333,N_2801,N_2404);
nor UO_334 (O_334,N_2267,N_2762);
or UO_335 (O_335,N_2488,N_2262);
and UO_336 (O_336,N_2152,N_2430);
or UO_337 (O_337,N_2233,N_2354);
and UO_338 (O_338,N_2363,N_2325);
nand UO_339 (O_339,N_2494,N_2406);
and UO_340 (O_340,N_2598,N_2147);
nand UO_341 (O_341,N_2941,N_2592);
and UO_342 (O_342,N_2383,N_2142);
and UO_343 (O_343,N_2459,N_2993);
or UO_344 (O_344,N_2779,N_2289);
nand UO_345 (O_345,N_2509,N_2411);
nor UO_346 (O_346,N_2156,N_2339);
xor UO_347 (O_347,N_2741,N_2565);
nor UO_348 (O_348,N_2909,N_2378);
or UO_349 (O_349,N_2257,N_2072);
nor UO_350 (O_350,N_2211,N_2292);
nor UO_351 (O_351,N_2632,N_2851);
nor UO_352 (O_352,N_2182,N_2026);
and UO_353 (O_353,N_2634,N_2389);
nand UO_354 (O_354,N_2666,N_2520);
nand UO_355 (O_355,N_2577,N_2680);
and UO_356 (O_356,N_2512,N_2596);
or UO_357 (O_357,N_2264,N_2431);
nor UO_358 (O_358,N_2471,N_2748);
or UO_359 (O_359,N_2804,N_2761);
nand UO_360 (O_360,N_2107,N_2416);
and UO_361 (O_361,N_2491,N_2866);
and UO_362 (O_362,N_2450,N_2498);
or UO_363 (O_363,N_2303,N_2857);
nand UO_364 (O_364,N_2712,N_2630);
nand UO_365 (O_365,N_2870,N_2096);
or UO_366 (O_366,N_2708,N_2042);
nor UO_367 (O_367,N_2931,N_2662);
nand UO_368 (O_368,N_2312,N_2125);
or UO_369 (O_369,N_2551,N_2370);
or UO_370 (O_370,N_2968,N_2628);
or UO_371 (O_371,N_2925,N_2329);
and UO_372 (O_372,N_2126,N_2237);
nand UO_373 (O_373,N_2781,N_2337);
nand UO_374 (O_374,N_2040,N_2228);
nor UO_375 (O_375,N_2311,N_2052);
nand UO_376 (O_376,N_2853,N_2041);
or UO_377 (O_377,N_2386,N_2246);
nand UO_378 (O_378,N_2652,N_2827);
and UO_379 (O_379,N_2633,N_2884);
nand UO_380 (O_380,N_2522,N_2828);
and UO_381 (O_381,N_2243,N_2672);
nand UO_382 (O_382,N_2000,N_2953);
xor UO_383 (O_383,N_2215,N_2813);
nor UO_384 (O_384,N_2795,N_2291);
or UO_385 (O_385,N_2595,N_2538);
nand UO_386 (O_386,N_2812,N_2883);
nor UO_387 (O_387,N_2003,N_2568);
or UO_388 (O_388,N_2952,N_2286);
and UO_389 (O_389,N_2780,N_2497);
or UO_390 (O_390,N_2518,N_2202);
or UO_391 (O_391,N_2322,N_2806);
and UO_392 (O_392,N_2376,N_2750);
and UO_393 (O_393,N_2280,N_2876);
and UO_394 (O_394,N_2225,N_2197);
nand UO_395 (O_395,N_2500,N_2692);
nor UO_396 (O_396,N_2483,N_2545);
nor UO_397 (O_397,N_2332,N_2943);
nor UO_398 (O_398,N_2216,N_2047);
nand UO_399 (O_399,N_2428,N_2092);
nor UO_400 (O_400,N_2678,N_2317);
and UO_401 (O_401,N_2531,N_2412);
nor UO_402 (O_402,N_2646,N_2030);
nor UO_403 (O_403,N_2180,N_2529);
nand UO_404 (O_404,N_2849,N_2230);
nor UO_405 (O_405,N_2271,N_2709);
nand UO_406 (O_406,N_2559,N_2907);
and UO_407 (O_407,N_2274,N_2995);
xor UO_408 (O_408,N_2417,N_2046);
and UO_409 (O_409,N_2321,N_2240);
nand UO_410 (O_410,N_2078,N_2740);
or UO_411 (O_411,N_2503,N_2038);
nor UO_412 (O_412,N_2423,N_2402);
or UO_413 (O_413,N_2667,N_2010);
xnor UO_414 (O_414,N_2583,N_2978);
nor UO_415 (O_415,N_2681,N_2984);
or UO_416 (O_416,N_2805,N_2977);
and UO_417 (O_417,N_2025,N_2958);
nand UO_418 (O_418,N_2623,N_2409);
nor UO_419 (O_419,N_2744,N_2527);
nand UO_420 (O_420,N_2170,N_2734);
nand UO_421 (O_421,N_2808,N_2063);
and UO_422 (O_422,N_2621,N_2461);
or UO_423 (O_423,N_2189,N_2477);
and UO_424 (O_424,N_2715,N_2764);
and UO_425 (O_425,N_2368,N_2660);
xor UO_426 (O_426,N_2464,N_2515);
or UO_427 (O_427,N_2732,N_2543);
and UO_428 (O_428,N_2331,N_2166);
nand UO_429 (O_429,N_2023,N_2963);
and UO_430 (O_430,N_2251,N_2075);
nor UO_431 (O_431,N_2171,N_2004);
nor UO_432 (O_432,N_2283,N_2258);
or UO_433 (O_433,N_2105,N_2664);
nor UO_434 (O_434,N_2591,N_2342);
and UO_435 (O_435,N_2051,N_2868);
nand UO_436 (O_436,N_2528,N_2788);
nor UO_437 (O_437,N_2706,N_2365);
xnor UO_438 (O_438,N_2606,N_2612);
and UO_439 (O_439,N_2050,N_2861);
nor UO_440 (O_440,N_2867,N_2594);
or UO_441 (O_441,N_2266,N_2542);
nand UO_442 (O_442,N_2445,N_2556);
nand UO_443 (O_443,N_2227,N_2532);
and UO_444 (O_444,N_2983,N_2167);
and UO_445 (O_445,N_2831,N_2643);
or UO_446 (O_446,N_2586,N_2704);
or UO_447 (O_447,N_2756,N_2084);
nand UO_448 (O_448,N_2845,N_2137);
xor UO_449 (O_449,N_2534,N_2298);
or UO_450 (O_450,N_2463,N_2109);
or UO_451 (O_451,N_2915,N_2212);
nor UO_452 (O_452,N_2749,N_2918);
nand UO_453 (O_453,N_2986,N_2705);
or UO_454 (O_454,N_2174,N_2645);
nand UO_455 (O_455,N_2770,N_2309);
or UO_456 (O_456,N_2186,N_2511);
nand UO_457 (O_457,N_2155,N_2809);
and UO_458 (O_458,N_2499,N_2890);
or UO_459 (O_459,N_2763,N_2076);
and UO_460 (O_460,N_2536,N_2675);
nor UO_461 (O_461,N_2841,N_2248);
and UO_462 (O_462,N_2671,N_2276);
or UO_463 (O_463,N_2350,N_2504);
nor UO_464 (O_464,N_2964,N_2434);
nand UO_465 (O_465,N_2939,N_2934);
and UO_466 (O_466,N_2982,N_2083);
and UO_467 (O_467,N_2090,N_2714);
or UO_468 (O_468,N_2093,N_2466);
nand UO_469 (O_469,N_2684,N_2919);
and UO_470 (O_470,N_2693,N_2811);
nand UO_471 (O_471,N_2578,N_2893);
xnor UO_472 (O_472,N_2758,N_2256);
or UO_473 (O_473,N_2892,N_2379);
nor UO_474 (O_474,N_2833,N_2848);
xor UO_475 (O_475,N_2486,N_2426);
or UO_476 (O_476,N_2489,N_2647);
nor UO_477 (O_477,N_2439,N_2351);
nand UO_478 (O_478,N_2852,N_2563);
xor UO_479 (O_479,N_2720,N_2012);
nand UO_480 (O_480,N_2585,N_2238);
nor UO_481 (O_481,N_2810,N_2195);
nand UO_482 (O_482,N_2566,N_2838);
and UO_483 (O_483,N_2989,N_2338);
or UO_484 (O_484,N_2629,N_2793);
nor UO_485 (O_485,N_2481,N_2476);
nand UO_486 (O_486,N_2273,N_2996);
nor UO_487 (O_487,N_2597,N_2783);
and UO_488 (O_488,N_2917,N_2427);
nor UO_489 (O_489,N_2079,N_2387);
or UO_490 (O_490,N_2187,N_2553);
or UO_491 (O_491,N_2085,N_2131);
and UO_492 (O_492,N_2625,N_2921);
nand UO_493 (O_493,N_2403,N_2546);
nand UO_494 (O_494,N_2394,N_2661);
nor UO_495 (O_495,N_2896,N_2582);
and UO_496 (O_496,N_2158,N_2524);
and UO_497 (O_497,N_2049,N_2911);
nor UO_498 (O_498,N_2649,N_2874);
and UO_499 (O_499,N_2731,N_2962);
endmodule