module basic_3000_30000_3500_25_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_757,In_2250);
xnor U1 (N_1,In_968,In_700);
and U2 (N_2,In_2414,In_1753);
nor U3 (N_3,In_1885,In_2962);
nand U4 (N_4,In_1303,In_231);
xor U5 (N_5,In_829,In_1049);
nor U6 (N_6,In_1427,In_2629);
nor U7 (N_7,In_2760,In_1412);
nor U8 (N_8,In_1369,In_2136);
and U9 (N_9,In_1139,In_891);
and U10 (N_10,In_2910,In_917);
nor U11 (N_11,In_1969,In_2905);
xnor U12 (N_12,In_2087,In_296);
or U13 (N_13,In_1506,In_2398);
nand U14 (N_14,In_1663,In_2065);
xor U15 (N_15,In_262,In_2954);
or U16 (N_16,In_1065,In_2953);
nand U17 (N_17,In_885,In_2188);
or U18 (N_18,In_1757,In_247);
and U19 (N_19,In_513,In_1224);
and U20 (N_20,In_168,In_651);
xnor U21 (N_21,In_59,In_2444);
and U22 (N_22,In_1936,In_1256);
xnor U23 (N_23,In_1615,In_1881);
and U24 (N_24,In_850,In_1105);
xnor U25 (N_25,In_2125,In_1522);
and U26 (N_26,In_1561,In_2082);
and U27 (N_27,In_2283,In_2);
nand U28 (N_28,In_684,In_268);
and U29 (N_29,In_1916,In_1542);
nand U30 (N_30,In_196,In_855);
and U31 (N_31,In_2940,In_1622);
nor U32 (N_32,In_2636,In_1212);
nor U33 (N_33,In_1767,In_2004);
and U34 (N_34,In_1651,In_2854);
nor U35 (N_35,In_1305,In_2086);
nand U36 (N_36,In_1203,In_665);
nand U37 (N_37,In_1094,In_324);
and U38 (N_38,In_400,In_1964);
nand U39 (N_39,In_449,In_1490);
nor U40 (N_40,In_531,In_1543);
and U41 (N_41,In_1196,In_2981);
nand U42 (N_42,In_1967,In_1457);
nor U43 (N_43,In_2064,In_24);
and U44 (N_44,In_2840,In_1314);
nor U45 (N_45,In_1980,In_1341);
or U46 (N_46,In_1052,In_1778);
or U47 (N_47,In_462,In_1416);
xnor U48 (N_48,In_1045,In_2624);
or U49 (N_49,In_1388,In_1353);
xnor U50 (N_50,In_2189,In_3);
and U51 (N_51,In_2134,In_1640);
or U52 (N_52,In_893,In_2117);
or U53 (N_53,In_1735,In_1905);
and U54 (N_54,In_1315,In_2479);
and U55 (N_55,In_75,In_2697);
and U56 (N_56,In_790,In_2102);
nand U57 (N_57,In_2865,In_2616);
nand U58 (N_58,In_2140,In_2617);
nor U59 (N_59,In_1050,In_2835);
nor U60 (N_60,In_1951,In_249);
or U61 (N_61,In_876,In_1039);
and U62 (N_62,In_2655,In_2313);
nor U63 (N_63,In_125,In_521);
and U64 (N_64,In_213,In_570);
xor U65 (N_65,In_2589,In_289);
or U66 (N_66,In_874,In_1373);
xnor U67 (N_67,In_2463,In_2280);
nand U68 (N_68,In_2847,In_190);
nand U69 (N_69,In_2586,In_2787);
or U70 (N_70,In_317,In_336);
and U71 (N_71,In_661,In_706);
nand U72 (N_72,In_1425,In_1365);
nand U73 (N_73,In_2105,In_1245);
or U74 (N_74,In_1176,In_1344);
and U75 (N_75,In_142,In_2817);
nor U76 (N_76,In_2752,In_2789);
nor U77 (N_77,In_1555,In_747);
and U78 (N_78,In_2135,In_1940);
or U79 (N_79,In_2264,In_2206);
and U80 (N_80,In_206,In_1813);
xor U81 (N_81,In_1226,In_1471);
xor U82 (N_82,In_89,In_2505);
xor U83 (N_83,In_1582,In_2773);
nor U84 (N_84,In_226,In_1335);
xor U85 (N_85,In_631,In_1265);
nand U86 (N_86,In_2424,In_2942);
nor U87 (N_87,In_1264,In_610);
nand U88 (N_88,In_2420,In_1031);
nor U89 (N_89,In_1509,In_554);
xor U90 (N_90,In_345,In_2454);
nand U91 (N_91,In_920,In_1111);
and U92 (N_92,In_2349,In_1467);
nand U93 (N_93,In_1316,In_1703);
nor U94 (N_94,In_1678,In_2862);
nor U95 (N_95,In_2811,In_1680);
or U96 (N_96,In_2709,In_1498);
nor U97 (N_97,In_1701,In_322);
or U98 (N_98,In_2019,In_2266);
or U99 (N_99,In_2897,In_2470);
or U100 (N_100,In_2520,In_1963);
nor U101 (N_101,In_380,In_781);
and U102 (N_102,In_722,In_1710);
and U103 (N_103,In_2648,In_2031);
and U104 (N_104,In_783,In_1646);
or U105 (N_105,In_2385,In_1355);
and U106 (N_106,In_995,In_1871);
or U107 (N_107,In_2016,In_755);
nor U108 (N_108,In_1170,In_2177);
or U109 (N_109,In_1510,In_312);
nand U110 (N_110,In_2001,In_373);
and U111 (N_111,In_1658,In_50);
and U112 (N_112,In_2929,In_143);
nand U113 (N_113,In_692,In_2603);
nand U114 (N_114,In_1290,In_364);
nor U115 (N_115,In_1590,In_1751);
and U116 (N_116,In_1802,In_1763);
or U117 (N_117,In_843,In_814);
nand U118 (N_118,In_2724,In_1733);
or U119 (N_119,In_915,In_2602);
or U120 (N_120,In_545,In_1852);
and U121 (N_121,In_2795,In_150);
and U122 (N_122,In_2083,In_622);
xor U123 (N_123,In_977,In_2687);
nor U124 (N_124,In_2978,In_2614);
xor U125 (N_125,In_798,In_2372);
nand U126 (N_126,In_2890,In_2407);
or U127 (N_127,In_1462,In_64);
or U128 (N_128,In_2791,In_523);
or U129 (N_129,In_477,In_2492);
nand U130 (N_130,In_2654,In_2023);
nand U131 (N_131,In_1319,In_340);
nand U132 (N_132,In_2464,In_2036);
or U133 (N_133,In_1461,In_333);
and U134 (N_134,In_2491,In_0);
nor U135 (N_135,In_1879,In_152);
nor U136 (N_136,In_679,In_384);
xor U137 (N_137,In_522,In_2236);
or U138 (N_138,In_245,In_1565);
xor U139 (N_139,In_1248,In_1278);
nand U140 (N_140,In_2826,In_2156);
or U141 (N_141,In_1609,In_391);
nand U142 (N_142,In_2904,In_2934);
nor U143 (N_143,In_2566,In_147);
and U144 (N_144,In_1076,In_2625);
nand U145 (N_145,In_546,In_2776);
xnor U146 (N_146,In_2048,In_241);
nand U147 (N_147,In_1433,In_2375);
and U148 (N_148,In_1676,In_1306);
xnor U149 (N_149,In_744,In_1333);
or U150 (N_150,In_1473,In_547);
nor U151 (N_151,In_2252,In_2144);
and U152 (N_152,In_383,In_1151);
nand U153 (N_153,In_375,In_680);
and U154 (N_154,In_445,In_1845);
nand U155 (N_155,In_2549,In_2815);
nor U156 (N_156,In_2432,In_2494);
nor U157 (N_157,In_2692,In_1086);
nor U158 (N_158,In_549,In_2063);
and U159 (N_159,In_868,In_1659);
and U160 (N_160,In_2119,In_359);
and U161 (N_161,In_261,In_1928);
nand U162 (N_162,In_1689,In_1028);
and U163 (N_163,In_34,In_2751);
and U164 (N_164,In_1470,In_2389);
and U165 (N_165,In_371,In_1357);
or U166 (N_166,In_1516,In_1674);
and U167 (N_167,In_858,In_114);
xor U168 (N_168,In_1075,In_1064);
and U169 (N_169,In_2154,In_1550);
xnor U170 (N_170,In_860,In_2311);
and U171 (N_171,In_1882,In_1304);
nor U172 (N_172,In_2886,In_2255);
xnor U173 (N_173,In_2796,In_2115);
nor U174 (N_174,In_1019,In_1015);
xnor U175 (N_175,In_2576,In_507);
nand U176 (N_176,In_2476,In_848);
or U177 (N_177,In_431,In_991);
or U178 (N_178,In_2294,In_616);
xor U179 (N_179,In_1154,In_2440);
or U180 (N_180,In_1125,In_765);
xor U181 (N_181,In_458,In_43);
or U182 (N_182,In_1095,In_1268);
or U183 (N_183,In_1818,In_1588);
nand U184 (N_184,In_2238,In_159);
nand U185 (N_185,In_2686,In_1418);
nand U186 (N_186,In_1374,In_767);
nor U187 (N_187,In_560,In_2717);
or U188 (N_188,In_2081,In_973);
nor U189 (N_189,In_758,In_903);
xor U190 (N_190,In_444,In_1349);
xor U191 (N_191,In_1791,In_869);
nand U192 (N_192,In_376,In_558);
nor U193 (N_193,In_688,In_826);
and U194 (N_194,In_1518,In_2816);
nor U195 (N_195,In_20,In_1548);
and U196 (N_196,In_2225,In_1205);
xor U197 (N_197,In_2714,In_2926);
and U198 (N_198,In_2633,In_2969);
xor U199 (N_199,In_2998,In_704);
nor U200 (N_200,In_2682,In_2911);
xnor U201 (N_201,In_2319,In_2438);
or U202 (N_202,In_1157,In_2670);
nand U203 (N_203,In_1901,In_2679);
xnor U204 (N_204,In_2169,In_2310);
and U205 (N_205,In_129,In_1497);
or U206 (N_206,In_577,In_585);
or U207 (N_207,In_2155,In_1839);
nand U208 (N_208,In_1758,In_926);
xor U209 (N_209,In_2247,In_225);
xor U210 (N_210,In_153,In_1721);
nand U211 (N_211,In_1382,In_1864);
nand U212 (N_212,In_1445,In_2078);
nand U213 (N_213,In_890,In_2199);
or U214 (N_214,In_420,In_1079);
nand U215 (N_215,In_2095,In_1488);
xor U216 (N_216,In_2705,In_481);
or U217 (N_217,In_2075,In_556);
xor U218 (N_218,In_974,In_1141);
nand U219 (N_219,In_177,In_101);
and U220 (N_220,In_2191,In_234);
nor U221 (N_221,In_1089,In_2837);
and U222 (N_222,In_901,In_1260);
nor U223 (N_223,In_248,In_2415);
nor U224 (N_224,In_986,In_1559);
nor U225 (N_225,In_1,In_1456);
nand U226 (N_226,In_1796,In_1665);
and U227 (N_227,In_339,In_2631);
xor U228 (N_228,In_9,In_1232);
nand U229 (N_229,In_600,In_955);
or U230 (N_230,In_1503,In_818);
nor U231 (N_231,In_1444,In_2500);
nand U232 (N_232,In_5,In_985);
xor U233 (N_233,In_1742,In_221);
nor U234 (N_234,In_1432,In_1287);
and U235 (N_235,In_2957,In_151);
nand U236 (N_236,In_1515,In_1848);
and U237 (N_237,In_620,In_1006);
or U238 (N_238,In_697,In_2834);
and U239 (N_239,In_2259,In_1184);
or U240 (N_240,In_708,In_2809);
or U241 (N_241,In_808,In_87);
xor U242 (N_242,In_542,In_1464);
xnor U243 (N_243,In_243,In_2781);
nand U244 (N_244,In_2404,In_634);
xor U245 (N_245,In_228,In_2582);
and U246 (N_246,In_1116,In_2345);
xnor U247 (N_247,In_1391,In_2057);
nand U248 (N_248,In_2366,In_1326);
xor U249 (N_249,In_1952,In_2202);
nand U250 (N_250,In_2059,In_629);
and U251 (N_251,In_2277,In_2232);
nand U252 (N_252,In_1715,In_354);
xnor U253 (N_253,In_760,In_837);
nor U254 (N_254,In_828,In_2484);
xor U255 (N_255,In_402,In_2813);
nor U256 (N_256,In_2040,In_124);
or U257 (N_257,In_2026,In_635);
xnor U258 (N_258,In_1716,In_1599);
xor U259 (N_259,In_726,In_658);
nor U260 (N_260,In_1544,In_2888);
nand U261 (N_261,In_579,In_1586);
nand U262 (N_262,In_275,In_2858);
nand U263 (N_263,In_1135,In_2783);
and U264 (N_264,In_779,In_2009);
and U265 (N_265,In_127,In_173);
nand U266 (N_266,In_2873,In_1091);
xor U267 (N_267,In_290,In_2234);
nand U268 (N_268,In_847,In_2380);
xnor U269 (N_269,In_1942,In_1857);
nand U270 (N_270,In_11,In_67);
nand U271 (N_271,In_1199,In_7);
nor U272 (N_272,In_1907,In_1730);
xor U273 (N_273,In_136,In_1085);
nand U274 (N_274,In_126,In_305);
or U275 (N_275,In_2567,In_1821);
xor U276 (N_276,In_699,In_1902);
or U277 (N_277,In_300,In_348);
xor U278 (N_278,In_2068,In_1521);
or U279 (N_279,In_807,In_2980);
or U280 (N_280,In_2007,In_925);
and U281 (N_281,In_517,In_1016);
xnor U282 (N_282,In_718,In_389);
nand U283 (N_283,In_1422,In_1572);
nor U284 (N_284,In_1043,In_2371);
nor U285 (N_285,In_993,In_46);
nor U286 (N_286,In_854,In_2473);
or U287 (N_287,In_181,In_2565);
nor U288 (N_288,In_2110,In_550);
or U289 (N_289,In_668,In_1954);
nor U290 (N_290,In_2033,In_2486);
nor U291 (N_291,In_1576,In_1823);
or U292 (N_292,In_1745,In_482);
nor U293 (N_293,In_484,In_411);
nand U294 (N_294,In_2577,In_548);
nand U295 (N_295,In_2098,In_2894);
nand U296 (N_296,In_2992,In_592);
and U297 (N_297,In_38,In_2666);
xor U298 (N_298,In_2925,In_1876);
nor U299 (N_299,In_625,In_2373);
xnor U300 (N_300,In_1691,In_2109);
nor U301 (N_301,In_1153,In_2275);
nand U302 (N_302,In_1280,In_672);
or U303 (N_303,In_514,In_2558);
nor U304 (N_304,In_335,In_266);
and U305 (N_305,In_37,In_1222);
nand U306 (N_306,In_2005,In_2584);
xnor U307 (N_307,In_1711,In_1114);
and U308 (N_308,In_2922,In_475);
or U309 (N_309,In_1322,In_2782);
or U310 (N_310,In_1941,In_1884);
or U311 (N_311,In_541,In_2580);
or U312 (N_312,In_2443,In_2300);
nor U313 (N_313,In_797,In_2128);
and U314 (N_314,In_1886,In_1552);
xor U315 (N_315,In_180,In_1334);
nor U316 (N_316,In_1389,In_1443);
nor U317 (N_317,In_2235,In_582);
nand U318 (N_318,In_2270,In_1413);
xor U319 (N_319,In_1181,In_2222);
nand U320 (N_320,In_2561,In_2506);
nor U321 (N_321,In_1460,In_2691);
xnor U322 (N_322,In_1829,In_2229);
xor U323 (N_323,In_1513,In_1168);
or U324 (N_324,In_2619,In_737);
xnor U325 (N_325,In_2877,In_2657);
nand U326 (N_326,In_1889,In_883);
nor U327 (N_327,In_2284,In_1414);
xor U328 (N_328,In_2611,In_1430);
nand U329 (N_329,In_1025,In_374);
xnor U330 (N_330,In_1475,In_134);
nand U331 (N_331,In_1794,In_2778);
nand U332 (N_332,In_738,In_1209);
nand U333 (N_333,In_1810,In_1229);
nand U334 (N_334,In_689,In_1048);
or U335 (N_335,In_442,In_1044);
xor U336 (N_336,In_615,In_1734);
or U337 (N_337,In_1466,In_1771);
or U338 (N_338,In_1854,In_1899);
and U339 (N_339,In_2193,In_2299);
nand U340 (N_340,In_2659,In_1243);
nor U341 (N_341,In_2052,In_1227);
nor U342 (N_342,In_105,In_2866);
and U343 (N_343,In_2356,In_361);
nand U344 (N_344,In_69,In_932);
nor U345 (N_345,In_809,In_2729);
xor U346 (N_346,In_2133,In_1396);
nand U347 (N_347,In_2995,In_2278);
nor U348 (N_348,In_1956,In_2210);
xor U349 (N_349,In_2839,In_341);
nand U350 (N_350,In_77,In_1566);
or U351 (N_351,In_954,In_2743);
or U352 (N_352,In_2151,In_1997);
nor U353 (N_353,In_1429,In_293);
and U354 (N_354,In_80,In_1712);
xnor U355 (N_355,In_2485,In_1449);
nand U356 (N_356,In_632,In_2599);
nor U357 (N_357,In_2955,In_1982);
or U358 (N_358,In_2996,In_441);
nor U359 (N_359,In_1769,In_1600);
and U360 (N_360,In_1077,In_992);
or U361 (N_361,In_2216,In_1138);
nor U362 (N_362,In_1054,In_408);
nor U363 (N_363,In_763,In_1595);
or U364 (N_364,In_1536,In_2528);
nor U365 (N_365,In_1923,In_1180);
nand U366 (N_366,In_1423,In_1874);
nor U367 (N_367,In_1150,In_1237);
nor U368 (N_368,In_1491,In_1128);
and U369 (N_369,In_857,In_313);
xor U370 (N_370,In_392,In_2254);
nor U371 (N_371,In_1267,In_2792);
xor U372 (N_372,In_79,In_1896);
and U373 (N_373,In_2935,In_2120);
or U374 (N_374,In_2806,In_969);
nor U375 (N_375,In_2411,In_2100);
xnor U376 (N_376,In_1005,In_109);
nand U377 (N_377,In_2564,In_395);
nor U378 (N_378,In_1008,In_2032);
nand U379 (N_379,In_396,In_2219);
and U380 (N_380,In_769,In_583);
nor U381 (N_381,In_880,In_1579);
or U382 (N_382,In_315,In_1235);
or U383 (N_383,In_1539,In_1762);
xor U384 (N_384,In_2784,In_1623);
nand U385 (N_385,In_2658,In_1189);
nand U386 (N_386,In_1645,In_2157);
nor U387 (N_387,In_676,In_2051);
and U388 (N_388,In_1681,In_2829);
and U389 (N_389,In_417,In_878);
xor U390 (N_390,In_1293,In_2342);
nand U391 (N_391,In_85,In_1883);
xor U392 (N_392,In_2667,In_1069);
nor U393 (N_393,In_2725,In_1722);
xor U394 (N_394,In_1055,In_832);
or U395 (N_395,In_1981,In_674);
or U396 (N_396,In_1792,In_730);
xor U397 (N_397,In_1909,In_1131);
or U398 (N_398,In_1009,In_1807);
or U399 (N_399,In_2977,In_285);
nand U400 (N_400,In_1805,In_2598);
xnor U401 (N_401,In_2112,In_1024);
or U402 (N_402,In_1350,In_2161);
and U403 (N_403,In_1773,In_2742);
or U404 (N_404,In_637,In_1347);
and U405 (N_405,In_2439,In_2685);
xor U406 (N_406,In_2863,In_533);
nand U407 (N_407,In_1148,In_618);
or U408 (N_408,In_2993,In_2632);
and U409 (N_409,In_1641,In_2469);
nor U410 (N_410,In_2146,In_95);
and U411 (N_411,In_1754,In_645);
or U412 (N_412,In_2848,In_2634);
and U413 (N_413,In_1931,In_2646);
or U414 (N_414,In_308,In_935);
or U415 (N_415,In_2029,In_2258);
nor U416 (N_416,In_158,In_1338);
or U417 (N_417,In_536,In_2271);
or U418 (N_418,In_716,In_1352);
nand U419 (N_419,In_2983,In_782);
nor U420 (N_420,In_530,In_330);
and U421 (N_421,In_1271,In_2218);
nand U422 (N_422,In_1819,In_2551);
and U423 (N_423,In_117,In_1696);
nor U424 (N_424,In_197,In_1560);
or U425 (N_425,In_2308,In_1398);
nand U426 (N_426,In_2333,In_1632);
and U427 (N_427,In_820,In_47);
nand U428 (N_428,In_2012,In_1144);
or U429 (N_429,In_96,In_555);
and U430 (N_430,In_283,In_1842);
and U431 (N_431,In_695,In_2895);
and U432 (N_432,In_756,In_478);
or U433 (N_433,In_8,In_2325);
and U434 (N_434,In_1832,In_2241);
xnor U435 (N_435,In_1327,In_2088);
nor U436 (N_436,In_1062,In_2712);
nand U437 (N_437,In_465,In_123);
xor U438 (N_438,In_1119,In_1826);
and U439 (N_439,In_2604,In_569);
or U440 (N_440,In_1693,In_989);
xnor U441 (N_441,In_2159,In_1809);
nor U442 (N_442,In_1814,In_2923);
or U443 (N_443,In_1752,In_703);
and U444 (N_444,In_2510,In_2930);
or U445 (N_445,In_1018,In_666);
or U446 (N_446,In_1567,In_719);
nor U447 (N_447,In_578,In_1906);
nand U448 (N_448,In_771,In_951);
nand U449 (N_449,In_1359,In_496);
xnor U450 (N_450,In_1156,In_2312);
nor U451 (N_451,In_18,In_2129);
xnor U452 (N_452,In_1482,In_1354);
or U453 (N_453,In_930,In_1589);
nand U454 (N_454,In_2903,In_916);
nor U455 (N_455,In_591,In_342);
nand U456 (N_456,In_2391,In_1007);
and U457 (N_457,In_2041,In_659);
or U458 (N_458,In_259,In_2101);
nand U459 (N_459,In_1859,In_2212);
xor U460 (N_460,In_2823,In_835);
nor U461 (N_461,In_1415,In_1861);
and U462 (N_462,In_386,In_1073);
nor U463 (N_463,In_156,In_120);
nor U464 (N_464,In_270,In_884);
nand U465 (N_465,In_537,In_853);
and U466 (N_466,In_2422,In_1336);
nor U467 (N_467,In_709,In_1393);
nand U468 (N_468,In_2513,In_2539);
xor U469 (N_469,In_2537,In_2797);
and U470 (N_470,In_2606,In_2749);
and U471 (N_471,In_1295,In_2887);
xnor U472 (N_472,In_2689,In_2351);
xor U473 (N_473,In_2713,In_372);
xnor U474 (N_474,In_1933,In_2365);
xnor U475 (N_475,In_1106,In_1123);
nand U476 (N_476,In_1262,In_2295);
nor U477 (N_477,In_1512,In_98);
xor U478 (N_478,In_2741,In_673);
xor U479 (N_479,In_183,In_2880);
xnor U480 (N_480,In_598,In_310);
and U481 (N_481,In_2845,In_1013);
and U482 (N_482,In_2593,In_1568);
or U483 (N_483,In_1634,In_975);
xor U484 (N_484,In_1833,In_960);
nand U485 (N_485,In_1058,In_1387);
xor U486 (N_486,In_1455,In_238);
xnor U487 (N_487,In_1581,In_1765);
xnor U488 (N_488,In_1434,In_406);
nand U489 (N_489,In_2961,In_1083);
nor U490 (N_490,In_2248,In_1244);
nor U491 (N_491,In_1010,In_2084);
and U492 (N_492,In_2419,In_1481);
nand U493 (N_493,In_2597,In_979);
xor U494 (N_494,In_2379,In_233);
nand U495 (N_495,In_525,In_1738);
nor U496 (N_496,In_2754,In_1596);
nor U497 (N_497,In_2164,In_1628);
or U498 (N_498,In_2803,In_1719);
and U499 (N_499,In_1962,In_1863);
xor U500 (N_500,In_2770,In_316);
and U501 (N_501,In_2615,In_2757);
and U502 (N_502,In_1937,In_922);
or U503 (N_503,In_440,In_2960);
and U504 (N_504,In_2437,In_2677);
nor U505 (N_505,In_2292,In_2529);
nor U506 (N_506,In_1837,In_2286);
nand U507 (N_507,In_907,In_470);
nor U508 (N_508,In_2856,In_966);
nand U509 (N_509,In_112,In_1210);
xnor U510 (N_510,In_185,In_349);
nand U511 (N_511,In_63,In_2445);
and U512 (N_512,In_1672,In_2511);
or U513 (N_513,In_1152,In_1783);
nor U514 (N_514,In_1939,In_2341);
nand U515 (N_515,In_732,In_303);
nand U516 (N_516,In_949,In_236);
nor U517 (N_517,In_2570,In_1190);
nor U518 (N_518,In_55,In_1965);
and U519 (N_519,In_2545,In_1760);
nand U520 (N_520,In_387,In_1146);
nand U521 (N_521,In_2322,In_2400);
nand U522 (N_522,In_2799,In_2710);
xor U523 (N_523,In_1324,In_1617);
or U524 (N_524,In_2131,In_999);
xnor U525 (N_525,In_686,In_2896);
xor U526 (N_526,In_1652,In_861);
nand U527 (N_527,In_1790,In_191);
nor U528 (N_528,In_1263,In_267);
or U529 (N_529,In_1988,In_603);
nand U530 (N_530,In_2337,In_870);
and U531 (N_531,In_2509,In_1092);
and U532 (N_532,In_84,In_1911);
or U533 (N_533,In_2060,In_1729);
xor U534 (N_534,In_1577,In_1774);
nor U535 (N_535,In_2653,In_334);
xnor U536 (N_536,In_1277,In_1384);
and U537 (N_537,In_2257,In_362);
and U538 (N_538,In_1014,In_2986);
or U539 (N_539,In_415,In_1921);
xor U540 (N_540,In_1585,In_2828);
nand U541 (N_541,In_1112,In_1811);
and U542 (N_542,In_590,In_1915);
xor U543 (N_543,In_1526,In_2718);
or U544 (N_544,In_2167,In_1584);
and U545 (N_545,In_896,In_1356);
nor U546 (N_546,In_1472,In_717);
nand U547 (N_547,In_2386,In_1294);
xnor U548 (N_548,In_795,In_1858);
xnor U549 (N_549,In_1872,In_1409);
nor U550 (N_550,In_2071,In_2711);
and U551 (N_551,In_1545,In_1328);
nand U552 (N_552,In_2174,In_1242);
or U553 (N_553,In_1637,In_1286);
nor U554 (N_554,In_1817,In_1435);
nand U555 (N_555,In_2786,In_492);
xnor U556 (N_556,In_865,In_83);
xor U557 (N_557,In_2912,In_1970);
and U558 (N_558,In_2050,In_353);
nand U559 (N_559,In_1053,In_959);
or U560 (N_560,In_1675,In_2726);
nor U561 (N_561,In_2466,In_1991);
or U562 (N_562,In_1563,In_1908);
or U563 (N_563,In_2552,In_2243);
nor U564 (N_564,In_451,In_2074);
and U565 (N_565,In_1593,In_2303);
and U566 (N_566,In_2282,In_483);
nor U567 (N_567,In_1841,In_1012);
and U568 (N_568,In_1583,In_899);
or U569 (N_569,In_56,In_1097);
xor U570 (N_570,In_1179,In_851);
nand U571 (N_571,In_427,In_806);
nor U572 (N_572,In_239,In_1218);
and U573 (N_573,In_2425,In_2186);
nor U574 (N_574,In_2298,In_360);
and U575 (N_575,In_54,In_326);
or U576 (N_576,In_2198,In_2630);
xor U577 (N_577,In_2950,In_1362);
and U578 (N_578,In_2163,In_2039);
xnor U579 (N_579,In_1161,In_1531);
and U580 (N_580,In_2690,In_2546);
xor U581 (N_581,In_2124,In_446);
or U582 (N_582,In_1977,In_2532);
and U583 (N_583,In_2173,In_1713);
xor U584 (N_584,In_710,In_2364);
nor U585 (N_585,In_2762,In_1298);
xor U586 (N_586,In_1194,In_2952);
and U587 (N_587,In_2972,In_2975);
nor U588 (N_588,In_2798,In_2272);
nand U589 (N_589,In_2671,In_971);
or U590 (N_590,In_2442,In_138);
and U591 (N_591,In_1770,In_1147);
nor U592 (N_592,In_2637,In_1558);
and U593 (N_593,In_904,In_1063);
and U594 (N_594,In_2381,In_1281);
xor U595 (N_595,In_1348,In_439);
xor U596 (N_596,In_199,In_1912);
nand U597 (N_597,In_1891,In_2387);
nand U598 (N_598,In_2855,In_943);
and U599 (N_599,In_611,In_751);
or U600 (N_600,In_113,In_2111);
nor U601 (N_601,In_377,In_2673);
xor U602 (N_602,In_532,In_2650);
xor U603 (N_603,In_394,In_2182);
nand U604 (N_604,In_2967,In_379);
nor U605 (N_605,In_1642,In_830);
nor U606 (N_606,In_871,In_931);
nor U607 (N_607,In_1633,In_1297);
and U608 (N_608,In_1996,In_1132);
or U609 (N_609,In_984,In_1381);
or U610 (N_610,In_654,In_1337);
and U611 (N_611,In_1447,In_187);
nor U612 (N_612,In_1164,In_2769);
nand U613 (N_613,In_2426,In_251);
nand U614 (N_614,In_1725,In_1797);
xnor U615 (N_615,In_1999,In_260);
xnor U616 (N_616,In_459,In_1120);
nand U617 (N_617,In_2675,In_862);
xor U618 (N_618,In_486,In_833);
and U619 (N_619,In_2719,In_222);
nand U620 (N_620,In_1220,In_2478);
and U621 (N_621,In_1061,In_2859);
xnor U622 (N_622,In_165,In_2203);
nand U623 (N_623,In_1332,In_1175);
or U624 (N_624,In_29,In_1279);
or U625 (N_625,In_946,In_1824);
nand U626 (N_626,In_2536,In_456);
xor U627 (N_627,In_253,In_627);
nand U628 (N_628,In_1679,In_2519);
nor U629 (N_629,In_543,In_2142);
or U630 (N_630,In_1463,In_1033);
nor U631 (N_631,In_2507,In_2260);
xor U632 (N_632,In_1660,In_2958);
and U633 (N_633,In_1619,In_21);
or U634 (N_634,In_2590,In_1668);
nand U635 (N_635,In_1825,In_2660);
and U636 (N_636,In_2046,In_278);
nand U637 (N_637,In_224,In_2104);
nor U638 (N_638,In_184,In_286);
and U639 (N_639,In_1975,In_352);
and U640 (N_640,In_2253,In_1291);
xor U641 (N_641,In_2497,In_437);
or U642 (N_642,In_1484,In_2827);
xnor U643 (N_643,In_2338,In_1714);
nor U644 (N_644,In_81,In_332);
nand U645 (N_645,In_331,In_276);
and U646 (N_646,In_2641,In_1786);
and U647 (N_647,In_1777,In_1607);
or U648 (N_648,In_1431,In_207);
nand U649 (N_649,In_1302,In_2327);
nand U650 (N_650,In_2394,In_155);
and U651 (N_651,In_594,In_728);
xnor U652 (N_652,In_2841,In_1844);
or U653 (N_653,In_2273,In_742);
or U654 (N_654,In_2518,In_786);
nand U655 (N_655,In_1610,In_801);
nor U656 (N_656,In_2618,In_2780);
and U657 (N_657,In_1525,In_501);
nand U658 (N_658,In_898,In_2462);
nor U659 (N_659,In_209,In_92);
or U660 (N_660,In_944,In_160);
nand U661 (N_661,In_2578,In_1866);
nand U662 (N_662,In_526,In_587);
and U663 (N_663,In_540,In_1873);
or U664 (N_664,In_2833,In_1587);
xnor U665 (N_665,In_397,In_490);
nand U666 (N_666,In_6,In_480);
or U667 (N_667,In_983,In_2239);
xor U668 (N_668,In_174,In_2217);
and U669 (N_669,In_2452,In_2968);
nor U670 (N_670,In_509,In_2810);
or U671 (N_671,In_1036,In_2832);
xor U672 (N_672,In_2096,In_1323);
nand U673 (N_673,In_229,In_754);
nand U674 (N_674,In_2044,In_2916);
nand U675 (N_675,In_2985,In_2883);
xnor U676 (N_676,In_2368,In_1974);
and U677 (N_677,In_469,In_1897);
nand U678 (N_678,In_2644,In_2976);
nand U679 (N_679,In_1605,In_621);
and U680 (N_680,In_2402,In_552);
nor U681 (N_681,In_2588,In_172);
nand U682 (N_682,In_2204,In_1822);
nor U683 (N_683,In_17,In_140);
nand U684 (N_684,In_1478,In_2885);
or U685 (N_685,In_2099,In_2879);
nor U686 (N_686,In_952,In_1638);
or U687 (N_687,In_2964,In_72);
or U688 (N_688,In_60,In_2825);
and U689 (N_689,In_913,In_2680);
nor U690 (N_690,In_381,In_1236);
or U691 (N_691,In_595,In_1124);
nand U692 (N_692,In_434,In_2612);
or U693 (N_693,In_2676,In_2489);
nor U694 (N_694,In_329,In_2963);
and U695 (N_695,In_2465,In_1417);
or U696 (N_696,In_284,In_2158);
nand U697 (N_697,In_1173,In_888);
xnor U698 (N_698,In_2213,In_1292);
nor U699 (N_699,In_2475,In_1784);
and U700 (N_700,In_867,In_2263);
nor U701 (N_701,In_2384,In_16);
nand U702 (N_702,In_626,In_1917);
nand U703 (N_703,In_304,In_720);
xnor U704 (N_704,In_1920,In_777);
and U705 (N_705,In_1214,In_2073);
and U706 (N_706,In_2022,In_1072);
or U707 (N_707,In_1958,In_436);
or U708 (N_708,In_2768,In_1875);
nor U709 (N_709,In_68,In_1410);
nor U710 (N_710,In_1100,In_2647);
or U711 (N_711,In_1137,In_713);
nand U712 (N_712,In_368,In_2287);
nand U713 (N_713,In_2195,In_1492);
nor U714 (N_714,In_1274,In_1925);
nor U715 (N_715,In_2920,In_1272);
xnor U716 (N_716,In_1042,In_2251);
xor U717 (N_717,In_2047,In_1215);
xnor U718 (N_718,In_908,In_121);
and U719 (N_719,In_1557,In_1201);
or U720 (N_720,In_460,In_244);
and U721 (N_721,In_2200,In_1188);
or U722 (N_722,In_15,In_1913);
nand U723 (N_723,In_524,In_2196);
or U724 (N_724,In_1307,In_1538);
xnor U725 (N_725,In_1766,In_299);
nor U726 (N_726,In_1300,In_2496);
nor U727 (N_727,In_2148,In_343);
or U728 (N_728,In_1479,In_2559);
xnor U729 (N_729,In_821,In_1330);
nor U730 (N_730,In_1360,In_2053);
nor U731 (N_731,In_1318,In_838);
nor U732 (N_732,In_967,In_1635);
nand U733 (N_733,In_2409,In_912);
xor U734 (N_734,In_671,In_2984);
xor U735 (N_735,In_281,In_1439);
or U736 (N_736,In_2664,In_2030);
and U737 (N_737,In_257,In_2696);
or U738 (N_738,In_2455,In_370);
or U739 (N_739,In_2688,In_796);
and U740 (N_740,In_2843,In_565);
and U741 (N_741,In_1204,In_2870);
nand U742 (N_742,In_2607,In_2413);
xor U743 (N_743,In_2149,In_424);
xnor U744 (N_744,In_650,In_2533);
and U745 (N_745,In_761,In_1643);
nor U746 (N_746,In_982,In_1495);
nand U747 (N_747,In_1068,In_770);
nor U748 (N_748,In_823,In_800);
and U749 (N_749,In_2736,In_2525);
nor U750 (N_750,In_2802,In_502);
xor U751 (N_751,In_2579,In_2747);
xor U752 (N_752,In_2830,In_2861);
or U753 (N_753,In_170,In_794);
xnor U754 (N_754,In_279,In_2092);
nand U755 (N_755,In_419,In_314);
xnor U756 (N_756,In_2921,In_500);
nand U757 (N_757,In_2764,In_2428);
nor U758 (N_758,In_551,In_49);
xor U759 (N_759,In_220,In_2321);
nor U760 (N_760,In_562,In_2850);
or U761 (N_761,In_2318,In_735);
nor U762 (N_762,In_2853,In_108);
nor U763 (N_763,In_1726,In_2317);
or U764 (N_764,In_232,In_1592);
or U765 (N_765,In_2392,In_948);
xor U766 (N_766,In_2669,In_1629);
nand U767 (N_767,In_2575,In_2521);
xnor U768 (N_768,In_2187,In_2274);
xnor U769 (N_769,In_2358,In_1476);
xnor U770 (N_770,In_132,In_1504);
nand U771 (N_771,In_508,In_574);
nand U772 (N_772,In_288,In_799);
nor U773 (N_773,In_839,In_2973);
xnor U774 (N_774,In_2237,In_1661);
nor U775 (N_775,In_2395,In_2722);
xnor U776 (N_776,In_1747,In_1570);
nand U777 (N_777,In_1207,In_1904);
and U778 (N_778,In_1505,In_2909);
and U779 (N_779,In_2211,In_1578);
or U780 (N_780,In_1707,In_1741);
or U781 (N_781,In_2336,In_295);
nand U782 (N_782,In_1612,In_271);
nor U783 (N_783,In_1247,In_2765);
or U784 (N_784,In_1968,In_664);
nor U785 (N_785,In_1507,In_1165);
nor U786 (N_786,In_1708,In_2571);
xor U787 (N_787,In_1601,In_499);
nand U788 (N_788,In_586,In_2899);
nand U789 (N_789,In_2544,In_252);
nand U790 (N_790,In_2399,In_2171);
or U791 (N_791,In_1167,In_687);
nand U792 (N_792,In_2107,In_2061);
nor U793 (N_793,In_793,In_235);
and U794 (N_794,In_2153,In_1556);
and U795 (N_795,In_1755,In_1995);
and U796 (N_796,In_201,In_115);
and U797 (N_797,In_819,In_1890);
nor U798 (N_798,In_217,In_1685);
and U799 (N_799,In_1549,In_2249);
nor U800 (N_800,In_1017,In_1407);
xnor U801 (N_801,In_1059,In_1892);
nand U802 (N_802,In_1452,In_88);
and U803 (N_803,In_1074,In_2042);
nand U804 (N_804,In_263,In_1801);
xor U805 (N_805,In_2328,In_846);
or U806 (N_806,In_628,In_1799);
nor U807 (N_807,In_2917,In_1296);
xor U808 (N_808,In_2594,In_825);
and U809 (N_809,In_1528,In_1945);
xor U810 (N_810,In_775,In_725);
and U811 (N_811,In_1694,In_1759);
or U812 (N_812,In_2062,In_2763);
or U813 (N_813,In_2623,In_538);
nand U814 (N_814,In_997,In_2836);
nand U815 (N_815,In_1614,In_1030);
nor U816 (N_816,In_1787,In_2555);
nand U817 (N_817,In_1219,In_2091);
and U818 (N_818,In_2388,In_2662);
and U819 (N_819,In_2893,In_93);
or U820 (N_820,In_1385,In_321);
and U821 (N_821,In_656,In_784);
and U822 (N_822,In_2244,In_2801);
nor U823 (N_823,In_2548,In_1878);
and U824 (N_824,In_443,In_1772);
nand U825 (N_825,In_2693,In_2150);
xnor U826 (N_826,In_2499,In_2755);
nor U827 (N_827,In_1978,In_1397);
nor U828 (N_828,In_1090,In_1172);
xor U829 (N_829,In_2530,In_1731);
xnor U830 (N_830,In_535,In_1880);
xnor U831 (N_831,In_972,In_1034);
and U832 (N_832,In_292,In_58);
and U833 (N_833,In_473,In_906);
or U834 (N_834,In_1411,In_2731);
xnor U835 (N_835,In_2208,In_1406);
or U836 (N_836,In_736,In_457);
nand U837 (N_837,In_534,In_2305);
nor U838 (N_838,In_418,In_472);
nor U839 (N_839,In_2335,In_2891);
nand U840 (N_840,In_575,In_1392);
nand U841 (N_841,In_2138,In_2483);
and U842 (N_842,In_1211,In_2256);
and U843 (N_843,In_642,In_905);
nand U844 (N_844,In_2227,In_2495);
or U845 (N_845,In_1107,In_2613);
or U846 (N_846,In_778,In_189);
nor U847 (N_847,In_2936,In_2943);
xor U848 (N_848,In_1155,In_1339);
nor U849 (N_849,In_1573,In_2735);
xor U850 (N_850,In_1309,In_216);
nor U851 (N_851,In_2201,In_2435);
and U852 (N_852,In_25,In_423);
or U853 (N_853,In_144,In_294);
or U854 (N_854,In_1225,In_1692);
nor U855 (N_855,In_2639,In_1060);
nand U856 (N_856,In_2114,In_269);
nor U857 (N_857,In_1066,In_2055);
nor U858 (N_858,In_2852,In_254);
xor U859 (N_859,In_2951,In_963);
xnor U860 (N_860,In_2000,In_836);
or U861 (N_861,In_1519,In_2010);
nand U862 (N_862,In_2352,In_407);
nor U863 (N_863,In_2774,In_1644);
and U864 (N_864,In_849,In_2753);
and U865 (N_865,In_28,In_2034);
and U866 (N_866,In_573,In_1368);
xnor U867 (N_867,In_1142,In_1372);
nor U868 (N_868,In_82,In_1193);
xor U869 (N_869,In_1914,In_1580);
or U870 (N_870,In_1598,In_1020);
xor U871 (N_871,In_2516,In_1284);
and U872 (N_872,In_1718,In_1989);
xnor U873 (N_873,In_1764,In_45);
xnor U874 (N_874,In_12,In_2340);
and U875 (N_875,In_2304,In_1604);
or U876 (N_876,In_2585,In_2307);
xor U877 (N_877,In_1924,In_2876);
nand U878 (N_878,In_2185,In_2192);
and U879 (N_879,In_2906,In_2744);
and U880 (N_880,In_1325,In_2106);
nand U881 (N_881,In_2290,In_1122);
nand U882 (N_882,In_2554,In_2472);
and U883 (N_883,In_2332,In_1468);
or U884 (N_884,In_2459,In_2025);
and U885 (N_885,In_1399,In_2181);
nand U886 (N_886,In_1535,In_2416);
nand U887 (N_887,In_2547,In_2289);
nor U888 (N_888,In_553,In_1736);
and U889 (N_889,In_604,In_2293);
xnor U890 (N_890,In_1234,In_162);
nor U891 (N_891,In_2179,In_1541);
xor U892 (N_892,In_1217,In_1440);
nor U893 (N_893,In_1983,In_2355);
nor U894 (N_894,In_559,In_593);
nand U895 (N_895,In_1547,In_1450);
xor U896 (N_896,In_2583,In_219);
or U897 (N_897,In_2344,In_1047);
nor U898 (N_898,In_1021,In_2541);
xnor U899 (N_899,In_2941,In_624);
nand U900 (N_900,In_1943,In_148);
or U901 (N_901,In_1948,In_927);
xnor U902 (N_902,In_1994,In_2436);
nor U903 (N_903,In_1990,In_2035);
nand U904 (N_904,In_2427,In_2461);
and U905 (N_905,In_369,In_1394);
nand U906 (N_906,In_1251,In_435);
or U907 (N_907,In_1998,In_788);
nor U908 (N_908,In_2066,In_1465);
nand U909 (N_909,In_657,In_2223);
and U910 (N_910,In_2089,In_2775);
nand U911 (N_911,In_167,In_205);
or U912 (N_912,In_563,In_2875);
and U913 (N_913,In_544,In_416);
xnor U914 (N_914,In_1611,In_2230);
or U915 (N_915,In_2020,In_2515);
xor U916 (N_916,In_319,In_2246);
nor U917 (N_917,In_2716,In_2557);
and U918 (N_918,In_2397,In_504);
xor U919 (N_919,In_1254,In_42);
xor U920 (N_920,In_2343,In_1815);
xor U921 (N_921,In_1266,In_1739);
nand U922 (N_922,In_1149,In_1458);
nor U923 (N_923,In_964,In_2132);
nor U924 (N_924,In_2457,In_2456);
xor U925 (N_925,In_2183,In_1918);
or U926 (N_926,In_2919,In_571);
xnor U927 (N_927,In_2730,In_1174);
or U928 (N_928,In_2401,In_996);
nor U929 (N_929,In_1793,In_1239);
xnor U930 (N_930,In_2820,In_2527);
nor U931 (N_931,In_2531,In_2868);
or U932 (N_932,In_2938,In_539);
nand U933 (N_933,In_53,In_723);
nand U934 (N_934,In_57,In_264);
nor U935 (N_935,In_448,In_889);
nor U936 (N_936,In_2864,In_1159);
nand U937 (N_937,In_1185,In_211);
or U938 (N_938,In_2989,In_2596);
or U939 (N_939,In_1276,In_2160);
and U940 (N_940,In_280,In_2807);
xnor U941 (N_941,In_588,In_745);
xor U942 (N_942,In_2651,In_161);
or U943 (N_943,In_875,In_2446);
nor U944 (N_944,In_1195,In_663);
or U945 (N_945,In_1597,In_2370);
or U946 (N_946,In_1233,In_506);
nor U947 (N_947,In_1843,In_1944);
or U948 (N_948,In_2965,In_1749);
nand U949 (N_949,In_2932,In_337);
nor U950 (N_950,In_1117,In_759);
nand U951 (N_951,In_227,In_608);
nand U952 (N_952,In_2842,In_350);
xnor U953 (N_953,In_1919,In_99);
nand U954 (N_954,In_325,In_363);
and U955 (N_955,In_2077,In_2622);
nor U956 (N_956,In_1249,In_2573);
xnor U957 (N_957,In_2502,In_1682);
xnor U958 (N_958,In_2918,In_655);
nand U959 (N_959,In_2846,In_2482);
nor U960 (N_960,In_2882,In_1756);
nor U961 (N_961,In_919,In_1575);
or U962 (N_962,In_576,In_1084);
nor U963 (N_963,In_218,In_685);
nor U964 (N_964,In_2788,In_1957);
xnor U965 (N_965,In_2620,In_202);
xnor U966 (N_966,In_2309,In_644);
nand U967 (N_967,In_2665,In_1534);
xnor U968 (N_968,In_1768,In_2233);
or U969 (N_969,In_1363,In_2014);
nor U970 (N_970,In_2405,In_256);
xor U971 (N_971,In_2649,In_1514);
xnor U972 (N_972,In_282,In_566);
nor U973 (N_973,In_636,In_1571);
xor U974 (N_974,In_2638,In_2878);
nor U975 (N_975,In_1699,In_1057);
and U976 (N_976,In_463,In_772);
nor U977 (N_977,In_1867,In_512);
and U978 (N_978,In_2592,In_1140);
nand U979 (N_979,In_1489,In_2471);
and U980 (N_980,In_844,In_1004);
nand U981 (N_981,In_2357,In_1101);
and U982 (N_982,In_2450,In_1177);
nor U983 (N_983,In_2522,In_297);
nor U984 (N_984,In_2487,In_994);
nand U985 (N_985,In_2699,In_2987);
and U986 (N_986,In_306,In_2141);
and U987 (N_987,In_1684,In_2999);
nor U988 (N_988,In_90,In_2015);
nor U989 (N_989,In_2600,In_1093);
and U990 (N_990,In_78,In_1653);
xor U991 (N_991,In_1893,In_910);
nand U992 (N_992,In_2130,In_1000);
xor U993 (N_993,In_188,In_746);
or U994 (N_994,In_1029,In_911);
and U995 (N_995,In_2139,In_2197);
and U996 (N_996,In_1537,In_2113);
or U997 (N_997,In_214,In_1098);
xnor U998 (N_998,In_945,In_1022);
xnor U999 (N_999,In_640,In_65);
or U1000 (N_1000,In_203,In_30);
or U1001 (N_1001,In_4,In_2214);
nand U1002 (N_1002,In_727,In_928);
xnor U1003 (N_1003,In_2268,In_2860);
or U1004 (N_1004,In_1345,In_2205);
and U1005 (N_1005,In_886,In_2838);
xor U1006 (N_1006,In_2123,In_953);
nand U1007 (N_1007,In_612,In_866);
nor U1008 (N_1008,In_471,In_164);
and U1009 (N_1009,In_2207,In_1553);
and U1010 (N_1010,In_157,In_614);
xor U1011 (N_1011,In_2377,In_237);
nand U1012 (N_1012,In_250,In_23);
nor U1013 (N_1013,In_887,In_1448);
and U1014 (N_1014,In_1836,In_711);
nand U1015 (N_1015,In_31,In_2024);
nand U1016 (N_1016,In_1127,In_1828);
nor U1017 (N_1017,In_2190,In_1540);
and U1018 (N_1018,In_1023,In_1441);
or U1019 (N_1019,In_2279,In_2324);
or U1020 (N_1020,In_1780,In_2431);
nand U1021 (N_1021,In_1926,In_2694);
nor U1022 (N_1022,In_1200,In_2901);
or U1023 (N_1023,In_731,In_494);
nor U1024 (N_1024,In_811,In_1746);
nand U1025 (N_1025,In_2626,In_1082);
nor U1026 (N_1026,In_1087,In_1554);
nor U1027 (N_1027,In_320,In_2176);
and U1028 (N_1028,In_1380,In_2746);
nor U1029 (N_1029,In_2732,In_1282);
xor U1030 (N_1030,In_1546,In_1183);
and U1031 (N_1031,In_1477,In_1070);
xnor U1032 (N_1032,In_503,In_230);
xnor U1033 (N_1033,In_1621,In_1130);
nand U1034 (N_1034,In_1900,In_1104);
nor U1035 (N_1035,In_1955,In_1198);
nand U1036 (N_1036,In_2011,In_2708);
nand U1037 (N_1037,In_204,In_581);
or U1038 (N_1038,In_2076,In_107);
or U1039 (N_1039,In_1240,In_1402);
nor U1040 (N_1040,In_2701,In_14);
nor U1041 (N_1041,In_1310,In_2824);
or U1042 (N_1042,In_2330,In_662);
and U1043 (N_1043,In_724,In_242);
or U1044 (N_1044,In_774,In_327);
nand U1045 (N_1045,In_1795,In_2226);
or U1046 (N_1046,In_195,In_2143);
nor U1047 (N_1047,In_748,In_2448);
xnor U1048 (N_1048,In_429,In_2572);
nand U1049 (N_1049,In_401,In_2944);
or U1050 (N_1050,In_1231,In_2794);
xnor U1051 (N_1051,In_1032,In_792);
or U1052 (N_1052,In_1493,In_2946);
xnor U1053 (N_1053,In_863,In_382);
xnor U1054 (N_1054,In_768,In_2209);
nor U1055 (N_1055,In_1761,In_1483);
or U1056 (N_1056,In_467,In_2902);
nand U1057 (N_1057,In_62,In_1569);
xnor U1058 (N_1058,In_957,In_1202);
or U1059 (N_1059,In_879,In_1358);
nor U1060 (N_1060,In_1511,In_2281);
or U1061 (N_1061,In_2003,In_1379);
nand U1062 (N_1062,In_2334,In_962);
and U1063 (N_1063,In_1250,In_1647);
nor U1064 (N_1064,In_497,In_1312);
nor U1065 (N_1065,In_2808,In_1667);
xnor U1066 (N_1066,In_652,In_2881);
and U1067 (N_1067,In_1850,In_1261);
nor U1068 (N_1068,In_1308,In_681);
nand U1069 (N_1069,In_430,In_856);
xnor U1070 (N_1070,In_2966,In_102);
or U1071 (N_1071,In_1529,In_1562);
nor U1072 (N_1072,In_733,In_753);
xnor U1073 (N_1073,In_2715,In_1608);
or U1074 (N_1074,In_1451,In_2683);
nand U1075 (N_1075,In_2043,In_1273);
and U1076 (N_1076,In_2359,In_1289);
nand U1077 (N_1077,In_1789,In_2982);
and U1078 (N_1078,In_2441,In_128);
xor U1079 (N_1079,In_2329,In_76);
xor U1080 (N_1080,In_2406,In_605);
nor U1081 (N_1081,In_1228,In_2937);
and U1082 (N_1082,In_163,In_1624);
xor U1083 (N_1083,In_106,In_139);
nor U1084 (N_1084,In_1631,In_2080);
xnor U1085 (N_1085,In_2122,In_1648);
and U1086 (N_1086,In_1499,In_2021);
nand U1087 (N_1087,In_2777,In_1946);
or U1088 (N_1088,In_178,In_1027);
nand U1089 (N_1089,In_2514,In_568);
nor U1090 (N_1090,In_2166,In_2997);
or U1091 (N_1091,In_2417,In_2991);
nand U1092 (N_1092,In_669,In_131);
or U1093 (N_1093,In_1171,In_1740);
nand U1094 (N_1094,In_721,In_694);
nand U1095 (N_1095,In_302,In_2678);
xnor U1096 (N_1096,In_2376,In_1935);
or U1097 (N_1097,In_1331,In_1532);
nor U1098 (N_1098,In_529,In_613);
or U1099 (N_1099,In_965,In_1480);
xnor U1100 (N_1100,In_273,In_881);
or U1101 (N_1101,In_2058,In_1317);
nor U1102 (N_1102,In_2265,In_1037);
nand U1103 (N_1103,In_606,In_2948);
xnor U1104 (N_1104,In_2430,In_488);
nand U1105 (N_1105,In_1705,In_1808);
nor U1106 (N_1106,In_2970,In_859);
and U1107 (N_1107,In_773,In_2285);
nand U1108 (N_1108,In_2320,In_648);
and U1109 (N_1109,In_208,In_1947);
xor U1110 (N_1110,In_2543,In_1437);
nand U1111 (N_1111,In_1080,In_2605);
nor U1112 (N_1112,In_200,In_2913);
or U1113 (N_1113,In_824,In_1376);
and U1114 (N_1114,In_464,In_2550);
and U1115 (N_1115,In_2421,In_1446);
xnor U1116 (N_1116,In_2412,In_2362);
or U1117 (N_1117,In_1800,In_841);
and U1118 (N_1118,In_1744,In_1865);
and U1119 (N_1119,In_1840,In_1834);
or U1120 (N_1120,In_2740,In_2049);
and U1121 (N_1121,In_1494,In_2553);
or U1122 (N_1122,In_827,In_2093);
and U1123 (N_1123,In_2704,In_1737);
or U1124 (N_1124,In_894,In_1846);
and U1125 (N_1125,In_1856,In_2542);
or U1126 (N_1126,In_998,In_510);
and U1127 (N_1127,In_939,In_1959);
and U1128 (N_1128,In_1574,In_1669);
xnor U1129 (N_1129,In_1847,In_2339);
xor U1130 (N_1130,In_791,In_1438);
or U1131 (N_1131,In_1985,In_619);
and U1132 (N_1132,In_1496,In_347);
and U1133 (N_1133,In_1626,In_1252);
nor U1134 (N_1134,In_2812,In_1602);
or U1135 (N_1135,In_2028,In_1798);
and U1136 (N_1136,In_145,In_1377);
xor U1137 (N_1137,In_1894,In_2423);
xor U1138 (N_1138,In_1088,In_714);
and U1139 (N_1139,In_2645,In_450);
nand U1140 (N_1140,In_2045,In_617);
nand U1141 (N_1141,In_2396,In_48);
nand U1142 (N_1142,In_776,In_2353);
nand U1143 (N_1143,In_2194,In_13);
nand U1144 (N_1144,In_1953,In_176);
nand U1145 (N_1145,In_1781,In_691);
or U1146 (N_1146,In_2361,In_1099);
nand U1147 (N_1147,In_1664,In_1695);
xor U1148 (N_1148,In_2474,In_2939);
nor U1149 (N_1149,In_1487,In_766);
and U1150 (N_1150,In_1927,In_1704);
nor U1151 (N_1151,In_1343,In_1855);
and U1152 (N_1152,In_1346,In_498);
xnor U1153 (N_1153,In_1727,In_2302);
and U1154 (N_1154,In_1748,In_764);
xnor U1155 (N_1155,In_2601,In_638);
or U1156 (N_1156,In_398,In_2276);
nor U1157 (N_1157,In_2116,In_1986);
or U1158 (N_1158,In_27,In_840);
nand U1159 (N_1159,In_2652,In_2079);
or U1160 (N_1160,In_1830,In_1408);
or U1161 (N_1161,In_2591,In_1831);
nor U1162 (N_1162,In_2627,In_852);
nor U1163 (N_1163,In_527,In_2988);
or U1164 (N_1164,In_2956,In_2504);
or U1165 (N_1165,In_154,In_988);
or U1166 (N_1166,In_97,In_1163);
nand U1167 (N_1167,In_1697,In_2449);
nor U1168 (N_1168,In_365,In_2560);
xnor U1169 (N_1169,In_1853,In_2994);
nor U1170 (N_1170,In_1421,In_1078);
nand U1171 (N_1171,In_2750,In_2700);
and U1172 (N_1172,In_1002,In_2928);
nor U1173 (N_1173,In_1903,In_900);
xnor U1174 (N_1174,In_487,In_2628);
or U1175 (N_1175,In_1067,In_2262);
nand U1176 (N_1176,In_73,In_940);
nor U1177 (N_1177,In_712,In_873);
nor U1178 (N_1178,In_810,In_787);
nand U1179 (N_1179,In_1403,In_2297);
xor U1180 (N_1180,In_1145,In_1383);
and U1181 (N_1181,In_1671,In_1400);
xnor U1182 (N_1182,In_1603,In_1390);
or U1183 (N_1183,In_2175,In_938);
or U1184 (N_1184,In_980,In_2844);
and U1185 (N_1185,In_1720,In_2017);
xnor U1186 (N_1186,In_422,In_2493);
xnor U1187 (N_1187,In_902,In_2127);
and U1188 (N_1188,In_1993,In_1804);
nand U1189 (N_1189,In_750,In_1367);
nor U1190 (N_1190,In_2296,In_240);
or U1191 (N_1191,In_1275,In_1657);
nand U1192 (N_1192,In_1096,In_2526);
or U1193 (N_1193,In_715,In_2674);
xnor U1194 (N_1194,In_2108,In_2945);
nor U1195 (N_1195,In_2315,In_2884);
and U1196 (N_1196,In_1404,In_1001);
or U1197 (N_1197,In_194,In_1625);
xor U1198 (N_1198,In_816,In_2924);
nor U1199 (N_1199,In_1594,In_2540);
xnor U1200 (N_1200,N_160,In_2178);
nand U1201 (N_1201,In_1246,In_1342);
or U1202 (N_1202,N_599,N_81);
or U1203 (N_1203,N_504,In_2090);
or U1204 (N_1204,N_867,N_782);
or U1205 (N_1205,N_687,N_302);
and U1206 (N_1206,In_1216,N_366);
xor U1207 (N_1207,In_1192,N_532);
xnor U1208 (N_1208,N_702,N_669);
xor U1209 (N_1209,In_596,In_66);
and U1210 (N_1210,In_2512,In_186);
nor U1211 (N_1211,In_705,In_2288);
nor U1212 (N_1212,In_1966,In_2523);
or U1213 (N_1213,N_353,In_495);
nor U1214 (N_1214,N_730,N_995);
xnor U1215 (N_1215,N_817,N_246);
xor U1216 (N_1216,In_2503,In_258);
nor U1217 (N_1217,N_421,N_483);
or U1218 (N_1218,In_2458,In_2656);
nor U1219 (N_1219,N_398,In_1241);
and U1220 (N_1220,N_454,N_845);
and U1221 (N_1221,In_1109,N_462);
xor U1222 (N_1222,N_864,In_2869);
and U1223 (N_1223,In_246,N_701);
nand U1224 (N_1224,N_139,In_1869);
or U1225 (N_1225,N_666,N_191);
nand U1226 (N_1226,N_261,N_382);
xnor U1227 (N_1227,N_871,In_1375);
nand U1228 (N_1228,N_451,N_120);
or U1229 (N_1229,N_1052,N_99);
or U1230 (N_1230,N_314,N_329);
nor U1231 (N_1231,N_1070,In_803);
and U1232 (N_1232,In_937,In_2534);
xor U1233 (N_1233,In_1115,N_912);
nand U1234 (N_1234,N_1112,N_1002);
or U1235 (N_1235,N_40,In_2756);
and U1236 (N_1236,N_835,In_1158);
nand U1237 (N_1237,N_904,N_1072);
or U1238 (N_1238,In_1776,N_965);
or U1239 (N_1239,N_16,In_116);
xnor U1240 (N_1240,N_638,In_2224);
xor U1241 (N_1241,N_719,In_2261);
nor U1242 (N_1242,N_981,N_954);
and U1243 (N_1243,N_430,N_1049);
or U1244 (N_1244,N_596,In_36);
or U1245 (N_1245,N_976,N_1120);
or U1246 (N_1246,In_52,In_414);
xnor U1247 (N_1247,N_1163,N_791);
or U1248 (N_1248,In_2382,N_647);
nand U1249 (N_1249,In_2152,N_43);
nand U1250 (N_1250,N_998,N_873);
nor U1251 (N_1251,N_502,In_358);
nor U1252 (N_1252,N_259,N_569);
or U1253 (N_1253,In_2907,N_1177);
xor U1254 (N_1254,N_380,N_222);
nor U1255 (N_1255,In_1321,In_2215);
nand U1256 (N_1256,N_515,N_722);
nand U1257 (N_1257,N_1160,N_994);
and U1258 (N_1258,N_455,N_622);
nand U1259 (N_1259,N_834,N_882);
xnor U1260 (N_1260,N_452,N_399);
xor U1261 (N_1261,N_181,N_343);
and U1262 (N_1262,In_698,N_1044);
xnor U1263 (N_1263,N_793,N_768);
or U1264 (N_1264,N_582,N_943);
or U1265 (N_1265,N_264,N_615);
nand U1266 (N_1266,N_1,N_339);
nand U1267 (N_1267,N_975,N_748);
xnor U1268 (N_1268,In_2793,N_1111);
and U1269 (N_1269,N_223,In_804);
xor U1270 (N_1270,In_51,N_500);
and U1271 (N_1271,In_468,In_1502);
or U1272 (N_1272,In_357,N_86);
or U1273 (N_1273,In_1673,N_471);
nand U1274 (N_1274,In_1698,In_2785);
and U1275 (N_1275,N_270,N_870);
and U1276 (N_1276,N_1176,N_449);
nand U1277 (N_1277,N_1089,In_1187);
and U1278 (N_1278,In_2070,N_999);
xnor U1279 (N_1279,In_61,In_1929);
nor U1280 (N_1280,N_276,In_1500);
xnor U1281 (N_1281,In_528,N_378);
nand U1282 (N_1282,N_1050,In_1782);
or U1283 (N_1283,N_77,N_1100);
xnor U1284 (N_1284,N_36,In_1533);
nor U1285 (N_1285,N_485,N_1033);
xor U1286 (N_1286,In_976,N_62);
and U1287 (N_1287,N_589,N_1189);
nand U1288 (N_1288,N_224,N_699);
and U1289 (N_1289,N_88,N_128);
nor U1290 (N_1290,N_394,N_1198);
or U1291 (N_1291,N_73,N_584);
or U1292 (N_1292,N_671,N_1062);
xor U1293 (N_1293,N_374,N_266);
and U1294 (N_1294,In_805,In_1785);
or U1295 (N_1295,N_113,N_738);
and U1296 (N_1296,In_356,N_881);
nand U1297 (N_1297,N_244,N_918);
xnor U1298 (N_1298,In_1688,N_923);
and U1299 (N_1299,In_40,N_764);
nand U1300 (N_1300,In_1877,N_591);
nor U1301 (N_1301,N_733,N_587);
xor U1302 (N_1302,N_1084,In_2569);
xor U1303 (N_1303,N_635,In_643);
or U1304 (N_1304,In_323,In_1860);
or U1305 (N_1305,In_812,N_880);
and U1306 (N_1306,In_864,N_324);
nor U1307 (N_1307,N_650,In_35);
nor U1308 (N_1308,In_941,In_1003);
nand U1309 (N_1309,In_1709,In_1530);
or U1310 (N_1310,In_2433,In_842);
and U1311 (N_1311,N_356,In_1208);
xor U1312 (N_1312,In_70,N_872);
and U1313 (N_1313,In_2927,In_2037);
xor U1314 (N_1314,N_108,In_2517);
xor U1315 (N_1315,N_54,N_204);
nor U1316 (N_1316,In_1666,N_1031);
nand U1317 (N_1317,N_595,N_375);
xnor U1318 (N_1318,N_1180,In_1453);
and U1319 (N_1319,N_773,N_30);
and U1320 (N_1320,N_879,N_728);
or U1321 (N_1321,In_298,In_1870);
or U1322 (N_1322,In_2242,In_584);
nor U1323 (N_1323,N_1173,In_877);
xor U1324 (N_1324,In_1026,N_305);
and U1325 (N_1325,N_1028,N_875);
nor U1326 (N_1326,N_1011,In_518);
xnor U1327 (N_1327,N_39,N_1166);
nor U1328 (N_1328,N_1104,N_150);
xnor U1329 (N_1329,N_754,N_1135);
and U1330 (N_1330,N_291,N_713);
or U1331 (N_1331,N_654,In_1654);
nor U1332 (N_1332,N_933,N_422);
or U1333 (N_1333,In_1687,N_323);
and U1334 (N_1334,N_1014,N_1136);
xor U1335 (N_1335,In_817,N_1192);
and U1336 (N_1336,N_55,N_397);
nand U1337 (N_1337,N_388,N_1106);
or U1338 (N_1338,N_1199,In_378);
nor U1339 (N_1339,N_752,N_275);
nand U1340 (N_1340,N_783,N_673);
or U1341 (N_1341,N_288,N_556);
and U1342 (N_1342,In_1950,N_993);
and U1343 (N_1343,In_2137,In_432);
nand U1344 (N_1344,In_1700,N_517);
and U1345 (N_1345,N_693,N_403);
and U1346 (N_1346,In_1285,N_564);
xor U1347 (N_1347,In_2621,N_652);
xnor U1348 (N_1348,N_1172,N_1156);
nor U1349 (N_1349,N_306,N_670);
nor U1350 (N_1350,N_292,In_2727);
xor U1351 (N_1351,N_865,N_427);
or U1352 (N_1352,In_2538,In_1113);
nor U1353 (N_1353,In_2038,In_2804);
nor U1354 (N_1354,In_2595,N_174);
xnor U1355 (N_1355,N_828,N_957);
nand U1356 (N_1356,N_620,N_257);
xnor U1357 (N_1357,N_405,N_467);
and U1358 (N_1358,In_1166,N_117);
xnor U1359 (N_1359,In_1160,N_641);
or U1360 (N_1360,N_1035,N_262);
and U1361 (N_1361,N_802,N_804);
or U1362 (N_1362,In_2681,N_123);
or U1363 (N_1363,In_1649,In_2643);
xor U1364 (N_1364,In_179,In_403);
nor U1365 (N_1365,N_659,N_1041);
or U1366 (N_1366,In_399,N_1167);
nor U1367 (N_1367,N_66,N_481);
nor U1368 (N_1368,N_736,N_816);
and U1369 (N_1369,N_268,N_1138);
nor U1370 (N_1370,In_2772,In_1898);
nor U1371 (N_1371,In_1636,N_110);
xnor U1372 (N_1372,In_1803,N_526);
nor U1373 (N_1373,In_2008,In_1743);
nand U1374 (N_1374,N_94,N_1107);
and U1375 (N_1375,N_11,In_1724);
nand U1376 (N_1376,In_2346,N_617);
or U1377 (N_1377,N_971,N_586);
and U1378 (N_1378,N_235,In_1011);
and U1379 (N_1379,N_778,N_445);
nor U1380 (N_1380,N_157,In_882);
nand U1381 (N_1381,In_2831,In_122);
and U1382 (N_1382,N_206,N_1094);
and U1383 (N_1383,In_86,N_285);
nand U1384 (N_1384,N_632,N_920);
or U1385 (N_1385,In_780,In_344);
nor U1386 (N_1386,N_103,N_333);
or U1387 (N_1387,N_968,N_508);
and U1388 (N_1388,N_861,N_938);
and U1389 (N_1389,N_898,N_1145);
and U1390 (N_1390,N_249,N_1001);
nor U1391 (N_1391,N_482,In_307);
nor U1392 (N_1392,N_487,In_26);
or U1393 (N_1393,N_739,In_2410);
xnor U1394 (N_1394,N_169,N_274);
and U1395 (N_1395,N_195,N_1130);
nand U1396 (N_1396,N_646,N_136);
nor U1397 (N_1397,N_948,N_46);
xnor U1398 (N_1398,N_400,In_2900);
xnor U1399 (N_1399,In_210,N_147);
nor U1400 (N_1400,N_714,N_829);
nor U1401 (N_1401,N_218,N_831);
nand U1402 (N_1402,In_1606,N_688);
and U1403 (N_1403,N_255,N_37);
or U1404 (N_1404,N_325,N_964);
or U1405 (N_1405,N_740,N_958);
and U1406 (N_1406,In_2767,N_900);
nor U1407 (N_1407,In_649,In_2684);
or U1408 (N_1408,N_886,In_2720);
nand U1409 (N_1409,N_51,N_548);
xnor U1410 (N_1410,N_827,N_242);
nand U1411 (N_1411,In_287,N_196);
nor U1412 (N_1412,N_769,In_1238);
xor U1413 (N_1413,In_2481,N_417);
nand U1414 (N_1414,N_784,N_844);
and U1415 (N_1415,N_1165,In_2103);
nor U1416 (N_1416,In_602,In_572);
xor U1417 (N_1417,N_734,N_364);
xor U1418 (N_1418,In_1961,N_735);
nor U1419 (N_1419,N_1054,N_580);
and U1420 (N_1420,In_291,In_2228);
xnor U1421 (N_1421,In_1419,N_499);
nor U1422 (N_1422,N_603,N_818);
nor U1423 (N_1423,N_685,In_1887);
or U1424 (N_1424,N_168,N_220);
nand U1425 (N_1425,In_2468,N_840);
or U1426 (N_1426,N_199,In_1486);
nand U1427 (N_1427,N_210,In_895);
nand U1428 (N_1428,N_205,In_32);
nor U1429 (N_1429,In_1987,N_284);
xnor U1430 (N_1430,N_917,N_707);
and U1431 (N_1431,N_572,In_1270);
xor U1432 (N_1432,N_749,In_1551);
and U1433 (N_1433,In_1683,In_2702);
and U1434 (N_1434,N_496,N_408);
nor U1435 (N_1435,N_522,N_830);
nor U1436 (N_1436,N_423,N_667);
or U1437 (N_1437,N_858,N_248);
xor U1438 (N_1438,N_35,N_1093);
nand U1439 (N_1439,N_428,N_294);
nor U1440 (N_1440,N_1197,N_521);
nor U1441 (N_1441,In_1191,N_1042);
nand U1442 (N_1442,N_145,In_351);
or U1443 (N_1443,In_762,N_212);
or U1444 (N_1444,N_989,N_955);
or U1445 (N_1445,N_1046,In_1706);
nor U1446 (N_1446,N_1127,In_1046);
xnor U1447 (N_1447,N_348,In_897);
or U1448 (N_1448,In_1102,N_1003);
or U1449 (N_1449,N_1187,In_2147);
nand U1450 (N_1450,N_71,N_1150);
and U1451 (N_1451,N_686,N_878);
and U1452 (N_1452,In_2018,N_772);
or U1453 (N_1453,N_100,In_1169);
and U1454 (N_1454,In_942,N_1096);
nor U1455 (N_1455,N_712,N_672);
nor U1456 (N_1456,N_345,N_661);
or U1457 (N_1457,N_849,N_890);
xor U1458 (N_1458,N_273,N_524);
nor U1459 (N_1459,In_2556,N_1038);
nor U1460 (N_1460,N_497,N_407);
xnor U1461 (N_1461,N_1015,N_729);
nor U1462 (N_1462,In_1827,N_1051);
nor U1463 (N_1463,N_997,In_2006);
nor U1464 (N_1464,In_1269,N_527);
nor U1465 (N_1465,N_133,In_1949);
nand U1466 (N_1466,N_59,N_1139);
nor U1467 (N_1467,N_961,In_277);
nand U1468 (N_1468,N_21,In_479);
nand U1469 (N_1469,N_1109,N_156);
and U1470 (N_1470,N_935,N_990);
or U1471 (N_1471,N_799,In_2347);
xnor U1472 (N_1472,N_1058,In_1143);
xnor U1473 (N_1473,N_540,N_1085);
or U1474 (N_1474,N_553,In_1351);
and U1475 (N_1475,N_444,N_1018);
and U1476 (N_1476,N_316,N_1076);
and U1477 (N_1477,In_2915,In_474);
xor U1478 (N_1478,In_1103,N_230);
and U1479 (N_1479,In_413,In_2245);
nand U1480 (N_1480,N_87,In_2145);
or U1481 (N_1481,N_613,N_1114);
and U1482 (N_1482,N_393,N_1005);
and U1483 (N_1483,In_1630,N_950);
and U1484 (N_1484,N_796,N_822);
xor U1485 (N_1485,N_490,N_811);
nor U1486 (N_1486,N_1040,N_1190);
xor U1487 (N_1487,In_1851,N_1128);
nand U1488 (N_1488,N_947,N_1142);
nor U1489 (N_1489,In_2447,In_1723);
xor U1490 (N_1490,N_897,In_1591);
xor U1491 (N_1491,In_255,In_1820);
and U1492 (N_1492,N_69,In_393);
or U1493 (N_1493,In_1972,N_575);
and U1494 (N_1494,N_1153,N_583);
or U1495 (N_1495,N_89,In_682);
and U1496 (N_1496,N_215,In_1523);
xor U1497 (N_1497,In_561,N_1086);
or U1498 (N_1498,N_863,In_2563);
nand U1499 (N_1499,N_543,N_727);
nand U1500 (N_1500,N_511,N_328);
nor U1501 (N_1501,N_1095,In_1775);
or U1502 (N_1502,N_1023,N_327);
or U1503 (N_1503,In_1835,N_760);
xnor U1504 (N_1504,N_109,N_578);
xnor U1505 (N_1505,In_872,N_1077);
or U1506 (N_1506,In_1126,In_2707);
xor U1507 (N_1507,N_124,N_234);
nand U1508 (N_1508,N_724,N_982);
xnor U1509 (N_1509,N_624,N_544);
nand U1510 (N_1510,In_1960,N_286);
or U1511 (N_1511,N_555,N_547);
xor U1512 (N_1512,In_1788,N_1055);
nand U1513 (N_1513,In_2822,In_2085);
nand U1514 (N_1514,N_194,N_446);
xor U1515 (N_1515,In_1436,In_2054);
nor U1516 (N_1516,In_2761,In_133);
and U1517 (N_1517,N_237,N_902);
or U1518 (N_1518,N_792,In_2723);
or U1519 (N_1519,In_2301,In_2695);
nor U1520 (N_1520,In_1133,N_49);
nand U1521 (N_1521,N_869,N_163);
or U1522 (N_1522,N_833,In_2933);
and U1523 (N_1523,N_579,N_370);
nor U1524 (N_1524,N_585,In_1370);
xnor U1525 (N_1525,N_1144,N_634);
nor U1526 (N_1526,N_211,In_118);
nor U1527 (N_1527,N_885,N_576);
nand U1528 (N_1528,N_131,In_2871);
nand U1529 (N_1529,N_1182,N_1008);
nand U1530 (N_1530,In_2766,N_1140);
xor U1531 (N_1531,In_1527,N_1073);
nand U1532 (N_1532,N_936,N_172);
nor U1533 (N_1533,N_402,N_1191);
or U1534 (N_1534,In_1816,In_1938);
or U1535 (N_1535,N_1091,N_1045);
nand U1536 (N_1536,N_1117,In_2672);
or U1537 (N_1537,N_921,N_637);
xnor U1538 (N_1538,N_6,N_926);
nand U1539 (N_1539,N_1057,N_705);
xor U1540 (N_1540,N_653,In_1401);
or U1541 (N_1541,In_2849,N_299);
or U1542 (N_1542,In_520,N_821);
nor U1543 (N_1543,N_1066,N_358);
nor U1544 (N_1544,N_91,In_1520);
xnor U1545 (N_1545,N_192,In_366);
or U1546 (N_1546,N_552,In_10);
nand U1547 (N_1547,In_1283,N_254);
nor U1548 (N_1548,N_594,In_2914);
and U1549 (N_1549,In_707,In_2460);
xnor U1550 (N_1550,N_491,In_1056);
nand U1551 (N_1551,N_1168,In_921);
nor U1552 (N_1552,N_330,N_910);
nand U1553 (N_1553,N_1185,N_847);
nor U1554 (N_1554,N_605,In_1702);
nor U1555 (N_1555,N_520,N_866);
xor U1556 (N_1556,N_777,N_992);
nand U1557 (N_1557,N_352,In_918);
and U1558 (N_1558,In_2403,N_533);
nor U1559 (N_1559,N_484,N_309);
xor U1560 (N_1560,N_310,N_1159);
and U1561 (N_1561,N_1092,N_34);
nor U1562 (N_1562,In_990,In_2172);
nand U1563 (N_1563,N_618,N_95);
nand U1564 (N_1564,N_281,N_265);
nand U1565 (N_1565,In_485,In_1976);
nand U1566 (N_1566,N_813,In_653);
xor U1567 (N_1567,N_241,N_751);
nor U1568 (N_1568,N_604,N_726);
and U1569 (N_1569,N_381,In_1118);
xor U1570 (N_1570,In_2072,In_141);
xnor U1571 (N_1571,N_465,N_282);
nand U1572 (N_1572,N_801,N_290);
and U1573 (N_1573,N_38,N_560);
or U1574 (N_1574,N_794,N_848);
nand U1575 (N_1575,N_1157,N_107);
xor U1576 (N_1576,N_621,N_806);
xor U1577 (N_1577,N_283,N_1119);
and U1578 (N_1578,N_1088,N_563);
and U1579 (N_1579,N_689,N_628);
or U1580 (N_1580,N_14,N_922);
and U1581 (N_1581,N_308,In_2490);
nand U1582 (N_1582,In_564,N_437);
and U1583 (N_1583,N_410,N_477);
or U1584 (N_1584,In_702,N_721);
nor U1585 (N_1585,N_140,N_342);
xor U1586 (N_1586,N_93,N_72);
xnor U1587 (N_1587,N_814,N_453);
or U1588 (N_1588,N_789,In_223);
nor U1589 (N_1589,In_956,In_1650);
or U1590 (N_1590,In_412,In_2067);
and U1591 (N_1591,In_2867,N_747);
nor U1592 (N_1592,In_2819,In_2118);
nand U1593 (N_1593,N_256,N_1030);
nand U1594 (N_1594,In_111,N_984);
nor U1595 (N_1595,In_1221,N_0);
or U1596 (N_1596,N_159,N_297);
or U1597 (N_1597,In_729,N_495);
nor U1598 (N_1598,N_153,N_611);
or U1599 (N_1599,N_279,N_1059);
nand U1600 (N_1600,N_1053,In_740);
xor U1601 (N_1601,In_2748,N_494);
or U1602 (N_1602,N_565,N_27);
xnor U1603 (N_1603,In_2323,N_676);
and U1604 (N_1604,N_385,N_1026);
nand U1605 (N_1605,N_529,In_734);
and U1606 (N_1606,N_326,N_44);
xor U1607 (N_1607,N_208,N_1056);
nor U1608 (N_1608,N_643,N_1069);
xor U1609 (N_1609,N_919,In_601);
and U1610 (N_1610,N_807,In_1779);
and U1611 (N_1611,In_2931,In_696);
and U1612 (N_1612,N_67,In_149);
nand U1613 (N_1613,N_966,In_567);
nand U1614 (N_1614,N_797,In_2393);
nand U1615 (N_1615,N_505,N_319);
nand U1616 (N_1616,In_2326,N_190);
nor U1617 (N_1617,In_749,In_272);
or U1618 (N_1618,N_1024,In_2949);
nand U1619 (N_1619,N_226,N_447);
nand U1620 (N_1620,In_589,N_790);
or U1621 (N_1621,N_629,N_606);
nor U1622 (N_1622,In_743,N_636);
nor U1623 (N_1623,N_365,N_602);
or U1624 (N_1624,N_28,N_404);
nand U1625 (N_1625,N_221,N_130);
nand U1626 (N_1626,In_1134,In_425);
or U1627 (N_1627,N_1075,In_2350);
or U1628 (N_1628,N_1132,N_351);
nor U1629 (N_1629,In_491,N_1151);
xnor U1630 (N_1630,N_680,N_271);
or U1631 (N_1631,N_568,In_683);
or U1632 (N_1632,N_825,N_937);
nor U1633 (N_1633,In_923,In_834);
xor U1634 (N_1634,In_193,In_2640);
or U1635 (N_1635,In_599,N_1013);
or U1636 (N_1636,N_1020,In_2635);
and U1637 (N_1637,N_280,In_476);
nor U1638 (N_1638,N_229,In_641);
and U1639 (N_1639,N_144,N_57);
nor U1640 (N_1640,N_625,N_362);
xnor U1641 (N_1641,N_173,In_404);
or U1642 (N_1642,In_1213,In_2453);
xor U1643 (N_1643,N_842,In_752);
or U1644 (N_1644,N_367,N_859);
and U1645 (N_1645,N_703,N_903);
nor U1646 (N_1646,N_1000,N_750);
or U1647 (N_1647,In_1313,In_1838);
nand U1648 (N_1648,N_389,N_985);
or U1649 (N_1649,N_1186,N_909);
nand U1650 (N_1650,N_941,N_972);
nor U1651 (N_1651,N_468,N_774);
nor U1652 (N_1652,N_64,N_1036);
nor U1653 (N_1653,In_388,N_126);
xnor U1654 (N_1654,N_476,In_1910);
nor U1655 (N_1655,N_90,In_1485);
nand U1656 (N_1656,In_110,N_313);
xor U1657 (N_1657,N_247,N_68);
and U1658 (N_1658,N_812,N_376);
nand U1659 (N_1659,In_822,In_2508);
nand U1660 (N_1660,In_367,N_83);
and U1661 (N_1661,In_2069,In_802);
nor U1662 (N_1662,In_2739,N_597);
or U1663 (N_1663,N_186,N_631);
and U1664 (N_1664,N_1090,In_2221);
and U1665 (N_1665,N_457,In_2805);
and U1666 (N_1666,N_787,In_2180);
nand U1667 (N_1667,In_1613,N_470);
nand U1668 (N_1668,N_781,N_409);
or U1669 (N_1669,N_369,N_3);
nor U1670 (N_1670,In_1258,N_690);
or U1671 (N_1671,N_45,N_762);
or U1672 (N_1672,N_655,N_47);
and U1673 (N_1673,N_1006,N_354);
or U1674 (N_1674,N_331,N_26);
nand U1675 (N_1675,N_295,In_701);
and U1676 (N_1676,N_820,N_127);
or U1677 (N_1677,N_1115,N_1147);
nor U1678 (N_1678,N_359,In_2610);
nor U1679 (N_1679,N_856,N_278);
or U1680 (N_1680,In_175,N_289);
nor U1681 (N_1681,N_58,N_207);
and U1682 (N_1682,N_657,In_670);
nor U1683 (N_1683,N_542,In_1299);
and U1684 (N_1684,N_826,N_303);
nand U1685 (N_1685,N_709,In_2498);
or U1686 (N_1686,N_75,N_927);
nand U1687 (N_1687,N_1032,N_70);
and U1688 (N_1688,N_1068,N_1061);
xnor U1689 (N_1689,In_137,N_969);
and U1690 (N_1690,N_925,In_2418);
xnor U1691 (N_1691,In_1971,In_2056);
nand U1692 (N_1692,In_2316,N_1101);
nor U1693 (N_1693,In_182,In_1895);
xnor U1694 (N_1694,N_945,In_1517);
or U1695 (N_1695,N_805,In_947);
or U1696 (N_1696,N_433,N_486);
or U1697 (N_1697,N_24,In_1686);
or U1698 (N_1698,N_612,N_236);
or U1699 (N_1699,N_779,In_678);
nand U1700 (N_1700,In_1428,N_570);
nor U1701 (N_1701,N_355,In_1616);
xor U1702 (N_1702,N_135,N_554);
xor U1703 (N_1703,N_1078,N_932);
xnor U1704 (N_1704,N_610,In_453);
or U1705 (N_1705,N_1010,In_2524);
nor U1706 (N_1706,In_677,N_665);
nand U1707 (N_1707,N_121,N_25);
nor U1708 (N_1708,In_2990,In_950);
nor U1709 (N_1709,N_755,N_415);
xnor U1710 (N_1710,N_1118,In_2002);
nand U1711 (N_1711,N_1082,N_346);
or U1712 (N_1712,In_2608,N_883);
nor U1713 (N_1713,In_2354,N_891);
and U1714 (N_1714,In_1992,In_516);
or U1715 (N_1715,N_1125,N_488);
or U1716 (N_1716,N_383,N_48);
or U1717 (N_1717,N_301,In_2698);
or U1718 (N_1718,N_341,N_7);
and U1719 (N_1719,N_668,N_8);
nand U1720 (N_1720,N_913,N_691);
xnor U1721 (N_1721,In_1288,N_498);
and U1722 (N_1722,In_1984,N_166);
xnor U1723 (N_1723,N_1105,N_238);
and U1724 (N_1724,N_846,N_823);
or U1725 (N_1725,N_737,In_2220);
nand U1726 (N_1726,In_1564,N_837);
xor U1727 (N_1727,In_2892,N_183);
or U1728 (N_1728,N_1080,N_179);
or U1729 (N_1729,N_84,N_175);
nor U1730 (N_1730,In_1340,N_1021);
and U1731 (N_1731,N_798,N_377);
and U1732 (N_1732,In_511,N_396);
and U1733 (N_1733,In_519,In_1849);
nand U1734 (N_1734,N_164,N_122);
nand U1735 (N_1735,N_766,N_559);
xor U1736 (N_1736,N_105,N_116);
or U1737 (N_1737,N_1143,In_2974);
and U1738 (N_1738,N_908,N_843);
nor U1739 (N_1739,N_1162,In_1677);
xor U1740 (N_1740,N_536,N_340);
xnor U1741 (N_1741,N_928,N_267);
xnor U1742 (N_1742,N_137,N_627);
and U1743 (N_1743,N_17,In_1420);
nand U1744 (N_1744,In_2094,N_65);
nor U1745 (N_1745,N_19,In_2501);
or U1746 (N_1746,In_961,N_272);
nand U1747 (N_1747,N_677,In_166);
and U1748 (N_1748,N_360,In_1035);
xnor U1749 (N_1749,N_874,In_675);
xnor U1750 (N_1750,N_700,In_2314);
and U1751 (N_1751,N_639,N_616);
and U1752 (N_1752,N_475,N_79);
or U1753 (N_1753,N_887,N_1116);
or U1754 (N_1754,N_56,N_456);
nor U1755 (N_1755,In_2779,N_431);
and U1756 (N_1756,N_862,In_1371);
nor U1757 (N_1757,N_151,In_646);
and U1758 (N_1758,In_785,N_710);
nand U1759 (N_1759,N_836,In_2661);
nor U1760 (N_1760,In_633,N_277);
xnor U1761 (N_1761,N_15,N_307);
xor U1762 (N_1762,In_1257,N_518);
or U1763 (N_1763,N_649,N_97);
or U1764 (N_1764,N_414,N_217);
xnor U1765 (N_1765,In_2383,In_1979);
or U1766 (N_1766,In_301,In_660);
nor U1767 (N_1767,N_300,In_1110);
or U1768 (N_1768,In_2759,N_630);
and U1769 (N_1769,N_82,N_788);
and U1770 (N_1770,N_1074,In_355);
nor U1771 (N_1771,N_20,N_899);
nand U1772 (N_1772,N_371,In_1329);
xor U1773 (N_1773,In_2535,N_780);
and U1774 (N_1774,In_1301,N_104);
nor U1775 (N_1775,In_1934,In_2363);
nand U1776 (N_1776,N_549,In_1469);
xnor U1777 (N_1777,N_269,N_379);
nand U1778 (N_1778,In_607,N_18);
or U1779 (N_1779,N_744,N_696);
or U1780 (N_1780,In_311,N_1048);
xor U1781 (N_1781,In_813,In_1973);
and U1782 (N_1782,N_1170,N_1131);
or U1783 (N_1783,N_986,In_741);
nand U1784 (N_1784,In_2734,N_537);
nand U1785 (N_1785,N_525,N_441);
xnor U1786 (N_1786,N_391,N_197);
and U1787 (N_1787,N_503,In_2429);
xor U1788 (N_1788,N_893,N_1154);
or U1789 (N_1789,N_96,N_1141);
nand U1790 (N_1790,In_2231,N_763);
nor U1791 (N_1791,N_233,In_1656);
nor U1792 (N_1792,N_895,N_562);
and U1793 (N_1793,N_979,In_2733);
nand U1794 (N_1794,N_940,In_274);
and U1795 (N_1795,N_347,In_1690);
xnor U1796 (N_1796,N_853,In_639);
nor U1797 (N_1797,In_171,In_1868);
nor U1798 (N_1798,In_455,In_1442);
or U1799 (N_1799,N_854,N_809);
and U1800 (N_1800,N_1171,N_1029);
or U1801 (N_1801,N_1043,N_1194);
nor U1802 (N_1802,In_461,In_580);
xor U1803 (N_1803,N_142,N_440);
nor U1804 (N_1804,N_581,N_996);
nor U1805 (N_1805,N_63,N_138);
nand U1806 (N_1806,N_170,N_74);
xor U1807 (N_1807,N_1158,N_715);
nand U1808 (N_1808,N_795,In_2369);
nand U1809 (N_1809,In_2184,N_1065);
and U1810 (N_1810,N_1017,N_258);
or U1811 (N_1811,N_474,N_78);
nor U1812 (N_1812,In_2851,N_930);
nor U1813 (N_1813,N_492,N_232);
and U1814 (N_1814,N_571,N_171);
and U1815 (N_1815,N_761,In_2408);
nor U1816 (N_1816,N_149,In_1618);
nand U1817 (N_1817,N_1146,N_227);
or U1818 (N_1818,In_1627,In_2947);
and U1819 (N_1819,In_2291,N_557);
xnor U1820 (N_1820,N_711,N_681);
nor U1821 (N_1821,In_41,N_460);
nand U1822 (N_1822,N_479,N_13);
nor U1823 (N_1823,In_1071,N_970);
nor U1824 (N_1824,N_439,N_425);
or U1825 (N_1825,In_1424,N_450);
nand U1826 (N_1826,In_1670,N_253);
or U1827 (N_1827,In_328,In_1121);
and U1828 (N_1828,N_52,N_245);
xor U1829 (N_1829,N_911,In_909);
nor U1830 (N_1830,N_839,In_1364);
and U1831 (N_1831,N_785,N_1184);
nand U1832 (N_1832,N_395,N_832);
or U1833 (N_1833,In_421,N_601);
or U1834 (N_1834,N_401,N_694);
and U1835 (N_1835,N_448,N_438);
or U1836 (N_1836,In_1361,In_215);
nand U1837 (N_1837,N_112,In_104);
xnor U1838 (N_1838,In_489,N_501);
xnor U1839 (N_1839,In_2889,N_771);
or U1840 (N_1840,N_651,In_505);
xnor U1841 (N_1841,In_1038,In_169);
nand U1842 (N_1842,N_12,In_1620);
and U1843 (N_1843,N_623,In_2477);
nand U1844 (N_1844,In_2728,In_2488);
xnor U1845 (N_1845,In_1728,N_459);
nand U1846 (N_1846,In_103,N_706);
and U1847 (N_1847,N_1183,N_1129);
and U1848 (N_1848,N_419,In_1386);
nor U1849 (N_1849,N_952,N_411);
nor U1850 (N_1850,N_368,In_693);
and U1851 (N_1851,N_42,In_146);
or U1852 (N_1852,N_593,In_2097);
xnor U1853 (N_1853,In_2165,N_683);
xnor U1854 (N_1854,N_810,N_384);
xnor U1855 (N_1855,N_412,N_600);
or U1856 (N_1856,N_723,N_929);
nor U1857 (N_1857,In_385,N_519);
nor U1858 (N_1858,N_682,N_1103);
nor U1859 (N_1859,In_2703,N_541);
nor U1860 (N_1860,In_1040,N_478);
nand U1861 (N_1861,N_1037,N_658);
nor U1862 (N_1862,In_346,N_119);
nor U1863 (N_1863,N_531,N_363);
and U1864 (N_1864,N_155,N_1148);
and U1865 (N_1865,N_588,In_338);
nor U1866 (N_1866,N_1034,N_420);
or U1867 (N_1867,In_2790,In_2480);
nand U1868 (N_1868,N_298,N_5);
nand U1869 (N_1869,N_263,N_956);
or U1870 (N_1870,In_1255,In_19);
nor U1871 (N_1871,In_690,N_225);
or U1872 (N_1872,In_2170,N_535);
nand U1873 (N_1873,N_1016,N_332);
and U1874 (N_1874,In_970,In_2360);
and U1875 (N_1875,N_214,In_1378);
and U1876 (N_1876,N_534,N_745);
nor U1877 (N_1877,N_551,In_1508);
and U1878 (N_1878,In_2908,N_1175);
or U1879 (N_1879,In_2162,In_623);
and U1880 (N_1880,In_2872,N_857);
nand U1881 (N_1881,N_894,In_1474);
nand U1882 (N_1882,N_590,N_513);
nand U1883 (N_1883,In_91,N_435);
nand U1884 (N_1884,N_1009,In_1655);
and U1885 (N_1885,In_815,N_732);
and U1886 (N_1886,In_1806,N_901);
and U1887 (N_1887,N_1098,N_296);
nor U1888 (N_1888,N_426,N_767);
or U1889 (N_1889,N_1087,N_198);
nand U1890 (N_1890,N_697,N_905);
nand U1891 (N_1891,N_480,N_931);
nand U1892 (N_1892,In_515,N_387);
xor U1893 (N_1893,N_318,N_60);
nand U1894 (N_1894,N_143,N_50);
nand U1895 (N_1895,In_1366,N_592);
nor U1896 (N_1896,In_2267,N_201);
or U1897 (N_1897,In_739,N_915);
and U1898 (N_1898,In_2758,N_640);
nand U1899 (N_1899,In_2959,In_2331);
and U1900 (N_1900,In_1162,N_720);
and U1901 (N_1901,N_188,In_1320);
xnor U1902 (N_1902,In_2367,N_538);
and U1903 (N_1903,N_1004,N_974);
or U1904 (N_1904,In_405,N_656);
nor U1905 (N_1905,In_2771,N_158);
xnor U1906 (N_1906,N_200,N_493);
xnor U1907 (N_1907,N_41,N_775);
nand U1908 (N_1908,N_31,N_203);
nor U1909 (N_1909,In_1230,N_10);
xor U1910 (N_1910,N_1071,N_959);
or U1911 (N_1911,N_1178,N_663);
or U1912 (N_1912,N_608,N_489);
and U1913 (N_1913,N_9,N_988);
and U1914 (N_1914,In_410,N_182);
nor U1915 (N_1915,In_934,In_667);
and U1916 (N_1916,In_1405,In_1922);
or U1917 (N_1917,N_889,In_1182);
nand U1918 (N_1918,N_704,In_1888);
and U1919 (N_1919,N_1027,N_413);
xor U1920 (N_1920,N_1022,In_390);
and U1921 (N_1921,N_934,In_135);
nor U1922 (N_1922,N_106,In_1108);
xor U1923 (N_1923,N_692,N_1019);
xor U1924 (N_1924,In_2348,In_1186);
nand U1925 (N_1925,N_841,N_577);
and U1926 (N_1926,N_980,N_176);
xor U1927 (N_1927,In_130,N_573);
nand U1928 (N_1928,In_33,In_1812);
nor U1929 (N_1929,N_101,N_824);
nor U1930 (N_1930,N_434,N_154);
nor U1931 (N_1931,N_287,N_1133);
nor U1932 (N_1932,N_418,N_293);
nor U1933 (N_1933,N_357,In_2390);
and U1934 (N_1934,N_546,In_845);
and U1935 (N_1935,N_759,N_662);
nor U1936 (N_1936,In_428,In_1426);
xor U1937 (N_1937,N_507,N_209);
and U1938 (N_1938,N_416,N_219);
xor U1939 (N_1939,N_1047,N_260);
nor U1940 (N_1940,N_1181,In_2737);
xor U1941 (N_1941,N_1102,N_1108);
xor U1942 (N_1942,N_963,In_1136);
and U1943 (N_1943,N_178,N_946);
or U1944 (N_1944,In_318,N_252);
nand U1945 (N_1945,N_725,N_320);
or U1946 (N_1946,N_906,In_2738);
and U1947 (N_1947,N_896,N_888);
nor U1948 (N_1948,In_119,In_647);
nand U1949 (N_1949,In_924,N_466);
xnor U1950 (N_1950,N_731,N_148);
xor U1951 (N_1951,In_2574,N_758);
nor U1952 (N_1952,N_916,In_447);
nor U1953 (N_1953,N_660,In_1223);
or U1954 (N_1954,In_831,N_819);
and U1955 (N_1955,In_597,N_202);
nor U1956 (N_1956,In_1454,In_1524);
xor U1957 (N_1957,N_1169,N_469);
xnor U1958 (N_1958,N_32,In_1081);
and U1959 (N_1959,In_1932,N_1063);
and U1960 (N_1960,N_962,N_372);
xnor U1961 (N_1961,In_2374,N_852);
xor U1962 (N_1962,N_185,N_523);
and U1963 (N_1963,N_1193,N_770);
xor U1964 (N_1964,In_1178,In_1129);
xor U1965 (N_1965,N_1097,N_216);
and U1966 (N_1966,N_180,In_1501);
nor U1967 (N_1967,N_162,N_803);
nor U1968 (N_1968,N_33,In_914);
and U1969 (N_1969,N_776,In_1206);
nor U1970 (N_1970,N_619,N_1149);
and U1971 (N_1971,N_876,In_44);
nor U1972 (N_1972,In_493,N_228);
nand U1973 (N_1973,N_115,N_321);
xnor U1974 (N_1974,N_386,N_574);
xnor U1975 (N_1975,N_167,N_392);
and U1976 (N_1976,N_53,N_22);
xor U1977 (N_1977,In_409,N_1123);
and U1978 (N_1978,In_192,N_815);
or U1979 (N_1979,N_1121,In_1639);
xor U1980 (N_1980,N_165,N_684);
and U1981 (N_1981,N_808,N_1137);
and U1982 (N_1982,In_309,N_1134);
or U1983 (N_1983,N_1174,In_1253);
nor U1984 (N_1984,N_757,N_29);
xnor U1985 (N_1985,N_92,In_2800);
nand U1986 (N_1986,N_80,N_1064);
or U1987 (N_1987,In_2587,N_951);
xor U1988 (N_1988,N_860,N_967);
nand U1989 (N_1989,N_344,N_98);
nand U1990 (N_1990,N_765,In_438);
or U1991 (N_1991,N_977,N_464);
and U1992 (N_1992,N_424,In_2434);
nand U1993 (N_1993,In_2121,In_2568);
nor U1994 (N_1994,N_1164,N_509);
nor U1995 (N_1995,N_373,In_1930);
nor U1996 (N_1996,N_558,N_61);
xor U1997 (N_1997,In_212,In_2562);
nor U1998 (N_1998,N_545,N_742);
nand U1999 (N_1999,N_1152,N_1110);
nand U2000 (N_2000,N_23,N_1196);
nand U2001 (N_2001,In_2857,N_1161);
and U2002 (N_2002,In_1662,N_1195);
or U2003 (N_2003,N_1126,N_1122);
xnor U2004 (N_2004,In_2668,In_958);
nand U2005 (N_2005,N_213,N_125);
xor U2006 (N_2006,N_1188,N_550);
nor U2007 (N_2007,In_2126,N_1007);
nand U2008 (N_2008,N_516,In_2027);
nor U2009 (N_2009,In_265,N_675);
xnor U2010 (N_2010,N_978,N_716);
nand U2011 (N_2011,In_74,In_981);
nand U2012 (N_2012,N_111,N_800);
and U2013 (N_2013,N_892,N_1179);
xor U2014 (N_2014,N_877,N_187);
and U2015 (N_2015,In_2874,N_626);
or U2016 (N_2016,N_1099,N_753);
xor U2017 (N_2017,In_2818,In_433);
or U2018 (N_2018,N_114,N_991);
or U2019 (N_2019,In_2168,In_2642);
nor U2020 (N_2020,In_2821,N_924);
and U2021 (N_2021,In_2378,N_1155);
xor U2022 (N_2022,In_2269,In_71);
nor U2023 (N_2023,N_786,N_461);
or U2024 (N_2024,N_1113,N_695);
or U2025 (N_2025,N_949,N_746);
nand U2026 (N_2026,N_1081,In_2898);
and U2027 (N_2027,N_193,N_614);
nor U2028 (N_2028,N_506,N_458);
nand U2029 (N_2029,N_134,N_1067);
nand U2030 (N_2030,N_645,N_1025);
or U2031 (N_2031,N_609,N_708);
or U2032 (N_2032,N_189,In_1197);
xnor U2033 (N_2033,N_472,N_250);
nor U2034 (N_2034,N_850,N_907);
or U2035 (N_2035,N_251,N_1060);
and U2036 (N_2036,N_851,In_1717);
or U2037 (N_2037,In_2706,N_304);
nand U2038 (N_2038,N_129,N_855);
nor U2039 (N_2039,N_960,N_336);
xnor U2040 (N_2040,N_436,In_2814);
nor U2041 (N_2041,N_2,In_933);
nor U2042 (N_2042,N_648,N_674);
and U2043 (N_2043,N_1083,N_349);
and U2044 (N_2044,N_315,N_334);
xnor U2045 (N_2045,N_184,N_231);
and U2046 (N_2046,In_100,N_561);
and U2047 (N_2047,N_717,N_530);
and U2048 (N_2048,N_642,N_914);
xnor U2049 (N_2049,N_678,N_607);
and U2050 (N_2050,N_361,N_335);
nor U2051 (N_2051,N_146,N_442);
nand U2052 (N_2052,N_161,N_510);
and U2053 (N_2053,N_406,N_514);
or U2054 (N_2054,N_432,In_1311);
or U2055 (N_2055,N_239,N_1012);
nand U2056 (N_2056,N_633,N_756);
xor U2057 (N_2057,N_152,N_4);
or U2058 (N_2058,N_743,N_102);
nand U2059 (N_2059,In_94,N_1124);
xnor U2060 (N_2060,In_2240,N_1039);
xor U2061 (N_2061,In_2663,N_567);
and U2062 (N_2062,N_644,N_942);
and U2063 (N_2063,In_936,In_466);
or U2064 (N_2064,N_337,N_566);
and U2065 (N_2065,In_1750,N_939);
or U2066 (N_2066,N_322,In_1862);
xnor U2067 (N_2067,N_429,N_698);
xor U2068 (N_2068,In_1259,N_240);
nor U2069 (N_2069,N_338,In_1732);
or U2070 (N_2070,In_630,N_718);
or U2071 (N_2071,N_473,In_1041);
xor U2072 (N_2072,In_2467,N_664);
nor U2073 (N_2073,N_944,In_39);
or U2074 (N_2074,N_973,N_443);
or U2075 (N_2075,N_528,In_609);
xor U2076 (N_2076,N_312,In_426);
and U2077 (N_2077,In_557,N_76);
nand U2078 (N_2078,In_2979,N_1079);
and U2079 (N_2079,In_892,In_2581);
nor U2080 (N_2080,N_463,In_2609);
nor U2081 (N_2081,N_350,In_452);
or U2082 (N_2082,N_838,N_679);
xnor U2083 (N_2083,In_987,N_987);
nor U2084 (N_2084,N_983,In_789);
xor U2085 (N_2085,N_118,N_85);
and U2086 (N_2086,N_177,In_2745);
or U2087 (N_2087,N_741,In_978);
and U2088 (N_2088,N_598,In_929);
or U2089 (N_2089,In_1395,N_243);
or U2090 (N_2090,In_2451,N_512);
nor U2091 (N_2091,In_2013,N_953);
nand U2092 (N_2092,N_317,In_1051);
nand U2093 (N_2093,N_311,N_141);
nand U2094 (N_2094,N_539,N_884);
nand U2095 (N_2095,In_2971,N_390);
nor U2096 (N_2096,N_132,In_454);
xor U2097 (N_2097,In_1459,In_198);
or U2098 (N_2098,In_2306,N_868);
and U2099 (N_2099,In_2721,In_22);
nand U2100 (N_2100,N_551,In_2301);
xor U2101 (N_2101,N_49,N_448);
nor U2102 (N_2102,N_157,In_2168);
nand U2103 (N_2103,N_755,In_1690);
or U2104 (N_2104,N_1029,In_2054);
nand U2105 (N_2105,N_360,In_1238);
xnor U2106 (N_2106,In_785,N_284);
nand U2107 (N_2107,N_51,N_957);
nor U2108 (N_2108,N_970,N_482);
or U2109 (N_2109,N_379,N_32);
nand U2110 (N_2110,N_1180,N_287);
and U2111 (N_2111,N_1137,N_621);
nor U2112 (N_2112,N_1053,N_465);
or U2113 (N_2113,N_218,In_2433);
xnor U2114 (N_2114,N_5,N_23);
and U2115 (N_2115,N_1191,N_1130);
nor U2116 (N_2116,In_602,In_1424);
nor U2117 (N_2117,N_617,N_818);
xor U2118 (N_2118,N_392,N_558);
nor U2119 (N_2119,N_545,N_767);
nor U2120 (N_2120,In_455,N_227);
and U2121 (N_2121,N_973,N_609);
nand U2122 (N_2122,N_1100,In_897);
nor U2123 (N_2123,N_723,N_371);
xnor U2124 (N_2124,N_355,N_3);
or U2125 (N_2125,N_327,N_1092);
nand U2126 (N_2126,N_179,N_1129);
and U2127 (N_2127,In_2346,N_938);
nand U2128 (N_2128,N_348,N_961);
nor U2129 (N_2129,In_485,N_195);
nor U2130 (N_2130,N_465,N_852);
or U2131 (N_2131,In_734,In_2165);
and U2132 (N_2132,N_34,In_1370);
and U2133 (N_2133,N_480,In_2556);
or U2134 (N_2134,N_493,N_994);
nor U2135 (N_2135,N_551,N_1001);
or U2136 (N_2136,N_986,In_1375);
or U2137 (N_2137,In_1551,N_636);
nor U2138 (N_2138,N_780,N_326);
nand U2139 (N_2139,N_632,N_886);
nor U2140 (N_2140,N_257,N_92);
and U2141 (N_2141,N_1105,N_1137);
nand U2142 (N_2142,In_1788,In_909);
nor U2143 (N_2143,N_556,N_417);
or U2144 (N_2144,N_818,N_1010);
and U2145 (N_2145,In_1253,In_2002);
and U2146 (N_2146,N_205,N_52);
or U2147 (N_2147,In_941,In_981);
nor U2148 (N_2148,In_1011,N_975);
nor U2149 (N_2149,N_807,N_339);
or U2150 (N_2150,N_1098,N_185);
nand U2151 (N_2151,N_51,In_2027);
and U2152 (N_2152,N_387,In_409);
or U2153 (N_2153,N_896,In_987);
nand U2154 (N_2154,N_1118,N_1026);
or U2155 (N_2155,N_823,N_344);
and U2156 (N_2156,In_212,N_684);
nand U2157 (N_2157,In_2085,N_759);
xor U2158 (N_2158,In_2503,N_1173);
nor U2159 (N_2159,In_2374,N_283);
and U2160 (N_2160,In_740,In_1683);
xor U2161 (N_2161,N_1018,In_2090);
or U2162 (N_2162,N_1196,In_2006);
nor U2163 (N_2163,In_1630,N_418);
nor U2164 (N_2164,In_468,N_1152);
or U2165 (N_2165,N_8,N_1159);
xnor U2166 (N_2166,N_784,N_949);
xor U2167 (N_2167,In_749,N_105);
xnor U2168 (N_2168,N_840,In_2288);
xnor U2169 (N_2169,N_1122,N_260);
xnor U2170 (N_2170,N_94,N_795);
and U2171 (N_2171,N_221,N_413);
or U2172 (N_2172,In_432,N_239);
or U2173 (N_2173,N_9,N_1124);
xnor U2174 (N_2174,In_2267,N_351);
nand U2175 (N_2175,In_933,N_1123);
or U2176 (N_2176,N_288,N_770);
and U2177 (N_2177,N_311,N_389);
or U2178 (N_2178,In_1109,In_1454);
and U2179 (N_2179,N_922,N_511);
xnor U2180 (N_2180,N_495,N_1176);
and U2181 (N_2181,N_699,N_879);
nand U2182 (N_2182,N_1199,In_1564);
nor U2183 (N_2183,In_698,In_171);
and U2184 (N_2184,N_195,In_749);
nand U2185 (N_2185,In_2734,N_337);
or U2186 (N_2186,N_1196,In_2971);
nor U2187 (N_2187,N_45,N_37);
and U2188 (N_2188,N_1129,N_844);
nand U2189 (N_2189,In_1639,In_2990);
nor U2190 (N_2190,N_345,N_1044);
and U2191 (N_2191,N_866,N_519);
xnor U2192 (N_2192,In_831,N_807);
nor U2193 (N_2193,N_96,N_1122);
nor U2194 (N_2194,N_250,N_1185);
xor U2195 (N_2195,In_609,N_397);
xor U2196 (N_2196,N_314,In_1081);
xor U2197 (N_2197,N_1035,In_2871);
nand U2198 (N_2198,N_439,N_985);
xnor U2199 (N_2199,N_786,In_2458);
or U2200 (N_2200,In_2524,N_228);
nand U2201 (N_2201,N_1132,N_1175);
or U2202 (N_2202,In_32,N_126);
xor U2203 (N_2203,N_712,In_2085);
xnor U2204 (N_2204,In_1654,N_1045);
xor U2205 (N_2205,N_743,N_691);
xor U2206 (N_2206,In_1564,In_2508);
nor U2207 (N_2207,N_1174,In_2346);
nor U2208 (N_2208,N_123,N_1048);
nor U2209 (N_2209,N_234,N_1095);
nand U2210 (N_2210,N_880,N_931);
xor U2211 (N_2211,In_51,N_1072);
nand U2212 (N_2212,N_892,N_1178);
and U2213 (N_2213,N_128,N_386);
or U2214 (N_2214,In_924,N_733);
or U2215 (N_2215,N_502,In_291);
or U2216 (N_2216,N_1025,N_27);
xor U2217 (N_2217,In_2306,N_1157);
nand U2218 (N_2218,N_336,N_814);
xor U2219 (N_2219,In_1371,In_1688);
nand U2220 (N_2220,In_2738,N_1010);
xor U2221 (N_2221,In_2501,In_1820);
nor U2222 (N_2222,In_66,N_1068);
nor U2223 (N_2223,N_288,In_822);
nand U2224 (N_2224,N_630,N_522);
and U2225 (N_2225,In_1386,In_198);
or U2226 (N_2226,N_1036,N_815);
nand U2227 (N_2227,N_1119,In_1785);
nand U2228 (N_2228,In_2737,N_120);
xnor U2229 (N_2229,N_25,N_1157);
or U2230 (N_2230,N_1119,N_1023);
or U2231 (N_2231,In_2242,N_717);
nand U2232 (N_2232,N_375,N_621);
nand U2233 (N_2233,N_20,In_2069);
xor U2234 (N_2234,N_617,In_707);
nor U2235 (N_2235,N_1011,In_2738);
xor U2236 (N_2236,N_329,In_596);
nand U2237 (N_2237,N_764,In_897);
xnor U2238 (N_2238,N_795,In_1270);
xnor U2239 (N_2239,N_429,In_277);
or U2240 (N_2240,In_2447,N_851);
or U2241 (N_2241,N_358,N_301);
or U2242 (N_2242,In_643,N_660);
xnor U2243 (N_2243,N_437,In_2538);
nor U2244 (N_2244,N_72,N_819);
and U2245 (N_2245,In_914,N_559);
nor U2246 (N_2246,In_179,N_34);
nor U2247 (N_2247,N_357,In_1938);
nand U2248 (N_2248,N_567,N_1010);
or U2249 (N_2249,N_106,N_687);
and U2250 (N_2250,In_71,N_486);
and U2251 (N_2251,In_1961,N_173);
or U2252 (N_2252,N_891,N_683);
and U2253 (N_2253,N_277,In_1401);
and U2254 (N_2254,N_98,In_1378);
or U2255 (N_2255,N_766,N_872);
nor U2256 (N_2256,In_990,In_1743);
and U2257 (N_2257,N_57,In_1639);
or U2258 (N_2258,In_2301,N_707);
and U2259 (N_2259,In_2793,N_521);
nand U2260 (N_2260,N_476,N_495);
xnor U2261 (N_2261,N_410,N_702);
xor U2262 (N_2262,N_1038,In_328);
xor U2263 (N_2263,N_422,N_746);
nor U2264 (N_2264,In_338,In_2979);
or U2265 (N_2265,In_580,In_1938);
nand U2266 (N_2266,In_357,N_1172);
and U2267 (N_2267,N_364,In_1630);
and U2268 (N_2268,N_269,N_1085);
or U2269 (N_2269,N_48,N_436);
nand U2270 (N_2270,N_1147,N_454);
xor U2271 (N_2271,N_450,In_1340);
and U2272 (N_2272,N_982,N_472);
nor U2273 (N_2273,In_2698,N_272);
or U2274 (N_2274,In_1108,N_625);
or U2275 (N_2275,N_1092,In_2172);
or U2276 (N_2276,In_1253,N_477);
nand U2277 (N_2277,In_351,N_906);
xnor U2278 (N_2278,In_1929,N_406);
or U2279 (N_2279,In_2793,In_39);
and U2280 (N_2280,In_272,In_1115);
nor U2281 (N_2281,In_1442,N_1076);
xnor U2282 (N_2282,N_462,In_1040);
xor U2283 (N_2283,N_131,In_1670);
nand U2284 (N_2284,N_126,N_1120);
xnor U2285 (N_2285,In_198,N_630);
xor U2286 (N_2286,N_746,In_1666);
nand U2287 (N_2287,N_731,N_1033);
or U2288 (N_2288,N_694,N_403);
xnor U2289 (N_2289,N_768,In_2610);
or U2290 (N_2290,N_842,N_107);
nor U2291 (N_2291,N_963,N_723);
nor U2292 (N_2292,N_446,N_826);
nor U2293 (N_2293,In_2867,N_235);
xnor U2294 (N_2294,N_758,N_227);
and U2295 (N_2295,In_1246,N_278);
or U2296 (N_2296,N_252,N_19);
nor U2297 (N_2297,In_2672,N_118);
nor U2298 (N_2298,In_1424,In_1606);
nor U2299 (N_2299,In_520,N_132);
nor U2300 (N_2300,In_653,N_1039);
nor U2301 (N_2301,N_178,N_485);
nand U2302 (N_2302,In_179,In_1930);
nor U2303 (N_2303,In_2734,N_542);
xor U2304 (N_2304,N_109,N_326);
and U2305 (N_2305,N_55,N_273);
xnor U2306 (N_2306,N_2,N_817);
and U2307 (N_2307,N_278,In_609);
nand U2308 (N_2308,In_2346,N_172);
or U2309 (N_2309,N_664,In_2556);
or U2310 (N_2310,N_166,N_727);
nand U2311 (N_2311,N_1051,N_348);
nor U2312 (N_2312,N_474,In_1420);
nor U2313 (N_2313,N_701,N_1025);
or U2314 (N_2314,N_832,In_2772);
nor U2315 (N_2315,In_2569,N_225);
nand U2316 (N_2316,In_2642,N_926);
or U2317 (N_2317,N_278,In_505);
xnor U2318 (N_2318,N_22,N_142);
nand U2319 (N_2319,In_2707,N_853);
and U2320 (N_2320,N_620,N_1047);
nor U2321 (N_2321,N_379,N_317);
or U2322 (N_2322,N_476,In_485);
or U2323 (N_2323,N_838,In_1134);
nor U2324 (N_2324,N_286,In_1620);
or U2325 (N_2325,In_2314,N_989);
or U2326 (N_2326,In_2242,In_309);
and U2327 (N_2327,In_19,In_660);
xnor U2328 (N_2328,N_394,N_968);
nand U2329 (N_2329,N_571,N_666);
nand U2330 (N_2330,In_2759,In_1527);
or U2331 (N_2331,In_678,N_867);
xnor U2332 (N_2332,N_76,In_2538);
or U2333 (N_2333,In_1501,In_476);
and U2334 (N_2334,In_1869,N_559);
nor U2335 (N_2335,N_134,N_791);
or U2336 (N_2336,N_1006,N_332);
xor U2337 (N_2337,N_852,In_2363);
and U2338 (N_2338,In_528,N_1075);
nand U2339 (N_2339,In_2974,N_624);
xor U2340 (N_2340,In_701,N_678);
nand U2341 (N_2341,N_696,N_587);
nor U2342 (N_2342,N_146,N_853);
nand U2343 (N_2343,N_466,N_410);
and U2344 (N_2344,N_449,N_702);
nor U2345 (N_2345,N_1140,N_326);
nor U2346 (N_2346,N_1139,In_298);
or U2347 (N_2347,N_53,In_2184);
nand U2348 (N_2348,N_746,N_542);
nand U2349 (N_2349,N_1060,In_1230);
nand U2350 (N_2350,In_2090,N_1196);
or U2351 (N_2351,In_942,In_607);
nor U2352 (N_2352,In_19,N_1180);
and U2353 (N_2353,N_781,N_403);
nand U2354 (N_2354,N_1039,N_434);
nand U2355 (N_2355,N_535,N_369);
and U2356 (N_2356,N_376,In_1930);
nand U2357 (N_2357,In_1186,N_1131);
nor U2358 (N_2358,In_2587,N_190);
xor U2359 (N_2359,In_1655,N_797);
and U2360 (N_2360,In_40,N_35);
nor U2361 (N_2361,N_543,N_883);
or U2362 (N_2362,N_86,In_1041);
xor U2363 (N_2363,N_511,N_843);
nor U2364 (N_2364,N_966,In_1129);
nand U2365 (N_2365,N_483,N_1140);
xnor U2366 (N_2366,N_283,In_1806);
or U2367 (N_2367,N_371,N_160);
and U2368 (N_2368,N_288,N_435);
or U2369 (N_2369,N_489,N_1066);
or U2370 (N_2370,N_501,N_558);
or U2371 (N_2371,N_1056,In_2067);
and U2372 (N_2372,N_330,In_2306);
nand U2373 (N_2373,N_234,N_811);
or U2374 (N_2374,N_230,N_958);
nor U2375 (N_2375,N_51,In_461);
nand U2376 (N_2376,In_584,In_182);
xnor U2377 (N_2377,N_172,N_174);
nor U2378 (N_2378,In_351,N_461);
and U2379 (N_2379,N_36,N_276);
and U2380 (N_2380,In_1690,In_1166);
nand U2381 (N_2381,N_776,In_515);
and U2382 (N_2382,In_116,N_488);
nand U2383 (N_2383,In_432,In_356);
nand U2384 (N_2384,N_183,N_683);
and U2385 (N_2385,N_97,In_2524);
and U2386 (N_2386,In_683,N_877);
xnor U2387 (N_2387,N_520,In_2508);
nand U2388 (N_2388,N_1125,N_351);
or U2389 (N_2389,N_922,N_789);
and U2390 (N_2390,In_414,N_285);
nor U2391 (N_2391,In_493,In_2706);
nand U2392 (N_2392,N_1025,N_1151);
xor U2393 (N_2393,In_1887,In_2267);
and U2394 (N_2394,N_1178,N_392);
or U2395 (N_2395,N_28,In_2907);
or U2396 (N_2396,N_1047,N_251);
xnor U2397 (N_2397,N_655,N_1119);
xor U2398 (N_2398,N_990,N_622);
nor U2399 (N_2399,N_20,N_571);
xnor U2400 (N_2400,N_1674,N_1698);
or U2401 (N_2401,N_1491,N_1310);
or U2402 (N_2402,N_1495,N_2243);
xor U2403 (N_2403,N_1224,N_1581);
or U2404 (N_2404,N_1549,N_2035);
or U2405 (N_2405,N_2022,N_1213);
nand U2406 (N_2406,N_1919,N_1514);
and U2407 (N_2407,N_1616,N_1667);
xor U2408 (N_2408,N_2359,N_2394);
xnor U2409 (N_2409,N_2048,N_1364);
nor U2410 (N_2410,N_1947,N_1992);
or U2411 (N_2411,N_2121,N_2315);
and U2412 (N_2412,N_2361,N_1650);
xor U2413 (N_2413,N_1524,N_1681);
xor U2414 (N_2414,N_2202,N_1417);
xor U2415 (N_2415,N_1365,N_2137);
and U2416 (N_2416,N_1265,N_1436);
xor U2417 (N_2417,N_2319,N_1571);
and U2418 (N_2418,N_1857,N_2061);
nor U2419 (N_2419,N_1932,N_2024);
or U2420 (N_2420,N_1915,N_2172);
nor U2421 (N_2421,N_1295,N_1880);
and U2422 (N_2422,N_1411,N_2264);
nor U2423 (N_2423,N_2195,N_1718);
nor U2424 (N_2424,N_1999,N_1447);
xor U2425 (N_2425,N_1225,N_1207);
xnor U2426 (N_2426,N_2377,N_1774);
or U2427 (N_2427,N_2108,N_2041);
nor U2428 (N_2428,N_1872,N_2118);
nand U2429 (N_2429,N_1676,N_1652);
nor U2430 (N_2430,N_1744,N_1507);
and U2431 (N_2431,N_2102,N_1541);
xor U2432 (N_2432,N_1559,N_1734);
nor U2433 (N_2433,N_1501,N_1474);
nor U2434 (N_2434,N_1697,N_1901);
nand U2435 (N_2435,N_1771,N_1457);
nor U2436 (N_2436,N_2020,N_1463);
xor U2437 (N_2437,N_1211,N_1287);
xnor U2438 (N_2438,N_1424,N_1658);
nand U2439 (N_2439,N_1831,N_2381);
and U2440 (N_2440,N_2105,N_1728);
xor U2441 (N_2441,N_2258,N_2182);
nand U2442 (N_2442,N_1439,N_1939);
xor U2443 (N_2443,N_2331,N_1819);
or U2444 (N_2444,N_1952,N_2047);
and U2445 (N_2445,N_2357,N_2200);
nor U2446 (N_2446,N_2310,N_1407);
nor U2447 (N_2447,N_2327,N_2301);
nor U2448 (N_2448,N_1512,N_2360);
xnor U2449 (N_2449,N_2274,N_2367);
nor U2450 (N_2450,N_1725,N_1714);
nor U2451 (N_2451,N_1742,N_1889);
nand U2452 (N_2452,N_1982,N_1375);
nor U2453 (N_2453,N_1597,N_1309);
or U2454 (N_2454,N_2294,N_1875);
nor U2455 (N_2455,N_1660,N_1589);
nand U2456 (N_2456,N_1285,N_2368);
nor U2457 (N_2457,N_1325,N_1200);
xor U2458 (N_2458,N_2006,N_2343);
xnor U2459 (N_2459,N_1591,N_1927);
nand U2460 (N_2460,N_1551,N_2208);
and U2461 (N_2461,N_1790,N_1839);
nand U2462 (N_2462,N_2144,N_1260);
nor U2463 (N_2463,N_2322,N_1866);
or U2464 (N_2464,N_1764,N_1894);
xnor U2465 (N_2465,N_1754,N_1973);
xnor U2466 (N_2466,N_1640,N_1232);
nand U2467 (N_2467,N_1523,N_2211);
and U2468 (N_2468,N_1532,N_1777);
or U2469 (N_2469,N_1422,N_1203);
nor U2470 (N_2470,N_2028,N_1689);
xnor U2471 (N_2471,N_2250,N_2193);
and U2472 (N_2472,N_1922,N_1553);
nor U2473 (N_2473,N_1712,N_1311);
and U2474 (N_2474,N_2371,N_2189);
nand U2475 (N_2475,N_2127,N_1598);
xnor U2476 (N_2476,N_1482,N_1497);
xor U2477 (N_2477,N_2037,N_1477);
nand U2478 (N_2478,N_1829,N_1958);
nor U2479 (N_2479,N_2308,N_1427);
nand U2480 (N_2480,N_1432,N_1678);
nand U2481 (N_2481,N_2186,N_2387);
nor U2482 (N_2482,N_1420,N_1705);
nand U2483 (N_2483,N_1394,N_2054);
nor U2484 (N_2484,N_1582,N_2346);
nand U2485 (N_2485,N_1277,N_1624);
and U2486 (N_2486,N_2194,N_2318);
nand U2487 (N_2487,N_1851,N_2109);
xor U2488 (N_2488,N_1242,N_2052);
and U2489 (N_2489,N_2192,N_1672);
nand U2490 (N_2490,N_2207,N_2071);
xor U2491 (N_2491,N_2075,N_2154);
nor U2492 (N_2492,N_2266,N_1960);
nand U2493 (N_2493,N_1812,N_1655);
nand U2494 (N_2494,N_1446,N_2043);
nor U2495 (N_2495,N_1994,N_1703);
nor U2496 (N_2496,N_1273,N_2215);
nor U2497 (N_2497,N_1679,N_1910);
xnor U2498 (N_2498,N_2003,N_1688);
nand U2499 (N_2499,N_1649,N_2130);
xnor U2500 (N_2500,N_1269,N_2333);
nor U2501 (N_2501,N_2117,N_2352);
xnor U2502 (N_2502,N_1465,N_1349);
and U2503 (N_2503,N_2085,N_2285);
nand U2504 (N_2504,N_1564,N_1770);
and U2505 (N_2505,N_1896,N_2252);
nand U2506 (N_2506,N_2302,N_2027);
nor U2507 (N_2507,N_1493,N_1330);
and U2508 (N_2508,N_1879,N_1271);
nor U2509 (N_2509,N_1617,N_1805);
or U2510 (N_2510,N_1724,N_1266);
and U2511 (N_2511,N_2222,N_1782);
nand U2512 (N_2512,N_1909,N_2067);
and U2513 (N_2513,N_2083,N_1270);
or U2514 (N_2514,N_1443,N_1802);
nor U2515 (N_2515,N_1510,N_1248);
nor U2516 (N_2516,N_1558,N_2004);
xnor U2517 (N_2517,N_2279,N_1766);
and U2518 (N_2518,N_1838,N_1205);
xnor U2519 (N_2519,N_1995,N_2198);
or U2520 (N_2520,N_1907,N_1721);
and U2521 (N_2521,N_1942,N_2009);
nor U2522 (N_2522,N_2389,N_1586);
xnor U2523 (N_2523,N_1404,N_1540);
nor U2524 (N_2524,N_2213,N_1595);
nand U2525 (N_2525,N_1292,N_1428);
nor U2526 (N_2526,N_1405,N_2374);
nor U2527 (N_2527,N_2380,N_1733);
nand U2528 (N_2528,N_1353,N_1560);
xnor U2529 (N_2529,N_2175,N_2087);
and U2530 (N_2530,N_2058,N_1302);
xor U2531 (N_2531,N_1326,N_2183);
and U2532 (N_2532,N_1344,N_2397);
or U2533 (N_2533,N_1904,N_1578);
nor U2534 (N_2534,N_1367,N_2265);
nand U2535 (N_2535,N_1717,N_1882);
nand U2536 (N_2536,N_1884,N_1487);
nor U2537 (N_2537,N_1971,N_2206);
and U2538 (N_2538,N_2365,N_2016);
xor U2539 (N_2539,N_1221,N_2219);
nand U2540 (N_2540,N_1410,N_1833);
or U2541 (N_2541,N_1625,N_2057);
xnor U2542 (N_2542,N_1788,N_1228);
nand U2543 (N_2543,N_1740,N_2214);
xnor U2544 (N_2544,N_1888,N_1425);
nor U2545 (N_2545,N_2307,N_1779);
or U2546 (N_2546,N_1263,N_1637);
xor U2547 (N_2547,N_1303,N_1609);
nand U2548 (N_2548,N_1227,N_2291);
xor U2549 (N_2549,N_1281,N_1464);
or U2550 (N_2550,N_1210,N_2148);
and U2551 (N_2551,N_1669,N_2204);
nor U2552 (N_2552,N_2078,N_1408);
nor U2553 (N_2553,N_1562,N_1935);
nand U2554 (N_2554,N_2312,N_1409);
nor U2555 (N_2555,N_2014,N_1731);
nand U2556 (N_2556,N_1216,N_1602);
and U2557 (N_2557,N_1715,N_2306);
nor U2558 (N_2558,N_2018,N_1557);
or U2559 (N_2559,N_1887,N_1906);
and U2560 (N_2560,N_2284,N_1352);
and U2561 (N_2561,N_2034,N_1478);
nor U2562 (N_2562,N_1944,N_1504);
or U2563 (N_2563,N_1950,N_2349);
xnor U2564 (N_2564,N_1778,N_1822);
nor U2565 (N_2565,N_1686,N_1677);
and U2566 (N_2566,N_2293,N_1521);
xor U2567 (N_2567,N_1253,N_2277);
nand U2568 (N_2568,N_1750,N_1945);
xnor U2569 (N_2569,N_1238,N_1614);
xor U2570 (N_2570,N_2382,N_1985);
and U2571 (N_2571,N_1418,N_2229);
and U2572 (N_2572,N_2228,N_1671);
and U2573 (N_2573,N_1461,N_1986);
nor U2574 (N_2574,N_1575,N_2069);
nor U2575 (N_2575,N_2303,N_2158);
xnor U2576 (N_2576,N_1351,N_2248);
nand U2577 (N_2577,N_1648,N_1403);
xor U2578 (N_2578,N_2205,N_2399);
xnor U2579 (N_2579,N_1892,N_1923);
xor U2580 (N_2580,N_2116,N_1948);
nor U2581 (N_2581,N_1545,N_1389);
nor U2582 (N_2582,N_1834,N_1605);
nor U2583 (N_2583,N_1955,N_2029);
or U2584 (N_2584,N_1479,N_2000);
nor U2585 (N_2585,N_1444,N_2039);
nor U2586 (N_2586,N_1716,N_1296);
nor U2587 (N_2587,N_2131,N_2155);
and U2588 (N_2588,N_1918,N_1555);
nand U2589 (N_2589,N_2090,N_1241);
nor U2590 (N_2590,N_1594,N_1630);
xnor U2591 (N_2591,N_1746,N_1550);
xor U2592 (N_2592,N_1247,N_1612);
nor U2593 (N_2593,N_2030,N_1621);
or U2594 (N_2594,N_1662,N_1996);
or U2595 (N_2595,N_1818,N_2120);
and U2596 (N_2596,N_1385,N_1204);
or U2597 (N_2597,N_2230,N_1930);
and U2598 (N_2598,N_1406,N_1758);
or U2599 (N_2599,N_2050,N_1755);
xor U2600 (N_2600,N_2084,N_1291);
or U2601 (N_2601,N_1828,N_1651);
nor U2602 (N_2602,N_1267,N_2281);
nand U2603 (N_2603,N_1951,N_1704);
nand U2604 (N_2604,N_1587,N_1864);
and U2605 (N_2605,N_1636,N_2336);
nand U2606 (N_2606,N_1334,N_2358);
and U2607 (N_2607,N_1577,N_1552);
nor U2608 (N_2608,N_1978,N_1530);
nor U2609 (N_2609,N_1329,N_2031);
and U2610 (N_2610,N_1868,N_1264);
and U2611 (N_2611,N_2356,N_2385);
nor U2612 (N_2612,N_1230,N_1469);
nand U2613 (N_2613,N_1460,N_2282);
nand U2614 (N_2614,N_1869,N_1747);
or U2615 (N_2615,N_2073,N_1272);
and U2616 (N_2616,N_2151,N_2095);
nor U2617 (N_2617,N_1438,N_2236);
nand U2618 (N_2618,N_2077,N_1664);
and U2619 (N_2619,N_1807,N_1974);
xor U2620 (N_2620,N_1471,N_1539);
or U2621 (N_2621,N_1261,N_1252);
nor U2622 (N_2622,N_1765,N_1933);
nand U2623 (N_2623,N_1223,N_2150);
nor U2624 (N_2624,N_2044,N_1572);
nand U2625 (N_2625,N_2383,N_1596);
and U2626 (N_2626,N_2156,N_1583);
nor U2627 (N_2627,N_1492,N_1769);
nand U2628 (N_2628,N_1941,N_1361);
or U2629 (N_2629,N_1376,N_1903);
xor U2630 (N_2630,N_2386,N_1354);
xor U2631 (N_2631,N_1599,N_1244);
or U2632 (N_2632,N_2142,N_2096);
xnor U2633 (N_2633,N_1984,N_1484);
nand U2634 (N_2634,N_1339,N_2159);
or U2635 (N_2635,N_1761,N_1600);
nor U2636 (N_2636,N_1250,N_1610);
nor U2637 (N_2637,N_1396,N_1897);
or U2638 (N_2638,N_1350,N_1543);
xor U2639 (N_2639,N_1706,N_1623);
and U2640 (N_2640,N_1297,N_1258);
or U2641 (N_2641,N_1360,N_2124);
nand U2642 (N_2642,N_2176,N_2045);
and U2643 (N_2643,N_1229,N_1423);
nor U2644 (N_2644,N_2099,N_2168);
or U2645 (N_2645,N_2246,N_1319);
and U2646 (N_2646,N_1519,N_1803);
and U2647 (N_2647,N_1659,N_1707);
nor U2648 (N_2648,N_2326,N_1816);
nor U2649 (N_2649,N_2086,N_1964);
or U2650 (N_2650,N_1215,N_1848);
and U2651 (N_2651,N_2316,N_1647);
and U2652 (N_2652,N_1231,N_2002);
xnor U2653 (N_2653,N_1787,N_1893);
nand U2654 (N_2654,N_1201,N_1826);
xnor U2655 (N_2655,N_1914,N_1379);
and U2656 (N_2656,N_2296,N_1535);
nand U2657 (N_2657,N_1499,N_2321);
nor U2658 (N_2658,N_2342,N_1874);
and U2659 (N_2659,N_2170,N_1214);
nor U2660 (N_2660,N_2049,N_1324);
xor U2661 (N_2661,N_1276,N_2239);
nand U2662 (N_2662,N_1369,N_1837);
nor U2663 (N_2663,N_1956,N_2276);
xnor U2664 (N_2664,N_1937,N_1318);
nand U2665 (N_2665,N_2169,N_1800);
nand U2666 (N_2666,N_1488,N_1794);
nand U2667 (N_2667,N_2253,N_1862);
nand U2668 (N_2668,N_2259,N_1395);
and U2669 (N_2669,N_1590,N_1462);
or U2670 (N_2670,N_2060,N_1926);
nor U2671 (N_2671,N_1431,N_2221);
xor U2672 (N_2672,N_2390,N_2132);
or U2673 (N_2673,N_1437,N_1502);
and U2674 (N_2674,N_1568,N_2079);
nand U2675 (N_2675,N_2227,N_1348);
and U2676 (N_2676,N_2181,N_1619);
xor U2677 (N_2677,N_1891,N_1286);
nor U2678 (N_2678,N_2335,N_1305);
nor U2679 (N_2679,N_1574,N_1554);
nand U2680 (N_2680,N_1936,N_1283);
xnor U2681 (N_2681,N_2249,N_2298);
nand U2682 (N_2682,N_2074,N_1454);
xnor U2683 (N_2683,N_1452,N_2262);
and U2684 (N_2684,N_1399,N_1653);
and U2685 (N_2685,N_1966,N_1314);
nor U2686 (N_2686,N_2015,N_1569);
or U2687 (N_2687,N_2313,N_1852);
and U2688 (N_2688,N_2149,N_1346);
or U2689 (N_2689,N_2097,N_1480);
nand U2690 (N_2690,N_1262,N_2345);
xor U2691 (N_2691,N_1856,N_2210);
or U2692 (N_2692,N_1998,N_1929);
and U2693 (N_2693,N_1824,N_2010);
or U2694 (N_2694,N_1692,N_2395);
nand U2695 (N_2695,N_1990,N_1799);
or U2696 (N_2696,N_1520,N_1741);
nand U2697 (N_2697,N_1206,N_1827);
or U2698 (N_2698,N_1924,N_2042);
xor U2699 (N_2699,N_2234,N_2070);
xnor U2700 (N_2700,N_1255,N_2201);
nand U2701 (N_2701,N_2292,N_1810);
xnor U2702 (N_2702,N_2147,N_1538);
nand U2703 (N_2703,N_1335,N_1342);
nand U2704 (N_2704,N_2379,N_1673);
or U2705 (N_2705,N_1748,N_1371);
nor U2706 (N_2706,N_1953,N_2072);
nor U2707 (N_2707,N_1784,N_2232);
nand U2708 (N_2708,N_2287,N_1737);
or U2709 (N_2709,N_1969,N_1912);
or U2710 (N_2710,N_2165,N_1976);
and U2711 (N_2711,N_2263,N_1668);
nor U2712 (N_2712,N_2290,N_2059);
xor U2713 (N_2713,N_1392,N_1202);
nor U2714 (N_2714,N_1208,N_2295);
xnor U2715 (N_2715,N_1975,N_2033);
nand U2716 (N_2716,N_1735,N_1886);
or U2717 (N_2717,N_2173,N_1486);
xnor U2718 (N_2718,N_2026,N_2375);
nor U2719 (N_2719,N_2089,N_2111);
xnor U2720 (N_2720,N_1435,N_1300);
or U2721 (N_2721,N_1282,N_1817);
and U2722 (N_2722,N_2320,N_1328);
nor U2723 (N_2723,N_2091,N_2348);
xor U2724 (N_2724,N_1475,N_1413);
and U2725 (N_2725,N_2212,N_2012);
nand U2726 (N_2726,N_1393,N_1633);
or U2727 (N_2727,N_1957,N_1792);
and U2728 (N_2728,N_1380,N_1307);
nor U2729 (N_2729,N_1383,N_1726);
nor U2730 (N_2730,N_1290,N_2261);
xnor U2731 (N_2731,N_1759,N_2330);
nor U2732 (N_2732,N_1845,N_2063);
or U2733 (N_2733,N_2216,N_1357);
and U2734 (N_2734,N_1615,N_1727);
nand U2735 (N_2735,N_1791,N_1738);
xor U2736 (N_2736,N_2220,N_2001);
xnor U2737 (N_2737,N_2135,N_1280);
nand U2738 (N_2738,N_1513,N_1752);
or U2739 (N_2739,N_1226,N_1340);
nor U2740 (N_2740,N_1949,N_1878);
xor U2741 (N_2741,N_1254,N_1983);
or U2742 (N_2742,N_1751,N_2324);
and U2743 (N_2743,N_1338,N_1279);
or U2744 (N_2744,N_1972,N_2092);
or U2745 (N_2745,N_1533,N_1299);
and U2746 (N_2746,N_1516,N_1362);
nor U2747 (N_2747,N_1565,N_1573);
or U2748 (N_2748,N_1821,N_1606);
nand U2749 (N_2749,N_2209,N_1666);
or U2750 (N_2750,N_1940,N_2280);
nor U2751 (N_2751,N_1327,N_2325);
nand U2752 (N_2752,N_2025,N_1331);
nand U2753 (N_2753,N_1494,N_2235);
nor U2754 (N_2754,N_1527,N_1576);
xor U2755 (N_2755,N_1531,N_1858);
and U2756 (N_2756,N_1278,N_2145);
xnor U2757 (N_2757,N_1968,N_2217);
or U2758 (N_2758,N_1908,N_2272);
nand U2759 (N_2759,N_1696,N_1489);
and U2760 (N_2760,N_1785,N_2143);
nand U2761 (N_2761,N_1243,N_2338);
xor U2762 (N_2762,N_1308,N_1854);
xnor U2763 (N_2763,N_1274,N_1959);
xnor U2764 (N_2764,N_2373,N_1702);
nor U2765 (N_2765,N_2218,N_1762);
nor U2766 (N_2766,N_2184,N_1517);
nor U2767 (N_2767,N_2032,N_1592);
and U2768 (N_2768,N_1401,N_2317);
nor U2769 (N_2769,N_1453,N_1629);
or U2770 (N_2770,N_1928,N_2370);
nand U2771 (N_2771,N_1775,N_1685);
nor U2772 (N_2772,N_2133,N_2203);
xor U2773 (N_2773,N_1256,N_1511);
nor U2774 (N_2774,N_1781,N_1840);
nand U2775 (N_2775,N_2340,N_1222);
and U2776 (N_2776,N_1467,N_1789);
or U2777 (N_2777,N_1895,N_1626);
nand U2778 (N_2778,N_1859,N_2115);
nand U2779 (N_2779,N_1806,N_2013);
xnor U2780 (N_2780,N_1776,N_2019);
xor U2781 (N_2781,N_2392,N_1289);
and U2782 (N_2782,N_2056,N_1301);
nand U2783 (N_2783,N_1402,N_2119);
or U2784 (N_2784,N_1341,N_1808);
nor U2785 (N_2785,N_1320,N_1240);
or U2786 (N_2786,N_1701,N_1743);
xor U2787 (N_2787,N_1963,N_1865);
and U2788 (N_2788,N_1470,N_1835);
or U2789 (N_2789,N_2093,N_2231);
or U2790 (N_2790,N_1451,N_2372);
and U2791 (N_2791,N_1783,N_1312);
nor U2792 (N_2792,N_1506,N_1275);
and U2793 (N_2793,N_1757,N_1796);
and U2794 (N_2794,N_2286,N_2337);
or U2795 (N_2795,N_1710,N_2196);
or U2796 (N_2796,N_2100,N_1529);
nor U2797 (N_2797,N_2341,N_1313);
xor U2798 (N_2798,N_2157,N_1580);
nor U2799 (N_2799,N_2134,N_1322);
and U2800 (N_2800,N_2354,N_1694);
nor U2801 (N_2801,N_1607,N_1217);
xnor U2802 (N_2802,N_2167,N_2297);
xor U2803 (N_2803,N_1246,N_1426);
nor U2804 (N_2804,N_2136,N_2362);
nand U2805 (N_2805,N_1245,N_1618);
or U2806 (N_2806,N_2023,N_2188);
nor U2807 (N_2807,N_1561,N_1695);
and U2808 (N_2808,N_1989,N_2081);
nand U2809 (N_2809,N_1306,N_2129);
and U2810 (N_2810,N_1873,N_2398);
nor U2811 (N_2811,N_1219,N_2139);
nor U2812 (N_2812,N_1472,N_2347);
nand U2813 (N_2813,N_2021,N_2256);
nor U2814 (N_2814,N_2241,N_2122);
and U2815 (N_2815,N_1547,N_1323);
nand U2816 (N_2816,N_2068,N_1525);
nor U2817 (N_2817,N_1683,N_2114);
and U2818 (N_2818,N_1358,N_1925);
nand U2819 (N_2819,N_1356,N_1294);
or U2820 (N_2820,N_1670,N_1251);
or U2821 (N_2821,N_1466,N_1793);
xor U2822 (N_2822,N_2244,N_2269);
and U2823 (N_2823,N_1509,N_2177);
nand U2824 (N_2824,N_2275,N_2128);
nor U2825 (N_2825,N_2160,N_1981);
nor U2826 (N_2826,N_1459,N_2270);
and U2827 (N_2827,N_2199,N_1642);
nor U2828 (N_2828,N_1212,N_1237);
or U2829 (N_2829,N_2245,N_1378);
or U2830 (N_2830,N_2353,N_1760);
and U2831 (N_2831,N_1730,N_2350);
nor U2832 (N_2832,N_2055,N_1987);
xnor U2833 (N_2833,N_1434,N_1913);
nor U2834 (N_2834,N_2088,N_1400);
and U2835 (N_2835,N_1421,N_1387);
nand U2836 (N_2836,N_2125,N_1911);
nor U2837 (N_2837,N_2267,N_2066);
xnor U2838 (N_2838,N_1699,N_1693);
and U2839 (N_2839,N_1566,N_1804);
xor U2840 (N_2840,N_2240,N_1458);
xnor U2841 (N_2841,N_1900,N_2179);
or U2842 (N_2842,N_1795,N_2251);
xnor U2843 (N_2843,N_2005,N_1259);
nor U2844 (N_2844,N_1544,N_1898);
or U2845 (N_2845,N_1797,N_1815);
xnor U2846 (N_2846,N_2299,N_1366);
nand U2847 (N_2847,N_1780,N_2110);
xnor U2848 (N_2848,N_2036,N_2314);
and U2849 (N_2849,N_1820,N_1801);
and U2850 (N_2850,N_1977,N_1496);
and U2851 (N_2851,N_2378,N_2393);
or U2852 (N_2852,N_1965,N_1415);
xnor U2853 (N_2853,N_1548,N_1390);
and U2854 (N_2854,N_1508,N_2164);
and U2855 (N_2855,N_2094,N_2053);
xor U2856 (N_2856,N_1691,N_1768);
or U2857 (N_2857,N_2141,N_2300);
and U2858 (N_2858,N_2007,N_2366);
nor U2859 (N_2859,N_1233,N_1388);
xnor U2860 (N_2860,N_1485,N_1877);
nand U2861 (N_2861,N_1481,N_1680);
nand U2862 (N_2862,N_1931,N_2185);
nor U2863 (N_2863,N_1773,N_1883);
nand U2864 (N_2864,N_2233,N_1736);
nand U2865 (N_2865,N_1249,N_2396);
and U2866 (N_2866,N_1628,N_1384);
nand U2867 (N_2867,N_1359,N_2344);
nand U2868 (N_2868,N_2082,N_2112);
nor U2869 (N_2869,N_2339,N_2101);
nand U2870 (N_2870,N_1841,N_2046);
or U2871 (N_2871,N_1811,N_1430);
nor U2872 (N_2872,N_1946,N_1528);
or U2873 (N_2873,N_1753,N_1732);
xnor U2874 (N_2874,N_2268,N_1885);
and U2875 (N_2875,N_1368,N_1518);
xnor U2876 (N_2876,N_2166,N_1473);
xor U2877 (N_2877,N_2311,N_2328);
nand U2878 (N_2878,N_2334,N_1515);
xnor U2879 (N_2879,N_1962,N_1814);
and U2880 (N_2880,N_1700,N_1445);
and U2881 (N_2881,N_1347,N_1345);
xor U2882 (N_2882,N_1961,N_2305);
nor U2883 (N_2883,N_1288,N_1522);
nand U2884 (N_2884,N_1611,N_1209);
nor U2885 (N_2885,N_2329,N_2288);
nand U2886 (N_2886,N_2038,N_1382);
or U2887 (N_2887,N_1656,N_1416);
or U2888 (N_2888,N_1620,N_1284);
nand U2889 (N_2889,N_2161,N_1321);
xor U2890 (N_2890,N_1970,N_2040);
nand U2891 (N_2891,N_1483,N_1690);
nand U2892 (N_2892,N_1863,N_1997);
nor U2893 (N_2893,N_2309,N_1468);
nor U2894 (N_2894,N_1682,N_1870);
nor U2895 (N_2895,N_1316,N_1739);
or U2896 (N_2896,N_2237,N_2107);
or U2897 (N_2897,N_1567,N_1967);
nor U2898 (N_2898,N_1268,N_2351);
or U2899 (N_2899,N_2098,N_2171);
nor U2900 (N_2900,N_1632,N_2355);
and U2901 (N_2901,N_1905,N_2376);
and U2902 (N_2902,N_1825,N_2224);
and U2903 (N_2903,N_2113,N_2146);
nor U2904 (N_2904,N_1593,N_1684);
nand U2905 (N_2905,N_1920,N_1442);
nor U2906 (N_2906,N_1317,N_1336);
nor U2907 (N_2907,N_2106,N_1343);
and U2908 (N_2908,N_1490,N_1234);
nand U2909 (N_2909,N_2242,N_2104);
nor U2910 (N_2910,N_2180,N_1476);
nand U2911 (N_2911,N_1844,N_1546);
and U2912 (N_2912,N_1934,N_2278);
xor U2913 (N_2913,N_1298,N_1239);
nor U2914 (N_2914,N_1832,N_2363);
xor U2915 (N_2915,N_1503,N_1709);
nand U2916 (N_2916,N_2388,N_1397);
nor U2917 (N_2917,N_1980,N_1603);
nor U2918 (N_2918,N_1441,N_2260);
or U2919 (N_2919,N_1823,N_1236);
nand U2920 (N_2920,N_1333,N_1988);
xnor U2921 (N_2921,N_1654,N_1722);
nor U2922 (N_2922,N_1556,N_1993);
nor U2923 (N_2923,N_2011,N_1645);
nor U2924 (N_2924,N_1355,N_1377);
nand U2925 (N_2925,N_1720,N_1861);
nor U2926 (N_2926,N_1381,N_2369);
xnor U2927 (N_2927,N_1938,N_1646);
and U2928 (N_2928,N_1842,N_1304);
xor U2929 (N_2929,N_2190,N_2153);
nand U2930 (N_2930,N_1860,N_1849);
xnor U2931 (N_2931,N_1635,N_1657);
or U2932 (N_2932,N_1585,N_2238);
or U2933 (N_2933,N_1398,N_2247);
and U2934 (N_2934,N_2051,N_1235);
or U2935 (N_2935,N_1916,N_1579);
nand U2936 (N_2936,N_1448,N_2289);
and U2937 (N_2937,N_1786,N_1846);
or U2938 (N_2938,N_1631,N_1745);
nand U2939 (N_2939,N_1526,N_1363);
and U2940 (N_2940,N_2162,N_2271);
or U2941 (N_2941,N_2273,N_2138);
nand U2942 (N_2942,N_1850,N_1450);
or U2943 (N_2943,N_2062,N_2123);
or U2944 (N_2944,N_1412,N_1767);
and U2945 (N_2945,N_1729,N_1534);
xnor U2946 (N_2946,N_1723,N_1373);
nor U2947 (N_2947,N_1876,N_1853);
xnor U2948 (N_2948,N_1372,N_1627);
xnor U2949 (N_2949,N_1537,N_1386);
or U2950 (N_2950,N_1542,N_1644);
and U2951 (N_2951,N_1991,N_1337);
nor U2952 (N_2952,N_1843,N_2391);
nand U2953 (N_2953,N_1608,N_2163);
nor U2954 (N_2954,N_1749,N_1756);
or U2955 (N_2955,N_1641,N_1429);
and U2956 (N_2956,N_1663,N_1687);
nor U2957 (N_2957,N_1881,N_1370);
xor U2958 (N_2958,N_2254,N_1708);
nand U2959 (N_2959,N_2174,N_1563);
nand U2960 (N_2960,N_1634,N_1661);
and U2961 (N_2961,N_1638,N_1440);
xnor U2962 (N_2962,N_2323,N_1954);
xnor U2963 (N_2963,N_1713,N_1293);
nor U2964 (N_2964,N_1622,N_1798);
nand U2965 (N_2965,N_1433,N_1711);
and U2966 (N_2966,N_1763,N_2255);
and U2967 (N_2967,N_2178,N_2283);
or U2968 (N_2968,N_1719,N_1257);
or U2969 (N_2969,N_1419,N_2065);
and U2970 (N_2970,N_1772,N_1601);
xor U2971 (N_2971,N_1639,N_2257);
and U2972 (N_2972,N_1570,N_1917);
nor U2973 (N_2973,N_2187,N_1836);
or U2974 (N_2974,N_2225,N_1505);
xnor U2975 (N_2975,N_1500,N_1921);
and U2976 (N_2976,N_1943,N_1899);
nor U2977 (N_2977,N_1830,N_1449);
or U2978 (N_2978,N_1890,N_2080);
or U2979 (N_2979,N_2197,N_1588);
xor U2980 (N_2980,N_1979,N_1455);
xor U2981 (N_2981,N_2140,N_1536);
nor U2982 (N_2982,N_2223,N_1871);
nor U2983 (N_2983,N_1218,N_2017);
or U2984 (N_2984,N_2064,N_2364);
and U2985 (N_2985,N_2304,N_2384);
nand U2986 (N_2986,N_2076,N_1374);
or U2987 (N_2987,N_1584,N_1675);
nor U2988 (N_2988,N_1613,N_1332);
nand U2989 (N_2989,N_1220,N_1902);
and U2990 (N_2990,N_1456,N_1867);
nor U2991 (N_2991,N_2126,N_2226);
nand U2992 (N_2992,N_1498,N_1809);
nand U2993 (N_2993,N_2152,N_2008);
nor U2994 (N_2994,N_1855,N_2191);
and U2995 (N_2995,N_1847,N_1414);
nand U2996 (N_2996,N_1604,N_1391);
or U2997 (N_2997,N_2332,N_1315);
or U2998 (N_2998,N_1643,N_1813);
nand U2999 (N_2999,N_2103,N_1665);
nor U3000 (N_3000,N_1203,N_1653);
or U3001 (N_3001,N_1865,N_1476);
and U3002 (N_3002,N_1771,N_1510);
nand U3003 (N_3003,N_2195,N_1545);
or U3004 (N_3004,N_2129,N_1686);
or U3005 (N_3005,N_1270,N_1468);
nand U3006 (N_3006,N_1590,N_1541);
and U3007 (N_3007,N_1904,N_2089);
nand U3008 (N_3008,N_1937,N_1551);
nand U3009 (N_3009,N_2171,N_1368);
or U3010 (N_3010,N_1546,N_1333);
nor U3011 (N_3011,N_2203,N_1603);
xnor U3012 (N_3012,N_1245,N_1262);
and U3013 (N_3013,N_2205,N_1678);
or U3014 (N_3014,N_1462,N_2097);
xor U3015 (N_3015,N_1667,N_1839);
xor U3016 (N_3016,N_1786,N_2360);
nor U3017 (N_3017,N_1937,N_1851);
xnor U3018 (N_3018,N_1838,N_1430);
nor U3019 (N_3019,N_1372,N_1526);
or U3020 (N_3020,N_1221,N_1516);
xor U3021 (N_3021,N_2380,N_1745);
or U3022 (N_3022,N_1837,N_1429);
xor U3023 (N_3023,N_1914,N_1714);
nor U3024 (N_3024,N_1780,N_1262);
nor U3025 (N_3025,N_1587,N_1847);
nor U3026 (N_3026,N_2368,N_1689);
nand U3027 (N_3027,N_2173,N_2086);
or U3028 (N_3028,N_1949,N_1972);
and U3029 (N_3029,N_2221,N_1315);
nand U3030 (N_3030,N_1571,N_1618);
nand U3031 (N_3031,N_1927,N_1349);
nand U3032 (N_3032,N_1254,N_1974);
and U3033 (N_3033,N_2393,N_1814);
or U3034 (N_3034,N_2382,N_2178);
xor U3035 (N_3035,N_1954,N_2016);
xnor U3036 (N_3036,N_1293,N_2323);
nand U3037 (N_3037,N_1419,N_1905);
xor U3038 (N_3038,N_1648,N_1911);
nand U3039 (N_3039,N_2375,N_1693);
nor U3040 (N_3040,N_1348,N_1489);
or U3041 (N_3041,N_1203,N_2263);
nor U3042 (N_3042,N_1634,N_2238);
xor U3043 (N_3043,N_2302,N_1673);
nand U3044 (N_3044,N_2065,N_1448);
nor U3045 (N_3045,N_1665,N_2276);
and U3046 (N_3046,N_1836,N_1799);
nor U3047 (N_3047,N_1425,N_1230);
or U3048 (N_3048,N_1221,N_1730);
nor U3049 (N_3049,N_1579,N_2198);
nor U3050 (N_3050,N_1223,N_1420);
and U3051 (N_3051,N_1768,N_2253);
xor U3052 (N_3052,N_2037,N_1338);
or U3053 (N_3053,N_2213,N_1738);
nand U3054 (N_3054,N_1926,N_1419);
nor U3055 (N_3055,N_2117,N_2317);
nor U3056 (N_3056,N_2327,N_1742);
xor U3057 (N_3057,N_1842,N_1638);
nand U3058 (N_3058,N_2279,N_1442);
nand U3059 (N_3059,N_1639,N_1987);
or U3060 (N_3060,N_2221,N_1368);
nand U3061 (N_3061,N_1911,N_1281);
xnor U3062 (N_3062,N_1207,N_1234);
xnor U3063 (N_3063,N_1740,N_1579);
xnor U3064 (N_3064,N_2068,N_1756);
and U3065 (N_3065,N_1249,N_1683);
or U3066 (N_3066,N_1514,N_1539);
nor U3067 (N_3067,N_1657,N_1540);
or U3068 (N_3068,N_1378,N_1389);
xnor U3069 (N_3069,N_1940,N_1373);
nor U3070 (N_3070,N_1351,N_1664);
nand U3071 (N_3071,N_1554,N_1789);
nand U3072 (N_3072,N_1714,N_2010);
or U3073 (N_3073,N_1575,N_1204);
xor U3074 (N_3074,N_1313,N_2049);
and U3075 (N_3075,N_1470,N_2273);
xor U3076 (N_3076,N_1502,N_1429);
xnor U3077 (N_3077,N_1271,N_1405);
nor U3078 (N_3078,N_2161,N_1655);
and U3079 (N_3079,N_2101,N_2209);
or U3080 (N_3080,N_2120,N_1568);
nor U3081 (N_3081,N_1931,N_2117);
or U3082 (N_3082,N_1285,N_2048);
nor U3083 (N_3083,N_1547,N_2045);
nand U3084 (N_3084,N_2367,N_1561);
nand U3085 (N_3085,N_2293,N_1952);
and U3086 (N_3086,N_2152,N_2393);
or U3087 (N_3087,N_2162,N_1869);
and U3088 (N_3088,N_2354,N_1328);
xor U3089 (N_3089,N_1680,N_2394);
nand U3090 (N_3090,N_1442,N_1670);
nor U3091 (N_3091,N_1582,N_2255);
xnor U3092 (N_3092,N_1640,N_1246);
or U3093 (N_3093,N_2115,N_2324);
and U3094 (N_3094,N_1453,N_1270);
xor U3095 (N_3095,N_1341,N_2255);
nand U3096 (N_3096,N_1965,N_1499);
nand U3097 (N_3097,N_1473,N_1726);
xnor U3098 (N_3098,N_1741,N_1333);
or U3099 (N_3099,N_2371,N_2139);
and U3100 (N_3100,N_1688,N_1235);
and U3101 (N_3101,N_2206,N_1478);
nand U3102 (N_3102,N_2002,N_2204);
xor U3103 (N_3103,N_2149,N_1381);
xnor U3104 (N_3104,N_1455,N_2210);
nand U3105 (N_3105,N_1926,N_1587);
nor U3106 (N_3106,N_1372,N_1301);
or U3107 (N_3107,N_1360,N_1805);
or U3108 (N_3108,N_1899,N_1333);
or U3109 (N_3109,N_1644,N_2368);
or U3110 (N_3110,N_1266,N_1616);
nor U3111 (N_3111,N_2331,N_1902);
nor U3112 (N_3112,N_1205,N_2053);
nor U3113 (N_3113,N_1482,N_2069);
nand U3114 (N_3114,N_1329,N_1635);
and U3115 (N_3115,N_1409,N_2207);
xor U3116 (N_3116,N_1509,N_2150);
nor U3117 (N_3117,N_1630,N_1671);
or U3118 (N_3118,N_2020,N_1407);
or U3119 (N_3119,N_1889,N_1841);
or U3120 (N_3120,N_1913,N_1986);
and U3121 (N_3121,N_2103,N_1886);
or U3122 (N_3122,N_1641,N_1385);
and U3123 (N_3123,N_1466,N_2384);
nand U3124 (N_3124,N_2390,N_1968);
xnor U3125 (N_3125,N_2213,N_2057);
or U3126 (N_3126,N_1463,N_1782);
nand U3127 (N_3127,N_1648,N_1429);
nand U3128 (N_3128,N_1291,N_2007);
nand U3129 (N_3129,N_1766,N_2082);
or U3130 (N_3130,N_1462,N_1503);
xor U3131 (N_3131,N_1786,N_2193);
nor U3132 (N_3132,N_2023,N_1670);
xor U3133 (N_3133,N_2258,N_1396);
nand U3134 (N_3134,N_1449,N_1698);
nand U3135 (N_3135,N_1537,N_2332);
or U3136 (N_3136,N_1539,N_2380);
xor U3137 (N_3137,N_2318,N_2061);
nor U3138 (N_3138,N_1918,N_1484);
nand U3139 (N_3139,N_1644,N_1405);
and U3140 (N_3140,N_2049,N_1635);
nand U3141 (N_3141,N_1816,N_1579);
or U3142 (N_3142,N_1460,N_1942);
xnor U3143 (N_3143,N_1563,N_1468);
xor U3144 (N_3144,N_1463,N_2169);
nor U3145 (N_3145,N_2365,N_1660);
nor U3146 (N_3146,N_1523,N_1593);
and U3147 (N_3147,N_1350,N_1965);
and U3148 (N_3148,N_1701,N_1285);
nand U3149 (N_3149,N_1675,N_2127);
xnor U3150 (N_3150,N_1986,N_1423);
and U3151 (N_3151,N_1699,N_2369);
nand U3152 (N_3152,N_1462,N_1744);
nor U3153 (N_3153,N_2292,N_2124);
nand U3154 (N_3154,N_1542,N_2344);
or U3155 (N_3155,N_2048,N_1760);
nand U3156 (N_3156,N_1473,N_1559);
xor U3157 (N_3157,N_1823,N_1547);
or U3158 (N_3158,N_1407,N_1761);
nand U3159 (N_3159,N_1791,N_1642);
nor U3160 (N_3160,N_1890,N_1789);
xnor U3161 (N_3161,N_1390,N_1785);
and U3162 (N_3162,N_2364,N_1863);
nand U3163 (N_3163,N_1952,N_1443);
and U3164 (N_3164,N_2057,N_1392);
and U3165 (N_3165,N_1700,N_2239);
nand U3166 (N_3166,N_1839,N_1724);
and U3167 (N_3167,N_2220,N_2246);
xor U3168 (N_3168,N_2240,N_1658);
nor U3169 (N_3169,N_1744,N_2140);
nand U3170 (N_3170,N_1968,N_1316);
nand U3171 (N_3171,N_1763,N_1395);
or U3172 (N_3172,N_1737,N_1374);
nor U3173 (N_3173,N_2157,N_1557);
and U3174 (N_3174,N_1428,N_1982);
nor U3175 (N_3175,N_2185,N_1531);
and U3176 (N_3176,N_1343,N_2375);
xnor U3177 (N_3177,N_2009,N_1312);
nand U3178 (N_3178,N_1718,N_1844);
and U3179 (N_3179,N_2202,N_1407);
or U3180 (N_3180,N_2107,N_2252);
xnor U3181 (N_3181,N_1951,N_1783);
or U3182 (N_3182,N_1804,N_2374);
xnor U3183 (N_3183,N_1383,N_1628);
nor U3184 (N_3184,N_1560,N_2292);
or U3185 (N_3185,N_1798,N_1875);
nand U3186 (N_3186,N_1492,N_1962);
and U3187 (N_3187,N_1734,N_1598);
nand U3188 (N_3188,N_1234,N_1841);
nor U3189 (N_3189,N_1857,N_2055);
nand U3190 (N_3190,N_1310,N_1450);
nand U3191 (N_3191,N_1862,N_2027);
nor U3192 (N_3192,N_1713,N_2293);
and U3193 (N_3193,N_1269,N_1971);
nor U3194 (N_3194,N_1541,N_1237);
nand U3195 (N_3195,N_2147,N_1986);
xnor U3196 (N_3196,N_2247,N_1511);
or U3197 (N_3197,N_1609,N_1889);
nor U3198 (N_3198,N_1302,N_2142);
nor U3199 (N_3199,N_1593,N_2021);
or U3200 (N_3200,N_2032,N_1744);
xnor U3201 (N_3201,N_2008,N_2169);
or U3202 (N_3202,N_1516,N_1259);
or U3203 (N_3203,N_1759,N_1261);
nand U3204 (N_3204,N_2339,N_1591);
or U3205 (N_3205,N_1272,N_1776);
xnor U3206 (N_3206,N_2266,N_2004);
nor U3207 (N_3207,N_2140,N_1257);
nor U3208 (N_3208,N_2204,N_1457);
nand U3209 (N_3209,N_1368,N_1884);
or U3210 (N_3210,N_2227,N_1410);
xor U3211 (N_3211,N_1486,N_2131);
xnor U3212 (N_3212,N_2169,N_1472);
xor U3213 (N_3213,N_2138,N_1249);
and U3214 (N_3214,N_2239,N_1612);
or U3215 (N_3215,N_1848,N_1846);
nor U3216 (N_3216,N_1822,N_2398);
nand U3217 (N_3217,N_2240,N_1660);
nor U3218 (N_3218,N_1648,N_1274);
nand U3219 (N_3219,N_1882,N_1374);
or U3220 (N_3220,N_1941,N_1407);
nor U3221 (N_3221,N_1360,N_2133);
xor U3222 (N_3222,N_2239,N_1883);
or U3223 (N_3223,N_1874,N_1780);
xor U3224 (N_3224,N_1839,N_1494);
nand U3225 (N_3225,N_1659,N_1589);
xor U3226 (N_3226,N_1996,N_1839);
and U3227 (N_3227,N_1395,N_1418);
nand U3228 (N_3228,N_2379,N_1270);
or U3229 (N_3229,N_1780,N_1543);
and U3230 (N_3230,N_1765,N_1676);
or U3231 (N_3231,N_1422,N_2329);
nor U3232 (N_3232,N_1223,N_1957);
nor U3233 (N_3233,N_1631,N_1527);
xor U3234 (N_3234,N_1903,N_1631);
and U3235 (N_3235,N_1919,N_1869);
or U3236 (N_3236,N_1942,N_1909);
and U3237 (N_3237,N_1837,N_2257);
nand U3238 (N_3238,N_1251,N_2267);
and U3239 (N_3239,N_1276,N_1699);
or U3240 (N_3240,N_2342,N_1240);
nand U3241 (N_3241,N_1858,N_1703);
nand U3242 (N_3242,N_1860,N_2348);
xnor U3243 (N_3243,N_2342,N_2261);
or U3244 (N_3244,N_2375,N_1715);
and U3245 (N_3245,N_1967,N_2075);
nand U3246 (N_3246,N_2048,N_1822);
or U3247 (N_3247,N_1384,N_1915);
and U3248 (N_3248,N_1988,N_1804);
and U3249 (N_3249,N_1635,N_1971);
nor U3250 (N_3250,N_2076,N_1826);
and U3251 (N_3251,N_1473,N_1806);
and U3252 (N_3252,N_2218,N_1702);
xor U3253 (N_3253,N_2351,N_1779);
nand U3254 (N_3254,N_1343,N_1283);
xor U3255 (N_3255,N_1371,N_1990);
nor U3256 (N_3256,N_2230,N_2102);
nor U3257 (N_3257,N_2174,N_2160);
nor U3258 (N_3258,N_2104,N_2034);
xor U3259 (N_3259,N_1277,N_1514);
or U3260 (N_3260,N_1351,N_1594);
xor U3261 (N_3261,N_2106,N_2347);
nor U3262 (N_3262,N_1738,N_1357);
and U3263 (N_3263,N_1350,N_2273);
nor U3264 (N_3264,N_1345,N_2202);
nor U3265 (N_3265,N_2336,N_2379);
xor U3266 (N_3266,N_2008,N_1949);
or U3267 (N_3267,N_2218,N_1250);
and U3268 (N_3268,N_1514,N_1210);
or U3269 (N_3269,N_2097,N_2398);
and U3270 (N_3270,N_2119,N_2336);
or U3271 (N_3271,N_1842,N_1578);
nand U3272 (N_3272,N_1947,N_1750);
nor U3273 (N_3273,N_2046,N_1449);
xor U3274 (N_3274,N_1260,N_2351);
and U3275 (N_3275,N_2367,N_2286);
xor U3276 (N_3276,N_1920,N_2149);
and U3277 (N_3277,N_2361,N_1448);
xnor U3278 (N_3278,N_1556,N_2088);
and U3279 (N_3279,N_1858,N_2064);
nand U3280 (N_3280,N_1253,N_2355);
xor U3281 (N_3281,N_2157,N_1527);
or U3282 (N_3282,N_1911,N_1407);
nand U3283 (N_3283,N_2085,N_2105);
and U3284 (N_3284,N_2219,N_1765);
nor U3285 (N_3285,N_2238,N_1225);
or U3286 (N_3286,N_1520,N_2002);
nor U3287 (N_3287,N_1464,N_1552);
xor U3288 (N_3288,N_1775,N_1809);
xnor U3289 (N_3289,N_1488,N_1866);
xnor U3290 (N_3290,N_2073,N_1844);
nor U3291 (N_3291,N_1361,N_1381);
nand U3292 (N_3292,N_1911,N_2066);
or U3293 (N_3293,N_2326,N_1833);
xnor U3294 (N_3294,N_2227,N_1541);
xor U3295 (N_3295,N_1476,N_1665);
and U3296 (N_3296,N_1866,N_1967);
or U3297 (N_3297,N_2376,N_2086);
nor U3298 (N_3298,N_2202,N_2359);
xnor U3299 (N_3299,N_2113,N_2212);
or U3300 (N_3300,N_2116,N_2276);
xnor U3301 (N_3301,N_2132,N_1609);
and U3302 (N_3302,N_1688,N_1494);
or U3303 (N_3303,N_1889,N_1276);
xnor U3304 (N_3304,N_2307,N_1327);
or U3305 (N_3305,N_1434,N_1321);
nand U3306 (N_3306,N_1976,N_1554);
xnor U3307 (N_3307,N_2160,N_2080);
nand U3308 (N_3308,N_1411,N_1822);
nand U3309 (N_3309,N_1985,N_1773);
or U3310 (N_3310,N_1206,N_1564);
xnor U3311 (N_3311,N_1362,N_1847);
and U3312 (N_3312,N_1266,N_1820);
xnor U3313 (N_3313,N_1244,N_1364);
nand U3314 (N_3314,N_2258,N_1788);
nor U3315 (N_3315,N_1983,N_1666);
and U3316 (N_3316,N_1669,N_1889);
nand U3317 (N_3317,N_2343,N_1340);
nand U3318 (N_3318,N_2278,N_1834);
nand U3319 (N_3319,N_1327,N_1547);
and U3320 (N_3320,N_1635,N_1560);
nor U3321 (N_3321,N_1953,N_1619);
or U3322 (N_3322,N_2190,N_1719);
and U3323 (N_3323,N_1539,N_2089);
and U3324 (N_3324,N_1589,N_1852);
nand U3325 (N_3325,N_1632,N_1656);
nand U3326 (N_3326,N_1648,N_2207);
nand U3327 (N_3327,N_1969,N_1920);
or U3328 (N_3328,N_2076,N_1387);
nor U3329 (N_3329,N_2367,N_2392);
nand U3330 (N_3330,N_1508,N_1645);
nor U3331 (N_3331,N_1880,N_1485);
nor U3332 (N_3332,N_1939,N_1391);
and U3333 (N_3333,N_1924,N_1202);
nand U3334 (N_3334,N_2140,N_1957);
xnor U3335 (N_3335,N_1560,N_1882);
or U3336 (N_3336,N_1814,N_2306);
xor U3337 (N_3337,N_1613,N_1965);
nor U3338 (N_3338,N_1877,N_2323);
or U3339 (N_3339,N_2074,N_1798);
nand U3340 (N_3340,N_1784,N_1908);
and U3341 (N_3341,N_1865,N_1419);
nor U3342 (N_3342,N_1583,N_2186);
nor U3343 (N_3343,N_2133,N_1213);
nand U3344 (N_3344,N_1724,N_1817);
or U3345 (N_3345,N_1580,N_1747);
nand U3346 (N_3346,N_2043,N_2314);
and U3347 (N_3347,N_2062,N_2047);
or U3348 (N_3348,N_1467,N_2238);
nand U3349 (N_3349,N_1284,N_1521);
and U3350 (N_3350,N_1519,N_1851);
or U3351 (N_3351,N_2162,N_1434);
xor U3352 (N_3352,N_2270,N_1787);
nor U3353 (N_3353,N_1767,N_1690);
and U3354 (N_3354,N_1415,N_1413);
nor U3355 (N_3355,N_1670,N_1977);
xnor U3356 (N_3356,N_1526,N_1575);
nand U3357 (N_3357,N_1259,N_1750);
and U3358 (N_3358,N_2241,N_1798);
nor U3359 (N_3359,N_1387,N_2191);
xnor U3360 (N_3360,N_1223,N_2024);
or U3361 (N_3361,N_1940,N_2156);
nor U3362 (N_3362,N_2290,N_1555);
xor U3363 (N_3363,N_1354,N_1932);
and U3364 (N_3364,N_1761,N_2060);
xor U3365 (N_3365,N_1436,N_2083);
nand U3366 (N_3366,N_1446,N_1213);
xnor U3367 (N_3367,N_2355,N_2131);
nor U3368 (N_3368,N_2292,N_1283);
or U3369 (N_3369,N_1650,N_2250);
and U3370 (N_3370,N_1623,N_2005);
nor U3371 (N_3371,N_1651,N_2086);
or U3372 (N_3372,N_2380,N_1678);
xor U3373 (N_3373,N_1683,N_2138);
and U3374 (N_3374,N_1569,N_1435);
nand U3375 (N_3375,N_1746,N_1774);
and U3376 (N_3376,N_2301,N_2292);
nor U3377 (N_3377,N_1244,N_2361);
nand U3378 (N_3378,N_1244,N_1752);
nor U3379 (N_3379,N_1969,N_1762);
or U3380 (N_3380,N_2259,N_1922);
nand U3381 (N_3381,N_1772,N_1864);
or U3382 (N_3382,N_1976,N_1278);
xor U3383 (N_3383,N_2374,N_1505);
nand U3384 (N_3384,N_1465,N_2004);
xor U3385 (N_3385,N_1451,N_1635);
nand U3386 (N_3386,N_1399,N_1551);
xnor U3387 (N_3387,N_1655,N_1360);
xor U3388 (N_3388,N_1586,N_1902);
or U3389 (N_3389,N_1766,N_2056);
nor U3390 (N_3390,N_1633,N_1805);
and U3391 (N_3391,N_1287,N_1350);
nand U3392 (N_3392,N_1424,N_1233);
nand U3393 (N_3393,N_2187,N_2034);
nand U3394 (N_3394,N_1819,N_1492);
nand U3395 (N_3395,N_1238,N_1413);
and U3396 (N_3396,N_2133,N_1290);
or U3397 (N_3397,N_1585,N_1716);
or U3398 (N_3398,N_1732,N_1306);
and U3399 (N_3399,N_1422,N_1796);
xnor U3400 (N_3400,N_2028,N_1739);
and U3401 (N_3401,N_1367,N_1541);
nor U3402 (N_3402,N_2127,N_1728);
xnor U3403 (N_3403,N_1756,N_1315);
or U3404 (N_3404,N_1817,N_1842);
xnor U3405 (N_3405,N_2134,N_1799);
nand U3406 (N_3406,N_2201,N_1783);
or U3407 (N_3407,N_1461,N_2316);
nor U3408 (N_3408,N_2377,N_1605);
and U3409 (N_3409,N_1459,N_1765);
nor U3410 (N_3410,N_2278,N_1781);
or U3411 (N_3411,N_1208,N_1666);
and U3412 (N_3412,N_1555,N_1634);
nand U3413 (N_3413,N_1985,N_1574);
and U3414 (N_3414,N_2295,N_1532);
xor U3415 (N_3415,N_1326,N_1889);
xnor U3416 (N_3416,N_2330,N_1291);
xor U3417 (N_3417,N_1675,N_1301);
nand U3418 (N_3418,N_2167,N_2015);
nand U3419 (N_3419,N_1342,N_1716);
xor U3420 (N_3420,N_1286,N_2300);
nand U3421 (N_3421,N_1618,N_1651);
nand U3422 (N_3422,N_1571,N_1790);
nor U3423 (N_3423,N_1204,N_1647);
or U3424 (N_3424,N_1797,N_2019);
and U3425 (N_3425,N_1773,N_2224);
or U3426 (N_3426,N_1729,N_1517);
xnor U3427 (N_3427,N_2241,N_2395);
and U3428 (N_3428,N_1880,N_2058);
or U3429 (N_3429,N_1581,N_1429);
nor U3430 (N_3430,N_1555,N_2229);
or U3431 (N_3431,N_2057,N_2193);
nand U3432 (N_3432,N_2289,N_1871);
and U3433 (N_3433,N_2250,N_1510);
and U3434 (N_3434,N_1249,N_1606);
and U3435 (N_3435,N_1533,N_2079);
nor U3436 (N_3436,N_1571,N_2120);
xor U3437 (N_3437,N_1368,N_1598);
nand U3438 (N_3438,N_1466,N_1491);
and U3439 (N_3439,N_1807,N_1455);
nor U3440 (N_3440,N_2201,N_1578);
nor U3441 (N_3441,N_1557,N_1865);
and U3442 (N_3442,N_2343,N_1578);
nand U3443 (N_3443,N_1410,N_1313);
nor U3444 (N_3444,N_1875,N_1770);
xnor U3445 (N_3445,N_1806,N_1784);
xor U3446 (N_3446,N_1496,N_1904);
nand U3447 (N_3447,N_1489,N_2332);
and U3448 (N_3448,N_1675,N_1795);
nand U3449 (N_3449,N_1307,N_1644);
xor U3450 (N_3450,N_1893,N_2328);
and U3451 (N_3451,N_1882,N_2338);
or U3452 (N_3452,N_2183,N_1534);
xor U3453 (N_3453,N_1773,N_1651);
nor U3454 (N_3454,N_1446,N_1657);
or U3455 (N_3455,N_2154,N_1339);
nand U3456 (N_3456,N_2309,N_1835);
and U3457 (N_3457,N_1800,N_2211);
xor U3458 (N_3458,N_1494,N_1265);
nor U3459 (N_3459,N_1509,N_1557);
and U3460 (N_3460,N_1844,N_2288);
nor U3461 (N_3461,N_1943,N_2336);
and U3462 (N_3462,N_1705,N_1713);
and U3463 (N_3463,N_2368,N_1327);
nor U3464 (N_3464,N_2205,N_1282);
nor U3465 (N_3465,N_2001,N_2343);
nor U3466 (N_3466,N_2175,N_1487);
xnor U3467 (N_3467,N_2281,N_2395);
nand U3468 (N_3468,N_2297,N_2394);
nand U3469 (N_3469,N_1400,N_2227);
and U3470 (N_3470,N_2140,N_1616);
nor U3471 (N_3471,N_2266,N_2283);
or U3472 (N_3472,N_1382,N_1641);
nand U3473 (N_3473,N_1523,N_1915);
xnor U3474 (N_3474,N_1900,N_1706);
or U3475 (N_3475,N_1809,N_1474);
and U3476 (N_3476,N_2267,N_1238);
or U3477 (N_3477,N_1686,N_1222);
and U3478 (N_3478,N_1761,N_1614);
nand U3479 (N_3479,N_2078,N_1870);
and U3480 (N_3480,N_1623,N_1703);
or U3481 (N_3481,N_1353,N_1291);
xnor U3482 (N_3482,N_1383,N_1519);
or U3483 (N_3483,N_1849,N_1616);
nor U3484 (N_3484,N_1642,N_1647);
nor U3485 (N_3485,N_1757,N_1946);
and U3486 (N_3486,N_1861,N_2234);
nor U3487 (N_3487,N_1390,N_2204);
and U3488 (N_3488,N_1498,N_2088);
xnor U3489 (N_3489,N_2032,N_1970);
and U3490 (N_3490,N_2284,N_1662);
nand U3491 (N_3491,N_1685,N_1786);
nor U3492 (N_3492,N_2225,N_2031);
nand U3493 (N_3493,N_1643,N_2012);
and U3494 (N_3494,N_1299,N_1975);
nand U3495 (N_3495,N_2125,N_2153);
and U3496 (N_3496,N_1235,N_2209);
xor U3497 (N_3497,N_1468,N_2092);
xnor U3498 (N_3498,N_1238,N_1370);
nor U3499 (N_3499,N_1901,N_1731);
and U3500 (N_3500,N_2382,N_1210);
xor U3501 (N_3501,N_1406,N_2117);
nor U3502 (N_3502,N_1595,N_1561);
nand U3503 (N_3503,N_1531,N_2110);
or U3504 (N_3504,N_2140,N_1255);
and U3505 (N_3505,N_1349,N_2094);
nor U3506 (N_3506,N_1222,N_2048);
nand U3507 (N_3507,N_2224,N_2235);
nor U3508 (N_3508,N_2331,N_2390);
nand U3509 (N_3509,N_1332,N_1818);
nand U3510 (N_3510,N_1868,N_1496);
and U3511 (N_3511,N_2221,N_1422);
or U3512 (N_3512,N_2114,N_2293);
xnor U3513 (N_3513,N_2307,N_1994);
xor U3514 (N_3514,N_1639,N_1463);
or U3515 (N_3515,N_1850,N_1897);
or U3516 (N_3516,N_1672,N_2062);
and U3517 (N_3517,N_1706,N_1566);
or U3518 (N_3518,N_2184,N_1558);
xor U3519 (N_3519,N_1251,N_1269);
or U3520 (N_3520,N_1305,N_2175);
and U3521 (N_3521,N_1769,N_1246);
nor U3522 (N_3522,N_2057,N_1668);
xor U3523 (N_3523,N_1621,N_2174);
nand U3524 (N_3524,N_1353,N_1417);
nand U3525 (N_3525,N_1955,N_2098);
nor U3526 (N_3526,N_1733,N_1777);
xnor U3527 (N_3527,N_1674,N_2164);
and U3528 (N_3528,N_1600,N_2021);
nor U3529 (N_3529,N_2351,N_1917);
nand U3530 (N_3530,N_1677,N_2130);
nor U3531 (N_3531,N_1701,N_2137);
nor U3532 (N_3532,N_1868,N_2062);
or U3533 (N_3533,N_2069,N_2228);
and U3534 (N_3534,N_1507,N_1834);
and U3535 (N_3535,N_1778,N_2107);
nand U3536 (N_3536,N_1575,N_1555);
nand U3537 (N_3537,N_2204,N_1472);
and U3538 (N_3538,N_1967,N_2158);
nor U3539 (N_3539,N_1299,N_2046);
nor U3540 (N_3540,N_2068,N_2273);
nand U3541 (N_3541,N_1475,N_2175);
nor U3542 (N_3542,N_2189,N_1779);
nand U3543 (N_3543,N_1587,N_1207);
and U3544 (N_3544,N_1337,N_1387);
or U3545 (N_3545,N_1346,N_1738);
xor U3546 (N_3546,N_2161,N_1279);
nand U3547 (N_3547,N_2033,N_1720);
or U3548 (N_3548,N_1838,N_1954);
nor U3549 (N_3549,N_1559,N_1952);
nor U3550 (N_3550,N_1983,N_2103);
or U3551 (N_3551,N_2058,N_2316);
and U3552 (N_3552,N_1711,N_1801);
nor U3553 (N_3553,N_1547,N_2238);
and U3554 (N_3554,N_2018,N_1976);
xor U3555 (N_3555,N_1691,N_2205);
nand U3556 (N_3556,N_1321,N_2252);
nor U3557 (N_3557,N_1270,N_1705);
nor U3558 (N_3558,N_1420,N_1303);
and U3559 (N_3559,N_1601,N_1752);
or U3560 (N_3560,N_2185,N_1527);
nand U3561 (N_3561,N_1864,N_1820);
or U3562 (N_3562,N_2176,N_2201);
or U3563 (N_3563,N_2224,N_2230);
nor U3564 (N_3564,N_1776,N_1200);
and U3565 (N_3565,N_1949,N_1303);
or U3566 (N_3566,N_1654,N_1239);
or U3567 (N_3567,N_1953,N_1529);
xnor U3568 (N_3568,N_1491,N_2161);
nor U3569 (N_3569,N_1930,N_1678);
or U3570 (N_3570,N_1516,N_1457);
nand U3571 (N_3571,N_1454,N_2137);
nand U3572 (N_3572,N_2177,N_2368);
nor U3573 (N_3573,N_1878,N_1278);
and U3574 (N_3574,N_1523,N_1618);
and U3575 (N_3575,N_1518,N_1514);
nand U3576 (N_3576,N_1701,N_1245);
nand U3577 (N_3577,N_2361,N_1295);
and U3578 (N_3578,N_1250,N_1873);
or U3579 (N_3579,N_2103,N_1711);
nand U3580 (N_3580,N_2103,N_1637);
nand U3581 (N_3581,N_2384,N_2282);
nor U3582 (N_3582,N_1929,N_1345);
xor U3583 (N_3583,N_2036,N_1216);
or U3584 (N_3584,N_1961,N_1951);
xnor U3585 (N_3585,N_2344,N_1358);
nand U3586 (N_3586,N_1828,N_1866);
xor U3587 (N_3587,N_1990,N_1619);
xnor U3588 (N_3588,N_2107,N_2185);
nand U3589 (N_3589,N_1257,N_1640);
or U3590 (N_3590,N_1949,N_2264);
or U3591 (N_3591,N_1562,N_2379);
nor U3592 (N_3592,N_2182,N_2041);
nand U3593 (N_3593,N_1718,N_2038);
and U3594 (N_3594,N_2022,N_1594);
xor U3595 (N_3595,N_1862,N_2024);
or U3596 (N_3596,N_1851,N_1473);
and U3597 (N_3597,N_1541,N_2356);
xor U3598 (N_3598,N_1366,N_1480);
xor U3599 (N_3599,N_1740,N_1355);
nand U3600 (N_3600,N_3014,N_2784);
xor U3601 (N_3601,N_3324,N_2610);
and U3602 (N_3602,N_3454,N_2446);
xnor U3603 (N_3603,N_3372,N_3436);
nor U3604 (N_3604,N_2663,N_3159);
or U3605 (N_3605,N_2647,N_3556);
nor U3606 (N_3606,N_2580,N_3345);
xor U3607 (N_3607,N_3318,N_2637);
or U3608 (N_3608,N_2703,N_2570);
or U3609 (N_3609,N_2559,N_3511);
nand U3610 (N_3610,N_2970,N_2615);
xor U3611 (N_3611,N_2917,N_2674);
nor U3612 (N_3612,N_3252,N_2984);
nor U3613 (N_3613,N_2470,N_2788);
nor U3614 (N_3614,N_3148,N_3138);
and U3615 (N_3615,N_2937,N_3288);
nand U3616 (N_3616,N_2652,N_2881);
xor U3617 (N_3617,N_3027,N_2489);
xor U3618 (N_3618,N_3041,N_3243);
and U3619 (N_3619,N_3172,N_3430);
nand U3620 (N_3620,N_3572,N_3522);
xnor U3621 (N_3621,N_2665,N_3595);
and U3622 (N_3622,N_2825,N_3245);
xnor U3623 (N_3623,N_2473,N_2497);
and U3624 (N_3624,N_2946,N_2588);
xnor U3625 (N_3625,N_3200,N_3329);
nor U3626 (N_3626,N_3587,N_3507);
nand U3627 (N_3627,N_2648,N_2622);
nor U3628 (N_3628,N_3249,N_2577);
or U3629 (N_3629,N_3122,N_3232);
and U3630 (N_3630,N_3520,N_3567);
nor U3631 (N_3631,N_2625,N_2947);
and U3632 (N_3632,N_3256,N_2523);
or U3633 (N_3633,N_3362,N_2491);
or U3634 (N_3634,N_2675,N_3540);
xnor U3635 (N_3635,N_2505,N_3559);
nor U3636 (N_3636,N_3361,N_3493);
nand U3637 (N_3637,N_3353,N_2716);
nand U3638 (N_3638,N_3450,N_3498);
or U3639 (N_3639,N_3301,N_2530);
nand U3640 (N_3640,N_2520,N_3218);
xnor U3641 (N_3641,N_2488,N_2850);
nor U3642 (N_3642,N_3577,N_2687);
and U3643 (N_3643,N_3016,N_3055);
nor U3644 (N_3644,N_2453,N_2644);
nand U3645 (N_3645,N_2441,N_2713);
nor U3646 (N_3646,N_2790,N_2954);
nor U3647 (N_3647,N_2636,N_3585);
xor U3648 (N_3648,N_2434,N_3512);
xnor U3649 (N_3649,N_2705,N_2902);
nand U3650 (N_3650,N_2410,N_2775);
or U3651 (N_3651,N_2933,N_3561);
nand U3652 (N_3652,N_2742,N_2465);
nand U3653 (N_3653,N_2961,N_3352);
or U3654 (N_3654,N_3338,N_2678);
and U3655 (N_3655,N_3149,N_3410);
nand U3656 (N_3656,N_2493,N_2681);
nand U3657 (N_3657,N_3461,N_3371);
nor U3658 (N_3658,N_3581,N_3596);
nand U3659 (N_3659,N_2621,N_3568);
or U3660 (N_3660,N_3356,N_2824);
nor U3661 (N_3661,N_2847,N_2859);
or U3662 (N_3662,N_2765,N_3081);
xor U3663 (N_3663,N_3107,N_2720);
xor U3664 (N_3664,N_2511,N_2481);
or U3665 (N_3665,N_2799,N_3445);
and U3666 (N_3666,N_2758,N_3396);
or U3667 (N_3667,N_3384,N_3059);
or U3668 (N_3668,N_3150,N_3173);
nand U3669 (N_3669,N_2971,N_2948);
nand U3670 (N_3670,N_2899,N_2557);
nor U3671 (N_3671,N_2731,N_2952);
nor U3672 (N_3672,N_2585,N_2736);
xor U3673 (N_3673,N_2506,N_3255);
xor U3674 (N_3674,N_3291,N_3294);
nor U3675 (N_3675,N_2502,N_2684);
nor U3676 (N_3676,N_2438,N_3437);
nor U3677 (N_3677,N_2592,N_2867);
xnor U3678 (N_3678,N_2963,N_2760);
and U3679 (N_3679,N_3012,N_3504);
xor U3680 (N_3680,N_2762,N_2564);
and U3681 (N_3681,N_2873,N_2466);
and U3682 (N_3682,N_3115,N_2806);
xnor U3683 (N_3683,N_2459,N_2938);
xor U3684 (N_3684,N_2476,N_3278);
and U3685 (N_3685,N_3474,N_2912);
nand U3686 (N_3686,N_3388,N_3290);
nand U3687 (N_3687,N_3598,N_2953);
nand U3688 (N_3688,N_2818,N_2500);
nand U3689 (N_3689,N_2890,N_2604);
xor U3690 (N_3690,N_3141,N_2794);
nor U3691 (N_3691,N_3413,N_2729);
or U3692 (N_3692,N_2608,N_3316);
or U3693 (N_3693,N_2853,N_2940);
xor U3694 (N_3694,N_3536,N_2628);
nor U3695 (N_3695,N_2981,N_2693);
xnor U3696 (N_3696,N_2649,N_2682);
or U3697 (N_3697,N_3344,N_3404);
or U3698 (N_3698,N_2650,N_3216);
nor U3699 (N_3699,N_2416,N_2694);
nand U3700 (N_3700,N_2802,N_3281);
xor U3701 (N_3701,N_2719,N_2659);
nor U3702 (N_3702,N_3578,N_2602);
nand U3703 (N_3703,N_3346,N_3307);
and U3704 (N_3704,N_2535,N_3331);
nor U3705 (N_3705,N_3298,N_2992);
xnor U3706 (N_3706,N_3054,N_3189);
xor U3707 (N_3707,N_3032,N_3201);
xor U3708 (N_3708,N_3087,N_3002);
and U3709 (N_3709,N_2436,N_2852);
or U3710 (N_3710,N_2748,N_2668);
nand U3711 (N_3711,N_2797,N_3072);
and U3712 (N_3712,N_3280,N_2885);
or U3713 (N_3713,N_3276,N_3000);
nor U3714 (N_3714,N_2586,N_3181);
nor U3715 (N_3715,N_3078,N_3211);
or U3716 (N_3716,N_2814,N_3408);
nor U3717 (N_3717,N_2988,N_3406);
nand U3718 (N_3718,N_2638,N_2642);
or U3719 (N_3719,N_2995,N_2712);
and U3720 (N_3720,N_2914,N_2891);
nand U3721 (N_3721,N_3576,N_2974);
and U3722 (N_3722,N_2425,N_3239);
or U3723 (N_3723,N_2986,N_3038);
or U3724 (N_3724,N_2728,N_3099);
or U3725 (N_3725,N_3530,N_2996);
xor U3726 (N_3726,N_2723,N_2629);
or U3727 (N_3727,N_3472,N_3357);
nand U3728 (N_3728,N_3349,N_3185);
xnor U3729 (N_3729,N_3351,N_3386);
and U3730 (N_3730,N_3541,N_3348);
or U3731 (N_3731,N_2490,N_3036);
or U3732 (N_3732,N_2851,N_3263);
nor U3733 (N_3733,N_2420,N_2838);
or U3734 (N_3734,N_2471,N_2671);
or U3735 (N_3735,N_3193,N_2451);
xor U3736 (N_3736,N_3224,N_2896);
nor U3737 (N_3737,N_3492,N_2931);
and U3738 (N_3738,N_2534,N_3594);
or U3739 (N_3739,N_3420,N_3519);
xor U3740 (N_3740,N_2627,N_2739);
and U3741 (N_3741,N_3171,N_3202);
nor U3742 (N_3742,N_2479,N_3476);
and U3743 (N_3743,N_2526,N_3487);
nor U3744 (N_3744,N_3505,N_3451);
or U3745 (N_3745,N_3253,N_2759);
or U3746 (N_3746,N_2879,N_3550);
or U3747 (N_3747,N_3187,N_3254);
nand U3748 (N_3748,N_2764,N_3111);
or U3749 (N_3749,N_3135,N_2524);
xnor U3750 (N_3750,N_2672,N_2596);
and U3751 (N_3751,N_2576,N_2777);
nand U3752 (N_3752,N_2973,N_2443);
or U3753 (N_3753,N_3025,N_2866);
or U3754 (N_3754,N_3154,N_2882);
xor U3755 (N_3755,N_2406,N_3031);
xnor U3756 (N_3756,N_2911,N_3593);
nor U3757 (N_3757,N_2903,N_3240);
or U3758 (N_3758,N_2613,N_3570);
or U3759 (N_3759,N_3395,N_2486);
nor U3760 (N_3760,N_3162,N_3580);
nand U3761 (N_3761,N_3447,N_3573);
xnor U3762 (N_3762,N_3340,N_2427);
xnor U3763 (N_3763,N_3066,N_3082);
nand U3764 (N_3764,N_2755,N_3365);
or U3765 (N_3765,N_3260,N_3106);
and U3766 (N_3766,N_2733,N_3019);
or U3767 (N_3767,N_3426,N_3199);
or U3768 (N_3768,N_2454,N_2780);
nand U3769 (N_3769,N_3063,N_2558);
and U3770 (N_3770,N_3177,N_3155);
and U3771 (N_3771,N_3328,N_3207);
and U3772 (N_3772,N_3175,N_2413);
nor U3773 (N_3773,N_3157,N_2856);
nor U3774 (N_3774,N_3167,N_2985);
nor U3775 (N_3775,N_3174,N_3514);
nor U3776 (N_3776,N_3494,N_3070);
and U3777 (N_3777,N_3442,N_2993);
and U3778 (N_3778,N_3553,N_2521);
xnor U3779 (N_3779,N_2964,N_3277);
nand U3780 (N_3780,N_2670,N_3179);
or U3781 (N_3781,N_3557,N_2785);
or U3782 (N_3782,N_3247,N_2673);
xnor U3783 (N_3783,N_2793,N_2783);
xnor U3784 (N_3784,N_2766,N_2792);
and U3785 (N_3785,N_3008,N_2480);
and U3786 (N_3786,N_2706,N_3315);
and U3787 (N_3787,N_3131,N_2710);
and U3788 (N_3788,N_3168,N_2848);
nand U3789 (N_3789,N_3283,N_3385);
nor U3790 (N_3790,N_2540,N_3412);
and U3791 (N_3791,N_3160,N_3104);
or U3792 (N_3792,N_2464,N_3035);
and U3793 (N_3793,N_2907,N_2469);
nor U3794 (N_3794,N_3496,N_2715);
nand U3795 (N_3795,N_2424,N_3061);
xor U3796 (N_3796,N_2855,N_2400);
xnor U3797 (N_3797,N_3421,N_3533);
or U3798 (N_3798,N_2640,N_2515);
xor U3799 (N_3799,N_3342,N_2707);
and U3800 (N_3800,N_3021,N_3432);
or U3801 (N_3801,N_3416,N_2979);
nor U3802 (N_3802,N_2639,N_2876);
and U3803 (N_3803,N_2661,N_2959);
xor U3804 (N_3804,N_3210,N_3304);
and U3805 (N_3805,N_2417,N_3562);
and U3806 (N_3806,N_3490,N_2485);
and U3807 (N_3807,N_3275,N_3102);
nand U3808 (N_3808,N_3369,N_2768);
or U3809 (N_3809,N_3323,N_3013);
or U3810 (N_3810,N_3268,N_2495);
xor U3811 (N_3811,N_2928,N_3480);
and U3812 (N_3812,N_2732,N_2776);
xor U3813 (N_3813,N_2655,N_2677);
nand U3814 (N_3814,N_3523,N_3435);
or U3815 (N_3815,N_2428,N_3332);
nor U3816 (N_3816,N_3428,N_2704);
xnor U3817 (N_3817,N_3214,N_3591);
xnor U3818 (N_3818,N_3129,N_2698);
xor U3819 (N_3819,N_3484,N_3321);
nor U3820 (N_3820,N_2738,N_3105);
nor U3821 (N_3821,N_3191,N_3552);
or U3822 (N_3822,N_2810,N_2967);
nand U3823 (N_3823,N_2965,N_3588);
and U3824 (N_3824,N_3402,N_2927);
and U3825 (N_3825,N_3560,N_2617);
nand U3826 (N_3826,N_3192,N_3397);
nor U3827 (N_3827,N_3479,N_3023);
or U3828 (N_3828,N_3212,N_3103);
or U3829 (N_3829,N_3271,N_2426);
or U3830 (N_3830,N_3320,N_2412);
or U3831 (N_3831,N_3441,N_3548);
or U3832 (N_3832,N_3250,N_3544);
nor U3833 (N_3833,N_3265,N_2932);
nand U3834 (N_3834,N_2421,N_2737);
nor U3835 (N_3835,N_2916,N_3225);
and U3836 (N_3836,N_3266,N_2843);
or U3837 (N_3837,N_3091,N_2997);
nor U3838 (N_3838,N_3554,N_2669);
and U3839 (N_3839,N_3438,N_3090);
nand U3840 (N_3840,N_2895,N_2624);
nor U3841 (N_3841,N_3095,N_3382);
nand U3842 (N_3842,N_3322,N_2800);
and U3843 (N_3843,N_3183,N_2711);
xnor U3844 (N_3844,N_2977,N_2607);
nor U3845 (N_3845,N_3546,N_2442);
or U3846 (N_3846,N_3046,N_2423);
or U3847 (N_3847,N_2846,N_2975);
nand U3848 (N_3848,N_2960,N_2508);
or U3849 (N_3849,N_2990,N_3146);
xor U3850 (N_3850,N_3444,N_2578);
xor U3851 (N_3851,N_2600,N_3236);
nor U3852 (N_3852,N_3267,N_2878);
nor U3853 (N_3853,N_2498,N_3020);
xor U3854 (N_3854,N_2612,N_3333);
or U3855 (N_3855,N_3161,N_3488);
nor U3856 (N_3856,N_3040,N_3228);
nand U3857 (N_3857,N_2407,N_2516);
and U3858 (N_3858,N_3312,N_3350);
nand U3859 (N_3859,N_3467,N_2791);
xor U3860 (N_3860,N_2877,N_2849);
or U3861 (N_3861,N_2823,N_2708);
or U3862 (N_3862,N_2982,N_2543);
nor U3863 (N_3863,N_3062,N_2718);
and U3864 (N_3864,N_3469,N_3394);
and U3865 (N_3865,N_3478,N_2656);
or U3866 (N_3866,N_3547,N_2864);
or U3867 (N_3867,N_3528,N_2531);
and U3868 (N_3868,N_3269,N_3376);
nand U3869 (N_3869,N_3094,N_2819);
nand U3870 (N_3870,N_3389,N_2680);
or U3871 (N_3871,N_3354,N_2808);
nor U3872 (N_3872,N_3489,N_2956);
or U3873 (N_3873,N_3116,N_3153);
and U3874 (N_3874,N_2512,N_2821);
xor U3875 (N_3875,N_3071,N_3303);
nand U3876 (N_3876,N_2835,N_2841);
nand U3877 (N_3877,N_3525,N_2957);
nand U3878 (N_3878,N_2528,N_3423);
and U3879 (N_3879,N_2976,N_2870);
and U3880 (N_3880,N_3089,N_3110);
nand U3881 (N_3881,N_2654,N_2437);
nor U3882 (N_3882,N_2595,N_2830);
nand U3883 (N_3883,N_2462,N_2880);
and U3884 (N_3884,N_2779,N_3213);
nor U3885 (N_3885,N_2583,N_2468);
and U3886 (N_3886,N_2483,N_3198);
xnor U3887 (N_3887,N_3571,N_3400);
nand U3888 (N_3888,N_2561,N_2422);
xor U3889 (N_3889,N_2450,N_2894);
or U3890 (N_3890,N_3176,N_3539);
or U3891 (N_3891,N_2549,N_2641);
nand U3892 (N_3892,N_2845,N_3123);
and U3893 (N_3893,N_3024,N_2653);
nor U3894 (N_3894,N_3196,N_2862);
nand U3895 (N_3895,N_2721,N_2919);
or U3896 (N_3896,N_2941,N_2539);
nor U3897 (N_3897,N_3076,N_3433);
nor U3898 (N_3898,N_2532,N_3381);
nand U3899 (N_3899,N_3093,N_2522);
and U3900 (N_3900,N_3453,N_2909);
nand U3901 (N_3901,N_3206,N_3403);
or U3902 (N_3902,N_3001,N_2966);
xor U3903 (N_3903,N_3030,N_2789);
or U3904 (N_3904,N_2701,N_3182);
or U3905 (N_3905,N_3518,N_3419);
nand U3906 (N_3906,N_2743,N_2717);
or U3907 (N_3907,N_3347,N_3314);
or U3908 (N_3908,N_3446,N_3424);
xnor U3909 (N_3909,N_2751,N_2457);
and U3910 (N_3910,N_2913,N_3050);
or U3911 (N_3911,N_2553,N_2805);
xor U3912 (N_3912,N_3513,N_2472);
xnor U3913 (N_3913,N_2439,N_2685);
and U3914 (N_3914,N_3343,N_3590);
xor U3915 (N_3915,N_3434,N_3471);
xor U3916 (N_3916,N_3380,N_3537);
nor U3917 (N_3917,N_3109,N_3085);
and U3918 (N_3918,N_3440,N_2552);
nor U3919 (N_3919,N_2904,N_2513);
nand U3920 (N_3920,N_3586,N_3056);
nand U3921 (N_3921,N_3482,N_3052);
nor U3922 (N_3922,N_2690,N_3235);
or U3923 (N_3923,N_2501,N_2906);
xor U3924 (N_3924,N_3248,N_3169);
and U3925 (N_3925,N_3259,N_3355);
and U3926 (N_3926,N_3118,N_3405);
or U3927 (N_3927,N_3462,N_2892);
and U3928 (N_3928,N_3067,N_3459);
nand U3929 (N_3929,N_3186,N_3287);
xor U3930 (N_3930,N_3065,N_2924);
and U3931 (N_3931,N_2419,N_3464);
xnor U3932 (N_3932,N_2795,N_3417);
nor U3933 (N_3933,N_3073,N_2440);
nand U3934 (N_3934,N_3373,N_2546);
or U3935 (N_3935,N_3485,N_2562);
nand U3936 (N_3936,N_3306,N_2749);
nand U3937 (N_3937,N_3156,N_3292);
and U3938 (N_3938,N_2725,N_3526);
nor U3939 (N_3939,N_3374,N_2730);
and U3940 (N_3940,N_3575,N_2828);
nor U3941 (N_3941,N_3257,N_2918);
nand U3942 (N_3942,N_3084,N_3535);
and U3943 (N_3943,N_2429,N_3483);
nor U3944 (N_3944,N_3449,N_3368);
and U3945 (N_3945,N_2839,N_3299);
xor U3946 (N_3946,N_3241,N_3297);
and U3947 (N_3947,N_2571,N_2939);
or U3948 (N_3948,N_2935,N_2778);
xor U3949 (N_3949,N_2555,N_2537);
and U3950 (N_3950,N_3140,N_2905);
and U3951 (N_3951,N_3295,N_3286);
or U3952 (N_3952,N_2514,N_2955);
nor U3953 (N_3953,N_2989,N_3517);
nand U3954 (N_3954,N_2858,N_2575);
xnor U3955 (N_3955,N_2781,N_3165);
or U3956 (N_3956,N_3439,N_3583);
nand U3957 (N_3957,N_2598,N_2633);
xor U3958 (N_3958,N_3555,N_3363);
nand U3959 (N_3959,N_2475,N_3010);
nor U3960 (N_3960,N_3142,N_2817);
xnor U3961 (N_3961,N_3034,N_2645);
nand U3962 (N_3962,N_2944,N_3538);
nor U3963 (N_3963,N_3407,N_3452);
nand U3964 (N_3964,N_2616,N_3282);
nor U3965 (N_3965,N_3326,N_2623);
and U3966 (N_3966,N_3222,N_3330);
nand U3967 (N_3967,N_2474,N_2499);
nand U3968 (N_3968,N_2603,N_2609);
and U3969 (N_3969,N_2746,N_3060);
nor U3970 (N_3970,N_3506,N_2837);
xor U3971 (N_3971,N_2854,N_3113);
nand U3972 (N_3972,N_2509,N_2761);
and U3973 (N_3973,N_2614,N_3220);
and U3974 (N_3974,N_3499,N_3477);
nor U3975 (N_3975,N_2809,N_2869);
and U3976 (N_3976,N_3144,N_3579);
and U3977 (N_3977,N_2734,N_3049);
and U3978 (N_3978,N_2811,N_2714);
nand U3979 (N_3979,N_2942,N_3051);
and U3980 (N_3980,N_3455,N_2525);
nand U3981 (N_3981,N_3221,N_2772);
nor U3982 (N_3982,N_2435,N_2548);
and U3983 (N_3983,N_3017,N_2695);
or U3984 (N_3984,N_2709,N_2807);
nor U3985 (N_3985,N_3188,N_2574);
nor U3986 (N_3986,N_3005,N_2518);
nor U3987 (N_3987,N_2753,N_3582);
nor U3988 (N_3988,N_3527,N_3180);
xnor U3989 (N_3989,N_3043,N_3231);
and U3990 (N_3990,N_3549,N_3486);
xnor U3991 (N_3991,N_3378,N_3133);
and U3992 (N_3992,N_3006,N_2556);
nor U3993 (N_3993,N_3475,N_2415);
or U3994 (N_3994,N_3392,N_3279);
nor U3995 (N_3995,N_3597,N_2563);
nor U3996 (N_3996,N_3443,N_2875);
and U3997 (N_3997,N_2740,N_3425);
nor U3998 (N_3998,N_3132,N_2455);
or U3999 (N_3999,N_2782,N_3531);
and U4000 (N_4000,N_2492,N_2527);
or U4001 (N_4001,N_3003,N_2840);
and U4002 (N_4002,N_2925,N_3308);
and U4003 (N_4003,N_2494,N_3429);
and U4004 (N_4004,N_2599,N_3246);
xor U4005 (N_4005,N_2626,N_3075);
nand U4006 (N_4006,N_3042,N_2930);
nand U4007 (N_4007,N_3127,N_3170);
nor U4008 (N_4008,N_3028,N_3305);
and U4009 (N_4009,N_3463,N_3334);
or U4010 (N_4010,N_2547,N_2484);
or U4011 (N_4011,N_2408,N_3227);
and U4012 (N_4012,N_2831,N_2832);
or U4013 (N_4013,N_2994,N_2517);
nand U4014 (N_4014,N_2651,N_2888);
xor U4015 (N_4015,N_2447,N_2667);
and U4016 (N_4016,N_2874,N_2972);
nand U4017 (N_4017,N_2536,N_2402);
xor U4018 (N_4018,N_2724,N_3285);
nand U4019 (N_4019,N_2541,N_2886);
or U4020 (N_4020,N_3501,N_3097);
xnor U4021 (N_4021,N_3015,N_2544);
nand U4022 (N_4022,N_3273,N_3543);
and U4023 (N_4023,N_3390,N_3151);
nand U4024 (N_4024,N_2605,N_2431);
nor U4025 (N_4025,N_2752,N_2632);
nand U4026 (N_4026,N_2722,N_2568);
xnor U4027 (N_4027,N_3377,N_2448);
nor U4028 (N_4028,N_2773,N_3074);
xor U4029 (N_4029,N_2949,N_2691);
xor U4030 (N_4030,N_2444,N_3164);
or U4031 (N_4031,N_3190,N_2504);
nand U4032 (N_4032,N_3112,N_3229);
and U4033 (N_4033,N_3058,N_3163);
nor U4034 (N_4034,N_3311,N_2664);
nor U4035 (N_4035,N_3018,N_2987);
xor U4036 (N_4036,N_3509,N_2920);
or U4037 (N_4037,N_3589,N_2702);
and U4038 (N_4038,N_2487,N_2834);
or U4039 (N_4039,N_2815,N_3126);
xor U4040 (N_4040,N_3237,N_3367);
nand U4041 (N_4041,N_2496,N_2767);
nor U4042 (N_4042,N_2958,N_2757);
or U4043 (N_4043,N_2635,N_2796);
or U4044 (N_4044,N_2798,N_2538);
or U4045 (N_4045,N_2978,N_3409);
xnor U4046 (N_4046,N_2590,N_2433);
and U4047 (N_4047,N_3044,N_2950);
nor U4048 (N_4048,N_2692,N_2573);
and U4049 (N_4049,N_2774,N_3128);
xor U4050 (N_4050,N_2786,N_3542);
and U4051 (N_4051,N_3574,N_3375);
xnor U4052 (N_4052,N_2969,N_2943);
nand U4053 (N_4053,N_3096,N_2827);
and U4054 (N_4054,N_2582,N_3230);
and U4055 (N_4055,N_3566,N_2620);
and U4056 (N_4056,N_2545,N_3391);
nor U4057 (N_4057,N_2884,N_3491);
or U4058 (N_4058,N_3364,N_3209);
or U4059 (N_4059,N_3336,N_3398);
or U4060 (N_4060,N_2688,N_2936);
nor U4061 (N_4061,N_3497,N_3510);
nor U4062 (N_4062,N_3166,N_2897);
or U4063 (N_4063,N_2630,N_3007);
nand U4064 (N_4064,N_3223,N_3532);
or U4065 (N_4065,N_3244,N_2581);
xor U4066 (N_4066,N_3158,N_2910);
and U4067 (N_4067,N_2611,N_2606);
nand U4068 (N_4068,N_3251,N_2565);
or U4069 (N_4069,N_2529,N_3335);
nor U4070 (N_4070,N_2833,N_3119);
or U4071 (N_4071,N_3360,N_2926);
nand U4072 (N_4072,N_2769,N_3339);
nor U4073 (N_4073,N_2923,N_2883);
nor U4074 (N_4074,N_2787,N_2631);
and U4075 (N_4075,N_2822,N_3592);
or U4076 (N_4076,N_3465,N_2991);
or U4077 (N_4077,N_2550,N_3011);
or U4078 (N_4078,N_3068,N_2458);
or U4079 (N_4079,N_2763,N_3137);
or U4080 (N_4080,N_3466,N_2999);
nor U4081 (N_4081,N_2567,N_3379);
xnor U4082 (N_4082,N_3057,N_3048);
or U4083 (N_4083,N_2747,N_3515);
and U4084 (N_4084,N_2510,N_2584);
xnor U4085 (N_4085,N_2893,N_2801);
nor U4086 (N_4086,N_3366,N_2754);
nor U4087 (N_4087,N_3327,N_2860);
and U4088 (N_4088,N_3088,N_2657);
xnor U4089 (N_4089,N_2900,N_2403);
and U4090 (N_4090,N_3117,N_3022);
or U4091 (N_4091,N_3293,N_3310);
nor U4092 (N_4092,N_2934,N_2962);
xnor U4093 (N_4093,N_3470,N_3313);
nor U4094 (N_4094,N_2643,N_3125);
and U4095 (N_4095,N_3080,N_3242);
nand U4096 (N_4096,N_3309,N_3145);
xor U4097 (N_4097,N_2658,N_2829);
or U4098 (N_4098,N_3370,N_2519);
xnor U4099 (N_4099,N_2872,N_3234);
or U4100 (N_4100,N_3258,N_2735);
nand U4101 (N_4101,N_2618,N_2898);
or U4102 (N_4102,N_2619,N_2533);
or U4103 (N_4103,N_2414,N_3205);
and U4104 (N_4104,N_3124,N_3130);
or U4105 (N_4105,N_3284,N_3238);
xor U4106 (N_4106,N_2467,N_3383);
or U4107 (N_4107,N_2411,N_2591);
xor U4108 (N_4108,N_3300,N_3195);
or U4109 (N_4109,N_2820,N_3508);
nand U4110 (N_4110,N_2579,N_3194);
nand U4111 (N_4111,N_2634,N_3184);
xor U4112 (N_4112,N_2861,N_2889);
nor U4113 (N_4113,N_3564,N_3457);
xnor U4114 (N_4114,N_2686,N_3233);
and U4115 (N_4115,N_3414,N_3516);
and U4116 (N_4116,N_3108,N_2868);
and U4117 (N_4117,N_3411,N_3521);
nor U4118 (N_4118,N_3270,N_3359);
or U4119 (N_4119,N_3204,N_2554);
nand U4120 (N_4120,N_3261,N_2401);
or U4121 (N_4121,N_3468,N_2745);
xor U4122 (N_4122,N_2998,N_3460);
xor U4123 (N_4123,N_2812,N_2901);
or U4124 (N_4124,N_2503,N_2660);
nand U4125 (N_4125,N_3178,N_3431);
and U4126 (N_4126,N_3458,N_2405);
and U4127 (N_4127,N_3083,N_3502);
nand U4128 (N_4128,N_3387,N_2418);
nand U4129 (N_4129,N_3296,N_3029);
xnor U4130 (N_4130,N_2662,N_2922);
or U4131 (N_4131,N_3534,N_2507);
nand U4132 (N_4132,N_2813,N_2741);
or U4133 (N_4133,N_2915,N_2569);
xor U4134 (N_4134,N_3114,N_3358);
and U4135 (N_4135,N_2836,N_3341);
or U4136 (N_4136,N_3274,N_2542);
or U4137 (N_4137,N_3422,N_3495);
nor U4138 (N_4138,N_2980,N_2945);
and U4139 (N_4139,N_2983,N_3026);
xor U4140 (N_4140,N_3053,N_3101);
or U4141 (N_4141,N_3481,N_3121);
xnor U4142 (N_4142,N_3337,N_2593);
nand U4143 (N_4143,N_2771,N_2461);
xor U4144 (N_4144,N_2460,N_3529);
xor U4145 (N_4145,N_2560,N_2482);
or U4146 (N_4146,N_2676,N_2750);
or U4147 (N_4147,N_2551,N_3037);
and U4148 (N_4148,N_3100,N_2587);
and U4149 (N_4149,N_3064,N_2842);
or U4150 (N_4150,N_3563,N_3558);
xnor U4151 (N_4151,N_2756,N_2696);
nand U4152 (N_4152,N_3226,N_3456);
xor U4153 (N_4153,N_2683,N_2445);
or U4154 (N_4154,N_3565,N_3503);
nor U4155 (N_4155,N_3136,N_3427);
and U4156 (N_4156,N_2477,N_2449);
nand U4157 (N_4157,N_3418,N_3039);
nor U4158 (N_4158,N_3545,N_3317);
or U4159 (N_4159,N_2597,N_2646);
and U4160 (N_4160,N_3319,N_2968);
xnor U4161 (N_4161,N_3524,N_2432);
or U4162 (N_4162,N_3120,N_3147);
nand U4163 (N_4163,N_3033,N_3092);
nand U4164 (N_4164,N_3215,N_3009);
xnor U4165 (N_4165,N_3069,N_3289);
nor U4166 (N_4166,N_2744,N_2456);
nand U4167 (N_4167,N_2863,N_2951);
and U4168 (N_4168,N_3302,N_2404);
xnor U4169 (N_4169,N_3473,N_2770);
nor U4170 (N_4170,N_2726,N_3401);
nand U4171 (N_4171,N_2430,N_2727);
and U4172 (N_4172,N_3264,N_2572);
nor U4173 (N_4173,N_3599,N_3551);
or U4174 (N_4174,N_3152,N_2594);
nand U4175 (N_4175,N_3098,N_2929);
nand U4176 (N_4176,N_3272,N_2804);
xor U4177 (N_4177,N_2700,N_3004);
nor U4178 (N_4178,N_2908,N_2887);
or U4179 (N_4179,N_2871,N_2697);
xnor U4180 (N_4180,N_2566,N_2478);
or U4181 (N_4181,N_3584,N_3393);
and U4182 (N_4182,N_3143,N_3134);
xnor U4183 (N_4183,N_2463,N_3086);
nand U4184 (N_4184,N_3217,N_2679);
nor U4185 (N_4185,N_2666,N_2689);
and U4186 (N_4186,N_2589,N_2826);
or U4187 (N_4187,N_3325,N_2699);
and U4188 (N_4188,N_3047,N_3399);
or U4189 (N_4189,N_3208,N_3448);
nor U4190 (N_4190,N_3197,N_3569);
xor U4191 (N_4191,N_3262,N_3219);
and U4192 (N_4192,N_2921,N_3079);
and U4193 (N_4193,N_2409,N_3077);
xor U4194 (N_4194,N_3139,N_2865);
nor U4195 (N_4195,N_2601,N_2844);
or U4196 (N_4196,N_3203,N_2816);
nand U4197 (N_4197,N_3415,N_2803);
xor U4198 (N_4198,N_2857,N_3500);
or U4199 (N_4199,N_2452,N_3045);
nor U4200 (N_4200,N_3527,N_3436);
xor U4201 (N_4201,N_2999,N_2625);
xor U4202 (N_4202,N_3148,N_3356);
nor U4203 (N_4203,N_2724,N_3045);
and U4204 (N_4204,N_2434,N_2593);
or U4205 (N_4205,N_2686,N_3599);
xnor U4206 (N_4206,N_2953,N_3517);
xnor U4207 (N_4207,N_3201,N_2617);
and U4208 (N_4208,N_2959,N_3120);
nand U4209 (N_4209,N_2836,N_2986);
nor U4210 (N_4210,N_3596,N_2924);
and U4211 (N_4211,N_3528,N_3392);
and U4212 (N_4212,N_2515,N_3444);
nand U4213 (N_4213,N_3136,N_3152);
nor U4214 (N_4214,N_3348,N_2769);
or U4215 (N_4215,N_3460,N_3389);
and U4216 (N_4216,N_3429,N_2645);
nand U4217 (N_4217,N_2704,N_3299);
or U4218 (N_4218,N_2873,N_2491);
or U4219 (N_4219,N_2751,N_3136);
nor U4220 (N_4220,N_3070,N_2822);
or U4221 (N_4221,N_3349,N_3150);
xor U4222 (N_4222,N_3139,N_2461);
or U4223 (N_4223,N_3435,N_2910);
and U4224 (N_4224,N_3086,N_2617);
nor U4225 (N_4225,N_3466,N_2930);
and U4226 (N_4226,N_3554,N_3490);
nor U4227 (N_4227,N_2745,N_2688);
or U4228 (N_4228,N_2794,N_3273);
nand U4229 (N_4229,N_2710,N_2582);
nand U4230 (N_4230,N_2951,N_2463);
xor U4231 (N_4231,N_3535,N_3019);
or U4232 (N_4232,N_2833,N_2850);
nand U4233 (N_4233,N_3236,N_3308);
nand U4234 (N_4234,N_2585,N_3072);
nor U4235 (N_4235,N_3399,N_3311);
xnor U4236 (N_4236,N_2635,N_3406);
nor U4237 (N_4237,N_2411,N_3531);
xor U4238 (N_4238,N_3599,N_2788);
and U4239 (N_4239,N_3042,N_2916);
nand U4240 (N_4240,N_3557,N_2666);
nor U4241 (N_4241,N_3331,N_3365);
and U4242 (N_4242,N_2836,N_2955);
and U4243 (N_4243,N_2581,N_3074);
nor U4244 (N_4244,N_3163,N_2430);
or U4245 (N_4245,N_3573,N_2531);
nor U4246 (N_4246,N_3102,N_3089);
nand U4247 (N_4247,N_3418,N_2934);
nor U4248 (N_4248,N_3423,N_3429);
nand U4249 (N_4249,N_2641,N_2938);
and U4250 (N_4250,N_3410,N_2980);
nor U4251 (N_4251,N_2413,N_3424);
nand U4252 (N_4252,N_2525,N_3068);
xor U4253 (N_4253,N_2818,N_2415);
nor U4254 (N_4254,N_3144,N_3578);
nor U4255 (N_4255,N_2712,N_3169);
xor U4256 (N_4256,N_3235,N_3491);
xor U4257 (N_4257,N_2597,N_2552);
and U4258 (N_4258,N_2990,N_2704);
or U4259 (N_4259,N_2706,N_3261);
nand U4260 (N_4260,N_2660,N_2694);
nor U4261 (N_4261,N_2618,N_2984);
or U4262 (N_4262,N_2902,N_3262);
or U4263 (N_4263,N_3160,N_2559);
and U4264 (N_4264,N_2819,N_3034);
xnor U4265 (N_4265,N_2413,N_3423);
and U4266 (N_4266,N_2493,N_2458);
xor U4267 (N_4267,N_3253,N_3353);
nor U4268 (N_4268,N_3381,N_2477);
and U4269 (N_4269,N_2839,N_3348);
nand U4270 (N_4270,N_2842,N_2779);
nand U4271 (N_4271,N_3358,N_2702);
nand U4272 (N_4272,N_3472,N_2674);
nor U4273 (N_4273,N_3216,N_2591);
xnor U4274 (N_4274,N_2824,N_3229);
xnor U4275 (N_4275,N_3232,N_3521);
and U4276 (N_4276,N_3046,N_2616);
and U4277 (N_4277,N_2664,N_2621);
or U4278 (N_4278,N_3532,N_2658);
nand U4279 (N_4279,N_2838,N_2664);
nand U4280 (N_4280,N_3103,N_2750);
and U4281 (N_4281,N_2943,N_3387);
nor U4282 (N_4282,N_2477,N_2404);
nor U4283 (N_4283,N_3261,N_2439);
xor U4284 (N_4284,N_2720,N_2532);
nand U4285 (N_4285,N_2845,N_2573);
or U4286 (N_4286,N_3263,N_3254);
nor U4287 (N_4287,N_2680,N_2976);
nand U4288 (N_4288,N_2576,N_3278);
xnor U4289 (N_4289,N_2412,N_2773);
and U4290 (N_4290,N_2616,N_3559);
xnor U4291 (N_4291,N_3353,N_3269);
nand U4292 (N_4292,N_3041,N_3451);
or U4293 (N_4293,N_2777,N_2803);
and U4294 (N_4294,N_2934,N_2446);
xor U4295 (N_4295,N_3133,N_3426);
xor U4296 (N_4296,N_2740,N_3012);
or U4297 (N_4297,N_2808,N_2583);
nand U4298 (N_4298,N_3579,N_3431);
nand U4299 (N_4299,N_2462,N_3203);
xnor U4300 (N_4300,N_3568,N_2917);
nand U4301 (N_4301,N_2755,N_2568);
xnor U4302 (N_4302,N_2526,N_2831);
nor U4303 (N_4303,N_2595,N_2607);
or U4304 (N_4304,N_3413,N_2433);
nor U4305 (N_4305,N_3183,N_3233);
xnor U4306 (N_4306,N_2522,N_3194);
xor U4307 (N_4307,N_3046,N_2500);
and U4308 (N_4308,N_3030,N_2931);
nor U4309 (N_4309,N_2452,N_3257);
xnor U4310 (N_4310,N_3352,N_2425);
and U4311 (N_4311,N_3585,N_3021);
xnor U4312 (N_4312,N_3397,N_3405);
xnor U4313 (N_4313,N_2799,N_3231);
nor U4314 (N_4314,N_3151,N_2786);
nor U4315 (N_4315,N_3315,N_3408);
nor U4316 (N_4316,N_3151,N_3538);
nand U4317 (N_4317,N_2899,N_2677);
or U4318 (N_4318,N_2794,N_2572);
xnor U4319 (N_4319,N_2670,N_2654);
nand U4320 (N_4320,N_2604,N_2705);
nand U4321 (N_4321,N_2757,N_3485);
and U4322 (N_4322,N_2790,N_2514);
nand U4323 (N_4323,N_2873,N_2865);
or U4324 (N_4324,N_3564,N_3526);
and U4325 (N_4325,N_3203,N_2738);
nand U4326 (N_4326,N_2504,N_3119);
and U4327 (N_4327,N_2991,N_2844);
nor U4328 (N_4328,N_2475,N_3030);
and U4329 (N_4329,N_3134,N_3093);
nor U4330 (N_4330,N_2780,N_2613);
and U4331 (N_4331,N_3246,N_3440);
xnor U4332 (N_4332,N_3204,N_3039);
and U4333 (N_4333,N_2540,N_2923);
and U4334 (N_4334,N_3051,N_2925);
and U4335 (N_4335,N_3013,N_2665);
or U4336 (N_4336,N_2926,N_2744);
or U4337 (N_4337,N_2897,N_3468);
xnor U4338 (N_4338,N_2754,N_2512);
nor U4339 (N_4339,N_3543,N_2735);
or U4340 (N_4340,N_3239,N_2707);
nand U4341 (N_4341,N_2923,N_2935);
and U4342 (N_4342,N_2853,N_2976);
nand U4343 (N_4343,N_2511,N_2664);
nand U4344 (N_4344,N_2952,N_2594);
nor U4345 (N_4345,N_3402,N_2559);
and U4346 (N_4346,N_2981,N_3005);
or U4347 (N_4347,N_3117,N_2995);
or U4348 (N_4348,N_3534,N_2759);
xnor U4349 (N_4349,N_3574,N_2641);
nand U4350 (N_4350,N_2912,N_2811);
nand U4351 (N_4351,N_3259,N_3105);
or U4352 (N_4352,N_2763,N_3444);
or U4353 (N_4353,N_2856,N_2710);
nand U4354 (N_4354,N_2964,N_2697);
xnor U4355 (N_4355,N_2498,N_2990);
xor U4356 (N_4356,N_2946,N_3348);
and U4357 (N_4357,N_2534,N_2452);
nor U4358 (N_4358,N_2909,N_3294);
nand U4359 (N_4359,N_2457,N_2476);
nand U4360 (N_4360,N_3353,N_2674);
and U4361 (N_4361,N_3399,N_2496);
and U4362 (N_4362,N_2529,N_3472);
or U4363 (N_4363,N_2554,N_2925);
and U4364 (N_4364,N_2822,N_2764);
and U4365 (N_4365,N_2539,N_2414);
or U4366 (N_4366,N_2897,N_2483);
or U4367 (N_4367,N_3536,N_2544);
and U4368 (N_4368,N_2936,N_3483);
nand U4369 (N_4369,N_2412,N_3251);
nand U4370 (N_4370,N_3553,N_3079);
or U4371 (N_4371,N_3029,N_3171);
or U4372 (N_4372,N_3084,N_2832);
xor U4373 (N_4373,N_2886,N_3182);
and U4374 (N_4374,N_3498,N_2801);
xnor U4375 (N_4375,N_2990,N_3240);
and U4376 (N_4376,N_2718,N_2595);
xnor U4377 (N_4377,N_2973,N_2794);
nor U4378 (N_4378,N_2893,N_2423);
or U4379 (N_4379,N_3149,N_3373);
or U4380 (N_4380,N_2503,N_3160);
xnor U4381 (N_4381,N_2864,N_3349);
xnor U4382 (N_4382,N_3341,N_2501);
nor U4383 (N_4383,N_3191,N_3020);
or U4384 (N_4384,N_2981,N_3022);
or U4385 (N_4385,N_2746,N_3359);
nand U4386 (N_4386,N_3419,N_3196);
nand U4387 (N_4387,N_3586,N_3595);
nand U4388 (N_4388,N_2586,N_2770);
and U4389 (N_4389,N_3367,N_3005);
nand U4390 (N_4390,N_2837,N_2665);
nand U4391 (N_4391,N_2963,N_3127);
and U4392 (N_4392,N_3578,N_3492);
or U4393 (N_4393,N_2468,N_2993);
or U4394 (N_4394,N_3264,N_2646);
nor U4395 (N_4395,N_2446,N_2667);
nand U4396 (N_4396,N_3086,N_3473);
nor U4397 (N_4397,N_3557,N_3095);
nor U4398 (N_4398,N_2821,N_3393);
or U4399 (N_4399,N_3128,N_3266);
xnor U4400 (N_4400,N_3363,N_3361);
xor U4401 (N_4401,N_3074,N_3479);
and U4402 (N_4402,N_3504,N_2689);
nand U4403 (N_4403,N_2819,N_2540);
nand U4404 (N_4404,N_3004,N_3546);
or U4405 (N_4405,N_3170,N_2862);
nand U4406 (N_4406,N_3314,N_3007);
nor U4407 (N_4407,N_3574,N_3277);
and U4408 (N_4408,N_3500,N_3263);
and U4409 (N_4409,N_3073,N_3064);
xnor U4410 (N_4410,N_3062,N_2721);
nand U4411 (N_4411,N_3431,N_2583);
xnor U4412 (N_4412,N_3274,N_3345);
xnor U4413 (N_4413,N_3100,N_2406);
or U4414 (N_4414,N_2939,N_3522);
or U4415 (N_4415,N_2698,N_2448);
xor U4416 (N_4416,N_2697,N_3336);
nand U4417 (N_4417,N_2831,N_3469);
nand U4418 (N_4418,N_3416,N_3321);
and U4419 (N_4419,N_3495,N_2419);
xnor U4420 (N_4420,N_2659,N_3312);
xor U4421 (N_4421,N_3133,N_3030);
xnor U4422 (N_4422,N_3501,N_3480);
and U4423 (N_4423,N_2510,N_2994);
or U4424 (N_4424,N_2420,N_2581);
nor U4425 (N_4425,N_3432,N_3134);
and U4426 (N_4426,N_2853,N_3473);
nand U4427 (N_4427,N_2850,N_2659);
and U4428 (N_4428,N_2713,N_2470);
nand U4429 (N_4429,N_2752,N_2606);
or U4430 (N_4430,N_3478,N_3294);
nor U4431 (N_4431,N_3361,N_2578);
nor U4432 (N_4432,N_3467,N_3510);
nand U4433 (N_4433,N_3351,N_3293);
or U4434 (N_4434,N_2529,N_2917);
xnor U4435 (N_4435,N_2614,N_3404);
xnor U4436 (N_4436,N_3364,N_2676);
and U4437 (N_4437,N_2553,N_2599);
or U4438 (N_4438,N_2414,N_3283);
and U4439 (N_4439,N_3363,N_2853);
nand U4440 (N_4440,N_3052,N_2782);
nand U4441 (N_4441,N_2425,N_2565);
nor U4442 (N_4442,N_3414,N_2546);
nand U4443 (N_4443,N_2438,N_3521);
nor U4444 (N_4444,N_3288,N_3130);
or U4445 (N_4445,N_3258,N_3066);
xnor U4446 (N_4446,N_3342,N_3349);
nand U4447 (N_4447,N_3018,N_3030);
xnor U4448 (N_4448,N_3350,N_2434);
nand U4449 (N_4449,N_2993,N_3033);
and U4450 (N_4450,N_3549,N_3492);
xor U4451 (N_4451,N_3585,N_2491);
nand U4452 (N_4452,N_3466,N_2733);
or U4453 (N_4453,N_2542,N_3149);
nand U4454 (N_4454,N_2817,N_2547);
and U4455 (N_4455,N_2989,N_3401);
nor U4456 (N_4456,N_3184,N_3113);
and U4457 (N_4457,N_3408,N_3484);
nand U4458 (N_4458,N_3097,N_2864);
xnor U4459 (N_4459,N_3094,N_3400);
or U4460 (N_4460,N_3038,N_2546);
nor U4461 (N_4461,N_2490,N_3346);
xnor U4462 (N_4462,N_2938,N_2792);
nand U4463 (N_4463,N_2967,N_3451);
xnor U4464 (N_4464,N_2473,N_3203);
xnor U4465 (N_4465,N_2943,N_2584);
nor U4466 (N_4466,N_3573,N_2503);
nor U4467 (N_4467,N_2899,N_3505);
xor U4468 (N_4468,N_3357,N_3490);
and U4469 (N_4469,N_2414,N_2893);
xor U4470 (N_4470,N_2736,N_2856);
nor U4471 (N_4471,N_2410,N_3445);
and U4472 (N_4472,N_2852,N_2430);
nor U4473 (N_4473,N_3018,N_3042);
xnor U4474 (N_4474,N_3538,N_2614);
or U4475 (N_4475,N_2719,N_3513);
and U4476 (N_4476,N_2597,N_2530);
or U4477 (N_4477,N_3468,N_2911);
nor U4478 (N_4478,N_2810,N_2938);
or U4479 (N_4479,N_2959,N_3242);
or U4480 (N_4480,N_2774,N_3008);
and U4481 (N_4481,N_2475,N_3143);
or U4482 (N_4482,N_3297,N_3242);
or U4483 (N_4483,N_3155,N_3570);
and U4484 (N_4484,N_3216,N_3258);
nand U4485 (N_4485,N_3129,N_3476);
xor U4486 (N_4486,N_3114,N_3579);
xnor U4487 (N_4487,N_3005,N_2836);
nor U4488 (N_4488,N_2846,N_2425);
xnor U4489 (N_4489,N_2760,N_2642);
nor U4490 (N_4490,N_2790,N_2753);
nor U4491 (N_4491,N_2458,N_3454);
or U4492 (N_4492,N_3397,N_3269);
nand U4493 (N_4493,N_2688,N_3446);
or U4494 (N_4494,N_3396,N_2623);
nor U4495 (N_4495,N_3328,N_2866);
or U4496 (N_4496,N_2876,N_2434);
nor U4497 (N_4497,N_3357,N_3579);
and U4498 (N_4498,N_3537,N_3305);
and U4499 (N_4499,N_2742,N_3033);
nor U4500 (N_4500,N_3153,N_2959);
nand U4501 (N_4501,N_2596,N_3407);
and U4502 (N_4502,N_3420,N_3384);
xnor U4503 (N_4503,N_3287,N_3227);
nor U4504 (N_4504,N_3314,N_3110);
xor U4505 (N_4505,N_2453,N_2971);
nor U4506 (N_4506,N_2771,N_2899);
and U4507 (N_4507,N_2872,N_3084);
or U4508 (N_4508,N_3479,N_2527);
xnor U4509 (N_4509,N_3031,N_2803);
and U4510 (N_4510,N_3564,N_2793);
nor U4511 (N_4511,N_3243,N_3391);
or U4512 (N_4512,N_3131,N_2909);
nor U4513 (N_4513,N_3594,N_3048);
and U4514 (N_4514,N_2884,N_2653);
nand U4515 (N_4515,N_3481,N_3107);
and U4516 (N_4516,N_3468,N_2636);
nand U4517 (N_4517,N_2794,N_2595);
xnor U4518 (N_4518,N_3426,N_2777);
and U4519 (N_4519,N_2996,N_2589);
nor U4520 (N_4520,N_2975,N_2721);
or U4521 (N_4521,N_3226,N_2734);
and U4522 (N_4522,N_3016,N_3070);
and U4523 (N_4523,N_2529,N_2619);
nor U4524 (N_4524,N_2772,N_3524);
and U4525 (N_4525,N_2628,N_3425);
and U4526 (N_4526,N_3512,N_2877);
nor U4527 (N_4527,N_3073,N_2666);
nand U4528 (N_4528,N_2589,N_3467);
nor U4529 (N_4529,N_3196,N_2563);
and U4530 (N_4530,N_3201,N_2757);
and U4531 (N_4531,N_3464,N_2529);
and U4532 (N_4532,N_2656,N_2834);
or U4533 (N_4533,N_2485,N_2872);
nor U4534 (N_4534,N_2477,N_2695);
xor U4535 (N_4535,N_3126,N_2911);
and U4536 (N_4536,N_3312,N_3136);
nor U4537 (N_4537,N_2872,N_2997);
nor U4538 (N_4538,N_3011,N_3115);
xor U4539 (N_4539,N_3466,N_2862);
nor U4540 (N_4540,N_3283,N_2643);
nand U4541 (N_4541,N_3526,N_2927);
or U4542 (N_4542,N_2769,N_3306);
xnor U4543 (N_4543,N_3348,N_2694);
or U4544 (N_4544,N_2425,N_2490);
nor U4545 (N_4545,N_3469,N_3162);
xnor U4546 (N_4546,N_2827,N_3308);
nand U4547 (N_4547,N_3411,N_3112);
nand U4548 (N_4548,N_2402,N_2572);
or U4549 (N_4549,N_2990,N_3253);
and U4550 (N_4550,N_2920,N_3027);
or U4551 (N_4551,N_2783,N_2599);
or U4552 (N_4552,N_2605,N_2479);
and U4553 (N_4553,N_2479,N_3383);
nor U4554 (N_4554,N_2741,N_2861);
and U4555 (N_4555,N_3041,N_2966);
and U4556 (N_4556,N_2743,N_3330);
xnor U4557 (N_4557,N_3381,N_3065);
nand U4558 (N_4558,N_3446,N_2776);
nor U4559 (N_4559,N_3114,N_2923);
xor U4560 (N_4560,N_3248,N_3285);
nand U4561 (N_4561,N_2577,N_2526);
or U4562 (N_4562,N_3335,N_3118);
nor U4563 (N_4563,N_2820,N_3104);
or U4564 (N_4564,N_3318,N_2835);
nand U4565 (N_4565,N_2864,N_2944);
xor U4566 (N_4566,N_2678,N_2898);
nor U4567 (N_4567,N_3565,N_3354);
nor U4568 (N_4568,N_2578,N_2825);
nor U4569 (N_4569,N_3269,N_3033);
nor U4570 (N_4570,N_2609,N_2589);
xor U4571 (N_4571,N_2737,N_2859);
and U4572 (N_4572,N_3450,N_2502);
nor U4573 (N_4573,N_3264,N_2961);
or U4574 (N_4574,N_3105,N_2797);
or U4575 (N_4575,N_3020,N_2552);
nor U4576 (N_4576,N_3035,N_2703);
or U4577 (N_4577,N_2542,N_3378);
nand U4578 (N_4578,N_3006,N_3202);
xnor U4579 (N_4579,N_3149,N_3309);
or U4580 (N_4580,N_3255,N_2978);
and U4581 (N_4581,N_2820,N_2590);
nor U4582 (N_4582,N_3216,N_2704);
nand U4583 (N_4583,N_3193,N_2637);
nand U4584 (N_4584,N_2952,N_3117);
nor U4585 (N_4585,N_3508,N_2507);
nand U4586 (N_4586,N_3426,N_2423);
or U4587 (N_4587,N_3056,N_3583);
xor U4588 (N_4588,N_2771,N_2919);
or U4589 (N_4589,N_2582,N_3388);
nand U4590 (N_4590,N_3412,N_2509);
xnor U4591 (N_4591,N_2988,N_2942);
xnor U4592 (N_4592,N_2521,N_2548);
or U4593 (N_4593,N_3114,N_3313);
xnor U4594 (N_4594,N_3335,N_2549);
xor U4595 (N_4595,N_2499,N_3327);
xnor U4596 (N_4596,N_3130,N_3171);
and U4597 (N_4597,N_3435,N_2953);
nor U4598 (N_4598,N_3125,N_3487);
xnor U4599 (N_4599,N_2429,N_2886);
or U4600 (N_4600,N_3092,N_2440);
nand U4601 (N_4601,N_3046,N_2732);
nand U4602 (N_4602,N_2664,N_3519);
and U4603 (N_4603,N_3034,N_3596);
and U4604 (N_4604,N_2597,N_3117);
xor U4605 (N_4605,N_3200,N_2730);
xor U4606 (N_4606,N_3138,N_2446);
or U4607 (N_4607,N_2767,N_3389);
nand U4608 (N_4608,N_2781,N_2733);
or U4609 (N_4609,N_3062,N_3356);
or U4610 (N_4610,N_3329,N_2629);
and U4611 (N_4611,N_2616,N_3200);
nor U4612 (N_4612,N_3241,N_2424);
nor U4613 (N_4613,N_3183,N_3044);
and U4614 (N_4614,N_2751,N_3040);
and U4615 (N_4615,N_2537,N_2657);
nand U4616 (N_4616,N_3515,N_3539);
or U4617 (N_4617,N_3433,N_3337);
nand U4618 (N_4618,N_3347,N_2576);
nand U4619 (N_4619,N_3585,N_2702);
nand U4620 (N_4620,N_3535,N_2558);
or U4621 (N_4621,N_2479,N_3059);
nand U4622 (N_4622,N_2536,N_3008);
or U4623 (N_4623,N_2926,N_2757);
nor U4624 (N_4624,N_3033,N_2488);
and U4625 (N_4625,N_2835,N_3230);
xnor U4626 (N_4626,N_2562,N_2900);
or U4627 (N_4627,N_2761,N_3196);
or U4628 (N_4628,N_3122,N_3115);
and U4629 (N_4629,N_2763,N_3072);
nand U4630 (N_4630,N_3000,N_2812);
and U4631 (N_4631,N_2502,N_3312);
or U4632 (N_4632,N_2827,N_3536);
xor U4633 (N_4633,N_3242,N_2547);
nand U4634 (N_4634,N_2459,N_2718);
nor U4635 (N_4635,N_2777,N_3580);
or U4636 (N_4636,N_2627,N_3225);
nor U4637 (N_4637,N_2641,N_3224);
or U4638 (N_4638,N_3472,N_3243);
or U4639 (N_4639,N_3408,N_2425);
nand U4640 (N_4640,N_2905,N_2670);
nor U4641 (N_4641,N_3492,N_3588);
nor U4642 (N_4642,N_2816,N_3590);
nand U4643 (N_4643,N_2604,N_2833);
nand U4644 (N_4644,N_3091,N_3041);
nand U4645 (N_4645,N_3358,N_3315);
and U4646 (N_4646,N_2724,N_3222);
or U4647 (N_4647,N_3209,N_3210);
nor U4648 (N_4648,N_2475,N_2677);
nand U4649 (N_4649,N_2603,N_3198);
or U4650 (N_4650,N_2735,N_3303);
or U4651 (N_4651,N_3084,N_3530);
nand U4652 (N_4652,N_2725,N_3576);
nand U4653 (N_4653,N_2417,N_2671);
or U4654 (N_4654,N_3329,N_2435);
xnor U4655 (N_4655,N_3277,N_3457);
xnor U4656 (N_4656,N_2884,N_3234);
xor U4657 (N_4657,N_2973,N_3170);
xnor U4658 (N_4658,N_3577,N_2530);
and U4659 (N_4659,N_2404,N_2838);
or U4660 (N_4660,N_2857,N_3215);
nand U4661 (N_4661,N_2498,N_3023);
and U4662 (N_4662,N_3313,N_3257);
nor U4663 (N_4663,N_3117,N_2723);
or U4664 (N_4664,N_2493,N_2603);
nor U4665 (N_4665,N_3113,N_3144);
or U4666 (N_4666,N_3506,N_3209);
and U4667 (N_4667,N_2490,N_3050);
nor U4668 (N_4668,N_3114,N_2779);
and U4669 (N_4669,N_2446,N_2986);
or U4670 (N_4670,N_3062,N_2512);
nand U4671 (N_4671,N_2960,N_2455);
nand U4672 (N_4672,N_3386,N_3213);
xnor U4673 (N_4673,N_2551,N_2850);
nand U4674 (N_4674,N_2752,N_2767);
xnor U4675 (N_4675,N_2834,N_3410);
nand U4676 (N_4676,N_2929,N_2734);
nand U4677 (N_4677,N_3524,N_2494);
nor U4678 (N_4678,N_2750,N_3083);
nor U4679 (N_4679,N_2970,N_2781);
nor U4680 (N_4680,N_2927,N_3148);
xor U4681 (N_4681,N_2744,N_2604);
or U4682 (N_4682,N_2887,N_2964);
nor U4683 (N_4683,N_2880,N_2825);
xor U4684 (N_4684,N_3583,N_3308);
nor U4685 (N_4685,N_2542,N_3043);
nor U4686 (N_4686,N_2648,N_3243);
or U4687 (N_4687,N_2984,N_2651);
nand U4688 (N_4688,N_3531,N_2852);
and U4689 (N_4689,N_3025,N_2875);
and U4690 (N_4690,N_3409,N_3332);
nand U4691 (N_4691,N_2589,N_2782);
nor U4692 (N_4692,N_3273,N_3510);
or U4693 (N_4693,N_3054,N_3169);
nand U4694 (N_4694,N_2850,N_3528);
or U4695 (N_4695,N_2861,N_2664);
xnor U4696 (N_4696,N_3569,N_2502);
xor U4697 (N_4697,N_2523,N_2475);
nand U4698 (N_4698,N_2866,N_3135);
nand U4699 (N_4699,N_3361,N_2735);
xor U4700 (N_4700,N_3402,N_3204);
or U4701 (N_4701,N_3592,N_3304);
and U4702 (N_4702,N_3449,N_2987);
nor U4703 (N_4703,N_2957,N_2557);
nand U4704 (N_4704,N_3328,N_3577);
xnor U4705 (N_4705,N_3574,N_3490);
nand U4706 (N_4706,N_2626,N_3004);
nand U4707 (N_4707,N_2708,N_3433);
nor U4708 (N_4708,N_2853,N_2662);
and U4709 (N_4709,N_2554,N_2775);
nor U4710 (N_4710,N_2514,N_2804);
nor U4711 (N_4711,N_3008,N_2888);
xnor U4712 (N_4712,N_3070,N_2796);
nand U4713 (N_4713,N_3422,N_2532);
xnor U4714 (N_4714,N_2941,N_3400);
and U4715 (N_4715,N_2978,N_3488);
and U4716 (N_4716,N_2930,N_2940);
nand U4717 (N_4717,N_2636,N_3143);
nor U4718 (N_4718,N_2445,N_3236);
nor U4719 (N_4719,N_3227,N_2667);
nor U4720 (N_4720,N_2961,N_3007);
nand U4721 (N_4721,N_2476,N_2721);
nand U4722 (N_4722,N_2777,N_3378);
and U4723 (N_4723,N_3186,N_3216);
or U4724 (N_4724,N_2915,N_3466);
xnor U4725 (N_4725,N_2525,N_2693);
nand U4726 (N_4726,N_3470,N_3116);
and U4727 (N_4727,N_3258,N_3106);
and U4728 (N_4728,N_2925,N_2795);
nand U4729 (N_4729,N_2617,N_3120);
xnor U4730 (N_4730,N_2547,N_3352);
nor U4731 (N_4731,N_2799,N_3117);
nand U4732 (N_4732,N_3310,N_3314);
or U4733 (N_4733,N_2509,N_2430);
nand U4734 (N_4734,N_2971,N_2861);
or U4735 (N_4735,N_2534,N_3194);
or U4736 (N_4736,N_3158,N_3024);
and U4737 (N_4737,N_3341,N_2977);
and U4738 (N_4738,N_3028,N_3434);
or U4739 (N_4739,N_3075,N_2916);
nand U4740 (N_4740,N_2658,N_3306);
nand U4741 (N_4741,N_2501,N_3070);
nand U4742 (N_4742,N_3333,N_2693);
or U4743 (N_4743,N_2562,N_2811);
and U4744 (N_4744,N_2867,N_2703);
or U4745 (N_4745,N_3009,N_2798);
and U4746 (N_4746,N_3119,N_3394);
nor U4747 (N_4747,N_3177,N_3516);
xnor U4748 (N_4748,N_2411,N_2596);
nor U4749 (N_4749,N_2805,N_2643);
nor U4750 (N_4750,N_3138,N_3424);
or U4751 (N_4751,N_3271,N_3211);
nor U4752 (N_4752,N_3583,N_3386);
nor U4753 (N_4753,N_3388,N_2866);
nor U4754 (N_4754,N_3305,N_3211);
nand U4755 (N_4755,N_3310,N_2879);
nand U4756 (N_4756,N_2952,N_2891);
nand U4757 (N_4757,N_2437,N_2430);
and U4758 (N_4758,N_2915,N_2962);
xnor U4759 (N_4759,N_2806,N_3173);
nor U4760 (N_4760,N_3346,N_2541);
and U4761 (N_4761,N_2407,N_2645);
xor U4762 (N_4762,N_3337,N_3330);
or U4763 (N_4763,N_3443,N_2990);
xor U4764 (N_4764,N_3590,N_2782);
xnor U4765 (N_4765,N_3083,N_3521);
nand U4766 (N_4766,N_3399,N_3290);
or U4767 (N_4767,N_3333,N_2535);
nand U4768 (N_4768,N_3362,N_2720);
or U4769 (N_4769,N_3222,N_3500);
xnor U4770 (N_4770,N_3383,N_2973);
or U4771 (N_4771,N_2448,N_2518);
or U4772 (N_4772,N_3205,N_2453);
or U4773 (N_4773,N_2518,N_2642);
xnor U4774 (N_4774,N_2672,N_2568);
xor U4775 (N_4775,N_2514,N_2982);
xnor U4776 (N_4776,N_2800,N_2864);
nand U4777 (N_4777,N_2953,N_2859);
and U4778 (N_4778,N_3228,N_3596);
nor U4779 (N_4779,N_3005,N_3022);
xnor U4780 (N_4780,N_2983,N_2776);
and U4781 (N_4781,N_2695,N_2886);
nor U4782 (N_4782,N_2816,N_2695);
or U4783 (N_4783,N_3466,N_2614);
or U4784 (N_4784,N_2981,N_3361);
nand U4785 (N_4785,N_3470,N_3024);
or U4786 (N_4786,N_3286,N_3155);
nand U4787 (N_4787,N_2589,N_2786);
xnor U4788 (N_4788,N_3439,N_3540);
or U4789 (N_4789,N_3411,N_2646);
nand U4790 (N_4790,N_3316,N_2704);
nand U4791 (N_4791,N_2716,N_2700);
or U4792 (N_4792,N_3075,N_2868);
or U4793 (N_4793,N_2617,N_3044);
nor U4794 (N_4794,N_3287,N_2707);
nand U4795 (N_4795,N_2562,N_2736);
nand U4796 (N_4796,N_2509,N_3463);
and U4797 (N_4797,N_3368,N_2843);
or U4798 (N_4798,N_2689,N_3275);
nor U4799 (N_4799,N_3392,N_3530);
nand U4800 (N_4800,N_3703,N_4784);
nor U4801 (N_4801,N_3689,N_3721);
and U4802 (N_4802,N_4709,N_4086);
nor U4803 (N_4803,N_4555,N_4250);
or U4804 (N_4804,N_4616,N_3962);
or U4805 (N_4805,N_4262,N_4290);
or U4806 (N_4806,N_3883,N_3771);
or U4807 (N_4807,N_4780,N_4260);
nand U4808 (N_4808,N_4622,N_4657);
nand U4809 (N_4809,N_4381,N_4289);
or U4810 (N_4810,N_4793,N_4462);
or U4811 (N_4811,N_3914,N_4229);
nand U4812 (N_4812,N_3978,N_4483);
or U4813 (N_4813,N_4062,N_3670);
xor U4814 (N_4814,N_4016,N_3902);
and U4815 (N_4815,N_4702,N_4334);
and U4816 (N_4816,N_3744,N_4195);
and U4817 (N_4817,N_4478,N_4190);
or U4818 (N_4818,N_4186,N_4496);
or U4819 (N_4819,N_4614,N_4067);
and U4820 (N_4820,N_4365,N_3822);
xor U4821 (N_4821,N_4569,N_3851);
nor U4822 (N_4822,N_4233,N_4448);
or U4823 (N_4823,N_4258,N_4751);
nor U4824 (N_4824,N_4240,N_4690);
or U4825 (N_4825,N_4563,N_4313);
or U4826 (N_4826,N_4304,N_4630);
nand U4827 (N_4827,N_3873,N_4459);
xor U4828 (N_4828,N_4161,N_4577);
or U4829 (N_4829,N_3664,N_4201);
or U4830 (N_4830,N_4378,N_4032);
or U4831 (N_4831,N_3789,N_3903);
nor U4832 (N_4832,N_3956,N_4398);
and U4833 (N_4833,N_4532,N_3706);
xnor U4834 (N_4834,N_4183,N_4714);
or U4835 (N_4835,N_3616,N_3986);
and U4836 (N_4836,N_3880,N_4036);
or U4837 (N_4837,N_4404,N_3815);
or U4838 (N_4838,N_4627,N_3623);
nor U4839 (N_4839,N_3655,N_3724);
nor U4840 (N_4840,N_4232,N_3723);
nand U4841 (N_4841,N_3869,N_4344);
xnor U4842 (N_4842,N_3989,N_4674);
or U4843 (N_4843,N_4643,N_4668);
xor U4844 (N_4844,N_4533,N_4150);
xor U4845 (N_4845,N_4468,N_3842);
nand U4846 (N_4846,N_3625,N_4717);
nand U4847 (N_4847,N_4427,N_4184);
xor U4848 (N_4848,N_4299,N_4571);
or U4849 (N_4849,N_3618,N_3942);
and U4850 (N_4850,N_3933,N_4601);
or U4851 (N_4851,N_4442,N_4768);
nor U4852 (N_4852,N_3887,N_3839);
nor U4853 (N_4853,N_4343,N_3997);
xor U4854 (N_4854,N_3982,N_4306);
nor U4855 (N_4855,N_4749,N_3940);
nand U4856 (N_4856,N_4742,N_3761);
nand U4857 (N_4857,N_3961,N_3938);
nand U4858 (N_4858,N_4659,N_3969);
and U4859 (N_4859,N_4409,N_3679);
nand U4860 (N_4860,N_4118,N_4175);
and U4861 (N_4861,N_4314,N_4537);
nand U4862 (N_4862,N_4082,N_4417);
or U4863 (N_4863,N_4511,N_4598);
nand U4864 (N_4864,N_4697,N_3926);
and U4865 (N_4865,N_4239,N_4738);
xor U4866 (N_4866,N_3830,N_3620);
nor U4867 (N_4867,N_4222,N_4341);
nand U4868 (N_4868,N_4715,N_4597);
and U4869 (N_4869,N_4434,N_3888);
and U4870 (N_4870,N_4154,N_4582);
or U4871 (N_4871,N_3717,N_4047);
xor U4872 (N_4872,N_4642,N_3973);
nand U4873 (N_4873,N_4469,N_4028);
nand U4874 (N_4874,N_4531,N_4429);
xor U4875 (N_4875,N_4733,N_3751);
nand U4876 (N_4876,N_3658,N_4633);
xnor U4877 (N_4877,N_3635,N_3649);
and U4878 (N_4878,N_3777,N_3954);
and U4879 (N_4879,N_3811,N_4333);
or U4880 (N_4880,N_4441,N_4599);
and U4881 (N_4881,N_3629,N_4631);
xor U4882 (N_4882,N_3638,N_3661);
nor U4883 (N_4883,N_4484,N_4710);
xor U4884 (N_4884,N_4579,N_3798);
or U4885 (N_4885,N_4741,N_4688);
and U4886 (N_4886,N_3829,N_3603);
xor U4887 (N_4887,N_4358,N_4416);
nor U4888 (N_4888,N_4595,N_3824);
or U4889 (N_4889,N_3628,N_4042);
nor U4890 (N_4890,N_4237,N_4162);
and U4891 (N_4891,N_3781,N_3801);
xnor U4892 (N_4892,N_3901,N_4449);
nand U4893 (N_4893,N_3944,N_4330);
nor U4894 (N_4894,N_4522,N_3684);
nand U4895 (N_4895,N_4506,N_4782);
nand U4896 (N_4896,N_4747,N_3810);
or U4897 (N_4897,N_4009,N_4744);
xnor U4898 (N_4898,N_4193,N_3736);
and U4899 (N_4899,N_4084,N_3610);
nor U4900 (N_4900,N_4074,N_4263);
and U4901 (N_4901,N_4406,N_4624);
nand U4902 (N_4902,N_3785,N_4418);
and U4903 (N_4903,N_4320,N_4148);
nand U4904 (N_4904,N_3674,N_4603);
or U4905 (N_4905,N_3870,N_4346);
and U4906 (N_4906,N_4165,N_3720);
nand U4907 (N_4907,N_4374,N_4310);
and U4908 (N_4908,N_4251,N_3795);
nor U4909 (N_4909,N_4058,N_3890);
xor U4910 (N_4910,N_4583,N_4700);
and U4911 (N_4911,N_4575,N_4167);
nor U4912 (N_4912,N_3714,N_4559);
and U4913 (N_4913,N_4670,N_4094);
xor U4914 (N_4914,N_3860,N_4737);
nand U4915 (N_4915,N_4644,N_3974);
xor U4916 (N_4916,N_4705,N_3841);
nor U4917 (N_4917,N_4486,N_3945);
nor U4918 (N_4918,N_4281,N_4127);
or U4919 (N_4919,N_4109,N_4408);
xnor U4920 (N_4920,N_4147,N_4463);
xnor U4921 (N_4921,N_4097,N_3791);
xor U4922 (N_4922,N_3696,N_3899);
xor U4923 (N_4923,N_4133,N_4671);
and U4924 (N_4924,N_4128,N_4101);
nor U4925 (N_4925,N_3763,N_4301);
nand U4926 (N_4926,N_4116,N_4022);
nor U4927 (N_4927,N_4662,N_4460);
nor U4928 (N_4928,N_3906,N_4187);
nand U4929 (N_4929,N_4445,N_4266);
nor U4930 (N_4930,N_4725,N_4581);
and U4931 (N_4931,N_4777,N_4092);
or U4932 (N_4932,N_3701,N_3951);
or U4933 (N_4933,N_4479,N_4695);
and U4934 (N_4934,N_4321,N_4414);
xor U4935 (N_4935,N_4179,N_4376);
or U4936 (N_4936,N_4159,N_3650);
and U4937 (N_4937,N_4748,N_3636);
xor U4938 (N_4938,N_3931,N_4057);
or U4939 (N_4939,N_3715,N_4399);
nor U4940 (N_4940,N_4040,N_4099);
or U4941 (N_4941,N_4061,N_4206);
and U4942 (N_4942,N_3915,N_4396);
or U4943 (N_4943,N_4231,N_3900);
xnor U4944 (N_4944,N_4561,N_4795);
nand U4945 (N_4945,N_4353,N_4403);
or U4946 (N_4946,N_3921,N_3957);
or U4947 (N_4947,N_4509,N_4743);
nand U4948 (N_4948,N_4589,N_4072);
and U4949 (N_4949,N_4491,N_4523);
and U4950 (N_4950,N_4540,N_3773);
or U4951 (N_4951,N_3834,N_3621);
or U4952 (N_4952,N_3964,N_3927);
nor U4953 (N_4953,N_4004,N_4323);
nor U4954 (N_4954,N_3632,N_3686);
xor U4955 (N_4955,N_4080,N_3861);
and U4956 (N_4956,N_3600,N_3939);
nor U4957 (N_4957,N_3608,N_3754);
nand U4958 (N_4958,N_4536,N_3960);
nor U4959 (N_4959,N_3971,N_4046);
and U4960 (N_4960,N_4108,N_4730);
nand U4961 (N_4961,N_4421,N_4703);
xnor U4962 (N_4962,N_4055,N_4636);
and U4963 (N_4963,N_4005,N_4146);
nand U4964 (N_4964,N_4329,N_4543);
xnor U4965 (N_4965,N_4213,N_4174);
xor U4966 (N_4966,N_4664,N_4349);
or U4967 (N_4967,N_4497,N_4166);
or U4968 (N_4968,N_3672,N_4485);
nand U4969 (N_4969,N_4384,N_4584);
and U4970 (N_4970,N_3687,N_3980);
xnor U4971 (N_4971,N_4767,N_4255);
or U4972 (N_4972,N_3683,N_4656);
or U4973 (N_4973,N_3845,N_3749);
or U4974 (N_4974,N_4124,N_4752);
nand U4975 (N_4975,N_4593,N_3750);
xnor U4976 (N_4976,N_4017,N_4401);
or U4977 (N_4977,N_4711,N_4424);
and U4978 (N_4978,N_3802,N_4140);
xor U4979 (N_4979,N_4574,N_4171);
or U4980 (N_4980,N_4367,N_4254);
nor U4981 (N_4981,N_3924,N_3659);
nand U4982 (N_4982,N_4006,N_3646);
nor U4983 (N_4983,N_3850,N_4775);
xor U4984 (N_4984,N_3866,N_4447);
and U4985 (N_4985,N_4383,N_4771);
xor U4986 (N_4986,N_4214,N_4692);
nand U4987 (N_4987,N_4432,N_4450);
xor U4988 (N_4988,N_4189,N_3837);
nand U4989 (N_4989,N_4235,N_4655);
or U4990 (N_4990,N_3871,N_4617);
xor U4991 (N_4991,N_4436,N_4437);
xnor U4992 (N_4992,N_4488,N_4219);
or U4993 (N_4993,N_3775,N_4490);
nor U4994 (N_4994,N_3808,N_3746);
and U4995 (N_4995,N_3748,N_4267);
or U4996 (N_4996,N_4474,N_4694);
nor U4997 (N_4997,N_4269,N_4528);
or U4998 (N_4998,N_4168,N_3996);
nor U4999 (N_4999,N_4699,N_4363);
or U5000 (N_5000,N_4691,N_3694);
xor U5001 (N_5001,N_3799,N_4209);
or U5002 (N_5002,N_3709,N_4362);
nor U5003 (N_5003,N_4088,N_4008);
nor U5004 (N_5004,N_3642,N_3886);
or U5005 (N_5005,N_3657,N_4562);
or U5006 (N_5006,N_4407,N_4188);
nor U5007 (N_5007,N_3852,N_3963);
or U5008 (N_5008,N_4014,N_4081);
or U5009 (N_5009,N_4298,N_3897);
nor U5010 (N_5010,N_3735,N_3784);
nand U5011 (N_5011,N_4173,N_4719);
nand U5012 (N_5012,N_4316,N_4212);
xnor U5013 (N_5013,N_4785,N_4535);
nand U5014 (N_5014,N_4024,N_3865);
nor U5015 (N_5015,N_4618,N_3609);
and U5016 (N_5016,N_4023,N_4020);
nor U5017 (N_5017,N_3946,N_3738);
xor U5018 (N_5018,N_3849,N_3611);
xnor U5019 (N_5019,N_3966,N_4202);
and U5020 (N_5020,N_4294,N_3624);
and U5021 (N_5021,N_4292,N_4610);
and U5022 (N_5022,N_4735,N_4572);
nand U5023 (N_5023,N_3941,N_3947);
and U5024 (N_5024,N_4380,N_4591);
and U5025 (N_5025,N_4707,N_4324);
xnor U5026 (N_5026,N_3698,N_4275);
nor U5027 (N_5027,N_4736,N_4625);
and U5028 (N_5028,N_3937,N_3695);
xor U5029 (N_5029,N_4286,N_4033);
nor U5030 (N_5030,N_4120,N_3949);
nand U5031 (N_5031,N_4687,N_4477);
nand U5032 (N_5032,N_3640,N_4600);
xor U5033 (N_5033,N_4514,N_4044);
and U5034 (N_5034,N_4273,N_4221);
nand U5035 (N_5035,N_4370,N_3772);
nand U5036 (N_5036,N_4287,N_4745);
xnor U5037 (N_5037,N_4282,N_4753);
and U5038 (N_5038,N_4686,N_3627);
and U5039 (N_5039,N_4180,N_4673);
nor U5040 (N_5040,N_4181,N_3797);
or U5041 (N_5041,N_3745,N_3923);
or U5042 (N_5042,N_3615,N_4428);
nor U5043 (N_5043,N_4327,N_3668);
or U5044 (N_5044,N_4556,N_3848);
and U5045 (N_5045,N_4170,N_4666);
xor U5046 (N_5046,N_3863,N_4520);
or U5047 (N_5047,N_4051,N_3948);
xor U5048 (N_5048,N_4345,N_3836);
nand U5049 (N_5049,N_3958,N_4297);
nand U5050 (N_5050,N_3663,N_4645);
nand U5051 (N_5051,N_4143,N_4243);
nand U5052 (N_5052,N_4355,N_4245);
and U5053 (N_5053,N_4356,N_4456);
nor U5054 (N_5054,N_4728,N_3809);
and U5055 (N_5055,N_3652,N_4669);
nand U5056 (N_5056,N_3952,N_4724);
nand U5057 (N_5057,N_4592,N_4368);
nor U5058 (N_5058,N_4156,N_4546);
and U5059 (N_5059,N_4198,N_3794);
and U5060 (N_5060,N_3855,N_3867);
nor U5061 (N_5061,N_4492,N_4142);
xnor U5062 (N_5062,N_4003,N_4137);
nor U5063 (N_5063,N_3700,N_4420);
and U5064 (N_5064,N_4204,N_4185);
nor U5065 (N_5065,N_4056,N_4538);
nand U5066 (N_5066,N_4471,N_4089);
and U5067 (N_5067,N_4604,N_3828);
xnor U5068 (N_5068,N_4034,N_4236);
nand U5069 (N_5069,N_4696,N_4394);
xnor U5070 (N_5070,N_4387,N_4721);
nor U5071 (N_5071,N_4426,N_4586);
or U5072 (N_5072,N_4757,N_4620);
nand U5073 (N_5073,N_3666,N_3846);
xnor U5074 (N_5074,N_4435,N_4663);
nand U5075 (N_5075,N_3677,N_4015);
or U5076 (N_5076,N_4489,N_4508);
and U5077 (N_5077,N_4457,N_4288);
and U5078 (N_5078,N_4544,N_3968);
nand U5079 (N_5079,N_4410,N_3730);
and U5080 (N_5080,N_3651,N_3874);
or U5081 (N_5081,N_4425,N_4279);
and U5082 (N_5082,N_4125,N_4672);
or U5083 (N_5083,N_4641,N_3985);
and U5084 (N_5084,N_4103,N_3719);
and U5085 (N_5085,N_4493,N_4763);
and U5086 (N_5086,N_3739,N_3818);
and U5087 (N_5087,N_4280,N_4596);
or U5088 (N_5088,N_4481,N_4734);
xnor U5089 (N_5089,N_3734,N_3764);
nand U5090 (N_5090,N_3722,N_3741);
nor U5091 (N_5091,N_4684,N_3639);
or U5092 (N_5092,N_4482,N_4566);
or U5093 (N_5093,N_3742,N_4712);
xnor U5094 (N_5094,N_4698,N_3780);
nor U5095 (N_5095,N_4131,N_4059);
nand U5096 (N_5096,N_4634,N_4602);
xnor U5097 (N_5097,N_3792,N_3820);
or U5098 (N_5098,N_4789,N_3733);
nand U5099 (N_5099,N_3909,N_4111);
xnor U5100 (N_5100,N_4652,N_4038);
or U5101 (N_5101,N_4302,N_4379);
or U5102 (N_5102,N_4066,N_4011);
nor U5103 (N_5103,N_4770,N_4585);
nand U5104 (N_5104,N_3929,N_4075);
and U5105 (N_5105,N_3859,N_4665);
and U5106 (N_5106,N_4053,N_3619);
xor U5107 (N_5107,N_4007,N_4242);
nand U5108 (N_5108,N_3778,N_4386);
nand U5109 (N_5109,N_4529,N_4400);
or U5110 (N_5110,N_4761,N_4208);
and U5111 (N_5111,N_4605,N_3987);
nand U5112 (N_5112,N_4513,N_4340);
xnor U5113 (N_5113,N_4274,N_3911);
nand U5114 (N_5114,N_3782,N_4326);
or U5115 (N_5115,N_4613,N_4608);
or U5116 (N_5116,N_4590,N_4031);
or U5117 (N_5117,N_3894,N_4203);
xor U5118 (N_5118,N_4534,N_4247);
or U5119 (N_5119,N_3613,N_4225);
and U5120 (N_5120,N_4578,N_4682);
or U5121 (N_5121,N_4256,N_4164);
xnor U5122 (N_5122,N_4551,N_4218);
and U5123 (N_5123,N_4706,N_4681);
and U5124 (N_5124,N_3796,N_4648);
xor U5125 (N_5125,N_3970,N_3835);
or U5126 (N_5126,N_4319,N_4683);
or U5127 (N_5127,N_4458,N_4762);
nand U5128 (N_5128,N_4226,N_4200);
and U5129 (N_5129,N_4303,N_4115);
nand U5130 (N_5130,N_3918,N_4550);
nor U5131 (N_5131,N_4758,N_4253);
nor U5132 (N_5132,N_4352,N_3605);
nand U5133 (N_5133,N_4160,N_4035);
and U5134 (N_5134,N_4507,N_4070);
xnor U5135 (N_5135,N_4693,N_3710);
nor U5136 (N_5136,N_4078,N_4157);
xor U5137 (N_5137,N_4013,N_4238);
nor U5138 (N_5138,N_4021,N_4678);
and U5139 (N_5139,N_4077,N_3752);
xnor U5140 (N_5140,N_3727,N_4444);
nor U5141 (N_5141,N_3898,N_3800);
or U5142 (N_5142,N_4653,N_3882);
nor U5143 (N_5143,N_4076,N_4739);
xnor U5144 (N_5144,N_4679,N_4126);
and U5145 (N_5145,N_4799,N_4788);
nand U5146 (N_5146,N_4361,N_4440);
nor U5147 (N_5147,N_4083,N_4638);
nand U5148 (N_5148,N_4339,N_3704);
nor U5149 (N_5149,N_3743,N_4272);
or U5150 (N_5150,N_3606,N_4252);
xor U5151 (N_5151,N_3707,N_3648);
xnor U5152 (N_5152,N_4141,N_4558);
nor U5153 (N_5153,N_4647,N_3607);
or U5154 (N_5154,N_4454,N_4772);
or U5155 (N_5155,N_3920,N_4177);
or U5156 (N_5156,N_4750,N_4397);
and U5157 (N_5157,N_4373,N_4246);
nor U5158 (N_5158,N_4623,N_3943);
or U5159 (N_5159,N_4332,N_3930);
xor U5160 (N_5160,N_4364,N_3998);
xor U5161 (N_5161,N_3602,N_4382);
xnor U5162 (N_5162,N_4139,N_3737);
and U5163 (N_5163,N_4755,N_4122);
nand U5164 (N_5164,N_4580,N_4270);
nor U5165 (N_5165,N_3669,N_4461);
nand U5166 (N_5166,N_4518,N_4661);
xnor U5167 (N_5167,N_4650,N_4307);
nand U5168 (N_5168,N_4132,N_3904);
or U5169 (N_5169,N_4037,N_4759);
nand U5170 (N_5170,N_3995,N_4443);
nand U5171 (N_5171,N_4110,N_4760);
nand U5172 (N_5172,N_4756,N_4106);
and U5173 (N_5173,N_3622,N_3612);
and U5174 (N_5174,N_4685,N_3817);
or U5175 (N_5175,N_4182,N_4431);
nor U5176 (N_5176,N_4594,N_4276);
nor U5177 (N_5177,N_4676,N_4611);
xnor U5178 (N_5178,N_4677,N_4729);
nand U5179 (N_5179,N_3807,N_3935);
and U5180 (N_5180,N_3641,N_4552);
nand U5181 (N_5181,N_4342,N_3774);
or U5182 (N_5182,N_3993,N_4722);
nor U5183 (N_5183,N_3731,N_4331);
nand U5184 (N_5184,N_4136,N_4646);
xnor U5185 (N_5185,N_4328,N_3975);
or U5186 (N_5186,N_4129,N_3831);
nand U5187 (N_5187,N_4029,N_4105);
and U5188 (N_5188,N_4501,N_3878);
or U5189 (N_5189,N_4158,N_3856);
and U5190 (N_5190,N_3601,N_4176);
xnor U5191 (N_5191,N_4568,N_3656);
nor U5192 (N_5192,N_4369,N_4787);
nand U5193 (N_5193,N_3647,N_3950);
and U5194 (N_5194,N_4530,N_3876);
or U5195 (N_5195,N_4192,N_4098);
nand U5196 (N_5196,N_4790,N_4405);
nand U5197 (N_5197,N_4588,N_4134);
nand U5198 (N_5198,N_4002,N_4639);
nand U5199 (N_5199,N_4152,N_4241);
nand U5200 (N_5200,N_4114,N_3881);
nand U5201 (N_5201,N_3857,N_3816);
nor U5202 (N_5202,N_4265,N_4216);
nor U5203 (N_5203,N_3988,N_4731);
nor U5204 (N_5204,N_3753,N_3765);
and U5205 (N_5205,N_4172,N_4095);
xnor U5206 (N_5206,N_4113,N_4567);
or U5207 (N_5207,N_3692,N_4701);
or U5208 (N_5208,N_3916,N_4227);
xnor U5209 (N_5209,N_3979,N_4740);
nor U5210 (N_5210,N_4505,N_4451);
and U5211 (N_5211,N_4001,N_3967);
or U5212 (N_5212,N_4197,N_4415);
or U5213 (N_5213,N_3643,N_4499);
nand U5214 (N_5214,N_3907,N_4145);
or U5215 (N_5215,N_4268,N_4487);
nand U5216 (N_5216,N_4065,N_3803);
and U5217 (N_5217,N_4654,N_3917);
nor U5218 (N_5218,N_3981,N_3875);
xor U5219 (N_5219,N_4271,N_3693);
or U5220 (N_5220,N_4660,N_4587);
nor U5221 (N_5221,N_4257,N_3932);
xnor U5222 (N_5222,N_4107,N_4718);
and U5223 (N_5223,N_4000,N_4234);
xnor U5224 (N_5224,N_3893,N_3631);
nor U5225 (N_5225,N_4210,N_3922);
or U5226 (N_5226,N_3726,N_3630);
nand U5227 (N_5227,N_3826,N_4178);
or U5228 (N_5228,N_4524,N_4554);
or U5229 (N_5229,N_4027,N_3814);
xor U5230 (N_5230,N_3756,N_3725);
and U5231 (N_5231,N_4781,N_3896);
nor U5232 (N_5232,N_4723,N_4091);
xor U5233 (N_5233,N_4539,N_4153);
nor U5234 (N_5234,N_3762,N_4317);
nand U5235 (N_5235,N_3991,N_4675);
nand U5236 (N_5236,N_4395,N_3959);
or U5237 (N_5237,N_4121,N_3729);
and U5238 (N_5238,N_4778,N_4632);
or U5239 (N_5239,N_4019,N_3705);
xor U5240 (N_5240,N_4629,N_4446);
and U5241 (N_5241,N_4073,N_4163);
or U5242 (N_5242,N_4064,N_3913);
and U5243 (N_5243,N_3766,N_3847);
and U5244 (N_5244,N_4309,N_4350);
nand U5245 (N_5245,N_4776,N_4104);
or U5246 (N_5246,N_3617,N_4635);
nand U5247 (N_5247,N_3892,N_4764);
nand U5248 (N_5248,N_4311,N_4264);
and U5249 (N_5249,N_3604,N_3858);
or U5250 (N_5250,N_4375,N_4389);
nand U5251 (N_5251,N_3790,N_4527);
nor U5252 (N_5252,N_4196,N_4102);
nand U5253 (N_5253,N_4494,N_4149);
or U5254 (N_5254,N_4798,N_4754);
nand U5255 (N_5255,N_3919,N_4796);
xor U5256 (N_5256,N_3644,N_4215);
or U5257 (N_5257,N_4285,N_4786);
nor U5258 (N_5258,N_4640,N_3864);
nor U5259 (N_5259,N_4371,N_4348);
nor U5260 (N_5260,N_3832,N_4607);
xor U5261 (N_5261,N_3972,N_4336);
xnor U5262 (N_5262,N_4144,N_3718);
xor U5263 (N_5263,N_4357,N_4473);
and U5264 (N_5264,N_4466,N_4068);
and U5265 (N_5265,N_3793,N_4773);
xor U5266 (N_5266,N_3977,N_4732);
nand U5267 (N_5267,N_3787,N_4689);
xor U5268 (N_5268,N_4422,N_4746);
nand U5269 (N_5269,N_3776,N_4402);
nor U5270 (N_5270,N_4284,N_3884);
xor U5271 (N_5271,N_4439,N_4480);
and U5272 (N_5272,N_3626,N_4549);
and U5273 (N_5273,N_4018,N_4708);
or U5274 (N_5274,N_4052,N_3844);
xor U5275 (N_5275,N_4069,N_3769);
nor U5276 (N_5276,N_4797,N_4465);
nand U5277 (N_5277,N_4049,N_4612);
or U5278 (N_5278,N_4423,N_4123);
nor U5279 (N_5279,N_4155,N_3877);
nor U5280 (N_5280,N_3680,N_3732);
nand U5281 (N_5281,N_3905,N_4351);
nor U5282 (N_5282,N_4726,N_4519);
nor U5283 (N_5283,N_3691,N_4335);
nor U5284 (N_5284,N_3685,N_4041);
nor U5285 (N_5285,N_3676,N_3712);
xnor U5286 (N_5286,N_3805,N_4570);
nor U5287 (N_5287,N_4769,N_3984);
or U5288 (N_5288,N_4609,N_4498);
nor U5289 (N_5289,N_3614,N_3667);
or U5290 (N_5290,N_4495,N_4512);
xnor U5291 (N_5291,N_4413,N_3825);
nor U5292 (N_5292,N_4347,N_3786);
xor U5293 (N_5293,N_3821,N_4223);
and U5294 (N_5294,N_3955,N_4194);
or U5295 (N_5295,N_4526,N_3740);
and U5296 (N_5296,N_4783,N_3660);
or U5297 (N_5297,N_3770,N_4564);
nor U5298 (N_5298,N_3925,N_3840);
nand U5299 (N_5299,N_4295,N_3889);
nand U5300 (N_5300,N_3999,N_3838);
or U5301 (N_5301,N_3936,N_4619);
xnor U5302 (N_5302,N_4792,N_3697);
nor U5303 (N_5303,N_4063,N_4050);
nor U5304 (N_5304,N_4322,N_3990);
xor U5305 (N_5305,N_4025,N_4517);
and U5306 (N_5306,N_4359,N_4278);
or U5307 (N_5307,N_4649,N_3690);
xor U5308 (N_5308,N_4300,N_4385);
or U5309 (N_5309,N_3953,N_4220);
nor U5310 (N_5310,N_3843,N_4026);
xnor U5311 (N_5311,N_4030,N_3665);
xor U5312 (N_5312,N_4651,N_4054);
xor U5313 (N_5313,N_4087,N_3662);
nor U5314 (N_5314,N_3833,N_4658);
or U5315 (N_5315,N_3992,N_3678);
or U5316 (N_5316,N_4704,N_4774);
or U5317 (N_5317,N_3759,N_4391);
xor U5318 (N_5318,N_4515,N_3912);
and U5319 (N_5319,N_3853,N_4765);
and U5320 (N_5320,N_4573,N_4779);
and U5321 (N_5321,N_4217,N_4291);
nand U5322 (N_5322,N_3965,N_4360);
xor U5323 (N_5323,N_4548,N_4043);
xnor U5324 (N_5324,N_3819,N_3645);
nor U5325 (N_5325,N_4547,N_4680);
and U5326 (N_5326,N_4377,N_3854);
xnor U5327 (N_5327,N_4438,N_4315);
and U5328 (N_5328,N_3716,N_3895);
nor U5329 (N_5329,N_3806,N_4261);
nand U5330 (N_5330,N_3868,N_3872);
or U5331 (N_5331,N_4553,N_4412);
or U5332 (N_5332,N_4545,N_4628);
or U5333 (N_5333,N_4071,N_4039);
or U5334 (N_5334,N_4557,N_4372);
nand U5335 (N_5335,N_4366,N_4713);
or U5336 (N_5336,N_4130,N_4338);
nand U5337 (N_5337,N_4606,N_3891);
xnor U5338 (N_5338,N_4010,N_4467);
or U5339 (N_5339,N_4393,N_4516);
and U5340 (N_5340,N_4521,N_4667);
and U5341 (N_5341,N_4791,N_4504);
nor U5342 (N_5342,N_4277,N_3994);
nor U5343 (N_5343,N_4259,N_4453);
xor U5344 (N_5344,N_3675,N_4093);
and U5345 (N_5345,N_4151,N_4727);
or U5346 (N_5346,N_4541,N_4112);
and U5347 (N_5347,N_3823,N_4060);
nor U5348 (N_5348,N_3928,N_3637);
or U5349 (N_5349,N_3673,N_4296);
xnor U5350 (N_5350,N_4433,N_3879);
nor U5351 (N_5351,N_4476,N_3681);
or U5352 (N_5352,N_4615,N_4502);
xnor U5353 (N_5353,N_4249,N_4475);
or U5354 (N_5354,N_3713,N_4135);
xnor U5355 (N_5355,N_4337,N_4205);
nor U5356 (N_5356,N_3910,N_4452);
nand U5357 (N_5357,N_4388,N_3758);
and U5358 (N_5358,N_4045,N_4305);
nor U5359 (N_5359,N_4079,N_3976);
and U5360 (N_5360,N_3779,N_4565);
or U5361 (N_5361,N_3767,N_3728);
or U5362 (N_5362,N_3755,N_4500);
and U5363 (N_5363,N_4472,N_4503);
nand U5364 (N_5364,N_4191,N_4794);
nand U5365 (N_5365,N_4621,N_4293);
and U5366 (N_5366,N_4211,N_4207);
nand U5367 (N_5367,N_3634,N_3885);
nor U5368 (N_5368,N_3757,N_4430);
nor U5369 (N_5369,N_4244,N_4766);
and U5370 (N_5370,N_4117,N_4325);
or U5371 (N_5371,N_4012,N_3788);
nand U5372 (N_5372,N_4510,N_4119);
xor U5373 (N_5373,N_4199,N_4390);
nor U5374 (N_5374,N_4096,N_4560);
and U5375 (N_5375,N_4455,N_3654);
and U5376 (N_5376,N_4248,N_4169);
nand U5377 (N_5377,N_4716,N_4283);
nor U5378 (N_5378,N_4228,N_3708);
or U5379 (N_5379,N_4576,N_3827);
xor U5380 (N_5380,N_4411,N_3702);
nand U5381 (N_5381,N_3688,N_4230);
xor U5382 (N_5382,N_4308,N_3699);
and U5383 (N_5383,N_4419,N_4464);
or U5384 (N_5384,N_3653,N_4090);
or U5385 (N_5385,N_4312,N_3934);
and U5386 (N_5386,N_4720,N_4542);
xnor U5387 (N_5387,N_3682,N_4100);
nand U5388 (N_5388,N_3783,N_4085);
and U5389 (N_5389,N_4048,N_3813);
or U5390 (N_5390,N_4626,N_3633);
nand U5391 (N_5391,N_4637,N_3983);
nand U5392 (N_5392,N_3747,N_3812);
and U5393 (N_5393,N_3711,N_3862);
and U5394 (N_5394,N_3768,N_3908);
or U5395 (N_5395,N_3804,N_4318);
and U5396 (N_5396,N_4392,N_4470);
and U5397 (N_5397,N_3760,N_4525);
nand U5398 (N_5398,N_4138,N_4224);
or U5399 (N_5399,N_4354,N_3671);
and U5400 (N_5400,N_3622,N_4516);
nand U5401 (N_5401,N_3958,N_4472);
nand U5402 (N_5402,N_4302,N_3738);
or U5403 (N_5403,N_3600,N_4038);
nand U5404 (N_5404,N_4457,N_4230);
or U5405 (N_5405,N_4649,N_4609);
xnor U5406 (N_5406,N_3859,N_4208);
xor U5407 (N_5407,N_4001,N_4534);
or U5408 (N_5408,N_4059,N_4577);
and U5409 (N_5409,N_4372,N_4325);
or U5410 (N_5410,N_4711,N_4071);
xnor U5411 (N_5411,N_4173,N_4400);
nor U5412 (N_5412,N_4441,N_4557);
or U5413 (N_5413,N_3672,N_4118);
xor U5414 (N_5414,N_3830,N_3812);
nor U5415 (N_5415,N_4030,N_4754);
xnor U5416 (N_5416,N_4606,N_4683);
or U5417 (N_5417,N_4706,N_4756);
nor U5418 (N_5418,N_4594,N_3920);
xnor U5419 (N_5419,N_4161,N_4406);
nand U5420 (N_5420,N_3640,N_4237);
and U5421 (N_5421,N_4329,N_4504);
nor U5422 (N_5422,N_3824,N_3621);
xnor U5423 (N_5423,N_3682,N_4231);
xnor U5424 (N_5424,N_4423,N_3823);
or U5425 (N_5425,N_4716,N_4155);
nand U5426 (N_5426,N_4591,N_4124);
or U5427 (N_5427,N_4663,N_4456);
xor U5428 (N_5428,N_4398,N_3841);
or U5429 (N_5429,N_3693,N_3663);
nand U5430 (N_5430,N_4785,N_3616);
nand U5431 (N_5431,N_3745,N_4254);
or U5432 (N_5432,N_3609,N_4043);
xnor U5433 (N_5433,N_3732,N_4396);
xnor U5434 (N_5434,N_3753,N_3744);
xor U5435 (N_5435,N_4039,N_4316);
nor U5436 (N_5436,N_4253,N_4246);
and U5437 (N_5437,N_4758,N_3856);
nor U5438 (N_5438,N_4523,N_3642);
nor U5439 (N_5439,N_4107,N_3849);
nand U5440 (N_5440,N_4508,N_4477);
nor U5441 (N_5441,N_4232,N_3775);
nand U5442 (N_5442,N_4761,N_4400);
xor U5443 (N_5443,N_3894,N_3669);
or U5444 (N_5444,N_4093,N_4705);
or U5445 (N_5445,N_4157,N_4319);
nor U5446 (N_5446,N_4364,N_3830);
nand U5447 (N_5447,N_4348,N_4285);
nand U5448 (N_5448,N_4401,N_4503);
nor U5449 (N_5449,N_4110,N_3822);
and U5450 (N_5450,N_4501,N_4776);
xnor U5451 (N_5451,N_4407,N_4099);
nand U5452 (N_5452,N_4021,N_4579);
nor U5453 (N_5453,N_4007,N_3657);
nor U5454 (N_5454,N_3894,N_4303);
and U5455 (N_5455,N_4139,N_4760);
nor U5456 (N_5456,N_3857,N_4625);
nand U5457 (N_5457,N_3732,N_4430);
xnor U5458 (N_5458,N_4112,N_3786);
and U5459 (N_5459,N_4295,N_4277);
nand U5460 (N_5460,N_4590,N_4193);
nand U5461 (N_5461,N_3984,N_4441);
or U5462 (N_5462,N_4281,N_4465);
nor U5463 (N_5463,N_3658,N_3951);
nand U5464 (N_5464,N_4725,N_4068);
nor U5465 (N_5465,N_4314,N_3602);
and U5466 (N_5466,N_4443,N_4278);
nand U5467 (N_5467,N_3758,N_3673);
nor U5468 (N_5468,N_4555,N_4068);
xor U5469 (N_5469,N_4574,N_4348);
xnor U5470 (N_5470,N_4344,N_4183);
nor U5471 (N_5471,N_3833,N_3962);
nand U5472 (N_5472,N_4463,N_4512);
nor U5473 (N_5473,N_4551,N_4293);
nor U5474 (N_5474,N_3615,N_3717);
and U5475 (N_5475,N_4503,N_4257);
and U5476 (N_5476,N_3720,N_4587);
nand U5477 (N_5477,N_3881,N_4580);
or U5478 (N_5478,N_3657,N_4548);
xnor U5479 (N_5479,N_3884,N_3851);
or U5480 (N_5480,N_4682,N_3812);
nand U5481 (N_5481,N_4077,N_3709);
nor U5482 (N_5482,N_4499,N_4274);
or U5483 (N_5483,N_4112,N_3795);
nand U5484 (N_5484,N_4635,N_3926);
nand U5485 (N_5485,N_3964,N_4374);
nor U5486 (N_5486,N_4482,N_3937);
nand U5487 (N_5487,N_3883,N_3671);
nand U5488 (N_5488,N_4242,N_4213);
and U5489 (N_5489,N_4516,N_4705);
and U5490 (N_5490,N_3796,N_3959);
and U5491 (N_5491,N_4380,N_3665);
and U5492 (N_5492,N_4512,N_3837);
or U5493 (N_5493,N_3743,N_4379);
or U5494 (N_5494,N_4248,N_4382);
nand U5495 (N_5495,N_3868,N_3983);
xor U5496 (N_5496,N_4424,N_4388);
and U5497 (N_5497,N_4056,N_3917);
and U5498 (N_5498,N_4085,N_4245);
nand U5499 (N_5499,N_4165,N_3679);
nor U5500 (N_5500,N_4699,N_4123);
nor U5501 (N_5501,N_4555,N_4702);
nand U5502 (N_5502,N_4219,N_3638);
xnor U5503 (N_5503,N_3908,N_4750);
nand U5504 (N_5504,N_3660,N_3746);
nand U5505 (N_5505,N_4282,N_4271);
xnor U5506 (N_5506,N_4020,N_4529);
xnor U5507 (N_5507,N_4663,N_4453);
or U5508 (N_5508,N_4012,N_4570);
xnor U5509 (N_5509,N_4549,N_3694);
or U5510 (N_5510,N_3941,N_4563);
nor U5511 (N_5511,N_4424,N_3833);
or U5512 (N_5512,N_4341,N_3740);
xnor U5513 (N_5513,N_4475,N_4639);
or U5514 (N_5514,N_4136,N_4160);
nor U5515 (N_5515,N_4116,N_4547);
or U5516 (N_5516,N_4301,N_4106);
and U5517 (N_5517,N_4777,N_4058);
xor U5518 (N_5518,N_4391,N_4709);
nor U5519 (N_5519,N_4777,N_3673);
xnor U5520 (N_5520,N_3875,N_4653);
nand U5521 (N_5521,N_3617,N_3731);
nand U5522 (N_5522,N_4149,N_4124);
xnor U5523 (N_5523,N_4665,N_4011);
nand U5524 (N_5524,N_3861,N_4439);
nand U5525 (N_5525,N_4773,N_4659);
nor U5526 (N_5526,N_4323,N_4411);
and U5527 (N_5527,N_4797,N_3814);
xnor U5528 (N_5528,N_4067,N_4039);
nand U5529 (N_5529,N_4753,N_4587);
xor U5530 (N_5530,N_3626,N_3624);
nor U5531 (N_5531,N_4632,N_4690);
and U5532 (N_5532,N_4486,N_4106);
or U5533 (N_5533,N_3641,N_4140);
or U5534 (N_5534,N_4341,N_3819);
nand U5535 (N_5535,N_4466,N_4528);
and U5536 (N_5536,N_4139,N_4119);
and U5537 (N_5537,N_4251,N_3787);
or U5538 (N_5538,N_3806,N_4565);
xnor U5539 (N_5539,N_4059,N_4588);
nor U5540 (N_5540,N_4763,N_3665);
nand U5541 (N_5541,N_3825,N_4426);
nand U5542 (N_5542,N_4007,N_4093);
or U5543 (N_5543,N_4313,N_3690);
nor U5544 (N_5544,N_4096,N_4555);
xor U5545 (N_5545,N_3714,N_4704);
nand U5546 (N_5546,N_4091,N_3617);
xnor U5547 (N_5547,N_4578,N_3779);
xor U5548 (N_5548,N_4739,N_3958);
and U5549 (N_5549,N_4651,N_4613);
xor U5550 (N_5550,N_4486,N_3886);
nand U5551 (N_5551,N_4391,N_4518);
nand U5552 (N_5552,N_4617,N_4603);
or U5553 (N_5553,N_4126,N_3823);
and U5554 (N_5554,N_3731,N_3957);
nand U5555 (N_5555,N_3644,N_4036);
nor U5556 (N_5556,N_3713,N_3799);
and U5557 (N_5557,N_3727,N_4529);
nand U5558 (N_5558,N_4725,N_3610);
or U5559 (N_5559,N_4215,N_3908);
or U5560 (N_5560,N_4609,N_3874);
xnor U5561 (N_5561,N_4320,N_3727);
nand U5562 (N_5562,N_3627,N_4694);
and U5563 (N_5563,N_3675,N_4275);
or U5564 (N_5564,N_4795,N_4474);
xnor U5565 (N_5565,N_3671,N_3687);
and U5566 (N_5566,N_4633,N_4776);
or U5567 (N_5567,N_4239,N_4236);
nor U5568 (N_5568,N_4000,N_4615);
and U5569 (N_5569,N_4317,N_4161);
or U5570 (N_5570,N_4662,N_4174);
or U5571 (N_5571,N_4645,N_3630);
nor U5572 (N_5572,N_3999,N_3855);
nand U5573 (N_5573,N_4624,N_4512);
nor U5574 (N_5574,N_3894,N_4606);
nand U5575 (N_5575,N_3696,N_3715);
nor U5576 (N_5576,N_4079,N_4226);
nor U5577 (N_5577,N_4203,N_3855);
and U5578 (N_5578,N_4360,N_4107);
and U5579 (N_5579,N_4396,N_3642);
nor U5580 (N_5580,N_4523,N_4104);
nor U5581 (N_5581,N_3966,N_3889);
nand U5582 (N_5582,N_3630,N_3954);
xor U5583 (N_5583,N_4084,N_3700);
or U5584 (N_5584,N_4749,N_3606);
nor U5585 (N_5585,N_4649,N_3754);
or U5586 (N_5586,N_4527,N_4469);
xnor U5587 (N_5587,N_4154,N_4326);
and U5588 (N_5588,N_4424,N_4764);
and U5589 (N_5589,N_4713,N_4179);
xnor U5590 (N_5590,N_4041,N_4543);
or U5591 (N_5591,N_4750,N_3645);
and U5592 (N_5592,N_3757,N_4364);
xor U5593 (N_5593,N_3728,N_4763);
nand U5594 (N_5594,N_3895,N_4487);
xor U5595 (N_5595,N_3676,N_3884);
nand U5596 (N_5596,N_3976,N_4570);
and U5597 (N_5597,N_4618,N_4467);
nand U5598 (N_5598,N_4168,N_4502);
nor U5599 (N_5599,N_4316,N_4406);
xnor U5600 (N_5600,N_4408,N_4335);
and U5601 (N_5601,N_3622,N_3994);
xnor U5602 (N_5602,N_4779,N_4061);
nor U5603 (N_5603,N_4324,N_4090);
or U5604 (N_5604,N_4204,N_4364);
or U5605 (N_5605,N_4459,N_4180);
nor U5606 (N_5606,N_3635,N_4079);
or U5607 (N_5607,N_4560,N_3953);
or U5608 (N_5608,N_4647,N_4039);
xnor U5609 (N_5609,N_4128,N_4320);
nand U5610 (N_5610,N_3996,N_4296);
nand U5611 (N_5611,N_4034,N_4202);
xnor U5612 (N_5612,N_4535,N_3676);
nor U5613 (N_5613,N_4347,N_4631);
or U5614 (N_5614,N_4541,N_3721);
nor U5615 (N_5615,N_4241,N_4763);
xnor U5616 (N_5616,N_4211,N_4296);
or U5617 (N_5617,N_4796,N_4116);
nor U5618 (N_5618,N_4705,N_4461);
or U5619 (N_5619,N_4648,N_3774);
nand U5620 (N_5620,N_4183,N_3735);
nor U5621 (N_5621,N_4124,N_4209);
xor U5622 (N_5622,N_3992,N_4665);
xor U5623 (N_5623,N_3751,N_3985);
or U5624 (N_5624,N_3880,N_4220);
or U5625 (N_5625,N_3612,N_4562);
nor U5626 (N_5626,N_3766,N_4176);
and U5627 (N_5627,N_3806,N_4641);
xnor U5628 (N_5628,N_4468,N_3720);
or U5629 (N_5629,N_4410,N_4645);
xor U5630 (N_5630,N_3979,N_4132);
and U5631 (N_5631,N_4564,N_4705);
nor U5632 (N_5632,N_3924,N_4626);
nor U5633 (N_5633,N_3962,N_3907);
and U5634 (N_5634,N_4130,N_4094);
xor U5635 (N_5635,N_3770,N_4011);
xor U5636 (N_5636,N_3817,N_4735);
or U5637 (N_5637,N_3985,N_3620);
or U5638 (N_5638,N_4567,N_4255);
or U5639 (N_5639,N_4205,N_4577);
xnor U5640 (N_5640,N_4198,N_3622);
and U5641 (N_5641,N_4025,N_4015);
nand U5642 (N_5642,N_3828,N_4495);
or U5643 (N_5643,N_3873,N_3803);
and U5644 (N_5644,N_3650,N_4124);
and U5645 (N_5645,N_4163,N_4482);
nor U5646 (N_5646,N_3820,N_3614);
and U5647 (N_5647,N_4337,N_4094);
nor U5648 (N_5648,N_3672,N_4464);
or U5649 (N_5649,N_4434,N_4344);
and U5650 (N_5650,N_4048,N_4410);
or U5651 (N_5651,N_4234,N_3966);
or U5652 (N_5652,N_4121,N_4104);
xor U5653 (N_5653,N_4585,N_3632);
and U5654 (N_5654,N_4282,N_4537);
nand U5655 (N_5655,N_4221,N_4654);
and U5656 (N_5656,N_4448,N_3686);
nand U5657 (N_5657,N_4408,N_3801);
and U5658 (N_5658,N_4433,N_4725);
nor U5659 (N_5659,N_4520,N_3627);
nor U5660 (N_5660,N_4318,N_4228);
nand U5661 (N_5661,N_4069,N_4376);
nand U5662 (N_5662,N_4590,N_4068);
xnor U5663 (N_5663,N_3948,N_4069);
and U5664 (N_5664,N_4166,N_3992);
or U5665 (N_5665,N_4190,N_3977);
nand U5666 (N_5666,N_4451,N_4788);
xnor U5667 (N_5667,N_3856,N_4358);
nand U5668 (N_5668,N_3656,N_4137);
xor U5669 (N_5669,N_4404,N_4394);
nor U5670 (N_5670,N_4328,N_4470);
xnor U5671 (N_5671,N_3724,N_4503);
xnor U5672 (N_5672,N_4179,N_3673);
xor U5673 (N_5673,N_3857,N_4611);
xnor U5674 (N_5674,N_4581,N_4288);
and U5675 (N_5675,N_3712,N_3822);
and U5676 (N_5676,N_3741,N_4041);
or U5677 (N_5677,N_3926,N_4630);
xnor U5678 (N_5678,N_4722,N_4050);
or U5679 (N_5679,N_3668,N_4108);
or U5680 (N_5680,N_4000,N_3949);
or U5681 (N_5681,N_4315,N_3775);
or U5682 (N_5682,N_4093,N_4573);
and U5683 (N_5683,N_4019,N_4472);
nor U5684 (N_5684,N_4288,N_3859);
nor U5685 (N_5685,N_4247,N_3723);
or U5686 (N_5686,N_3765,N_4313);
nor U5687 (N_5687,N_3872,N_4706);
or U5688 (N_5688,N_4558,N_3990);
xor U5689 (N_5689,N_3763,N_3765);
and U5690 (N_5690,N_3628,N_3709);
xor U5691 (N_5691,N_4637,N_3634);
or U5692 (N_5692,N_3974,N_4553);
nor U5693 (N_5693,N_3657,N_4117);
xor U5694 (N_5694,N_4119,N_3932);
or U5695 (N_5695,N_3626,N_4314);
nand U5696 (N_5696,N_4209,N_3794);
or U5697 (N_5697,N_4121,N_4285);
or U5698 (N_5698,N_4735,N_3930);
or U5699 (N_5699,N_4190,N_3748);
nand U5700 (N_5700,N_3704,N_4757);
nor U5701 (N_5701,N_4362,N_4798);
and U5702 (N_5702,N_4432,N_3916);
xor U5703 (N_5703,N_4542,N_3819);
nor U5704 (N_5704,N_3987,N_4563);
nand U5705 (N_5705,N_4652,N_4485);
or U5706 (N_5706,N_4386,N_4437);
nand U5707 (N_5707,N_4375,N_4784);
or U5708 (N_5708,N_4606,N_4179);
nor U5709 (N_5709,N_3876,N_4125);
nor U5710 (N_5710,N_4092,N_3918);
or U5711 (N_5711,N_3900,N_4415);
or U5712 (N_5712,N_4505,N_4308);
xnor U5713 (N_5713,N_3712,N_3886);
or U5714 (N_5714,N_4334,N_4290);
nand U5715 (N_5715,N_3727,N_3626);
and U5716 (N_5716,N_4643,N_4792);
nand U5717 (N_5717,N_4211,N_3754);
xor U5718 (N_5718,N_4498,N_3785);
xor U5719 (N_5719,N_4337,N_4537);
xor U5720 (N_5720,N_4680,N_4127);
xnor U5721 (N_5721,N_4239,N_4793);
nor U5722 (N_5722,N_4653,N_3842);
or U5723 (N_5723,N_4646,N_4757);
or U5724 (N_5724,N_4524,N_3884);
xnor U5725 (N_5725,N_4493,N_3672);
or U5726 (N_5726,N_4700,N_4246);
and U5727 (N_5727,N_4467,N_4056);
or U5728 (N_5728,N_3747,N_4712);
xnor U5729 (N_5729,N_3626,N_4028);
nor U5730 (N_5730,N_4078,N_4740);
or U5731 (N_5731,N_4481,N_4066);
or U5732 (N_5732,N_4647,N_4643);
nor U5733 (N_5733,N_4312,N_4783);
xnor U5734 (N_5734,N_4321,N_4663);
nor U5735 (N_5735,N_4777,N_3878);
nand U5736 (N_5736,N_4172,N_3616);
nor U5737 (N_5737,N_4721,N_4274);
and U5738 (N_5738,N_4481,N_3767);
nand U5739 (N_5739,N_3807,N_3964);
nand U5740 (N_5740,N_4510,N_4118);
nand U5741 (N_5741,N_4612,N_4796);
and U5742 (N_5742,N_4001,N_4283);
nand U5743 (N_5743,N_3913,N_4517);
or U5744 (N_5744,N_4379,N_4308);
and U5745 (N_5745,N_3964,N_4021);
xor U5746 (N_5746,N_3772,N_3734);
nor U5747 (N_5747,N_3946,N_4238);
or U5748 (N_5748,N_3724,N_4663);
xnor U5749 (N_5749,N_4106,N_4043);
nand U5750 (N_5750,N_4244,N_4484);
or U5751 (N_5751,N_3846,N_4086);
or U5752 (N_5752,N_4430,N_4273);
xnor U5753 (N_5753,N_4644,N_4583);
nand U5754 (N_5754,N_3778,N_3709);
or U5755 (N_5755,N_4373,N_4776);
or U5756 (N_5756,N_4377,N_3758);
xor U5757 (N_5757,N_4190,N_4464);
and U5758 (N_5758,N_4030,N_4012);
and U5759 (N_5759,N_3834,N_4705);
and U5760 (N_5760,N_3791,N_3722);
and U5761 (N_5761,N_4060,N_4109);
nand U5762 (N_5762,N_4739,N_3929);
nand U5763 (N_5763,N_4511,N_4758);
and U5764 (N_5764,N_4104,N_4135);
nor U5765 (N_5765,N_4674,N_3930);
nand U5766 (N_5766,N_3832,N_3950);
and U5767 (N_5767,N_4057,N_4664);
and U5768 (N_5768,N_3694,N_4208);
or U5769 (N_5769,N_3638,N_4280);
and U5770 (N_5770,N_4379,N_4626);
and U5771 (N_5771,N_4369,N_4593);
nor U5772 (N_5772,N_4325,N_3652);
xor U5773 (N_5773,N_4305,N_4193);
xnor U5774 (N_5774,N_3689,N_4566);
nand U5775 (N_5775,N_4434,N_4573);
nand U5776 (N_5776,N_4785,N_3965);
nand U5777 (N_5777,N_4681,N_4236);
or U5778 (N_5778,N_4320,N_3714);
nor U5779 (N_5779,N_4738,N_4649);
xor U5780 (N_5780,N_4061,N_4134);
or U5781 (N_5781,N_3616,N_4013);
xor U5782 (N_5782,N_3630,N_4796);
nor U5783 (N_5783,N_4460,N_4328);
or U5784 (N_5784,N_4594,N_4417);
or U5785 (N_5785,N_3992,N_3695);
xnor U5786 (N_5786,N_4240,N_4478);
nand U5787 (N_5787,N_4303,N_3676);
nor U5788 (N_5788,N_4505,N_4719);
and U5789 (N_5789,N_3995,N_4401);
nand U5790 (N_5790,N_4448,N_3806);
and U5791 (N_5791,N_4664,N_3842);
xor U5792 (N_5792,N_4303,N_4524);
xor U5793 (N_5793,N_4064,N_4445);
nand U5794 (N_5794,N_4794,N_3721);
nor U5795 (N_5795,N_3708,N_4034);
or U5796 (N_5796,N_3727,N_4263);
and U5797 (N_5797,N_3620,N_4709);
xnor U5798 (N_5798,N_3738,N_4756);
nand U5799 (N_5799,N_4320,N_4583);
or U5800 (N_5800,N_3938,N_3642);
nor U5801 (N_5801,N_4124,N_3662);
and U5802 (N_5802,N_4437,N_4535);
and U5803 (N_5803,N_4332,N_4431);
and U5804 (N_5804,N_4783,N_3953);
xor U5805 (N_5805,N_4054,N_3653);
or U5806 (N_5806,N_4044,N_3699);
and U5807 (N_5807,N_4668,N_3915);
xor U5808 (N_5808,N_4504,N_4736);
and U5809 (N_5809,N_3797,N_4632);
xor U5810 (N_5810,N_4642,N_3793);
and U5811 (N_5811,N_4413,N_4676);
or U5812 (N_5812,N_3636,N_4027);
nand U5813 (N_5813,N_4199,N_4056);
nor U5814 (N_5814,N_4648,N_4645);
nor U5815 (N_5815,N_3784,N_4474);
xnor U5816 (N_5816,N_3965,N_3957);
nor U5817 (N_5817,N_4668,N_4452);
nand U5818 (N_5818,N_4359,N_4772);
nand U5819 (N_5819,N_3682,N_3767);
nand U5820 (N_5820,N_4234,N_4212);
nor U5821 (N_5821,N_4039,N_4499);
xnor U5822 (N_5822,N_4680,N_4271);
and U5823 (N_5823,N_4750,N_3845);
nor U5824 (N_5824,N_4640,N_3734);
xnor U5825 (N_5825,N_4022,N_4707);
and U5826 (N_5826,N_4018,N_4151);
and U5827 (N_5827,N_4439,N_3973);
and U5828 (N_5828,N_3773,N_4103);
nand U5829 (N_5829,N_3784,N_3616);
or U5830 (N_5830,N_3978,N_4600);
xnor U5831 (N_5831,N_4298,N_4196);
and U5832 (N_5832,N_4131,N_3730);
nand U5833 (N_5833,N_3851,N_4108);
nor U5834 (N_5834,N_3609,N_4527);
nor U5835 (N_5835,N_4396,N_4455);
nand U5836 (N_5836,N_4793,N_4010);
nor U5837 (N_5837,N_3889,N_4278);
or U5838 (N_5838,N_3997,N_4219);
or U5839 (N_5839,N_4323,N_4518);
and U5840 (N_5840,N_4551,N_4170);
nor U5841 (N_5841,N_4741,N_3794);
nand U5842 (N_5842,N_4511,N_4009);
and U5843 (N_5843,N_4280,N_4734);
or U5844 (N_5844,N_4288,N_3618);
nor U5845 (N_5845,N_4588,N_4346);
nor U5846 (N_5846,N_3935,N_3852);
or U5847 (N_5847,N_3899,N_3684);
nand U5848 (N_5848,N_4475,N_4665);
and U5849 (N_5849,N_3656,N_4151);
xor U5850 (N_5850,N_4741,N_3814);
nor U5851 (N_5851,N_4463,N_4429);
xnor U5852 (N_5852,N_4669,N_4675);
or U5853 (N_5853,N_4619,N_3741);
nand U5854 (N_5854,N_4088,N_3801);
or U5855 (N_5855,N_4785,N_4201);
nand U5856 (N_5856,N_3971,N_3724);
and U5857 (N_5857,N_4763,N_4338);
and U5858 (N_5858,N_4396,N_4016);
nand U5859 (N_5859,N_4710,N_4084);
nand U5860 (N_5860,N_4486,N_4714);
nand U5861 (N_5861,N_4572,N_4579);
xnor U5862 (N_5862,N_3956,N_3821);
nor U5863 (N_5863,N_4000,N_4372);
nor U5864 (N_5864,N_4067,N_4594);
or U5865 (N_5865,N_4043,N_3943);
nor U5866 (N_5866,N_4561,N_4238);
xnor U5867 (N_5867,N_3998,N_4163);
nand U5868 (N_5868,N_4561,N_4677);
and U5869 (N_5869,N_3799,N_4754);
and U5870 (N_5870,N_4637,N_4319);
xnor U5871 (N_5871,N_3952,N_4418);
xor U5872 (N_5872,N_4175,N_4434);
and U5873 (N_5873,N_4455,N_4413);
nor U5874 (N_5874,N_3692,N_3899);
and U5875 (N_5875,N_4663,N_4223);
and U5876 (N_5876,N_4636,N_4062);
or U5877 (N_5877,N_4687,N_4624);
or U5878 (N_5878,N_4001,N_4459);
nor U5879 (N_5879,N_3908,N_4024);
xnor U5880 (N_5880,N_4513,N_4147);
or U5881 (N_5881,N_4584,N_4520);
xor U5882 (N_5882,N_4385,N_4381);
nand U5883 (N_5883,N_4614,N_4440);
xnor U5884 (N_5884,N_4163,N_4318);
nor U5885 (N_5885,N_4411,N_4024);
nor U5886 (N_5886,N_3624,N_3748);
nor U5887 (N_5887,N_4540,N_4696);
and U5888 (N_5888,N_3664,N_4333);
nand U5889 (N_5889,N_4762,N_3906);
and U5890 (N_5890,N_4471,N_3914);
or U5891 (N_5891,N_3888,N_4314);
nor U5892 (N_5892,N_4786,N_3687);
or U5893 (N_5893,N_4157,N_3637);
or U5894 (N_5894,N_4796,N_4061);
and U5895 (N_5895,N_3985,N_4752);
and U5896 (N_5896,N_4058,N_4050);
nor U5897 (N_5897,N_4318,N_4213);
xnor U5898 (N_5898,N_4437,N_3698);
or U5899 (N_5899,N_4019,N_4757);
nor U5900 (N_5900,N_4658,N_3955);
or U5901 (N_5901,N_3855,N_3993);
nand U5902 (N_5902,N_4361,N_4592);
nor U5903 (N_5903,N_4673,N_4415);
or U5904 (N_5904,N_4304,N_3800);
nand U5905 (N_5905,N_4162,N_4404);
nand U5906 (N_5906,N_4122,N_4137);
and U5907 (N_5907,N_3649,N_4115);
xnor U5908 (N_5908,N_4581,N_3620);
nand U5909 (N_5909,N_4421,N_4478);
nand U5910 (N_5910,N_4292,N_4694);
xnor U5911 (N_5911,N_4233,N_3845);
xor U5912 (N_5912,N_4369,N_3682);
nor U5913 (N_5913,N_4225,N_3625);
xnor U5914 (N_5914,N_4053,N_4158);
nor U5915 (N_5915,N_4002,N_4621);
and U5916 (N_5916,N_3709,N_4775);
and U5917 (N_5917,N_4701,N_3911);
and U5918 (N_5918,N_4514,N_4515);
xor U5919 (N_5919,N_4096,N_4636);
and U5920 (N_5920,N_3865,N_3920);
nor U5921 (N_5921,N_4193,N_3870);
nor U5922 (N_5922,N_4050,N_4222);
and U5923 (N_5923,N_4022,N_4052);
xnor U5924 (N_5924,N_4087,N_4272);
nand U5925 (N_5925,N_4745,N_3706);
and U5926 (N_5926,N_3884,N_3756);
nand U5927 (N_5927,N_4599,N_4203);
nand U5928 (N_5928,N_3610,N_4719);
and U5929 (N_5929,N_3956,N_4476);
xnor U5930 (N_5930,N_4574,N_4139);
nand U5931 (N_5931,N_3933,N_4259);
nand U5932 (N_5932,N_3730,N_4657);
nor U5933 (N_5933,N_3849,N_4644);
xor U5934 (N_5934,N_4621,N_4179);
nand U5935 (N_5935,N_4128,N_3956);
or U5936 (N_5936,N_4620,N_4414);
xnor U5937 (N_5937,N_4381,N_4520);
nand U5938 (N_5938,N_3932,N_3823);
nor U5939 (N_5939,N_3648,N_4154);
xnor U5940 (N_5940,N_4478,N_3976);
and U5941 (N_5941,N_3688,N_4620);
or U5942 (N_5942,N_4173,N_3877);
nand U5943 (N_5943,N_3868,N_4588);
nand U5944 (N_5944,N_4526,N_4416);
nor U5945 (N_5945,N_4341,N_3858);
nand U5946 (N_5946,N_4224,N_3995);
xnor U5947 (N_5947,N_3721,N_4427);
nor U5948 (N_5948,N_4360,N_4003);
and U5949 (N_5949,N_3661,N_3901);
nor U5950 (N_5950,N_4721,N_3752);
nor U5951 (N_5951,N_3682,N_3732);
xnor U5952 (N_5952,N_4482,N_3840);
nand U5953 (N_5953,N_4685,N_3789);
nor U5954 (N_5954,N_4072,N_4607);
and U5955 (N_5955,N_4429,N_3795);
or U5956 (N_5956,N_4385,N_4255);
and U5957 (N_5957,N_4108,N_4081);
nor U5958 (N_5958,N_3815,N_4417);
xnor U5959 (N_5959,N_3843,N_4101);
nor U5960 (N_5960,N_3604,N_4551);
nor U5961 (N_5961,N_4127,N_3889);
nand U5962 (N_5962,N_3636,N_4291);
nand U5963 (N_5963,N_3733,N_3676);
nand U5964 (N_5964,N_4791,N_4347);
nand U5965 (N_5965,N_4390,N_3843);
nor U5966 (N_5966,N_4118,N_3877);
and U5967 (N_5967,N_3908,N_4212);
or U5968 (N_5968,N_4466,N_4579);
or U5969 (N_5969,N_3912,N_4432);
nand U5970 (N_5970,N_4110,N_3718);
or U5971 (N_5971,N_3724,N_4796);
nor U5972 (N_5972,N_4355,N_3629);
nand U5973 (N_5973,N_4496,N_4095);
and U5974 (N_5974,N_3896,N_4770);
nand U5975 (N_5975,N_4331,N_3774);
and U5976 (N_5976,N_4224,N_3628);
nor U5977 (N_5977,N_4294,N_4206);
and U5978 (N_5978,N_4724,N_4436);
or U5979 (N_5979,N_4786,N_4663);
xnor U5980 (N_5980,N_4440,N_4252);
xor U5981 (N_5981,N_3868,N_4349);
or U5982 (N_5982,N_3910,N_4789);
and U5983 (N_5983,N_4759,N_4096);
nor U5984 (N_5984,N_4341,N_3769);
nor U5985 (N_5985,N_3726,N_4260);
or U5986 (N_5986,N_4692,N_4209);
nor U5987 (N_5987,N_4410,N_3926);
or U5988 (N_5988,N_3814,N_4086);
nor U5989 (N_5989,N_4234,N_4487);
and U5990 (N_5990,N_4783,N_3820);
and U5991 (N_5991,N_4691,N_3600);
nor U5992 (N_5992,N_3842,N_4367);
nand U5993 (N_5993,N_4013,N_4039);
nor U5994 (N_5994,N_4298,N_4099);
or U5995 (N_5995,N_4094,N_4310);
nor U5996 (N_5996,N_3650,N_4216);
nand U5997 (N_5997,N_4220,N_3860);
or U5998 (N_5998,N_4718,N_4211);
nor U5999 (N_5999,N_3859,N_4160);
xor U6000 (N_6000,N_5691,N_5169);
xor U6001 (N_6001,N_5493,N_5092);
nor U6002 (N_6002,N_5708,N_5772);
xor U6003 (N_6003,N_5023,N_5693);
nand U6004 (N_6004,N_5378,N_5653);
nor U6005 (N_6005,N_5070,N_5208);
or U6006 (N_6006,N_4906,N_5381);
or U6007 (N_6007,N_5600,N_5610);
xor U6008 (N_6008,N_4990,N_5048);
nand U6009 (N_6009,N_5407,N_5699);
nand U6010 (N_6010,N_5064,N_5826);
nand U6011 (N_6011,N_5509,N_5710);
nand U6012 (N_6012,N_5814,N_5951);
and U6013 (N_6013,N_5686,N_5081);
xor U6014 (N_6014,N_4863,N_5244);
xnor U6015 (N_6015,N_5120,N_4827);
nand U6016 (N_6016,N_5227,N_5611);
nor U6017 (N_6017,N_5884,N_5148);
or U6018 (N_6018,N_5361,N_4851);
nor U6019 (N_6019,N_5957,N_5987);
xnor U6020 (N_6020,N_5088,N_5910);
and U6021 (N_6021,N_5541,N_5272);
xor U6022 (N_6022,N_5179,N_5485);
or U6023 (N_6023,N_5624,N_5923);
or U6024 (N_6024,N_5406,N_5977);
nor U6025 (N_6025,N_4888,N_5968);
nand U6026 (N_6026,N_5477,N_4992);
nand U6027 (N_6027,N_4875,N_5038);
xor U6028 (N_6028,N_4911,N_5303);
nand U6029 (N_6029,N_5906,N_5344);
nand U6030 (N_6030,N_5238,N_5062);
nor U6031 (N_6031,N_5734,N_5770);
xnor U6032 (N_6032,N_5758,N_5841);
and U6033 (N_6033,N_4847,N_5755);
nor U6034 (N_6034,N_5197,N_5199);
and U6035 (N_6035,N_5393,N_5126);
nor U6036 (N_6036,N_5830,N_5265);
or U6037 (N_6037,N_5704,N_5207);
xnor U6038 (N_6038,N_5049,N_5454);
or U6039 (N_6039,N_5270,N_5877);
and U6040 (N_6040,N_5836,N_5616);
nor U6041 (N_6041,N_5763,N_5443);
nor U6042 (N_6042,N_5325,N_5993);
xor U6043 (N_6043,N_5964,N_4874);
xnor U6044 (N_6044,N_4948,N_5803);
nor U6045 (N_6045,N_4993,N_5740);
or U6046 (N_6046,N_4935,N_5479);
or U6047 (N_6047,N_5465,N_5472);
nor U6048 (N_6048,N_5625,N_5421);
nor U6049 (N_6049,N_5480,N_5404);
or U6050 (N_6050,N_4933,N_5398);
xnor U6051 (N_6051,N_5347,N_4833);
and U6052 (N_6052,N_4811,N_5895);
xor U6053 (N_6053,N_5522,N_5683);
xor U6054 (N_6054,N_4969,N_5969);
and U6055 (N_6055,N_5562,N_4867);
nand U6056 (N_6056,N_5947,N_4994);
or U6057 (N_6057,N_5596,N_4858);
xor U6058 (N_6058,N_5688,N_5333);
nand U6059 (N_6059,N_5310,N_5748);
nand U6060 (N_6060,N_5150,N_5698);
or U6061 (N_6061,N_5323,N_5921);
and U6062 (N_6062,N_5824,N_4836);
nand U6063 (N_6063,N_4802,N_5722);
nor U6064 (N_6064,N_5457,N_5429);
and U6065 (N_6065,N_5582,N_4953);
nor U6066 (N_6066,N_5619,N_5340);
or U6067 (N_6067,N_5453,N_5022);
and U6068 (N_6068,N_5556,N_5955);
xnor U6069 (N_6069,N_5263,N_5324);
nor U6070 (N_6070,N_4879,N_5223);
xor U6071 (N_6071,N_4983,N_5782);
or U6072 (N_6072,N_5145,N_5471);
nand U6073 (N_6073,N_4849,N_5042);
or U6074 (N_6074,N_5954,N_4958);
nor U6075 (N_6075,N_5487,N_4869);
and U6076 (N_6076,N_5300,N_5591);
and U6077 (N_6077,N_4936,N_4856);
nor U6078 (N_6078,N_5133,N_5245);
xor U6079 (N_6079,N_5114,N_5853);
nor U6080 (N_6080,N_5422,N_5383);
nor U6081 (N_6081,N_4823,N_5897);
nor U6082 (N_6082,N_5900,N_5700);
xor U6083 (N_6083,N_5010,N_5336);
and U6084 (N_6084,N_5871,N_5858);
nor U6085 (N_6085,N_5638,N_5003);
or U6086 (N_6086,N_5848,N_4954);
nand U6087 (N_6087,N_5380,N_5416);
nor U6088 (N_6088,N_5075,N_5140);
and U6089 (N_6089,N_5297,N_5459);
nor U6090 (N_6090,N_5400,N_5119);
nand U6091 (N_6091,N_5766,N_5159);
or U6092 (N_6092,N_4821,N_5484);
and U6093 (N_6093,N_5850,N_4889);
nor U6094 (N_6094,N_5759,N_5090);
and U6095 (N_6095,N_4808,N_5952);
xor U6096 (N_6096,N_5640,N_5233);
and U6097 (N_6097,N_5202,N_5170);
or U6098 (N_6098,N_5681,N_5019);
nor U6099 (N_6099,N_5634,N_4899);
nand U6100 (N_6100,N_5321,N_5741);
and U6101 (N_6101,N_5052,N_5934);
xor U6102 (N_6102,N_5156,N_5697);
nor U6103 (N_6103,N_5521,N_5108);
nor U6104 (N_6104,N_5054,N_5801);
and U6105 (N_6105,N_5603,N_5372);
and U6106 (N_6106,N_5561,N_5373);
or U6107 (N_6107,N_5256,N_5221);
nor U6108 (N_6108,N_5639,N_5889);
xnor U6109 (N_6109,N_5797,N_5878);
and U6110 (N_6110,N_4918,N_5503);
and U6111 (N_6111,N_5255,N_5513);
xnor U6112 (N_6112,N_5891,N_5130);
xnor U6113 (N_6113,N_5425,N_5219);
and U6114 (N_6114,N_5819,N_5061);
or U6115 (N_6115,N_5492,N_5044);
nand U6116 (N_6116,N_5099,N_4868);
nor U6117 (N_6117,N_4854,N_5559);
nor U6118 (N_6118,N_5185,N_5342);
or U6119 (N_6119,N_5621,N_5399);
nand U6120 (N_6120,N_5124,N_5553);
xnor U6121 (N_6121,N_4925,N_5916);
nand U6122 (N_6122,N_5362,N_4982);
xnor U6123 (N_6123,N_5334,N_5395);
xor U6124 (N_6124,N_5448,N_5384);
xor U6125 (N_6125,N_5235,N_4944);
nor U6126 (N_6126,N_5294,N_5312);
and U6127 (N_6127,N_4842,N_5657);
and U6128 (N_6128,N_5112,N_5974);
nor U6129 (N_6129,N_5230,N_5776);
nand U6130 (N_6130,N_5804,N_5439);
xor U6131 (N_6131,N_5139,N_5098);
or U6132 (N_6132,N_5931,N_4805);
and U6133 (N_6133,N_5643,N_5847);
or U6134 (N_6134,N_5811,N_5873);
or U6135 (N_6135,N_5534,N_5765);
nor U6136 (N_6136,N_5569,N_5390);
and U6137 (N_6137,N_5168,N_5842);
nand U6138 (N_6138,N_5915,N_4934);
or U6139 (N_6139,N_5205,N_4887);
nand U6140 (N_6140,N_5147,N_5536);
or U6141 (N_6141,N_4861,N_5835);
or U6142 (N_6142,N_4980,N_5960);
nor U6143 (N_6143,N_5231,N_5991);
or U6144 (N_6144,N_5876,N_5946);
nor U6145 (N_6145,N_5412,N_5537);
and U6146 (N_6146,N_5790,N_5045);
nand U6147 (N_6147,N_5583,N_5618);
nor U6148 (N_6148,N_5307,N_5469);
and U6149 (N_6149,N_5176,N_4882);
nor U6150 (N_6150,N_5106,N_5261);
nor U6151 (N_6151,N_5374,N_5706);
nor U6152 (N_6152,N_5359,N_5507);
or U6153 (N_6153,N_5608,N_5142);
nand U6154 (N_6154,N_5967,N_5579);
nand U6155 (N_6155,N_5935,N_4891);
or U6156 (N_6156,N_4813,N_5500);
xor U6157 (N_6157,N_5978,N_5291);
nand U6158 (N_6158,N_5654,N_4902);
nand U6159 (N_6159,N_5214,N_5146);
nor U6160 (N_6160,N_5409,N_4840);
nand U6161 (N_6161,N_5958,N_4981);
and U6162 (N_6162,N_5014,N_4873);
and U6163 (N_6163,N_5744,N_5411);
nand U6164 (N_6164,N_5091,N_4951);
or U6165 (N_6165,N_4913,N_5547);
and U6166 (N_6166,N_5277,N_4921);
nand U6167 (N_6167,N_4926,N_5832);
or U6168 (N_6168,N_4815,N_5438);
and U6169 (N_6169,N_5129,N_4897);
nor U6170 (N_6170,N_5149,N_5375);
or U6171 (N_6171,N_5599,N_5386);
nor U6172 (N_6172,N_5226,N_5316);
nor U6173 (N_6173,N_4924,N_5434);
nor U6174 (N_6174,N_4991,N_5423);
nand U6175 (N_6175,N_5845,N_5442);
nor U6176 (N_6176,N_5201,N_5745);
xor U6177 (N_6177,N_5834,N_5035);
nand U6178 (N_6178,N_5414,N_5497);
xnor U6179 (N_6179,N_5545,N_5036);
nand U6180 (N_6180,N_5100,N_5396);
xnor U6181 (N_6181,N_5539,N_5357);
nand U6182 (N_6182,N_5026,N_5578);
and U6183 (N_6183,N_5079,N_5919);
or U6184 (N_6184,N_5341,N_5808);
and U6185 (N_6185,N_5376,N_5723);
nand U6186 (N_6186,N_5086,N_5180);
and U6187 (N_6187,N_5874,N_5320);
and U6188 (N_6188,N_5592,N_5703);
and U6189 (N_6189,N_5444,N_5240);
xor U6190 (N_6190,N_5028,N_5128);
xnor U6191 (N_6191,N_5016,N_5615);
or U6192 (N_6192,N_4930,N_5138);
nor U6193 (N_6193,N_5143,N_5495);
nand U6194 (N_6194,N_5486,N_5410);
nand U6195 (N_6195,N_4905,N_5462);
or U6196 (N_6196,N_5679,N_5292);
and U6197 (N_6197,N_5468,N_5437);
or U6198 (N_6198,N_5807,N_4973);
nor U6199 (N_6199,N_5769,N_5566);
and U6200 (N_6200,N_5996,N_5440);
xnor U6201 (N_6201,N_5800,N_5555);
xor U6202 (N_6202,N_5046,N_4986);
xnor U6203 (N_6203,N_5785,N_5560);
or U6204 (N_6204,N_5109,N_5531);
xnor U6205 (N_6205,N_5152,N_5286);
xor U6206 (N_6206,N_4855,N_5525);
or U6207 (N_6207,N_5856,N_5154);
and U6208 (N_6208,N_5609,N_5224);
nor U6209 (N_6209,N_5945,N_4883);
and U6210 (N_6210,N_5354,N_5949);
or U6211 (N_6211,N_5379,N_4949);
xnor U6212 (N_6212,N_4878,N_5356);
nor U6213 (N_6213,N_5264,N_5481);
or U6214 (N_6214,N_5505,N_5163);
and U6215 (N_6215,N_4987,N_5476);
xor U6216 (N_6216,N_5001,N_5458);
or U6217 (N_6217,N_5215,N_5980);
xnor U6218 (N_6218,N_5450,N_4970);
nand U6219 (N_6219,N_5222,N_5266);
xor U6220 (N_6220,N_5933,N_5118);
and U6221 (N_6221,N_5095,N_5254);
and U6222 (N_6222,N_5217,N_5456);
or U6223 (N_6223,N_4929,N_4803);
nand U6224 (N_6224,N_5455,N_5134);
nor U6225 (N_6225,N_4885,N_5859);
or U6226 (N_6226,N_5709,N_5794);
nand U6227 (N_6227,N_5588,N_5177);
and U6228 (N_6228,N_5466,N_5346);
and U6229 (N_6229,N_5234,N_5651);
xnor U6230 (N_6230,N_5183,N_5554);
and U6231 (N_6231,N_5287,N_5549);
nor U6232 (N_6232,N_5072,N_5849);
nor U6233 (N_6233,N_4907,N_5115);
nor U6234 (N_6234,N_5664,N_5311);
and U6235 (N_6235,N_4846,N_5085);
nand U6236 (N_6236,N_5251,N_5025);
nand U6237 (N_6237,N_5273,N_4894);
or U6238 (N_6238,N_4912,N_5123);
xor U6239 (N_6239,N_4904,N_5632);
and U6240 (N_6240,N_5451,N_5293);
xnor U6241 (N_6241,N_5864,N_5792);
xnor U6242 (N_6242,N_5446,N_4910);
and U6243 (N_6243,N_5107,N_4942);
and U6244 (N_6244,N_4988,N_5220);
and U6245 (N_6245,N_5267,N_5546);
nor U6246 (N_6246,N_5418,N_5707);
or U6247 (N_6247,N_5461,N_5299);
nor U6248 (N_6248,N_5886,N_4938);
xnor U6249 (N_6249,N_5203,N_5812);
nor U6250 (N_6250,N_5844,N_4920);
or U6251 (N_6251,N_5358,N_5731);
xnor U6252 (N_6252,N_5966,N_5189);
nand U6253 (N_6253,N_5082,N_5512);
nor U6254 (N_6254,N_5447,N_5449);
or U6255 (N_6255,N_5866,N_5284);
nand U6256 (N_6256,N_5059,N_5097);
nand U6257 (N_6257,N_5051,N_5232);
xnor U6258 (N_6258,N_5714,N_5252);
or U6259 (N_6259,N_5726,N_5905);
and U6260 (N_6260,N_5058,N_4837);
nor U6261 (N_6261,N_5605,N_5777);
nand U6262 (N_6262,N_4892,N_5039);
nand U6263 (N_6263,N_5894,N_4826);
nor U6264 (N_6264,N_4848,N_5276);
and U6265 (N_6265,N_4985,N_5577);
and U6266 (N_6266,N_4996,N_5508);
nor U6267 (N_6267,N_5815,N_5065);
xor U6268 (N_6268,N_5870,N_5656);
nor U6269 (N_6269,N_4964,N_5313);
or U6270 (N_6270,N_4853,N_5288);
xnor U6271 (N_6271,N_5367,N_5424);
or U6272 (N_6272,N_5274,N_5696);
nand U6273 (N_6273,N_4886,N_5278);
or U6274 (N_6274,N_5676,N_5228);
nand U6275 (N_6275,N_5196,N_5793);
xnor U6276 (N_6276,N_5113,N_5524);
xor U6277 (N_6277,N_5435,N_4807);
and U6278 (N_6278,N_5925,N_5033);
nor U6279 (N_6279,N_5667,N_5784);
nand U6280 (N_6280,N_5490,N_5094);
xnor U6281 (N_6281,N_5913,N_5998);
or U6282 (N_6282,N_5918,N_5869);
or U6283 (N_6283,N_5198,N_5136);
and U6284 (N_6284,N_4974,N_5601);
nand U6285 (N_6285,N_5570,N_5822);
nor U6286 (N_6286,N_4943,N_4922);
nand U6287 (N_6287,N_5413,N_5965);
nand U6288 (N_6288,N_5786,N_5258);
xor U6289 (N_6289,N_4877,N_5305);
nor U6290 (N_6290,N_5861,N_5581);
xor U6291 (N_6291,N_5746,N_5247);
and U6292 (N_6292,N_4908,N_5496);
nand U6293 (N_6293,N_5067,N_5403);
xnor U6294 (N_6294,N_5780,N_4952);
and U6295 (N_6295,N_5105,N_5371);
xor U6296 (N_6296,N_5962,N_5749);
and U6297 (N_6297,N_4898,N_5474);
nand U6298 (N_6298,N_4862,N_4998);
nand U6299 (N_6299,N_4978,N_5355);
xnor U6300 (N_6300,N_5007,N_5733);
nor U6301 (N_6301,N_5066,N_5678);
nor U6302 (N_6302,N_5783,N_4828);
and U6303 (N_6303,N_5077,N_5074);
and U6304 (N_6304,N_5430,N_5903);
nor U6305 (N_6305,N_5926,N_5702);
or U6306 (N_6306,N_5999,N_5550);
nor U6307 (N_6307,N_5795,N_4997);
or U6308 (N_6308,N_5008,N_5103);
and U6309 (N_6309,N_5131,N_5408);
xnor U6310 (N_6310,N_4931,N_5337);
xor U6311 (N_6311,N_5050,N_5939);
xnor U6312 (N_6312,N_5250,N_5506);
or U6313 (N_6313,N_5805,N_5319);
nand U6314 (N_6314,N_5053,N_4844);
xnor U6315 (N_6315,N_5445,N_5433);
nand U6316 (N_6316,N_5104,N_5364);
xnor U6317 (N_6317,N_5768,N_5463);
nor U6318 (N_6318,N_5837,N_5349);
and U6319 (N_6319,N_5191,N_5595);
xor U6320 (N_6320,N_5902,N_5627);
nor U6321 (N_6321,N_4999,N_4966);
nand U6322 (N_6322,N_5719,N_4967);
nor U6323 (N_6323,N_5350,N_5761);
nand U6324 (N_6324,N_5006,N_5936);
and U6325 (N_6325,N_5881,N_4830);
and U6326 (N_6326,N_5175,N_5405);
nor U6327 (N_6327,N_5034,N_5630);
xor U6328 (N_6328,N_5865,N_5585);
and U6329 (N_6329,N_5190,N_5322);
nand U6330 (N_6330,N_5778,N_5872);
nand U6331 (N_6331,N_4901,N_5253);
or U6332 (N_6332,N_4820,N_5441);
nand U6333 (N_6333,N_5167,N_5574);
nand U6334 (N_6334,N_5799,N_5892);
nor U6335 (N_6335,N_5997,N_5165);
xnor U6336 (N_6336,N_5682,N_4832);
xnor U6337 (N_6337,N_5907,N_5432);
nor U6338 (N_6338,N_5739,N_5329);
nor U6339 (N_6339,N_4852,N_5060);
or U6340 (N_6340,N_5529,N_4838);
nand U6341 (N_6341,N_5984,N_4857);
nand U6342 (N_6342,N_4810,N_4939);
and U6343 (N_6343,N_5389,N_5348);
nand U6344 (N_6344,N_5211,N_5716);
xor U6345 (N_6345,N_5694,N_5188);
nand U6346 (N_6346,N_5880,N_5101);
and U6347 (N_6347,N_5132,N_5820);
xnor U6348 (N_6348,N_5774,N_4859);
or U6349 (N_6349,N_5622,N_5218);
nor U6350 (N_6350,N_5713,N_5518);
xnor U6351 (N_6351,N_4824,N_5426);
xor U6352 (N_6352,N_5580,N_5613);
nand U6353 (N_6353,N_5004,N_5764);
and U6354 (N_6354,N_5281,N_5717);
and U6355 (N_6355,N_5597,N_5677);
or U6356 (N_6356,N_5756,N_5773);
nor U6357 (N_6357,N_5540,N_5111);
nor U6358 (N_6358,N_5069,N_5666);
nand U6359 (N_6359,N_5690,N_4865);
or U6360 (N_6360,N_5182,N_5502);
nand U6361 (N_6361,N_5590,N_5102);
nand U6362 (N_6362,N_5879,N_5637);
nand U6363 (N_6363,N_5542,N_5575);
and U6364 (N_6364,N_5890,N_5332);
nor U6365 (N_6365,N_5551,N_5742);
nand U6366 (N_6366,N_5721,N_5377);
nor U6367 (N_6367,N_5331,N_4817);
nand U6368 (N_6368,N_5750,N_5598);
and U6369 (N_6369,N_5983,N_4860);
and U6370 (N_6370,N_5295,N_5576);
nor U6371 (N_6371,N_5887,N_5747);
and U6372 (N_6372,N_5526,N_5990);
nand U6373 (N_6373,N_5478,N_4835);
xnor U6374 (N_6374,N_5527,N_4834);
or U6375 (N_6375,N_5953,N_5161);
nor U6376 (N_6376,N_5096,N_5024);
or U6377 (N_6377,N_5635,N_4940);
nor U6378 (N_6378,N_5976,N_5544);
nor U6379 (N_6379,N_5922,N_5940);
and U6380 (N_6380,N_4839,N_5282);
and U6381 (N_6381,N_5840,N_5279);
nor U6382 (N_6382,N_5779,N_5283);
and U6383 (N_6383,N_5961,N_5909);
or U6384 (N_6384,N_5268,N_5280);
nor U6385 (N_6385,N_5736,N_4809);
nor U6386 (N_6386,N_5419,N_5116);
nand U6387 (N_6387,N_5631,N_5938);
nor U6388 (N_6388,N_5000,N_4977);
nor U6389 (N_6389,N_5854,N_5788);
nand U6390 (N_6390,N_5499,N_5246);
xor U6391 (N_6391,N_5941,N_5498);
or U6392 (N_6392,N_5633,N_5017);
and U6393 (N_6393,N_4818,N_5125);
and U6394 (N_6394,N_5924,N_4975);
xor U6395 (N_6395,N_4819,N_5791);
nor U6396 (N_6396,N_5920,N_5867);
and U6397 (N_6397,N_5855,N_5257);
nand U6398 (N_6398,N_5056,N_5083);
and U6399 (N_6399,N_4961,N_4822);
nand U6400 (N_6400,N_5078,N_5192);
nor U6401 (N_6401,N_5838,N_5728);
nor U6402 (N_6402,N_5589,N_5992);
or U6403 (N_6403,N_5904,N_5727);
nand U6404 (N_6404,N_5290,N_5370);
xnor U6405 (N_6405,N_5928,N_5301);
or U6406 (N_6406,N_5345,N_5898);
xor U6407 (N_6407,N_5420,N_5216);
nand U6408 (N_6408,N_5557,N_5645);
xor U6409 (N_6409,N_5612,N_5950);
nand U6410 (N_6410,N_4812,N_5084);
or U6411 (N_6411,N_5584,N_5628);
xnor U6412 (N_6412,N_4804,N_5360);
and U6413 (N_6413,N_4963,N_5564);
nor U6414 (N_6414,N_5339,N_4825);
and U6415 (N_6415,N_5173,N_5594);
nor U6416 (N_6416,N_5908,N_5771);
nand U6417 (N_6417,N_5157,N_4917);
and U6418 (N_6418,N_5186,N_5473);
xnor U6419 (N_6419,N_5650,N_5494);
and U6420 (N_6420,N_5937,N_5767);
nor U6421 (N_6421,N_5309,N_4923);
and U6422 (N_6422,N_5172,N_5729);
nor U6423 (N_6423,N_5184,N_5956);
xnor U6424 (N_6424,N_5981,N_4959);
nand U6425 (N_6425,N_5705,N_4946);
and U6426 (N_6426,N_4968,N_5718);
and U6427 (N_6427,N_5942,N_5818);
nor U6428 (N_6428,N_5885,N_5567);
and U6429 (N_6429,N_5827,N_5302);
and U6430 (N_6430,N_5047,N_5141);
and U6431 (N_6431,N_4829,N_4850);
or U6432 (N_6432,N_5239,N_5187);
and U6433 (N_6433,N_5388,N_5641);
and U6434 (N_6434,N_4884,N_5680);
nor U6435 (N_6435,N_5882,N_5151);
and U6436 (N_6436,N_5236,N_5911);
nor U6437 (N_6437,N_5068,N_5365);
xor U6438 (N_6438,N_5810,N_5787);
nand U6439 (N_6439,N_5673,N_5158);
or U6440 (N_6440,N_5225,N_5989);
nand U6441 (N_6441,N_5543,N_4831);
and U6442 (N_6442,N_5392,N_5027);
and U6443 (N_6443,N_5646,N_5135);
and U6444 (N_6444,N_5516,N_5644);
nand U6445 (N_6445,N_5649,N_5813);
or U6446 (N_6446,N_5757,N_5353);
and U6447 (N_6447,N_5760,N_5652);
or U6448 (N_6448,N_5394,N_5781);
or U6449 (N_6449,N_4937,N_5166);
nand U6450 (N_6450,N_5831,N_5262);
xor U6451 (N_6451,N_5366,N_5636);
nand U6452 (N_6452,N_5735,N_5009);
and U6453 (N_6453,N_5467,N_5213);
or U6454 (N_6454,N_4950,N_5668);
xor U6455 (N_6455,N_5972,N_5689);
or U6456 (N_6456,N_5171,N_5110);
or U6457 (N_6457,N_4890,N_5665);
nand U6458 (N_6458,N_5565,N_4976);
nor U6459 (N_6459,N_5401,N_5153);
nand U6460 (N_6460,N_4956,N_5662);
or U6461 (N_6461,N_5237,N_5762);
nor U6462 (N_6462,N_5315,N_5883);
nand U6463 (N_6463,N_5063,N_5982);
xnor U6464 (N_6464,N_5530,N_5510);
xor U6465 (N_6465,N_5368,N_5893);
nand U6466 (N_6466,N_4915,N_5671);
or U6467 (N_6467,N_4800,N_5573);
xor U6468 (N_6468,N_4871,N_5511);
xnor U6469 (N_6469,N_5675,N_4843);
nand U6470 (N_6470,N_5243,N_5117);
nand U6471 (N_6471,N_5846,N_5464);
nor U6472 (N_6472,N_5427,N_5021);
and U6473 (N_6473,N_5602,N_5642);
and U6474 (N_6474,N_5229,N_5672);
xnor U6475 (N_6475,N_5995,N_5285);
and U6476 (N_6476,N_5523,N_5482);
nor U6477 (N_6477,N_5314,N_5725);
nand U6478 (N_6478,N_5073,N_5971);
and U6479 (N_6479,N_5206,N_5796);
nand U6480 (N_6480,N_5970,N_5724);
or U6481 (N_6481,N_5712,N_5692);
xnor U6482 (N_6482,N_5730,N_5397);
or U6483 (N_6483,N_5715,N_5738);
xnor U6484 (N_6484,N_5020,N_5711);
or U6485 (N_6485,N_5041,N_5851);
xnor U6486 (N_6486,N_5743,N_4962);
and U6487 (N_6487,N_5617,N_5823);
nor U6488 (N_6488,N_5071,N_4845);
nor U6489 (N_6489,N_5080,N_5387);
nand U6490 (N_6490,N_5658,N_5164);
and U6491 (N_6491,N_5012,N_4941);
xor U6492 (N_6492,N_4955,N_4881);
nor U6493 (N_6493,N_4972,N_5127);
nand U6494 (N_6494,N_5018,N_4896);
or U6495 (N_6495,N_5687,N_5944);
and U6496 (N_6496,N_5002,N_5737);
xor U6497 (N_6497,N_4984,N_5289);
or U6498 (N_6498,N_4880,N_4806);
nor U6499 (N_6499,N_5514,N_5162);
or U6500 (N_6500,N_5087,N_5655);
nand U6501 (N_6501,N_5661,N_4927);
xnor U6502 (N_6502,N_5674,N_5695);
nand U6503 (N_6503,N_5629,N_5607);
nor U6504 (N_6504,N_5901,N_4979);
or U6505 (N_6505,N_5005,N_5057);
nor U6506 (N_6506,N_5043,N_5571);
or U6507 (N_6507,N_5015,N_5296);
nor U6508 (N_6508,N_5470,N_5896);
nand U6509 (N_6509,N_5488,N_5382);
nand U6510 (N_6510,N_5076,N_5520);
nand U6511 (N_6511,N_5195,N_5857);
nor U6512 (N_6512,N_5417,N_5587);
nand U6513 (N_6513,N_5917,N_5011);
and U6514 (N_6514,N_5806,N_5860);
nor U6515 (N_6515,N_5306,N_5986);
or U6516 (N_6516,N_5475,N_5973);
xnor U6517 (N_6517,N_5528,N_5242);
nor U6518 (N_6518,N_5732,N_5568);
and U6519 (N_6519,N_5685,N_4960);
xnor U6520 (N_6520,N_5241,N_5308);
or U6521 (N_6521,N_4932,N_5888);
xnor U6522 (N_6522,N_4876,N_5269);
xnor U6523 (N_6523,N_5604,N_5912);
or U6524 (N_6524,N_5330,N_5660);
nand U6525 (N_6525,N_5817,N_5204);
nand U6526 (N_6526,N_5647,N_4870);
and U6527 (N_6527,N_4947,N_4971);
or U6528 (N_6528,N_5275,N_4816);
or U6529 (N_6529,N_5816,N_5775);
nor U6530 (N_6530,N_5614,N_5363);
nor U6531 (N_6531,N_5436,N_5535);
nand U6532 (N_6532,N_5318,N_5862);
and U6533 (N_6533,N_5248,N_5501);
xor U6534 (N_6534,N_5326,N_5930);
nand U6535 (N_6535,N_5875,N_4919);
nand U6536 (N_6536,N_5317,N_5963);
or U6537 (N_6537,N_5483,N_5352);
xnor U6538 (N_6538,N_5975,N_4995);
xnor U6539 (N_6539,N_4989,N_5402);
nand U6540 (N_6540,N_5552,N_4841);
xor U6541 (N_6541,N_5517,N_5751);
xor U6542 (N_6542,N_5979,N_5753);
nand U6543 (N_6543,N_5178,N_5863);
or U6544 (N_6544,N_5030,N_5328);
nand U6545 (N_6545,N_5985,N_5828);
or U6546 (N_6546,N_5338,N_5538);
and U6547 (N_6547,N_5193,N_5899);
xnor U6548 (N_6548,N_4903,N_4928);
and U6549 (N_6549,N_4909,N_5489);
xnor U6550 (N_6550,N_5606,N_5821);
nor U6551 (N_6551,N_5304,N_5428);
nor U6552 (N_6552,N_5259,N_5174);
or U6553 (N_6553,N_5663,N_5533);
or U6554 (N_6554,N_5031,N_5720);
xor U6555 (N_6555,N_5572,N_5122);
nor U6556 (N_6556,N_5548,N_4900);
nand U6557 (N_6557,N_5932,N_5137);
nor U6558 (N_6558,N_5648,N_5789);
and U6559 (N_6559,N_5620,N_5431);
xor U6560 (N_6560,N_5825,N_4814);
nand U6561 (N_6561,N_5089,N_5515);
or U6562 (N_6562,N_5504,N_5200);
or U6563 (N_6563,N_5943,N_4864);
nor U6564 (N_6564,N_5249,N_4895);
nor U6565 (N_6565,N_5032,N_5929);
xnor U6566 (N_6566,N_5988,N_5335);
nand U6567 (N_6567,N_5701,N_5040);
xnor U6568 (N_6568,N_5298,N_5829);
or U6569 (N_6569,N_5959,N_5563);
xnor U6570 (N_6570,N_5160,N_4965);
or U6571 (N_6571,N_5343,N_5532);
and U6572 (N_6572,N_5927,N_5948);
or U6573 (N_6573,N_5586,N_5210);
or U6574 (N_6574,N_5452,N_5914);
nor U6575 (N_6575,N_5852,N_5391);
or U6576 (N_6576,N_5093,N_5144);
xor U6577 (N_6577,N_5623,N_4957);
nand U6578 (N_6578,N_5194,N_5155);
xor U6579 (N_6579,N_5670,N_4916);
and U6580 (N_6580,N_4872,N_5351);
nand U6581 (N_6581,N_5271,N_5327);
nand U6582 (N_6582,N_5833,N_5037);
nor U6583 (N_6583,N_4866,N_4914);
and U6584 (N_6584,N_5839,N_5055);
and U6585 (N_6585,N_5593,N_5659);
xnor U6586 (N_6586,N_5385,N_5684);
nand U6587 (N_6587,N_5519,N_5029);
or U6588 (N_6588,N_5843,N_5669);
and U6589 (N_6589,N_5558,N_5369);
nor U6590 (N_6590,N_5013,N_5121);
and U6591 (N_6591,N_5260,N_5212);
or U6592 (N_6592,N_5754,N_5626);
and U6593 (N_6593,N_5491,N_4801);
or U6594 (N_6594,N_5752,N_5798);
nor U6595 (N_6595,N_4893,N_5994);
and U6596 (N_6596,N_5460,N_5868);
xor U6597 (N_6597,N_5181,N_5802);
or U6598 (N_6598,N_5209,N_5809);
or U6599 (N_6599,N_4945,N_5415);
nand U6600 (N_6600,N_5628,N_5629);
xnor U6601 (N_6601,N_5294,N_5578);
nand U6602 (N_6602,N_5822,N_5277);
nand U6603 (N_6603,N_5696,N_4876);
xnor U6604 (N_6604,N_5445,N_5289);
and U6605 (N_6605,N_5706,N_4839);
or U6606 (N_6606,N_5317,N_5926);
nor U6607 (N_6607,N_5975,N_5109);
and U6608 (N_6608,N_5730,N_5685);
xor U6609 (N_6609,N_5060,N_5360);
and U6610 (N_6610,N_5050,N_5009);
nor U6611 (N_6611,N_4949,N_5548);
or U6612 (N_6612,N_4897,N_5064);
and U6613 (N_6613,N_5159,N_5677);
or U6614 (N_6614,N_5427,N_5687);
nor U6615 (N_6615,N_5047,N_4990);
nand U6616 (N_6616,N_5378,N_5509);
and U6617 (N_6617,N_4843,N_5201);
nand U6618 (N_6618,N_5260,N_5836);
xor U6619 (N_6619,N_4855,N_5329);
xnor U6620 (N_6620,N_5488,N_5304);
or U6621 (N_6621,N_5408,N_5037);
or U6622 (N_6622,N_5095,N_5548);
and U6623 (N_6623,N_5542,N_5345);
and U6624 (N_6624,N_5615,N_5939);
nand U6625 (N_6625,N_5730,N_5178);
and U6626 (N_6626,N_5800,N_5502);
and U6627 (N_6627,N_4912,N_5904);
or U6628 (N_6628,N_5575,N_5041);
nand U6629 (N_6629,N_4973,N_5702);
or U6630 (N_6630,N_5896,N_5448);
xnor U6631 (N_6631,N_5921,N_5581);
xor U6632 (N_6632,N_4974,N_5573);
xor U6633 (N_6633,N_5222,N_5551);
nor U6634 (N_6634,N_5938,N_4833);
nand U6635 (N_6635,N_5454,N_5416);
and U6636 (N_6636,N_4979,N_5142);
or U6637 (N_6637,N_4923,N_5811);
nor U6638 (N_6638,N_5480,N_5253);
or U6639 (N_6639,N_5068,N_5718);
or U6640 (N_6640,N_5154,N_5327);
and U6641 (N_6641,N_5929,N_5968);
and U6642 (N_6642,N_5354,N_5546);
and U6643 (N_6643,N_5095,N_5854);
and U6644 (N_6644,N_4854,N_5536);
xor U6645 (N_6645,N_5686,N_5270);
and U6646 (N_6646,N_5500,N_5861);
nand U6647 (N_6647,N_5769,N_4805);
and U6648 (N_6648,N_5044,N_5900);
nor U6649 (N_6649,N_5150,N_4973);
xnor U6650 (N_6650,N_4950,N_5733);
and U6651 (N_6651,N_5139,N_5774);
and U6652 (N_6652,N_4946,N_5782);
xor U6653 (N_6653,N_4934,N_4855);
nor U6654 (N_6654,N_4824,N_4860);
nand U6655 (N_6655,N_5936,N_5958);
nand U6656 (N_6656,N_5216,N_4972);
nand U6657 (N_6657,N_5060,N_5763);
xnor U6658 (N_6658,N_5260,N_5980);
or U6659 (N_6659,N_5977,N_5215);
and U6660 (N_6660,N_4932,N_4812);
nand U6661 (N_6661,N_5700,N_5765);
nand U6662 (N_6662,N_5911,N_5907);
xor U6663 (N_6663,N_5953,N_5795);
or U6664 (N_6664,N_5848,N_5907);
xnor U6665 (N_6665,N_5281,N_4903);
nand U6666 (N_6666,N_5137,N_5354);
xor U6667 (N_6667,N_5725,N_5304);
nand U6668 (N_6668,N_4952,N_5793);
nand U6669 (N_6669,N_4942,N_5357);
xor U6670 (N_6670,N_5947,N_5083);
and U6671 (N_6671,N_5776,N_4986);
nor U6672 (N_6672,N_5323,N_5543);
nor U6673 (N_6673,N_5334,N_5483);
nor U6674 (N_6674,N_5518,N_5520);
xnor U6675 (N_6675,N_5367,N_5562);
or U6676 (N_6676,N_5385,N_5386);
nand U6677 (N_6677,N_5702,N_5843);
or U6678 (N_6678,N_5464,N_5199);
or U6679 (N_6679,N_5062,N_5903);
nand U6680 (N_6680,N_4819,N_5176);
nor U6681 (N_6681,N_5105,N_5647);
xnor U6682 (N_6682,N_5838,N_4834);
nor U6683 (N_6683,N_5024,N_5063);
xor U6684 (N_6684,N_5077,N_5774);
nand U6685 (N_6685,N_5289,N_5813);
nand U6686 (N_6686,N_5850,N_5950);
and U6687 (N_6687,N_5349,N_5047);
xnor U6688 (N_6688,N_5641,N_5956);
nor U6689 (N_6689,N_5045,N_5816);
xor U6690 (N_6690,N_5765,N_5341);
xor U6691 (N_6691,N_5408,N_5607);
or U6692 (N_6692,N_4923,N_5258);
or U6693 (N_6693,N_5617,N_5136);
or U6694 (N_6694,N_5814,N_4937);
nor U6695 (N_6695,N_5193,N_5448);
or U6696 (N_6696,N_5152,N_5505);
nor U6697 (N_6697,N_4939,N_5735);
nand U6698 (N_6698,N_5864,N_5506);
nor U6699 (N_6699,N_5009,N_5636);
and U6700 (N_6700,N_4998,N_5114);
or U6701 (N_6701,N_4805,N_4942);
or U6702 (N_6702,N_5850,N_4930);
and U6703 (N_6703,N_4963,N_5661);
and U6704 (N_6704,N_5719,N_4899);
and U6705 (N_6705,N_5734,N_5177);
nor U6706 (N_6706,N_5155,N_5616);
and U6707 (N_6707,N_5323,N_4835);
xor U6708 (N_6708,N_5654,N_5428);
nand U6709 (N_6709,N_5984,N_5771);
and U6710 (N_6710,N_5685,N_5595);
nor U6711 (N_6711,N_5276,N_5873);
xnor U6712 (N_6712,N_4847,N_5880);
xnor U6713 (N_6713,N_5764,N_5421);
nand U6714 (N_6714,N_5967,N_5624);
nand U6715 (N_6715,N_5029,N_5121);
nor U6716 (N_6716,N_4826,N_5557);
or U6717 (N_6717,N_5631,N_5612);
nor U6718 (N_6718,N_5870,N_5427);
or U6719 (N_6719,N_5667,N_5365);
nor U6720 (N_6720,N_5058,N_5818);
or U6721 (N_6721,N_5599,N_5929);
and U6722 (N_6722,N_5973,N_5581);
nand U6723 (N_6723,N_5891,N_5362);
xnor U6724 (N_6724,N_4913,N_4857);
xor U6725 (N_6725,N_4988,N_5387);
xnor U6726 (N_6726,N_5334,N_5339);
nor U6727 (N_6727,N_5816,N_4845);
and U6728 (N_6728,N_5151,N_5161);
and U6729 (N_6729,N_4904,N_5602);
nor U6730 (N_6730,N_5811,N_5766);
and U6731 (N_6731,N_5065,N_5943);
or U6732 (N_6732,N_5090,N_5419);
and U6733 (N_6733,N_5386,N_5803);
nand U6734 (N_6734,N_5450,N_5716);
or U6735 (N_6735,N_5090,N_4958);
nor U6736 (N_6736,N_4982,N_5419);
and U6737 (N_6737,N_5165,N_5886);
or U6738 (N_6738,N_5459,N_5842);
xnor U6739 (N_6739,N_5717,N_5523);
xnor U6740 (N_6740,N_5726,N_4813);
nor U6741 (N_6741,N_5886,N_5487);
nand U6742 (N_6742,N_5949,N_4827);
and U6743 (N_6743,N_5298,N_4959);
nor U6744 (N_6744,N_5872,N_5504);
or U6745 (N_6745,N_5620,N_5302);
or U6746 (N_6746,N_4988,N_5276);
or U6747 (N_6747,N_5900,N_5564);
xnor U6748 (N_6748,N_4921,N_5653);
xnor U6749 (N_6749,N_5459,N_5661);
and U6750 (N_6750,N_5229,N_5396);
or U6751 (N_6751,N_5659,N_5460);
or U6752 (N_6752,N_4936,N_5347);
nand U6753 (N_6753,N_5115,N_5825);
xor U6754 (N_6754,N_5493,N_5274);
nor U6755 (N_6755,N_5265,N_5214);
xnor U6756 (N_6756,N_5886,N_5393);
xnor U6757 (N_6757,N_4821,N_5864);
or U6758 (N_6758,N_5562,N_5492);
nand U6759 (N_6759,N_5435,N_5507);
nor U6760 (N_6760,N_5444,N_5684);
or U6761 (N_6761,N_4830,N_5753);
or U6762 (N_6762,N_5984,N_4955);
nand U6763 (N_6763,N_5032,N_4971);
and U6764 (N_6764,N_5245,N_5606);
nor U6765 (N_6765,N_5075,N_4898);
xor U6766 (N_6766,N_5458,N_5331);
or U6767 (N_6767,N_5531,N_4966);
or U6768 (N_6768,N_5564,N_5336);
xnor U6769 (N_6769,N_4965,N_5271);
xor U6770 (N_6770,N_5002,N_5053);
nor U6771 (N_6771,N_5465,N_5933);
or U6772 (N_6772,N_5816,N_5755);
xor U6773 (N_6773,N_5977,N_5893);
and U6774 (N_6774,N_5698,N_4835);
and U6775 (N_6775,N_5356,N_5857);
nor U6776 (N_6776,N_5261,N_5846);
nand U6777 (N_6777,N_4884,N_5826);
xnor U6778 (N_6778,N_5928,N_4845);
xor U6779 (N_6779,N_5017,N_5292);
nand U6780 (N_6780,N_5067,N_4862);
nand U6781 (N_6781,N_5652,N_5626);
nand U6782 (N_6782,N_5186,N_4981);
nor U6783 (N_6783,N_5401,N_4800);
or U6784 (N_6784,N_5085,N_5241);
nand U6785 (N_6785,N_5748,N_5920);
nor U6786 (N_6786,N_5337,N_5143);
xor U6787 (N_6787,N_5518,N_5971);
or U6788 (N_6788,N_5073,N_5049);
and U6789 (N_6789,N_5869,N_4974);
nand U6790 (N_6790,N_5931,N_5688);
nor U6791 (N_6791,N_4956,N_5688);
or U6792 (N_6792,N_5032,N_4989);
nand U6793 (N_6793,N_5030,N_5327);
or U6794 (N_6794,N_5587,N_5277);
or U6795 (N_6795,N_5650,N_5457);
xnor U6796 (N_6796,N_5412,N_5179);
and U6797 (N_6797,N_5490,N_5614);
nand U6798 (N_6798,N_5920,N_5908);
nor U6799 (N_6799,N_5495,N_5425);
nor U6800 (N_6800,N_4975,N_4976);
nor U6801 (N_6801,N_5010,N_5722);
and U6802 (N_6802,N_4959,N_5346);
nand U6803 (N_6803,N_4867,N_5078);
nor U6804 (N_6804,N_5163,N_5708);
nand U6805 (N_6805,N_5157,N_4884);
and U6806 (N_6806,N_5415,N_5619);
and U6807 (N_6807,N_4849,N_4883);
nand U6808 (N_6808,N_5262,N_5695);
nor U6809 (N_6809,N_5856,N_5014);
nor U6810 (N_6810,N_4942,N_5589);
xor U6811 (N_6811,N_5981,N_5155);
xor U6812 (N_6812,N_5572,N_5751);
nand U6813 (N_6813,N_5991,N_5877);
or U6814 (N_6814,N_5641,N_5099);
and U6815 (N_6815,N_5856,N_5438);
nor U6816 (N_6816,N_5344,N_5389);
and U6817 (N_6817,N_5745,N_5344);
nand U6818 (N_6818,N_4984,N_5288);
nor U6819 (N_6819,N_5576,N_5985);
nand U6820 (N_6820,N_4955,N_5618);
nor U6821 (N_6821,N_5557,N_5013);
xnor U6822 (N_6822,N_5646,N_5991);
and U6823 (N_6823,N_5157,N_5872);
nand U6824 (N_6824,N_5664,N_4902);
or U6825 (N_6825,N_4848,N_5933);
nand U6826 (N_6826,N_5377,N_5666);
or U6827 (N_6827,N_5940,N_4908);
xnor U6828 (N_6828,N_5354,N_5197);
xor U6829 (N_6829,N_5827,N_5448);
xor U6830 (N_6830,N_5395,N_5392);
nor U6831 (N_6831,N_5263,N_5372);
nor U6832 (N_6832,N_5013,N_5814);
xnor U6833 (N_6833,N_4880,N_5734);
nor U6834 (N_6834,N_5395,N_5637);
and U6835 (N_6835,N_5703,N_5314);
nor U6836 (N_6836,N_5875,N_5294);
nor U6837 (N_6837,N_5970,N_5865);
nor U6838 (N_6838,N_4935,N_5101);
and U6839 (N_6839,N_5432,N_5187);
or U6840 (N_6840,N_5936,N_5976);
nor U6841 (N_6841,N_5658,N_5957);
and U6842 (N_6842,N_5840,N_5652);
and U6843 (N_6843,N_5825,N_5827);
xnor U6844 (N_6844,N_5467,N_5132);
xor U6845 (N_6845,N_5618,N_5520);
or U6846 (N_6846,N_5298,N_5593);
xor U6847 (N_6847,N_5978,N_5497);
nor U6848 (N_6848,N_5687,N_5554);
nor U6849 (N_6849,N_5521,N_4941);
and U6850 (N_6850,N_5070,N_4970);
nand U6851 (N_6851,N_5635,N_5072);
or U6852 (N_6852,N_5999,N_4814);
xnor U6853 (N_6853,N_5260,N_4882);
and U6854 (N_6854,N_5394,N_5370);
nand U6855 (N_6855,N_5687,N_5368);
nor U6856 (N_6856,N_5826,N_5731);
nand U6857 (N_6857,N_5513,N_5589);
nor U6858 (N_6858,N_5975,N_5000);
nand U6859 (N_6859,N_5317,N_5986);
xor U6860 (N_6860,N_4814,N_5357);
nor U6861 (N_6861,N_5472,N_4824);
and U6862 (N_6862,N_5849,N_5867);
and U6863 (N_6863,N_5118,N_5144);
nor U6864 (N_6864,N_5428,N_5536);
and U6865 (N_6865,N_5602,N_4980);
and U6866 (N_6866,N_5967,N_5130);
xnor U6867 (N_6867,N_4906,N_5857);
nor U6868 (N_6868,N_5461,N_4811);
xor U6869 (N_6869,N_5262,N_5959);
or U6870 (N_6870,N_5028,N_5628);
nor U6871 (N_6871,N_5478,N_5940);
or U6872 (N_6872,N_5498,N_5037);
xor U6873 (N_6873,N_4954,N_5235);
and U6874 (N_6874,N_5555,N_5112);
xor U6875 (N_6875,N_5576,N_4854);
or U6876 (N_6876,N_5924,N_5903);
or U6877 (N_6877,N_5856,N_5876);
nand U6878 (N_6878,N_4802,N_5578);
xor U6879 (N_6879,N_4982,N_5128);
nand U6880 (N_6880,N_4823,N_5658);
nor U6881 (N_6881,N_5271,N_5526);
and U6882 (N_6882,N_5625,N_5131);
and U6883 (N_6883,N_5009,N_5384);
and U6884 (N_6884,N_5566,N_5803);
and U6885 (N_6885,N_5237,N_5156);
or U6886 (N_6886,N_5426,N_5652);
nand U6887 (N_6887,N_5312,N_5651);
xor U6888 (N_6888,N_4990,N_4963);
nand U6889 (N_6889,N_5581,N_4820);
nor U6890 (N_6890,N_5861,N_5614);
nor U6891 (N_6891,N_4814,N_5411);
or U6892 (N_6892,N_4968,N_4815);
nand U6893 (N_6893,N_5295,N_5143);
nand U6894 (N_6894,N_5949,N_5476);
and U6895 (N_6895,N_5858,N_5598);
nand U6896 (N_6896,N_5688,N_5113);
nor U6897 (N_6897,N_5713,N_5945);
or U6898 (N_6898,N_5282,N_4856);
nor U6899 (N_6899,N_5045,N_5724);
xnor U6900 (N_6900,N_5002,N_5596);
nor U6901 (N_6901,N_5630,N_5014);
nand U6902 (N_6902,N_5673,N_5208);
nor U6903 (N_6903,N_5498,N_5103);
and U6904 (N_6904,N_5757,N_5334);
nand U6905 (N_6905,N_4829,N_5838);
nand U6906 (N_6906,N_5120,N_5195);
or U6907 (N_6907,N_5141,N_5334);
or U6908 (N_6908,N_5965,N_4981);
nand U6909 (N_6909,N_4925,N_5705);
nor U6910 (N_6910,N_5247,N_5345);
nand U6911 (N_6911,N_4970,N_5924);
nand U6912 (N_6912,N_4957,N_5361);
and U6913 (N_6913,N_4935,N_5693);
xor U6914 (N_6914,N_5863,N_5785);
xor U6915 (N_6915,N_5573,N_5232);
or U6916 (N_6916,N_5492,N_5320);
and U6917 (N_6917,N_5797,N_5142);
or U6918 (N_6918,N_5589,N_5073);
nand U6919 (N_6919,N_5508,N_5090);
nand U6920 (N_6920,N_5978,N_4936);
and U6921 (N_6921,N_5091,N_4962);
xnor U6922 (N_6922,N_5333,N_5050);
nand U6923 (N_6923,N_4967,N_5641);
xor U6924 (N_6924,N_5395,N_5973);
or U6925 (N_6925,N_5958,N_4812);
nor U6926 (N_6926,N_4899,N_4812);
and U6927 (N_6927,N_5692,N_5106);
and U6928 (N_6928,N_5647,N_5962);
nor U6929 (N_6929,N_5795,N_5733);
xor U6930 (N_6930,N_5186,N_5354);
xor U6931 (N_6931,N_4981,N_5944);
nand U6932 (N_6932,N_5579,N_4835);
nand U6933 (N_6933,N_5398,N_5931);
nor U6934 (N_6934,N_5678,N_5795);
nor U6935 (N_6935,N_5697,N_5373);
xor U6936 (N_6936,N_5326,N_5112);
xor U6937 (N_6937,N_4990,N_4945);
nand U6938 (N_6938,N_5528,N_5794);
nor U6939 (N_6939,N_5536,N_5205);
and U6940 (N_6940,N_5024,N_5268);
or U6941 (N_6941,N_5572,N_4801);
or U6942 (N_6942,N_5278,N_5183);
and U6943 (N_6943,N_5959,N_5667);
xnor U6944 (N_6944,N_5316,N_5381);
or U6945 (N_6945,N_5759,N_5360);
or U6946 (N_6946,N_5084,N_5656);
xnor U6947 (N_6947,N_5006,N_5220);
xnor U6948 (N_6948,N_5442,N_5717);
xor U6949 (N_6949,N_5354,N_5863);
nand U6950 (N_6950,N_5385,N_4941);
and U6951 (N_6951,N_4943,N_5352);
or U6952 (N_6952,N_5791,N_5355);
and U6953 (N_6953,N_5848,N_5317);
nand U6954 (N_6954,N_5577,N_4971);
nand U6955 (N_6955,N_5389,N_5127);
xnor U6956 (N_6956,N_5813,N_4803);
and U6957 (N_6957,N_5355,N_5693);
or U6958 (N_6958,N_5115,N_5087);
nor U6959 (N_6959,N_5814,N_5789);
nor U6960 (N_6960,N_4818,N_5902);
nand U6961 (N_6961,N_5350,N_5365);
and U6962 (N_6962,N_5197,N_5013);
and U6963 (N_6963,N_4846,N_5539);
xor U6964 (N_6964,N_5676,N_4938);
xnor U6965 (N_6965,N_5652,N_5261);
nor U6966 (N_6966,N_5144,N_5264);
and U6967 (N_6967,N_4899,N_4828);
or U6968 (N_6968,N_5548,N_5241);
or U6969 (N_6969,N_5433,N_5039);
nand U6970 (N_6970,N_4963,N_5868);
xnor U6971 (N_6971,N_5407,N_5313);
and U6972 (N_6972,N_5757,N_5965);
nor U6973 (N_6973,N_5616,N_5839);
and U6974 (N_6974,N_5436,N_5720);
nor U6975 (N_6975,N_5125,N_5182);
nand U6976 (N_6976,N_5803,N_5115);
xnor U6977 (N_6977,N_5482,N_5645);
or U6978 (N_6978,N_4957,N_5451);
and U6979 (N_6979,N_5778,N_5695);
nor U6980 (N_6980,N_5673,N_5589);
and U6981 (N_6981,N_5712,N_5306);
or U6982 (N_6982,N_5936,N_4849);
or U6983 (N_6983,N_5914,N_5073);
xnor U6984 (N_6984,N_5584,N_5131);
and U6985 (N_6985,N_5607,N_5854);
xor U6986 (N_6986,N_4964,N_5629);
xnor U6987 (N_6987,N_5805,N_5657);
or U6988 (N_6988,N_5033,N_5735);
and U6989 (N_6989,N_5619,N_5416);
and U6990 (N_6990,N_5304,N_5649);
and U6991 (N_6991,N_4818,N_5311);
and U6992 (N_6992,N_4866,N_5233);
or U6993 (N_6993,N_4802,N_5998);
nand U6994 (N_6994,N_5590,N_5137);
or U6995 (N_6995,N_5075,N_5485);
and U6996 (N_6996,N_4862,N_5079);
xnor U6997 (N_6997,N_5758,N_4935);
nand U6998 (N_6998,N_5526,N_5815);
and U6999 (N_6999,N_4882,N_5809);
nor U7000 (N_7000,N_5903,N_5800);
and U7001 (N_7001,N_5512,N_5485);
and U7002 (N_7002,N_4867,N_4861);
or U7003 (N_7003,N_5151,N_5864);
nand U7004 (N_7004,N_5924,N_5969);
nand U7005 (N_7005,N_5528,N_4976);
nor U7006 (N_7006,N_5183,N_4897);
nand U7007 (N_7007,N_5381,N_4928);
and U7008 (N_7008,N_5846,N_4871);
and U7009 (N_7009,N_5964,N_4807);
and U7010 (N_7010,N_5837,N_5625);
nor U7011 (N_7011,N_5178,N_5542);
or U7012 (N_7012,N_5856,N_5955);
nor U7013 (N_7013,N_5437,N_4856);
and U7014 (N_7014,N_5268,N_5694);
nand U7015 (N_7015,N_5087,N_5976);
xor U7016 (N_7016,N_5605,N_4944);
nand U7017 (N_7017,N_5633,N_5817);
nand U7018 (N_7018,N_5907,N_4831);
nand U7019 (N_7019,N_4948,N_5308);
nor U7020 (N_7020,N_5773,N_5441);
or U7021 (N_7021,N_5699,N_5363);
nand U7022 (N_7022,N_5101,N_5895);
and U7023 (N_7023,N_5205,N_5478);
or U7024 (N_7024,N_5235,N_5926);
and U7025 (N_7025,N_4929,N_5431);
nand U7026 (N_7026,N_5232,N_4964);
xnor U7027 (N_7027,N_5072,N_5906);
or U7028 (N_7028,N_5505,N_5726);
nor U7029 (N_7029,N_5005,N_5365);
xnor U7030 (N_7030,N_5487,N_5894);
nor U7031 (N_7031,N_5840,N_5894);
nor U7032 (N_7032,N_5076,N_5237);
xor U7033 (N_7033,N_4805,N_5838);
and U7034 (N_7034,N_5112,N_5168);
xnor U7035 (N_7035,N_5332,N_5625);
nand U7036 (N_7036,N_4911,N_4916);
or U7037 (N_7037,N_5029,N_5497);
and U7038 (N_7038,N_5499,N_5461);
xnor U7039 (N_7039,N_5471,N_5727);
or U7040 (N_7040,N_5419,N_5955);
nor U7041 (N_7041,N_5946,N_4820);
nand U7042 (N_7042,N_5947,N_5844);
nand U7043 (N_7043,N_5170,N_5776);
nor U7044 (N_7044,N_4945,N_5174);
nor U7045 (N_7045,N_4958,N_5114);
or U7046 (N_7046,N_4818,N_5931);
nor U7047 (N_7047,N_5715,N_4997);
nand U7048 (N_7048,N_5477,N_5558);
and U7049 (N_7049,N_5314,N_5571);
nor U7050 (N_7050,N_5522,N_4863);
nor U7051 (N_7051,N_5950,N_5677);
nand U7052 (N_7052,N_5950,N_5598);
and U7053 (N_7053,N_4941,N_5488);
nor U7054 (N_7054,N_4866,N_4922);
or U7055 (N_7055,N_5237,N_5523);
xor U7056 (N_7056,N_5204,N_5834);
or U7057 (N_7057,N_5675,N_5792);
or U7058 (N_7058,N_5826,N_5554);
and U7059 (N_7059,N_5649,N_5893);
and U7060 (N_7060,N_5926,N_5919);
nand U7061 (N_7061,N_5576,N_4928);
nor U7062 (N_7062,N_5696,N_5784);
nor U7063 (N_7063,N_5612,N_5712);
nand U7064 (N_7064,N_5533,N_4950);
xnor U7065 (N_7065,N_5324,N_5255);
xnor U7066 (N_7066,N_5589,N_5429);
xor U7067 (N_7067,N_5734,N_4891);
or U7068 (N_7068,N_5336,N_4920);
nor U7069 (N_7069,N_5308,N_4832);
and U7070 (N_7070,N_4967,N_4908);
or U7071 (N_7071,N_4939,N_5922);
and U7072 (N_7072,N_4882,N_4814);
xnor U7073 (N_7073,N_5198,N_5810);
nand U7074 (N_7074,N_5216,N_5829);
nand U7075 (N_7075,N_5143,N_5991);
nand U7076 (N_7076,N_5242,N_4878);
or U7077 (N_7077,N_5843,N_5453);
or U7078 (N_7078,N_5658,N_5645);
nand U7079 (N_7079,N_5446,N_4858);
xnor U7080 (N_7080,N_5251,N_5821);
xor U7081 (N_7081,N_5803,N_5303);
or U7082 (N_7082,N_5656,N_5158);
or U7083 (N_7083,N_5500,N_5546);
nor U7084 (N_7084,N_5121,N_5555);
xnor U7085 (N_7085,N_5834,N_5581);
nor U7086 (N_7086,N_5305,N_5016);
and U7087 (N_7087,N_5410,N_5630);
or U7088 (N_7088,N_5233,N_5458);
and U7089 (N_7089,N_5258,N_5241);
xor U7090 (N_7090,N_5730,N_5193);
or U7091 (N_7091,N_5510,N_5552);
or U7092 (N_7092,N_5388,N_5166);
nand U7093 (N_7093,N_5470,N_5258);
or U7094 (N_7094,N_5737,N_5717);
and U7095 (N_7095,N_4821,N_4876);
and U7096 (N_7096,N_5243,N_5432);
nor U7097 (N_7097,N_5983,N_5531);
xnor U7098 (N_7098,N_5165,N_5499);
or U7099 (N_7099,N_5052,N_5430);
xor U7100 (N_7100,N_5368,N_5101);
nor U7101 (N_7101,N_5095,N_5733);
xnor U7102 (N_7102,N_5793,N_5853);
and U7103 (N_7103,N_5548,N_5832);
and U7104 (N_7104,N_5774,N_4985);
nor U7105 (N_7105,N_4811,N_5308);
nor U7106 (N_7106,N_5700,N_5298);
nand U7107 (N_7107,N_5427,N_5239);
nor U7108 (N_7108,N_5756,N_4955);
or U7109 (N_7109,N_5843,N_5671);
nor U7110 (N_7110,N_5499,N_5620);
and U7111 (N_7111,N_5412,N_5545);
nand U7112 (N_7112,N_5325,N_5368);
nor U7113 (N_7113,N_5516,N_5522);
nor U7114 (N_7114,N_5010,N_5801);
xor U7115 (N_7115,N_5206,N_5546);
nor U7116 (N_7116,N_5158,N_5724);
or U7117 (N_7117,N_5505,N_5774);
nand U7118 (N_7118,N_5536,N_5466);
xor U7119 (N_7119,N_5161,N_5576);
and U7120 (N_7120,N_5660,N_4842);
nand U7121 (N_7121,N_5492,N_5866);
nor U7122 (N_7122,N_5682,N_5177);
nand U7123 (N_7123,N_5424,N_5669);
xnor U7124 (N_7124,N_5388,N_5850);
nand U7125 (N_7125,N_5949,N_4821);
nand U7126 (N_7126,N_5863,N_5015);
nor U7127 (N_7127,N_5069,N_5727);
xnor U7128 (N_7128,N_5584,N_5776);
nor U7129 (N_7129,N_5478,N_5021);
nand U7130 (N_7130,N_5437,N_5184);
nor U7131 (N_7131,N_4811,N_5437);
xnor U7132 (N_7132,N_5257,N_5073);
and U7133 (N_7133,N_5389,N_5300);
xnor U7134 (N_7134,N_5077,N_5628);
nor U7135 (N_7135,N_5928,N_5473);
and U7136 (N_7136,N_4942,N_5068);
nor U7137 (N_7137,N_5913,N_5311);
nand U7138 (N_7138,N_5943,N_5776);
nor U7139 (N_7139,N_5728,N_5067);
xnor U7140 (N_7140,N_5036,N_4896);
nand U7141 (N_7141,N_5097,N_5789);
nand U7142 (N_7142,N_5932,N_5886);
xor U7143 (N_7143,N_4850,N_5728);
or U7144 (N_7144,N_5523,N_5104);
and U7145 (N_7145,N_4839,N_5869);
or U7146 (N_7146,N_5671,N_5158);
or U7147 (N_7147,N_5987,N_5519);
or U7148 (N_7148,N_5827,N_5097);
xnor U7149 (N_7149,N_5436,N_5399);
nor U7150 (N_7150,N_5027,N_5329);
nor U7151 (N_7151,N_5203,N_5603);
nor U7152 (N_7152,N_5146,N_5319);
nor U7153 (N_7153,N_4876,N_5598);
nor U7154 (N_7154,N_5059,N_5011);
nand U7155 (N_7155,N_5072,N_5529);
nor U7156 (N_7156,N_5060,N_5544);
xor U7157 (N_7157,N_5140,N_5270);
nor U7158 (N_7158,N_5137,N_4882);
nor U7159 (N_7159,N_4854,N_5367);
and U7160 (N_7160,N_5648,N_4899);
or U7161 (N_7161,N_5925,N_5171);
and U7162 (N_7162,N_5007,N_5476);
nand U7163 (N_7163,N_5579,N_5683);
nor U7164 (N_7164,N_5931,N_4978);
and U7165 (N_7165,N_4840,N_5772);
and U7166 (N_7166,N_4975,N_5054);
nand U7167 (N_7167,N_5537,N_5255);
nand U7168 (N_7168,N_5416,N_5045);
nor U7169 (N_7169,N_5164,N_5688);
nand U7170 (N_7170,N_5913,N_5955);
or U7171 (N_7171,N_4992,N_4960);
nand U7172 (N_7172,N_5533,N_4801);
or U7173 (N_7173,N_4902,N_5674);
xnor U7174 (N_7174,N_4916,N_5401);
and U7175 (N_7175,N_5772,N_5967);
nor U7176 (N_7176,N_5293,N_5084);
xor U7177 (N_7177,N_5155,N_5908);
xor U7178 (N_7178,N_4870,N_4873);
nand U7179 (N_7179,N_5223,N_5957);
nand U7180 (N_7180,N_5519,N_5852);
and U7181 (N_7181,N_5535,N_5963);
xor U7182 (N_7182,N_5886,N_5035);
xor U7183 (N_7183,N_5904,N_5443);
nand U7184 (N_7184,N_4944,N_5700);
nor U7185 (N_7185,N_5152,N_4891);
or U7186 (N_7186,N_4875,N_5851);
or U7187 (N_7187,N_5440,N_5289);
xor U7188 (N_7188,N_5122,N_5435);
nand U7189 (N_7189,N_5189,N_5103);
and U7190 (N_7190,N_5872,N_5373);
nor U7191 (N_7191,N_5898,N_4965);
or U7192 (N_7192,N_5139,N_4969);
xor U7193 (N_7193,N_5898,N_5715);
or U7194 (N_7194,N_5001,N_5359);
or U7195 (N_7195,N_5462,N_5379);
nor U7196 (N_7196,N_5263,N_5013);
or U7197 (N_7197,N_4966,N_5592);
xor U7198 (N_7198,N_5624,N_5876);
nor U7199 (N_7199,N_5849,N_5376);
nand U7200 (N_7200,N_7067,N_6755);
xnor U7201 (N_7201,N_6491,N_6948);
nor U7202 (N_7202,N_7160,N_7085);
and U7203 (N_7203,N_6459,N_6537);
and U7204 (N_7204,N_6250,N_6388);
and U7205 (N_7205,N_6791,N_6690);
nor U7206 (N_7206,N_6618,N_6142);
or U7207 (N_7207,N_6958,N_6034);
nand U7208 (N_7208,N_6259,N_6538);
xnor U7209 (N_7209,N_7163,N_6296);
and U7210 (N_7210,N_6310,N_6037);
and U7211 (N_7211,N_6432,N_6545);
xor U7212 (N_7212,N_6004,N_6005);
nor U7213 (N_7213,N_6705,N_6245);
xor U7214 (N_7214,N_6743,N_7165);
nand U7215 (N_7215,N_6445,N_7097);
nand U7216 (N_7216,N_6264,N_6685);
or U7217 (N_7217,N_6756,N_6154);
or U7218 (N_7218,N_6372,N_6344);
nor U7219 (N_7219,N_6483,N_6986);
nor U7220 (N_7220,N_7025,N_6125);
xor U7221 (N_7221,N_6510,N_6455);
nand U7222 (N_7222,N_6437,N_6658);
or U7223 (N_7223,N_6373,N_6974);
nor U7224 (N_7224,N_6069,N_6908);
and U7225 (N_7225,N_6119,N_7117);
xor U7226 (N_7226,N_6914,N_6687);
nand U7227 (N_7227,N_6443,N_6744);
and U7228 (N_7228,N_7141,N_6527);
and U7229 (N_7229,N_6570,N_7140);
or U7230 (N_7230,N_7170,N_6939);
xnor U7231 (N_7231,N_6955,N_6394);
nor U7232 (N_7232,N_6674,N_6118);
or U7233 (N_7233,N_6329,N_6506);
xor U7234 (N_7234,N_6447,N_6707);
or U7235 (N_7235,N_6297,N_6286);
and U7236 (N_7236,N_6775,N_6615);
or U7237 (N_7237,N_6417,N_6068);
and U7238 (N_7238,N_6768,N_6970);
and U7239 (N_7239,N_7068,N_6151);
and U7240 (N_7240,N_6162,N_6559);
nor U7241 (N_7241,N_6608,N_6697);
nor U7242 (N_7242,N_6099,N_6196);
nand U7243 (N_7243,N_7038,N_6864);
and U7244 (N_7244,N_6623,N_6214);
or U7245 (N_7245,N_7056,N_7114);
xnor U7246 (N_7246,N_6021,N_6737);
or U7247 (N_7247,N_6924,N_6129);
nor U7248 (N_7248,N_7126,N_6513);
nand U7249 (N_7249,N_7033,N_6473);
nand U7250 (N_7250,N_6503,N_7177);
and U7251 (N_7251,N_7057,N_6035);
or U7252 (N_7252,N_6979,N_6838);
and U7253 (N_7253,N_7020,N_6255);
and U7254 (N_7254,N_6167,N_6841);
nor U7255 (N_7255,N_6633,N_6348);
nand U7256 (N_7256,N_6891,N_6702);
and U7257 (N_7257,N_6379,N_6457);
xor U7258 (N_7258,N_6141,N_6071);
xnor U7259 (N_7259,N_6689,N_7146);
nand U7260 (N_7260,N_6806,N_6391);
nand U7261 (N_7261,N_7030,N_6186);
and U7262 (N_7262,N_6507,N_6552);
or U7263 (N_7263,N_7094,N_6161);
nor U7264 (N_7264,N_6012,N_6664);
nand U7265 (N_7265,N_7148,N_6577);
nor U7266 (N_7266,N_7019,N_6486);
or U7267 (N_7267,N_6845,N_6913);
nor U7268 (N_7268,N_6518,N_6074);
or U7269 (N_7269,N_7046,N_6382);
nor U7270 (N_7270,N_6342,N_6993);
nor U7271 (N_7271,N_6801,N_6941);
and U7272 (N_7272,N_6336,N_6421);
xnor U7273 (N_7273,N_6580,N_6778);
nand U7274 (N_7274,N_6856,N_6754);
and U7275 (N_7275,N_6999,N_6758);
and U7276 (N_7276,N_6761,N_6059);
nand U7277 (N_7277,N_6399,N_6526);
xor U7278 (N_7278,N_6197,N_6370);
nor U7279 (N_7279,N_6194,N_7198);
and U7280 (N_7280,N_6848,N_6530);
and U7281 (N_7281,N_6672,N_7110);
nand U7282 (N_7282,N_6149,N_6403);
nand U7283 (N_7283,N_6456,N_6516);
and U7284 (N_7284,N_7039,N_7086);
nand U7285 (N_7285,N_6726,N_6639);
nand U7286 (N_7286,N_6077,N_6810);
nand U7287 (N_7287,N_6590,N_6277);
nor U7288 (N_7288,N_6772,N_6779);
or U7289 (N_7289,N_6681,N_6079);
nor U7290 (N_7290,N_6206,N_6086);
or U7291 (N_7291,N_6193,N_6968);
nand U7292 (N_7292,N_6102,N_6834);
nand U7293 (N_7293,N_6495,N_6216);
or U7294 (N_7294,N_6989,N_6072);
nor U7295 (N_7295,N_6635,N_6492);
nand U7296 (N_7296,N_6256,N_7109);
nor U7297 (N_7297,N_6450,N_6660);
nand U7298 (N_7298,N_6562,N_6292);
nor U7299 (N_7299,N_6897,N_6043);
nand U7300 (N_7300,N_6863,N_6797);
nand U7301 (N_7301,N_7069,N_6138);
nor U7302 (N_7302,N_6900,N_6928);
nor U7303 (N_7303,N_6606,N_6793);
xor U7304 (N_7304,N_6564,N_6667);
or U7305 (N_7305,N_7169,N_6759);
or U7306 (N_7306,N_6232,N_6578);
nand U7307 (N_7307,N_6637,N_6930);
xnor U7308 (N_7308,N_6223,N_7121);
and U7309 (N_7309,N_6422,N_6089);
nor U7310 (N_7310,N_6936,N_6610);
xnor U7311 (N_7311,N_6584,N_7051);
nor U7312 (N_7312,N_6994,N_6725);
or U7313 (N_7313,N_6877,N_6872);
nand U7314 (N_7314,N_7176,N_6740);
nand U7315 (N_7315,N_6682,N_6628);
nor U7316 (N_7316,N_6619,N_6494);
xor U7317 (N_7317,N_6460,N_6343);
and U7318 (N_7318,N_7136,N_7037);
nor U7319 (N_7319,N_6497,N_6651);
nor U7320 (N_7320,N_7096,N_6818);
xnor U7321 (N_7321,N_6082,N_6463);
nand U7322 (N_7322,N_6890,N_7042);
and U7323 (N_7323,N_6446,N_7090);
xor U7324 (N_7324,N_6056,N_6547);
or U7325 (N_7325,N_6222,N_7137);
xor U7326 (N_7326,N_6094,N_6305);
xor U7327 (N_7327,N_6829,N_7074);
and U7328 (N_7328,N_6464,N_6385);
and U7329 (N_7329,N_6550,N_6147);
xnor U7330 (N_7330,N_6183,N_6815);
and U7331 (N_7331,N_6345,N_7076);
xor U7332 (N_7332,N_6291,N_6646);
and U7333 (N_7333,N_6111,N_7027);
and U7334 (N_7334,N_6185,N_6971);
xor U7335 (N_7335,N_6231,N_6531);
nand U7336 (N_7336,N_7166,N_7159);
nor U7337 (N_7337,N_6704,N_7167);
nor U7338 (N_7338,N_6551,N_6749);
nand U7339 (N_7339,N_7082,N_6398);
xnor U7340 (N_7340,N_6662,N_6467);
xnor U7341 (N_7341,N_6716,N_7119);
nor U7342 (N_7342,N_6541,N_7129);
or U7343 (N_7343,N_6055,N_7062);
nand U7344 (N_7344,N_6107,N_6332);
nor U7345 (N_7345,N_7059,N_6881);
nand U7346 (N_7346,N_6995,N_6721);
nor U7347 (N_7347,N_6517,N_6076);
nand U7348 (N_7348,N_6224,N_7063);
and U7349 (N_7349,N_6040,N_7023);
and U7350 (N_7350,N_7111,N_6324);
nand U7351 (N_7351,N_6713,N_6790);
nor U7352 (N_7352,N_6101,N_7084);
and U7353 (N_7353,N_6925,N_6935);
nor U7354 (N_7354,N_6949,N_6670);
or U7355 (N_7355,N_6880,N_6709);
or U7356 (N_7356,N_6816,N_6299);
and U7357 (N_7357,N_6805,N_6582);
xnor U7358 (N_7358,N_6053,N_7132);
and U7359 (N_7359,N_6817,N_6006);
nand U7360 (N_7360,N_6823,N_6278);
nor U7361 (N_7361,N_6603,N_6039);
xor U7362 (N_7362,N_7006,N_6630);
nand U7363 (N_7363,N_6188,N_6252);
or U7364 (N_7364,N_6613,N_6514);
xor U7365 (N_7365,N_7104,N_6227);
xor U7366 (N_7366,N_6802,N_7026);
or U7367 (N_7367,N_7099,N_6334);
nor U7368 (N_7368,N_6712,N_6202);
nor U7369 (N_7369,N_6840,N_6532);
or U7370 (N_7370,N_7072,N_6770);
or U7371 (N_7371,N_6498,N_6504);
nor U7372 (N_7372,N_7107,N_6632);
and U7373 (N_7373,N_6990,N_6279);
xnor U7374 (N_7374,N_6352,N_6569);
or U7375 (N_7375,N_6395,N_6042);
xnor U7376 (N_7376,N_7066,N_6274);
nor U7377 (N_7377,N_6301,N_7016);
xnor U7378 (N_7378,N_7055,N_6338);
and U7379 (N_7379,N_6942,N_7183);
or U7380 (N_7380,N_6431,N_6835);
nor U7381 (N_7381,N_6905,N_6918);
nand U7382 (N_7382,N_6262,N_6475);
nor U7383 (N_7383,N_6747,N_7199);
nor U7384 (N_7384,N_6139,N_6558);
nand U7385 (N_7385,N_6548,N_6016);
nand U7386 (N_7386,N_7149,N_6060);
nand U7387 (N_7387,N_6915,N_7155);
nor U7388 (N_7388,N_6057,N_6952);
and U7389 (N_7389,N_6302,N_6380);
and U7390 (N_7390,N_7007,N_6542);
and U7391 (N_7391,N_7182,N_6170);
nand U7392 (N_7392,N_6819,N_6409);
nor U7393 (N_7393,N_7088,N_6003);
and U7394 (N_7394,N_6921,N_7049);
and U7395 (N_7395,N_6316,N_6917);
nor U7396 (N_7396,N_6397,N_6742);
nor U7397 (N_7397,N_7188,N_7075);
or U7398 (N_7398,N_6017,N_6160);
nand U7399 (N_7399,N_6937,N_6378);
or U7400 (N_7400,N_6244,N_6826);
xnor U7401 (N_7401,N_6620,N_7186);
or U7402 (N_7402,N_6782,N_6947);
xnor U7403 (N_7403,N_6462,N_6315);
or U7404 (N_7404,N_7191,N_6824);
nor U7405 (N_7405,N_6831,N_6751);
xor U7406 (N_7406,N_6307,N_6728);
and U7407 (N_7407,N_7010,N_6052);
and U7408 (N_7408,N_6317,N_6535);
xor U7409 (N_7409,N_6563,N_7180);
or U7410 (N_7410,N_6965,N_6178);
nor U7411 (N_7411,N_6466,N_6873);
nand U7412 (N_7412,N_6152,N_6238);
nand U7413 (N_7413,N_6988,N_6860);
nand U7414 (N_7414,N_6587,N_6182);
or U7415 (N_7415,N_6136,N_7053);
xnor U7416 (N_7416,N_6954,N_7179);
nand U7417 (N_7417,N_6982,N_7095);
and U7418 (N_7418,N_6127,N_6512);
or U7419 (N_7419,N_6703,N_6677);
and U7420 (N_7420,N_6389,N_7047);
xnor U7421 (N_7421,N_6258,N_6496);
or U7422 (N_7422,N_6075,N_6717);
nand U7423 (N_7423,N_7135,N_6124);
or U7424 (N_7424,N_6589,N_6083);
nor U7425 (N_7425,N_7018,N_6131);
xnor U7426 (N_7426,N_7080,N_6321);
xnor U7427 (N_7427,N_6276,N_6351);
xor U7428 (N_7428,N_6561,N_6919);
or U7429 (N_7429,N_6922,N_6521);
xor U7430 (N_7430,N_6876,N_6146);
or U7431 (N_7431,N_6493,N_6041);
nor U7432 (N_7432,N_6953,N_6711);
or U7433 (N_7433,N_7154,N_7138);
or U7434 (N_7434,N_6235,N_6522);
nor U7435 (N_7435,N_6879,N_6001);
nor U7436 (N_7436,N_7061,N_6031);
and U7437 (N_7437,N_6028,N_6275);
nor U7438 (N_7438,N_6122,N_6465);
nand U7439 (N_7439,N_7194,N_6659);
nor U7440 (N_7440,N_6842,N_6555);
xnor U7441 (N_7441,N_6416,N_7197);
nand U7442 (N_7442,N_6413,N_6789);
nor U7443 (N_7443,N_6850,N_6708);
nand U7444 (N_7444,N_7078,N_6964);
xor U7445 (N_7445,N_6368,N_6081);
xor U7446 (N_7446,N_6356,N_6354);
or U7447 (N_7447,N_6734,N_6428);
nor U7448 (N_7448,N_6715,N_6358);
nand U7449 (N_7449,N_6710,N_6427);
or U7450 (N_7450,N_7040,N_6113);
nand U7451 (N_7451,N_6172,N_6184);
nor U7452 (N_7452,N_6596,N_6412);
and U7453 (N_7453,N_6341,N_6597);
nand U7454 (N_7454,N_6500,N_6192);
or U7455 (N_7455,N_6116,N_6987);
or U7456 (N_7456,N_6696,N_6629);
or U7457 (N_7457,N_6753,N_6067);
and U7458 (N_7458,N_6218,N_6733);
or U7459 (N_7459,N_6085,N_6926);
xnor U7460 (N_7460,N_6643,N_6163);
nor U7461 (N_7461,N_7125,N_6804);
nand U7462 (N_7462,N_6836,N_6261);
xor U7463 (N_7463,N_6212,N_6866);
nor U7464 (N_7464,N_6803,N_6130);
nor U7465 (N_7465,N_6631,N_6858);
nor U7466 (N_7466,N_6731,N_6454);
nor U7467 (N_7467,N_6396,N_6406);
nor U7468 (N_7468,N_6158,N_6036);
nand U7469 (N_7469,N_6168,N_6825);
or U7470 (N_7470,N_7014,N_6911);
nand U7471 (N_7471,N_6951,N_6730);
or U7472 (N_7472,N_6963,N_6812);
nor U7473 (N_7473,N_6155,N_7131);
nor U7474 (N_7474,N_6884,N_6174);
nor U7475 (N_7475,N_6795,N_6644);
nor U7476 (N_7476,N_7113,N_6050);
or U7477 (N_7477,N_7174,N_6846);
nor U7478 (N_7478,N_6794,N_6843);
and U7479 (N_7479,N_6066,N_6273);
nand U7480 (N_7480,N_6854,N_6022);
xnor U7481 (N_7481,N_7036,N_7116);
nor U7482 (N_7482,N_6665,N_6219);
or U7483 (N_7483,N_6923,N_6785);
nor U7484 (N_7484,N_6451,N_6691);
and U7485 (N_7485,N_6407,N_6528);
xnor U7486 (N_7486,N_6833,N_6722);
or U7487 (N_7487,N_6110,N_6430);
xor U7488 (N_7488,N_7017,N_6799);
and U7489 (N_7489,N_7065,N_6909);
and U7490 (N_7490,N_6199,N_6938);
or U7491 (N_7491,N_6899,N_6080);
nand U7492 (N_7492,N_7060,N_6384);
and U7493 (N_7493,N_6047,N_6934);
and U7494 (N_7494,N_6857,N_6894);
nor U7495 (N_7495,N_6752,N_6573);
nand U7496 (N_7496,N_6969,N_6353);
or U7497 (N_7497,N_6485,N_6400);
nand U7498 (N_7498,N_6330,N_6242);
or U7499 (N_7499,N_6777,N_6870);
and U7500 (N_7500,N_6204,N_7081);
nor U7501 (N_7501,N_6706,N_6061);
or U7502 (N_7502,N_6693,N_6088);
xor U7503 (N_7503,N_6200,N_6729);
or U7504 (N_7504,N_6318,N_6191);
and U7505 (N_7505,N_7175,N_6019);
nor U7506 (N_7506,N_6673,N_6381);
or U7507 (N_7507,N_6015,N_6410);
nand U7508 (N_7508,N_6612,N_6166);
nor U7509 (N_7509,N_7127,N_6335);
xor U7510 (N_7510,N_7003,N_6807);
nor U7511 (N_7511,N_6676,N_7031);
nand U7512 (N_7512,N_7000,N_6888);
nor U7513 (N_7513,N_6977,N_6581);
xor U7514 (N_7514,N_6333,N_6616);
and U7515 (N_7515,N_6904,N_6211);
nand U7516 (N_7516,N_7112,N_6246);
or U7517 (N_7517,N_6470,N_6363);
nor U7518 (N_7518,N_6627,N_6482);
nand U7519 (N_7519,N_6675,N_6861);
and U7520 (N_7520,N_6203,N_6320);
nor U7521 (N_7521,N_6796,N_6226);
or U7522 (N_7522,N_6105,N_6414);
nand U7523 (N_7523,N_6046,N_7077);
nor U7524 (N_7524,N_6390,N_6476);
and U7525 (N_7525,N_6653,N_6362);
or U7526 (N_7526,N_6699,N_7091);
nand U7527 (N_7527,N_6018,N_6376);
xnor U7528 (N_7528,N_6134,N_7013);
nand U7529 (N_7529,N_6720,N_6121);
nand U7530 (N_7530,N_6120,N_6975);
or U7531 (N_7531,N_7064,N_7098);
and U7532 (N_7532,N_6602,N_6959);
or U7533 (N_7533,N_6903,N_6209);
xor U7534 (N_7534,N_6073,N_6750);
nor U7535 (N_7535,N_7143,N_6095);
or U7536 (N_7536,N_6985,N_6821);
nand U7537 (N_7537,N_6657,N_6221);
nor U7538 (N_7538,N_6290,N_7071);
or U7539 (N_7539,N_6966,N_6087);
nand U7540 (N_7540,N_6405,N_6489);
or U7541 (N_7541,N_6260,N_6718);
nor U7542 (N_7542,N_6383,N_6109);
and U7543 (N_7543,N_6601,N_7073);
and U7544 (N_7544,N_6453,N_6798);
nor U7545 (N_7545,N_6566,N_7008);
or U7546 (N_7546,N_6350,N_7157);
and U7547 (N_7547,N_6229,N_6640);
or U7548 (N_7548,N_6669,N_6851);
xnor U7549 (N_7549,N_6169,N_6100);
xor U7550 (N_7550,N_6940,N_6641);
nor U7551 (N_7551,N_6236,N_7173);
nor U7552 (N_7552,N_7139,N_6280);
and U7553 (N_7553,N_6666,N_6038);
nand U7554 (N_7554,N_6661,N_6401);
xnor U7555 (N_7555,N_6654,N_7058);
nand U7556 (N_7556,N_6327,N_6441);
nand U7557 (N_7557,N_6386,N_6165);
xnor U7558 (N_7558,N_6853,N_6591);
or U7559 (N_7559,N_6625,N_6474);
nand U7560 (N_7560,N_7022,N_6906);
and U7561 (N_7561,N_6123,N_6887);
nor U7562 (N_7562,N_6347,N_6240);
xnor U7563 (N_7563,N_6855,N_7128);
nand U7564 (N_7564,N_6180,N_6418);
and U7565 (N_7565,N_6254,N_6931);
nand U7566 (N_7566,N_6271,N_7134);
xnor U7567 (N_7567,N_6502,N_7041);
nand U7568 (N_7568,N_6153,N_6642);
nand U7569 (N_7569,N_6698,N_6896);
and U7570 (N_7570,N_6294,N_6668);
and U7571 (N_7571,N_6472,N_6961);
and U7572 (N_7572,N_6179,N_6108);
nor U7573 (N_7573,N_6738,N_6267);
nand U7574 (N_7574,N_6164,N_7103);
or U7575 (N_7575,N_6735,N_6839);
nor U7576 (N_7576,N_6295,N_6187);
and U7577 (N_7577,N_6800,N_6883);
nor U7578 (N_7578,N_6576,N_6852);
nor U7579 (N_7579,N_6686,N_6084);
xnor U7580 (N_7580,N_6402,N_6634);
xnor U7581 (N_7581,N_6714,N_6544);
xnor U7582 (N_7582,N_6269,N_6889);
xor U7583 (N_7583,N_6933,N_6371);
and U7584 (N_7584,N_6828,N_6478);
nand U7585 (N_7585,N_7193,N_7102);
or U7586 (N_7586,N_6013,N_7192);
xor U7587 (N_7587,N_6727,N_6063);
nand U7588 (N_7588,N_6723,N_6827);
nand U7589 (N_7589,N_6765,N_6377);
nand U7590 (N_7590,N_6792,N_7153);
or U7591 (N_7591,N_6030,N_6499);
nand U7592 (N_7592,N_6739,N_6468);
and U7593 (N_7593,N_6461,N_6878);
nor U7594 (N_7594,N_7009,N_6181);
nand U7595 (N_7595,N_6375,N_6257);
and U7596 (N_7596,N_6220,N_6306);
or U7597 (N_7597,N_6272,N_6048);
xnor U7598 (N_7598,N_6957,N_6543);
nor U7599 (N_7599,N_6189,N_7028);
nand U7600 (N_7600,N_6593,N_6239);
nor U7601 (N_7601,N_7161,N_6051);
or U7602 (N_7602,N_6869,N_7124);
nand U7603 (N_7603,N_7079,N_6679);
nor U7604 (N_7604,N_6173,N_7002);
nor U7605 (N_7605,N_6976,N_6448);
nand U7606 (N_7606,N_7151,N_6764);
xor U7607 (N_7607,N_6511,N_7012);
nand U7608 (N_7608,N_6599,N_6298);
or U7609 (N_7609,N_6215,N_6145);
xor U7610 (N_7610,N_7184,N_6359);
and U7611 (N_7611,N_6207,N_6745);
and U7612 (N_7612,N_6594,N_6984);
and U7613 (N_7613,N_7152,N_6374);
or U7614 (N_7614,N_7162,N_6732);
nor U7615 (N_7615,N_6614,N_6692);
nor U7616 (N_7616,N_6546,N_6773);
nor U7617 (N_7617,N_6871,N_6556);
xor U7618 (N_7618,N_6766,N_6103);
nor U7619 (N_7619,N_7147,N_6477);
nand U7620 (N_7620,N_6501,N_6434);
and U7621 (N_7621,N_6217,N_6268);
or U7622 (N_7622,N_6960,N_6565);
or U7623 (N_7623,N_6978,N_7122);
nor U7624 (N_7624,N_6647,N_6595);
or U7625 (N_7625,N_7144,N_6426);
and U7626 (N_7626,N_6010,N_6253);
nor U7627 (N_7627,N_6355,N_6266);
nor U7628 (N_7628,N_6519,N_6944);
nor U7629 (N_7629,N_7189,N_6655);
xor U7630 (N_7630,N_6787,N_6956);
xnor U7631 (N_7631,N_6763,N_6009);
nand U7632 (N_7632,N_6652,N_6062);
and U7633 (N_7633,N_6762,N_6190);
and U7634 (N_7634,N_6916,N_6746);
nor U7635 (N_7635,N_6780,N_6176);
and U7636 (N_7636,N_6201,N_6438);
nor U7637 (N_7637,N_6424,N_6283);
nor U7638 (N_7638,N_6104,N_7171);
nand U7639 (N_7639,N_6213,N_6748);
nand U7640 (N_7640,N_6439,N_6011);
and U7641 (N_7641,N_6621,N_7106);
xnor U7642 (N_7642,N_6932,N_6509);
nor U7643 (N_7643,N_6736,N_6319);
nor U7644 (N_7644,N_6425,N_7005);
xor U7645 (N_7645,N_6484,N_6281);
nand U7646 (N_7646,N_6487,N_6322);
and U7647 (N_7647,N_6044,N_6210);
or U7648 (N_7648,N_6490,N_6325);
or U7649 (N_7649,N_7048,N_6366);
nor U7650 (N_7650,N_6032,N_7045);
and U7651 (N_7651,N_6524,N_7001);
and U7652 (N_7652,N_6609,N_6300);
or U7653 (N_7653,N_6549,N_6263);
nor U7654 (N_7654,N_6349,N_6198);
nand U7655 (N_7655,N_6090,N_7108);
nor U7656 (N_7656,N_6536,N_6440);
or U7657 (N_7657,N_7089,N_6404);
xnor U7658 (N_7658,N_6808,N_7185);
or U7659 (N_7659,N_7145,N_6065);
or U7660 (N_7660,N_6859,N_6694);
nand U7661 (N_7661,N_7195,N_6868);
nor U7662 (N_7662,N_7050,N_6901);
or U7663 (N_7663,N_6328,N_6572);
nor U7664 (N_7664,N_6997,N_6771);
or U7665 (N_7665,N_6892,N_6156);
or U7666 (N_7666,N_6135,N_6684);
and U7667 (N_7667,N_6249,N_6205);
nor U7668 (N_7668,N_6649,N_7100);
xor U7669 (N_7669,N_6093,N_7190);
xnor U7670 (N_7670,N_6568,N_6023);
or U7671 (N_7671,N_7092,N_6811);
xor U7672 (N_7672,N_6867,N_6064);
or U7673 (N_7673,N_6907,N_6420);
or U7674 (N_7674,N_7044,N_6137);
and U7675 (N_7675,N_6678,N_6814);
or U7676 (N_7676,N_6505,N_6605);
xnor U7677 (N_7677,N_7181,N_6567);
nor U7678 (N_7678,N_6600,N_6479);
or U7679 (N_7679,N_6337,N_6049);
nor U7680 (N_7680,N_7004,N_6645);
or U7681 (N_7681,N_6973,N_6893);
xnor U7682 (N_7682,N_6361,N_6525);
and U7683 (N_7683,N_7093,N_6444);
or U7684 (N_7684,N_6289,N_6683);
nor U7685 (N_7685,N_7052,N_6045);
and U7686 (N_7686,N_6774,N_6981);
xor U7687 (N_7687,N_7158,N_6784);
nand U7688 (N_7688,N_6326,N_6106);
and U7689 (N_7689,N_6874,N_7133);
or U7690 (N_7690,N_6419,N_6837);
nand U7691 (N_7691,N_7070,N_6027);
or U7692 (N_7692,N_6323,N_6574);
and U7693 (N_7693,N_6607,N_6885);
nor U7694 (N_7694,N_6533,N_6962);
nor U7695 (N_7695,N_6304,N_6025);
and U7696 (N_7696,N_6636,N_6515);
and U7697 (N_7697,N_6387,N_6225);
nor U7698 (N_7698,N_6054,N_6847);
nand U7699 (N_7699,N_6508,N_6767);
xnor U7700 (N_7700,N_6688,N_6007);
xor U7701 (N_7701,N_6002,N_6534);
or U7702 (N_7702,N_6912,N_6622);
nand U7703 (N_7703,N_6996,N_6140);
and U7704 (N_7704,N_6776,N_7130);
nand U7705 (N_7705,N_6592,N_6862);
xor U7706 (N_7706,N_6875,N_6442);
and U7707 (N_7707,N_6849,N_6098);
nand U7708 (N_7708,N_6171,N_6458);
and U7709 (N_7709,N_6014,N_6331);
nor U7710 (N_7710,N_6029,N_6671);
or U7711 (N_7711,N_6312,N_6367);
and U7712 (N_7712,N_6126,N_6150);
and U7713 (N_7713,N_6243,N_6365);
nor U7714 (N_7714,N_6809,N_6364);
nor U7715 (N_7715,N_7172,N_6540);
nor U7716 (N_7716,N_6781,N_6314);
xnor U7717 (N_7717,N_7021,N_7120);
and U7718 (N_7718,N_6339,N_7115);
or U7719 (N_7719,N_6423,N_6133);
xnor U7720 (N_7720,N_6539,N_6346);
nor U7721 (N_7721,N_7087,N_6309);
xor U7722 (N_7722,N_6436,N_6719);
nand U7723 (N_7723,N_6265,N_6992);
nor U7724 (N_7724,N_6251,N_6950);
nor U7725 (N_7725,N_6557,N_6411);
xor U7726 (N_7726,N_6293,N_6820);
xor U7727 (N_7727,N_6991,N_6143);
nand U7728 (N_7728,N_6132,N_6270);
nand U7729 (N_7729,N_6695,N_6757);
xor U7730 (N_7730,N_6741,N_6844);
nand U7731 (N_7731,N_6488,N_6117);
nor U7732 (N_7732,N_7187,N_6284);
xnor U7733 (N_7733,N_6026,N_6783);
or U7734 (N_7734,N_6234,N_6241);
xnor U7735 (N_7735,N_6638,N_7123);
or U7736 (N_7736,N_6865,N_6096);
or U7737 (N_7737,N_6020,N_6583);
nand U7738 (N_7738,N_6929,N_7043);
nor U7739 (N_7739,N_6128,N_6760);
or U7740 (N_7740,N_6033,N_6313);
or U7741 (N_7741,N_7034,N_7015);
nand U7742 (N_7742,N_6175,N_6115);
nand U7743 (N_7743,N_7142,N_6920);
and U7744 (N_7744,N_7101,N_6148);
nand U7745 (N_7745,N_6228,N_6700);
or U7746 (N_7746,N_6701,N_6480);
or U7747 (N_7747,N_6788,N_7032);
nand U7748 (N_7748,N_6946,N_6972);
or U7749 (N_7749,N_6288,N_6481);
nor U7750 (N_7750,N_6617,N_6248);
or U7751 (N_7751,N_6469,N_6998);
nor U7752 (N_7752,N_6575,N_6680);
nand U7753 (N_7753,N_6650,N_6311);
and U7754 (N_7754,N_6247,N_6392);
or U7755 (N_7755,N_7011,N_6433);
nand U7756 (N_7756,N_6097,N_7024);
nor U7757 (N_7757,N_6452,N_6832);
or U7758 (N_7758,N_6000,N_6611);
xor U7759 (N_7759,N_6091,N_6624);
and U7760 (N_7760,N_6285,N_7164);
nand U7761 (N_7761,N_6895,N_6769);
nor U7762 (N_7762,N_6598,N_6282);
xnor U7763 (N_7763,N_7156,N_6571);
nand U7764 (N_7764,N_6070,N_6980);
nor U7765 (N_7765,N_6114,N_6553);
or U7766 (N_7766,N_6588,N_6579);
nor U7767 (N_7767,N_7150,N_6024);
or U7768 (N_7768,N_7168,N_6177);
nand U7769 (N_7769,N_6435,N_6663);
nor U7770 (N_7770,N_6983,N_6092);
or U7771 (N_7771,N_6078,N_6340);
xnor U7772 (N_7772,N_6360,N_6554);
or U7773 (N_7773,N_6886,N_7178);
xnor U7774 (N_7774,N_6112,N_6058);
and U7775 (N_7775,N_7196,N_6648);
and U7776 (N_7776,N_6560,N_6357);
nor U7777 (N_7777,N_6429,N_6230);
and U7778 (N_7778,N_6303,N_6523);
xor U7779 (N_7779,N_6626,N_6471);
xor U7780 (N_7780,N_6786,N_6945);
nor U7781 (N_7781,N_6830,N_6415);
xnor U7782 (N_7782,N_7035,N_6159);
xnor U7783 (N_7783,N_6393,N_6529);
xor U7784 (N_7784,N_6237,N_6656);
xnor U7785 (N_7785,N_7105,N_6195);
nor U7786 (N_7786,N_7083,N_6208);
or U7787 (N_7787,N_6408,N_6822);
nor U7788 (N_7788,N_6585,N_6157);
or U7789 (N_7789,N_6287,N_6520);
and U7790 (N_7790,N_7029,N_7054);
nor U7791 (N_7791,N_6008,N_6144);
nand U7792 (N_7792,N_6449,N_6902);
nor U7793 (N_7793,N_6967,N_6882);
nor U7794 (N_7794,N_6586,N_6813);
and U7795 (N_7795,N_6724,N_6308);
nor U7796 (N_7796,N_6369,N_6910);
or U7797 (N_7797,N_6604,N_6927);
and U7798 (N_7798,N_6898,N_7118);
or U7799 (N_7799,N_6233,N_6943);
nand U7800 (N_7800,N_6627,N_6691);
or U7801 (N_7801,N_6881,N_6270);
or U7802 (N_7802,N_7127,N_6983);
xnor U7803 (N_7803,N_6405,N_6368);
and U7804 (N_7804,N_6880,N_6122);
xor U7805 (N_7805,N_6709,N_6464);
and U7806 (N_7806,N_6674,N_6091);
and U7807 (N_7807,N_6402,N_6926);
and U7808 (N_7808,N_6029,N_6188);
or U7809 (N_7809,N_6159,N_7053);
xor U7810 (N_7810,N_6751,N_6091);
and U7811 (N_7811,N_6812,N_7047);
nor U7812 (N_7812,N_6992,N_6430);
nor U7813 (N_7813,N_6480,N_6576);
xor U7814 (N_7814,N_7043,N_6123);
nor U7815 (N_7815,N_6515,N_6949);
nor U7816 (N_7816,N_6091,N_6773);
or U7817 (N_7817,N_6479,N_6339);
xnor U7818 (N_7818,N_6372,N_6206);
xor U7819 (N_7819,N_6727,N_7125);
and U7820 (N_7820,N_6517,N_6992);
and U7821 (N_7821,N_6631,N_6379);
or U7822 (N_7822,N_6387,N_6767);
or U7823 (N_7823,N_6895,N_6403);
xor U7824 (N_7824,N_7082,N_7076);
nor U7825 (N_7825,N_6219,N_6384);
xor U7826 (N_7826,N_6666,N_6132);
xor U7827 (N_7827,N_7086,N_6653);
nor U7828 (N_7828,N_6836,N_6699);
xnor U7829 (N_7829,N_6912,N_6883);
and U7830 (N_7830,N_6909,N_6421);
xnor U7831 (N_7831,N_6378,N_6584);
and U7832 (N_7832,N_6933,N_6281);
nor U7833 (N_7833,N_7029,N_6610);
nand U7834 (N_7834,N_6345,N_7017);
or U7835 (N_7835,N_6007,N_6841);
or U7836 (N_7836,N_6062,N_7169);
nand U7837 (N_7837,N_6293,N_6393);
nand U7838 (N_7838,N_6769,N_7179);
nand U7839 (N_7839,N_6513,N_7037);
nor U7840 (N_7840,N_6618,N_6670);
nand U7841 (N_7841,N_6338,N_6699);
xnor U7842 (N_7842,N_6976,N_6895);
and U7843 (N_7843,N_7162,N_6374);
or U7844 (N_7844,N_6144,N_6215);
xnor U7845 (N_7845,N_6315,N_6433);
nor U7846 (N_7846,N_6821,N_6430);
nand U7847 (N_7847,N_6389,N_6442);
or U7848 (N_7848,N_6327,N_6268);
nor U7849 (N_7849,N_7042,N_7017);
nor U7850 (N_7850,N_6150,N_6192);
nand U7851 (N_7851,N_6567,N_7103);
nand U7852 (N_7852,N_7152,N_6189);
or U7853 (N_7853,N_6836,N_6163);
nor U7854 (N_7854,N_6134,N_6266);
or U7855 (N_7855,N_6155,N_6014);
and U7856 (N_7856,N_6993,N_6490);
xor U7857 (N_7857,N_6367,N_6999);
nand U7858 (N_7858,N_6130,N_6992);
and U7859 (N_7859,N_6693,N_6230);
nor U7860 (N_7860,N_6972,N_6855);
or U7861 (N_7861,N_6156,N_6721);
or U7862 (N_7862,N_7192,N_6162);
nand U7863 (N_7863,N_6294,N_7124);
and U7864 (N_7864,N_7141,N_7061);
or U7865 (N_7865,N_6335,N_6127);
nand U7866 (N_7866,N_6991,N_6119);
nor U7867 (N_7867,N_7192,N_6829);
or U7868 (N_7868,N_6372,N_6731);
nor U7869 (N_7869,N_6242,N_6176);
and U7870 (N_7870,N_6318,N_6837);
or U7871 (N_7871,N_6646,N_6429);
xor U7872 (N_7872,N_6913,N_6401);
nor U7873 (N_7873,N_6427,N_6021);
nand U7874 (N_7874,N_6122,N_6613);
nor U7875 (N_7875,N_6330,N_7110);
and U7876 (N_7876,N_6917,N_7171);
nor U7877 (N_7877,N_6314,N_6841);
and U7878 (N_7878,N_6999,N_6941);
nand U7879 (N_7879,N_6513,N_6508);
xnor U7880 (N_7880,N_7118,N_6084);
nor U7881 (N_7881,N_6664,N_6067);
nor U7882 (N_7882,N_7105,N_6527);
nor U7883 (N_7883,N_7195,N_6639);
nor U7884 (N_7884,N_6322,N_6158);
and U7885 (N_7885,N_6220,N_6974);
nor U7886 (N_7886,N_6600,N_6499);
and U7887 (N_7887,N_6204,N_6870);
xor U7888 (N_7888,N_6916,N_6390);
nor U7889 (N_7889,N_6860,N_6529);
nor U7890 (N_7890,N_6625,N_6129);
or U7891 (N_7891,N_6709,N_6786);
nor U7892 (N_7892,N_6021,N_6091);
and U7893 (N_7893,N_6177,N_6765);
nand U7894 (N_7894,N_7026,N_6484);
nor U7895 (N_7895,N_6123,N_6299);
and U7896 (N_7896,N_7185,N_6613);
nand U7897 (N_7897,N_7173,N_6241);
and U7898 (N_7898,N_7027,N_6508);
nor U7899 (N_7899,N_6807,N_7118);
nand U7900 (N_7900,N_7159,N_7176);
and U7901 (N_7901,N_6198,N_6418);
nor U7902 (N_7902,N_6549,N_6816);
and U7903 (N_7903,N_6042,N_6076);
xnor U7904 (N_7904,N_6802,N_6113);
xnor U7905 (N_7905,N_6798,N_6161);
and U7906 (N_7906,N_6296,N_6889);
or U7907 (N_7907,N_7170,N_6883);
and U7908 (N_7908,N_6352,N_7093);
xnor U7909 (N_7909,N_7002,N_6965);
and U7910 (N_7910,N_6490,N_6453);
and U7911 (N_7911,N_6106,N_6980);
and U7912 (N_7912,N_6040,N_6404);
xor U7913 (N_7913,N_6401,N_7158);
and U7914 (N_7914,N_6929,N_6862);
xnor U7915 (N_7915,N_6471,N_7094);
or U7916 (N_7916,N_6499,N_7179);
nor U7917 (N_7917,N_6927,N_6889);
and U7918 (N_7918,N_6635,N_6819);
or U7919 (N_7919,N_6718,N_6633);
nor U7920 (N_7920,N_7041,N_6592);
nand U7921 (N_7921,N_6988,N_6024);
and U7922 (N_7922,N_6076,N_6037);
xnor U7923 (N_7923,N_6670,N_7159);
and U7924 (N_7924,N_6357,N_7010);
and U7925 (N_7925,N_6091,N_6167);
or U7926 (N_7926,N_6137,N_7023);
or U7927 (N_7927,N_7193,N_6457);
and U7928 (N_7928,N_6747,N_6230);
xnor U7929 (N_7929,N_6419,N_6803);
xnor U7930 (N_7930,N_6370,N_6825);
xor U7931 (N_7931,N_6342,N_6466);
nand U7932 (N_7932,N_6818,N_6559);
nand U7933 (N_7933,N_6000,N_6480);
and U7934 (N_7934,N_6159,N_6285);
or U7935 (N_7935,N_6617,N_6622);
xnor U7936 (N_7936,N_7088,N_6942);
nand U7937 (N_7937,N_6524,N_6478);
nand U7938 (N_7938,N_7000,N_7106);
nor U7939 (N_7939,N_6095,N_6838);
nor U7940 (N_7940,N_6461,N_6524);
or U7941 (N_7941,N_6521,N_6287);
nand U7942 (N_7942,N_6574,N_7103);
nor U7943 (N_7943,N_6994,N_6670);
nor U7944 (N_7944,N_6415,N_6567);
and U7945 (N_7945,N_7112,N_6636);
and U7946 (N_7946,N_6042,N_6459);
xnor U7947 (N_7947,N_6186,N_6512);
xnor U7948 (N_7948,N_6635,N_6599);
or U7949 (N_7949,N_6390,N_6299);
nor U7950 (N_7950,N_7068,N_6730);
nor U7951 (N_7951,N_6956,N_6822);
nand U7952 (N_7952,N_6962,N_7038);
nor U7953 (N_7953,N_6944,N_6323);
xnor U7954 (N_7954,N_6924,N_6693);
nor U7955 (N_7955,N_6295,N_6944);
xnor U7956 (N_7956,N_6619,N_6291);
nand U7957 (N_7957,N_6865,N_7088);
or U7958 (N_7958,N_6126,N_6614);
nor U7959 (N_7959,N_6977,N_6415);
nand U7960 (N_7960,N_7120,N_7088);
nor U7961 (N_7961,N_7085,N_6031);
or U7962 (N_7962,N_7180,N_6051);
or U7963 (N_7963,N_6282,N_6487);
or U7964 (N_7964,N_7086,N_6689);
nand U7965 (N_7965,N_6622,N_6270);
nand U7966 (N_7966,N_6908,N_6129);
and U7967 (N_7967,N_6077,N_6005);
xnor U7968 (N_7968,N_7159,N_6553);
or U7969 (N_7969,N_6566,N_6527);
and U7970 (N_7970,N_6516,N_6842);
nor U7971 (N_7971,N_6066,N_6434);
or U7972 (N_7972,N_6757,N_6228);
and U7973 (N_7973,N_6890,N_6578);
nand U7974 (N_7974,N_6454,N_6571);
xor U7975 (N_7975,N_6865,N_7017);
or U7976 (N_7976,N_6639,N_7076);
nor U7977 (N_7977,N_6996,N_6166);
and U7978 (N_7978,N_6115,N_6196);
xor U7979 (N_7979,N_6910,N_6043);
nor U7980 (N_7980,N_6796,N_6175);
nand U7981 (N_7981,N_6900,N_6873);
xnor U7982 (N_7982,N_6685,N_6625);
and U7983 (N_7983,N_6307,N_6184);
or U7984 (N_7984,N_6109,N_6973);
and U7985 (N_7985,N_6401,N_6076);
and U7986 (N_7986,N_6388,N_6725);
nand U7987 (N_7987,N_6216,N_6050);
nand U7988 (N_7988,N_6607,N_6029);
or U7989 (N_7989,N_7111,N_6016);
nand U7990 (N_7990,N_6806,N_6886);
xor U7991 (N_7991,N_6979,N_6656);
nor U7992 (N_7992,N_6622,N_6698);
nand U7993 (N_7993,N_7006,N_6038);
nand U7994 (N_7994,N_6585,N_6190);
or U7995 (N_7995,N_6545,N_6802);
nand U7996 (N_7996,N_7153,N_6102);
and U7997 (N_7997,N_6011,N_6184);
nand U7998 (N_7998,N_6644,N_6117);
xnor U7999 (N_7999,N_6903,N_6333);
nor U8000 (N_8000,N_6922,N_6641);
nor U8001 (N_8001,N_6592,N_6473);
xnor U8002 (N_8002,N_6167,N_6615);
nor U8003 (N_8003,N_6923,N_6842);
and U8004 (N_8004,N_6715,N_6637);
or U8005 (N_8005,N_6681,N_7188);
or U8006 (N_8006,N_7144,N_6853);
nand U8007 (N_8007,N_6243,N_6982);
and U8008 (N_8008,N_6645,N_6278);
nand U8009 (N_8009,N_6872,N_6886);
xor U8010 (N_8010,N_6122,N_6809);
xor U8011 (N_8011,N_6913,N_6359);
xnor U8012 (N_8012,N_6777,N_6847);
xor U8013 (N_8013,N_6049,N_7190);
nand U8014 (N_8014,N_6812,N_6490);
nor U8015 (N_8015,N_6014,N_6716);
nor U8016 (N_8016,N_6992,N_6086);
nor U8017 (N_8017,N_6041,N_6391);
nand U8018 (N_8018,N_6228,N_7175);
xor U8019 (N_8019,N_6966,N_6770);
and U8020 (N_8020,N_6692,N_7083);
nor U8021 (N_8021,N_7133,N_6571);
nor U8022 (N_8022,N_6013,N_6319);
nor U8023 (N_8023,N_6010,N_7130);
and U8024 (N_8024,N_6192,N_6110);
nor U8025 (N_8025,N_6316,N_6350);
nand U8026 (N_8026,N_6533,N_6310);
nand U8027 (N_8027,N_6773,N_7031);
or U8028 (N_8028,N_7038,N_6268);
xnor U8029 (N_8029,N_7083,N_7158);
or U8030 (N_8030,N_6737,N_6517);
xor U8031 (N_8031,N_6712,N_6721);
xnor U8032 (N_8032,N_6719,N_6758);
xor U8033 (N_8033,N_6659,N_6290);
xnor U8034 (N_8034,N_6642,N_6442);
nand U8035 (N_8035,N_6554,N_6250);
or U8036 (N_8036,N_6900,N_6872);
and U8037 (N_8037,N_6142,N_6755);
nand U8038 (N_8038,N_6090,N_7007);
and U8039 (N_8039,N_6310,N_7001);
or U8040 (N_8040,N_6208,N_6913);
or U8041 (N_8041,N_7091,N_6319);
or U8042 (N_8042,N_6923,N_6292);
nand U8043 (N_8043,N_6756,N_6669);
nand U8044 (N_8044,N_6461,N_7195);
and U8045 (N_8045,N_6827,N_6062);
and U8046 (N_8046,N_6765,N_6188);
or U8047 (N_8047,N_6537,N_6474);
xnor U8048 (N_8048,N_6022,N_6159);
nor U8049 (N_8049,N_6541,N_6718);
or U8050 (N_8050,N_6353,N_6165);
nor U8051 (N_8051,N_6291,N_6634);
or U8052 (N_8052,N_6242,N_6299);
xor U8053 (N_8053,N_6183,N_6627);
nor U8054 (N_8054,N_6411,N_6100);
nor U8055 (N_8055,N_6658,N_6297);
and U8056 (N_8056,N_7163,N_6619);
nor U8057 (N_8057,N_6358,N_6169);
or U8058 (N_8058,N_6496,N_7171);
or U8059 (N_8059,N_6762,N_7183);
and U8060 (N_8060,N_6077,N_6418);
or U8061 (N_8061,N_6583,N_6464);
nor U8062 (N_8062,N_6433,N_6425);
nor U8063 (N_8063,N_6652,N_7184);
nand U8064 (N_8064,N_6972,N_6341);
and U8065 (N_8065,N_6496,N_6419);
nor U8066 (N_8066,N_6779,N_6990);
or U8067 (N_8067,N_6981,N_6897);
and U8068 (N_8068,N_6258,N_6740);
xor U8069 (N_8069,N_7146,N_7114);
xor U8070 (N_8070,N_6462,N_6341);
nor U8071 (N_8071,N_6295,N_6103);
nand U8072 (N_8072,N_6052,N_6013);
xor U8073 (N_8073,N_6714,N_7192);
xnor U8074 (N_8074,N_6648,N_6922);
xnor U8075 (N_8075,N_6280,N_6014);
or U8076 (N_8076,N_6036,N_6787);
xor U8077 (N_8077,N_7076,N_7166);
xor U8078 (N_8078,N_6335,N_6700);
nand U8079 (N_8079,N_7148,N_6425);
xor U8080 (N_8080,N_6747,N_7154);
nor U8081 (N_8081,N_6791,N_6426);
nand U8082 (N_8082,N_6341,N_6374);
nor U8083 (N_8083,N_6385,N_6355);
nor U8084 (N_8084,N_7059,N_6253);
and U8085 (N_8085,N_6399,N_6589);
or U8086 (N_8086,N_6877,N_6532);
nor U8087 (N_8087,N_7193,N_6911);
or U8088 (N_8088,N_7169,N_7010);
xor U8089 (N_8089,N_6055,N_7183);
nand U8090 (N_8090,N_6807,N_6866);
nor U8091 (N_8091,N_6825,N_6378);
or U8092 (N_8092,N_6024,N_6440);
or U8093 (N_8093,N_6489,N_7103);
or U8094 (N_8094,N_7088,N_6392);
xor U8095 (N_8095,N_6886,N_6905);
nand U8096 (N_8096,N_7073,N_6632);
nand U8097 (N_8097,N_6777,N_6667);
nand U8098 (N_8098,N_6555,N_6692);
or U8099 (N_8099,N_7070,N_6007);
nand U8100 (N_8100,N_7115,N_6086);
xor U8101 (N_8101,N_6604,N_7184);
nor U8102 (N_8102,N_6326,N_6840);
or U8103 (N_8103,N_6152,N_6552);
xor U8104 (N_8104,N_6288,N_6045);
nand U8105 (N_8105,N_7058,N_6509);
nand U8106 (N_8106,N_6271,N_6813);
or U8107 (N_8107,N_6764,N_6411);
or U8108 (N_8108,N_6253,N_6693);
xor U8109 (N_8109,N_6389,N_6695);
nor U8110 (N_8110,N_6645,N_6789);
or U8111 (N_8111,N_6781,N_6518);
or U8112 (N_8112,N_6579,N_6136);
xor U8113 (N_8113,N_6788,N_7175);
nor U8114 (N_8114,N_6009,N_7165);
and U8115 (N_8115,N_6891,N_6578);
nor U8116 (N_8116,N_6646,N_6573);
nand U8117 (N_8117,N_6474,N_6379);
nand U8118 (N_8118,N_6566,N_7038);
nor U8119 (N_8119,N_6602,N_6245);
or U8120 (N_8120,N_6712,N_6374);
nor U8121 (N_8121,N_6453,N_6762);
or U8122 (N_8122,N_6898,N_6807);
xnor U8123 (N_8123,N_6598,N_6963);
and U8124 (N_8124,N_7190,N_6717);
and U8125 (N_8125,N_6561,N_6139);
or U8126 (N_8126,N_6000,N_6330);
xnor U8127 (N_8127,N_6240,N_6336);
nor U8128 (N_8128,N_6520,N_6664);
and U8129 (N_8129,N_7009,N_6706);
or U8130 (N_8130,N_6204,N_6132);
xnor U8131 (N_8131,N_6572,N_6862);
nor U8132 (N_8132,N_6555,N_6595);
nand U8133 (N_8133,N_6372,N_7046);
and U8134 (N_8134,N_6038,N_6395);
nand U8135 (N_8135,N_6743,N_6035);
and U8136 (N_8136,N_6494,N_6042);
nor U8137 (N_8137,N_6317,N_6809);
and U8138 (N_8138,N_6580,N_6824);
or U8139 (N_8139,N_6993,N_7013);
xnor U8140 (N_8140,N_6832,N_6820);
xor U8141 (N_8141,N_7033,N_7163);
nor U8142 (N_8142,N_6006,N_7098);
and U8143 (N_8143,N_7190,N_6589);
nor U8144 (N_8144,N_6605,N_6580);
nor U8145 (N_8145,N_6522,N_6621);
nand U8146 (N_8146,N_6520,N_6683);
xor U8147 (N_8147,N_6232,N_6354);
nand U8148 (N_8148,N_6039,N_7051);
nand U8149 (N_8149,N_6458,N_6490);
nor U8150 (N_8150,N_6246,N_6374);
and U8151 (N_8151,N_6074,N_6066);
and U8152 (N_8152,N_6543,N_6091);
xnor U8153 (N_8153,N_6911,N_6029);
and U8154 (N_8154,N_6156,N_6731);
nor U8155 (N_8155,N_6135,N_6354);
nand U8156 (N_8156,N_7021,N_6951);
or U8157 (N_8157,N_6057,N_7191);
nor U8158 (N_8158,N_6378,N_6587);
or U8159 (N_8159,N_6943,N_6983);
nor U8160 (N_8160,N_6034,N_6448);
or U8161 (N_8161,N_6278,N_6035);
or U8162 (N_8162,N_6101,N_6311);
xnor U8163 (N_8163,N_6122,N_6906);
or U8164 (N_8164,N_6763,N_7168);
nor U8165 (N_8165,N_6657,N_6304);
or U8166 (N_8166,N_6865,N_6779);
xnor U8167 (N_8167,N_6693,N_6709);
nand U8168 (N_8168,N_6958,N_6564);
or U8169 (N_8169,N_7022,N_6598);
nand U8170 (N_8170,N_6403,N_6900);
xor U8171 (N_8171,N_6297,N_6571);
xnor U8172 (N_8172,N_7117,N_7025);
xor U8173 (N_8173,N_6819,N_6937);
nand U8174 (N_8174,N_6156,N_6817);
nand U8175 (N_8175,N_6762,N_6805);
nor U8176 (N_8176,N_6429,N_7021);
nand U8177 (N_8177,N_6795,N_7006);
xor U8178 (N_8178,N_6258,N_6662);
nand U8179 (N_8179,N_6157,N_6493);
or U8180 (N_8180,N_6243,N_6730);
or U8181 (N_8181,N_6339,N_6899);
or U8182 (N_8182,N_6606,N_6751);
nor U8183 (N_8183,N_6932,N_6910);
and U8184 (N_8184,N_7194,N_6276);
nand U8185 (N_8185,N_6728,N_6053);
or U8186 (N_8186,N_6165,N_6371);
and U8187 (N_8187,N_6270,N_6238);
or U8188 (N_8188,N_7046,N_6388);
nor U8189 (N_8189,N_6722,N_6183);
nor U8190 (N_8190,N_6504,N_6929);
or U8191 (N_8191,N_6889,N_6612);
nor U8192 (N_8192,N_6075,N_6142);
or U8193 (N_8193,N_6936,N_6461);
nand U8194 (N_8194,N_6714,N_6308);
xnor U8195 (N_8195,N_6511,N_6609);
nand U8196 (N_8196,N_7063,N_6920);
xor U8197 (N_8197,N_6953,N_6658);
nand U8198 (N_8198,N_7101,N_6486);
nand U8199 (N_8199,N_7016,N_6909);
or U8200 (N_8200,N_7120,N_6456);
and U8201 (N_8201,N_6865,N_6316);
nand U8202 (N_8202,N_6644,N_7171);
xor U8203 (N_8203,N_6942,N_6015);
xnor U8204 (N_8204,N_6182,N_6455);
xor U8205 (N_8205,N_6694,N_6145);
or U8206 (N_8206,N_6630,N_7152);
xnor U8207 (N_8207,N_6394,N_6281);
nor U8208 (N_8208,N_6134,N_6396);
nor U8209 (N_8209,N_6221,N_6725);
and U8210 (N_8210,N_6211,N_6830);
nand U8211 (N_8211,N_6669,N_6822);
nor U8212 (N_8212,N_7045,N_6165);
nor U8213 (N_8213,N_6312,N_6162);
xor U8214 (N_8214,N_6467,N_6731);
nor U8215 (N_8215,N_6226,N_6243);
or U8216 (N_8216,N_6359,N_6533);
nor U8217 (N_8217,N_7131,N_6025);
xor U8218 (N_8218,N_6301,N_6540);
nor U8219 (N_8219,N_6706,N_6450);
nand U8220 (N_8220,N_6552,N_6108);
and U8221 (N_8221,N_6758,N_6398);
nand U8222 (N_8222,N_6237,N_6781);
nand U8223 (N_8223,N_6220,N_7060);
xnor U8224 (N_8224,N_6795,N_6500);
nand U8225 (N_8225,N_7119,N_6129);
nand U8226 (N_8226,N_6666,N_6530);
or U8227 (N_8227,N_6610,N_6513);
nand U8228 (N_8228,N_6006,N_6598);
or U8229 (N_8229,N_6166,N_6983);
or U8230 (N_8230,N_7152,N_6955);
and U8231 (N_8231,N_6150,N_6152);
xnor U8232 (N_8232,N_6077,N_6096);
nor U8233 (N_8233,N_6141,N_6955);
and U8234 (N_8234,N_6148,N_6207);
nand U8235 (N_8235,N_6492,N_6151);
nor U8236 (N_8236,N_6105,N_6769);
nor U8237 (N_8237,N_7197,N_6691);
xnor U8238 (N_8238,N_6516,N_6046);
nor U8239 (N_8239,N_6067,N_7190);
xor U8240 (N_8240,N_6382,N_6350);
nor U8241 (N_8241,N_7072,N_7004);
and U8242 (N_8242,N_6649,N_6766);
and U8243 (N_8243,N_6015,N_7031);
or U8244 (N_8244,N_7024,N_6957);
or U8245 (N_8245,N_6998,N_7063);
xor U8246 (N_8246,N_6791,N_6859);
or U8247 (N_8247,N_6147,N_6893);
nand U8248 (N_8248,N_7027,N_7039);
nand U8249 (N_8249,N_6785,N_6471);
and U8250 (N_8250,N_7121,N_6989);
xnor U8251 (N_8251,N_6797,N_7101);
nor U8252 (N_8252,N_6595,N_6756);
and U8253 (N_8253,N_6442,N_6035);
or U8254 (N_8254,N_6592,N_6728);
nand U8255 (N_8255,N_6379,N_6802);
nand U8256 (N_8256,N_6836,N_6567);
nor U8257 (N_8257,N_7192,N_7043);
and U8258 (N_8258,N_6449,N_6662);
nand U8259 (N_8259,N_6356,N_6592);
and U8260 (N_8260,N_6178,N_6650);
nor U8261 (N_8261,N_6243,N_6925);
or U8262 (N_8262,N_6880,N_6649);
or U8263 (N_8263,N_6050,N_6743);
xnor U8264 (N_8264,N_6748,N_6219);
nand U8265 (N_8265,N_6601,N_6094);
nand U8266 (N_8266,N_6460,N_6483);
nand U8267 (N_8267,N_6437,N_6131);
and U8268 (N_8268,N_6375,N_6484);
nand U8269 (N_8269,N_7052,N_7157);
nor U8270 (N_8270,N_6671,N_6487);
nand U8271 (N_8271,N_6727,N_6831);
nand U8272 (N_8272,N_6776,N_6312);
xnor U8273 (N_8273,N_6043,N_6067);
and U8274 (N_8274,N_6968,N_6507);
and U8275 (N_8275,N_6772,N_6590);
nor U8276 (N_8276,N_6153,N_6797);
xnor U8277 (N_8277,N_6318,N_6525);
and U8278 (N_8278,N_6917,N_6067);
and U8279 (N_8279,N_7022,N_6454);
nand U8280 (N_8280,N_6340,N_6012);
and U8281 (N_8281,N_6912,N_6499);
nand U8282 (N_8282,N_7015,N_6939);
nor U8283 (N_8283,N_6948,N_6143);
and U8284 (N_8284,N_6656,N_6446);
nand U8285 (N_8285,N_6463,N_6820);
and U8286 (N_8286,N_6428,N_6367);
nor U8287 (N_8287,N_6730,N_6394);
xnor U8288 (N_8288,N_6741,N_6085);
or U8289 (N_8289,N_6608,N_6193);
nor U8290 (N_8290,N_6236,N_6242);
nand U8291 (N_8291,N_6928,N_6013);
xnor U8292 (N_8292,N_6856,N_6303);
or U8293 (N_8293,N_6239,N_7106);
nor U8294 (N_8294,N_7125,N_6744);
nand U8295 (N_8295,N_6582,N_6472);
nor U8296 (N_8296,N_6969,N_6927);
nor U8297 (N_8297,N_6343,N_6976);
and U8298 (N_8298,N_6454,N_6374);
xnor U8299 (N_8299,N_6980,N_6088);
xnor U8300 (N_8300,N_6359,N_6165);
nand U8301 (N_8301,N_6856,N_6272);
nor U8302 (N_8302,N_6712,N_7096);
nor U8303 (N_8303,N_7115,N_6100);
nand U8304 (N_8304,N_7002,N_6255);
or U8305 (N_8305,N_6068,N_7099);
nor U8306 (N_8306,N_6561,N_6557);
nor U8307 (N_8307,N_6933,N_6495);
and U8308 (N_8308,N_6898,N_7190);
nor U8309 (N_8309,N_6023,N_6916);
and U8310 (N_8310,N_6732,N_6027);
nor U8311 (N_8311,N_6728,N_6692);
or U8312 (N_8312,N_6966,N_6011);
and U8313 (N_8313,N_6918,N_6797);
or U8314 (N_8314,N_6370,N_7029);
xnor U8315 (N_8315,N_7080,N_6746);
nor U8316 (N_8316,N_6168,N_6290);
xor U8317 (N_8317,N_7002,N_6565);
xnor U8318 (N_8318,N_6458,N_6397);
nand U8319 (N_8319,N_6343,N_6361);
nor U8320 (N_8320,N_7120,N_6735);
and U8321 (N_8321,N_6789,N_6177);
or U8322 (N_8322,N_7141,N_6706);
nor U8323 (N_8323,N_7155,N_6131);
nand U8324 (N_8324,N_6364,N_6700);
nand U8325 (N_8325,N_6499,N_6362);
and U8326 (N_8326,N_7052,N_6570);
nand U8327 (N_8327,N_6536,N_6056);
or U8328 (N_8328,N_6417,N_6137);
nor U8329 (N_8329,N_6944,N_6783);
nor U8330 (N_8330,N_7130,N_6955);
nor U8331 (N_8331,N_6696,N_6736);
or U8332 (N_8332,N_6323,N_6955);
xor U8333 (N_8333,N_6506,N_6331);
nand U8334 (N_8334,N_6196,N_6289);
and U8335 (N_8335,N_6571,N_6252);
xor U8336 (N_8336,N_6127,N_6306);
or U8337 (N_8337,N_6536,N_6064);
and U8338 (N_8338,N_6443,N_6501);
or U8339 (N_8339,N_6947,N_6245);
xnor U8340 (N_8340,N_6428,N_6317);
or U8341 (N_8341,N_6758,N_6231);
and U8342 (N_8342,N_6907,N_6868);
nor U8343 (N_8343,N_6016,N_6514);
nand U8344 (N_8344,N_6246,N_6300);
or U8345 (N_8345,N_6941,N_6888);
and U8346 (N_8346,N_6106,N_6440);
and U8347 (N_8347,N_6289,N_6392);
or U8348 (N_8348,N_7161,N_6555);
and U8349 (N_8349,N_6430,N_6280);
nor U8350 (N_8350,N_6076,N_6539);
nor U8351 (N_8351,N_6448,N_7137);
nor U8352 (N_8352,N_6192,N_6897);
or U8353 (N_8353,N_6205,N_6718);
and U8354 (N_8354,N_6125,N_6198);
xor U8355 (N_8355,N_6097,N_6661);
xor U8356 (N_8356,N_6831,N_7051);
or U8357 (N_8357,N_6001,N_7001);
nor U8358 (N_8358,N_6127,N_7131);
xor U8359 (N_8359,N_6817,N_7091);
nand U8360 (N_8360,N_6192,N_7195);
nor U8361 (N_8361,N_7169,N_6114);
xor U8362 (N_8362,N_6291,N_6339);
nand U8363 (N_8363,N_6943,N_6292);
nor U8364 (N_8364,N_7086,N_6005);
nand U8365 (N_8365,N_6273,N_6602);
nor U8366 (N_8366,N_6632,N_6055);
nand U8367 (N_8367,N_6605,N_6699);
and U8368 (N_8368,N_6433,N_6466);
xnor U8369 (N_8369,N_6414,N_6205);
nor U8370 (N_8370,N_6257,N_6384);
or U8371 (N_8371,N_6046,N_6125);
and U8372 (N_8372,N_6983,N_6522);
nand U8373 (N_8373,N_6952,N_6685);
and U8374 (N_8374,N_6701,N_6691);
nor U8375 (N_8375,N_6923,N_6729);
or U8376 (N_8376,N_6600,N_6101);
xnor U8377 (N_8377,N_6465,N_6625);
or U8378 (N_8378,N_6694,N_6366);
nand U8379 (N_8379,N_6259,N_6463);
and U8380 (N_8380,N_6471,N_6708);
or U8381 (N_8381,N_6167,N_6821);
nand U8382 (N_8382,N_6936,N_6914);
nand U8383 (N_8383,N_6757,N_6011);
and U8384 (N_8384,N_6928,N_6120);
and U8385 (N_8385,N_6000,N_6950);
nor U8386 (N_8386,N_6287,N_6917);
or U8387 (N_8387,N_6134,N_6537);
xnor U8388 (N_8388,N_6944,N_6706);
xnor U8389 (N_8389,N_6342,N_6908);
nand U8390 (N_8390,N_7072,N_6662);
nand U8391 (N_8391,N_7040,N_6728);
nand U8392 (N_8392,N_7103,N_7054);
nand U8393 (N_8393,N_6294,N_6351);
and U8394 (N_8394,N_6896,N_6845);
xnor U8395 (N_8395,N_6535,N_6746);
nand U8396 (N_8396,N_6133,N_6921);
and U8397 (N_8397,N_6156,N_6530);
and U8398 (N_8398,N_6971,N_6094);
and U8399 (N_8399,N_6013,N_6246);
nand U8400 (N_8400,N_8060,N_7268);
xor U8401 (N_8401,N_8294,N_7245);
nor U8402 (N_8402,N_7593,N_8343);
xor U8403 (N_8403,N_7940,N_7666);
nor U8404 (N_8404,N_8164,N_7614);
xnor U8405 (N_8405,N_7461,N_8175);
nand U8406 (N_8406,N_7440,N_7348);
nor U8407 (N_8407,N_8150,N_7454);
nand U8408 (N_8408,N_7627,N_7618);
nand U8409 (N_8409,N_7744,N_7356);
and U8410 (N_8410,N_8006,N_7370);
or U8411 (N_8411,N_7222,N_7916);
and U8412 (N_8412,N_7248,N_7223);
or U8413 (N_8413,N_7216,N_7421);
xnor U8414 (N_8414,N_7570,N_7922);
nand U8415 (N_8415,N_7761,N_7901);
nor U8416 (N_8416,N_8316,N_8122);
nand U8417 (N_8417,N_7990,N_7637);
nor U8418 (N_8418,N_7366,N_7480);
and U8419 (N_8419,N_7986,N_7798);
nand U8420 (N_8420,N_7596,N_7684);
nor U8421 (N_8421,N_7620,N_7696);
nand U8422 (N_8422,N_7908,N_8033);
nor U8423 (N_8423,N_7927,N_8095);
nor U8424 (N_8424,N_8102,N_8183);
nand U8425 (N_8425,N_7260,N_8074);
or U8426 (N_8426,N_7415,N_8010);
and U8427 (N_8427,N_8121,N_7210);
or U8428 (N_8428,N_7401,N_7318);
and U8429 (N_8429,N_8061,N_8073);
nor U8430 (N_8430,N_7780,N_7668);
nor U8431 (N_8431,N_7595,N_7544);
xor U8432 (N_8432,N_7285,N_7450);
and U8433 (N_8433,N_7751,N_7388);
and U8434 (N_8434,N_8237,N_8177);
or U8435 (N_8435,N_8200,N_7592);
nor U8436 (N_8436,N_8382,N_7675);
nand U8437 (N_8437,N_8390,N_7951);
nor U8438 (N_8438,N_7509,N_8236);
nand U8439 (N_8439,N_8002,N_8340);
nand U8440 (N_8440,N_7293,N_8182);
and U8441 (N_8441,N_8344,N_7969);
or U8442 (N_8442,N_7612,N_7770);
and U8443 (N_8443,N_8181,N_8101);
nand U8444 (N_8444,N_8328,N_7959);
xnor U8445 (N_8445,N_7453,N_8283);
and U8446 (N_8446,N_7532,N_7385);
xnor U8447 (N_8447,N_8051,N_8077);
nand U8448 (N_8448,N_7903,N_7205);
nand U8449 (N_8449,N_7995,N_7752);
or U8450 (N_8450,N_7670,N_7275);
and U8451 (N_8451,N_8373,N_7781);
and U8452 (N_8452,N_7869,N_7563);
xor U8453 (N_8453,N_8362,N_7267);
xor U8454 (N_8454,N_7811,N_7204);
and U8455 (N_8455,N_8109,N_7394);
nand U8456 (N_8456,N_8368,N_8337);
and U8457 (N_8457,N_7526,N_7561);
or U8458 (N_8458,N_7419,N_7554);
xor U8459 (N_8459,N_7296,N_7452);
and U8460 (N_8460,N_7760,N_8364);
nor U8461 (N_8461,N_8313,N_7409);
or U8462 (N_8462,N_7517,N_8085);
or U8463 (N_8463,N_8205,N_7674);
xor U8464 (N_8464,N_8072,N_7954);
and U8465 (N_8465,N_7469,N_8385);
nand U8466 (N_8466,N_8046,N_7791);
nor U8467 (N_8467,N_7771,N_8090);
xnor U8468 (N_8468,N_8219,N_8172);
xnor U8469 (N_8469,N_7395,N_7787);
xor U8470 (N_8470,N_8030,N_8124);
xnor U8471 (N_8471,N_8015,N_7573);
xnor U8472 (N_8472,N_7477,N_7436);
xor U8473 (N_8473,N_7322,N_8342);
or U8474 (N_8474,N_7432,N_7439);
and U8475 (N_8475,N_7937,N_7442);
and U8476 (N_8476,N_7513,N_7677);
nand U8477 (N_8477,N_8230,N_7699);
or U8478 (N_8478,N_8055,N_7747);
nand U8479 (N_8479,N_7556,N_7690);
and U8480 (N_8480,N_7806,N_7819);
nor U8481 (N_8481,N_7785,N_7582);
xor U8482 (N_8482,N_8217,N_8301);
and U8483 (N_8483,N_8377,N_7730);
nor U8484 (N_8484,N_7283,N_7257);
and U8485 (N_8485,N_7343,N_7514);
nand U8486 (N_8486,N_7705,N_7769);
nand U8487 (N_8487,N_7736,N_8036);
nand U8488 (N_8488,N_7843,N_8207);
and U8489 (N_8489,N_7557,N_7217);
nor U8490 (N_8490,N_8267,N_7971);
nand U8491 (N_8491,N_7307,N_8174);
and U8492 (N_8492,N_7655,N_7679);
xor U8493 (N_8493,N_7202,N_7324);
xnor U8494 (N_8494,N_8140,N_7498);
nor U8495 (N_8495,N_7535,N_7817);
or U8496 (N_8496,N_7816,N_8263);
nor U8497 (N_8497,N_7979,N_8176);
or U8498 (N_8498,N_8312,N_7465);
xnor U8499 (N_8499,N_7212,N_8013);
xor U8500 (N_8500,N_7938,N_7398);
nor U8501 (N_8501,N_7972,N_7414);
nor U8502 (N_8502,N_7528,N_8078);
nand U8503 (N_8503,N_7422,N_7815);
and U8504 (N_8504,N_7200,N_7594);
and U8505 (N_8505,N_7209,N_8096);
or U8506 (N_8506,N_7659,N_8037);
nor U8507 (N_8507,N_8031,N_7968);
and U8508 (N_8508,N_8380,N_8272);
and U8509 (N_8509,N_7287,N_7728);
or U8510 (N_8510,N_8024,N_8259);
or U8511 (N_8511,N_7788,N_7871);
nor U8512 (N_8512,N_7255,N_8323);
or U8513 (N_8513,N_7753,N_7634);
xnor U8514 (N_8514,N_8163,N_7224);
xnor U8515 (N_8515,N_7221,N_7387);
and U8516 (N_8516,N_7338,N_8304);
or U8517 (N_8517,N_8022,N_8376);
or U8518 (N_8518,N_7958,N_8159);
and U8519 (N_8519,N_8322,N_8381);
or U8520 (N_8520,N_7404,N_8238);
and U8521 (N_8521,N_7720,N_8370);
xnor U8522 (N_8522,N_8110,N_7349);
xor U8523 (N_8523,N_7763,N_8201);
nand U8524 (N_8524,N_7591,N_7575);
nor U8525 (N_8525,N_8224,N_7650);
and U8526 (N_8526,N_7397,N_7369);
nand U8527 (N_8527,N_7892,N_7966);
xor U8528 (N_8528,N_8225,N_7604);
nor U8529 (N_8529,N_7437,N_7578);
xor U8530 (N_8530,N_7360,N_8288);
and U8531 (N_8531,N_7352,N_8129);
and U8532 (N_8532,N_7802,N_8114);
xor U8533 (N_8533,N_8251,N_7295);
nand U8534 (N_8534,N_7831,N_7213);
and U8535 (N_8535,N_7332,N_7503);
or U8536 (N_8536,N_8116,N_8011);
nand U8537 (N_8537,N_8269,N_8395);
nor U8538 (N_8538,N_8320,N_8143);
and U8539 (N_8539,N_7839,N_7701);
and U8540 (N_8540,N_7632,N_7873);
xnor U8541 (N_8541,N_7717,N_8093);
or U8542 (N_8542,N_7206,N_7269);
or U8543 (N_8543,N_8026,N_7740);
or U8544 (N_8544,N_7837,N_8260);
and U8545 (N_8545,N_8356,N_8324);
or U8546 (N_8546,N_7625,N_8311);
and U8547 (N_8547,N_7896,N_7499);
nand U8548 (N_8548,N_7842,N_7820);
xor U8549 (N_8549,N_8048,N_8349);
xor U8550 (N_8550,N_7691,N_7628);
nor U8551 (N_8551,N_7776,N_8128);
and U8552 (N_8552,N_7587,N_7361);
or U8553 (N_8553,N_7365,N_8388);
nor U8554 (N_8554,N_7919,N_8123);
nor U8555 (N_8555,N_7658,N_7247);
nand U8556 (N_8556,N_8242,N_7645);
and U8557 (N_8557,N_7639,N_8084);
and U8558 (N_8558,N_7660,N_7722);
nor U8559 (N_8559,N_7803,N_7235);
or U8560 (N_8560,N_7396,N_7610);
or U8561 (N_8561,N_8346,N_7836);
or U8562 (N_8562,N_7400,N_8218);
xor U8563 (N_8563,N_7755,N_8321);
xnor U8564 (N_8564,N_7850,N_7790);
nand U8565 (N_8565,N_7708,N_7764);
and U8566 (N_8566,N_8397,N_8276);
and U8567 (N_8567,N_8042,N_8020);
or U8568 (N_8568,N_7227,N_7795);
nand U8569 (N_8569,N_7801,N_8229);
and U8570 (N_8570,N_7583,N_7765);
and U8571 (N_8571,N_8087,N_8384);
and U8572 (N_8572,N_8365,N_7965);
or U8573 (N_8573,N_8266,N_7417);
xor U8574 (N_8574,N_8299,N_7832);
and U8575 (N_8575,N_7962,N_7783);
nor U8576 (N_8576,N_8287,N_7520);
and U8577 (N_8577,N_8393,N_7881);
and U8578 (N_8578,N_7997,N_8047);
xor U8579 (N_8579,N_7451,N_7784);
or U8580 (N_8580,N_7928,N_7745);
nor U8581 (N_8581,N_8155,N_8392);
and U8582 (N_8582,N_8310,N_7447);
nor U8583 (N_8583,N_7600,N_8290);
xor U8584 (N_8584,N_7923,N_7553);
nand U8585 (N_8585,N_7250,N_7762);
or U8586 (N_8586,N_7518,N_7462);
and U8587 (N_8587,N_7493,N_7229);
xor U8588 (N_8588,N_7936,N_7303);
or U8589 (N_8589,N_7737,N_7813);
or U8590 (N_8590,N_8043,N_7921);
and U8591 (N_8591,N_7256,N_8035);
and U8592 (N_8592,N_7848,N_7571);
or U8593 (N_8593,N_8070,N_8147);
nand U8594 (N_8594,N_8091,N_7527);
xor U8595 (N_8595,N_7363,N_7516);
nand U8596 (N_8596,N_7719,N_7758);
nand U8597 (N_8597,N_7335,N_8248);
nor U8598 (N_8598,N_7818,N_7569);
or U8599 (N_8599,N_8001,N_7925);
xor U8600 (N_8600,N_7512,N_7642);
nor U8601 (N_8601,N_7987,N_7471);
nor U8602 (N_8602,N_7550,N_7624);
nor U8603 (N_8603,N_8179,N_7314);
and U8604 (N_8604,N_7441,N_8256);
nand U8605 (N_8605,N_8214,N_7767);
or U8606 (N_8606,N_7808,N_7555);
xor U8607 (N_8607,N_7852,N_7716);
or U8608 (N_8608,N_7799,N_8394);
or U8609 (N_8609,N_7605,N_8160);
xnor U8610 (N_8610,N_8071,N_7264);
nand U8611 (N_8611,N_7431,N_8187);
and U8612 (N_8612,N_7733,N_7663);
nand U8613 (N_8613,N_8165,N_8371);
xor U8614 (N_8614,N_7756,N_7685);
and U8615 (N_8615,N_8297,N_7495);
or U8616 (N_8616,N_7941,N_7738);
or U8617 (N_8617,N_7702,N_7904);
nand U8618 (N_8618,N_8080,N_7239);
and U8619 (N_8619,N_7992,N_8277);
xnor U8620 (N_8620,N_7226,N_7282);
nor U8621 (N_8621,N_7304,N_7463);
and U8622 (N_8622,N_7861,N_7960);
and U8623 (N_8623,N_8271,N_7757);
nand U8624 (N_8624,N_8327,N_7934);
nor U8625 (N_8625,N_7621,N_7615);
or U8626 (N_8626,N_8148,N_7312);
and U8627 (N_8627,N_7878,N_7931);
nor U8628 (N_8628,N_7597,N_8076);
nor U8629 (N_8629,N_7448,N_8314);
nor U8630 (N_8630,N_7266,N_8292);
nor U8631 (N_8631,N_8386,N_7866);
xor U8632 (N_8632,N_8223,N_7492);
or U8633 (N_8633,N_7218,N_7497);
nor U8634 (N_8634,N_7609,N_7698);
nand U8635 (N_8635,N_8049,N_7484);
or U8636 (N_8636,N_7262,N_7487);
nor U8637 (N_8637,N_7598,N_7862);
xor U8638 (N_8638,N_7888,N_7301);
nor U8639 (N_8639,N_8065,N_8054);
or U8640 (N_8640,N_7891,N_7644);
nor U8641 (N_8641,N_7502,N_7917);
and U8642 (N_8642,N_7510,N_8202);
xnor U8643 (N_8643,N_8298,N_8185);
xnor U8644 (N_8644,N_8359,N_8246);
nor U8645 (N_8645,N_7809,N_7464);
or U8646 (N_8646,N_8302,N_7629);
xor U8647 (N_8647,N_7270,N_8142);
and U8648 (N_8648,N_7589,N_7623);
or U8649 (N_8649,N_8039,N_7542);
xnor U8650 (N_8650,N_7434,N_7723);
and U8651 (N_8651,N_7297,N_7418);
xnor U8652 (N_8652,N_7983,N_7576);
and U8653 (N_8653,N_8088,N_8336);
xor U8654 (N_8654,N_8106,N_7508);
nor U8655 (N_8655,N_8389,N_7661);
nor U8656 (N_8656,N_7333,N_7633);
nand U8657 (N_8657,N_8156,N_7898);
or U8658 (N_8658,N_8232,N_7856);
nor U8659 (N_8659,N_7294,N_7534);
or U8660 (N_8660,N_8146,N_7251);
xor U8661 (N_8661,N_8190,N_7299);
xor U8662 (N_8662,N_7559,N_7608);
xnor U8663 (N_8663,N_8289,N_7219);
xor U8664 (N_8664,N_8153,N_8097);
xnor U8665 (N_8665,N_7244,N_7793);
xor U8666 (N_8666,N_7680,N_8107);
and U8667 (N_8667,N_7329,N_8012);
xor U8668 (N_8668,N_8058,N_7313);
nand U8669 (N_8669,N_7883,N_8396);
and U8670 (N_8670,N_7796,N_7689);
nor U8671 (N_8671,N_7841,N_7511);
or U8672 (N_8672,N_7910,N_7496);
nor U8673 (N_8673,N_8014,N_7252);
xor U8674 (N_8674,N_8358,N_7727);
xor U8675 (N_8675,N_7773,N_7697);
nor U8676 (N_8676,N_7725,N_7789);
nor U8677 (N_8677,N_8045,N_7380);
or U8678 (N_8678,N_8275,N_7443);
and U8679 (N_8679,N_8333,N_8341);
xnor U8680 (N_8680,N_7807,N_7676);
xor U8681 (N_8681,N_8166,N_8279);
or U8682 (N_8682,N_7649,N_7868);
xor U8683 (N_8683,N_7834,N_7641);
nor U8684 (N_8684,N_7426,N_7741);
xor U8685 (N_8685,N_8374,N_7900);
xnor U8686 (N_8686,N_7838,N_7468);
xor U8687 (N_8687,N_7585,N_7336);
and U8688 (N_8688,N_8038,N_7408);
or U8689 (N_8689,N_7371,N_8119);
xnor U8690 (N_8690,N_8169,N_7353);
xor U8691 (N_8691,N_7444,N_7412);
nor U8692 (N_8692,N_7884,N_7522);
nand U8693 (N_8693,N_7999,N_8303);
xnor U8694 (N_8694,N_8353,N_7631);
nand U8695 (N_8695,N_8258,N_7381);
and U8696 (N_8696,N_7549,N_8383);
nand U8697 (N_8697,N_7375,N_7427);
and U8698 (N_8698,N_8352,N_7800);
xor U8699 (N_8699,N_7291,N_7607);
nor U8700 (N_8700,N_8239,N_7721);
nor U8701 (N_8701,N_7746,N_7918);
and U8702 (N_8702,N_7693,N_7358);
xor U8703 (N_8703,N_7930,N_8135);
nor U8704 (N_8704,N_8211,N_7331);
nand U8705 (N_8705,N_7568,N_8268);
xnor U8706 (N_8706,N_7538,N_7671);
nand U8707 (N_8707,N_8145,N_7488);
xor U8708 (N_8708,N_7935,N_7709);
nor U8709 (N_8709,N_8329,N_7779);
nand U8710 (N_8710,N_8008,N_7970);
and U8711 (N_8711,N_7909,N_7870);
nand U8712 (N_8712,N_7286,N_7533);
or U8713 (N_8713,N_7963,N_8189);
nor U8714 (N_8714,N_8162,N_8332);
xnor U8715 (N_8715,N_8180,N_8355);
nor U8716 (N_8716,N_8184,N_7984);
and U8717 (N_8717,N_7232,N_7695);
and U8718 (N_8718,N_7377,N_7616);
and U8719 (N_8719,N_7759,N_7390);
and U8720 (N_8720,N_7383,N_7207);
and U8721 (N_8721,N_7413,N_7425);
and U8722 (N_8722,N_7606,N_8305);
and U8723 (N_8723,N_7327,N_7265);
or U8724 (N_8724,N_7867,N_7749);
nor U8725 (N_8725,N_7473,N_8300);
or U8726 (N_8726,N_7334,N_7777);
xor U8727 (N_8727,N_7630,N_7998);
nor U8728 (N_8728,N_7411,N_7367);
or U8729 (N_8729,N_8228,N_7686);
and U8730 (N_8730,N_7640,N_7302);
nand U8731 (N_8731,N_7424,N_7812);
and U8732 (N_8732,N_8139,N_7638);
nand U8733 (N_8733,N_7500,N_7678);
nand U8734 (N_8734,N_7662,N_7912);
nand U8735 (N_8735,N_7466,N_7967);
nor U8736 (N_8736,N_8378,N_8204);
nand U8737 (N_8737,N_7844,N_7420);
xnor U8738 (N_8738,N_7525,N_7920);
nor U8739 (N_8739,N_7483,N_7316);
or U8740 (N_8740,N_7234,N_7459);
xor U8741 (N_8741,N_7939,N_7306);
and U8742 (N_8742,N_7775,N_7249);
or U8743 (N_8743,N_7961,N_7539);
nor U8744 (N_8744,N_7300,N_7545);
and U8745 (N_8745,N_7849,N_8278);
and U8746 (N_8746,N_7321,N_7687);
nor U8747 (N_8747,N_7399,N_7455);
nor U8748 (N_8748,N_7259,N_7855);
and U8749 (N_8749,N_8104,N_7541);
xnor U8750 (N_8750,N_7305,N_8210);
nor U8751 (N_8751,N_7991,N_8209);
and U8752 (N_8752,N_7731,N_8168);
or U8753 (N_8753,N_7292,N_7272);
xor U8754 (N_8754,N_8326,N_7362);
nor U8755 (N_8755,N_7797,N_8089);
nand U8756 (N_8756,N_7238,N_8354);
nand U8757 (N_8757,N_8379,N_7794);
nor U8758 (N_8758,N_7208,N_7735);
nor U8759 (N_8759,N_7964,N_7956);
nor U8760 (N_8760,N_7330,N_8363);
nor U8761 (N_8761,N_7824,N_7449);
or U8762 (N_8762,N_7847,N_8032);
nand U8763 (N_8763,N_7902,N_8003);
nand U8764 (N_8764,N_7558,N_7393);
or U8765 (N_8765,N_7364,N_7643);
or U8766 (N_8766,N_7458,N_7858);
or U8767 (N_8767,N_7707,N_7368);
xnor U8768 (N_8768,N_7669,N_7289);
and U8769 (N_8769,N_7882,N_8206);
or U8770 (N_8770,N_7985,N_7810);
and U8771 (N_8771,N_7233,N_7475);
nor U8772 (N_8772,N_7948,N_7308);
nand U8773 (N_8773,N_7851,N_8317);
or U8774 (N_8774,N_7344,N_8137);
and U8775 (N_8775,N_8281,N_8199);
and U8776 (N_8776,N_7590,N_8173);
xnor U8777 (N_8777,N_8094,N_7263);
xor U8778 (N_8778,N_8021,N_7872);
or U8779 (N_8779,N_7237,N_7976);
xnor U8780 (N_8780,N_8103,N_8132);
and U8781 (N_8781,N_7519,N_7230);
nand U8782 (N_8782,N_7750,N_7402);
nor U8783 (N_8783,N_7635,N_8118);
or U8784 (N_8784,N_7531,N_8331);
and U8785 (N_8785,N_7565,N_8027);
xor U8786 (N_8786,N_8309,N_8375);
or U8787 (N_8787,N_8138,N_7828);
nand U8788 (N_8788,N_8348,N_7537);
xor U8789 (N_8789,N_7281,N_7996);
nand U8790 (N_8790,N_7485,N_7506);
and U8791 (N_8791,N_7552,N_7899);
xnor U8792 (N_8792,N_8192,N_7864);
and U8793 (N_8793,N_7253,N_8064);
xnor U8794 (N_8794,N_8215,N_8330);
xnor U8795 (N_8795,N_7258,N_7857);
xnor U8796 (N_8796,N_7543,N_7350);
xor U8797 (N_8797,N_7949,N_7376);
or U8798 (N_8798,N_7656,N_8082);
and U8799 (N_8799,N_7374,N_8361);
nand U8800 (N_8800,N_8282,N_8068);
xnor U8801 (N_8801,N_7271,N_7739);
xor U8802 (N_8802,N_7284,N_8170);
nand U8803 (N_8803,N_7830,N_7490);
nor U8804 (N_8804,N_8178,N_7924);
and U8805 (N_8805,N_8391,N_7672);
xor U8806 (N_8806,N_8034,N_8280);
xnor U8807 (N_8807,N_8351,N_8018);
and U8808 (N_8808,N_8167,N_8325);
xor U8809 (N_8809,N_7584,N_7667);
and U8810 (N_8810,N_7827,N_7613);
nor U8811 (N_8811,N_7586,N_7724);
xnor U8812 (N_8812,N_7340,N_7505);
or U8813 (N_8813,N_7865,N_7973);
or U8814 (N_8814,N_8108,N_7579);
and U8815 (N_8815,N_8334,N_7386);
or U8816 (N_8816,N_7470,N_7472);
nor U8817 (N_8817,N_8235,N_7913);
nor U8818 (N_8818,N_7201,N_7845);
or U8819 (N_8819,N_7907,N_7435);
nor U8820 (N_8820,N_8157,N_8273);
nand U8821 (N_8821,N_7540,N_7982);
or U8822 (N_8822,N_8100,N_7885);
and U8823 (N_8823,N_7860,N_7391);
xor U8824 (N_8824,N_7354,N_7276);
or U8825 (N_8825,N_7599,N_7994);
or U8826 (N_8826,N_7430,N_7489);
nor U8827 (N_8827,N_7405,N_7880);
nor U8828 (N_8828,N_8253,N_8345);
and U8829 (N_8829,N_8366,N_7863);
nor U8830 (N_8830,N_7246,N_7562);
or U8831 (N_8831,N_7372,N_7311);
and U8832 (N_8832,N_7228,N_7407);
and U8833 (N_8833,N_7890,N_8113);
nor U8834 (N_8834,N_7974,N_7236);
and U8835 (N_8835,N_8291,N_7309);
nand U8836 (N_8836,N_7905,N_7476);
or U8837 (N_8837,N_8062,N_8293);
nor U8838 (N_8838,N_7345,N_7482);
or U8839 (N_8839,N_7273,N_7786);
or U8840 (N_8840,N_7945,N_8050);
and U8841 (N_8841,N_7879,N_8262);
and U8842 (N_8842,N_7357,N_8264);
nand U8843 (N_8843,N_8105,N_7942);
or U8844 (N_8844,N_8117,N_8339);
nor U8845 (N_8845,N_7242,N_7339);
or U8846 (N_8846,N_7700,N_7341);
and U8847 (N_8847,N_8086,N_7714);
nand U8848 (N_8848,N_7748,N_7530);
and U8849 (N_8849,N_8149,N_8231);
and U8850 (N_8850,N_8194,N_7854);
xor U8851 (N_8851,N_8357,N_7822);
and U8852 (N_8852,N_7328,N_8227);
or U8853 (N_8853,N_7766,N_7220);
nor U8854 (N_8854,N_8040,N_7529);
nand U8855 (N_8855,N_8240,N_7564);
and U8856 (N_8856,N_7946,N_7280);
nor U8857 (N_8857,N_7524,N_7551);
or U8858 (N_8858,N_7840,N_8274);
xor U8859 (N_8859,N_7782,N_7378);
or U8860 (N_8860,N_7325,N_7243);
and U8861 (N_8861,N_7950,N_7603);
nor U8862 (N_8862,N_7768,N_7955);
and U8863 (N_8863,N_8296,N_7647);
nor U8864 (N_8864,N_7211,N_8220);
xor U8865 (N_8865,N_8133,N_7975);
or U8866 (N_8866,N_7887,N_7536);
xnor U8867 (N_8867,N_7874,N_7980);
and U8868 (N_8868,N_7467,N_7479);
or U8869 (N_8869,N_7710,N_7823);
xor U8870 (N_8870,N_7320,N_8053);
and U8871 (N_8871,N_7428,N_8112);
or U8872 (N_8872,N_7754,N_7929);
nand U8873 (N_8873,N_7894,N_7711);
xnor U8874 (N_8874,N_7989,N_7826);
xor U8875 (N_8875,N_7392,N_7893);
and U8876 (N_8876,N_7445,N_7682);
or U8877 (N_8877,N_7486,N_8398);
nand U8878 (N_8878,N_7581,N_8136);
nand U8879 (N_8879,N_7792,N_7403);
or U8880 (N_8880,N_8284,N_7317);
xor U8881 (N_8881,N_7337,N_7410);
or U8882 (N_8882,N_7298,N_8007);
nand U8883 (N_8883,N_7384,N_7914);
nand U8884 (N_8884,N_8241,N_8261);
or U8885 (N_8885,N_8234,N_7947);
xor U8886 (N_8886,N_8017,N_7566);
xor U8887 (N_8887,N_8216,N_7713);
or U8888 (N_8888,N_7665,N_8052);
or U8889 (N_8889,N_7277,N_7704);
nor U8890 (N_8890,N_8069,N_7580);
nand U8891 (N_8891,N_7351,N_8127);
nor U8892 (N_8892,N_7743,N_7821);
xnor U8893 (N_8893,N_8196,N_8295);
xnor U8894 (N_8894,N_7619,N_7829);
nand U8895 (N_8895,N_7261,N_7895);
nor U8896 (N_8896,N_7932,N_8000);
and U8897 (N_8897,N_7323,N_7588);
nor U8898 (N_8898,N_7859,N_8099);
nand U8899 (N_8899,N_8250,N_7481);
nor U8900 (N_8900,N_7772,N_8360);
nand U8901 (N_8901,N_7523,N_7952);
xor U8902 (N_8902,N_7651,N_8023);
nor U8903 (N_8903,N_8092,N_8115);
or U8904 (N_8904,N_7636,N_7474);
xnor U8905 (N_8905,N_7359,N_7977);
xor U8906 (N_8906,N_8347,N_7933);
and U8907 (N_8907,N_8029,N_8212);
nand U8908 (N_8908,N_8213,N_7648);
or U8909 (N_8909,N_8016,N_7491);
and U8910 (N_8910,N_7373,N_7617);
nor U8911 (N_8911,N_8252,N_8233);
xnor U8912 (N_8912,N_8255,N_8126);
or U8913 (N_8913,N_7214,N_7897);
xor U8914 (N_8914,N_8083,N_8198);
or U8915 (N_8915,N_7915,N_8152);
and U8916 (N_8916,N_8285,N_7876);
or U8917 (N_8917,N_8221,N_7981);
nand U8918 (N_8918,N_8120,N_8203);
nor U8919 (N_8919,N_8191,N_7572);
xnor U8920 (N_8920,N_8208,N_7423);
nand U8921 (N_8921,N_8131,N_7547);
or U8922 (N_8922,N_8245,N_7877);
nand U8923 (N_8923,N_8247,N_7521);
xnor U8924 (N_8924,N_7231,N_7646);
xor U8925 (N_8925,N_7729,N_7993);
nand U8926 (N_8926,N_7664,N_7626);
xor U8927 (N_8927,N_7456,N_7622);
or U8928 (N_8928,N_8171,N_8154);
xnor U8929 (N_8929,N_7886,N_7577);
xor U8930 (N_8930,N_7382,N_8130);
nand U8931 (N_8931,N_7694,N_7241);
and U8932 (N_8932,N_7906,N_8270);
nor U8933 (N_8933,N_8161,N_8079);
nand U8934 (N_8934,N_8335,N_7657);
xor U8935 (N_8935,N_8041,N_7478);
nand U8936 (N_8936,N_8244,N_7310);
nor U8937 (N_8937,N_7718,N_7406);
and U8938 (N_8938,N_8286,N_8372);
and U8939 (N_8939,N_7602,N_7494);
and U8940 (N_8940,N_7438,N_8144);
and U8941 (N_8941,N_7326,N_8151);
or U8942 (N_8942,N_8265,N_8369);
nand U8943 (N_8943,N_8004,N_7688);
nor U8944 (N_8944,N_7853,N_7706);
and U8945 (N_8945,N_8387,N_7515);
and U8946 (N_8946,N_7319,N_7346);
nor U8947 (N_8947,N_8111,N_7653);
and U8948 (N_8948,N_7953,N_7548);
and U8949 (N_8949,N_8338,N_7279);
or U8950 (N_8950,N_7889,N_8009);
or U8951 (N_8951,N_7215,N_8195);
xor U8952 (N_8952,N_8005,N_7814);
or U8953 (N_8953,N_7944,N_7988);
xor U8954 (N_8954,N_7278,N_8044);
nand U8955 (N_8955,N_7846,N_8063);
nand U8956 (N_8956,N_7734,N_7457);
nand U8957 (N_8957,N_7567,N_7825);
xor U8958 (N_8958,N_7703,N_7433);
and U8959 (N_8959,N_7315,N_7957);
or U8960 (N_8960,N_7355,N_8318);
nor U8961 (N_8961,N_7460,N_7742);
nor U8962 (N_8962,N_8098,N_7429);
nor U8963 (N_8963,N_8134,N_8306);
and U8964 (N_8964,N_7835,N_8025);
and U8965 (N_8965,N_7254,N_8141);
nor U8966 (N_8966,N_8158,N_7225);
xnor U8967 (N_8967,N_7504,N_8059);
or U8968 (N_8968,N_7943,N_7681);
and U8969 (N_8969,N_7416,N_8226);
xnor U8970 (N_8970,N_8222,N_8188);
and U8971 (N_8971,N_7507,N_8028);
nor U8972 (N_8972,N_7774,N_8056);
xor U8973 (N_8973,N_7379,N_8243);
xnor U8974 (N_8974,N_8019,N_8125);
or U8975 (N_8975,N_8308,N_7673);
and U8976 (N_8976,N_7342,N_8186);
xor U8977 (N_8977,N_8193,N_8249);
nand U8978 (N_8978,N_7926,N_7652);
xnor U8979 (N_8979,N_8307,N_7875);
and U8980 (N_8980,N_7274,N_8254);
or U8981 (N_8981,N_7683,N_7546);
xor U8982 (N_8982,N_8350,N_8367);
and U8983 (N_8983,N_8319,N_7347);
nand U8984 (N_8984,N_8081,N_8066);
or U8985 (N_8985,N_7290,N_7778);
xor U8986 (N_8986,N_7240,N_7501);
nand U8987 (N_8987,N_7833,N_7732);
nand U8988 (N_8988,N_7978,N_7911);
xnor U8989 (N_8989,N_7611,N_7692);
and U8990 (N_8990,N_7654,N_7712);
nand U8991 (N_8991,N_8399,N_8315);
and U8992 (N_8992,N_7203,N_7288);
or U8993 (N_8993,N_7726,N_7715);
and U8994 (N_8994,N_7601,N_8075);
or U8995 (N_8995,N_7805,N_7389);
xor U8996 (N_8996,N_7446,N_8067);
nor U8997 (N_8997,N_8257,N_8057);
and U8998 (N_8998,N_8197,N_7574);
or U8999 (N_8999,N_7804,N_7560);
and U9000 (N_9000,N_8222,N_7339);
and U9001 (N_9001,N_7502,N_8078);
nor U9002 (N_9002,N_7964,N_7649);
or U9003 (N_9003,N_8323,N_7790);
or U9004 (N_9004,N_7508,N_7550);
nand U9005 (N_9005,N_7748,N_7841);
and U9006 (N_9006,N_8072,N_7747);
nor U9007 (N_9007,N_8200,N_7803);
nand U9008 (N_9008,N_7250,N_8242);
xnor U9009 (N_9009,N_7213,N_8140);
and U9010 (N_9010,N_7611,N_7749);
xnor U9011 (N_9011,N_7922,N_7907);
nand U9012 (N_9012,N_7785,N_7992);
nor U9013 (N_9013,N_7873,N_8358);
nand U9014 (N_9014,N_7800,N_7472);
nor U9015 (N_9015,N_7951,N_7872);
nor U9016 (N_9016,N_7525,N_7221);
nand U9017 (N_9017,N_7706,N_7700);
nand U9018 (N_9018,N_8046,N_7990);
nand U9019 (N_9019,N_8233,N_8018);
and U9020 (N_9020,N_8377,N_7563);
or U9021 (N_9021,N_7847,N_7369);
nor U9022 (N_9022,N_7558,N_7751);
and U9023 (N_9023,N_7913,N_7408);
nand U9024 (N_9024,N_7293,N_7970);
and U9025 (N_9025,N_7653,N_7813);
xnor U9026 (N_9026,N_7230,N_7274);
xor U9027 (N_9027,N_8237,N_8101);
nor U9028 (N_9028,N_8047,N_8168);
xor U9029 (N_9029,N_8130,N_8018);
or U9030 (N_9030,N_7652,N_8148);
nand U9031 (N_9031,N_8387,N_8148);
or U9032 (N_9032,N_8173,N_8375);
and U9033 (N_9033,N_7607,N_8346);
xnor U9034 (N_9034,N_7556,N_7840);
or U9035 (N_9035,N_7653,N_7788);
or U9036 (N_9036,N_7483,N_7806);
or U9037 (N_9037,N_7993,N_7771);
nor U9038 (N_9038,N_8229,N_8194);
or U9039 (N_9039,N_8151,N_7343);
or U9040 (N_9040,N_7637,N_7370);
or U9041 (N_9041,N_7539,N_7969);
and U9042 (N_9042,N_7776,N_8305);
nor U9043 (N_9043,N_7521,N_8283);
and U9044 (N_9044,N_8014,N_8049);
xnor U9045 (N_9045,N_7812,N_7425);
xor U9046 (N_9046,N_8262,N_7529);
nand U9047 (N_9047,N_7850,N_7246);
nor U9048 (N_9048,N_8116,N_7779);
nand U9049 (N_9049,N_8085,N_7343);
or U9050 (N_9050,N_7407,N_7351);
or U9051 (N_9051,N_7513,N_7501);
xnor U9052 (N_9052,N_7591,N_7951);
xor U9053 (N_9053,N_8195,N_7447);
and U9054 (N_9054,N_8147,N_7428);
nand U9055 (N_9055,N_8355,N_7850);
xor U9056 (N_9056,N_7387,N_7739);
and U9057 (N_9057,N_8306,N_8331);
and U9058 (N_9058,N_7231,N_7281);
nor U9059 (N_9059,N_7807,N_7328);
xor U9060 (N_9060,N_7626,N_7940);
nor U9061 (N_9061,N_7668,N_7628);
and U9062 (N_9062,N_7938,N_7972);
nand U9063 (N_9063,N_7273,N_7256);
or U9064 (N_9064,N_7980,N_7468);
or U9065 (N_9065,N_7417,N_8107);
or U9066 (N_9066,N_8378,N_8155);
and U9067 (N_9067,N_8155,N_7278);
nor U9068 (N_9068,N_7674,N_7763);
and U9069 (N_9069,N_7760,N_7922);
xnor U9070 (N_9070,N_8175,N_7223);
nand U9071 (N_9071,N_7682,N_8048);
nor U9072 (N_9072,N_8004,N_7890);
or U9073 (N_9073,N_8230,N_7914);
nand U9074 (N_9074,N_8307,N_7569);
nor U9075 (N_9075,N_8131,N_8028);
xnor U9076 (N_9076,N_7406,N_7937);
nand U9077 (N_9077,N_7918,N_7440);
or U9078 (N_9078,N_7576,N_7538);
xnor U9079 (N_9079,N_7444,N_7374);
and U9080 (N_9080,N_7366,N_7440);
xnor U9081 (N_9081,N_7575,N_7373);
nand U9082 (N_9082,N_7868,N_7450);
or U9083 (N_9083,N_8016,N_8168);
or U9084 (N_9084,N_7514,N_8183);
xor U9085 (N_9085,N_8094,N_8102);
nand U9086 (N_9086,N_8275,N_7762);
or U9087 (N_9087,N_7256,N_7258);
nor U9088 (N_9088,N_7994,N_7584);
xnor U9089 (N_9089,N_8048,N_7461);
nor U9090 (N_9090,N_8006,N_8115);
or U9091 (N_9091,N_7768,N_7751);
nand U9092 (N_9092,N_7262,N_7792);
or U9093 (N_9093,N_8249,N_8154);
nor U9094 (N_9094,N_7635,N_7904);
nor U9095 (N_9095,N_7794,N_7593);
and U9096 (N_9096,N_7669,N_7486);
or U9097 (N_9097,N_8112,N_7853);
xnor U9098 (N_9098,N_7493,N_8149);
xor U9099 (N_9099,N_7430,N_8227);
or U9100 (N_9100,N_8156,N_7316);
or U9101 (N_9101,N_7823,N_8209);
nand U9102 (N_9102,N_8101,N_7522);
xnor U9103 (N_9103,N_7314,N_7444);
xnor U9104 (N_9104,N_8165,N_7659);
nor U9105 (N_9105,N_8334,N_7943);
and U9106 (N_9106,N_7844,N_8325);
xor U9107 (N_9107,N_7708,N_7465);
nor U9108 (N_9108,N_8228,N_8307);
nor U9109 (N_9109,N_7379,N_7281);
nand U9110 (N_9110,N_7701,N_7761);
nand U9111 (N_9111,N_8303,N_8057);
and U9112 (N_9112,N_7828,N_7336);
nand U9113 (N_9113,N_7633,N_7693);
or U9114 (N_9114,N_8104,N_7717);
xnor U9115 (N_9115,N_7218,N_7466);
and U9116 (N_9116,N_7758,N_8363);
nor U9117 (N_9117,N_7488,N_8092);
nor U9118 (N_9118,N_8081,N_7463);
or U9119 (N_9119,N_8373,N_8392);
nand U9120 (N_9120,N_7959,N_7473);
and U9121 (N_9121,N_8033,N_8298);
nand U9122 (N_9122,N_7742,N_7948);
and U9123 (N_9123,N_7980,N_7401);
and U9124 (N_9124,N_7966,N_8085);
xnor U9125 (N_9125,N_7254,N_7501);
or U9126 (N_9126,N_7260,N_7620);
nor U9127 (N_9127,N_7929,N_7652);
or U9128 (N_9128,N_7605,N_7246);
and U9129 (N_9129,N_7485,N_8295);
nor U9130 (N_9130,N_7881,N_7738);
nand U9131 (N_9131,N_8330,N_7251);
nor U9132 (N_9132,N_7494,N_8087);
nor U9133 (N_9133,N_8027,N_7427);
nor U9134 (N_9134,N_7781,N_8096);
or U9135 (N_9135,N_7814,N_7944);
and U9136 (N_9136,N_7671,N_8041);
xnor U9137 (N_9137,N_8315,N_7426);
nor U9138 (N_9138,N_7364,N_7475);
nor U9139 (N_9139,N_7577,N_7822);
xor U9140 (N_9140,N_7354,N_7373);
nor U9141 (N_9141,N_8272,N_7544);
and U9142 (N_9142,N_7751,N_8238);
nor U9143 (N_9143,N_8217,N_7314);
and U9144 (N_9144,N_7822,N_7283);
and U9145 (N_9145,N_8006,N_7858);
nor U9146 (N_9146,N_7922,N_7201);
or U9147 (N_9147,N_8318,N_8125);
or U9148 (N_9148,N_8302,N_7900);
nor U9149 (N_9149,N_8125,N_7855);
xor U9150 (N_9150,N_7333,N_7937);
or U9151 (N_9151,N_7200,N_7674);
nand U9152 (N_9152,N_7532,N_7364);
and U9153 (N_9153,N_8147,N_8092);
and U9154 (N_9154,N_7376,N_8000);
nor U9155 (N_9155,N_7423,N_7875);
or U9156 (N_9156,N_7371,N_8236);
or U9157 (N_9157,N_7498,N_7379);
xnor U9158 (N_9158,N_7596,N_7832);
or U9159 (N_9159,N_7419,N_8094);
nor U9160 (N_9160,N_7670,N_7503);
and U9161 (N_9161,N_8266,N_7734);
nand U9162 (N_9162,N_7355,N_8173);
nand U9163 (N_9163,N_8044,N_7496);
xnor U9164 (N_9164,N_7285,N_8147);
xor U9165 (N_9165,N_8209,N_8234);
and U9166 (N_9166,N_7537,N_7385);
xnor U9167 (N_9167,N_8377,N_8351);
nand U9168 (N_9168,N_7397,N_8359);
xnor U9169 (N_9169,N_7795,N_7209);
nand U9170 (N_9170,N_7338,N_8257);
or U9171 (N_9171,N_7420,N_8195);
xor U9172 (N_9172,N_8232,N_7464);
xor U9173 (N_9173,N_8153,N_8187);
nor U9174 (N_9174,N_7523,N_8285);
nor U9175 (N_9175,N_8091,N_8396);
xor U9176 (N_9176,N_8252,N_8021);
xor U9177 (N_9177,N_8241,N_8096);
xnor U9178 (N_9178,N_7731,N_7373);
or U9179 (N_9179,N_7344,N_7723);
or U9180 (N_9180,N_7518,N_7812);
nand U9181 (N_9181,N_7790,N_7218);
or U9182 (N_9182,N_7862,N_7934);
and U9183 (N_9183,N_7994,N_7909);
nor U9184 (N_9184,N_7418,N_8241);
and U9185 (N_9185,N_8184,N_8254);
and U9186 (N_9186,N_7899,N_8218);
and U9187 (N_9187,N_7834,N_7730);
nand U9188 (N_9188,N_7284,N_8098);
nor U9189 (N_9189,N_8253,N_7773);
nor U9190 (N_9190,N_7431,N_7386);
or U9191 (N_9191,N_7624,N_7954);
xor U9192 (N_9192,N_7335,N_7476);
xor U9193 (N_9193,N_7447,N_7845);
nor U9194 (N_9194,N_7796,N_8000);
or U9195 (N_9195,N_8189,N_8362);
xnor U9196 (N_9196,N_7331,N_7249);
and U9197 (N_9197,N_7561,N_7514);
and U9198 (N_9198,N_7640,N_7486);
or U9199 (N_9199,N_7811,N_7896);
and U9200 (N_9200,N_7267,N_7756);
nor U9201 (N_9201,N_8382,N_7632);
nand U9202 (N_9202,N_7580,N_7298);
nand U9203 (N_9203,N_8107,N_7825);
or U9204 (N_9204,N_8247,N_7483);
or U9205 (N_9205,N_8278,N_8140);
or U9206 (N_9206,N_7763,N_7995);
nor U9207 (N_9207,N_7632,N_7317);
xnor U9208 (N_9208,N_8375,N_7206);
or U9209 (N_9209,N_7661,N_8393);
or U9210 (N_9210,N_7498,N_7327);
or U9211 (N_9211,N_7781,N_7275);
and U9212 (N_9212,N_8162,N_7353);
or U9213 (N_9213,N_7530,N_7808);
or U9214 (N_9214,N_7910,N_8358);
and U9215 (N_9215,N_7438,N_8061);
nor U9216 (N_9216,N_7311,N_7691);
xnor U9217 (N_9217,N_7928,N_7826);
xnor U9218 (N_9218,N_7237,N_7915);
and U9219 (N_9219,N_8331,N_8069);
or U9220 (N_9220,N_8239,N_7513);
or U9221 (N_9221,N_8084,N_7829);
and U9222 (N_9222,N_8246,N_7876);
and U9223 (N_9223,N_7729,N_8193);
and U9224 (N_9224,N_7793,N_8371);
or U9225 (N_9225,N_8392,N_8253);
nor U9226 (N_9226,N_7306,N_7600);
nor U9227 (N_9227,N_7298,N_7654);
nor U9228 (N_9228,N_7862,N_7704);
or U9229 (N_9229,N_7364,N_7379);
nor U9230 (N_9230,N_8193,N_7627);
and U9231 (N_9231,N_7864,N_8284);
xnor U9232 (N_9232,N_8220,N_7610);
and U9233 (N_9233,N_7274,N_8372);
and U9234 (N_9234,N_7269,N_8143);
nand U9235 (N_9235,N_7781,N_7305);
nand U9236 (N_9236,N_7385,N_7342);
xor U9237 (N_9237,N_7368,N_7613);
nor U9238 (N_9238,N_8098,N_7426);
nor U9239 (N_9239,N_7681,N_7865);
nor U9240 (N_9240,N_7716,N_7455);
nand U9241 (N_9241,N_7805,N_7621);
or U9242 (N_9242,N_7311,N_8229);
and U9243 (N_9243,N_7226,N_7796);
or U9244 (N_9244,N_8086,N_7824);
or U9245 (N_9245,N_7403,N_7275);
nand U9246 (N_9246,N_8142,N_7956);
nor U9247 (N_9247,N_7472,N_7689);
and U9248 (N_9248,N_7725,N_7444);
xor U9249 (N_9249,N_8169,N_8296);
nor U9250 (N_9250,N_8161,N_7308);
xor U9251 (N_9251,N_7381,N_7822);
nand U9252 (N_9252,N_7409,N_7786);
nand U9253 (N_9253,N_7504,N_8171);
nor U9254 (N_9254,N_8162,N_7923);
and U9255 (N_9255,N_7329,N_7673);
nor U9256 (N_9256,N_7376,N_7394);
nor U9257 (N_9257,N_8261,N_8378);
xnor U9258 (N_9258,N_7812,N_7474);
nand U9259 (N_9259,N_7865,N_7274);
or U9260 (N_9260,N_7266,N_8140);
or U9261 (N_9261,N_7500,N_7582);
and U9262 (N_9262,N_7284,N_7651);
xor U9263 (N_9263,N_7635,N_7993);
xor U9264 (N_9264,N_7536,N_7813);
nor U9265 (N_9265,N_8385,N_7369);
nand U9266 (N_9266,N_8351,N_7690);
and U9267 (N_9267,N_8323,N_7513);
nand U9268 (N_9268,N_7219,N_7489);
or U9269 (N_9269,N_7553,N_8070);
xnor U9270 (N_9270,N_7687,N_7468);
xnor U9271 (N_9271,N_7381,N_8286);
and U9272 (N_9272,N_7504,N_7871);
or U9273 (N_9273,N_7550,N_7580);
nor U9274 (N_9274,N_7479,N_7657);
nor U9275 (N_9275,N_8241,N_7221);
and U9276 (N_9276,N_7360,N_8027);
or U9277 (N_9277,N_8065,N_7631);
or U9278 (N_9278,N_7521,N_7532);
nand U9279 (N_9279,N_8170,N_8281);
nor U9280 (N_9280,N_7649,N_7228);
nor U9281 (N_9281,N_7901,N_7203);
xor U9282 (N_9282,N_7803,N_8314);
xnor U9283 (N_9283,N_7968,N_8164);
and U9284 (N_9284,N_7648,N_8237);
and U9285 (N_9285,N_7425,N_8024);
and U9286 (N_9286,N_7347,N_8246);
nor U9287 (N_9287,N_7551,N_7710);
and U9288 (N_9288,N_7979,N_7243);
xor U9289 (N_9289,N_8129,N_7785);
nand U9290 (N_9290,N_7470,N_8099);
xnor U9291 (N_9291,N_8220,N_8081);
xor U9292 (N_9292,N_8059,N_7443);
xor U9293 (N_9293,N_7477,N_7205);
nor U9294 (N_9294,N_7333,N_7928);
and U9295 (N_9295,N_7721,N_7714);
nand U9296 (N_9296,N_7592,N_8091);
xnor U9297 (N_9297,N_8056,N_7793);
nor U9298 (N_9298,N_7304,N_7657);
nand U9299 (N_9299,N_7387,N_7283);
or U9300 (N_9300,N_7980,N_7951);
nor U9301 (N_9301,N_7238,N_7309);
nor U9302 (N_9302,N_8168,N_7623);
and U9303 (N_9303,N_7238,N_8272);
or U9304 (N_9304,N_8232,N_8382);
nor U9305 (N_9305,N_8013,N_7433);
nand U9306 (N_9306,N_7406,N_8167);
nand U9307 (N_9307,N_7797,N_7289);
and U9308 (N_9308,N_8388,N_8379);
nand U9309 (N_9309,N_7275,N_7712);
or U9310 (N_9310,N_7814,N_7405);
and U9311 (N_9311,N_8050,N_7800);
nand U9312 (N_9312,N_8238,N_7440);
and U9313 (N_9313,N_7883,N_8213);
xor U9314 (N_9314,N_7413,N_7689);
nor U9315 (N_9315,N_7399,N_7716);
nor U9316 (N_9316,N_7572,N_7639);
or U9317 (N_9317,N_7266,N_7570);
nand U9318 (N_9318,N_7760,N_7299);
nand U9319 (N_9319,N_7996,N_7261);
xnor U9320 (N_9320,N_7569,N_7310);
nand U9321 (N_9321,N_7887,N_7781);
nand U9322 (N_9322,N_8387,N_7510);
nor U9323 (N_9323,N_7612,N_7663);
and U9324 (N_9324,N_8271,N_8161);
xnor U9325 (N_9325,N_7272,N_7207);
xor U9326 (N_9326,N_7564,N_7956);
xor U9327 (N_9327,N_7548,N_7801);
xor U9328 (N_9328,N_7789,N_7301);
nor U9329 (N_9329,N_8313,N_8226);
or U9330 (N_9330,N_7266,N_7944);
and U9331 (N_9331,N_7662,N_8264);
and U9332 (N_9332,N_7949,N_8009);
nor U9333 (N_9333,N_8352,N_8223);
nor U9334 (N_9334,N_8142,N_8023);
and U9335 (N_9335,N_8301,N_8336);
nand U9336 (N_9336,N_7630,N_7972);
nand U9337 (N_9337,N_7674,N_8046);
nor U9338 (N_9338,N_7340,N_7805);
or U9339 (N_9339,N_7286,N_7585);
nor U9340 (N_9340,N_7530,N_7235);
nor U9341 (N_9341,N_7310,N_7972);
nand U9342 (N_9342,N_7882,N_7913);
nor U9343 (N_9343,N_7343,N_7962);
xnor U9344 (N_9344,N_7306,N_8228);
nor U9345 (N_9345,N_7550,N_7326);
or U9346 (N_9346,N_7561,N_8083);
xnor U9347 (N_9347,N_7843,N_7330);
xor U9348 (N_9348,N_7381,N_7980);
nand U9349 (N_9349,N_7699,N_7908);
nor U9350 (N_9350,N_7217,N_7248);
nor U9351 (N_9351,N_7862,N_7463);
and U9352 (N_9352,N_7907,N_7792);
xnor U9353 (N_9353,N_7476,N_8042);
nand U9354 (N_9354,N_7496,N_8178);
or U9355 (N_9355,N_8306,N_8207);
nand U9356 (N_9356,N_7740,N_7316);
xor U9357 (N_9357,N_7622,N_7417);
or U9358 (N_9358,N_7845,N_7903);
nor U9359 (N_9359,N_8320,N_7720);
nor U9360 (N_9360,N_8253,N_8361);
nand U9361 (N_9361,N_7611,N_7348);
or U9362 (N_9362,N_7585,N_8167);
nor U9363 (N_9363,N_7304,N_8075);
and U9364 (N_9364,N_7210,N_7716);
nor U9365 (N_9365,N_8104,N_7662);
nor U9366 (N_9366,N_7275,N_8029);
nand U9367 (N_9367,N_7444,N_7778);
and U9368 (N_9368,N_7533,N_8379);
and U9369 (N_9369,N_7673,N_8298);
and U9370 (N_9370,N_7792,N_8122);
xor U9371 (N_9371,N_7916,N_7502);
nand U9372 (N_9372,N_8121,N_8056);
or U9373 (N_9373,N_8044,N_7464);
or U9374 (N_9374,N_7628,N_8240);
and U9375 (N_9375,N_8337,N_7758);
nor U9376 (N_9376,N_7278,N_7507);
nand U9377 (N_9377,N_8366,N_8117);
xnor U9378 (N_9378,N_8092,N_7979);
and U9379 (N_9379,N_7745,N_8257);
or U9380 (N_9380,N_7643,N_8292);
nor U9381 (N_9381,N_7831,N_7823);
xor U9382 (N_9382,N_8174,N_7431);
and U9383 (N_9383,N_8064,N_7952);
nand U9384 (N_9384,N_8107,N_7808);
nand U9385 (N_9385,N_7604,N_7822);
and U9386 (N_9386,N_7551,N_8026);
nand U9387 (N_9387,N_7257,N_8207);
xnor U9388 (N_9388,N_7914,N_8286);
and U9389 (N_9389,N_8303,N_7459);
and U9390 (N_9390,N_8042,N_7353);
or U9391 (N_9391,N_8155,N_7263);
and U9392 (N_9392,N_8394,N_7206);
xnor U9393 (N_9393,N_7915,N_8110);
nor U9394 (N_9394,N_8009,N_7342);
and U9395 (N_9395,N_7419,N_7364);
nand U9396 (N_9396,N_7983,N_7912);
nand U9397 (N_9397,N_8250,N_7741);
or U9398 (N_9398,N_7797,N_7445);
and U9399 (N_9399,N_7459,N_7496);
xor U9400 (N_9400,N_7500,N_8070);
xnor U9401 (N_9401,N_8259,N_8081);
nor U9402 (N_9402,N_7575,N_8300);
and U9403 (N_9403,N_7526,N_7820);
nor U9404 (N_9404,N_8215,N_7712);
nor U9405 (N_9405,N_7503,N_8025);
or U9406 (N_9406,N_8173,N_7870);
or U9407 (N_9407,N_8051,N_8397);
nand U9408 (N_9408,N_8078,N_7824);
xnor U9409 (N_9409,N_7627,N_7275);
xor U9410 (N_9410,N_7852,N_7609);
and U9411 (N_9411,N_7203,N_7271);
and U9412 (N_9412,N_8173,N_8216);
nor U9413 (N_9413,N_7369,N_7508);
nor U9414 (N_9414,N_7743,N_7986);
xnor U9415 (N_9415,N_8086,N_7741);
or U9416 (N_9416,N_8046,N_8374);
xor U9417 (N_9417,N_7571,N_7855);
nor U9418 (N_9418,N_7522,N_7922);
nand U9419 (N_9419,N_8095,N_7742);
or U9420 (N_9420,N_8129,N_7933);
and U9421 (N_9421,N_7731,N_8282);
nor U9422 (N_9422,N_7336,N_8001);
nand U9423 (N_9423,N_7439,N_7242);
and U9424 (N_9424,N_8061,N_7436);
xor U9425 (N_9425,N_7461,N_7592);
nand U9426 (N_9426,N_7590,N_8050);
nor U9427 (N_9427,N_7354,N_7754);
xnor U9428 (N_9428,N_8270,N_8083);
and U9429 (N_9429,N_7383,N_7546);
xor U9430 (N_9430,N_7773,N_7496);
nor U9431 (N_9431,N_7444,N_7247);
xnor U9432 (N_9432,N_7670,N_8391);
xor U9433 (N_9433,N_8109,N_7687);
nor U9434 (N_9434,N_7547,N_8175);
nor U9435 (N_9435,N_7519,N_7743);
or U9436 (N_9436,N_8221,N_7901);
xor U9437 (N_9437,N_8385,N_8070);
and U9438 (N_9438,N_7507,N_8158);
xor U9439 (N_9439,N_7626,N_7482);
or U9440 (N_9440,N_8322,N_7544);
xor U9441 (N_9441,N_7921,N_7294);
xor U9442 (N_9442,N_7351,N_8183);
and U9443 (N_9443,N_8132,N_7983);
nand U9444 (N_9444,N_8068,N_8303);
nand U9445 (N_9445,N_7906,N_7555);
xnor U9446 (N_9446,N_7817,N_7549);
xnor U9447 (N_9447,N_7843,N_8022);
nor U9448 (N_9448,N_8229,N_8370);
or U9449 (N_9449,N_7255,N_7865);
and U9450 (N_9450,N_8348,N_8374);
nor U9451 (N_9451,N_7766,N_8236);
nor U9452 (N_9452,N_7887,N_7588);
nand U9453 (N_9453,N_8377,N_7527);
nor U9454 (N_9454,N_8176,N_7860);
nand U9455 (N_9455,N_7978,N_8180);
and U9456 (N_9456,N_8108,N_7520);
nand U9457 (N_9457,N_7971,N_7322);
xor U9458 (N_9458,N_7445,N_7633);
nand U9459 (N_9459,N_8180,N_8280);
nand U9460 (N_9460,N_7918,N_8072);
or U9461 (N_9461,N_7407,N_7563);
xor U9462 (N_9462,N_7662,N_7710);
and U9463 (N_9463,N_7651,N_7908);
and U9464 (N_9464,N_8116,N_7573);
xnor U9465 (N_9465,N_7604,N_7306);
nor U9466 (N_9466,N_7682,N_7932);
nor U9467 (N_9467,N_7644,N_8254);
xnor U9468 (N_9468,N_7280,N_8308);
xor U9469 (N_9469,N_7817,N_7356);
nor U9470 (N_9470,N_8058,N_8117);
nand U9471 (N_9471,N_8380,N_8067);
nand U9472 (N_9472,N_7594,N_8304);
nor U9473 (N_9473,N_7257,N_7525);
nor U9474 (N_9474,N_8243,N_7737);
xor U9475 (N_9475,N_8004,N_7500);
nor U9476 (N_9476,N_8276,N_7329);
and U9477 (N_9477,N_7413,N_7648);
nor U9478 (N_9478,N_7212,N_7305);
or U9479 (N_9479,N_7805,N_8010);
and U9480 (N_9480,N_7896,N_8097);
or U9481 (N_9481,N_7662,N_8075);
xor U9482 (N_9482,N_7441,N_8144);
nor U9483 (N_9483,N_7429,N_7685);
and U9484 (N_9484,N_8385,N_7944);
xor U9485 (N_9485,N_8071,N_8362);
or U9486 (N_9486,N_7946,N_8089);
and U9487 (N_9487,N_7651,N_8089);
xnor U9488 (N_9488,N_7568,N_7812);
or U9489 (N_9489,N_7899,N_8134);
nor U9490 (N_9490,N_8136,N_7263);
and U9491 (N_9491,N_8304,N_7535);
or U9492 (N_9492,N_7746,N_7356);
and U9493 (N_9493,N_8219,N_7628);
or U9494 (N_9494,N_7465,N_8027);
and U9495 (N_9495,N_7496,N_7284);
nand U9496 (N_9496,N_7859,N_7246);
xor U9497 (N_9497,N_7750,N_8119);
or U9498 (N_9498,N_7665,N_8323);
or U9499 (N_9499,N_7536,N_7826);
nor U9500 (N_9500,N_7944,N_8380);
nand U9501 (N_9501,N_8201,N_7833);
or U9502 (N_9502,N_7985,N_8173);
and U9503 (N_9503,N_7936,N_7488);
xnor U9504 (N_9504,N_7436,N_7374);
or U9505 (N_9505,N_7417,N_7293);
nor U9506 (N_9506,N_7794,N_7729);
nand U9507 (N_9507,N_7937,N_7437);
and U9508 (N_9508,N_8024,N_7275);
nand U9509 (N_9509,N_7535,N_8102);
and U9510 (N_9510,N_7209,N_7232);
xor U9511 (N_9511,N_8219,N_8266);
nor U9512 (N_9512,N_7397,N_8283);
or U9513 (N_9513,N_7843,N_8162);
xnor U9514 (N_9514,N_7974,N_7899);
or U9515 (N_9515,N_7807,N_7727);
nor U9516 (N_9516,N_7762,N_7908);
xnor U9517 (N_9517,N_7665,N_7240);
and U9518 (N_9518,N_7201,N_7851);
xor U9519 (N_9519,N_8024,N_8157);
nor U9520 (N_9520,N_7565,N_7461);
or U9521 (N_9521,N_8031,N_7624);
and U9522 (N_9522,N_7882,N_8276);
and U9523 (N_9523,N_7764,N_7292);
xnor U9524 (N_9524,N_7933,N_8175);
nor U9525 (N_9525,N_7465,N_7821);
xor U9526 (N_9526,N_7935,N_8117);
xor U9527 (N_9527,N_7893,N_7617);
nand U9528 (N_9528,N_7235,N_8039);
nand U9529 (N_9529,N_7911,N_8141);
nand U9530 (N_9530,N_7699,N_7331);
nand U9531 (N_9531,N_8349,N_8061);
nor U9532 (N_9532,N_7632,N_7245);
or U9533 (N_9533,N_7402,N_7738);
nand U9534 (N_9534,N_7411,N_7894);
nor U9535 (N_9535,N_8213,N_8131);
nor U9536 (N_9536,N_7957,N_7509);
nand U9537 (N_9537,N_7915,N_7577);
nor U9538 (N_9538,N_8301,N_8143);
or U9539 (N_9539,N_8244,N_8117);
nand U9540 (N_9540,N_7653,N_7201);
and U9541 (N_9541,N_7377,N_7267);
and U9542 (N_9542,N_7753,N_8190);
nor U9543 (N_9543,N_8290,N_7893);
xor U9544 (N_9544,N_8258,N_7274);
nor U9545 (N_9545,N_7946,N_8244);
and U9546 (N_9546,N_7312,N_7372);
or U9547 (N_9547,N_8356,N_7718);
xor U9548 (N_9548,N_7467,N_7446);
nand U9549 (N_9549,N_7425,N_7281);
nor U9550 (N_9550,N_8242,N_8292);
nor U9551 (N_9551,N_7754,N_7383);
xor U9552 (N_9552,N_7893,N_8260);
and U9553 (N_9553,N_7676,N_7554);
nor U9554 (N_9554,N_7955,N_8234);
xor U9555 (N_9555,N_7717,N_7972);
or U9556 (N_9556,N_7388,N_7282);
nor U9557 (N_9557,N_8172,N_8320);
and U9558 (N_9558,N_7736,N_7838);
nand U9559 (N_9559,N_7987,N_7212);
or U9560 (N_9560,N_8127,N_7619);
nor U9561 (N_9561,N_7717,N_7701);
xnor U9562 (N_9562,N_7420,N_8082);
nor U9563 (N_9563,N_7855,N_8128);
or U9564 (N_9564,N_7812,N_7219);
and U9565 (N_9565,N_7482,N_7754);
nand U9566 (N_9566,N_8031,N_8138);
nor U9567 (N_9567,N_7609,N_7765);
or U9568 (N_9568,N_8076,N_8135);
nand U9569 (N_9569,N_8322,N_7465);
nor U9570 (N_9570,N_7607,N_7318);
and U9571 (N_9571,N_8199,N_8103);
xnor U9572 (N_9572,N_7324,N_7624);
nor U9573 (N_9573,N_7478,N_7835);
and U9574 (N_9574,N_8364,N_7527);
xor U9575 (N_9575,N_7585,N_7430);
xnor U9576 (N_9576,N_7499,N_7283);
and U9577 (N_9577,N_8104,N_7567);
or U9578 (N_9578,N_8064,N_7236);
nand U9579 (N_9579,N_8157,N_8075);
nand U9580 (N_9580,N_7593,N_7737);
nand U9581 (N_9581,N_7310,N_7840);
xor U9582 (N_9582,N_7648,N_7252);
and U9583 (N_9583,N_7285,N_7734);
and U9584 (N_9584,N_7536,N_7930);
xnor U9585 (N_9585,N_7852,N_7806);
xor U9586 (N_9586,N_7527,N_8192);
nand U9587 (N_9587,N_7247,N_7467);
or U9588 (N_9588,N_7984,N_7614);
and U9589 (N_9589,N_7947,N_8159);
or U9590 (N_9590,N_7955,N_7740);
or U9591 (N_9591,N_7638,N_8021);
or U9592 (N_9592,N_7444,N_7359);
or U9593 (N_9593,N_8004,N_8352);
nand U9594 (N_9594,N_7691,N_8267);
nand U9595 (N_9595,N_7742,N_7772);
xor U9596 (N_9596,N_7519,N_7233);
xor U9597 (N_9597,N_7857,N_8012);
xor U9598 (N_9598,N_7595,N_7211);
xnor U9599 (N_9599,N_7336,N_7410);
nand U9600 (N_9600,N_9103,N_9272);
nor U9601 (N_9601,N_8698,N_9134);
nand U9602 (N_9602,N_8679,N_9087);
nand U9603 (N_9603,N_8933,N_9198);
nand U9604 (N_9604,N_8978,N_8980);
nand U9605 (N_9605,N_8677,N_8651);
xor U9606 (N_9606,N_9305,N_9458);
nor U9607 (N_9607,N_9223,N_9069);
nor U9608 (N_9608,N_9238,N_8521);
nor U9609 (N_9609,N_8496,N_9130);
or U9610 (N_9610,N_8750,N_8645);
xnor U9611 (N_9611,N_8783,N_9581);
nand U9612 (N_9612,N_9232,N_8441);
nand U9613 (N_9613,N_9514,N_8658);
nand U9614 (N_9614,N_8424,N_8764);
or U9615 (N_9615,N_9189,N_9523);
and U9616 (N_9616,N_8778,N_9241);
and U9617 (N_9617,N_8553,N_8605);
nand U9618 (N_9618,N_8542,N_9403);
xor U9619 (N_9619,N_8788,N_9288);
and U9620 (N_9620,N_9294,N_9506);
or U9621 (N_9621,N_8505,N_8501);
or U9622 (N_9622,N_8884,N_9244);
nand U9623 (N_9623,N_9287,N_9290);
and U9624 (N_9624,N_9267,N_8408);
nand U9625 (N_9625,N_8723,N_8608);
xnor U9626 (N_9626,N_8599,N_8756);
nand U9627 (N_9627,N_8641,N_9599);
nor U9628 (N_9628,N_9121,N_9030);
or U9629 (N_9629,N_8481,N_8484);
or U9630 (N_9630,N_9058,N_9182);
nand U9631 (N_9631,N_9407,N_8759);
or U9632 (N_9632,N_9497,N_8771);
or U9633 (N_9633,N_9117,N_9071);
and U9634 (N_9634,N_8707,N_8949);
xor U9635 (N_9635,N_9574,N_9509);
and U9636 (N_9636,N_9227,N_9564);
xnor U9637 (N_9637,N_9469,N_8656);
xor U9638 (N_9638,N_9374,N_8425);
or U9639 (N_9639,N_9319,N_9229);
nor U9640 (N_9640,N_9107,N_8740);
nand U9641 (N_9641,N_8718,N_9116);
nand U9642 (N_9642,N_9304,N_9396);
and U9643 (N_9643,N_8811,N_8515);
and U9644 (N_9644,N_8513,N_8416);
nand U9645 (N_9645,N_9181,N_9500);
nor U9646 (N_9646,N_8734,N_9222);
nand U9647 (N_9647,N_9484,N_9490);
nand U9648 (N_9648,N_8816,N_9263);
nand U9649 (N_9649,N_9275,N_8598);
nand U9650 (N_9650,N_8455,N_9170);
nor U9651 (N_9651,N_9369,N_8660);
xnor U9652 (N_9652,N_8839,N_9334);
or U9653 (N_9653,N_9335,N_8937);
nor U9654 (N_9654,N_9445,N_9416);
or U9655 (N_9655,N_9342,N_8670);
xor U9656 (N_9656,N_9173,N_8886);
or U9657 (N_9657,N_8671,N_8668);
xnor U9658 (N_9658,N_9470,N_8572);
xor U9659 (N_9659,N_9346,N_9593);
nand U9660 (N_9660,N_9251,N_8556);
xnor U9661 (N_9661,N_9004,N_8986);
nand U9662 (N_9662,N_8433,N_8749);
nor U9663 (N_9663,N_8796,N_9177);
xnor U9664 (N_9664,N_8953,N_8638);
and U9665 (N_9665,N_9091,N_8554);
or U9666 (N_9666,N_9577,N_9115);
and U9667 (N_9667,N_8987,N_9329);
or U9668 (N_9668,N_9217,N_8571);
xnor U9669 (N_9669,N_8958,N_8557);
nor U9670 (N_9670,N_8813,N_8731);
or U9671 (N_9671,N_9277,N_9088);
nand U9672 (N_9672,N_9482,N_9373);
or U9673 (N_9673,N_9359,N_8857);
xnor U9674 (N_9674,N_8536,N_9518);
xor U9675 (N_9675,N_8842,N_9151);
nand U9676 (N_9676,N_9153,N_8498);
nor U9677 (N_9677,N_8402,N_9412);
xnor U9678 (N_9678,N_8517,N_9547);
nand U9679 (N_9679,N_8966,N_9344);
xor U9680 (N_9680,N_8997,N_8954);
nand U9681 (N_9681,N_9281,N_8792);
nor U9682 (N_9682,N_8843,N_8591);
or U9683 (N_9683,N_9269,N_9452);
nor U9684 (N_9684,N_8854,N_8473);
nor U9685 (N_9685,N_8904,N_9154);
or U9686 (N_9686,N_8637,N_9245);
and U9687 (N_9687,N_9527,N_8985);
nand U9688 (N_9688,N_9094,N_9074);
or U9689 (N_9689,N_8465,N_8873);
nor U9690 (N_9690,N_8782,N_9358);
and U9691 (N_9691,N_8472,N_8655);
or U9692 (N_9692,N_8931,N_8744);
nor U9693 (N_9693,N_9535,N_8624);
and U9694 (N_9694,N_8798,N_8566);
nor U9695 (N_9695,N_8838,N_9164);
and U9696 (N_9696,N_8634,N_8576);
and U9697 (N_9697,N_8715,N_8578);
nor U9698 (N_9698,N_9466,N_8661);
nor U9699 (N_9699,N_9278,N_9323);
nor U9700 (N_9700,N_9018,N_8494);
xnor U9701 (N_9701,N_9163,N_8528);
xnor U9702 (N_9702,N_9208,N_8550);
and U9703 (N_9703,N_9234,N_9333);
and U9704 (N_9704,N_9023,N_8866);
xnor U9705 (N_9705,N_8642,N_9253);
xor U9706 (N_9706,N_9427,N_9159);
or U9707 (N_9707,N_8999,N_8810);
or U9708 (N_9708,N_9356,N_8647);
and U9709 (N_9709,N_8486,N_9447);
nor U9710 (N_9710,N_9510,N_9276);
or U9711 (N_9711,N_9194,N_9420);
xnor U9712 (N_9712,N_9364,N_9226);
xnor U9713 (N_9713,N_8502,N_8631);
and U9714 (N_9714,N_9021,N_9465);
or U9715 (N_9715,N_9519,N_8864);
nor U9716 (N_9716,N_8547,N_8560);
or U9717 (N_9717,N_8574,N_9051);
nor U9718 (N_9718,N_9578,N_9195);
xnor U9719 (N_9719,N_8663,N_8940);
and U9720 (N_9720,N_9009,N_9001);
and U9721 (N_9721,N_8907,N_8575);
or U9722 (N_9722,N_9439,N_9136);
xor U9723 (N_9723,N_8922,N_9044);
nor U9724 (N_9724,N_9302,N_8834);
xor U9725 (N_9725,N_9491,N_9247);
nand U9726 (N_9726,N_9137,N_9256);
or U9727 (N_9727,N_8561,N_9179);
and U9728 (N_9728,N_8601,N_9594);
or U9729 (N_9729,N_9060,N_8785);
and U9730 (N_9730,N_9201,N_8879);
nand U9731 (N_9731,N_9083,N_9525);
nor U9732 (N_9732,N_8629,N_9589);
and U9733 (N_9733,N_9128,N_8511);
nand U9734 (N_9734,N_8950,N_8616);
xnor U9735 (N_9735,N_8431,N_8628);
nand U9736 (N_9736,N_8973,N_9119);
nand U9737 (N_9737,N_8483,N_8898);
and U9738 (N_9738,N_8943,N_8824);
xor U9739 (N_9739,N_9556,N_8935);
nor U9740 (N_9740,N_9230,N_9488);
or U9741 (N_9741,N_8452,N_9014);
nor U9742 (N_9742,N_9575,N_8835);
nand U9743 (N_9743,N_8475,N_8860);
or U9744 (N_9744,N_8509,N_9279);
and U9745 (N_9745,N_8758,N_8530);
and U9746 (N_9746,N_8972,N_8582);
nand U9747 (N_9747,N_9220,N_9029);
xor U9748 (N_9748,N_8529,N_9434);
nand U9749 (N_9749,N_9224,N_9101);
nand U9750 (N_9750,N_9282,N_9537);
nor U9751 (N_9751,N_9406,N_8769);
nand U9752 (N_9752,N_9444,N_9080);
or U9753 (N_9753,N_8714,N_9148);
nor U9754 (N_9754,N_9122,N_9025);
and U9755 (N_9755,N_9089,N_9096);
nand U9756 (N_9756,N_9493,N_8467);
or U9757 (N_9757,N_9554,N_8685);
nand U9758 (N_9758,N_9235,N_8666);
or U9759 (N_9759,N_9197,N_9546);
and U9760 (N_9760,N_8748,N_8533);
xor U9761 (N_9761,N_9111,N_8401);
nor U9762 (N_9762,N_9214,N_8704);
or U9763 (N_9763,N_8590,N_9125);
and U9764 (N_9764,N_8752,N_9487);
nor U9765 (N_9765,N_9039,N_8956);
nor U9766 (N_9766,N_8721,N_8900);
and U9767 (N_9767,N_9534,N_9242);
xor U9768 (N_9768,N_9363,N_9285);
xnor U9769 (N_9769,N_8817,N_8700);
or U9770 (N_9770,N_9280,N_9558);
nand U9771 (N_9771,N_9395,N_9399);
nand U9772 (N_9772,N_8490,N_9417);
xnor U9773 (N_9773,N_8623,N_8439);
nand U9774 (N_9774,N_9461,N_9050);
nor U9775 (N_9775,N_8770,N_9563);
nor U9776 (N_9776,N_9414,N_9544);
or U9777 (N_9777,N_9078,N_9565);
nor U9778 (N_9778,N_8797,N_8510);
or U9779 (N_9779,N_9320,N_9200);
nor U9780 (N_9780,N_8754,N_9202);
nand U9781 (N_9781,N_8829,N_8535);
or U9782 (N_9782,N_8418,N_9316);
nor U9783 (N_9783,N_9053,N_8837);
nor U9784 (N_9784,N_9375,N_9236);
and U9785 (N_9785,N_9105,N_8709);
or U9786 (N_9786,N_9569,N_9477);
and U9787 (N_9787,N_9585,N_8621);
nand U9788 (N_9788,N_8789,N_9587);
and U9789 (N_9789,N_9436,N_9433);
or U9790 (N_9790,N_8625,N_8890);
nand U9791 (N_9791,N_9503,N_8902);
xnor U9792 (N_9792,N_9120,N_9257);
nor U9793 (N_9793,N_9038,N_8516);
nand U9794 (N_9794,N_9057,N_8541);
or U9795 (N_9795,N_8603,N_8991);
and U9796 (N_9796,N_9144,N_8870);
nor U9797 (N_9797,N_8551,N_9501);
nand U9798 (N_9798,N_8844,N_9492);
or U9799 (N_9799,N_9258,N_9261);
nand U9800 (N_9800,N_8780,N_8805);
or U9801 (N_9801,N_8451,N_8876);
nand U9802 (N_9802,N_9552,N_9028);
or U9803 (N_9803,N_8703,N_9070);
xor U9804 (N_9804,N_8604,N_8945);
or U9805 (N_9805,N_8680,N_8400);
nand U9806 (N_9806,N_9349,N_8614);
nand U9807 (N_9807,N_9210,N_9521);
and U9808 (N_9808,N_8585,N_9560);
nor U9809 (N_9809,N_9306,N_8919);
or U9810 (N_9810,N_8894,N_9193);
nor U9811 (N_9811,N_8539,N_9212);
xor U9812 (N_9812,N_8428,N_9409);
nor U9813 (N_9813,N_9106,N_8653);
nand U9814 (N_9814,N_8440,N_8538);
and U9815 (N_9815,N_9048,N_9225);
and U9816 (N_9816,N_8442,N_9536);
and U9817 (N_9817,N_8468,N_9517);
and U9818 (N_9818,N_9024,N_9446);
or U9819 (N_9819,N_8983,N_8918);
nor U9820 (N_9820,N_8957,N_8588);
and U9821 (N_9821,N_9026,N_8643);
xnor U9822 (N_9822,N_9475,N_9459);
xor U9823 (N_9823,N_9215,N_8449);
and U9824 (N_9824,N_8544,N_8790);
nand U9825 (N_9825,N_9429,N_9331);
nand U9826 (N_9826,N_9318,N_9486);
nand U9827 (N_9827,N_8863,N_8742);
or U9828 (N_9828,N_8753,N_9324);
xor U9829 (N_9829,N_8522,N_8411);
nor U9830 (N_9830,N_8994,N_9478);
or U9831 (N_9831,N_8868,N_9408);
or U9832 (N_9832,N_8644,N_8888);
and U9833 (N_9833,N_8885,N_8491);
xnor U9834 (N_9834,N_8507,N_8567);
and U9835 (N_9835,N_9424,N_8760);
or U9836 (N_9836,N_8777,N_8447);
and U9837 (N_9837,N_9161,N_8775);
nand U9838 (N_9838,N_8579,N_9312);
xor U9839 (N_9839,N_9379,N_8892);
nand U9840 (N_9840,N_8595,N_8427);
xnor U9841 (N_9841,N_9557,N_8836);
xnor U9842 (N_9842,N_9207,N_9315);
nor U9843 (N_9843,N_9428,N_8664);
nor U9844 (N_9844,N_9528,N_9572);
nand U9845 (N_9845,N_9160,N_8801);
nand U9846 (N_9846,N_8974,N_9489);
nor U9847 (N_9847,N_9192,N_9171);
nand U9848 (N_9848,N_8955,N_9108);
or U9849 (N_9849,N_9314,N_9553);
nand U9850 (N_9850,N_9027,N_8909);
nor U9851 (N_9851,N_9249,N_9328);
or U9852 (N_9852,N_9046,N_8755);
xor U9853 (N_9853,N_8794,N_9545);
and U9854 (N_9854,N_8594,N_8746);
xnor U9855 (N_9855,N_9064,N_8524);
nand U9856 (N_9856,N_8687,N_8696);
or U9857 (N_9857,N_9457,N_9114);
and U9858 (N_9858,N_8606,N_9000);
nand U9859 (N_9859,N_9481,N_9451);
nand U9860 (N_9860,N_9296,N_9218);
xnor U9861 (N_9861,N_8968,N_8423);
xnor U9862 (N_9862,N_8725,N_9152);
and U9863 (N_9863,N_8480,N_9430);
or U9864 (N_9864,N_8701,N_9240);
nor U9865 (N_9865,N_9450,N_8877);
nand U9866 (N_9866,N_8406,N_9596);
nor U9867 (N_9867,N_8692,N_9321);
or U9868 (N_9868,N_8984,N_8667);
nand U9869 (N_9869,N_8512,N_9365);
or U9870 (N_9870,N_8657,N_9259);
nand U9871 (N_9871,N_8462,N_8706);
or U9872 (N_9872,N_8458,N_8932);
and U9873 (N_9873,N_8543,N_8745);
xnor U9874 (N_9874,N_8826,N_9549);
and U9875 (N_9875,N_9378,N_8518);
and U9876 (N_9876,N_8855,N_8683);
nand U9877 (N_9877,N_8640,N_9570);
or U9878 (N_9878,N_9271,N_9162);
nor U9879 (N_9879,N_8727,N_9471);
or U9880 (N_9880,N_8961,N_9502);
nand U9881 (N_9881,N_9006,N_8503);
nor U9882 (N_9882,N_8799,N_8930);
and U9883 (N_9883,N_9539,N_9135);
nand U9884 (N_9884,N_9262,N_8414);
nand U9885 (N_9885,N_8445,N_9190);
and U9886 (N_9886,N_9090,N_9100);
nor U9887 (N_9887,N_8874,N_8766);
and U9888 (N_9888,N_8823,N_8948);
and U9889 (N_9889,N_9499,N_8726);
xnor U9890 (N_9890,N_8534,N_9307);
xnor U9891 (N_9891,N_9464,N_9515);
xor U9892 (N_9892,N_8872,N_8691);
and U9893 (N_9893,N_9268,N_9016);
xnor U9894 (N_9894,N_8791,N_9308);
xor U9895 (N_9895,N_9309,N_9140);
and U9896 (N_9896,N_8548,N_9423);
xor U9897 (N_9897,N_8896,N_9448);
nand U9898 (N_9898,N_9310,N_9005);
or U9899 (N_9899,N_8850,N_8409);
nor U9900 (N_9900,N_8587,N_8415);
and U9901 (N_9901,N_8830,N_9054);
nor U9902 (N_9902,N_9150,N_8906);
and U9903 (N_9903,N_8403,N_8912);
xnor U9904 (N_9904,N_9205,N_9426);
xor U9905 (N_9905,N_9524,N_9180);
or U9906 (N_9906,N_9239,N_9084);
xor U9907 (N_9907,N_8537,N_8812);
nand U9908 (N_9908,N_8728,N_9332);
and U9909 (N_9909,N_9463,N_8674);
xnor U9910 (N_9910,N_9040,N_8962);
and U9911 (N_9911,N_8531,N_9008);
nor U9912 (N_9912,N_8800,N_9299);
nand U9913 (N_9913,N_9512,N_8546);
or U9914 (N_9914,N_9597,N_9325);
nor U9915 (N_9915,N_8916,N_8652);
or U9916 (N_9916,N_8584,N_8761);
xor U9917 (N_9917,N_9185,N_9383);
or U9918 (N_9918,N_9052,N_8928);
and U9919 (N_9919,N_8913,N_8713);
and U9920 (N_9920,N_9017,N_8814);
and U9921 (N_9921,N_9274,N_8432);
xnor U9922 (N_9922,N_9149,N_9246);
nand U9923 (N_9923,N_9522,N_8716);
nand U9924 (N_9924,N_9166,N_9206);
nand U9925 (N_9925,N_8632,N_9067);
xnor U9926 (N_9926,N_9400,N_9387);
and U9927 (N_9927,N_8577,N_9370);
nor U9928 (N_9928,N_9485,N_8508);
nand U9929 (N_9929,N_8471,N_8938);
nand U9930 (N_9930,N_9548,N_8695);
nand U9931 (N_9931,N_8689,N_9479);
or U9932 (N_9932,N_9203,N_9394);
xor U9933 (N_9933,N_8615,N_8880);
nand U9934 (N_9934,N_8699,N_9093);
xor U9935 (N_9935,N_8569,N_8434);
nand U9936 (N_9936,N_8887,N_9085);
nor U9937 (N_9937,N_9568,N_9583);
nor U9938 (N_9938,N_9063,N_9062);
or U9939 (N_9939,N_9442,N_9511);
nand U9940 (N_9940,N_8851,N_9550);
or U9941 (N_9941,N_9311,N_8732);
and U9942 (N_9942,N_8757,N_9449);
nand U9943 (N_9943,N_8952,N_9167);
nand U9944 (N_9944,N_9368,N_8453);
and U9945 (N_9945,N_8454,N_8417);
and U9946 (N_9946,N_9172,N_9209);
and U9947 (N_9947,N_9196,N_9443);
nand U9948 (N_9948,N_8446,N_9143);
xnor U9949 (N_9949,N_8977,N_9476);
xor U9950 (N_9950,N_8448,N_9291);
xor U9951 (N_9951,N_8840,N_8684);
nor U9952 (N_9952,N_8804,N_8422);
and U9953 (N_9953,N_8899,N_9384);
or U9954 (N_9954,N_8923,N_8784);
nand U9955 (N_9955,N_8404,N_8654);
or U9956 (N_9956,N_8852,N_9124);
and U9957 (N_9957,N_9388,N_8841);
or U9958 (N_9958,N_9327,N_9531);
or U9959 (N_9959,N_9494,N_8504);
or U9960 (N_9960,N_9595,N_8901);
xnor U9961 (N_9961,N_9131,N_8905);
and U9962 (N_9962,N_8622,N_9260);
and U9963 (N_9963,N_8920,N_9455);
xnor U9964 (N_9964,N_9072,N_8597);
and U9965 (N_9965,N_8589,N_9367);
nor U9966 (N_9966,N_9352,N_8482);
or U9967 (N_9967,N_9075,N_8506);
and U9968 (N_9968,N_9322,N_9123);
or U9969 (N_9969,N_9221,N_8881);
nor U9970 (N_9970,N_8822,N_8982);
nand U9971 (N_9971,N_8862,N_8741);
nand U9972 (N_9972,N_9007,N_9562);
nand U9973 (N_9973,N_9473,N_9382);
and U9974 (N_9974,N_8768,N_8564);
nand U9975 (N_9975,N_9187,N_9472);
xnor U9976 (N_9976,N_9013,N_8420);
and U9977 (N_9977,N_9112,N_9264);
xnor U9978 (N_9978,N_8438,N_8563);
xnor U9979 (N_9979,N_9022,N_8828);
or U9980 (N_9980,N_8871,N_8639);
nand U9981 (N_9981,N_9292,N_8618);
xor U9982 (N_9982,N_9086,N_8891);
and U9983 (N_9983,N_9147,N_8470);
and U9984 (N_9984,N_8650,N_9340);
nor U9985 (N_9985,N_8996,N_8437);
or U9986 (N_9986,N_9066,N_9460);
xor U9987 (N_9987,N_8743,N_9010);
nand U9988 (N_9988,N_8636,N_8845);
nand U9989 (N_9989,N_9339,N_9405);
or U9990 (N_9990,N_9081,N_8988);
nor U9991 (N_9991,N_8410,N_8568);
nor U9992 (N_9992,N_8690,N_9432);
and U9993 (N_9993,N_8519,N_8976);
or U9994 (N_9994,N_8773,N_9082);
nand U9995 (N_9995,N_9348,N_9033);
nand U9996 (N_9996,N_8929,N_8497);
nor U9997 (N_9997,N_9176,N_9002);
and U9998 (N_9998,N_8738,N_8693);
nor U9999 (N_9999,N_9252,N_9498);
and U10000 (N_10000,N_8489,N_8457);
or U10001 (N_10001,N_8648,N_8630);
nand U10002 (N_10002,N_8848,N_8586);
and U10003 (N_10003,N_9142,N_9297);
nand U10004 (N_10004,N_9538,N_8908);
nor U10005 (N_10005,N_9095,N_9483);
nor U10006 (N_10006,N_8751,N_8581);
nor U10007 (N_10007,N_8525,N_9055);
nor U10008 (N_10008,N_9178,N_9092);
xnor U10009 (N_10009,N_9118,N_8847);
or U10010 (N_10010,N_8477,N_8893);
and U10011 (N_10011,N_9141,N_8865);
nor U10012 (N_10012,N_9213,N_8802);
nand U10013 (N_10013,N_9061,N_8964);
nand U10014 (N_10014,N_9507,N_9059);
nor U10015 (N_10015,N_9104,N_8555);
xor U10016 (N_10016,N_8808,N_9590);
xor U10017 (N_10017,N_9211,N_9155);
nand U10018 (N_10018,N_9579,N_9169);
nor U10019 (N_10019,N_8914,N_8514);
nor U10020 (N_10020,N_9139,N_8611);
xor U10021 (N_10021,N_8552,N_9330);
nor U10022 (N_10022,N_9079,N_9377);
and U10023 (N_10023,N_9047,N_8479);
nand U10024 (N_10024,N_8619,N_9199);
or U10025 (N_10025,N_8910,N_9157);
nand U10026 (N_10026,N_8821,N_9273);
or U10027 (N_10027,N_8819,N_9065);
or U10028 (N_10028,N_9186,N_9425);
nand U10029 (N_10029,N_9165,N_8942);
xnor U10030 (N_10030,N_8675,N_9174);
or U10031 (N_10031,N_9540,N_9561);
xor U10032 (N_10032,N_9357,N_8610);
or U10033 (N_10033,N_9284,N_9003);
and U10034 (N_10034,N_8626,N_9015);
and U10035 (N_10035,N_9480,N_8459);
and U10036 (N_10036,N_9020,N_9376);
and U10037 (N_10037,N_8450,N_8846);
and U10038 (N_10038,N_9127,N_9301);
and U10039 (N_10039,N_8627,N_9043);
or U10040 (N_10040,N_8925,N_9248);
and U10041 (N_10041,N_9126,N_8412);
or U10042 (N_10042,N_8711,N_9391);
nand U10043 (N_10043,N_8736,N_8970);
and U10044 (N_10044,N_8815,N_9341);
or U10045 (N_10045,N_8831,N_9505);
nor U10046 (N_10046,N_8682,N_9073);
xor U10047 (N_10047,N_9295,N_8883);
nand U10048 (N_10048,N_9042,N_8488);
and U10049 (N_10049,N_8895,N_9468);
nand U10050 (N_10050,N_8774,N_9584);
xnor U10051 (N_10051,N_9317,N_8992);
nand U10052 (N_10052,N_9076,N_8795);
nor U10053 (N_10053,N_9467,N_9371);
or U10054 (N_10054,N_8776,N_8478);
nand U10055 (N_10055,N_9336,N_9049);
or U10056 (N_10056,N_9390,N_8833);
nand U10057 (N_10057,N_8593,N_8960);
nor U10058 (N_10058,N_8733,N_8921);
nand U10059 (N_10059,N_9437,N_8903);
nand U10060 (N_10060,N_9034,N_8662);
and U10061 (N_10061,N_9351,N_8969);
nor U10062 (N_10062,N_8686,N_8523);
nand U10063 (N_10063,N_8934,N_8936);
or U10064 (N_10064,N_8867,N_8803);
nor U10065 (N_10065,N_9591,N_8607);
nand U10066 (N_10066,N_9056,N_8767);
or U10067 (N_10067,N_8990,N_8540);
nand U10068 (N_10068,N_9133,N_9250);
or U10069 (N_10069,N_8924,N_8807);
xnor U10070 (N_10070,N_9381,N_9099);
nor U10071 (N_10071,N_8951,N_8613);
nand U10072 (N_10072,N_8620,N_8429);
xor U10073 (N_10073,N_8993,N_8878);
nor U10074 (N_10074,N_8672,N_9580);
and U10075 (N_10075,N_9254,N_9303);
and U10076 (N_10076,N_9019,N_9362);
xor U10077 (N_10077,N_9567,N_8998);
nand U10078 (N_10078,N_8419,N_9559);
xnor U10079 (N_10079,N_8806,N_9361);
xnor U10080 (N_10080,N_9401,N_8717);
and U10081 (N_10081,N_8875,N_8487);
xnor U10082 (N_10082,N_8612,N_9520);
and U10083 (N_10083,N_8712,N_8526);
and U10084 (N_10084,N_8436,N_8737);
nand U10085 (N_10085,N_8527,N_8747);
xnor U10086 (N_10086,N_8596,N_8793);
nand U10087 (N_10087,N_8981,N_9551);
nand U10088 (N_10088,N_9582,N_9233);
and U10089 (N_10089,N_8825,N_8832);
xor U10090 (N_10090,N_8444,N_9098);
xor U10091 (N_10091,N_8592,N_8710);
and U10092 (N_10092,N_9532,N_9421);
nor U10093 (N_10093,N_8915,N_9474);
nor U10094 (N_10094,N_9566,N_8602);
xnor U10095 (N_10095,N_9298,N_9516);
nand U10096 (N_10096,N_8772,N_8580);
xor U10097 (N_10097,N_9326,N_8724);
xor U10098 (N_10098,N_9102,N_8694);
or U10099 (N_10099,N_8730,N_9413);
or U10100 (N_10100,N_9453,N_9183);
xnor U10101 (N_10101,N_8941,N_8739);
nor U10102 (N_10102,N_8947,N_8967);
nor U10103 (N_10103,N_9542,N_9041);
and U10104 (N_10104,N_8633,N_8971);
nand U10105 (N_10105,N_8708,N_9228);
and U10106 (N_10106,N_8520,N_9353);
nand U10107 (N_10107,N_8702,N_8820);
nor U10108 (N_10108,N_8763,N_9191);
nand U10109 (N_10109,N_9168,N_9392);
or U10110 (N_10110,N_8927,N_8435);
and U10111 (N_10111,N_8430,N_9411);
nand U10112 (N_10112,N_9386,N_8659);
nand U10113 (N_10113,N_8705,N_8859);
and U10114 (N_10114,N_8476,N_8735);
or U10115 (N_10115,N_9265,N_8676);
nand U10116 (N_10116,N_8917,N_8649);
xor U10117 (N_10117,N_9216,N_9110);
xnor U10118 (N_10118,N_9270,N_9129);
nand U10119 (N_10119,N_8426,N_8697);
nand U10120 (N_10120,N_8617,N_8573);
xnor U10121 (N_10121,N_9533,N_8858);
or U10122 (N_10122,N_8600,N_8781);
xor U10123 (N_10123,N_9419,N_8562);
xnor U10124 (N_10124,N_9347,N_9415);
or U10125 (N_10125,N_8939,N_9571);
xnor U10126 (N_10126,N_8853,N_8583);
and U10127 (N_10127,N_8646,N_9389);
or U10128 (N_10128,N_8405,N_9219);
nor U10129 (N_10129,N_8665,N_8722);
nand U10130 (N_10130,N_9343,N_8989);
and U10131 (N_10131,N_9313,N_9158);
and U10132 (N_10132,N_8570,N_9109);
or U10133 (N_10133,N_8407,N_9045);
and U10134 (N_10134,N_9385,N_9592);
and U10135 (N_10135,N_8565,N_9293);
xor U10136 (N_10136,N_9508,N_9338);
and U10137 (N_10137,N_8673,N_9035);
nand U10138 (N_10138,N_8995,N_9418);
nor U10139 (N_10139,N_9266,N_9576);
nand U10140 (N_10140,N_9156,N_8500);
xor U10141 (N_10141,N_9350,N_9398);
or U10142 (N_10142,N_9526,N_9077);
nor U10143 (N_10143,N_9366,N_8786);
and U10144 (N_10144,N_8559,N_8499);
nor U10145 (N_10145,N_9012,N_8463);
or U10146 (N_10146,N_9573,N_9289);
and U10147 (N_10147,N_9036,N_8897);
xor U10148 (N_10148,N_8809,N_9372);
or U10149 (N_10149,N_8762,N_9037);
nor U10150 (N_10150,N_8493,N_9422);
nand U10151 (N_10151,N_9555,N_9068);
and U10152 (N_10152,N_8818,N_8979);
xor U10153 (N_10153,N_9175,N_9231);
nor U10154 (N_10154,N_9402,N_9454);
and U10155 (N_10155,N_9184,N_9255);
and U10156 (N_10156,N_9283,N_8856);
and U10157 (N_10157,N_8558,N_8959);
nand U10158 (N_10158,N_8545,N_8882);
and U10159 (N_10159,N_8926,N_8485);
nor U10160 (N_10160,N_8861,N_8719);
nor U10161 (N_10161,N_8787,N_9360);
nor U10162 (N_10162,N_9598,N_8889);
nand U10163 (N_10163,N_8669,N_8456);
xor U10164 (N_10164,N_8688,N_9462);
and U10165 (N_10165,N_9243,N_9355);
xor U10166 (N_10166,N_9300,N_9496);
nand U10167 (N_10167,N_9393,N_9495);
xnor U10168 (N_10168,N_8975,N_8495);
and U10169 (N_10169,N_8827,N_9031);
and U10170 (N_10170,N_9435,N_9146);
and U10171 (N_10171,N_9380,N_8549);
or U10172 (N_10172,N_8474,N_8460);
nand U10173 (N_10173,N_8944,N_9530);
or U10174 (N_10174,N_9145,N_9337);
xor U10175 (N_10175,N_8729,N_9504);
xor U10176 (N_10176,N_8609,N_9204);
and U10177 (N_10177,N_8681,N_9586);
xor U10178 (N_10178,N_8849,N_8461);
and U10179 (N_10179,N_8421,N_8532);
nand U10180 (N_10180,N_9541,N_9438);
nor U10181 (N_10181,N_9588,N_8466);
xnor U10182 (N_10182,N_9138,N_9441);
xnor U10183 (N_10183,N_8779,N_8635);
xnor U10184 (N_10184,N_9440,N_9410);
nor U10185 (N_10185,N_8869,N_9431);
nor U10186 (N_10186,N_8413,N_9345);
nand U10187 (N_10187,N_9456,N_9286);
or U10188 (N_10188,N_8946,N_8469);
or U10189 (N_10189,N_9397,N_9513);
or U10190 (N_10190,N_9097,N_9011);
nor U10191 (N_10191,N_9543,N_9032);
nor U10192 (N_10192,N_8765,N_8720);
nand U10193 (N_10193,N_9132,N_8678);
or U10194 (N_10194,N_8963,N_8443);
or U10195 (N_10195,N_9237,N_8965);
xnor U10196 (N_10196,N_9404,N_8464);
or U10197 (N_10197,N_9354,N_9188);
xor U10198 (N_10198,N_8911,N_8492);
or U10199 (N_10199,N_9113,N_9529);
xnor U10200 (N_10200,N_8468,N_8498);
nor U10201 (N_10201,N_9375,N_9586);
nand U10202 (N_10202,N_8694,N_8423);
xor U10203 (N_10203,N_8761,N_9126);
nor U10204 (N_10204,N_8628,N_8449);
xor U10205 (N_10205,N_8666,N_8814);
xnor U10206 (N_10206,N_8445,N_9121);
nor U10207 (N_10207,N_9422,N_9299);
nor U10208 (N_10208,N_8828,N_8671);
or U10209 (N_10209,N_9111,N_8779);
nand U10210 (N_10210,N_8662,N_9530);
xor U10211 (N_10211,N_8964,N_8974);
and U10212 (N_10212,N_9401,N_8642);
xor U10213 (N_10213,N_9510,N_8551);
nand U10214 (N_10214,N_8535,N_9277);
xor U10215 (N_10215,N_9199,N_8488);
and U10216 (N_10216,N_9291,N_9547);
or U10217 (N_10217,N_8494,N_8441);
nand U10218 (N_10218,N_9419,N_8851);
nor U10219 (N_10219,N_8505,N_8952);
nand U10220 (N_10220,N_9062,N_8770);
nand U10221 (N_10221,N_9064,N_8922);
and U10222 (N_10222,N_8493,N_8986);
xnor U10223 (N_10223,N_9072,N_8677);
nor U10224 (N_10224,N_8812,N_8977);
nor U10225 (N_10225,N_9006,N_9518);
xnor U10226 (N_10226,N_9189,N_9133);
nand U10227 (N_10227,N_8903,N_9115);
xnor U10228 (N_10228,N_8781,N_8861);
or U10229 (N_10229,N_9240,N_9472);
or U10230 (N_10230,N_9268,N_8418);
nor U10231 (N_10231,N_9155,N_9551);
and U10232 (N_10232,N_9117,N_8562);
xnor U10233 (N_10233,N_8493,N_8925);
xnor U10234 (N_10234,N_8850,N_8801);
nand U10235 (N_10235,N_8442,N_9336);
nand U10236 (N_10236,N_9122,N_9387);
nor U10237 (N_10237,N_9007,N_8738);
xor U10238 (N_10238,N_9273,N_8522);
nand U10239 (N_10239,N_8636,N_8882);
nor U10240 (N_10240,N_9072,N_8838);
and U10241 (N_10241,N_8403,N_9599);
xnor U10242 (N_10242,N_9136,N_8691);
or U10243 (N_10243,N_9153,N_9302);
nor U10244 (N_10244,N_9071,N_8454);
nor U10245 (N_10245,N_9299,N_8725);
and U10246 (N_10246,N_9262,N_9222);
or U10247 (N_10247,N_8491,N_9240);
xnor U10248 (N_10248,N_9337,N_9005);
xor U10249 (N_10249,N_9288,N_9399);
nand U10250 (N_10250,N_8663,N_8993);
and U10251 (N_10251,N_8667,N_8817);
xor U10252 (N_10252,N_9109,N_9320);
xnor U10253 (N_10253,N_8507,N_9455);
nor U10254 (N_10254,N_8725,N_8636);
or U10255 (N_10255,N_9438,N_8612);
nand U10256 (N_10256,N_9065,N_8446);
nor U10257 (N_10257,N_8701,N_9314);
nand U10258 (N_10258,N_8491,N_9166);
nand U10259 (N_10259,N_8993,N_9446);
and U10260 (N_10260,N_8689,N_9542);
nor U10261 (N_10261,N_9347,N_9555);
and U10262 (N_10262,N_9045,N_9356);
nor U10263 (N_10263,N_8812,N_9414);
or U10264 (N_10264,N_8976,N_9348);
or U10265 (N_10265,N_9281,N_8552);
nand U10266 (N_10266,N_8560,N_9353);
nor U10267 (N_10267,N_9340,N_9535);
nor U10268 (N_10268,N_9486,N_8902);
xor U10269 (N_10269,N_9368,N_8773);
or U10270 (N_10270,N_8589,N_9475);
or U10271 (N_10271,N_9393,N_9141);
and U10272 (N_10272,N_8745,N_8402);
nand U10273 (N_10273,N_9382,N_8559);
nor U10274 (N_10274,N_8758,N_8921);
and U10275 (N_10275,N_8915,N_9595);
xor U10276 (N_10276,N_9059,N_8436);
xor U10277 (N_10277,N_8682,N_9291);
xnor U10278 (N_10278,N_8635,N_9228);
xnor U10279 (N_10279,N_9515,N_9311);
and U10280 (N_10280,N_8649,N_9366);
xor U10281 (N_10281,N_8543,N_9237);
nor U10282 (N_10282,N_8761,N_8923);
nor U10283 (N_10283,N_9412,N_8667);
nor U10284 (N_10284,N_9577,N_9288);
or U10285 (N_10285,N_8622,N_9370);
nand U10286 (N_10286,N_8412,N_8935);
nor U10287 (N_10287,N_8911,N_8607);
nand U10288 (N_10288,N_8620,N_9040);
nor U10289 (N_10289,N_9433,N_9152);
or U10290 (N_10290,N_9302,N_8840);
xor U10291 (N_10291,N_8829,N_9050);
and U10292 (N_10292,N_8434,N_8759);
nor U10293 (N_10293,N_8972,N_8591);
xor U10294 (N_10294,N_8463,N_8603);
and U10295 (N_10295,N_8480,N_8878);
or U10296 (N_10296,N_8427,N_8619);
and U10297 (N_10297,N_9292,N_9204);
nor U10298 (N_10298,N_9099,N_8649);
xor U10299 (N_10299,N_8940,N_9271);
xor U10300 (N_10300,N_8449,N_8613);
nor U10301 (N_10301,N_9471,N_8582);
nand U10302 (N_10302,N_9508,N_9092);
xnor U10303 (N_10303,N_8802,N_8775);
nor U10304 (N_10304,N_8915,N_9504);
nand U10305 (N_10305,N_8866,N_8887);
nand U10306 (N_10306,N_9392,N_9483);
or U10307 (N_10307,N_8422,N_9385);
xnor U10308 (N_10308,N_9019,N_8921);
or U10309 (N_10309,N_9245,N_9090);
nand U10310 (N_10310,N_8631,N_8706);
or U10311 (N_10311,N_9158,N_8651);
nand U10312 (N_10312,N_9007,N_8945);
or U10313 (N_10313,N_9223,N_8443);
or U10314 (N_10314,N_8787,N_9537);
and U10315 (N_10315,N_9205,N_8651);
nor U10316 (N_10316,N_9027,N_8993);
and U10317 (N_10317,N_8685,N_9010);
and U10318 (N_10318,N_9546,N_9083);
nand U10319 (N_10319,N_8667,N_8738);
or U10320 (N_10320,N_8441,N_8421);
xnor U10321 (N_10321,N_9055,N_8683);
and U10322 (N_10322,N_9139,N_9453);
or U10323 (N_10323,N_9304,N_8452);
and U10324 (N_10324,N_8607,N_9164);
xor U10325 (N_10325,N_9174,N_8572);
xor U10326 (N_10326,N_8696,N_8803);
nand U10327 (N_10327,N_9127,N_9244);
or U10328 (N_10328,N_8539,N_8641);
nand U10329 (N_10329,N_8444,N_9565);
or U10330 (N_10330,N_8805,N_8637);
and U10331 (N_10331,N_8822,N_9129);
nor U10332 (N_10332,N_9579,N_8486);
xor U10333 (N_10333,N_9370,N_9340);
or U10334 (N_10334,N_9408,N_9339);
nand U10335 (N_10335,N_9272,N_8537);
and U10336 (N_10336,N_9425,N_9111);
xnor U10337 (N_10337,N_8507,N_9484);
nand U10338 (N_10338,N_8985,N_9155);
nor U10339 (N_10339,N_9456,N_9466);
nor U10340 (N_10340,N_9022,N_9328);
nor U10341 (N_10341,N_8711,N_8466);
xnor U10342 (N_10342,N_9215,N_8407);
or U10343 (N_10343,N_9443,N_8789);
nand U10344 (N_10344,N_8903,N_8662);
nand U10345 (N_10345,N_9402,N_8950);
nor U10346 (N_10346,N_8441,N_8833);
and U10347 (N_10347,N_9014,N_9513);
nand U10348 (N_10348,N_9387,N_9090);
nand U10349 (N_10349,N_8872,N_9238);
nand U10350 (N_10350,N_9449,N_8456);
nand U10351 (N_10351,N_9241,N_9156);
or U10352 (N_10352,N_9089,N_9143);
and U10353 (N_10353,N_9463,N_9567);
or U10354 (N_10354,N_9529,N_9559);
xor U10355 (N_10355,N_9208,N_9534);
nor U10356 (N_10356,N_9105,N_8764);
nand U10357 (N_10357,N_9028,N_8665);
nor U10358 (N_10358,N_8680,N_8637);
nor U10359 (N_10359,N_9007,N_8540);
or U10360 (N_10360,N_9136,N_8888);
xor U10361 (N_10361,N_9208,N_9044);
xor U10362 (N_10362,N_9350,N_9237);
xor U10363 (N_10363,N_8512,N_9154);
or U10364 (N_10364,N_9367,N_8774);
nor U10365 (N_10365,N_8834,N_8887);
nor U10366 (N_10366,N_9009,N_9205);
nand U10367 (N_10367,N_9229,N_8465);
xnor U10368 (N_10368,N_9480,N_9311);
nor U10369 (N_10369,N_8766,N_9275);
or U10370 (N_10370,N_8686,N_9283);
nand U10371 (N_10371,N_9385,N_9007);
or U10372 (N_10372,N_9430,N_9427);
or U10373 (N_10373,N_8644,N_8975);
nor U10374 (N_10374,N_9315,N_9560);
nand U10375 (N_10375,N_8774,N_8503);
and U10376 (N_10376,N_8737,N_8699);
nor U10377 (N_10377,N_8455,N_9487);
or U10378 (N_10378,N_8547,N_8847);
or U10379 (N_10379,N_9514,N_8437);
or U10380 (N_10380,N_9359,N_8689);
xor U10381 (N_10381,N_8424,N_9197);
nand U10382 (N_10382,N_8474,N_9525);
xnor U10383 (N_10383,N_8973,N_8854);
and U10384 (N_10384,N_9377,N_8544);
and U10385 (N_10385,N_9194,N_9066);
or U10386 (N_10386,N_8767,N_9354);
nor U10387 (N_10387,N_9509,N_8964);
nor U10388 (N_10388,N_9202,N_9152);
xor U10389 (N_10389,N_9422,N_9592);
and U10390 (N_10390,N_8462,N_9584);
nand U10391 (N_10391,N_8866,N_8459);
nor U10392 (N_10392,N_9179,N_8908);
nand U10393 (N_10393,N_8420,N_8919);
or U10394 (N_10394,N_9345,N_9477);
nand U10395 (N_10395,N_9460,N_9254);
and U10396 (N_10396,N_8454,N_8405);
nor U10397 (N_10397,N_9271,N_8830);
or U10398 (N_10398,N_9361,N_8924);
and U10399 (N_10399,N_8765,N_9112);
and U10400 (N_10400,N_9367,N_9354);
and U10401 (N_10401,N_9243,N_9159);
or U10402 (N_10402,N_9167,N_8621);
nand U10403 (N_10403,N_9525,N_9352);
and U10404 (N_10404,N_8648,N_8771);
nand U10405 (N_10405,N_9018,N_8892);
xnor U10406 (N_10406,N_9046,N_9477);
nor U10407 (N_10407,N_9154,N_8900);
xnor U10408 (N_10408,N_9544,N_9010);
nand U10409 (N_10409,N_9244,N_9594);
nor U10410 (N_10410,N_9563,N_9280);
nor U10411 (N_10411,N_9193,N_8950);
and U10412 (N_10412,N_8749,N_9003);
and U10413 (N_10413,N_8529,N_9373);
or U10414 (N_10414,N_8442,N_9507);
nor U10415 (N_10415,N_9351,N_9371);
or U10416 (N_10416,N_8613,N_8525);
nor U10417 (N_10417,N_9428,N_8421);
xnor U10418 (N_10418,N_8679,N_9109);
nor U10419 (N_10419,N_9132,N_8428);
nand U10420 (N_10420,N_9476,N_8883);
xnor U10421 (N_10421,N_8642,N_9338);
or U10422 (N_10422,N_9326,N_9012);
nor U10423 (N_10423,N_8949,N_9525);
nor U10424 (N_10424,N_9154,N_9312);
xor U10425 (N_10425,N_9451,N_9227);
nor U10426 (N_10426,N_8572,N_9451);
nor U10427 (N_10427,N_8787,N_8723);
and U10428 (N_10428,N_9443,N_9424);
xor U10429 (N_10429,N_8584,N_9425);
nand U10430 (N_10430,N_8509,N_9445);
nor U10431 (N_10431,N_9447,N_9420);
or U10432 (N_10432,N_9584,N_8938);
and U10433 (N_10433,N_8602,N_8533);
nor U10434 (N_10434,N_9258,N_9378);
xor U10435 (N_10435,N_8709,N_8471);
or U10436 (N_10436,N_8944,N_8551);
and U10437 (N_10437,N_8990,N_9584);
or U10438 (N_10438,N_9209,N_9099);
and U10439 (N_10439,N_8891,N_9295);
xnor U10440 (N_10440,N_9477,N_9563);
nand U10441 (N_10441,N_9140,N_9106);
nor U10442 (N_10442,N_9410,N_9280);
or U10443 (N_10443,N_9490,N_9146);
or U10444 (N_10444,N_9262,N_9363);
or U10445 (N_10445,N_8790,N_9497);
xnor U10446 (N_10446,N_9426,N_9528);
or U10447 (N_10447,N_9564,N_9006);
or U10448 (N_10448,N_8997,N_8472);
or U10449 (N_10449,N_9187,N_9388);
or U10450 (N_10450,N_9136,N_9089);
xnor U10451 (N_10451,N_8795,N_9020);
nand U10452 (N_10452,N_8880,N_8826);
nor U10453 (N_10453,N_8611,N_8606);
or U10454 (N_10454,N_8506,N_9497);
nand U10455 (N_10455,N_9281,N_9157);
or U10456 (N_10456,N_8759,N_8455);
or U10457 (N_10457,N_8476,N_9504);
and U10458 (N_10458,N_8860,N_8561);
nor U10459 (N_10459,N_9167,N_8495);
nand U10460 (N_10460,N_8685,N_9027);
and U10461 (N_10461,N_8914,N_9124);
xnor U10462 (N_10462,N_9394,N_9206);
or U10463 (N_10463,N_9533,N_8443);
and U10464 (N_10464,N_8567,N_9285);
nand U10465 (N_10465,N_9225,N_9052);
or U10466 (N_10466,N_9215,N_8527);
nand U10467 (N_10467,N_9484,N_9111);
and U10468 (N_10468,N_8700,N_9462);
or U10469 (N_10469,N_8918,N_8661);
nand U10470 (N_10470,N_8739,N_9078);
nor U10471 (N_10471,N_9009,N_8463);
and U10472 (N_10472,N_9440,N_9009);
nor U10473 (N_10473,N_9324,N_9087);
or U10474 (N_10474,N_8778,N_8674);
nand U10475 (N_10475,N_8788,N_9242);
and U10476 (N_10476,N_9216,N_9013);
and U10477 (N_10477,N_8668,N_8416);
nor U10478 (N_10478,N_9289,N_9527);
and U10479 (N_10479,N_9416,N_8629);
and U10480 (N_10480,N_8615,N_9207);
and U10481 (N_10481,N_8667,N_8793);
nand U10482 (N_10482,N_9107,N_9032);
nand U10483 (N_10483,N_8653,N_9037);
and U10484 (N_10484,N_9170,N_9402);
nor U10485 (N_10485,N_8535,N_8943);
nand U10486 (N_10486,N_8402,N_8896);
xnor U10487 (N_10487,N_9355,N_9172);
or U10488 (N_10488,N_9519,N_8678);
nand U10489 (N_10489,N_9262,N_9277);
and U10490 (N_10490,N_8502,N_9594);
nor U10491 (N_10491,N_9049,N_9280);
nor U10492 (N_10492,N_9473,N_9423);
or U10493 (N_10493,N_8946,N_8828);
or U10494 (N_10494,N_8759,N_8888);
and U10495 (N_10495,N_8738,N_8613);
or U10496 (N_10496,N_9506,N_8638);
nor U10497 (N_10497,N_8988,N_8514);
xnor U10498 (N_10498,N_9404,N_9384);
xor U10499 (N_10499,N_8990,N_9382);
xnor U10500 (N_10500,N_8504,N_8907);
or U10501 (N_10501,N_8598,N_8454);
xnor U10502 (N_10502,N_9081,N_8691);
or U10503 (N_10503,N_9340,N_8922);
and U10504 (N_10504,N_9388,N_8514);
and U10505 (N_10505,N_8608,N_8987);
xor U10506 (N_10506,N_8650,N_8780);
or U10507 (N_10507,N_9013,N_8698);
xnor U10508 (N_10508,N_8785,N_9053);
and U10509 (N_10509,N_8963,N_9072);
xnor U10510 (N_10510,N_9463,N_9299);
xnor U10511 (N_10511,N_8900,N_9524);
nand U10512 (N_10512,N_8918,N_9329);
nor U10513 (N_10513,N_9015,N_9443);
nor U10514 (N_10514,N_9554,N_8527);
xnor U10515 (N_10515,N_8688,N_9498);
nand U10516 (N_10516,N_8778,N_8642);
nand U10517 (N_10517,N_8492,N_8990);
nand U10518 (N_10518,N_8606,N_9096);
nand U10519 (N_10519,N_8965,N_8495);
nand U10520 (N_10520,N_9410,N_8734);
nor U10521 (N_10521,N_9432,N_8826);
and U10522 (N_10522,N_8415,N_8503);
xor U10523 (N_10523,N_8838,N_9555);
and U10524 (N_10524,N_8991,N_8459);
nand U10525 (N_10525,N_8499,N_9177);
or U10526 (N_10526,N_9121,N_8704);
and U10527 (N_10527,N_8577,N_9012);
or U10528 (N_10528,N_9458,N_8896);
and U10529 (N_10529,N_8455,N_8558);
and U10530 (N_10530,N_9435,N_9459);
nand U10531 (N_10531,N_9494,N_9364);
and U10532 (N_10532,N_9413,N_9232);
nand U10533 (N_10533,N_8779,N_9354);
nand U10534 (N_10534,N_8792,N_8459);
nor U10535 (N_10535,N_8654,N_8880);
nor U10536 (N_10536,N_8937,N_8648);
nand U10537 (N_10537,N_8421,N_9534);
xor U10538 (N_10538,N_8684,N_8874);
nand U10539 (N_10539,N_8836,N_9316);
nand U10540 (N_10540,N_9356,N_8537);
nor U10541 (N_10541,N_9011,N_9127);
nand U10542 (N_10542,N_8671,N_8542);
nand U10543 (N_10543,N_8724,N_9021);
nor U10544 (N_10544,N_8661,N_8532);
nand U10545 (N_10545,N_9053,N_9374);
and U10546 (N_10546,N_9410,N_9498);
and U10547 (N_10547,N_8703,N_8826);
and U10548 (N_10548,N_9102,N_9208);
nand U10549 (N_10549,N_9480,N_8725);
or U10550 (N_10550,N_8415,N_9174);
nand U10551 (N_10551,N_8764,N_8456);
nand U10552 (N_10552,N_9245,N_8804);
nand U10553 (N_10553,N_8759,N_9475);
xnor U10554 (N_10554,N_8921,N_8947);
and U10555 (N_10555,N_9161,N_8841);
or U10556 (N_10556,N_9485,N_8580);
nor U10557 (N_10557,N_8989,N_8522);
nand U10558 (N_10558,N_9348,N_8575);
xnor U10559 (N_10559,N_9168,N_9134);
or U10560 (N_10560,N_8562,N_8979);
nand U10561 (N_10561,N_9551,N_9073);
nor U10562 (N_10562,N_8821,N_8596);
xor U10563 (N_10563,N_8739,N_8499);
nand U10564 (N_10564,N_9080,N_9338);
nand U10565 (N_10565,N_8663,N_9344);
xor U10566 (N_10566,N_9312,N_9152);
nor U10567 (N_10567,N_9136,N_9489);
nor U10568 (N_10568,N_9037,N_9567);
and U10569 (N_10569,N_8580,N_8423);
nand U10570 (N_10570,N_9498,N_8431);
or U10571 (N_10571,N_9319,N_8878);
or U10572 (N_10572,N_8955,N_9511);
nor U10573 (N_10573,N_9069,N_9035);
nor U10574 (N_10574,N_8863,N_8445);
and U10575 (N_10575,N_8417,N_8868);
or U10576 (N_10576,N_9033,N_8553);
xnor U10577 (N_10577,N_9168,N_9342);
and U10578 (N_10578,N_8758,N_8427);
and U10579 (N_10579,N_9596,N_9282);
nand U10580 (N_10580,N_9452,N_9310);
nor U10581 (N_10581,N_9398,N_9525);
nor U10582 (N_10582,N_8438,N_9017);
or U10583 (N_10583,N_8945,N_9444);
xnor U10584 (N_10584,N_9046,N_9086);
nand U10585 (N_10585,N_8848,N_8934);
xnor U10586 (N_10586,N_8501,N_8629);
or U10587 (N_10587,N_8643,N_8756);
and U10588 (N_10588,N_8440,N_8812);
nand U10589 (N_10589,N_8741,N_8484);
or U10590 (N_10590,N_8573,N_9107);
xnor U10591 (N_10591,N_9225,N_8649);
xnor U10592 (N_10592,N_9509,N_8796);
nand U10593 (N_10593,N_8719,N_9223);
or U10594 (N_10594,N_8496,N_9280);
xnor U10595 (N_10595,N_9570,N_9059);
or U10596 (N_10596,N_8726,N_9462);
nand U10597 (N_10597,N_9487,N_9001);
nand U10598 (N_10598,N_9470,N_8663);
nor U10599 (N_10599,N_8423,N_8888);
or U10600 (N_10600,N_9375,N_8605);
xnor U10601 (N_10601,N_9287,N_9506);
nor U10602 (N_10602,N_8648,N_9490);
nor U10603 (N_10603,N_9298,N_8863);
nor U10604 (N_10604,N_9474,N_8926);
and U10605 (N_10605,N_8989,N_8967);
nor U10606 (N_10606,N_9207,N_9163);
or U10607 (N_10607,N_9309,N_8896);
or U10608 (N_10608,N_8944,N_9499);
or U10609 (N_10609,N_8899,N_9004);
nand U10610 (N_10610,N_9148,N_9430);
nor U10611 (N_10611,N_9156,N_8833);
and U10612 (N_10612,N_9118,N_9367);
and U10613 (N_10613,N_8756,N_8670);
nand U10614 (N_10614,N_9198,N_9237);
and U10615 (N_10615,N_8936,N_9095);
and U10616 (N_10616,N_9274,N_8555);
or U10617 (N_10617,N_8995,N_8450);
xnor U10618 (N_10618,N_8985,N_9188);
nand U10619 (N_10619,N_9548,N_9281);
nand U10620 (N_10620,N_8402,N_9447);
xor U10621 (N_10621,N_9366,N_8951);
or U10622 (N_10622,N_8891,N_9352);
xnor U10623 (N_10623,N_8828,N_9596);
or U10624 (N_10624,N_8436,N_9546);
nor U10625 (N_10625,N_8947,N_8754);
nor U10626 (N_10626,N_8849,N_8477);
and U10627 (N_10627,N_8734,N_8730);
and U10628 (N_10628,N_8835,N_9101);
nor U10629 (N_10629,N_9486,N_8764);
or U10630 (N_10630,N_8820,N_8538);
or U10631 (N_10631,N_8496,N_9480);
and U10632 (N_10632,N_8571,N_8678);
or U10633 (N_10633,N_8614,N_8456);
nor U10634 (N_10634,N_8514,N_9337);
xor U10635 (N_10635,N_8588,N_9206);
and U10636 (N_10636,N_9507,N_8413);
xor U10637 (N_10637,N_8663,N_9595);
and U10638 (N_10638,N_8942,N_9465);
and U10639 (N_10639,N_8507,N_8780);
and U10640 (N_10640,N_8781,N_8883);
xnor U10641 (N_10641,N_9012,N_8575);
nor U10642 (N_10642,N_9512,N_9075);
or U10643 (N_10643,N_9519,N_9016);
nand U10644 (N_10644,N_8678,N_8798);
nor U10645 (N_10645,N_8923,N_9270);
or U10646 (N_10646,N_9085,N_9506);
or U10647 (N_10647,N_9219,N_8731);
or U10648 (N_10648,N_9402,N_9346);
nor U10649 (N_10649,N_9060,N_8942);
xnor U10650 (N_10650,N_9122,N_9075);
xnor U10651 (N_10651,N_8730,N_9453);
nor U10652 (N_10652,N_9521,N_8487);
or U10653 (N_10653,N_8904,N_8935);
xor U10654 (N_10654,N_8936,N_8718);
and U10655 (N_10655,N_8759,N_8879);
or U10656 (N_10656,N_8925,N_9347);
or U10657 (N_10657,N_8784,N_8803);
nand U10658 (N_10658,N_9061,N_8710);
or U10659 (N_10659,N_9522,N_8870);
nand U10660 (N_10660,N_9585,N_8445);
and U10661 (N_10661,N_8493,N_9481);
and U10662 (N_10662,N_9577,N_9139);
and U10663 (N_10663,N_8745,N_9356);
xnor U10664 (N_10664,N_8573,N_9407);
xor U10665 (N_10665,N_9466,N_8737);
or U10666 (N_10666,N_9032,N_9169);
nand U10667 (N_10667,N_9234,N_9520);
or U10668 (N_10668,N_9519,N_9577);
or U10669 (N_10669,N_9130,N_9002);
or U10670 (N_10670,N_9252,N_8690);
or U10671 (N_10671,N_9503,N_8948);
and U10672 (N_10672,N_9116,N_8733);
nand U10673 (N_10673,N_9112,N_8967);
or U10674 (N_10674,N_8985,N_8634);
xnor U10675 (N_10675,N_9450,N_9139);
nand U10676 (N_10676,N_8673,N_9304);
or U10677 (N_10677,N_8975,N_8541);
or U10678 (N_10678,N_9236,N_8592);
nor U10679 (N_10679,N_8557,N_9207);
nand U10680 (N_10680,N_8792,N_8698);
and U10681 (N_10681,N_8634,N_8669);
xor U10682 (N_10682,N_9024,N_9215);
or U10683 (N_10683,N_9531,N_9139);
and U10684 (N_10684,N_8456,N_8659);
nand U10685 (N_10685,N_9424,N_8894);
nor U10686 (N_10686,N_8546,N_8820);
nor U10687 (N_10687,N_8861,N_8779);
nor U10688 (N_10688,N_8571,N_9009);
xor U10689 (N_10689,N_9372,N_8696);
and U10690 (N_10690,N_9486,N_9144);
xor U10691 (N_10691,N_9290,N_8951);
and U10692 (N_10692,N_9173,N_8975);
xnor U10693 (N_10693,N_8615,N_9345);
nor U10694 (N_10694,N_8532,N_8769);
or U10695 (N_10695,N_9409,N_8608);
and U10696 (N_10696,N_9415,N_9291);
nor U10697 (N_10697,N_9500,N_8433);
and U10698 (N_10698,N_9091,N_8544);
nor U10699 (N_10699,N_8979,N_9201);
or U10700 (N_10700,N_9052,N_8455);
xnor U10701 (N_10701,N_8415,N_8946);
and U10702 (N_10702,N_9022,N_9243);
or U10703 (N_10703,N_8654,N_8466);
nor U10704 (N_10704,N_8415,N_8698);
and U10705 (N_10705,N_8853,N_8889);
nand U10706 (N_10706,N_9450,N_8572);
nand U10707 (N_10707,N_8760,N_9433);
nor U10708 (N_10708,N_9055,N_8465);
or U10709 (N_10709,N_8901,N_9113);
and U10710 (N_10710,N_9171,N_9114);
and U10711 (N_10711,N_8802,N_9574);
nor U10712 (N_10712,N_9412,N_8628);
nand U10713 (N_10713,N_8419,N_8600);
nand U10714 (N_10714,N_8471,N_8856);
xnor U10715 (N_10715,N_8775,N_9243);
nor U10716 (N_10716,N_9466,N_9017);
xnor U10717 (N_10717,N_9499,N_9244);
xnor U10718 (N_10718,N_8429,N_8950);
nor U10719 (N_10719,N_8985,N_9013);
xnor U10720 (N_10720,N_9006,N_8550);
and U10721 (N_10721,N_8651,N_8709);
nand U10722 (N_10722,N_9071,N_9089);
nor U10723 (N_10723,N_9566,N_8799);
nand U10724 (N_10724,N_9148,N_9352);
xor U10725 (N_10725,N_8637,N_9333);
and U10726 (N_10726,N_9284,N_9038);
xor U10727 (N_10727,N_8596,N_9040);
nor U10728 (N_10728,N_8811,N_9022);
nor U10729 (N_10729,N_8897,N_8889);
nor U10730 (N_10730,N_8542,N_9046);
or U10731 (N_10731,N_9393,N_8624);
xor U10732 (N_10732,N_8534,N_9218);
xnor U10733 (N_10733,N_9307,N_8892);
and U10734 (N_10734,N_8693,N_9591);
nor U10735 (N_10735,N_9468,N_9254);
nand U10736 (N_10736,N_8589,N_9432);
nor U10737 (N_10737,N_8894,N_9014);
and U10738 (N_10738,N_9529,N_8857);
nand U10739 (N_10739,N_8875,N_9015);
and U10740 (N_10740,N_8826,N_9310);
nand U10741 (N_10741,N_8847,N_9557);
xor U10742 (N_10742,N_8535,N_8563);
xor U10743 (N_10743,N_8507,N_8855);
nor U10744 (N_10744,N_9083,N_8482);
nand U10745 (N_10745,N_9372,N_9473);
nand U10746 (N_10746,N_8609,N_8749);
nor U10747 (N_10747,N_9414,N_9340);
or U10748 (N_10748,N_8521,N_9188);
nand U10749 (N_10749,N_9144,N_9466);
nand U10750 (N_10750,N_8511,N_8964);
or U10751 (N_10751,N_9158,N_9144);
nand U10752 (N_10752,N_8624,N_9579);
or U10753 (N_10753,N_8659,N_9483);
or U10754 (N_10754,N_8574,N_9153);
nor U10755 (N_10755,N_9049,N_9219);
and U10756 (N_10756,N_9098,N_9000);
xor U10757 (N_10757,N_9483,N_9176);
and U10758 (N_10758,N_9183,N_8421);
and U10759 (N_10759,N_9133,N_9190);
and U10760 (N_10760,N_8913,N_9533);
xnor U10761 (N_10761,N_9366,N_9155);
nand U10762 (N_10762,N_8511,N_9228);
xor U10763 (N_10763,N_8489,N_8693);
or U10764 (N_10764,N_9263,N_8916);
xor U10765 (N_10765,N_8757,N_9122);
and U10766 (N_10766,N_9079,N_9341);
nor U10767 (N_10767,N_8973,N_9433);
xor U10768 (N_10768,N_8938,N_8724);
and U10769 (N_10769,N_9433,N_8902);
nand U10770 (N_10770,N_8677,N_8580);
xor U10771 (N_10771,N_9392,N_9399);
and U10772 (N_10772,N_9311,N_9571);
or U10773 (N_10773,N_9515,N_9057);
or U10774 (N_10774,N_9233,N_8489);
and U10775 (N_10775,N_9124,N_9300);
and U10776 (N_10776,N_9519,N_8616);
and U10777 (N_10777,N_8978,N_8502);
or U10778 (N_10778,N_9057,N_8643);
nor U10779 (N_10779,N_8865,N_9156);
xnor U10780 (N_10780,N_9052,N_8780);
and U10781 (N_10781,N_8411,N_8869);
xor U10782 (N_10782,N_9274,N_8580);
nand U10783 (N_10783,N_8507,N_9392);
xnor U10784 (N_10784,N_9235,N_8633);
nor U10785 (N_10785,N_8814,N_8678);
xnor U10786 (N_10786,N_8928,N_8805);
or U10787 (N_10787,N_8909,N_9248);
or U10788 (N_10788,N_8621,N_8422);
nand U10789 (N_10789,N_8535,N_8602);
and U10790 (N_10790,N_8941,N_8696);
or U10791 (N_10791,N_9222,N_9197);
and U10792 (N_10792,N_9063,N_9259);
or U10793 (N_10793,N_9499,N_8671);
or U10794 (N_10794,N_8867,N_8744);
xor U10795 (N_10795,N_9128,N_9359);
xnor U10796 (N_10796,N_9120,N_8572);
nand U10797 (N_10797,N_9231,N_9531);
or U10798 (N_10798,N_8631,N_8904);
nor U10799 (N_10799,N_8504,N_8849);
nand U10800 (N_10800,N_10359,N_9675);
nor U10801 (N_10801,N_9982,N_10505);
xnor U10802 (N_10802,N_10602,N_9799);
or U10803 (N_10803,N_10064,N_10315);
and U10804 (N_10804,N_9646,N_10186);
and U10805 (N_10805,N_9860,N_10516);
or U10806 (N_10806,N_10278,N_9838);
or U10807 (N_10807,N_10338,N_9644);
and U10808 (N_10808,N_10491,N_9876);
nand U10809 (N_10809,N_10349,N_9851);
or U10810 (N_10810,N_10449,N_10343);
nor U10811 (N_10811,N_9667,N_10564);
nor U10812 (N_10812,N_10334,N_10222);
xnor U10813 (N_10813,N_9928,N_10198);
and U10814 (N_10814,N_10237,N_9871);
or U10815 (N_10815,N_10748,N_9966);
and U10816 (N_10816,N_9955,N_10425);
and U10817 (N_10817,N_10525,N_10378);
or U10818 (N_10818,N_10632,N_10655);
xor U10819 (N_10819,N_10296,N_9770);
nand U10820 (N_10820,N_10780,N_10298);
nand U10821 (N_10821,N_10101,N_9768);
and U10822 (N_10822,N_10046,N_9886);
and U10823 (N_10823,N_10570,N_10319);
nor U10824 (N_10824,N_10039,N_9922);
nor U10825 (N_10825,N_9919,N_9954);
and U10826 (N_10826,N_10071,N_9730);
xor U10827 (N_10827,N_10756,N_10308);
nand U10828 (N_10828,N_10687,N_9752);
nand U10829 (N_10829,N_10156,N_10003);
or U10830 (N_10830,N_9834,N_10216);
and U10831 (N_10831,N_9936,N_10595);
nor U10832 (N_10832,N_10673,N_10382);
xor U10833 (N_10833,N_10138,N_10023);
nand U10834 (N_10834,N_10504,N_9638);
nand U10835 (N_10835,N_10514,N_9962);
nand U10836 (N_10836,N_10262,N_10354);
nor U10837 (N_10837,N_10478,N_9617);
or U10838 (N_10838,N_9804,N_10696);
xor U10839 (N_10839,N_10123,N_9968);
nor U10840 (N_10840,N_10412,N_9779);
xor U10841 (N_10841,N_9633,N_10347);
and U10842 (N_10842,N_10768,N_10289);
nand U10843 (N_10843,N_9864,N_9995);
xor U10844 (N_10844,N_10455,N_10117);
xor U10845 (N_10845,N_10456,N_10323);
or U10846 (N_10846,N_9607,N_9979);
nor U10847 (N_10847,N_10465,N_10436);
xor U10848 (N_10848,N_10145,N_9980);
xnor U10849 (N_10849,N_10453,N_9746);
nand U10850 (N_10850,N_10727,N_10684);
nor U10851 (N_10851,N_10473,N_10481);
nor U10852 (N_10852,N_10579,N_9636);
xnor U10853 (N_10853,N_10657,N_10600);
nor U10854 (N_10854,N_10243,N_9819);
nor U10855 (N_10855,N_10059,N_9679);
or U10856 (N_10856,N_10509,N_10085);
xor U10857 (N_10857,N_10053,N_9830);
xnor U10858 (N_10858,N_10075,N_10394);
nand U10859 (N_10859,N_10598,N_10726);
xor U10860 (N_10860,N_10745,N_10521);
nand U10861 (N_10861,N_10331,N_10231);
nor U10862 (N_10862,N_9678,N_10164);
nand U10863 (N_10863,N_10189,N_9845);
and U10864 (N_10864,N_10385,N_9662);
and U10865 (N_10865,N_10631,N_10017);
nand U10866 (N_10866,N_10662,N_10383);
nand U10867 (N_10867,N_10345,N_10470);
xor U10868 (N_10868,N_9665,N_10639);
and U10869 (N_10869,N_10523,N_10251);
xor U10870 (N_10870,N_10114,N_10041);
nor U10871 (N_10871,N_10152,N_10765);
nor U10872 (N_10872,N_10543,N_10499);
or U10873 (N_10873,N_10444,N_9726);
and U10874 (N_10874,N_10125,N_10739);
nand U10875 (N_10875,N_10176,N_10445);
nor U10876 (N_10876,N_10008,N_9977);
and U10877 (N_10877,N_9642,N_10356);
nor U10878 (N_10878,N_9647,N_10688);
or U10879 (N_10879,N_9902,N_9693);
nand U10880 (N_10880,N_9885,N_10160);
nand U10881 (N_10881,N_10734,N_9737);
and U10882 (N_10882,N_10577,N_10741);
and U10883 (N_10883,N_10510,N_10795);
nand U10884 (N_10884,N_10573,N_9811);
nor U10885 (N_10885,N_10058,N_10287);
nor U10886 (N_10886,N_10077,N_10400);
nor U10887 (N_10887,N_10433,N_10680);
and U10888 (N_10888,N_9970,N_10312);
nor U10889 (N_10889,N_10421,N_9916);
and U10890 (N_10890,N_9854,N_10515);
xor U10891 (N_10891,N_10363,N_10616);
nor U10892 (N_10892,N_10207,N_9703);
nand U10893 (N_10893,N_10401,N_10781);
and U10894 (N_10894,N_10789,N_10544);
xor U10895 (N_10895,N_9862,N_10572);
nor U10896 (N_10896,N_10099,N_10622);
and U10897 (N_10897,N_10667,N_10295);
and U10898 (N_10898,N_10321,N_9622);
or U10899 (N_10899,N_10614,N_10280);
or U10900 (N_10900,N_10173,N_9740);
nand U10901 (N_10901,N_10178,N_9610);
and U10902 (N_10902,N_9612,N_10530);
or U10903 (N_10903,N_10537,N_10568);
nand U10904 (N_10904,N_10764,N_9631);
nand U10905 (N_10905,N_9824,N_10605);
xnor U10906 (N_10906,N_10633,N_9975);
and U10907 (N_10907,N_10462,N_10518);
xor U10908 (N_10908,N_10601,N_10049);
or U10909 (N_10909,N_10731,N_10273);
and U10910 (N_10910,N_9701,N_10105);
nor U10911 (N_10911,N_10206,N_10387);
nor U10912 (N_10912,N_10221,N_10332);
nand U10913 (N_10913,N_10498,N_10552);
nand U10914 (N_10914,N_9791,N_10672);
nand U10915 (N_10915,N_10325,N_10092);
or U10916 (N_10916,N_9608,N_9805);
nor U10917 (N_10917,N_9844,N_10670);
nor U10918 (N_10918,N_10018,N_10150);
and U10919 (N_10919,N_10715,N_10259);
or U10920 (N_10920,N_10469,N_10047);
nand U10921 (N_10921,N_9933,N_10292);
or U10922 (N_10922,N_10584,N_9993);
or U10923 (N_10923,N_10426,N_10214);
nor U10924 (N_10924,N_9640,N_9648);
nand U10925 (N_10925,N_9857,N_10578);
xor U10926 (N_10926,N_10419,N_10035);
xor U10927 (N_10927,N_10226,N_10057);
nand U10928 (N_10928,N_9895,N_10265);
and U10929 (N_10929,N_9974,N_10586);
or U10930 (N_10930,N_9738,N_10648);
nor U10931 (N_10931,N_9664,N_10559);
or U10932 (N_10932,N_10428,N_10037);
xnor U10933 (N_10933,N_9956,N_10241);
xor U10934 (N_10934,N_9797,N_9786);
or U10935 (N_10935,N_10255,N_10420);
or U10936 (N_10936,N_9651,N_10617);
and U10937 (N_10937,N_10061,N_10458);
xnor U10938 (N_10938,N_9809,N_10116);
and U10939 (N_10939,N_9852,N_10095);
nor U10940 (N_10940,N_10471,N_10540);
or U10941 (N_10941,N_10233,N_9987);
nor U10942 (N_10942,N_10679,N_10341);
nor U10943 (N_10943,N_9963,N_10678);
and U10944 (N_10944,N_10148,N_10202);
nand U10945 (N_10945,N_9878,N_10333);
and U10946 (N_10946,N_9621,N_9721);
nor U10947 (N_10947,N_10107,N_9985);
or U10948 (N_10948,N_10266,N_9745);
and U10949 (N_10949,N_10740,N_10532);
and U10950 (N_10950,N_10682,N_9652);
and U10951 (N_10951,N_10188,N_10466);
xnor U10952 (N_10952,N_10630,N_9714);
nor U10953 (N_10953,N_10327,N_10585);
nor U10954 (N_10954,N_9867,N_9643);
nand U10955 (N_10955,N_10253,N_10100);
nand U10956 (N_10956,N_9835,N_9842);
nor U10957 (N_10957,N_9718,N_10264);
nand U10958 (N_10958,N_10318,N_9937);
nand U10959 (N_10959,N_10056,N_10257);
xnor U10960 (N_10960,N_9771,N_9912);
xor U10961 (N_10961,N_10369,N_10157);
and U10962 (N_10962,N_9778,N_10172);
xnor U10963 (N_10963,N_9847,N_9994);
nor U10964 (N_10964,N_10763,N_10162);
nor U10965 (N_10965,N_10083,N_10380);
or U10966 (N_10966,N_10081,N_10060);
and U10967 (N_10967,N_10699,N_10032);
and U10968 (N_10968,N_10635,N_9958);
nor U10969 (N_10969,N_10494,N_9641);
nand U10970 (N_10970,N_10155,N_10080);
or U10971 (N_10971,N_9817,N_10279);
nor U10972 (N_10972,N_9940,N_10574);
nand U10973 (N_10973,N_10301,N_10045);
and U10974 (N_10974,N_10762,N_9986);
nor U10975 (N_10975,N_9793,N_10171);
nand U10976 (N_10976,N_9783,N_10649);
and U10977 (N_10977,N_10429,N_10555);
or U10978 (N_10978,N_10604,N_10766);
xor U10979 (N_10979,N_10652,N_10424);
nor U10980 (N_10980,N_10608,N_10040);
or U10981 (N_10981,N_9932,N_10698);
nand U10982 (N_10982,N_9984,N_10399);
xor U10983 (N_10983,N_10344,N_10431);
xnor U10984 (N_10984,N_10275,N_10381);
or U10985 (N_10985,N_10026,N_10261);
nand U10986 (N_10986,N_10239,N_10755);
nand U10987 (N_10987,N_10238,N_10210);
nor U10988 (N_10988,N_10541,N_9736);
xor U10989 (N_10989,N_10036,N_9866);
or U10990 (N_10990,N_10685,N_10592);
or U10991 (N_10991,N_10025,N_10771);
or U10992 (N_10992,N_9808,N_10668);
and U10993 (N_10993,N_9654,N_9766);
nand U10994 (N_10994,N_10645,N_10563);
xnor U10995 (N_10995,N_10054,N_10192);
and U10996 (N_10996,N_10084,N_10713);
or U10997 (N_10997,N_10127,N_10693);
and U10998 (N_10998,N_9753,N_9723);
nor U10999 (N_10999,N_10671,N_9719);
xnor U11000 (N_11000,N_10194,N_10752);
and U11001 (N_11001,N_10597,N_10001);
and U11002 (N_11002,N_10277,N_10619);
nand U11003 (N_11003,N_10430,N_9749);
xnor U11004 (N_11004,N_10413,N_9700);
or U11005 (N_11005,N_10069,N_10550);
xor U11006 (N_11006,N_10451,N_9605);
nor U11007 (N_11007,N_9704,N_10720);
xor U11008 (N_11008,N_9780,N_10733);
nor U11009 (N_11009,N_10070,N_9861);
nand U11010 (N_11010,N_9814,N_9687);
xnor U11011 (N_11011,N_9903,N_10594);
nand U11012 (N_11012,N_10212,N_10772);
and U11013 (N_11013,N_10282,N_10722);
nor U11014 (N_11014,N_10367,N_10450);
nor U11015 (N_11015,N_10031,N_9840);
and U11016 (N_11016,N_9717,N_10408);
nand U11017 (N_11017,N_10492,N_10270);
xor U11018 (N_11018,N_10423,N_10154);
and U11019 (N_11019,N_10208,N_10588);
nand U11020 (N_11020,N_9725,N_9614);
or U11021 (N_11021,N_9875,N_9948);
xor U11022 (N_11022,N_9628,N_10417);
nor U11023 (N_11023,N_10744,N_10386);
nor U11024 (N_11024,N_10683,N_10476);
xnor U11025 (N_11025,N_10621,N_10180);
nand U11026 (N_11026,N_10131,N_9992);
or U11027 (N_11027,N_9934,N_10236);
or U11028 (N_11028,N_10593,N_10618);
nor U11029 (N_11029,N_9790,N_10747);
and U11030 (N_11030,N_10091,N_10474);
and U11031 (N_11031,N_9711,N_10034);
nor U11032 (N_11032,N_9829,N_10728);
nor U11033 (N_11033,N_9873,N_9757);
nor U11034 (N_11034,N_10260,N_9818);
xnor U11035 (N_11035,N_9708,N_10664);
or U11036 (N_11036,N_10751,N_9894);
and U11037 (N_11037,N_10551,N_10109);
and U11038 (N_11038,N_10336,N_10407);
or U11039 (N_11039,N_10288,N_10457);
nand U11040 (N_11040,N_9868,N_10256);
nor U11041 (N_11041,N_9619,N_10403);
or U11042 (N_11042,N_9705,N_10377);
xor U11043 (N_11043,N_9653,N_10330);
xnor U11044 (N_11044,N_9688,N_9685);
xnor U11045 (N_11045,N_9748,N_9759);
or U11046 (N_11046,N_10446,N_10524);
and U11047 (N_11047,N_10447,N_10785);
or U11048 (N_11048,N_9776,N_10258);
xnor U11049 (N_11049,N_9945,N_10501);
nor U11050 (N_11050,N_10783,N_10132);
nor U11051 (N_11051,N_9976,N_10374);
xor U11052 (N_11052,N_9800,N_10596);
nor U11053 (N_11053,N_10538,N_10010);
or U11054 (N_11054,N_9777,N_9645);
xor U11055 (N_11055,N_10159,N_10326);
and U11056 (N_11056,N_10181,N_10730);
nand U11057 (N_11057,N_10676,N_10545);
nor U11058 (N_11058,N_10486,N_9931);
and U11059 (N_11059,N_9858,N_10729);
nor U11060 (N_11060,N_9944,N_10587);
and U11061 (N_11061,N_9870,N_10314);
and U11062 (N_11062,N_10371,N_9850);
nor U11063 (N_11063,N_10389,N_10044);
nor U11064 (N_11064,N_10220,N_10767);
or U11065 (N_11065,N_10620,N_10792);
xor U11066 (N_11066,N_10463,N_10303);
nand U11067 (N_11067,N_10583,N_10439);
xnor U11068 (N_11068,N_10370,N_9695);
or U11069 (N_11069,N_9965,N_9889);
xnor U11070 (N_11070,N_9670,N_9739);
xnor U11071 (N_11071,N_9991,N_10115);
or U11072 (N_11072,N_9901,N_10711);
and U11073 (N_11073,N_10087,N_9689);
and U11074 (N_11074,N_10137,N_10638);
or U11075 (N_11075,N_10144,N_10348);
nand U11076 (N_11076,N_10777,N_9702);
xor U11077 (N_11077,N_10310,N_9639);
xor U11078 (N_11078,N_10111,N_10364);
or U11079 (N_11079,N_10717,N_10719);
xnor U11080 (N_11080,N_10788,N_9884);
nor U11081 (N_11081,N_10660,N_9796);
or U11082 (N_11082,N_9660,N_9942);
xor U11083 (N_11083,N_10472,N_9802);
or U11084 (N_11084,N_9773,N_10067);
nand U11085 (N_11085,N_10324,N_10461);
and U11086 (N_11086,N_9816,N_10448);
xor U11087 (N_11087,N_10272,N_9935);
nand U11088 (N_11088,N_10590,N_10391);
nor U11089 (N_11089,N_10218,N_10089);
nand U11090 (N_11090,N_9964,N_10654);
nor U11091 (N_11091,N_10666,N_10774);
nand U11092 (N_11092,N_10441,N_9686);
xnor U11093 (N_11093,N_10414,N_10760);
xnor U11094 (N_11094,N_10651,N_10142);
xnor U11095 (N_11095,N_9900,N_10168);
xor U11096 (N_11096,N_9656,N_10692);
and U11097 (N_11097,N_10368,N_10468);
xnor U11098 (N_11098,N_10710,N_9661);
nor U11099 (N_11099,N_10066,N_9904);
xor U11100 (N_11100,N_9715,N_9795);
nor U11101 (N_11101,N_10005,N_10533);
or U11102 (N_11102,N_9951,N_9839);
or U11103 (N_11103,N_10395,N_10042);
xor U11104 (N_11104,N_10422,N_10011);
or U11105 (N_11105,N_9673,N_10508);
and U11106 (N_11106,N_9697,N_9668);
nor U11107 (N_11107,N_10228,N_10103);
or U11108 (N_11108,N_10576,N_9843);
nor U11109 (N_11109,N_10475,N_10637);
xor U11110 (N_11110,N_10535,N_10675);
or U11111 (N_11111,N_10182,N_10106);
and U11112 (N_11112,N_10196,N_10285);
xor U11113 (N_11113,N_10124,N_10379);
and U11114 (N_11114,N_10249,N_10689);
nor U11115 (N_11115,N_10562,N_10108);
and U11116 (N_11116,N_9650,N_9957);
and U11117 (N_11117,N_9859,N_9890);
or U11118 (N_11118,N_10793,N_10665);
and U11119 (N_11119,N_10104,N_10140);
and U11120 (N_11120,N_9671,N_9659);
nor U11121 (N_11121,N_10133,N_10786);
nor U11122 (N_11122,N_9720,N_10418);
or U11123 (N_11123,N_10244,N_9727);
or U11124 (N_11124,N_10022,N_10187);
nor U11125 (N_11125,N_9891,N_10139);
nor U11126 (N_11126,N_10337,N_10043);
or U11127 (N_11127,N_9728,N_10183);
and U11128 (N_11128,N_9927,N_10358);
nor U11129 (N_11129,N_10293,N_9606);
xor U11130 (N_11130,N_9911,N_9680);
nand U11131 (N_11131,N_10234,N_9882);
xnor U11132 (N_11132,N_10388,N_9831);
nand U11133 (N_11133,N_10549,N_9774);
nand U11134 (N_11134,N_10758,N_9696);
or U11135 (N_11135,N_10063,N_9674);
and U11136 (N_11136,N_10128,N_9832);
nand U11137 (N_11137,N_10141,N_10704);
nor U11138 (N_11138,N_10415,N_10750);
nor U11139 (N_11139,N_9602,N_10406);
nand U11140 (N_11140,N_10749,N_10179);
xor U11141 (N_11141,N_10283,N_9812);
nor U11142 (N_11142,N_10575,N_10434);
or U11143 (N_11143,N_10607,N_9909);
and U11144 (N_11144,N_9960,N_10612);
nor U11145 (N_11145,N_9676,N_9732);
and U11146 (N_11146,N_10694,N_10489);
or U11147 (N_11147,N_9691,N_10610);
and U11148 (N_11148,N_9604,N_9813);
nand U11149 (N_11149,N_10790,N_10791);
nor U11150 (N_11150,N_9907,N_10294);
xor U11151 (N_11151,N_10490,N_10480);
nand U11152 (N_11152,N_10086,N_10297);
and U11153 (N_11153,N_10522,N_10496);
and U11154 (N_11154,N_10223,N_10440);
and U11155 (N_11155,N_10746,N_10134);
xor U11156 (N_11156,N_10517,N_9649);
and U11157 (N_11157,N_9755,N_10452);
nand U11158 (N_11158,N_10778,N_9655);
nor U11159 (N_11159,N_9879,N_10485);
and U11160 (N_11160,N_9751,N_9988);
or U11161 (N_11161,N_9952,N_10511);
nor U11162 (N_11162,N_10000,N_10165);
and U11163 (N_11163,N_10467,N_10002);
nor U11164 (N_11164,N_10073,N_10153);
nand U11165 (N_11165,N_10798,N_10690);
nand U11166 (N_11166,N_10360,N_10629);
and U11167 (N_11167,N_10613,N_10569);
xor U11168 (N_11168,N_10009,N_10703);
nand U11169 (N_11169,N_10546,N_10015);
nor U11170 (N_11170,N_10493,N_10691);
or U11171 (N_11171,N_9893,N_9863);
nor U11172 (N_11172,N_9999,N_10784);
nor U11173 (N_11173,N_10120,N_10442);
or U11174 (N_11174,N_9713,N_9915);
nand U11175 (N_11175,N_10136,N_9716);
nor U11176 (N_11176,N_10742,N_10102);
and U11177 (N_11177,N_9792,N_10735);
xnor U11178 (N_11178,N_9921,N_9669);
nor U11179 (N_11179,N_10506,N_10163);
or U11180 (N_11180,N_10623,N_9710);
nor U11181 (N_11181,N_9837,N_9760);
or U11182 (N_11182,N_10365,N_10030);
and U11183 (N_11183,N_10707,N_10700);
nor U11184 (N_11184,N_10513,N_10012);
nor U11185 (N_11185,N_9692,N_10460);
nand U11186 (N_11186,N_10024,N_10674);
and U11187 (N_11187,N_10254,N_10628);
nand U11188 (N_11188,N_9856,N_9972);
xor U11189 (N_11189,N_10299,N_10566);
xor U11190 (N_11190,N_10640,N_9694);
nand U11191 (N_11191,N_10737,N_9750);
nor U11192 (N_11192,N_10203,N_9618);
and U11193 (N_11193,N_10794,N_10232);
xnor U11194 (N_11194,N_9765,N_10464);
nand U11195 (N_11195,N_10659,N_10409);
xnor U11196 (N_11196,N_10329,N_10190);
and U11197 (N_11197,N_10484,N_10240);
nor U11198 (N_11198,N_10761,N_10384);
xnor U11199 (N_11199,N_10093,N_10328);
xor U11200 (N_11200,N_9990,N_10567);
or U11201 (N_11201,N_9941,N_10557);
nand U11202 (N_11202,N_10316,N_10055);
nor U11203 (N_11203,N_9848,N_10641);
nor U11204 (N_11204,N_10705,N_10305);
xor U11205 (N_11205,N_10065,N_9918);
nand U11206 (N_11206,N_10021,N_10129);
nor U11207 (N_11207,N_10677,N_10642);
nand U11208 (N_11208,N_9996,N_10571);
nor U11209 (N_11209,N_10714,N_9807);
xnor U11210 (N_11210,N_9741,N_10197);
nand U11211 (N_11211,N_9888,N_10224);
xnor U11212 (N_11212,N_10560,N_9729);
nor U11213 (N_11213,N_9761,N_9789);
or U11214 (N_11214,N_9634,N_9825);
xnor U11215 (N_11215,N_10161,N_10306);
nor U11216 (N_11216,N_9706,N_10591);
nor U11217 (N_11217,N_10779,N_10355);
and U11218 (N_11218,N_9923,N_10118);
and U11219 (N_11219,N_9758,N_10392);
xnor U11220 (N_11220,N_9600,N_9623);
or U11221 (N_11221,N_9828,N_10110);
xnor U11222 (N_11222,N_10527,N_10757);
nand U11223 (N_11223,N_10130,N_10169);
xnor U11224 (N_11224,N_10004,N_9763);
nor U11225 (N_11225,N_10151,N_9784);
or U11226 (N_11226,N_9754,N_10663);
nand U11227 (N_11227,N_9821,N_10146);
xor U11228 (N_11228,N_10437,N_9764);
xnor U11229 (N_11229,N_9981,N_10410);
xnor U11230 (N_11230,N_9767,N_9946);
nor U11231 (N_11231,N_10695,N_9961);
nand U11232 (N_11232,N_10443,N_9637);
or U11233 (N_11233,N_10398,N_10033);
or U11234 (N_11234,N_10732,N_9883);
nand U11235 (N_11235,N_9787,N_9910);
nor U11236 (N_11236,N_9827,N_9905);
nand U11237 (N_11237,N_9616,N_9969);
xnor U11238 (N_11238,N_10170,N_10606);
and U11239 (N_11239,N_9798,N_10211);
or U11240 (N_11240,N_10479,N_9925);
and U11241 (N_11241,N_10339,N_10770);
and U11242 (N_11242,N_9971,N_9892);
nor U11243 (N_11243,N_10227,N_10488);
and U11244 (N_11244,N_10028,N_9846);
xnor U11245 (N_11245,N_10534,N_10542);
and U11246 (N_11246,N_10121,N_10497);
nand U11247 (N_11247,N_10376,N_9724);
xor U11248 (N_11248,N_10661,N_10068);
nor U11249 (N_11249,N_10185,N_9899);
and U11250 (N_11250,N_10454,N_10507);
nand U11251 (N_11251,N_9872,N_9989);
nor U11252 (N_11252,N_10405,N_10304);
nor U11253 (N_11253,N_10404,N_10581);
xor U11254 (N_11254,N_10706,N_10529);
nand U11255 (N_11255,N_10502,N_10119);
xnor U11256 (N_11256,N_10352,N_10643);
nand U11257 (N_11257,N_9983,N_9603);
nand U11258 (N_11258,N_9836,N_10204);
nand U11259 (N_11259,N_9810,N_10038);
or U11260 (N_11260,N_10290,N_10708);
and U11261 (N_11261,N_10647,N_10754);
nand U11262 (N_11262,N_10094,N_10701);
nand U11263 (N_11263,N_10556,N_10531);
or U11264 (N_11264,N_9943,N_10200);
nand U11265 (N_11265,N_10702,N_9920);
nor U11266 (N_11266,N_9742,N_10561);
nand U11267 (N_11267,N_9806,N_10311);
nor U11268 (N_11268,N_10219,N_10235);
or U11269 (N_11269,N_10723,N_9896);
or U11270 (N_11270,N_10247,N_10014);
nor U11271 (N_11271,N_9906,N_9924);
xor U11272 (N_11272,N_9672,N_9914);
or U11273 (N_11273,N_10143,N_10477);
xor U11274 (N_11274,N_10252,N_10268);
and U11275 (N_11275,N_9801,N_10340);
nor U11276 (N_11276,N_9629,N_10191);
xor U11277 (N_11277,N_9908,N_10548);
nor U11278 (N_11278,N_10495,N_9769);
nand U11279 (N_11279,N_10193,N_10427);
and U11280 (N_11280,N_10175,N_10390);
nand U11281 (N_11281,N_10263,N_10113);
and U11282 (N_11282,N_10149,N_10624);
or U11283 (N_11283,N_10773,N_10438);
nor U11284 (N_11284,N_9627,N_10526);
nand U11285 (N_11285,N_10373,N_10709);
and U11286 (N_11286,N_10353,N_9815);
or U11287 (N_11287,N_10565,N_10372);
and U11288 (N_11288,N_10229,N_10603);
and U11289 (N_11289,N_10097,N_9998);
nand U11290 (N_11290,N_9917,N_9869);
nor U11291 (N_11291,N_10636,N_10724);
and U11292 (N_11292,N_9658,N_10242);
and U11293 (N_11293,N_10271,N_10459);
nor U11294 (N_11294,N_10027,N_9626);
xnor U11295 (N_11295,N_10656,N_9826);
nand U11296 (N_11296,N_9775,N_9849);
xnor U11297 (N_11297,N_10634,N_9820);
nor U11298 (N_11298,N_9913,N_10286);
and U11299 (N_11299,N_9632,N_10167);
nor U11300 (N_11300,N_10051,N_10366);
xor U11301 (N_11301,N_9735,N_9684);
or U11302 (N_11302,N_9743,N_10013);
xor U11303 (N_11303,N_10209,N_9953);
nand U11304 (N_11304,N_9877,N_10402);
xor U11305 (N_11305,N_10135,N_9756);
or U11306 (N_11306,N_10500,N_10697);
and U11307 (N_11307,N_10201,N_10393);
or U11308 (N_11308,N_10317,N_10082);
nor U11309 (N_11309,N_10487,N_10653);
or U11310 (N_11310,N_10250,N_10776);
or U11311 (N_11311,N_10300,N_10020);
nor U11312 (N_11312,N_10519,N_10029);
and U11313 (N_11313,N_10554,N_10246);
and U11314 (N_11314,N_9609,N_10599);
and U11315 (N_11315,N_10079,N_10313);
xnor U11316 (N_11316,N_10245,N_9666);
nand U11317 (N_11317,N_10320,N_10553);
or U11318 (N_11318,N_10225,N_9950);
nor U11319 (N_11319,N_10007,N_10177);
xnor U11320 (N_11320,N_10611,N_10205);
or U11321 (N_11321,N_10432,N_10625);
or U11322 (N_11322,N_10126,N_9803);
nor U11323 (N_11323,N_9707,N_10743);
or U11324 (N_11324,N_9625,N_10716);
nand U11325 (N_11325,N_9762,N_9897);
nor U11326 (N_11326,N_9613,N_10088);
nor U11327 (N_11327,N_9874,N_10052);
xnor U11328 (N_11328,N_10302,N_10650);
and U11329 (N_11329,N_9698,N_10346);
or U11330 (N_11330,N_9772,N_10158);
and U11331 (N_11331,N_9731,N_10520);
nand U11332 (N_11332,N_10686,N_10248);
nor U11333 (N_11333,N_10309,N_9938);
nand U11334 (N_11334,N_10284,N_9709);
nor U11335 (N_11335,N_10375,N_9929);
and U11336 (N_11336,N_10753,N_10725);
xor U11337 (N_11337,N_10626,N_9733);
nor U11338 (N_11338,N_10019,N_9611);
xnor U11339 (N_11339,N_10195,N_10062);
nand U11340 (N_11340,N_9690,N_10213);
nand U11341 (N_11341,N_9959,N_10539);
and U11342 (N_11342,N_10718,N_10646);
xor U11343 (N_11343,N_10357,N_9785);
nor U11344 (N_11344,N_9682,N_9939);
nand U11345 (N_11345,N_9782,N_9722);
or U11346 (N_11346,N_9833,N_10799);
nor U11347 (N_11347,N_9887,N_10721);
nor U11348 (N_11348,N_9699,N_10078);
and U11349 (N_11349,N_10609,N_10615);
xor U11350 (N_11350,N_10217,N_9788);
or U11351 (N_11351,N_10681,N_9881);
nand U11352 (N_11352,N_10589,N_10281);
xnor U11353 (N_11353,N_10361,N_9677);
nand U11354 (N_11354,N_9681,N_9926);
nor U11355 (N_11355,N_10076,N_10396);
and U11356 (N_11356,N_10072,N_10291);
nor U11357 (N_11357,N_9744,N_10351);
nand U11358 (N_11358,N_10335,N_10658);
or U11359 (N_11359,N_10016,N_9930);
and U11360 (N_11360,N_10547,N_10098);
and U11361 (N_11361,N_10644,N_10512);
nand U11362 (N_11362,N_10342,N_10147);
xnor U11363 (N_11363,N_10416,N_9601);
nand U11364 (N_11364,N_9657,N_9973);
or U11365 (N_11365,N_10269,N_10759);
xor U11366 (N_11366,N_10411,N_9615);
xor U11367 (N_11367,N_10276,N_10483);
xor U11368 (N_11368,N_9624,N_10582);
nand U11369 (N_11369,N_9898,N_10267);
or U11370 (N_11370,N_9880,N_10797);
xnor U11371 (N_11371,N_9734,N_10712);
and U11372 (N_11372,N_9747,N_10230);
xor U11373 (N_11373,N_10627,N_9967);
xor U11374 (N_11374,N_10184,N_10048);
nand U11375 (N_11375,N_10397,N_9949);
xor U11376 (N_11376,N_9865,N_9663);
xor U11377 (N_11377,N_10787,N_10050);
nand U11378 (N_11378,N_10580,N_9620);
or U11379 (N_11379,N_9997,N_10350);
xnor U11380 (N_11380,N_10174,N_9978);
nor U11381 (N_11381,N_10112,N_9841);
nor U11382 (N_11382,N_10274,N_10558);
nor U11383 (N_11383,N_10166,N_10074);
xnor U11384 (N_11384,N_9823,N_9683);
nor U11385 (N_11385,N_10122,N_9853);
nand U11386 (N_11386,N_9822,N_10006);
nand U11387 (N_11387,N_10435,N_10736);
nor U11388 (N_11388,N_9781,N_10738);
or U11389 (N_11389,N_10199,N_9947);
and U11390 (N_11390,N_10090,N_10536);
or U11391 (N_11391,N_10528,N_10796);
xor U11392 (N_11392,N_10775,N_10482);
xnor U11393 (N_11393,N_10769,N_9794);
or U11394 (N_11394,N_10096,N_10362);
xor U11395 (N_11395,N_10503,N_10782);
or U11396 (N_11396,N_10307,N_9855);
or U11397 (N_11397,N_9630,N_9635);
and U11398 (N_11398,N_9712,N_10215);
nand U11399 (N_11399,N_10322,N_10669);
nor U11400 (N_11400,N_9843,N_9763);
xnor U11401 (N_11401,N_10185,N_10108);
nand U11402 (N_11402,N_10366,N_10399);
nand U11403 (N_11403,N_10532,N_10698);
or U11404 (N_11404,N_10366,N_9891);
and U11405 (N_11405,N_10361,N_10196);
nand U11406 (N_11406,N_10432,N_10469);
or U11407 (N_11407,N_10108,N_10227);
nor U11408 (N_11408,N_10566,N_10360);
nor U11409 (N_11409,N_10672,N_10042);
xor U11410 (N_11410,N_10645,N_9999);
xnor U11411 (N_11411,N_9894,N_10253);
nand U11412 (N_11412,N_9958,N_9880);
or U11413 (N_11413,N_10779,N_9703);
nor U11414 (N_11414,N_10353,N_10463);
or U11415 (N_11415,N_10623,N_9678);
and U11416 (N_11416,N_10702,N_10716);
xnor U11417 (N_11417,N_10446,N_9821);
and U11418 (N_11418,N_9807,N_9901);
nand U11419 (N_11419,N_9726,N_9807);
nand U11420 (N_11420,N_10502,N_10278);
or U11421 (N_11421,N_10250,N_10385);
or U11422 (N_11422,N_9652,N_9887);
and U11423 (N_11423,N_10644,N_10613);
nand U11424 (N_11424,N_10506,N_10236);
or U11425 (N_11425,N_9913,N_9686);
nand U11426 (N_11426,N_9972,N_10044);
xor U11427 (N_11427,N_10471,N_10392);
nor U11428 (N_11428,N_9949,N_9845);
nor U11429 (N_11429,N_9685,N_10093);
or U11430 (N_11430,N_9957,N_10159);
xor U11431 (N_11431,N_10606,N_10107);
nand U11432 (N_11432,N_9855,N_10603);
and U11433 (N_11433,N_10270,N_10160);
and U11434 (N_11434,N_10104,N_9827);
xor U11435 (N_11435,N_10158,N_9820);
and U11436 (N_11436,N_10648,N_10737);
xor U11437 (N_11437,N_10797,N_10211);
xor U11438 (N_11438,N_10582,N_9616);
nand U11439 (N_11439,N_10581,N_9786);
nand U11440 (N_11440,N_10118,N_9981);
nor U11441 (N_11441,N_9810,N_9962);
xnor U11442 (N_11442,N_10643,N_10443);
nor U11443 (N_11443,N_9707,N_10428);
nor U11444 (N_11444,N_9777,N_10746);
and U11445 (N_11445,N_10159,N_10581);
xor U11446 (N_11446,N_10314,N_10132);
nor U11447 (N_11447,N_9923,N_10488);
and U11448 (N_11448,N_10012,N_9791);
nor U11449 (N_11449,N_10426,N_10570);
nand U11450 (N_11450,N_10232,N_10072);
nand U11451 (N_11451,N_9883,N_10434);
or U11452 (N_11452,N_10279,N_9865);
nor U11453 (N_11453,N_9709,N_10143);
nor U11454 (N_11454,N_10009,N_9641);
and U11455 (N_11455,N_10037,N_9965);
nor U11456 (N_11456,N_10040,N_10523);
or U11457 (N_11457,N_10327,N_10104);
nand U11458 (N_11458,N_10560,N_10026);
nand U11459 (N_11459,N_10065,N_9622);
nor U11460 (N_11460,N_10408,N_9908);
and U11461 (N_11461,N_10501,N_9921);
or U11462 (N_11462,N_10701,N_10099);
xor U11463 (N_11463,N_10791,N_10554);
nand U11464 (N_11464,N_10678,N_10280);
nand U11465 (N_11465,N_10132,N_10073);
and U11466 (N_11466,N_9874,N_9809);
or U11467 (N_11467,N_9684,N_9729);
or U11468 (N_11468,N_9935,N_10552);
or U11469 (N_11469,N_10370,N_10391);
xnor U11470 (N_11470,N_10349,N_10269);
nand U11471 (N_11471,N_9975,N_9721);
and U11472 (N_11472,N_10667,N_10414);
or U11473 (N_11473,N_10329,N_9767);
nor U11474 (N_11474,N_9880,N_10282);
nor U11475 (N_11475,N_10342,N_10571);
nand U11476 (N_11476,N_10355,N_9608);
xnor U11477 (N_11477,N_10761,N_10232);
nand U11478 (N_11478,N_10195,N_10297);
or U11479 (N_11479,N_10654,N_9822);
or U11480 (N_11480,N_9844,N_9758);
xnor U11481 (N_11481,N_10266,N_10699);
nand U11482 (N_11482,N_10006,N_10540);
nor U11483 (N_11483,N_9634,N_9987);
or U11484 (N_11484,N_10144,N_9898);
and U11485 (N_11485,N_9856,N_10411);
and U11486 (N_11486,N_10410,N_10082);
nand U11487 (N_11487,N_10782,N_9665);
and U11488 (N_11488,N_10568,N_9750);
nand U11489 (N_11489,N_10404,N_9723);
xor U11490 (N_11490,N_10639,N_9758);
nand U11491 (N_11491,N_10223,N_9858);
nand U11492 (N_11492,N_9812,N_10036);
xnor U11493 (N_11493,N_9938,N_10745);
and U11494 (N_11494,N_10641,N_9747);
xor U11495 (N_11495,N_10120,N_10108);
and U11496 (N_11496,N_10052,N_10697);
and U11497 (N_11497,N_10462,N_9967);
xnor U11498 (N_11498,N_10775,N_10401);
nand U11499 (N_11499,N_9693,N_10281);
nor U11500 (N_11500,N_10101,N_9774);
nand U11501 (N_11501,N_10569,N_10273);
nand U11502 (N_11502,N_9683,N_10626);
or U11503 (N_11503,N_10518,N_9788);
or U11504 (N_11504,N_10067,N_10707);
nor U11505 (N_11505,N_10647,N_10374);
or U11506 (N_11506,N_10460,N_10634);
and U11507 (N_11507,N_10177,N_10425);
or U11508 (N_11508,N_10468,N_10148);
nand U11509 (N_11509,N_10623,N_10520);
nor U11510 (N_11510,N_10717,N_10690);
or U11511 (N_11511,N_9622,N_10724);
nand U11512 (N_11512,N_10469,N_10712);
or U11513 (N_11513,N_10322,N_10760);
and U11514 (N_11514,N_10379,N_9968);
and U11515 (N_11515,N_10008,N_10406);
nand U11516 (N_11516,N_10160,N_10041);
xor U11517 (N_11517,N_10137,N_9820);
or U11518 (N_11518,N_10390,N_10413);
nand U11519 (N_11519,N_9920,N_9957);
nand U11520 (N_11520,N_10247,N_10236);
xor U11521 (N_11521,N_9868,N_10786);
nor U11522 (N_11522,N_10029,N_9670);
xnor U11523 (N_11523,N_10388,N_9961);
xnor U11524 (N_11524,N_10054,N_10464);
and U11525 (N_11525,N_9847,N_10450);
and U11526 (N_11526,N_10072,N_10754);
or U11527 (N_11527,N_9915,N_10050);
nand U11528 (N_11528,N_10272,N_10128);
xnor U11529 (N_11529,N_10672,N_9838);
xnor U11530 (N_11530,N_9685,N_9965);
nor U11531 (N_11531,N_10662,N_9685);
nand U11532 (N_11532,N_10235,N_10559);
or U11533 (N_11533,N_10382,N_10694);
xnor U11534 (N_11534,N_10035,N_9995);
xor U11535 (N_11535,N_10301,N_10185);
nand U11536 (N_11536,N_9790,N_10123);
and U11537 (N_11537,N_10559,N_9833);
and U11538 (N_11538,N_9860,N_9946);
xnor U11539 (N_11539,N_10470,N_10156);
and U11540 (N_11540,N_10365,N_9856);
and U11541 (N_11541,N_10301,N_10419);
nor U11542 (N_11542,N_10300,N_10070);
xor U11543 (N_11543,N_10637,N_10105);
or U11544 (N_11544,N_9705,N_10642);
or U11545 (N_11545,N_10178,N_10312);
or U11546 (N_11546,N_10100,N_10109);
nor U11547 (N_11547,N_10359,N_10286);
nor U11548 (N_11548,N_10568,N_10385);
or U11549 (N_11549,N_10456,N_10510);
nor U11550 (N_11550,N_9872,N_10624);
nand U11551 (N_11551,N_9764,N_10607);
and U11552 (N_11552,N_10215,N_9796);
nor U11553 (N_11553,N_10469,N_9907);
xnor U11554 (N_11554,N_9953,N_10449);
xnor U11555 (N_11555,N_10018,N_10281);
and U11556 (N_11556,N_10079,N_10661);
and U11557 (N_11557,N_10559,N_10345);
or U11558 (N_11558,N_10381,N_10694);
xnor U11559 (N_11559,N_10459,N_9714);
or U11560 (N_11560,N_9631,N_9902);
xnor U11561 (N_11561,N_9903,N_10088);
or U11562 (N_11562,N_10754,N_9887);
or U11563 (N_11563,N_9832,N_10213);
and U11564 (N_11564,N_10670,N_10164);
and U11565 (N_11565,N_9939,N_9600);
xor U11566 (N_11566,N_10499,N_10047);
and U11567 (N_11567,N_9923,N_10602);
or U11568 (N_11568,N_9873,N_9728);
xnor U11569 (N_11569,N_10714,N_9961);
or U11570 (N_11570,N_9662,N_10088);
nor U11571 (N_11571,N_10055,N_10079);
nand U11572 (N_11572,N_10022,N_10441);
nor U11573 (N_11573,N_9751,N_10578);
or U11574 (N_11574,N_10589,N_9707);
nand U11575 (N_11575,N_10385,N_10260);
nor U11576 (N_11576,N_10799,N_10592);
and U11577 (N_11577,N_9679,N_9753);
nor U11578 (N_11578,N_9616,N_10739);
and U11579 (N_11579,N_10728,N_10193);
and U11580 (N_11580,N_9746,N_10434);
nor U11581 (N_11581,N_9920,N_9893);
nor U11582 (N_11582,N_9607,N_10434);
and U11583 (N_11583,N_10362,N_10541);
nand U11584 (N_11584,N_9955,N_10111);
nand U11585 (N_11585,N_10043,N_9768);
nand U11586 (N_11586,N_10485,N_9813);
xnor U11587 (N_11587,N_9619,N_10443);
nor U11588 (N_11588,N_10665,N_10507);
and U11589 (N_11589,N_10435,N_9758);
and U11590 (N_11590,N_10550,N_10339);
or U11591 (N_11591,N_10493,N_10706);
or U11592 (N_11592,N_10727,N_10139);
nor U11593 (N_11593,N_9633,N_10318);
and U11594 (N_11594,N_10462,N_9819);
nor U11595 (N_11595,N_10701,N_10299);
nand U11596 (N_11596,N_10471,N_10272);
nand U11597 (N_11597,N_9953,N_9900);
xor U11598 (N_11598,N_10303,N_10594);
and U11599 (N_11599,N_10274,N_10164);
xor U11600 (N_11600,N_9755,N_9839);
nand U11601 (N_11601,N_9661,N_9935);
nand U11602 (N_11602,N_10026,N_10401);
or U11603 (N_11603,N_10641,N_10359);
nand U11604 (N_11604,N_10059,N_9938);
and U11605 (N_11605,N_10162,N_9999);
nand U11606 (N_11606,N_10666,N_10335);
nand U11607 (N_11607,N_10605,N_9634);
nand U11608 (N_11608,N_9671,N_10797);
nand U11609 (N_11609,N_10314,N_10467);
xnor U11610 (N_11610,N_10142,N_9660);
nor U11611 (N_11611,N_10248,N_9778);
and U11612 (N_11612,N_9607,N_9938);
xor U11613 (N_11613,N_10446,N_10290);
or U11614 (N_11614,N_9785,N_10069);
xor U11615 (N_11615,N_9643,N_9602);
xor U11616 (N_11616,N_9742,N_10154);
or U11617 (N_11617,N_9783,N_10601);
nor U11618 (N_11618,N_9950,N_10418);
or U11619 (N_11619,N_9786,N_10513);
nand U11620 (N_11620,N_10142,N_10679);
nor U11621 (N_11621,N_10019,N_9908);
xor U11622 (N_11622,N_9617,N_10342);
or U11623 (N_11623,N_10731,N_10142);
nand U11624 (N_11624,N_9636,N_9692);
xor U11625 (N_11625,N_9963,N_9895);
or U11626 (N_11626,N_10579,N_9996);
nand U11627 (N_11627,N_9819,N_10005);
nand U11628 (N_11628,N_9843,N_10199);
or U11629 (N_11629,N_9735,N_10589);
xnor U11630 (N_11630,N_9956,N_10752);
nor U11631 (N_11631,N_10375,N_10585);
and U11632 (N_11632,N_10112,N_10359);
and U11633 (N_11633,N_10037,N_10385);
and U11634 (N_11634,N_10663,N_10138);
or U11635 (N_11635,N_10657,N_10614);
or U11636 (N_11636,N_9824,N_10790);
nor U11637 (N_11637,N_9897,N_10223);
nand U11638 (N_11638,N_10104,N_10110);
xor U11639 (N_11639,N_10398,N_10704);
and U11640 (N_11640,N_10727,N_9665);
or U11641 (N_11641,N_10637,N_9958);
and U11642 (N_11642,N_10569,N_10486);
and U11643 (N_11643,N_9898,N_10782);
nand U11644 (N_11644,N_9801,N_10790);
nor U11645 (N_11645,N_10396,N_10328);
and U11646 (N_11646,N_9684,N_9867);
nor U11647 (N_11647,N_10767,N_10330);
nand U11648 (N_11648,N_10208,N_10619);
xor U11649 (N_11649,N_9951,N_9808);
or U11650 (N_11650,N_9640,N_9805);
or U11651 (N_11651,N_10016,N_10320);
nand U11652 (N_11652,N_9782,N_10569);
nor U11653 (N_11653,N_10161,N_10766);
and U11654 (N_11654,N_10357,N_10580);
xor U11655 (N_11655,N_10540,N_10259);
and U11656 (N_11656,N_9909,N_10700);
or U11657 (N_11657,N_9744,N_9919);
and U11658 (N_11658,N_10267,N_9600);
nand U11659 (N_11659,N_9626,N_9662);
and U11660 (N_11660,N_9761,N_10701);
nand U11661 (N_11661,N_10218,N_9807);
xor U11662 (N_11662,N_10371,N_10208);
nor U11663 (N_11663,N_10510,N_10284);
nand U11664 (N_11664,N_10755,N_10299);
or U11665 (N_11665,N_10597,N_10089);
xor U11666 (N_11666,N_10743,N_9794);
nand U11667 (N_11667,N_10653,N_10661);
and U11668 (N_11668,N_10171,N_10750);
nand U11669 (N_11669,N_10452,N_9920);
nand U11670 (N_11670,N_10221,N_10652);
nand U11671 (N_11671,N_10635,N_10013);
xnor U11672 (N_11672,N_10483,N_10753);
xnor U11673 (N_11673,N_10306,N_9923);
and U11674 (N_11674,N_10161,N_10171);
xnor U11675 (N_11675,N_9713,N_10071);
or U11676 (N_11676,N_10347,N_10064);
xnor U11677 (N_11677,N_10329,N_10772);
or U11678 (N_11678,N_10553,N_9909);
nor U11679 (N_11679,N_10641,N_10558);
nor U11680 (N_11680,N_9890,N_9794);
or U11681 (N_11681,N_10394,N_9928);
or U11682 (N_11682,N_10608,N_9744);
and U11683 (N_11683,N_9895,N_9998);
nand U11684 (N_11684,N_10062,N_10072);
nand U11685 (N_11685,N_9910,N_9827);
xnor U11686 (N_11686,N_10480,N_10688);
and U11687 (N_11687,N_9695,N_9650);
or U11688 (N_11688,N_10706,N_9999);
nand U11689 (N_11689,N_10104,N_9658);
nor U11690 (N_11690,N_10489,N_10663);
xnor U11691 (N_11691,N_9942,N_10586);
or U11692 (N_11692,N_10281,N_10297);
or U11693 (N_11693,N_9703,N_10028);
nor U11694 (N_11694,N_9752,N_9996);
and U11695 (N_11695,N_9939,N_10673);
or U11696 (N_11696,N_10764,N_10347);
xnor U11697 (N_11697,N_10343,N_9891);
nand U11698 (N_11698,N_10645,N_10045);
xnor U11699 (N_11699,N_9750,N_9700);
xor U11700 (N_11700,N_10778,N_10467);
or U11701 (N_11701,N_10665,N_9970);
nand U11702 (N_11702,N_10771,N_9620);
xnor U11703 (N_11703,N_10528,N_10081);
nand U11704 (N_11704,N_10276,N_10494);
nor U11705 (N_11705,N_10204,N_9987);
nor U11706 (N_11706,N_10420,N_10038);
xor U11707 (N_11707,N_9956,N_9704);
nor U11708 (N_11708,N_10305,N_9802);
xnor U11709 (N_11709,N_10363,N_10084);
and U11710 (N_11710,N_10781,N_10178);
or U11711 (N_11711,N_9685,N_9874);
xnor U11712 (N_11712,N_10532,N_9736);
nand U11713 (N_11713,N_10650,N_9900);
nand U11714 (N_11714,N_10266,N_10072);
nor U11715 (N_11715,N_9719,N_10609);
and U11716 (N_11716,N_10403,N_10567);
nor U11717 (N_11717,N_10029,N_10775);
nand U11718 (N_11718,N_10042,N_10464);
and U11719 (N_11719,N_10465,N_9793);
and U11720 (N_11720,N_9877,N_10417);
nand U11721 (N_11721,N_10776,N_10363);
nand U11722 (N_11722,N_10070,N_9892);
nor U11723 (N_11723,N_10179,N_9910);
nor U11724 (N_11724,N_10633,N_9613);
xnor U11725 (N_11725,N_9704,N_10047);
or U11726 (N_11726,N_10018,N_10283);
nor U11727 (N_11727,N_10798,N_10747);
or U11728 (N_11728,N_10470,N_9708);
or U11729 (N_11729,N_10073,N_9958);
or U11730 (N_11730,N_10409,N_10300);
xor U11731 (N_11731,N_10174,N_10290);
or U11732 (N_11732,N_9737,N_9796);
xnor U11733 (N_11733,N_9905,N_9746);
and U11734 (N_11734,N_9757,N_9989);
nand U11735 (N_11735,N_9798,N_10187);
and U11736 (N_11736,N_10759,N_9675);
or U11737 (N_11737,N_9604,N_10629);
nand U11738 (N_11738,N_9648,N_10206);
and U11739 (N_11739,N_10734,N_10126);
or U11740 (N_11740,N_9703,N_10120);
xnor U11741 (N_11741,N_10594,N_9796);
or U11742 (N_11742,N_10682,N_10166);
nor U11743 (N_11743,N_10016,N_9883);
xor U11744 (N_11744,N_9728,N_10061);
nand U11745 (N_11745,N_9946,N_9863);
and U11746 (N_11746,N_10223,N_10675);
nand U11747 (N_11747,N_10563,N_10698);
nor U11748 (N_11748,N_10421,N_10330);
and U11749 (N_11749,N_10166,N_9916);
nor U11750 (N_11750,N_10542,N_9605);
nor U11751 (N_11751,N_9645,N_10586);
and U11752 (N_11752,N_10721,N_10101);
nor U11753 (N_11753,N_9940,N_9798);
nand U11754 (N_11754,N_10638,N_10257);
xnor U11755 (N_11755,N_10704,N_10576);
and U11756 (N_11756,N_10132,N_10641);
nor U11757 (N_11757,N_9903,N_10452);
or U11758 (N_11758,N_10774,N_10153);
nand U11759 (N_11759,N_9644,N_10628);
and U11760 (N_11760,N_10760,N_10721);
nand U11761 (N_11761,N_10138,N_10048);
or U11762 (N_11762,N_9760,N_10501);
nand U11763 (N_11763,N_10016,N_10723);
nor U11764 (N_11764,N_10226,N_9698);
or U11765 (N_11765,N_9696,N_10656);
and U11766 (N_11766,N_9963,N_10149);
and U11767 (N_11767,N_10716,N_10437);
and U11768 (N_11768,N_10223,N_9891);
xnor U11769 (N_11769,N_10683,N_9989);
nand U11770 (N_11770,N_10331,N_9851);
or U11771 (N_11771,N_10612,N_9854);
xor U11772 (N_11772,N_10321,N_10718);
nand U11773 (N_11773,N_9656,N_9734);
and U11774 (N_11774,N_10607,N_10037);
or U11775 (N_11775,N_9929,N_9689);
nand U11776 (N_11776,N_9847,N_9960);
xnor U11777 (N_11777,N_10188,N_10632);
nand U11778 (N_11778,N_10765,N_9916);
nand U11779 (N_11779,N_10581,N_9674);
and U11780 (N_11780,N_9901,N_10631);
nor U11781 (N_11781,N_10298,N_10718);
or U11782 (N_11782,N_10329,N_9793);
nor U11783 (N_11783,N_9860,N_10589);
xnor U11784 (N_11784,N_9629,N_10589);
and U11785 (N_11785,N_10485,N_10658);
xnor U11786 (N_11786,N_10792,N_9994);
xnor U11787 (N_11787,N_10286,N_9880);
or U11788 (N_11788,N_10264,N_10129);
or U11789 (N_11789,N_10660,N_9768);
nor U11790 (N_11790,N_10500,N_9935);
xor U11791 (N_11791,N_9898,N_10747);
nand U11792 (N_11792,N_10584,N_10670);
nor U11793 (N_11793,N_10605,N_10143);
xor U11794 (N_11794,N_9687,N_9709);
and U11795 (N_11795,N_10761,N_9651);
xnor U11796 (N_11796,N_10625,N_10496);
nand U11797 (N_11797,N_9845,N_10569);
xor U11798 (N_11798,N_9805,N_9687);
and U11799 (N_11799,N_9656,N_9658);
xnor U11800 (N_11800,N_10422,N_10409);
nand U11801 (N_11801,N_10557,N_10727);
nor U11802 (N_11802,N_10319,N_10713);
xnor U11803 (N_11803,N_10056,N_10417);
or U11804 (N_11804,N_10167,N_10492);
xnor U11805 (N_11805,N_9663,N_10553);
and U11806 (N_11806,N_10154,N_9607);
xnor U11807 (N_11807,N_10388,N_9875);
xor U11808 (N_11808,N_10385,N_10649);
and U11809 (N_11809,N_10431,N_10626);
nand U11810 (N_11810,N_10754,N_9870);
and U11811 (N_11811,N_10515,N_10438);
and U11812 (N_11812,N_10210,N_9874);
nor U11813 (N_11813,N_9665,N_9929);
or U11814 (N_11814,N_10477,N_10502);
or U11815 (N_11815,N_9972,N_9676);
nor U11816 (N_11816,N_9871,N_9765);
xnor U11817 (N_11817,N_9947,N_9789);
nand U11818 (N_11818,N_10419,N_9603);
nor U11819 (N_11819,N_9964,N_9853);
nor U11820 (N_11820,N_10194,N_10567);
nor U11821 (N_11821,N_9712,N_9906);
nor U11822 (N_11822,N_10715,N_9991);
nand U11823 (N_11823,N_10023,N_10395);
nor U11824 (N_11824,N_9947,N_9974);
or U11825 (N_11825,N_9746,N_10244);
or U11826 (N_11826,N_10281,N_10005);
or U11827 (N_11827,N_9635,N_10615);
xor U11828 (N_11828,N_10539,N_9855);
nor U11829 (N_11829,N_9748,N_10695);
and U11830 (N_11830,N_9745,N_10601);
or U11831 (N_11831,N_9959,N_10050);
or U11832 (N_11832,N_10215,N_10592);
nor U11833 (N_11833,N_10696,N_9949);
xnor U11834 (N_11834,N_9982,N_10186);
nand U11835 (N_11835,N_10528,N_10295);
nand U11836 (N_11836,N_10704,N_10110);
or U11837 (N_11837,N_10464,N_9650);
or U11838 (N_11838,N_10764,N_10476);
nand U11839 (N_11839,N_10637,N_9603);
xor U11840 (N_11840,N_10296,N_9665);
nor U11841 (N_11841,N_9698,N_10602);
and U11842 (N_11842,N_10698,N_10237);
and U11843 (N_11843,N_10488,N_10411);
and U11844 (N_11844,N_9655,N_9715);
nand U11845 (N_11845,N_10044,N_10602);
nand U11846 (N_11846,N_10434,N_10711);
or U11847 (N_11847,N_10777,N_10078);
or U11848 (N_11848,N_10204,N_9918);
xor U11849 (N_11849,N_9699,N_9629);
or U11850 (N_11850,N_10506,N_9904);
xnor U11851 (N_11851,N_9802,N_9861);
or U11852 (N_11852,N_10704,N_9664);
xnor U11853 (N_11853,N_9878,N_10208);
nand U11854 (N_11854,N_9898,N_10041);
nor U11855 (N_11855,N_10387,N_10487);
and U11856 (N_11856,N_10476,N_9605);
nand U11857 (N_11857,N_10604,N_10222);
and U11858 (N_11858,N_10297,N_10309);
and U11859 (N_11859,N_9996,N_9747);
nand U11860 (N_11860,N_9754,N_10570);
nor U11861 (N_11861,N_10431,N_10524);
or U11862 (N_11862,N_10778,N_9731);
nand U11863 (N_11863,N_10537,N_10262);
nor U11864 (N_11864,N_10133,N_10597);
xnor U11865 (N_11865,N_10780,N_10254);
xor U11866 (N_11866,N_10664,N_10321);
xnor U11867 (N_11867,N_9783,N_9877);
nand U11868 (N_11868,N_10579,N_10082);
and U11869 (N_11869,N_10448,N_10624);
nand U11870 (N_11870,N_10711,N_10558);
nand U11871 (N_11871,N_10291,N_10606);
and U11872 (N_11872,N_9771,N_10788);
and U11873 (N_11873,N_10473,N_10693);
nand U11874 (N_11874,N_10220,N_9689);
or U11875 (N_11875,N_9718,N_9830);
or U11876 (N_11876,N_9960,N_10218);
or U11877 (N_11877,N_10693,N_10246);
and U11878 (N_11878,N_9637,N_10071);
nor U11879 (N_11879,N_10129,N_10195);
nor U11880 (N_11880,N_10130,N_9699);
nand U11881 (N_11881,N_10635,N_10052);
nand U11882 (N_11882,N_10482,N_10027);
xor U11883 (N_11883,N_10022,N_10773);
xor U11884 (N_11884,N_9946,N_9794);
and U11885 (N_11885,N_10388,N_9985);
xor U11886 (N_11886,N_9685,N_10476);
nor U11887 (N_11887,N_10470,N_10081);
xor U11888 (N_11888,N_10745,N_10328);
and U11889 (N_11889,N_10722,N_10176);
xnor U11890 (N_11890,N_9984,N_9866);
and U11891 (N_11891,N_10055,N_9739);
nand U11892 (N_11892,N_9723,N_10070);
xnor U11893 (N_11893,N_9772,N_10640);
or U11894 (N_11894,N_10142,N_10345);
or U11895 (N_11895,N_10450,N_10120);
and U11896 (N_11896,N_10396,N_10113);
nand U11897 (N_11897,N_10594,N_10531);
or U11898 (N_11898,N_10658,N_9616);
xnor U11899 (N_11899,N_10235,N_10458);
xor U11900 (N_11900,N_9920,N_9715);
or U11901 (N_11901,N_9927,N_10016);
nand U11902 (N_11902,N_10739,N_9804);
nand U11903 (N_11903,N_9783,N_10718);
and U11904 (N_11904,N_10663,N_10437);
xor U11905 (N_11905,N_9969,N_10521);
xor U11906 (N_11906,N_9623,N_10048);
xor U11907 (N_11907,N_9875,N_10569);
and U11908 (N_11908,N_10001,N_10173);
nor U11909 (N_11909,N_10476,N_10626);
nand U11910 (N_11910,N_10373,N_9762);
nor U11911 (N_11911,N_10664,N_10371);
nor U11912 (N_11912,N_10227,N_10373);
and U11913 (N_11913,N_9941,N_10327);
and U11914 (N_11914,N_10132,N_9689);
xor U11915 (N_11915,N_10464,N_10368);
nor U11916 (N_11916,N_10756,N_10469);
or U11917 (N_11917,N_9686,N_10779);
nand U11918 (N_11918,N_10101,N_10183);
nand U11919 (N_11919,N_10072,N_10677);
or U11920 (N_11920,N_9780,N_10021);
or U11921 (N_11921,N_10186,N_9745);
xor U11922 (N_11922,N_9685,N_10696);
and U11923 (N_11923,N_10240,N_10691);
nor U11924 (N_11924,N_9958,N_10466);
or U11925 (N_11925,N_10672,N_10353);
nor U11926 (N_11926,N_10413,N_10240);
or U11927 (N_11927,N_10185,N_10127);
xor U11928 (N_11928,N_10708,N_10002);
nor U11929 (N_11929,N_9680,N_10392);
and U11930 (N_11930,N_10534,N_10788);
and U11931 (N_11931,N_9999,N_9935);
xor U11932 (N_11932,N_10400,N_10614);
and U11933 (N_11933,N_10447,N_10387);
xnor U11934 (N_11934,N_10583,N_10379);
or U11935 (N_11935,N_10472,N_10304);
nor U11936 (N_11936,N_10510,N_9881);
nand U11937 (N_11937,N_10433,N_10759);
xnor U11938 (N_11938,N_9644,N_9714);
or U11939 (N_11939,N_10597,N_9958);
nand U11940 (N_11940,N_10228,N_9833);
or U11941 (N_11941,N_10492,N_9775);
and U11942 (N_11942,N_10651,N_9631);
and U11943 (N_11943,N_10788,N_9682);
and U11944 (N_11944,N_10725,N_10097);
xor U11945 (N_11945,N_9955,N_10284);
xor U11946 (N_11946,N_10055,N_10684);
nand U11947 (N_11947,N_10186,N_10299);
and U11948 (N_11948,N_10101,N_10404);
or U11949 (N_11949,N_10495,N_10660);
nor U11950 (N_11950,N_10058,N_9676);
and U11951 (N_11951,N_9730,N_10580);
nor U11952 (N_11952,N_9698,N_9962);
and U11953 (N_11953,N_9752,N_10446);
nor U11954 (N_11954,N_10645,N_10548);
nand U11955 (N_11955,N_10786,N_10379);
nor U11956 (N_11956,N_10354,N_9890);
and U11957 (N_11957,N_9660,N_10452);
and U11958 (N_11958,N_10725,N_10711);
nor U11959 (N_11959,N_10118,N_9643);
and U11960 (N_11960,N_10010,N_10307);
nand U11961 (N_11961,N_9790,N_10152);
nor U11962 (N_11962,N_10253,N_10490);
or U11963 (N_11963,N_10251,N_9623);
xor U11964 (N_11964,N_10196,N_9753);
nand U11965 (N_11965,N_9728,N_10621);
and U11966 (N_11966,N_9648,N_10243);
or U11967 (N_11967,N_9943,N_10626);
nor U11968 (N_11968,N_9760,N_9871);
and U11969 (N_11969,N_10328,N_9837);
or U11970 (N_11970,N_10384,N_9709);
xor U11971 (N_11971,N_10331,N_10754);
or U11972 (N_11972,N_9881,N_10529);
xnor U11973 (N_11973,N_10621,N_10224);
xor U11974 (N_11974,N_9827,N_10261);
nor U11975 (N_11975,N_9965,N_10614);
nor U11976 (N_11976,N_10590,N_9808);
nor U11977 (N_11977,N_9729,N_9626);
or U11978 (N_11978,N_10792,N_10114);
nor U11979 (N_11979,N_10221,N_10033);
and U11980 (N_11980,N_9704,N_9834);
or U11981 (N_11981,N_10653,N_9820);
or U11982 (N_11982,N_9630,N_10594);
nor U11983 (N_11983,N_10530,N_9903);
or U11984 (N_11984,N_10196,N_9826);
and U11985 (N_11985,N_9782,N_10402);
or U11986 (N_11986,N_10284,N_10317);
or U11987 (N_11987,N_9684,N_9694);
and U11988 (N_11988,N_9636,N_10740);
nand U11989 (N_11989,N_10082,N_10088);
or U11990 (N_11990,N_10589,N_10725);
and U11991 (N_11991,N_10483,N_9801);
nor U11992 (N_11992,N_9795,N_10692);
and U11993 (N_11993,N_10575,N_10648);
and U11994 (N_11994,N_9826,N_9928);
and U11995 (N_11995,N_10241,N_10229);
or U11996 (N_11996,N_9869,N_9975);
nand U11997 (N_11997,N_9745,N_10247);
or U11998 (N_11998,N_10479,N_9930);
nor U11999 (N_11999,N_9896,N_9696);
xor U12000 (N_12000,N_11583,N_11647);
or U12001 (N_12001,N_11851,N_11630);
and U12002 (N_12002,N_11992,N_10956);
and U12003 (N_12003,N_11748,N_11055);
xor U12004 (N_12004,N_11891,N_11920);
nor U12005 (N_12005,N_11935,N_10951);
or U12006 (N_12006,N_11423,N_11598);
or U12007 (N_12007,N_11167,N_11214);
xnor U12008 (N_12008,N_11464,N_10858);
nand U12009 (N_12009,N_11380,N_11028);
xnor U12010 (N_12010,N_11094,N_10846);
xor U12011 (N_12011,N_11868,N_11608);
nand U12012 (N_12012,N_10954,N_11073);
nor U12013 (N_12013,N_11922,N_11221);
nor U12014 (N_12014,N_11699,N_11930);
and U12015 (N_12015,N_11783,N_11714);
xnor U12016 (N_12016,N_11408,N_11189);
nand U12017 (N_12017,N_11373,N_10938);
nor U12018 (N_12018,N_10801,N_11774);
and U12019 (N_12019,N_11808,N_10897);
nor U12020 (N_12020,N_11792,N_11542);
and U12021 (N_12021,N_11599,N_11810);
nand U12022 (N_12022,N_11383,N_11601);
xor U12023 (N_12023,N_11365,N_10842);
nor U12024 (N_12024,N_11082,N_11220);
nor U12025 (N_12025,N_11689,N_11656);
or U12026 (N_12026,N_11275,N_11015);
xnor U12027 (N_12027,N_11024,N_11300);
nand U12028 (N_12028,N_10983,N_11159);
and U12029 (N_12029,N_10855,N_11097);
xor U12030 (N_12030,N_10918,N_11720);
nor U12031 (N_12031,N_11108,N_10882);
or U12032 (N_12032,N_11757,N_11861);
or U12033 (N_12033,N_11319,N_11512);
nor U12034 (N_12034,N_11865,N_10853);
xor U12035 (N_12035,N_11933,N_11048);
or U12036 (N_12036,N_11356,N_10915);
or U12037 (N_12037,N_11911,N_11118);
nor U12038 (N_12038,N_11923,N_11602);
xnor U12039 (N_12039,N_11832,N_11654);
xor U12040 (N_12040,N_11518,N_11660);
nor U12041 (N_12041,N_11676,N_11825);
xor U12042 (N_12042,N_11064,N_11467);
and U12043 (N_12043,N_11880,N_11270);
xnor U12044 (N_12044,N_10948,N_11716);
and U12045 (N_12045,N_11386,N_11404);
nor U12046 (N_12046,N_11709,N_11937);
and U12047 (N_12047,N_11560,N_11957);
xor U12048 (N_12048,N_10865,N_10850);
xnor U12049 (N_12049,N_11955,N_10848);
and U12050 (N_12050,N_11078,N_11162);
nand U12051 (N_12051,N_11492,N_11394);
nor U12052 (N_12052,N_11194,N_11201);
xor U12053 (N_12053,N_11322,N_11994);
nor U12054 (N_12054,N_11043,N_11762);
and U12055 (N_12055,N_11129,N_11781);
nor U12056 (N_12056,N_11860,N_10873);
nor U12057 (N_12057,N_11259,N_11795);
nand U12058 (N_12058,N_11068,N_11188);
and U12059 (N_12059,N_10917,N_11453);
nand U12060 (N_12060,N_11869,N_10978);
nand U12061 (N_12061,N_10970,N_11266);
nor U12062 (N_12062,N_11479,N_11369);
or U12063 (N_12063,N_11628,N_11023);
nand U12064 (N_12064,N_11669,N_11682);
or U12065 (N_12065,N_11537,N_11262);
or U12066 (N_12066,N_10941,N_10857);
or U12067 (N_12067,N_11848,N_11276);
nand U12068 (N_12068,N_10990,N_11744);
and U12069 (N_12069,N_11886,N_11085);
nor U12070 (N_12070,N_11375,N_11498);
or U12071 (N_12071,N_11847,N_11787);
nand U12072 (N_12072,N_11105,N_10867);
and U12073 (N_12073,N_11278,N_11508);
nand U12074 (N_12074,N_11501,N_10919);
or U12075 (N_12075,N_10987,N_10845);
nand U12076 (N_12076,N_11681,N_10875);
nand U12077 (N_12077,N_11874,N_10989);
xor U12078 (N_12078,N_11543,N_11326);
xor U12079 (N_12079,N_11791,N_11001);
nand U12080 (N_12080,N_10991,N_11496);
nand U12081 (N_12081,N_11577,N_11967);
and U12082 (N_12082,N_10922,N_11029);
and U12083 (N_12083,N_11587,N_11481);
xor U12084 (N_12084,N_11755,N_11605);
and U12085 (N_12085,N_11291,N_11663);
xnor U12086 (N_12086,N_11348,N_11251);
nand U12087 (N_12087,N_11160,N_11330);
nor U12088 (N_12088,N_10959,N_11113);
and U12089 (N_12089,N_11176,N_11741);
and U12090 (N_12090,N_11609,N_10843);
nor U12091 (N_12091,N_11797,N_11679);
and U12092 (N_12092,N_11405,N_11722);
and U12093 (N_12093,N_11511,N_11588);
nor U12094 (N_12094,N_10893,N_11149);
or U12095 (N_12095,N_11127,N_11554);
or U12096 (N_12096,N_11707,N_11364);
and U12097 (N_12097,N_10943,N_11416);
or U12098 (N_12098,N_11648,N_10981);
nor U12099 (N_12099,N_11273,N_11339);
and U12100 (N_12100,N_11528,N_11538);
or U12101 (N_12101,N_11455,N_11562);
and U12102 (N_12102,N_11968,N_11172);
or U12103 (N_12103,N_11604,N_10864);
or U12104 (N_12104,N_11711,N_11534);
or U12105 (N_12105,N_11314,N_11181);
xor U12106 (N_12106,N_10836,N_11017);
xnor U12107 (N_12107,N_11486,N_11510);
or U12108 (N_12108,N_11903,N_11777);
nor U12109 (N_12109,N_11051,N_11474);
xnor U12110 (N_12110,N_10929,N_11756);
xor U12111 (N_12111,N_11962,N_11209);
nor U12112 (N_12112,N_11739,N_11536);
or U12113 (N_12113,N_11087,N_11522);
nand U12114 (N_12114,N_11471,N_10886);
or U12115 (N_12115,N_11284,N_11288);
or U12116 (N_12116,N_11882,N_11858);
nor U12117 (N_12117,N_11584,N_10937);
or U12118 (N_12118,N_10820,N_10974);
and U12119 (N_12119,N_11135,N_11970);
nor U12120 (N_12120,N_10986,N_11378);
nand U12121 (N_12121,N_11089,N_11625);
nand U12122 (N_12122,N_11419,N_11845);
or U12123 (N_12123,N_10957,N_11204);
nor U12124 (N_12124,N_11140,N_11859);
nor U12125 (N_12125,N_10904,N_11008);
nor U12126 (N_12126,N_11460,N_11591);
or U12127 (N_12127,N_11828,N_11745);
or U12128 (N_12128,N_11547,N_11918);
or U12129 (N_12129,N_11377,N_11426);
or U12130 (N_12130,N_11523,N_11799);
or U12131 (N_12131,N_11134,N_11100);
nor U12132 (N_12132,N_11685,N_11264);
xnor U12133 (N_12133,N_10808,N_11837);
nor U12134 (N_12134,N_11086,N_11399);
nor U12135 (N_12135,N_11067,N_11713);
or U12136 (N_12136,N_11396,N_11084);
or U12137 (N_12137,N_11895,N_11506);
and U12138 (N_12138,N_11788,N_11246);
or U12139 (N_12139,N_10914,N_11873);
xor U12140 (N_12140,N_11296,N_11461);
and U12141 (N_12141,N_11458,N_11177);
nor U12142 (N_12142,N_11704,N_11030);
and U12143 (N_12143,N_11320,N_11947);
or U12144 (N_12144,N_11363,N_11574);
nand U12145 (N_12145,N_10913,N_11595);
or U12146 (N_12146,N_11727,N_11686);
and U12147 (N_12147,N_10976,N_11060);
nand U12148 (N_12148,N_11677,N_11803);
nand U12149 (N_12149,N_11907,N_11080);
nand U12150 (N_12150,N_10884,N_11042);
or U12151 (N_12151,N_10972,N_11179);
and U12152 (N_12152,N_10963,N_11710);
nand U12153 (N_12153,N_11842,N_11954);
or U12154 (N_12154,N_11995,N_11944);
nand U12155 (N_12155,N_11973,N_11693);
and U12156 (N_12156,N_11002,N_11462);
and U12157 (N_12157,N_11034,N_11431);
xnor U12158 (N_12158,N_11936,N_10924);
nand U12159 (N_12159,N_10926,N_11836);
and U12160 (N_12160,N_11312,N_11593);
and U12161 (N_12161,N_11374,N_10879);
nand U12162 (N_12162,N_10955,N_11611);
and U12163 (N_12163,N_11329,N_10979);
xnor U12164 (N_12164,N_11286,N_11432);
nand U12165 (N_12165,N_11645,N_11303);
nor U12166 (N_12166,N_11401,N_11564);
or U12167 (N_12167,N_11224,N_11589);
xnor U12168 (N_12168,N_10833,N_11126);
nand U12169 (N_12169,N_11892,N_11659);
and U12170 (N_12170,N_11387,N_11833);
nor U12171 (N_12171,N_11978,N_11991);
and U12172 (N_12172,N_10823,N_11996);
nor U12173 (N_12173,N_11767,N_10908);
nor U12174 (N_12174,N_11897,N_10909);
nand U12175 (N_12175,N_11768,N_11131);
nand U12176 (N_12176,N_11281,N_11723);
nand U12177 (N_12177,N_11195,N_11751);
nand U12178 (N_12178,N_11341,N_11505);
nand U12179 (N_12179,N_10999,N_11938);
and U12180 (N_12180,N_11899,N_11743);
nand U12181 (N_12181,N_11287,N_11603);
xnor U12182 (N_12182,N_11016,N_11184);
or U12183 (N_12183,N_11239,N_11697);
xnor U12184 (N_12184,N_11729,N_11249);
or U12185 (N_12185,N_11843,N_11446);
nand U12186 (N_12186,N_10898,N_11203);
nand U12187 (N_12187,N_10860,N_11227);
nor U12188 (N_12188,N_10852,N_11800);
or U12189 (N_12189,N_11893,N_11539);
or U12190 (N_12190,N_11207,N_11742);
nand U12191 (N_12191,N_11393,N_11457);
nand U12192 (N_12192,N_11726,N_11417);
nand U12193 (N_12193,N_11812,N_11411);
and U12194 (N_12194,N_11514,N_11494);
or U12195 (N_12195,N_11485,N_11785);
nand U12196 (N_12196,N_11620,N_11076);
nor U12197 (N_12197,N_11216,N_11237);
and U12198 (N_12198,N_11229,N_11305);
xor U12199 (N_12199,N_11888,N_11272);
nor U12200 (N_12200,N_10921,N_11403);
xnor U12201 (N_12201,N_11963,N_11894);
nor U12202 (N_12202,N_11489,N_10806);
nor U12203 (N_12203,N_11966,N_11794);
and U12204 (N_12204,N_11010,N_10835);
or U12205 (N_12205,N_11210,N_11213);
xnor U12206 (N_12206,N_11013,N_10807);
nor U12207 (N_12207,N_11548,N_11517);
and U12208 (N_12208,N_11703,N_11530);
and U12209 (N_12209,N_11324,N_10932);
xor U12210 (N_12210,N_11924,N_11032);
and U12211 (N_12211,N_11758,N_11362);
xor U12212 (N_12212,N_11946,N_11132);
xnor U12213 (N_12213,N_11580,N_11465);
nor U12214 (N_12214,N_10934,N_10911);
xor U12215 (N_12215,N_11083,N_11980);
nand U12216 (N_12216,N_11231,N_11174);
and U12217 (N_12217,N_10859,N_10838);
or U12218 (N_12218,N_11145,N_11077);
nand U12219 (N_12219,N_11804,N_10994);
or U12220 (N_12220,N_11052,N_11844);
nor U12221 (N_12221,N_11600,N_11503);
nor U12222 (N_12222,N_11635,N_11570);
nor U12223 (N_12223,N_11950,N_10993);
nor U12224 (N_12224,N_11949,N_11728);
and U12225 (N_12225,N_11056,N_11988);
nor U12226 (N_12226,N_10930,N_11355);
or U12227 (N_12227,N_10810,N_11306);
nand U12228 (N_12228,N_11345,N_11199);
nand U12229 (N_12229,N_11550,N_11391);
nor U12230 (N_12230,N_11765,N_11904);
or U12231 (N_12231,N_11119,N_11983);
nand U12232 (N_12232,N_11798,N_11629);
nand U12233 (N_12233,N_11137,N_11117);
or U12234 (N_12234,N_11336,N_11409);
and U12235 (N_12235,N_11876,N_11541);
and U12236 (N_12236,N_11071,N_10939);
nand U12237 (N_12237,N_11700,N_11932);
nor U12238 (N_12238,N_10878,N_10964);
nand U12239 (N_12239,N_11974,N_11525);
nand U12240 (N_12240,N_10856,N_11454);
nand U12241 (N_12241,N_11752,N_11053);
nand U12242 (N_12242,N_11096,N_11079);
and U12243 (N_12243,N_11780,N_11488);
nor U12244 (N_12244,N_11397,N_10803);
or U12245 (N_12245,N_11563,N_11658);
xnor U12246 (N_12246,N_11790,N_10984);
or U12247 (N_12247,N_11984,N_11524);
nand U12248 (N_12248,N_11243,N_11175);
xor U12249 (N_12249,N_11637,N_11219);
or U12250 (N_12250,N_11230,N_10899);
or U12251 (N_12251,N_11590,N_11680);
or U12252 (N_12252,N_11222,N_10923);
xor U12253 (N_12253,N_11597,N_11102);
nand U12254 (N_12254,N_11581,N_11621);
xor U12255 (N_12255,N_11657,N_11639);
or U12256 (N_12256,N_11821,N_11555);
xnor U12257 (N_12257,N_11725,N_11158);
xor U12258 (N_12258,N_11081,N_10805);
nand U12259 (N_12259,N_11116,N_10812);
or U12260 (N_12260,N_11552,N_11694);
and U12261 (N_12261,N_11687,N_11627);
nand U12262 (N_12262,N_11360,N_11665);
nor U12263 (N_12263,N_11255,N_11163);
or U12264 (N_12264,N_11823,N_11171);
nand U12265 (N_12265,N_11124,N_11025);
or U12266 (N_12266,N_10912,N_11826);
or U12267 (N_12267,N_11233,N_11338);
nor U12268 (N_12268,N_11395,N_10961);
nand U12269 (N_12269,N_11824,N_11141);
xnor U12270 (N_12270,N_11075,N_11817);
xor U12271 (N_12271,N_10834,N_10903);
xor U12272 (N_12272,N_11443,N_11340);
and U12273 (N_12273,N_11784,N_11573);
nor U12274 (N_12274,N_11003,N_11121);
nand U12275 (N_12275,N_11623,N_10829);
or U12276 (N_12276,N_11006,N_11989);
xnor U12277 (N_12277,N_11155,N_11244);
or U12278 (N_12278,N_11661,N_11749);
nor U12279 (N_12279,N_11835,N_11520);
xor U12280 (N_12280,N_10831,N_11939);
nand U12281 (N_12281,N_11425,N_11335);
nand U12282 (N_12282,N_11392,N_11011);
nor U12283 (N_12283,N_11532,N_11297);
nor U12284 (N_12284,N_11138,N_11265);
nor U12285 (N_12285,N_11301,N_10821);
xnor U12286 (N_12286,N_11381,N_11277);
xor U12287 (N_12287,N_11565,N_11066);
or U12288 (N_12288,N_10968,N_11200);
nor U12289 (N_12289,N_11434,N_10967);
nor U12290 (N_12290,N_11735,N_11822);
or U12291 (N_12291,N_10894,N_11917);
and U12292 (N_12292,N_11390,N_11279);
nor U12293 (N_12293,N_11830,N_11975);
and U12294 (N_12294,N_11971,N_10901);
or U12295 (N_12295,N_11410,N_10935);
or U12296 (N_12296,N_11688,N_11499);
xnor U12297 (N_12297,N_11317,N_11180);
and U12298 (N_12298,N_11065,N_11619);
xor U12299 (N_12299,N_11382,N_11695);
nor U12300 (N_12300,N_11667,N_10847);
nor U12301 (N_12301,N_10876,N_11849);
nor U12302 (N_12302,N_11986,N_11953);
nor U12303 (N_12303,N_11114,N_10871);
and U12304 (N_12304,N_11883,N_10815);
or U12305 (N_12305,N_10950,N_10969);
nor U12306 (N_12306,N_11857,N_11352);
or U12307 (N_12307,N_11979,N_11156);
nor U12308 (N_12308,N_11618,N_11906);
xor U12309 (N_12309,N_11225,N_11435);
nand U12310 (N_12310,N_11059,N_11846);
nand U12311 (N_12311,N_11106,N_10880);
xnor U12312 (N_12312,N_11579,N_11049);
or U12313 (N_12313,N_10851,N_11544);
nor U12314 (N_12314,N_11998,N_11109);
nand U12315 (N_12315,N_11981,N_10907);
nor U12316 (N_12316,N_11664,N_11092);
nand U12317 (N_12317,N_11128,N_11019);
nor U12318 (N_12318,N_10966,N_10872);
or U12319 (N_12319,N_11586,N_10940);
and U12320 (N_12320,N_10949,N_11235);
xnor U12321 (N_12321,N_11853,N_11351);
xor U12322 (N_12322,N_11307,N_11412);
xor U12323 (N_12323,N_11384,N_11027);
nand U12324 (N_12324,N_11640,N_11238);
xor U12325 (N_12325,N_10881,N_11746);
xor U12326 (N_12326,N_11232,N_11021);
xor U12327 (N_12327,N_11248,N_11805);
nor U12328 (N_12328,N_10804,N_11841);
nand U12329 (N_12329,N_11509,N_10952);
or U12330 (N_12330,N_11215,N_11031);
or U12331 (N_12331,N_11274,N_11942);
and U12332 (N_12332,N_11926,N_11678);
and U12333 (N_12333,N_11495,N_11368);
nand U12334 (N_12334,N_11125,N_11327);
nand U12335 (N_12335,N_11218,N_11941);
nand U12336 (N_12336,N_11014,N_11472);
nor U12337 (N_12337,N_10819,N_11234);
xor U12338 (N_12338,N_11890,N_11775);
xor U12339 (N_12339,N_11864,N_11643);
and U12340 (N_12340,N_11653,N_11101);
xor U12341 (N_12341,N_10892,N_11294);
nand U12342 (N_12342,N_11112,N_11072);
nor U12343 (N_12343,N_10927,N_11004);
or U12344 (N_12344,N_11298,N_11772);
and U12345 (N_12345,N_11371,N_11740);
nand U12346 (N_12346,N_11546,N_10887);
nor U12347 (N_12347,N_11925,N_10905);
nand U12348 (N_12348,N_11449,N_11931);
nand U12349 (N_12349,N_11183,N_11561);
or U12350 (N_12350,N_11424,N_11253);
nand U12351 (N_12351,N_11566,N_10985);
xnor U12352 (N_12352,N_11241,N_11582);
nand U12353 (N_12353,N_10802,N_11615);
nand U12354 (N_12354,N_11896,N_11263);
nor U12355 (N_12355,N_10866,N_11982);
and U12356 (N_12356,N_10925,N_10818);
nor U12357 (N_12357,N_11814,N_11650);
or U12358 (N_12358,N_11927,N_11107);
nand U12359 (N_12359,N_11347,N_11120);
nand U12360 (N_12360,N_10811,N_11045);
nor U12361 (N_12361,N_11884,N_11976);
or U12362 (N_12362,N_11507,N_11705);
nor U12363 (N_12363,N_11617,N_10869);
and U12364 (N_12364,N_11753,N_10861);
or U12365 (N_12365,N_11123,N_11407);
or U12366 (N_12366,N_11422,N_11044);
nand U12367 (N_12367,N_10916,N_11421);
nand U12368 (N_12368,N_11295,N_11267);
and U12369 (N_12369,N_11009,N_11228);
nand U12370 (N_12370,N_11690,N_11612);
nand U12371 (N_12371,N_11333,N_11683);
nand U12372 (N_12372,N_11456,N_11666);
nor U12373 (N_12373,N_11413,N_11437);
or U12374 (N_12374,N_11754,N_11737);
nor U12375 (N_12375,N_11929,N_11069);
and U12376 (N_12376,N_11719,N_10885);
nor U12377 (N_12377,N_11634,N_11182);
and U12378 (N_12378,N_11972,N_10971);
nor U12379 (N_12379,N_11477,N_11250);
xor U12380 (N_12380,N_11388,N_11299);
and U12381 (N_12381,N_11402,N_11557);
and U12382 (N_12382,N_11311,N_11773);
nand U12383 (N_12383,N_11959,N_10973);
nor U12384 (N_12384,N_11964,N_11304);
nor U12385 (N_12385,N_11448,N_11468);
or U12386 (N_12386,N_10888,N_11769);
and U12387 (N_12387,N_11838,N_11050);
and U12388 (N_12388,N_10975,N_11490);
xnor U12389 (N_12389,N_11576,N_11451);
or U12390 (N_12390,N_11875,N_11133);
and U12391 (N_12391,N_11631,N_11389);
xnor U12392 (N_12392,N_11855,N_11750);
xor U12393 (N_12393,N_11871,N_11342);
xor U12394 (N_12394,N_10928,N_11594);
nand U12395 (N_12395,N_11921,N_11475);
nor U12396 (N_12396,N_11000,N_11867);
xnor U12397 (N_12397,N_11254,N_11928);
and U12398 (N_12398,N_10832,N_10816);
or U12399 (N_12399,N_10946,N_11166);
or U12400 (N_12400,N_11436,N_11192);
or U12401 (N_12401,N_11771,N_11571);
or U12402 (N_12402,N_11271,N_11759);
and U12403 (N_12403,N_11041,N_11366);
nor U12404 (N_12404,N_11473,N_11961);
or U12405 (N_12405,N_11442,N_10817);
nand U12406 (N_12406,N_11318,N_11878);
xnor U12407 (N_12407,N_11385,N_11146);
nand U12408 (N_12408,N_11839,N_11951);
nor U12409 (N_12409,N_11807,N_11164);
or U12410 (N_12410,N_10814,N_11316);
xor U12411 (N_12411,N_11332,N_11139);
nor U12412 (N_12412,N_11840,N_10813);
nand U12413 (N_12413,N_10874,N_11684);
or U12414 (N_12414,N_10862,N_10824);
nand U12415 (N_12415,N_11104,N_11779);
nand U12416 (N_12416,N_11718,N_11872);
nand U12417 (N_12417,N_11018,N_10890);
nand U12418 (N_12418,N_11358,N_11881);
and U12419 (N_12419,N_11559,N_10995);
nand U12420 (N_12420,N_11236,N_11321);
and U12421 (N_12421,N_11062,N_11497);
or U12422 (N_12422,N_11208,N_11346);
and U12423 (N_12423,N_11242,N_11885);
xnor U12424 (N_12424,N_10910,N_10828);
xnor U12425 (N_12425,N_11433,N_11428);
or U12426 (N_12426,N_11913,N_10896);
nor U12427 (N_12427,N_11675,N_11724);
nor U12428 (N_12428,N_11103,N_11801);
nor U12429 (N_12429,N_11834,N_11914);
and U12430 (N_12430,N_11624,N_10849);
or U12431 (N_12431,N_11856,N_11061);
or U12432 (N_12432,N_11671,N_11877);
nand U12433 (N_12433,N_11802,N_11662);
nand U12434 (N_12434,N_10889,N_11247);
nor U12435 (N_12435,N_10841,N_10839);
or U12436 (N_12436,N_11952,N_11282);
nor U12437 (N_12437,N_11484,N_11353);
nor U12438 (N_12438,N_11551,N_10982);
xnor U12439 (N_12439,N_11793,N_11674);
and U12440 (N_12440,N_11379,N_11540);
nor U12441 (N_12441,N_11325,N_11022);
or U12442 (N_12442,N_11636,N_11429);
and U12443 (N_12443,N_11185,N_11870);
and U12444 (N_12444,N_11622,N_10830);
nor U12445 (N_12445,N_11111,N_11093);
nor U12446 (N_12446,N_11350,N_11202);
nor U12447 (N_12447,N_11691,N_11527);
nand U12448 (N_12448,N_11047,N_11285);
xnor U12449 (N_12449,N_11715,N_11596);
and U12450 (N_12450,N_11733,N_11500);
nand U12451 (N_12451,N_11058,N_11090);
and U12452 (N_12452,N_11673,N_11649);
and U12453 (N_12453,N_11493,N_11708);
nor U12454 (N_12454,N_10906,N_11398);
or U12455 (N_12455,N_11607,N_11901);
nand U12456 (N_12456,N_11161,N_11575);
or U12457 (N_12457,N_11879,N_11670);
nand U12458 (N_12458,N_11731,N_11651);
or U12459 (N_12459,N_10900,N_11909);
nand U12460 (N_12460,N_11212,N_11519);
nor U12461 (N_12461,N_11040,N_11110);
nor U12462 (N_12462,N_11313,N_11863);
and U12463 (N_12463,N_11960,N_10960);
or U12464 (N_12464,N_11887,N_11889);
xor U12465 (N_12465,N_11831,N_11323);
or U12466 (N_12466,N_11150,N_11337);
nand U12467 (N_12467,N_11290,N_11819);
and U12468 (N_12468,N_11761,N_11515);
nand U12469 (N_12469,N_11535,N_11652);
nor U12470 (N_12470,N_11706,N_11193);
nand U12471 (N_12471,N_11513,N_10870);
nand U12472 (N_12472,N_10844,N_10997);
nor U12473 (N_12473,N_11747,N_11736);
and U12474 (N_12474,N_11578,N_11148);
nand U12475 (N_12475,N_11007,N_11328);
or U12476 (N_12476,N_11796,N_11414);
or U12477 (N_12477,N_11070,N_11866);
xor U12478 (N_12478,N_11502,N_11459);
and U12479 (N_12479,N_11418,N_11668);
nor U12480 (N_12480,N_11349,N_11147);
or U12481 (N_12481,N_11440,N_11361);
xor U12482 (N_12482,N_10953,N_11898);
nor U12483 (N_12483,N_11260,N_11672);
xor U12484 (N_12484,N_11186,N_11144);
nor U12485 (N_12485,N_11430,N_11482);
or U12486 (N_12486,N_11463,N_11940);
xnor U12487 (N_12487,N_11122,N_11173);
xnor U12488 (N_12488,N_11191,N_10945);
or U12489 (N_12489,N_10958,N_10947);
nand U12490 (N_12490,N_11190,N_10931);
nor U12491 (N_12491,N_11533,N_11308);
nand U12492 (N_12492,N_11692,N_10998);
xnor U12493 (N_12493,N_11289,N_10895);
or U12494 (N_12494,N_11357,N_11447);
or U12495 (N_12495,N_11721,N_11655);
xor U12496 (N_12496,N_10920,N_11441);
nor U12497 (N_12497,N_11480,N_11354);
or U12498 (N_12498,N_11033,N_11789);
xnor U12499 (N_12499,N_11638,N_11256);
nor U12500 (N_12500,N_10933,N_11999);
nand U12501 (N_12501,N_11948,N_11919);
or U12502 (N_12502,N_11908,N_11526);
nand U12503 (N_12503,N_11763,N_11310);
nand U12504 (N_12504,N_11054,N_11099);
xor U12505 (N_12505,N_10837,N_10826);
nand U12506 (N_12506,N_11786,N_11445);
xnor U12507 (N_12507,N_11063,N_11343);
xor U12508 (N_12508,N_11730,N_11827);
or U12509 (N_12509,N_11035,N_10992);
xnor U12510 (N_12510,N_11717,N_11154);
xnor U12511 (N_12511,N_11038,N_11616);
nor U12512 (N_12512,N_11452,N_11257);
nor U12513 (N_12513,N_11626,N_11969);
and U12514 (N_12514,N_10854,N_11036);
or U12515 (N_12515,N_11206,N_11226);
nand U12516 (N_12516,N_11370,N_11037);
or U12517 (N_12517,N_11205,N_10988);
xnor U12518 (N_12518,N_11331,N_11558);
nor U12519 (N_12519,N_11197,N_11504);
or U12520 (N_12520,N_10942,N_11469);
nand U12521 (N_12521,N_11760,N_11606);
nand U12522 (N_12522,N_11487,N_11261);
nor U12523 (N_12523,N_11905,N_11698);
xor U12524 (N_12524,N_11439,N_11592);
nand U12525 (N_12525,N_11223,N_11211);
nor U12526 (N_12526,N_11444,N_11198);
nor U12527 (N_12527,N_11309,N_11633);
and U12528 (N_12528,N_11993,N_11269);
nand U12529 (N_12529,N_11491,N_11142);
and U12530 (N_12530,N_11902,N_11466);
nand U12531 (N_12531,N_11642,N_11151);
nor U12532 (N_12532,N_11240,N_10936);
xnor U12533 (N_12533,N_10827,N_10944);
xor U12534 (N_12534,N_11153,N_11367);
and U12535 (N_12535,N_11531,N_11567);
nand U12536 (N_12536,N_11529,N_10962);
xor U12537 (N_12537,N_11816,N_11420);
nand U12538 (N_12538,N_11545,N_11696);
xor U12539 (N_12539,N_11292,N_10840);
or U12540 (N_12540,N_11702,N_11977);
xor U12541 (N_12541,N_11157,N_11427);
nand U12542 (N_12542,N_11829,N_10977);
nand U12543 (N_12543,N_11738,N_11169);
and U12544 (N_12544,N_11585,N_11813);
nor U12545 (N_12545,N_11315,N_11569);
and U12546 (N_12546,N_11406,N_11302);
nand U12547 (N_12547,N_11088,N_10809);
xor U12548 (N_12548,N_11987,N_11012);
nand U12549 (N_12549,N_11641,N_11258);
or U12550 (N_12550,N_11701,N_11470);
nand U12551 (N_12551,N_11372,N_11990);
nand U12552 (N_12552,N_10996,N_11900);
nand U12553 (N_12553,N_11334,N_11170);
or U12554 (N_12554,N_11130,N_11811);
nand U12555 (N_12555,N_11136,N_11850);
nor U12556 (N_12556,N_11178,N_10902);
nand U12557 (N_12557,N_11252,N_11483);
or U12558 (N_12558,N_11644,N_11782);
or U12559 (N_12559,N_11516,N_11818);
or U12560 (N_12560,N_11521,N_11280);
or U12561 (N_12561,N_11965,N_11806);
nor U12562 (N_12562,N_10965,N_11268);
nor U12563 (N_12563,N_11074,N_11553);
xor U12564 (N_12564,N_11026,N_11187);
nor U12565 (N_12565,N_11934,N_11572);
xnor U12566 (N_12566,N_11165,N_11734);
and U12567 (N_12567,N_10822,N_11293);
or U12568 (N_12568,N_11852,N_11776);
nand U12569 (N_12569,N_11005,N_10883);
xor U12570 (N_12570,N_11958,N_11196);
nand U12571 (N_12571,N_11997,N_11376);
xnor U12572 (N_12572,N_11614,N_11820);
or U12573 (N_12573,N_11046,N_11712);
nor U12574 (N_12574,N_11400,N_10868);
or U12575 (N_12575,N_11912,N_11778);
and U12576 (N_12576,N_11152,N_11943);
xnor U12577 (N_12577,N_11985,N_11115);
and U12578 (N_12578,N_11020,N_11770);
nand U12579 (N_12579,N_11143,N_11168);
nand U12580 (N_12580,N_11764,N_10863);
nor U12581 (N_12581,N_11646,N_11415);
nand U12582 (N_12582,N_11910,N_11450);
nor U12583 (N_12583,N_11568,N_11438);
and U12584 (N_12584,N_11478,N_11613);
nand U12585 (N_12585,N_10825,N_11862);
or U12586 (N_12586,N_10877,N_11854);
nor U12587 (N_12587,N_10980,N_11057);
nand U12588 (N_12588,N_11217,N_11039);
or U12589 (N_12589,N_11095,N_11809);
nor U12590 (N_12590,N_11359,N_11915);
and U12591 (N_12591,N_11815,N_11091);
nor U12592 (N_12592,N_11766,N_11283);
or U12593 (N_12593,N_11632,N_11098);
or U12594 (N_12594,N_11549,N_11610);
or U12595 (N_12595,N_11344,N_11916);
nand U12596 (N_12596,N_11556,N_11245);
and U12597 (N_12597,N_10891,N_11945);
or U12598 (N_12598,N_11732,N_10800);
and U12599 (N_12599,N_11956,N_11476);
xor U12600 (N_12600,N_11459,N_11022);
xnor U12601 (N_12601,N_11366,N_11175);
or U12602 (N_12602,N_11576,N_11617);
xor U12603 (N_12603,N_11864,N_10936);
nand U12604 (N_12604,N_11308,N_10951);
nor U12605 (N_12605,N_11343,N_11987);
xnor U12606 (N_12606,N_11188,N_11191);
nand U12607 (N_12607,N_11853,N_11373);
and U12608 (N_12608,N_11316,N_11648);
nand U12609 (N_12609,N_11648,N_11751);
and U12610 (N_12610,N_11443,N_11150);
nor U12611 (N_12611,N_11713,N_11403);
and U12612 (N_12612,N_11875,N_11581);
or U12613 (N_12613,N_11820,N_11644);
xnor U12614 (N_12614,N_11142,N_11671);
or U12615 (N_12615,N_10836,N_11764);
xor U12616 (N_12616,N_10950,N_11021);
or U12617 (N_12617,N_11064,N_11824);
nand U12618 (N_12618,N_10887,N_11304);
and U12619 (N_12619,N_11813,N_11426);
and U12620 (N_12620,N_10868,N_11439);
xnor U12621 (N_12621,N_10979,N_11904);
xor U12622 (N_12622,N_11729,N_10926);
and U12623 (N_12623,N_11687,N_11113);
or U12624 (N_12624,N_11265,N_11246);
nor U12625 (N_12625,N_11149,N_11792);
and U12626 (N_12626,N_10933,N_11179);
nand U12627 (N_12627,N_11394,N_11081);
nand U12628 (N_12628,N_11109,N_11165);
and U12629 (N_12629,N_11186,N_10932);
and U12630 (N_12630,N_11164,N_11385);
or U12631 (N_12631,N_11269,N_11040);
nand U12632 (N_12632,N_10866,N_11765);
xor U12633 (N_12633,N_11949,N_11545);
and U12634 (N_12634,N_10900,N_11573);
xor U12635 (N_12635,N_11555,N_11794);
nor U12636 (N_12636,N_11913,N_11049);
xor U12637 (N_12637,N_10939,N_10921);
nand U12638 (N_12638,N_11504,N_10843);
or U12639 (N_12639,N_10855,N_11481);
nand U12640 (N_12640,N_11393,N_11281);
nand U12641 (N_12641,N_11578,N_11313);
nor U12642 (N_12642,N_10831,N_11585);
nor U12643 (N_12643,N_11277,N_11901);
and U12644 (N_12644,N_11461,N_11820);
nand U12645 (N_12645,N_11819,N_11019);
nand U12646 (N_12646,N_10985,N_11581);
nor U12647 (N_12647,N_11372,N_11417);
or U12648 (N_12648,N_11016,N_11252);
and U12649 (N_12649,N_11799,N_11986);
nand U12650 (N_12650,N_11638,N_11907);
nor U12651 (N_12651,N_11812,N_11049);
or U12652 (N_12652,N_11483,N_10839);
xor U12653 (N_12653,N_11461,N_10847);
nor U12654 (N_12654,N_11821,N_11497);
and U12655 (N_12655,N_11633,N_11508);
and U12656 (N_12656,N_11805,N_11025);
xor U12657 (N_12657,N_11956,N_11335);
xnor U12658 (N_12658,N_11168,N_10994);
and U12659 (N_12659,N_11842,N_11278);
and U12660 (N_12660,N_10859,N_11053);
or U12661 (N_12661,N_11736,N_11490);
xor U12662 (N_12662,N_11984,N_11489);
nand U12663 (N_12663,N_11390,N_11885);
nor U12664 (N_12664,N_10983,N_10896);
nor U12665 (N_12665,N_11149,N_10860);
or U12666 (N_12666,N_11468,N_11672);
and U12667 (N_12667,N_10981,N_11695);
and U12668 (N_12668,N_11092,N_11294);
or U12669 (N_12669,N_11697,N_11818);
nand U12670 (N_12670,N_10890,N_11251);
xor U12671 (N_12671,N_11749,N_11388);
or U12672 (N_12672,N_11109,N_11077);
and U12673 (N_12673,N_11558,N_11423);
xnor U12674 (N_12674,N_11728,N_11140);
nor U12675 (N_12675,N_11409,N_11123);
nor U12676 (N_12676,N_11317,N_11042);
nand U12677 (N_12677,N_10911,N_11927);
nor U12678 (N_12678,N_11406,N_11207);
or U12679 (N_12679,N_10962,N_11033);
nand U12680 (N_12680,N_11545,N_11736);
nor U12681 (N_12681,N_11021,N_11857);
nor U12682 (N_12682,N_10992,N_11077);
nand U12683 (N_12683,N_11405,N_11842);
and U12684 (N_12684,N_10801,N_11826);
xnor U12685 (N_12685,N_11887,N_11400);
or U12686 (N_12686,N_11015,N_10867);
or U12687 (N_12687,N_11466,N_11069);
and U12688 (N_12688,N_11323,N_11918);
nand U12689 (N_12689,N_11743,N_10869);
nor U12690 (N_12690,N_10985,N_11708);
nand U12691 (N_12691,N_11450,N_11092);
and U12692 (N_12692,N_11025,N_11159);
nand U12693 (N_12693,N_11018,N_11188);
nand U12694 (N_12694,N_11641,N_11614);
nand U12695 (N_12695,N_11680,N_11319);
or U12696 (N_12696,N_10990,N_11341);
xor U12697 (N_12697,N_11409,N_10880);
or U12698 (N_12698,N_11986,N_11577);
xnor U12699 (N_12699,N_11628,N_11131);
nand U12700 (N_12700,N_11782,N_11955);
and U12701 (N_12701,N_11173,N_10892);
nor U12702 (N_12702,N_10995,N_10965);
nand U12703 (N_12703,N_11112,N_11616);
nor U12704 (N_12704,N_11932,N_11375);
nor U12705 (N_12705,N_11709,N_11138);
xor U12706 (N_12706,N_10964,N_11236);
and U12707 (N_12707,N_11418,N_11482);
xor U12708 (N_12708,N_10990,N_11460);
or U12709 (N_12709,N_11560,N_11632);
xor U12710 (N_12710,N_11369,N_11445);
nor U12711 (N_12711,N_11471,N_11159);
nand U12712 (N_12712,N_11802,N_11806);
nand U12713 (N_12713,N_11123,N_11098);
and U12714 (N_12714,N_11886,N_11565);
nor U12715 (N_12715,N_10941,N_11885);
and U12716 (N_12716,N_10880,N_11046);
nand U12717 (N_12717,N_11093,N_11815);
nand U12718 (N_12718,N_10992,N_11028);
and U12719 (N_12719,N_11888,N_10903);
xor U12720 (N_12720,N_11583,N_11147);
and U12721 (N_12721,N_11242,N_11251);
xnor U12722 (N_12722,N_11630,N_11901);
nor U12723 (N_12723,N_11427,N_11658);
or U12724 (N_12724,N_10952,N_11708);
xnor U12725 (N_12725,N_11486,N_11065);
nand U12726 (N_12726,N_11800,N_11771);
nand U12727 (N_12727,N_10806,N_11143);
or U12728 (N_12728,N_10884,N_11074);
or U12729 (N_12729,N_11270,N_11366);
nand U12730 (N_12730,N_10899,N_11321);
xor U12731 (N_12731,N_11718,N_10825);
or U12732 (N_12732,N_11728,N_11875);
and U12733 (N_12733,N_11686,N_11064);
nand U12734 (N_12734,N_11416,N_11204);
xnor U12735 (N_12735,N_11066,N_11735);
nor U12736 (N_12736,N_11921,N_10908);
and U12737 (N_12737,N_11597,N_11082);
or U12738 (N_12738,N_11849,N_11028);
nor U12739 (N_12739,N_11946,N_11804);
xnor U12740 (N_12740,N_11193,N_11596);
and U12741 (N_12741,N_11421,N_10931);
and U12742 (N_12742,N_10872,N_11458);
nand U12743 (N_12743,N_10951,N_11479);
and U12744 (N_12744,N_11751,N_11600);
and U12745 (N_12745,N_11835,N_10801);
nor U12746 (N_12746,N_10878,N_11238);
xnor U12747 (N_12747,N_11833,N_10854);
xor U12748 (N_12748,N_10948,N_11190);
nor U12749 (N_12749,N_11098,N_11922);
nand U12750 (N_12750,N_11287,N_11552);
nand U12751 (N_12751,N_11598,N_11519);
and U12752 (N_12752,N_10883,N_11788);
xnor U12753 (N_12753,N_11068,N_11667);
nand U12754 (N_12754,N_11914,N_11609);
xor U12755 (N_12755,N_11986,N_11154);
nor U12756 (N_12756,N_11775,N_11005);
and U12757 (N_12757,N_11590,N_10812);
nor U12758 (N_12758,N_10890,N_11010);
or U12759 (N_12759,N_11702,N_10843);
or U12760 (N_12760,N_10817,N_10940);
and U12761 (N_12761,N_11074,N_11940);
and U12762 (N_12762,N_11636,N_11784);
and U12763 (N_12763,N_11440,N_11405);
xnor U12764 (N_12764,N_11127,N_11501);
nor U12765 (N_12765,N_10808,N_11546);
and U12766 (N_12766,N_11808,N_11114);
nor U12767 (N_12767,N_11149,N_11577);
nand U12768 (N_12768,N_11534,N_11397);
or U12769 (N_12769,N_11764,N_11474);
nand U12770 (N_12770,N_11212,N_11447);
xnor U12771 (N_12771,N_11737,N_11656);
nand U12772 (N_12772,N_11373,N_10887);
xor U12773 (N_12773,N_11032,N_11236);
nand U12774 (N_12774,N_10834,N_11132);
or U12775 (N_12775,N_11386,N_11269);
nand U12776 (N_12776,N_11149,N_11108);
nor U12777 (N_12777,N_11238,N_10827);
and U12778 (N_12778,N_11293,N_11945);
nor U12779 (N_12779,N_10886,N_11032);
and U12780 (N_12780,N_11620,N_11511);
and U12781 (N_12781,N_11015,N_11004);
nand U12782 (N_12782,N_11851,N_11464);
nand U12783 (N_12783,N_11326,N_10863);
xor U12784 (N_12784,N_11115,N_11231);
or U12785 (N_12785,N_11432,N_10880);
or U12786 (N_12786,N_11216,N_11392);
nand U12787 (N_12787,N_11041,N_11312);
and U12788 (N_12788,N_11603,N_11806);
nand U12789 (N_12789,N_10933,N_11029);
nand U12790 (N_12790,N_11832,N_11680);
and U12791 (N_12791,N_10994,N_11538);
nand U12792 (N_12792,N_11489,N_10930);
xor U12793 (N_12793,N_10941,N_11207);
and U12794 (N_12794,N_11053,N_11506);
nand U12795 (N_12795,N_10937,N_11694);
nor U12796 (N_12796,N_11020,N_11084);
nand U12797 (N_12797,N_11342,N_11994);
nand U12798 (N_12798,N_11810,N_11036);
or U12799 (N_12799,N_10894,N_11664);
and U12800 (N_12800,N_11806,N_11332);
or U12801 (N_12801,N_11429,N_11821);
nor U12802 (N_12802,N_11022,N_11326);
xnor U12803 (N_12803,N_11100,N_11449);
and U12804 (N_12804,N_11391,N_11707);
and U12805 (N_12805,N_11597,N_11214);
nor U12806 (N_12806,N_11512,N_10822);
xor U12807 (N_12807,N_11564,N_11173);
xnor U12808 (N_12808,N_11113,N_11580);
nor U12809 (N_12809,N_11063,N_10998);
nand U12810 (N_12810,N_11023,N_11334);
xnor U12811 (N_12811,N_11944,N_11205);
xor U12812 (N_12812,N_11456,N_11105);
and U12813 (N_12813,N_11712,N_11114);
xor U12814 (N_12814,N_11776,N_10986);
or U12815 (N_12815,N_11559,N_11791);
nand U12816 (N_12816,N_11120,N_11249);
nor U12817 (N_12817,N_11305,N_11379);
nor U12818 (N_12818,N_11520,N_11794);
nand U12819 (N_12819,N_11202,N_11456);
or U12820 (N_12820,N_11359,N_11772);
and U12821 (N_12821,N_10983,N_11289);
and U12822 (N_12822,N_11431,N_11225);
nand U12823 (N_12823,N_11800,N_11500);
nor U12824 (N_12824,N_10977,N_11422);
and U12825 (N_12825,N_11218,N_10893);
nand U12826 (N_12826,N_11600,N_11784);
or U12827 (N_12827,N_11260,N_11130);
or U12828 (N_12828,N_11576,N_11218);
or U12829 (N_12829,N_11154,N_11800);
or U12830 (N_12830,N_11431,N_11732);
and U12831 (N_12831,N_11503,N_11519);
nand U12832 (N_12832,N_10944,N_11259);
nand U12833 (N_12833,N_10945,N_11261);
or U12834 (N_12834,N_11911,N_11448);
or U12835 (N_12835,N_11911,N_11224);
and U12836 (N_12836,N_11656,N_11454);
nor U12837 (N_12837,N_11756,N_11019);
nor U12838 (N_12838,N_11524,N_11214);
xor U12839 (N_12839,N_11683,N_11230);
and U12840 (N_12840,N_11807,N_11312);
xnor U12841 (N_12841,N_11624,N_11702);
nand U12842 (N_12842,N_11524,N_11498);
nor U12843 (N_12843,N_11468,N_11308);
or U12844 (N_12844,N_11999,N_11994);
xor U12845 (N_12845,N_11977,N_11692);
or U12846 (N_12846,N_10940,N_11236);
nor U12847 (N_12847,N_11554,N_11668);
xnor U12848 (N_12848,N_11179,N_10856);
nor U12849 (N_12849,N_11880,N_11777);
or U12850 (N_12850,N_11860,N_11024);
nand U12851 (N_12851,N_11617,N_11355);
and U12852 (N_12852,N_11665,N_10807);
and U12853 (N_12853,N_11457,N_11029);
and U12854 (N_12854,N_10904,N_11692);
or U12855 (N_12855,N_11164,N_10809);
or U12856 (N_12856,N_11503,N_11167);
nand U12857 (N_12857,N_10969,N_11679);
and U12858 (N_12858,N_10956,N_11548);
or U12859 (N_12859,N_11899,N_10988);
nand U12860 (N_12860,N_11270,N_11482);
xnor U12861 (N_12861,N_10833,N_11067);
and U12862 (N_12862,N_11400,N_11288);
nor U12863 (N_12863,N_10823,N_11750);
nor U12864 (N_12864,N_11284,N_10810);
and U12865 (N_12865,N_11158,N_11372);
and U12866 (N_12866,N_10884,N_11417);
xnor U12867 (N_12867,N_11592,N_11312);
nor U12868 (N_12868,N_11609,N_10884);
and U12869 (N_12869,N_11482,N_11425);
or U12870 (N_12870,N_10862,N_11519);
nor U12871 (N_12871,N_11722,N_11116);
or U12872 (N_12872,N_10869,N_11073);
xnor U12873 (N_12873,N_11621,N_10881);
or U12874 (N_12874,N_11282,N_11426);
nand U12875 (N_12875,N_11129,N_11991);
or U12876 (N_12876,N_11496,N_10879);
or U12877 (N_12877,N_11576,N_11380);
and U12878 (N_12878,N_11292,N_11038);
xor U12879 (N_12879,N_10921,N_11241);
or U12880 (N_12880,N_11752,N_11039);
and U12881 (N_12881,N_11193,N_11170);
xnor U12882 (N_12882,N_11924,N_11245);
nand U12883 (N_12883,N_11513,N_11967);
xor U12884 (N_12884,N_11675,N_11656);
and U12885 (N_12885,N_11425,N_11695);
nand U12886 (N_12886,N_10895,N_11069);
or U12887 (N_12887,N_11915,N_11463);
nand U12888 (N_12888,N_10951,N_11257);
and U12889 (N_12889,N_11278,N_11908);
and U12890 (N_12890,N_11816,N_11263);
or U12891 (N_12891,N_11049,N_11773);
nor U12892 (N_12892,N_11616,N_11016);
and U12893 (N_12893,N_11587,N_11450);
and U12894 (N_12894,N_11325,N_11313);
and U12895 (N_12895,N_11582,N_10998);
or U12896 (N_12896,N_11500,N_11707);
xnor U12897 (N_12897,N_11051,N_11964);
nor U12898 (N_12898,N_10975,N_11897);
xnor U12899 (N_12899,N_10816,N_11554);
or U12900 (N_12900,N_11688,N_11220);
nor U12901 (N_12901,N_11524,N_11394);
xnor U12902 (N_12902,N_11894,N_10910);
xnor U12903 (N_12903,N_11326,N_11458);
or U12904 (N_12904,N_11734,N_10897);
nor U12905 (N_12905,N_10988,N_11766);
or U12906 (N_12906,N_11779,N_11250);
nand U12907 (N_12907,N_11614,N_11659);
and U12908 (N_12908,N_11528,N_11646);
and U12909 (N_12909,N_11108,N_11200);
nand U12910 (N_12910,N_11182,N_11924);
xor U12911 (N_12911,N_11257,N_11552);
and U12912 (N_12912,N_11565,N_11341);
xor U12913 (N_12913,N_10838,N_11050);
or U12914 (N_12914,N_11792,N_11152);
nand U12915 (N_12915,N_11089,N_10808);
and U12916 (N_12916,N_11601,N_10852);
xor U12917 (N_12917,N_11113,N_11856);
nand U12918 (N_12918,N_11785,N_11764);
nor U12919 (N_12919,N_11152,N_11814);
nand U12920 (N_12920,N_11350,N_11018);
xnor U12921 (N_12921,N_11085,N_11191);
xor U12922 (N_12922,N_11113,N_11752);
and U12923 (N_12923,N_11604,N_11326);
and U12924 (N_12924,N_11340,N_11737);
and U12925 (N_12925,N_11479,N_11153);
or U12926 (N_12926,N_10882,N_11474);
nor U12927 (N_12927,N_11881,N_11534);
nand U12928 (N_12928,N_10855,N_11463);
and U12929 (N_12929,N_11650,N_11850);
xor U12930 (N_12930,N_11772,N_11237);
nor U12931 (N_12931,N_11107,N_10835);
and U12932 (N_12932,N_11442,N_11049);
and U12933 (N_12933,N_11104,N_11690);
xor U12934 (N_12934,N_11139,N_11861);
xor U12935 (N_12935,N_11306,N_11966);
and U12936 (N_12936,N_11004,N_11145);
xor U12937 (N_12937,N_11266,N_11570);
xnor U12938 (N_12938,N_11238,N_10997);
nand U12939 (N_12939,N_11817,N_10914);
nand U12940 (N_12940,N_10850,N_11675);
nand U12941 (N_12941,N_10971,N_10824);
nor U12942 (N_12942,N_11438,N_11878);
or U12943 (N_12943,N_10940,N_11727);
or U12944 (N_12944,N_11832,N_11502);
xnor U12945 (N_12945,N_11988,N_11340);
and U12946 (N_12946,N_11335,N_11272);
xnor U12947 (N_12947,N_11442,N_11191);
xnor U12948 (N_12948,N_11957,N_11689);
nand U12949 (N_12949,N_11891,N_10955);
xor U12950 (N_12950,N_11256,N_11849);
and U12951 (N_12951,N_11920,N_11613);
nand U12952 (N_12952,N_11024,N_11700);
or U12953 (N_12953,N_11336,N_11108);
and U12954 (N_12954,N_11292,N_11205);
and U12955 (N_12955,N_11372,N_11439);
xor U12956 (N_12956,N_11448,N_11404);
or U12957 (N_12957,N_11338,N_11245);
xnor U12958 (N_12958,N_11717,N_11121);
xnor U12959 (N_12959,N_11334,N_11401);
xor U12960 (N_12960,N_11163,N_11398);
xor U12961 (N_12961,N_11716,N_11343);
nand U12962 (N_12962,N_10993,N_11888);
or U12963 (N_12963,N_11671,N_10984);
nand U12964 (N_12964,N_11953,N_11178);
nand U12965 (N_12965,N_11017,N_11312);
and U12966 (N_12966,N_10997,N_10977);
nor U12967 (N_12967,N_10915,N_10841);
nand U12968 (N_12968,N_11986,N_11811);
or U12969 (N_12969,N_10871,N_11280);
and U12970 (N_12970,N_11917,N_11723);
nor U12971 (N_12971,N_10886,N_11072);
nor U12972 (N_12972,N_11228,N_11527);
or U12973 (N_12973,N_11186,N_10992);
xor U12974 (N_12974,N_10810,N_11876);
nor U12975 (N_12975,N_11253,N_11258);
or U12976 (N_12976,N_11083,N_11813);
or U12977 (N_12977,N_11623,N_11048);
xnor U12978 (N_12978,N_11555,N_11231);
xnor U12979 (N_12979,N_11630,N_11718);
xnor U12980 (N_12980,N_10829,N_11258);
and U12981 (N_12981,N_11926,N_11514);
or U12982 (N_12982,N_11089,N_11861);
or U12983 (N_12983,N_11247,N_11181);
or U12984 (N_12984,N_11865,N_11540);
or U12985 (N_12985,N_11557,N_11718);
xnor U12986 (N_12986,N_10971,N_11428);
or U12987 (N_12987,N_11546,N_11631);
nor U12988 (N_12988,N_11215,N_11942);
nor U12989 (N_12989,N_11432,N_11327);
nand U12990 (N_12990,N_11650,N_11979);
xnor U12991 (N_12991,N_11485,N_10804);
xor U12992 (N_12992,N_10887,N_10830);
or U12993 (N_12993,N_11788,N_11994);
or U12994 (N_12994,N_11534,N_11087);
nand U12995 (N_12995,N_11812,N_11382);
or U12996 (N_12996,N_11447,N_11637);
and U12997 (N_12997,N_11731,N_10880);
nand U12998 (N_12998,N_11506,N_11937);
or U12999 (N_12999,N_11921,N_11209);
or U13000 (N_13000,N_11244,N_11673);
nor U13001 (N_13001,N_11151,N_11979);
xor U13002 (N_13002,N_10855,N_10880);
nor U13003 (N_13003,N_11950,N_10912);
and U13004 (N_13004,N_11121,N_10867);
xor U13005 (N_13005,N_11107,N_11945);
and U13006 (N_13006,N_11258,N_11526);
nand U13007 (N_13007,N_11770,N_10815);
xnor U13008 (N_13008,N_11037,N_11481);
nand U13009 (N_13009,N_11772,N_11552);
nand U13010 (N_13010,N_11345,N_10898);
nand U13011 (N_13011,N_11785,N_11864);
nor U13012 (N_13012,N_11515,N_10952);
nand U13013 (N_13013,N_11179,N_11616);
nor U13014 (N_13014,N_11163,N_11947);
xnor U13015 (N_13015,N_11170,N_11068);
nor U13016 (N_13016,N_11155,N_11200);
nand U13017 (N_13017,N_10973,N_11565);
and U13018 (N_13018,N_11609,N_11812);
xor U13019 (N_13019,N_11591,N_11195);
nand U13020 (N_13020,N_11276,N_11317);
nand U13021 (N_13021,N_11961,N_10832);
or U13022 (N_13022,N_10860,N_11221);
xor U13023 (N_13023,N_11016,N_11775);
or U13024 (N_13024,N_11088,N_11190);
xnor U13025 (N_13025,N_11679,N_11626);
and U13026 (N_13026,N_10893,N_10849);
or U13027 (N_13027,N_11225,N_11837);
and U13028 (N_13028,N_11888,N_11819);
and U13029 (N_13029,N_11534,N_11242);
and U13030 (N_13030,N_11920,N_11633);
nor U13031 (N_13031,N_10857,N_11235);
xor U13032 (N_13032,N_11992,N_11747);
nand U13033 (N_13033,N_11552,N_11479);
and U13034 (N_13034,N_11060,N_11231);
xnor U13035 (N_13035,N_11944,N_10884);
nor U13036 (N_13036,N_11305,N_11740);
xnor U13037 (N_13037,N_11963,N_10874);
or U13038 (N_13038,N_11469,N_11543);
xor U13039 (N_13039,N_11653,N_11549);
or U13040 (N_13040,N_11862,N_11913);
nor U13041 (N_13041,N_11214,N_11663);
or U13042 (N_13042,N_11007,N_10965);
nand U13043 (N_13043,N_11571,N_11029);
nand U13044 (N_13044,N_11379,N_11280);
nor U13045 (N_13045,N_11402,N_11462);
xnor U13046 (N_13046,N_11200,N_11470);
nand U13047 (N_13047,N_11214,N_11026);
and U13048 (N_13048,N_11119,N_11904);
nand U13049 (N_13049,N_11378,N_11705);
nand U13050 (N_13050,N_11341,N_11874);
or U13051 (N_13051,N_11226,N_11616);
or U13052 (N_13052,N_10865,N_11490);
nor U13053 (N_13053,N_11489,N_11429);
xor U13054 (N_13054,N_11778,N_11120);
and U13055 (N_13055,N_11040,N_11925);
nand U13056 (N_13056,N_11466,N_10914);
or U13057 (N_13057,N_10824,N_11394);
and U13058 (N_13058,N_10927,N_11996);
and U13059 (N_13059,N_10897,N_11613);
and U13060 (N_13060,N_11918,N_10814);
and U13061 (N_13061,N_11102,N_11754);
or U13062 (N_13062,N_10965,N_11739);
nor U13063 (N_13063,N_11229,N_11513);
or U13064 (N_13064,N_11774,N_11585);
xor U13065 (N_13065,N_11772,N_11304);
and U13066 (N_13066,N_10905,N_11973);
and U13067 (N_13067,N_11566,N_10802);
or U13068 (N_13068,N_11307,N_11837);
or U13069 (N_13069,N_10997,N_11572);
nand U13070 (N_13070,N_11979,N_11688);
and U13071 (N_13071,N_11530,N_11456);
nand U13072 (N_13072,N_11022,N_11461);
nand U13073 (N_13073,N_11398,N_11961);
and U13074 (N_13074,N_10802,N_11743);
or U13075 (N_13075,N_11541,N_11107);
xor U13076 (N_13076,N_11727,N_11220);
xor U13077 (N_13077,N_11432,N_11394);
nand U13078 (N_13078,N_11522,N_11650);
xor U13079 (N_13079,N_10934,N_11790);
nand U13080 (N_13080,N_11825,N_10896);
or U13081 (N_13081,N_11601,N_11587);
nand U13082 (N_13082,N_11530,N_11845);
and U13083 (N_13083,N_11159,N_11693);
or U13084 (N_13084,N_11529,N_10819);
nor U13085 (N_13085,N_11484,N_11415);
and U13086 (N_13086,N_11129,N_11564);
nor U13087 (N_13087,N_11510,N_11779);
or U13088 (N_13088,N_11042,N_11213);
and U13089 (N_13089,N_10932,N_11662);
nand U13090 (N_13090,N_11179,N_11721);
xor U13091 (N_13091,N_11348,N_11959);
nor U13092 (N_13092,N_11843,N_10910);
nand U13093 (N_13093,N_11161,N_10990);
nor U13094 (N_13094,N_11573,N_10878);
or U13095 (N_13095,N_11246,N_11150);
xnor U13096 (N_13096,N_11725,N_10886);
or U13097 (N_13097,N_11697,N_10907);
nand U13098 (N_13098,N_11503,N_11255);
nor U13099 (N_13099,N_11144,N_11872);
or U13100 (N_13100,N_11492,N_11435);
or U13101 (N_13101,N_11276,N_11036);
xor U13102 (N_13102,N_11656,N_11998);
and U13103 (N_13103,N_11247,N_11214);
or U13104 (N_13104,N_11128,N_11356);
or U13105 (N_13105,N_11940,N_11890);
nor U13106 (N_13106,N_11488,N_10831);
and U13107 (N_13107,N_11224,N_11256);
nand U13108 (N_13108,N_11257,N_11993);
nand U13109 (N_13109,N_10853,N_11850);
and U13110 (N_13110,N_10895,N_11040);
or U13111 (N_13111,N_10906,N_10974);
xnor U13112 (N_13112,N_11831,N_11340);
or U13113 (N_13113,N_10911,N_11250);
and U13114 (N_13114,N_11170,N_10986);
or U13115 (N_13115,N_11778,N_11198);
and U13116 (N_13116,N_11686,N_11618);
nand U13117 (N_13117,N_11325,N_11404);
and U13118 (N_13118,N_11129,N_11346);
and U13119 (N_13119,N_10829,N_11659);
nand U13120 (N_13120,N_11026,N_11538);
nand U13121 (N_13121,N_10840,N_11374);
nand U13122 (N_13122,N_11270,N_11138);
nand U13123 (N_13123,N_11981,N_10939);
and U13124 (N_13124,N_11131,N_11759);
xor U13125 (N_13125,N_11597,N_11514);
and U13126 (N_13126,N_11263,N_11650);
or U13127 (N_13127,N_11524,N_11710);
or U13128 (N_13128,N_11794,N_11455);
nand U13129 (N_13129,N_11452,N_11170);
nand U13130 (N_13130,N_10883,N_11051);
xnor U13131 (N_13131,N_11675,N_11403);
nand U13132 (N_13132,N_11626,N_11946);
and U13133 (N_13133,N_11306,N_11597);
xor U13134 (N_13134,N_10880,N_11702);
nand U13135 (N_13135,N_11911,N_11252);
xnor U13136 (N_13136,N_10844,N_11470);
and U13137 (N_13137,N_11597,N_11189);
xor U13138 (N_13138,N_11356,N_11850);
and U13139 (N_13139,N_11624,N_11504);
xor U13140 (N_13140,N_11732,N_11615);
nand U13141 (N_13141,N_11539,N_11854);
xor U13142 (N_13142,N_11490,N_11924);
nand U13143 (N_13143,N_11990,N_11700);
or U13144 (N_13144,N_11339,N_11514);
nand U13145 (N_13145,N_10934,N_11165);
and U13146 (N_13146,N_10961,N_11948);
nor U13147 (N_13147,N_11741,N_11411);
and U13148 (N_13148,N_11448,N_11062);
and U13149 (N_13149,N_11138,N_11407);
and U13150 (N_13150,N_11441,N_11137);
or U13151 (N_13151,N_10972,N_10939);
or U13152 (N_13152,N_11003,N_10932);
nand U13153 (N_13153,N_10927,N_11203);
nor U13154 (N_13154,N_11961,N_11489);
nor U13155 (N_13155,N_11756,N_11861);
nor U13156 (N_13156,N_11582,N_11876);
nand U13157 (N_13157,N_11440,N_11446);
and U13158 (N_13158,N_11985,N_11398);
xor U13159 (N_13159,N_11676,N_11527);
or U13160 (N_13160,N_11143,N_11884);
or U13161 (N_13161,N_11377,N_11063);
and U13162 (N_13162,N_11851,N_10884);
nor U13163 (N_13163,N_11777,N_11028);
or U13164 (N_13164,N_10996,N_11658);
nor U13165 (N_13165,N_10805,N_11089);
and U13166 (N_13166,N_11517,N_11519);
or U13167 (N_13167,N_11742,N_11300);
xnor U13168 (N_13168,N_11839,N_10821);
and U13169 (N_13169,N_11291,N_11236);
nand U13170 (N_13170,N_11585,N_11765);
xor U13171 (N_13171,N_11979,N_11434);
and U13172 (N_13172,N_11856,N_10821);
nor U13173 (N_13173,N_11607,N_11239);
nor U13174 (N_13174,N_11583,N_11680);
or U13175 (N_13175,N_11698,N_11049);
xor U13176 (N_13176,N_11672,N_11433);
xor U13177 (N_13177,N_11012,N_11503);
xor U13178 (N_13178,N_11784,N_11408);
xor U13179 (N_13179,N_11507,N_11445);
nand U13180 (N_13180,N_11863,N_11061);
xor U13181 (N_13181,N_11949,N_11745);
and U13182 (N_13182,N_11451,N_11589);
nand U13183 (N_13183,N_11216,N_11579);
or U13184 (N_13184,N_11461,N_11995);
nand U13185 (N_13185,N_11044,N_11370);
and U13186 (N_13186,N_11785,N_11032);
or U13187 (N_13187,N_10885,N_11117);
nand U13188 (N_13188,N_11750,N_11881);
or U13189 (N_13189,N_11971,N_10899);
nand U13190 (N_13190,N_11769,N_11727);
or U13191 (N_13191,N_11930,N_10942);
and U13192 (N_13192,N_11508,N_10925);
nor U13193 (N_13193,N_11229,N_11409);
xnor U13194 (N_13194,N_11501,N_11475);
or U13195 (N_13195,N_11561,N_11052);
nand U13196 (N_13196,N_11172,N_11885);
nand U13197 (N_13197,N_10821,N_10936);
and U13198 (N_13198,N_11009,N_11314);
xnor U13199 (N_13199,N_11545,N_11886);
or U13200 (N_13200,N_13177,N_12542);
or U13201 (N_13201,N_12778,N_12565);
nor U13202 (N_13202,N_12659,N_12388);
or U13203 (N_13203,N_12651,N_13089);
or U13204 (N_13204,N_13170,N_12309);
xor U13205 (N_13205,N_12324,N_12256);
xor U13206 (N_13206,N_12394,N_12128);
nand U13207 (N_13207,N_12684,N_12197);
xnor U13208 (N_13208,N_12531,N_12698);
and U13209 (N_13209,N_12906,N_12902);
xnor U13210 (N_13210,N_12610,N_12200);
nand U13211 (N_13211,N_12494,N_13025);
xor U13212 (N_13212,N_13032,N_12119);
nand U13213 (N_13213,N_13001,N_13061);
xor U13214 (N_13214,N_12836,N_13048);
and U13215 (N_13215,N_12399,N_12796);
and U13216 (N_13216,N_13059,N_12598);
xor U13217 (N_13217,N_12093,N_12992);
nor U13218 (N_13218,N_12439,N_12467);
nor U13219 (N_13219,N_12122,N_12697);
and U13220 (N_13220,N_12535,N_12809);
xor U13221 (N_13221,N_13005,N_12843);
or U13222 (N_13222,N_12340,N_13006);
xor U13223 (N_13223,N_12749,N_12295);
or U13224 (N_13224,N_13069,N_12202);
nand U13225 (N_13225,N_12244,N_12035);
xor U13226 (N_13226,N_12383,N_12515);
and U13227 (N_13227,N_12743,N_12053);
xor U13228 (N_13228,N_12374,N_12660);
nor U13229 (N_13229,N_12553,N_13159);
xor U13230 (N_13230,N_13096,N_12036);
nand U13231 (N_13231,N_12502,N_12260);
nor U13232 (N_13232,N_12290,N_13045);
nand U13233 (N_13233,N_12678,N_12158);
xor U13234 (N_13234,N_13003,N_13126);
xnor U13235 (N_13235,N_12069,N_12418);
nor U13236 (N_13236,N_12603,N_12821);
xnor U13237 (N_13237,N_12478,N_12692);
nor U13238 (N_13238,N_12572,N_12832);
and U13239 (N_13239,N_12996,N_12788);
or U13240 (N_13240,N_12852,N_12914);
nand U13241 (N_13241,N_12875,N_12322);
nor U13242 (N_13242,N_12503,N_12304);
nor U13243 (N_13243,N_13109,N_12686);
nor U13244 (N_13244,N_12928,N_12756);
nor U13245 (N_13245,N_12163,N_12674);
nand U13246 (N_13246,N_12168,N_12916);
and U13247 (N_13247,N_12228,N_13152);
xor U13248 (N_13248,N_12261,N_12373);
nand U13249 (N_13249,N_12380,N_12777);
and U13250 (N_13250,N_12847,N_12386);
or U13251 (N_13251,N_12953,N_12646);
xnor U13252 (N_13252,N_12900,N_12537);
nand U13253 (N_13253,N_12766,N_13018);
or U13254 (N_13254,N_12129,N_12084);
nor U13255 (N_13255,N_12140,N_12614);
or U13256 (N_13256,N_12316,N_12658);
and U13257 (N_13257,N_12799,N_13033);
xnor U13258 (N_13258,N_13141,N_13078);
or U13259 (N_13259,N_12476,N_12496);
xnor U13260 (N_13260,N_12811,N_12030);
nor U13261 (N_13261,N_12428,N_12438);
or U13262 (N_13262,N_12520,N_12637);
and U13263 (N_13263,N_12074,N_13062);
or U13264 (N_13264,N_12980,N_12219);
or U13265 (N_13265,N_12301,N_12525);
nor U13266 (N_13266,N_12206,N_13042);
or U13267 (N_13267,N_12020,N_12458);
or U13268 (N_13268,N_12818,N_12524);
xnor U13269 (N_13269,N_12712,N_12576);
nand U13270 (N_13270,N_12861,N_13066);
xnor U13271 (N_13271,N_12628,N_12761);
nand U13272 (N_13272,N_12465,N_12689);
and U13273 (N_13273,N_12544,N_13028);
and U13274 (N_13274,N_12123,N_12946);
nand U13275 (N_13275,N_12078,N_13154);
and U13276 (N_13276,N_12456,N_12250);
or U13277 (N_13277,N_12680,N_12048);
and U13278 (N_13278,N_13172,N_12564);
nand U13279 (N_13279,N_12822,N_12556);
nor U13280 (N_13280,N_12973,N_12594);
nand U13281 (N_13281,N_12839,N_13083);
or U13282 (N_13282,N_13110,N_12785);
xnor U13283 (N_13283,N_12014,N_13081);
xnor U13284 (N_13284,N_12563,N_13161);
and U13285 (N_13285,N_12171,N_13046);
nand U13286 (N_13286,N_12247,N_12733);
nand U13287 (N_13287,N_13142,N_12714);
nand U13288 (N_13288,N_12487,N_12349);
xnor U13289 (N_13289,N_13073,N_12488);
or U13290 (N_13290,N_12612,N_12462);
xnor U13291 (N_13291,N_13180,N_12229);
nor U13292 (N_13292,N_12237,N_12509);
nor U13293 (N_13293,N_12242,N_13162);
nand U13294 (N_13294,N_12470,N_13144);
and U13295 (N_13295,N_13104,N_12518);
nand U13296 (N_13296,N_12688,N_12676);
and U13297 (N_13297,N_12949,N_13027);
xnor U13298 (N_13298,N_12210,N_12963);
nor U13299 (N_13299,N_12956,N_12609);
and U13300 (N_13300,N_13071,N_13056);
nand U13301 (N_13301,N_12960,N_12728);
xnor U13302 (N_13302,N_12006,N_13074);
or U13303 (N_13303,N_12273,N_12246);
and U13304 (N_13304,N_13135,N_12395);
nand U13305 (N_13305,N_12073,N_12067);
and U13306 (N_13306,N_12241,N_12480);
or U13307 (N_13307,N_12055,N_12501);
or U13308 (N_13308,N_12408,N_12879);
and U13309 (N_13309,N_12725,N_12049);
nand U13310 (N_13310,N_12357,N_12224);
nand U13311 (N_13311,N_12816,N_12367);
xnor U13312 (N_13312,N_12338,N_12891);
and U13313 (N_13313,N_12829,N_13125);
nor U13314 (N_13314,N_12271,N_13002);
nand U13315 (N_13315,N_12257,N_12846);
nor U13316 (N_13316,N_12924,N_12411);
nand U13317 (N_13317,N_12884,N_12457);
and U13318 (N_13318,N_12893,N_13167);
and U13319 (N_13319,N_12072,N_13053);
or U13320 (N_13320,N_12189,N_12767);
or U13321 (N_13321,N_12016,N_12300);
or U13322 (N_13322,N_13097,N_12166);
or U13323 (N_13323,N_12560,N_13166);
or U13324 (N_13324,N_13014,N_12987);
nor U13325 (N_13325,N_12514,N_12033);
xnor U13326 (N_13326,N_12280,N_12505);
xor U13327 (N_13327,N_13191,N_12976);
or U13328 (N_13328,N_13124,N_12499);
xor U13329 (N_13329,N_12274,N_12003);
or U13330 (N_13330,N_12876,N_12240);
xor U13331 (N_13331,N_12389,N_12826);
and U13332 (N_13332,N_12112,N_12474);
and U13333 (N_13333,N_13108,N_12360);
or U13334 (N_13334,N_12056,N_12508);
or U13335 (N_13335,N_13060,N_12732);
xor U13336 (N_13336,N_12957,N_12729);
nor U13337 (N_13337,N_12387,N_12406);
nand U13338 (N_13338,N_13149,N_12500);
and U13339 (N_13339,N_12699,N_12691);
or U13340 (N_13340,N_13130,N_12423);
nor U13341 (N_13341,N_13143,N_12989);
or U13342 (N_13342,N_12995,N_12291);
and U13343 (N_13343,N_12253,N_12342);
xor U13344 (N_13344,N_13175,N_13009);
or U13345 (N_13345,N_12621,N_12705);
xor U13346 (N_13346,N_12741,N_12550);
xnor U13347 (N_13347,N_12090,N_13179);
nor U13348 (N_13348,N_12028,N_12626);
or U13349 (N_13349,N_12466,N_12100);
nor U13350 (N_13350,N_12968,N_12413);
nor U13351 (N_13351,N_13016,N_12567);
and U13352 (N_13352,N_13065,N_12484);
xnor U13353 (N_13353,N_13119,N_12682);
nand U13354 (N_13354,N_13127,N_12232);
nor U13355 (N_13355,N_12283,N_12787);
nand U13356 (N_13356,N_12314,N_12407);
nor U13357 (N_13357,N_13008,N_12401);
and U13358 (N_13358,N_13120,N_12604);
nand U13359 (N_13359,N_13037,N_12235);
xnor U13360 (N_13360,N_12529,N_12588);
xnor U13361 (N_13361,N_12139,N_12675);
nor U13362 (N_13362,N_12715,N_12752);
nand U13363 (N_13363,N_12753,N_12286);
nor U13364 (N_13364,N_12402,N_12475);
xnor U13365 (N_13365,N_12404,N_12898);
and U13366 (N_13366,N_13076,N_13072);
xor U13367 (N_13367,N_12942,N_13171);
nor U13368 (N_13368,N_12784,N_12866);
or U13369 (N_13369,N_12670,N_12482);
xor U13370 (N_13370,N_12765,N_12323);
and U13371 (N_13371,N_13139,N_12211);
and U13372 (N_13372,N_12432,N_12317);
and U13373 (N_13373,N_13041,N_12736);
xnor U13374 (N_13374,N_12547,N_12216);
nor U13375 (N_13375,N_13090,N_13117);
xnor U13376 (N_13376,N_12521,N_12881);
xnor U13377 (N_13377,N_13055,N_12591);
nor U13378 (N_13378,N_12062,N_12723);
nand U13379 (N_13379,N_12585,N_12516);
nor U13380 (N_13380,N_13093,N_12647);
nor U13381 (N_13381,N_12935,N_12779);
nor U13382 (N_13382,N_12243,N_12539);
xnor U13383 (N_13383,N_13088,N_12026);
nand U13384 (N_13384,N_12764,N_12650);
or U13385 (N_13385,N_12264,N_12932);
nand U13386 (N_13386,N_12353,N_12763);
and U13387 (N_13387,N_12583,N_12306);
nand U13388 (N_13388,N_12417,N_12114);
and U13389 (N_13389,N_12589,N_12640);
nand U13390 (N_13390,N_12042,N_12889);
nor U13391 (N_13391,N_12512,N_12176);
nand U13392 (N_13392,N_13102,N_13106);
xnor U13393 (N_13393,N_12955,N_12904);
or U13394 (N_13394,N_12436,N_12800);
xor U13395 (N_13395,N_12143,N_12566);
nand U13396 (N_13396,N_12440,N_12052);
or U13397 (N_13397,N_12558,N_12864);
xor U13398 (N_13398,N_12807,N_12277);
and U13399 (N_13399,N_12022,N_12377);
xor U13400 (N_13400,N_12701,N_12043);
and U13401 (N_13401,N_12592,N_12984);
nand U13402 (N_13402,N_13052,N_12136);
xnor U13403 (N_13403,N_13121,N_12593);
or U13404 (N_13404,N_12089,N_12419);
xnor U13405 (N_13405,N_12517,N_12160);
xnor U13406 (N_13406,N_12446,N_12275);
and U13407 (N_13407,N_12638,N_12065);
nand U13408 (N_13408,N_12281,N_12708);
nand U13409 (N_13409,N_12308,N_12454);
and U13410 (N_13410,N_12352,N_12803);
nand U13411 (N_13411,N_12101,N_12635);
or U13412 (N_13412,N_13186,N_12874);
and U13413 (N_13413,N_13075,N_12047);
or U13414 (N_13414,N_12532,N_12919);
nor U13415 (N_13415,N_12813,N_12941);
or U13416 (N_13416,N_12109,N_12471);
or U13417 (N_13417,N_12815,N_13169);
nand U13418 (N_13418,N_12262,N_12248);
nor U13419 (N_13419,N_12013,N_12814);
xnor U13420 (N_13420,N_12227,N_12721);
xnor U13421 (N_13421,N_12088,N_13000);
xor U13422 (N_13422,N_12840,N_12382);
or U13423 (N_13423,N_12718,N_12180);
nand U13424 (N_13424,N_12617,N_12769);
xnor U13425 (N_13425,N_12961,N_12978);
xor U13426 (N_13426,N_12622,N_12944);
xor U13427 (N_13427,N_13123,N_12590);
and U13428 (N_13428,N_12981,N_12152);
nor U13429 (N_13429,N_13151,N_12245);
or U13430 (N_13430,N_12213,N_12343);
nand U13431 (N_13431,N_12607,N_12605);
nand U13432 (N_13432,N_12234,N_12722);
xnor U13433 (N_13433,N_12613,N_12318);
and U13434 (N_13434,N_12606,N_13147);
nand U13435 (N_13435,N_12648,N_12249);
nor U13436 (N_13436,N_12937,N_12707);
and U13437 (N_13437,N_12231,N_12634);
nand U13438 (N_13438,N_12410,N_12744);
xor U13439 (N_13439,N_12018,N_12007);
nor U13440 (N_13440,N_12666,N_12742);
or U13441 (N_13441,N_12844,N_12597);
or U13442 (N_13442,N_12325,N_13155);
or U13443 (N_13443,N_12378,N_12444);
and U13444 (N_13444,N_12005,N_12392);
nand U13445 (N_13445,N_12877,N_12104);
xor U13446 (N_13446,N_12878,N_13190);
and U13447 (N_13447,N_13193,N_12327);
nand U13448 (N_13448,N_12381,N_12194);
or U13449 (N_13449,N_13031,N_12278);
nor U13450 (N_13450,N_12690,N_12319);
nor U13451 (N_13451,N_12203,N_12046);
xnor U13452 (N_13452,N_12188,N_12132);
nand U13453 (N_13453,N_12734,N_12655);
xor U13454 (N_13454,N_12762,N_13101);
xnor U13455 (N_13455,N_13015,N_12017);
nor U13456 (N_13456,N_13021,N_12582);
xnor U13457 (N_13457,N_12099,N_12633);
and U13458 (N_13458,N_12060,N_12999);
nor U13459 (N_13459,N_12930,N_12536);
nor U13460 (N_13460,N_12958,N_12954);
and U13461 (N_13461,N_12414,N_12857);
or U13462 (N_13462,N_12464,N_12196);
and U13463 (N_13463,N_12661,N_13136);
nand U13464 (N_13464,N_12385,N_12431);
and U13465 (N_13465,N_12596,N_12801);
nand U13466 (N_13466,N_12156,N_12170);
or U13467 (N_13467,N_12871,N_12894);
or U13468 (N_13468,N_12483,N_12365);
nor U13469 (N_13469,N_12002,N_12449);
and U13470 (N_13470,N_12333,N_12872);
nand U13471 (N_13471,N_12341,N_12581);
nand U13472 (N_13472,N_12486,N_12102);
xor U13473 (N_13473,N_12182,N_12681);
nand U13474 (N_13474,N_12573,N_12058);
or U13475 (N_13475,N_12882,N_13067);
xnor U13476 (N_13476,N_12397,N_12922);
and U13477 (N_13477,N_12673,N_12790);
nor U13478 (N_13478,N_13020,N_12795);
nor U13479 (N_13479,N_12662,N_12023);
or U13480 (N_13480,N_12491,N_13098);
nor U13481 (N_13481,N_12667,N_12294);
xor U13482 (N_13482,N_13131,N_12208);
xnor U13483 (N_13483,N_12791,N_12071);
or U13484 (N_13484,N_12972,N_12453);
nor U13485 (N_13485,N_12223,N_12636);
and U13486 (N_13486,N_12059,N_12504);
nor U13487 (N_13487,N_12773,N_13118);
nand U13488 (N_13488,N_12199,N_12015);
and U13489 (N_13489,N_12868,N_13050);
and U13490 (N_13490,N_12175,N_12950);
nor U13491 (N_13491,N_12201,N_12463);
or U13492 (N_13492,N_12094,N_12631);
nor U13493 (N_13493,N_12110,N_12405);
xor U13494 (N_13494,N_12739,N_13091);
and U13495 (N_13495,N_12144,N_12848);
and U13496 (N_13496,N_12757,N_13156);
nor U13497 (N_13497,N_12083,N_12918);
xnor U13498 (N_13498,N_12947,N_12997);
xor U13499 (N_13499,N_12311,N_12901);
nand U13500 (N_13500,N_12452,N_12629);
xor U13501 (N_13501,N_12971,N_12975);
nor U13502 (N_13502,N_12019,N_12735);
nand U13503 (N_13503,N_12489,N_12555);
xor U13504 (N_13504,N_12511,N_12165);
and U13505 (N_13505,N_12936,N_12103);
nand U13506 (N_13506,N_12962,N_13133);
or U13507 (N_13507,N_12082,N_12285);
or U13508 (N_13508,N_12967,N_12321);
nand U13509 (N_13509,N_12299,N_12117);
or U13510 (N_13510,N_12044,N_12251);
xor U13511 (N_13511,N_13138,N_13168);
nor U13512 (N_13512,N_12979,N_12912);
nor U13513 (N_13513,N_13182,N_12768);
nand U13514 (N_13514,N_12153,N_12448);
xor U13515 (N_13515,N_12421,N_12643);
nand U13516 (N_13516,N_12266,N_12789);
nor U13517 (N_13517,N_12724,N_12284);
xnor U13518 (N_13518,N_12347,N_12845);
nor U13519 (N_13519,N_12616,N_12081);
nor U13520 (N_13520,N_12649,N_12671);
and U13521 (N_13521,N_12468,N_12226);
and U13522 (N_13522,N_12400,N_12061);
nand U13523 (N_13523,N_12398,N_13087);
nor U13524 (N_13524,N_13030,N_12632);
xor U13525 (N_13525,N_12159,N_12664);
nor U13526 (N_13526,N_12376,N_12738);
nand U13527 (N_13527,N_12513,N_12481);
and U13528 (N_13528,N_12255,N_12442);
xor U13529 (N_13529,N_12982,N_13044);
nand U13530 (N_13530,N_12630,N_12838);
nor U13531 (N_13531,N_12372,N_12012);
nor U13532 (N_13532,N_12328,N_12187);
nand U13533 (N_13533,N_12862,N_12164);
or U13534 (N_13534,N_12653,N_12288);
nand U13535 (N_13535,N_12694,N_13107);
and U13536 (N_13536,N_12620,N_12469);
or U13537 (N_13537,N_12704,N_12776);
and U13538 (N_13538,N_13082,N_12174);
nand U13539 (N_13539,N_12786,N_13058);
nand U13540 (N_13540,N_12781,N_12087);
or U13541 (N_13541,N_13176,N_12435);
nand U13542 (N_13542,N_12125,N_13051);
xor U13543 (N_13543,N_12254,N_12568);
xnor U13544 (N_13544,N_12934,N_12369);
nand U13545 (N_13545,N_12966,N_12549);
or U13546 (N_13546,N_12824,N_12625);
and U13547 (N_13547,N_12375,N_12575);
nand U13548 (N_13548,N_12079,N_13174);
nand U13549 (N_13549,N_12326,N_12222);
and U13550 (N_13550,N_12867,N_12820);
nor U13551 (N_13551,N_12032,N_12805);
nand U13552 (N_13552,N_12485,N_12427);
nor U13553 (N_13553,N_12225,N_13199);
or U13554 (N_13554,N_12988,N_12420);
nand U13555 (N_13555,N_12070,N_12917);
or U13556 (N_13556,N_13111,N_13100);
and U13557 (N_13557,N_12905,N_12970);
or U13558 (N_13558,N_12080,N_12746);
nor U13559 (N_13559,N_12652,N_12296);
nand U13560 (N_13560,N_12391,N_12677);
and U13561 (N_13561,N_12259,N_13068);
xor U13562 (N_13562,N_13145,N_12146);
nand U13563 (N_13563,N_13039,N_12086);
xor U13564 (N_13564,N_12075,N_12915);
and U13565 (N_13565,N_12747,N_12931);
or U13566 (N_13566,N_12195,N_12335);
nand U13567 (N_13567,N_12137,N_13084);
xor U13568 (N_13568,N_12759,N_12880);
nor U13569 (N_13569,N_12717,N_12679);
or U13570 (N_13570,N_12772,N_12939);
nor U13571 (N_13571,N_12092,N_12498);
and U13572 (N_13572,N_12430,N_12379);
nand U13573 (N_13573,N_12533,N_13164);
or U13574 (N_13574,N_12644,N_12490);
xnor U13575 (N_13575,N_12068,N_12619);
or U13576 (N_13576,N_12368,N_12951);
and U13577 (N_13577,N_12804,N_12695);
or U13578 (N_13578,N_12337,N_12434);
or U13579 (N_13579,N_12134,N_12720);
and U13580 (N_13580,N_12716,N_12774);
and U13581 (N_13581,N_13024,N_12238);
and U13582 (N_13582,N_13077,N_12329);
xnor U13583 (N_13583,N_12272,N_12538);
or U13584 (N_13584,N_12150,N_12279);
and U13585 (N_13585,N_12310,N_12657);
nand U13586 (N_13586,N_12863,N_12854);
nand U13587 (N_13587,N_12645,N_12320);
or U13588 (N_13588,N_12554,N_12797);
and U13589 (N_13589,N_12236,N_12359);
and U13590 (N_13590,N_12370,N_12943);
nand U13591 (N_13591,N_12817,N_12010);
or U13592 (N_13592,N_12473,N_12856);
nor U13593 (N_13593,N_13063,N_12045);
or U13594 (N_13594,N_13047,N_12570);
and U13595 (N_13595,N_13064,N_12599);
and U13596 (N_13596,N_12771,N_12571);
and U13597 (N_13597,N_13004,N_12731);
nor U13598 (N_13598,N_12133,N_12713);
and U13599 (N_13599,N_12853,N_12172);
xor U13600 (N_13600,N_12252,N_12595);
and U13601 (N_13601,N_12031,N_12750);
nand U13602 (N_13602,N_12233,N_12025);
xor U13603 (N_13603,N_12908,N_12579);
nor U13604 (N_13604,N_13010,N_12526);
and U13605 (N_13605,N_12276,N_13013);
xnor U13606 (N_13606,N_12332,N_12883);
xor U13607 (N_13607,N_12287,N_12063);
nor U13608 (N_13608,N_12642,N_12230);
and U13609 (N_13609,N_12696,N_12293);
nand U13610 (N_13610,N_12522,N_12095);
and U13611 (N_13611,N_12663,N_12263);
xor U13612 (N_13612,N_12841,N_12561);
xor U13613 (N_13613,N_12760,N_12859);
nand U13614 (N_13614,N_12798,N_12860);
or U13615 (N_13615,N_12969,N_12130);
and U13616 (N_13616,N_13029,N_12748);
or U13617 (N_13617,N_12828,N_12001);
and U13618 (N_13618,N_12910,N_12183);
nand U13619 (N_13619,N_12220,N_12192);
xnor U13620 (N_13620,N_12145,N_12447);
and U13621 (N_13621,N_12618,N_12039);
and U13622 (N_13622,N_12363,N_12008);
and U13623 (N_13623,N_12141,N_12161);
nor U13624 (N_13624,N_12580,N_12437);
and U13625 (N_13625,N_13094,N_12135);
nand U13626 (N_13626,N_12895,N_13160);
xnor U13627 (N_13627,N_12569,N_12298);
and U13628 (N_13628,N_13019,N_12412);
and U13629 (N_13629,N_12993,N_12451);
xor U13630 (N_13630,N_12366,N_12974);
and U13631 (N_13631,N_12602,N_12097);
nand U13632 (N_13632,N_12885,N_12706);
and U13633 (N_13633,N_12115,N_12506);
and U13634 (N_13634,N_12641,N_12959);
or U13635 (N_13635,N_12433,N_12710);
nor U13636 (N_13636,N_12355,N_12051);
nand U13637 (N_13637,N_12948,N_12921);
nand U13638 (N_13638,N_12054,N_13178);
nand U13639 (N_13639,N_13132,N_13023);
nand U13640 (N_13640,N_12038,N_12892);
xor U13641 (N_13641,N_12390,N_13129);
and U13642 (N_13642,N_12755,N_12835);
nor U13643 (N_13643,N_13103,N_12207);
nor U13644 (N_13644,N_12615,N_12098);
nand U13645 (N_13645,N_12887,N_12205);
nand U13646 (N_13646,N_13092,N_12173);
and U13647 (N_13647,N_12855,N_12445);
nand U13648 (N_13648,N_12184,N_12827);
nor U13649 (N_13649,N_12000,N_12810);
nand U13650 (N_13650,N_13185,N_12940);
xnor U13651 (N_13651,N_12780,N_12169);
and U13652 (N_13652,N_12282,N_12998);
nor U13653 (N_13653,N_13183,N_13113);
xnor U13654 (N_13654,N_12218,N_12890);
nand U13655 (N_13655,N_12510,N_12672);
nand U13656 (N_13656,N_12587,N_12315);
or U13657 (N_13657,N_12945,N_12990);
xor U13658 (N_13658,N_12191,N_12040);
nand U13659 (N_13659,N_12964,N_12108);
or U13660 (N_13660,N_12024,N_12770);
or U13661 (N_13661,N_12562,N_12426);
xor U13662 (N_13662,N_13049,N_12190);
nand U13663 (N_13663,N_12792,N_12345);
xnor U13664 (N_13664,N_13086,N_12351);
nand U13665 (N_13665,N_12106,N_13192);
xnor U13666 (N_13666,N_12425,N_12808);
nand U13667 (N_13667,N_13194,N_12292);
and U13668 (N_13668,N_13150,N_13112);
nor U13669 (N_13669,N_12782,N_13038);
nand U13670 (N_13670,N_12837,N_12198);
nand U13671 (N_13671,N_12923,N_12214);
xor U13672 (N_13672,N_12396,N_12111);
or U13673 (N_13673,N_12209,N_12541);
nor U13674 (N_13674,N_13079,N_12842);
and U13675 (N_13675,N_12711,N_12823);
and U13676 (N_13676,N_12364,N_12584);
nor U13677 (N_13677,N_12600,N_12911);
nand U13678 (N_13678,N_12507,N_12066);
nor U13679 (N_13679,N_12416,N_13189);
or U13680 (N_13680,N_12472,N_13134);
nor U13681 (N_13681,N_12105,N_12793);
and U13682 (N_13682,N_12107,N_12545);
xor U13683 (N_13683,N_13054,N_12669);
xnor U13684 (N_13684,N_13158,N_12965);
xnor U13685 (N_13685,N_13012,N_12151);
or U13686 (N_13686,N_12331,N_12443);
and U13687 (N_13687,N_12334,N_12096);
and U13688 (N_13688,N_12179,N_12009);
xor U13689 (N_13689,N_12534,N_12021);
xnor U13690 (N_13690,N_12034,N_12873);
nand U13691 (N_13691,N_12687,N_12346);
or U13692 (N_13692,N_12574,N_12269);
xnor U13693 (N_13693,N_13140,N_12167);
nand U13694 (N_13694,N_12819,N_13197);
xor U13695 (N_13695,N_12217,N_13181);
nand U13696 (N_13696,N_12985,N_12858);
nor U13697 (N_13697,N_13163,N_12177);
xnor U13698 (N_13698,N_12116,N_12830);
and U13699 (N_13699,N_12656,N_13116);
or U13700 (N_13700,N_12952,N_13022);
and U13701 (N_13701,N_12727,N_12806);
xnor U13702 (N_13702,N_12127,N_12181);
or U13703 (N_13703,N_12730,N_12121);
nor U13704 (N_13704,N_12703,N_12429);
xor U13705 (N_13705,N_12654,N_12869);
or U13706 (N_13706,N_13105,N_12193);
nand U13707 (N_13707,N_12783,N_12693);
or U13708 (N_13708,N_12977,N_13165);
and U13709 (N_13709,N_12737,N_12495);
or U13710 (N_13710,N_13196,N_12551);
xnor U13711 (N_13711,N_12639,N_13137);
nand U13712 (N_13712,N_12812,N_12577);
and U13713 (N_13713,N_12986,N_12064);
xnor U13714 (N_13714,N_13017,N_12124);
xor U13715 (N_13715,N_12126,N_12702);
nor U13716 (N_13716,N_12851,N_12348);
nor U13717 (N_13717,N_13195,N_12624);
nand U13718 (N_13718,N_12091,N_12384);
or U13719 (N_13719,N_13187,N_13153);
xor U13720 (N_13720,N_12076,N_12623);
xnor U13721 (N_13721,N_13146,N_12330);
or U13722 (N_13722,N_12896,N_12350);
xnor U13723 (N_13723,N_12523,N_12258);
nand U13724 (N_13724,N_12268,N_12305);
nor U13725 (N_13725,N_12265,N_12037);
or U13726 (N_13726,N_12909,N_12888);
nand U13727 (N_13727,N_12886,N_12289);
nand U13728 (N_13728,N_12004,N_12492);
nor U13729 (N_13729,N_12403,N_12926);
and U13730 (N_13730,N_12994,N_12307);
nor U13731 (N_13731,N_12215,N_12559);
and U13732 (N_13732,N_12239,N_12897);
and U13733 (N_13733,N_12938,N_12611);
nand U13734 (N_13734,N_12354,N_13114);
xnor U13735 (N_13735,N_12751,N_12540);
nor U13736 (N_13736,N_12528,N_13095);
nand U13737 (N_13737,N_12186,N_12455);
nor U13738 (N_13738,N_12460,N_12543);
nor U13739 (N_13739,N_12927,N_13034);
or U13740 (N_13740,N_12794,N_12131);
nor U13741 (N_13741,N_12719,N_12221);
xnor U13742 (N_13742,N_13036,N_13026);
nand U13743 (N_13743,N_12149,N_12907);
nor U13744 (N_13744,N_12700,N_13070);
nand U13745 (N_13745,N_12709,N_12683);
or U13746 (N_13746,N_12185,N_13115);
xor U13747 (N_13747,N_12450,N_13099);
or U13748 (N_13748,N_12297,N_13148);
nor U13749 (N_13749,N_12527,N_12913);
xor U13750 (N_13750,N_12057,N_12409);
or U13751 (N_13751,N_12849,N_12371);
or U13752 (N_13752,N_12050,N_12077);
and U13753 (N_13753,N_12356,N_13007);
xnor U13754 (N_13754,N_12155,N_12461);
nand U13755 (N_13755,N_12303,N_13173);
nand U13756 (N_13756,N_12336,N_12339);
nand U13757 (N_13757,N_12740,N_12027);
nand U13758 (N_13758,N_12586,N_13085);
xnor U13759 (N_13759,N_12393,N_12212);
or U13760 (N_13760,N_12627,N_13080);
nand U13761 (N_13761,N_12178,N_12903);
or U13762 (N_13762,N_12833,N_12557);
nor U13763 (N_13763,N_12138,N_12608);
nor U13764 (N_13764,N_12118,N_12493);
and U13765 (N_13765,N_13128,N_12011);
xor U13766 (N_13766,N_12415,N_12204);
nor U13767 (N_13767,N_13122,N_12479);
nand U13768 (N_13768,N_12441,N_12775);
nor U13769 (N_13769,N_12358,N_12142);
and U13770 (N_13770,N_12685,N_12548);
or U13771 (N_13771,N_12665,N_12422);
nor U13772 (N_13772,N_13184,N_13035);
nor U13773 (N_13773,N_12530,N_12552);
nand U13774 (N_13774,N_12459,N_12758);
nand U13775 (N_13775,N_12313,N_12147);
nand U13776 (N_13776,N_12933,N_12578);
nand U13777 (N_13777,N_13043,N_12668);
or U13778 (N_13778,N_12154,N_12344);
and U13779 (N_13779,N_12834,N_12925);
nand U13780 (N_13780,N_12361,N_13040);
or U13781 (N_13781,N_12312,N_13011);
or U13782 (N_13782,N_12929,N_12267);
xnor U13783 (N_13783,N_12270,N_12870);
xor U13784 (N_13784,N_12920,N_12362);
nor U13785 (N_13785,N_13157,N_12899);
and U13786 (N_13786,N_12424,N_12754);
or U13787 (N_13787,N_12983,N_12302);
and U13788 (N_13788,N_12519,N_12120);
xor U13789 (N_13789,N_12726,N_12546);
nand U13790 (N_13790,N_12802,N_13188);
xor U13791 (N_13791,N_13198,N_12831);
or U13792 (N_13792,N_12497,N_12162);
nor U13793 (N_13793,N_12113,N_12825);
xnor U13794 (N_13794,N_12085,N_12991);
and U13795 (N_13795,N_12601,N_12157);
nor U13796 (N_13796,N_12850,N_12865);
xor U13797 (N_13797,N_12745,N_12148);
or U13798 (N_13798,N_12041,N_12477);
xor U13799 (N_13799,N_12029,N_13057);
nand U13800 (N_13800,N_13190,N_12827);
nand U13801 (N_13801,N_12357,N_12514);
or U13802 (N_13802,N_12776,N_12675);
xnor U13803 (N_13803,N_12974,N_12878);
nor U13804 (N_13804,N_13028,N_12989);
or U13805 (N_13805,N_12123,N_12652);
nor U13806 (N_13806,N_12421,N_12192);
or U13807 (N_13807,N_12289,N_12421);
nand U13808 (N_13808,N_12823,N_12480);
or U13809 (N_13809,N_12173,N_12056);
and U13810 (N_13810,N_12570,N_12036);
nand U13811 (N_13811,N_12938,N_12812);
or U13812 (N_13812,N_12870,N_12063);
and U13813 (N_13813,N_13071,N_13198);
nor U13814 (N_13814,N_12062,N_12884);
and U13815 (N_13815,N_13153,N_13017);
nor U13816 (N_13816,N_12576,N_12910);
nand U13817 (N_13817,N_13114,N_12607);
nor U13818 (N_13818,N_12241,N_12313);
nand U13819 (N_13819,N_12453,N_12694);
or U13820 (N_13820,N_13112,N_12077);
or U13821 (N_13821,N_13043,N_12969);
nand U13822 (N_13822,N_12235,N_12015);
or U13823 (N_13823,N_12652,N_12129);
and U13824 (N_13824,N_12113,N_12227);
nand U13825 (N_13825,N_13090,N_12096);
or U13826 (N_13826,N_12525,N_12695);
nand U13827 (N_13827,N_12417,N_12884);
or U13828 (N_13828,N_12627,N_12054);
and U13829 (N_13829,N_13199,N_13151);
and U13830 (N_13830,N_13028,N_13183);
or U13831 (N_13831,N_12487,N_12709);
and U13832 (N_13832,N_12980,N_12765);
and U13833 (N_13833,N_13066,N_13027);
xnor U13834 (N_13834,N_12493,N_12470);
and U13835 (N_13835,N_12459,N_12356);
and U13836 (N_13836,N_12381,N_12587);
xnor U13837 (N_13837,N_12395,N_12454);
and U13838 (N_13838,N_12404,N_13009);
nand U13839 (N_13839,N_12417,N_12201);
and U13840 (N_13840,N_12736,N_12978);
xor U13841 (N_13841,N_12579,N_12586);
xnor U13842 (N_13842,N_12287,N_12174);
nor U13843 (N_13843,N_12765,N_12518);
or U13844 (N_13844,N_12250,N_12442);
xor U13845 (N_13845,N_12512,N_12934);
or U13846 (N_13846,N_12786,N_12419);
nor U13847 (N_13847,N_12276,N_12988);
nor U13848 (N_13848,N_12847,N_12051);
or U13849 (N_13849,N_12186,N_12913);
or U13850 (N_13850,N_12098,N_12535);
and U13851 (N_13851,N_12512,N_12769);
nor U13852 (N_13852,N_12635,N_12410);
or U13853 (N_13853,N_12506,N_12800);
nor U13854 (N_13854,N_12099,N_13081);
nor U13855 (N_13855,N_13045,N_12517);
or U13856 (N_13856,N_12543,N_12820);
or U13857 (N_13857,N_12778,N_13038);
and U13858 (N_13858,N_13006,N_12304);
xnor U13859 (N_13859,N_12301,N_12981);
and U13860 (N_13860,N_12394,N_12519);
xor U13861 (N_13861,N_12913,N_13079);
or U13862 (N_13862,N_12770,N_12487);
and U13863 (N_13863,N_12735,N_12421);
nor U13864 (N_13864,N_13070,N_12396);
or U13865 (N_13865,N_12373,N_12237);
and U13866 (N_13866,N_12643,N_12063);
nor U13867 (N_13867,N_12035,N_12721);
xnor U13868 (N_13868,N_12481,N_12696);
and U13869 (N_13869,N_12381,N_12148);
xnor U13870 (N_13870,N_12255,N_12365);
xor U13871 (N_13871,N_12906,N_12670);
nor U13872 (N_13872,N_12745,N_12790);
xor U13873 (N_13873,N_12238,N_12105);
and U13874 (N_13874,N_12541,N_12184);
or U13875 (N_13875,N_12143,N_12684);
nor U13876 (N_13876,N_12272,N_12172);
nand U13877 (N_13877,N_12727,N_12359);
and U13878 (N_13878,N_13193,N_12091);
and U13879 (N_13879,N_12340,N_12184);
nand U13880 (N_13880,N_12714,N_13000);
or U13881 (N_13881,N_13098,N_13124);
or U13882 (N_13882,N_12801,N_13164);
or U13883 (N_13883,N_12955,N_12634);
xor U13884 (N_13884,N_12992,N_12003);
nor U13885 (N_13885,N_12062,N_12840);
nand U13886 (N_13886,N_12365,N_12942);
and U13887 (N_13887,N_13157,N_12153);
or U13888 (N_13888,N_12358,N_12168);
or U13889 (N_13889,N_12561,N_12153);
nand U13890 (N_13890,N_12375,N_12675);
or U13891 (N_13891,N_13129,N_12029);
nor U13892 (N_13892,N_12882,N_13187);
nor U13893 (N_13893,N_13090,N_12465);
nand U13894 (N_13894,N_12518,N_12845);
xnor U13895 (N_13895,N_12875,N_13074);
nor U13896 (N_13896,N_12209,N_12339);
or U13897 (N_13897,N_12316,N_12199);
xor U13898 (N_13898,N_12698,N_13162);
nand U13899 (N_13899,N_12197,N_12740);
and U13900 (N_13900,N_13031,N_12806);
or U13901 (N_13901,N_12418,N_12085);
nor U13902 (N_13902,N_12664,N_12443);
and U13903 (N_13903,N_12940,N_12512);
nor U13904 (N_13904,N_12823,N_12991);
or U13905 (N_13905,N_12461,N_12905);
nand U13906 (N_13906,N_13001,N_12170);
nand U13907 (N_13907,N_12422,N_12815);
or U13908 (N_13908,N_12525,N_12171);
nand U13909 (N_13909,N_12053,N_12548);
nand U13910 (N_13910,N_12292,N_12985);
nand U13911 (N_13911,N_13179,N_12701);
and U13912 (N_13912,N_12894,N_13112);
nor U13913 (N_13913,N_12680,N_12070);
and U13914 (N_13914,N_12268,N_12272);
nor U13915 (N_13915,N_12861,N_12772);
or U13916 (N_13916,N_12023,N_12081);
or U13917 (N_13917,N_12110,N_12303);
nor U13918 (N_13918,N_12698,N_12798);
nand U13919 (N_13919,N_12336,N_13072);
or U13920 (N_13920,N_12266,N_12384);
xnor U13921 (N_13921,N_13033,N_13030);
nand U13922 (N_13922,N_13163,N_12282);
xnor U13923 (N_13923,N_12617,N_12228);
or U13924 (N_13924,N_12405,N_12013);
and U13925 (N_13925,N_12371,N_12770);
and U13926 (N_13926,N_12884,N_12086);
or U13927 (N_13927,N_12094,N_12535);
xor U13928 (N_13928,N_12526,N_12325);
or U13929 (N_13929,N_12398,N_13126);
nand U13930 (N_13930,N_13119,N_12587);
and U13931 (N_13931,N_13115,N_12434);
nand U13932 (N_13932,N_12564,N_12551);
nor U13933 (N_13933,N_12004,N_12203);
or U13934 (N_13934,N_12622,N_12461);
or U13935 (N_13935,N_12088,N_12941);
nor U13936 (N_13936,N_12727,N_12579);
xor U13937 (N_13937,N_12243,N_12769);
xnor U13938 (N_13938,N_12947,N_12108);
nor U13939 (N_13939,N_12221,N_12173);
and U13940 (N_13940,N_12800,N_12533);
nand U13941 (N_13941,N_12342,N_12475);
xor U13942 (N_13942,N_12984,N_12275);
xor U13943 (N_13943,N_13153,N_12743);
xor U13944 (N_13944,N_12898,N_12243);
xor U13945 (N_13945,N_12023,N_12939);
xnor U13946 (N_13946,N_12562,N_12376);
xor U13947 (N_13947,N_12594,N_12936);
and U13948 (N_13948,N_12149,N_12595);
and U13949 (N_13949,N_12586,N_13165);
or U13950 (N_13950,N_13155,N_12166);
and U13951 (N_13951,N_12069,N_12971);
xor U13952 (N_13952,N_12584,N_12665);
or U13953 (N_13953,N_13196,N_12835);
and U13954 (N_13954,N_12848,N_12324);
and U13955 (N_13955,N_12654,N_12477);
and U13956 (N_13956,N_13141,N_12289);
or U13957 (N_13957,N_13037,N_12507);
or U13958 (N_13958,N_12543,N_13006);
nor U13959 (N_13959,N_12132,N_12230);
xor U13960 (N_13960,N_12663,N_12894);
nor U13961 (N_13961,N_12768,N_12444);
and U13962 (N_13962,N_12165,N_13186);
and U13963 (N_13963,N_12306,N_12410);
xor U13964 (N_13964,N_12551,N_12607);
xor U13965 (N_13965,N_12032,N_12408);
nor U13966 (N_13966,N_13078,N_13092);
nand U13967 (N_13967,N_13194,N_12497);
and U13968 (N_13968,N_12730,N_12137);
xor U13969 (N_13969,N_12233,N_12344);
nand U13970 (N_13970,N_12937,N_13132);
nor U13971 (N_13971,N_13108,N_12337);
nor U13972 (N_13972,N_12230,N_12122);
nand U13973 (N_13973,N_12447,N_12942);
nor U13974 (N_13974,N_12838,N_13131);
nand U13975 (N_13975,N_12679,N_13019);
nor U13976 (N_13976,N_12372,N_12468);
xor U13977 (N_13977,N_12456,N_13150);
nand U13978 (N_13978,N_12949,N_12085);
nand U13979 (N_13979,N_12288,N_13143);
or U13980 (N_13980,N_12982,N_12251);
xor U13981 (N_13981,N_12762,N_12664);
nand U13982 (N_13982,N_12174,N_12437);
nor U13983 (N_13983,N_12204,N_12319);
nand U13984 (N_13984,N_12475,N_12457);
nor U13985 (N_13985,N_12172,N_12781);
nand U13986 (N_13986,N_12627,N_12921);
or U13987 (N_13987,N_12716,N_13090);
or U13988 (N_13988,N_12639,N_12221);
xnor U13989 (N_13989,N_12701,N_12310);
and U13990 (N_13990,N_13161,N_12119);
nor U13991 (N_13991,N_12138,N_13171);
nor U13992 (N_13992,N_12512,N_12529);
and U13993 (N_13993,N_12487,N_12499);
and U13994 (N_13994,N_12553,N_13000);
xor U13995 (N_13995,N_12344,N_12921);
xnor U13996 (N_13996,N_12074,N_12807);
nor U13997 (N_13997,N_12727,N_13052);
and U13998 (N_13998,N_13101,N_12444);
nand U13999 (N_13999,N_12802,N_12236);
and U14000 (N_14000,N_12601,N_12559);
nor U14001 (N_14001,N_12048,N_12103);
nor U14002 (N_14002,N_12133,N_12361);
xnor U14003 (N_14003,N_13112,N_12952);
xnor U14004 (N_14004,N_12532,N_12859);
nand U14005 (N_14005,N_12833,N_13002);
or U14006 (N_14006,N_12035,N_12927);
nand U14007 (N_14007,N_12781,N_12911);
or U14008 (N_14008,N_13039,N_12179);
nor U14009 (N_14009,N_12699,N_13156);
xor U14010 (N_14010,N_12327,N_12790);
and U14011 (N_14011,N_12276,N_12531);
xnor U14012 (N_14012,N_12937,N_12725);
nand U14013 (N_14013,N_13004,N_12311);
and U14014 (N_14014,N_12016,N_12288);
nor U14015 (N_14015,N_12729,N_12882);
nand U14016 (N_14016,N_12537,N_12005);
nand U14017 (N_14017,N_12964,N_12257);
xnor U14018 (N_14018,N_12248,N_13112);
xor U14019 (N_14019,N_12984,N_12530);
or U14020 (N_14020,N_13177,N_12932);
nor U14021 (N_14021,N_12546,N_13164);
nor U14022 (N_14022,N_12488,N_13189);
nand U14023 (N_14023,N_12087,N_12551);
xor U14024 (N_14024,N_12239,N_12021);
or U14025 (N_14025,N_12191,N_12764);
or U14026 (N_14026,N_12444,N_12991);
nand U14027 (N_14027,N_12759,N_12215);
or U14028 (N_14028,N_12774,N_12075);
nor U14029 (N_14029,N_12681,N_12979);
nand U14030 (N_14030,N_13102,N_13143);
xnor U14031 (N_14031,N_12761,N_12959);
xnor U14032 (N_14032,N_13126,N_13103);
and U14033 (N_14033,N_12514,N_12898);
nor U14034 (N_14034,N_12369,N_12585);
and U14035 (N_14035,N_12675,N_12650);
nor U14036 (N_14036,N_12682,N_13105);
xnor U14037 (N_14037,N_12618,N_12621);
and U14038 (N_14038,N_12155,N_12615);
or U14039 (N_14039,N_12833,N_12839);
or U14040 (N_14040,N_12419,N_12307);
xor U14041 (N_14041,N_13003,N_12840);
nand U14042 (N_14042,N_13037,N_12349);
and U14043 (N_14043,N_13049,N_12069);
nand U14044 (N_14044,N_13082,N_12419);
nor U14045 (N_14045,N_12552,N_12064);
xor U14046 (N_14046,N_12685,N_12862);
and U14047 (N_14047,N_12722,N_12329);
xor U14048 (N_14048,N_12658,N_13047);
and U14049 (N_14049,N_13049,N_12684);
nand U14050 (N_14050,N_12758,N_12552);
or U14051 (N_14051,N_12566,N_12024);
xor U14052 (N_14052,N_12393,N_12737);
nand U14053 (N_14053,N_12546,N_12450);
xnor U14054 (N_14054,N_12414,N_12671);
nand U14055 (N_14055,N_12886,N_12086);
nand U14056 (N_14056,N_12241,N_12454);
nor U14057 (N_14057,N_13181,N_13042);
nor U14058 (N_14058,N_12581,N_12478);
nand U14059 (N_14059,N_13133,N_12723);
nand U14060 (N_14060,N_12418,N_13019);
xnor U14061 (N_14061,N_12891,N_12311);
xnor U14062 (N_14062,N_12193,N_12125);
nand U14063 (N_14063,N_13074,N_13090);
nor U14064 (N_14064,N_12063,N_12640);
nand U14065 (N_14065,N_12665,N_12171);
nand U14066 (N_14066,N_12458,N_13130);
and U14067 (N_14067,N_12057,N_12323);
and U14068 (N_14068,N_12283,N_12323);
or U14069 (N_14069,N_12744,N_12168);
xor U14070 (N_14070,N_12785,N_12268);
or U14071 (N_14071,N_12906,N_12507);
nor U14072 (N_14072,N_13110,N_12870);
nand U14073 (N_14073,N_12881,N_12055);
and U14074 (N_14074,N_12598,N_12745);
or U14075 (N_14075,N_12886,N_13177);
or U14076 (N_14076,N_13185,N_12374);
nand U14077 (N_14077,N_13041,N_12571);
nor U14078 (N_14078,N_12997,N_12611);
and U14079 (N_14079,N_12159,N_13196);
and U14080 (N_14080,N_12554,N_12104);
xnor U14081 (N_14081,N_13024,N_12726);
xor U14082 (N_14082,N_12755,N_12055);
or U14083 (N_14083,N_12400,N_12623);
nor U14084 (N_14084,N_12228,N_13146);
nor U14085 (N_14085,N_12567,N_12351);
xnor U14086 (N_14086,N_13179,N_12502);
or U14087 (N_14087,N_12172,N_13174);
nand U14088 (N_14088,N_12396,N_12067);
or U14089 (N_14089,N_12431,N_12056);
nand U14090 (N_14090,N_12260,N_13174);
and U14091 (N_14091,N_12141,N_12520);
and U14092 (N_14092,N_12927,N_12392);
nand U14093 (N_14093,N_12794,N_12888);
nand U14094 (N_14094,N_12667,N_13147);
nor U14095 (N_14095,N_13139,N_12518);
and U14096 (N_14096,N_13123,N_12613);
xor U14097 (N_14097,N_12892,N_13133);
and U14098 (N_14098,N_12509,N_13184);
nand U14099 (N_14099,N_12581,N_13163);
or U14100 (N_14100,N_13005,N_12543);
or U14101 (N_14101,N_12223,N_12824);
nor U14102 (N_14102,N_13123,N_12683);
nor U14103 (N_14103,N_12941,N_12763);
and U14104 (N_14104,N_12628,N_13028);
or U14105 (N_14105,N_12994,N_12541);
nor U14106 (N_14106,N_12916,N_12906);
nand U14107 (N_14107,N_12570,N_12630);
xnor U14108 (N_14108,N_12913,N_12492);
nor U14109 (N_14109,N_12176,N_12302);
and U14110 (N_14110,N_12059,N_12149);
nor U14111 (N_14111,N_13114,N_12651);
xor U14112 (N_14112,N_12945,N_12201);
or U14113 (N_14113,N_12345,N_12404);
and U14114 (N_14114,N_12265,N_12710);
nor U14115 (N_14115,N_12861,N_13120);
xor U14116 (N_14116,N_13101,N_13138);
nor U14117 (N_14117,N_12366,N_12764);
nand U14118 (N_14118,N_12937,N_12221);
nor U14119 (N_14119,N_12695,N_13007);
nand U14120 (N_14120,N_12425,N_12475);
or U14121 (N_14121,N_12660,N_13065);
xnor U14122 (N_14122,N_13075,N_12888);
nor U14123 (N_14123,N_12077,N_12467);
xnor U14124 (N_14124,N_12734,N_13097);
xnor U14125 (N_14125,N_12133,N_13088);
nand U14126 (N_14126,N_12705,N_13079);
xnor U14127 (N_14127,N_12209,N_12438);
or U14128 (N_14128,N_12690,N_13109);
nor U14129 (N_14129,N_12489,N_12870);
xnor U14130 (N_14130,N_12491,N_12240);
xnor U14131 (N_14131,N_13179,N_12533);
xnor U14132 (N_14132,N_12735,N_12750);
nand U14133 (N_14133,N_12124,N_12047);
xnor U14134 (N_14134,N_12344,N_13107);
and U14135 (N_14135,N_12789,N_12759);
xor U14136 (N_14136,N_12333,N_12881);
or U14137 (N_14137,N_12545,N_12212);
xnor U14138 (N_14138,N_12533,N_12400);
xor U14139 (N_14139,N_12130,N_12424);
or U14140 (N_14140,N_12534,N_12423);
or U14141 (N_14141,N_12906,N_12883);
nand U14142 (N_14142,N_12557,N_12702);
xnor U14143 (N_14143,N_12692,N_12971);
xor U14144 (N_14144,N_12471,N_12207);
xnor U14145 (N_14145,N_12485,N_12030);
nor U14146 (N_14146,N_12378,N_12296);
and U14147 (N_14147,N_12932,N_12018);
nor U14148 (N_14148,N_12988,N_12695);
nand U14149 (N_14149,N_12010,N_12180);
nor U14150 (N_14150,N_12217,N_12541);
xnor U14151 (N_14151,N_12429,N_13068);
xnor U14152 (N_14152,N_12797,N_12096);
nand U14153 (N_14153,N_12425,N_12703);
xnor U14154 (N_14154,N_12643,N_12342);
or U14155 (N_14155,N_12122,N_12633);
and U14156 (N_14156,N_12075,N_12090);
xnor U14157 (N_14157,N_13136,N_12448);
xor U14158 (N_14158,N_12755,N_13197);
nor U14159 (N_14159,N_12618,N_13089);
xnor U14160 (N_14160,N_12428,N_12224);
nor U14161 (N_14161,N_12452,N_12478);
nand U14162 (N_14162,N_12743,N_12927);
and U14163 (N_14163,N_12105,N_12858);
or U14164 (N_14164,N_12159,N_12991);
and U14165 (N_14165,N_12803,N_12655);
and U14166 (N_14166,N_12522,N_12405);
xor U14167 (N_14167,N_12373,N_13128);
or U14168 (N_14168,N_13010,N_12656);
nand U14169 (N_14169,N_12305,N_12952);
nor U14170 (N_14170,N_12089,N_12360);
or U14171 (N_14171,N_12742,N_13151);
or U14172 (N_14172,N_12728,N_12262);
and U14173 (N_14173,N_12593,N_12292);
nor U14174 (N_14174,N_12176,N_12149);
xor U14175 (N_14175,N_12819,N_13059);
nor U14176 (N_14176,N_12972,N_12495);
xor U14177 (N_14177,N_12704,N_12458);
and U14178 (N_14178,N_13029,N_12863);
nor U14179 (N_14179,N_13047,N_12971);
xor U14180 (N_14180,N_12740,N_13105);
nor U14181 (N_14181,N_12998,N_13041);
or U14182 (N_14182,N_12983,N_12519);
nor U14183 (N_14183,N_13025,N_12944);
nand U14184 (N_14184,N_12140,N_12194);
nand U14185 (N_14185,N_12281,N_12851);
nor U14186 (N_14186,N_12812,N_12400);
nor U14187 (N_14187,N_12451,N_12559);
or U14188 (N_14188,N_12125,N_12605);
nor U14189 (N_14189,N_13032,N_12615);
and U14190 (N_14190,N_12450,N_12097);
and U14191 (N_14191,N_12106,N_13017);
or U14192 (N_14192,N_12173,N_13015);
xnor U14193 (N_14193,N_13025,N_12188);
and U14194 (N_14194,N_12962,N_12285);
xnor U14195 (N_14195,N_12496,N_12102);
nor U14196 (N_14196,N_13136,N_12033);
nor U14197 (N_14197,N_12887,N_12244);
xor U14198 (N_14198,N_13123,N_12549);
or U14199 (N_14199,N_12259,N_12795);
nand U14200 (N_14200,N_12518,N_12854);
xor U14201 (N_14201,N_12016,N_12568);
nand U14202 (N_14202,N_12870,N_12268);
nand U14203 (N_14203,N_12405,N_12544);
and U14204 (N_14204,N_12751,N_12591);
or U14205 (N_14205,N_12278,N_12219);
nor U14206 (N_14206,N_12248,N_12107);
nor U14207 (N_14207,N_12546,N_12129);
nand U14208 (N_14208,N_12421,N_12096);
and U14209 (N_14209,N_13198,N_13082);
or U14210 (N_14210,N_12563,N_12529);
nor U14211 (N_14211,N_12822,N_13026);
or U14212 (N_14212,N_12557,N_12171);
and U14213 (N_14213,N_12697,N_13123);
nand U14214 (N_14214,N_12212,N_12927);
nor U14215 (N_14215,N_13082,N_13181);
and U14216 (N_14216,N_12370,N_12619);
and U14217 (N_14217,N_13081,N_12855);
and U14218 (N_14218,N_12663,N_12122);
or U14219 (N_14219,N_12200,N_12668);
nand U14220 (N_14220,N_12273,N_12163);
nor U14221 (N_14221,N_12090,N_13181);
xor U14222 (N_14222,N_12995,N_12768);
nor U14223 (N_14223,N_12577,N_12660);
nand U14224 (N_14224,N_12721,N_12645);
nor U14225 (N_14225,N_12938,N_13167);
nor U14226 (N_14226,N_12134,N_12806);
nand U14227 (N_14227,N_13194,N_12520);
xnor U14228 (N_14228,N_13110,N_12129);
or U14229 (N_14229,N_12429,N_12005);
nor U14230 (N_14230,N_12518,N_12701);
nor U14231 (N_14231,N_13049,N_12575);
or U14232 (N_14232,N_13167,N_12481);
nor U14233 (N_14233,N_13117,N_12004);
or U14234 (N_14234,N_12881,N_12291);
xnor U14235 (N_14235,N_12926,N_12832);
nand U14236 (N_14236,N_12614,N_12981);
and U14237 (N_14237,N_12467,N_12746);
xor U14238 (N_14238,N_12766,N_12448);
nand U14239 (N_14239,N_12394,N_12645);
nor U14240 (N_14240,N_12847,N_13150);
nor U14241 (N_14241,N_12804,N_12161);
nor U14242 (N_14242,N_12499,N_13101);
xnor U14243 (N_14243,N_12211,N_12026);
nand U14244 (N_14244,N_12991,N_12245);
and U14245 (N_14245,N_13168,N_12399);
or U14246 (N_14246,N_12187,N_12246);
nor U14247 (N_14247,N_12834,N_13104);
and U14248 (N_14248,N_12892,N_12979);
nor U14249 (N_14249,N_12866,N_12125);
and U14250 (N_14250,N_12962,N_12268);
or U14251 (N_14251,N_12715,N_12981);
or U14252 (N_14252,N_12996,N_13114);
and U14253 (N_14253,N_12423,N_12629);
nand U14254 (N_14254,N_12587,N_12648);
or U14255 (N_14255,N_12712,N_12941);
and U14256 (N_14256,N_12413,N_12470);
and U14257 (N_14257,N_13126,N_12819);
and U14258 (N_14258,N_13044,N_12560);
xor U14259 (N_14259,N_12103,N_12090);
nor U14260 (N_14260,N_12680,N_12223);
and U14261 (N_14261,N_12230,N_12278);
or U14262 (N_14262,N_12808,N_12020);
or U14263 (N_14263,N_12416,N_13053);
or U14264 (N_14264,N_12561,N_12910);
and U14265 (N_14265,N_13125,N_12635);
nor U14266 (N_14266,N_13010,N_12930);
or U14267 (N_14267,N_12641,N_12973);
nand U14268 (N_14268,N_13054,N_12214);
or U14269 (N_14269,N_12555,N_12209);
nand U14270 (N_14270,N_12912,N_12412);
or U14271 (N_14271,N_12737,N_12415);
xor U14272 (N_14272,N_12909,N_12179);
xnor U14273 (N_14273,N_12572,N_12681);
or U14274 (N_14274,N_12686,N_12184);
nand U14275 (N_14275,N_13001,N_12895);
xor U14276 (N_14276,N_12926,N_12955);
and U14277 (N_14277,N_12366,N_12915);
xnor U14278 (N_14278,N_12649,N_12688);
and U14279 (N_14279,N_12615,N_13141);
nand U14280 (N_14280,N_12043,N_13186);
nand U14281 (N_14281,N_13076,N_12141);
xnor U14282 (N_14282,N_12049,N_13125);
or U14283 (N_14283,N_13142,N_13072);
nor U14284 (N_14284,N_12162,N_12211);
or U14285 (N_14285,N_12625,N_12526);
nand U14286 (N_14286,N_12445,N_12795);
nand U14287 (N_14287,N_12104,N_12670);
and U14288 (N_14288,N_12910,N_12954);
and U14289 (N_14289,N_13106,N_13072);
and U14290 (N_14290,N_13068,N_12468);
xnor U14291 (N_14291,N_12384,N_12702);
or U14292 (N_14292,N_13188,N_13050);
or U14293 (N_14293,N_12185,N_13129);
xor U14294 (N_14294,N_12089,N_13019);
or U14295 (N_14295,N_13152,N_13125);
or U14296 (N_14296,N_12457,N_13123);
nor U14297 (N_14297,N_12931,N_12000);
or U14298 (N_14298,N_12492,N_12398);
nand U14299 (N_14299,N_12884,N_12130);
nand U14300 (N_14300,N_12195,N_12685);
nor U14301 (N_14301,N_12126,N_13059);
nor U14302 (N_14302,N_13026,N_12030);
xor U14303 (N_14303,N_12258,N_13029);
nand U14304 (N_14304,N_12215,N_12275);
nor U14305 (N_14305,N_12675,N_12684);
xor U14306 (N_14306,N_12328,N_12823);
nor U14307 (N_14307,N_12427,N_12928);
nand U14308 (N_14308,N_13171,N_12754);
nand U14309 (N_14309,N_13072,N_12603);
xor U14310 (N_14310,N_12049,N_12305);
xor U14311 (N_14311,N_12019,N_12272);
nand U14312 (N_14312,N_12169,N_12858);
nor U14313 (N_14313,N_12661,N_13185);
or U14314 (N_14314,N_12583,N_13173);
nand U14315 (N_14315,N_12534,N_12078);
or U14316 (N_14316,N_12118,N_12097);
nor U14317 (N_14317,N_12790,N_12457);
nand U14318 (N_14318,N_12228,N_12290);
xnor U14319 (N_14319,N_12380,N_12602);
nor U14320 (N_14320,N_12907,N_12252);
and U14321 (N_14321,N_12320,N_12396);
or U14322 (N_14322,N_12496,N_12003);
xnor U14323 (N_14323,N_12159,N_12794);
xnor U14324 (N_14324,N_12278,N_12254);
nand U14325 (N_14325,N_12830,N_12893);
and U14326 (N_14326,N_13137,N_12421);
or U14327 (N_14327,N_12977,N_12093);
nand U14328 (N_14328,N_12454,N_13052);
xor U14329 (N_14329,N_12762,N_12139);
and U14330 (N_14330,N_13076,N_12929);
nor U14331 (N_14331,N_12487,N_12398);
nand U14332 (N_14332,N_12023,N_12015);
or U14333 (N_14333,N_13161,N_12743);
and U14334 (N_14334,N_12249,N_12673);
nor U14335 (N_14335,N_12343,N_12011);
xor U14336 (N_14336,N_12583,N_13072);
nor U14337 (N_14337,N_12787,N_12649);
nor U14338 (N_14338,N_12500,N_12699);
nor U14339 (N_14339,N_13197,N_12796);
and U14340 (N_14340,N_12993,N_13102);
and U14341 (N_14341,N_13198,N_12765);
nand U14342 (N_14342,N_13047,N_12837);
xor U14343 (N_14343,N_12624,N_12198);
nand U14344 (N_14344,N_12842,N_12957);
nor U14345 (N_14345,N_12771,N_12343);
xor U14346 (N_14346,N_12697,N_12654);
nand U14347 (N_14347,N_12117,N_12413);
or U14348 (N_14348,N_13002,N_12104);
xnor U14349 (N_14349,N_12187,N_12997);
nand U14350 (N_14350,N_12038,N_12756);
nand U14351 (N_14351,N_12502,N_12361);
nand U14352 (N_14352,N_12296,N_12893);
and U14353 (N_14353,N_12166,N_12321);
nor U14354 (N_14354,N_12953,N_12050);
and U14355 (N_14355,N_12628,N_12355);
and U14356 (N_14356,N_12842,N_12868);
nor U14357 (N_14357,N_12670,N_12184);
nand U14358 (N_14358,N_12751,N_12451);
nand U14359 (N_14359,N_12545,N_12594);
nor U14360 (N_14360,N_12586,N_13055);
or U14361 (N_14361,N_12970,N_12992);
xnor U14362 (N_14362,N_13060,N_12142);
nand U14363 (N_14363,N_12962,N_12849);
and U14364 (N_14364,N_12984,N_12128);
xor U14365 (N_14365,N_12781,N_12675);
xnor U14366 (N_14366,N_12623,N_12310);
nand U14367 (N_14367,N_12508,N_12903);
xor U14368 (N_14368,N_12279,N_13152);
xor U14369 (N_14369,N_12030,N_12691);
nand U14370 (N_14370,N_12984,N_12082);
nor U14371 (N_14371,N_12194,N_13101);
nor U14372 (N_14372,N_12003,N_12189);
xnor U14373 (N_14373,N_12391,N_12521);
xor U14374 (N_14374,N_12843,N_12883);
nand U14375 (N_14375,N_12241,N_12237);
and U14376 (N_14376,N_12589,N_12416);
and U14377 (N_14377,N_12041,N_12401);
xor U14378 (N_14378,N_12314,N_12885);
and U14379 (N_14379,N_12021,N_12539);
and U14380 (N_14380,N_12472,N_12779);
nand U14381 (N_14381,N_12430,N_12402);
and U14382 (N_14382,N_12163,N_12296);
xnor U14383 (N_14383,N_12850,N_12422);
nand U14384 (N_14384,N_12219,N_12623);
or U14385 (N_14385,N_12904,N_12598);
nand U14386 (N_14386,N_12264,N_12843);
and U14387 (N_14387,N_12185,N_12899);
nand U14388 (N_14388,N_12041,N_12376);
or U14389 (N_14389,N_12525,N_13007);
nand U14390 (N_14390,N_12026,N_13128);
or U14391 (N_14391,N_12689,N_12255);
or U14392 (N_14392,N_13198,N_12562);
nand U14393 (N_14393,N_12844,N_12821);
and U14394 (N_14394,N_12326,N_12454);
or U14395 (N_14395,N_12294,N_12824);
and U14396 (N_14396,N_12178,N_12372);
and U14397 (N_14397,N_12923,N_12006);
or U14398 (N_14398,N_12094,N_12666);
nor U14399 (N_14399,N_12537,N_12066);
or U14400 (N_14400,N_13345,N_14207);
nand U14401 (N_14401,N_13596,N_14338);
nand U14402 (N_14402,N_13661,N_13419);
or U14403 (N_14403,N_14156,N_13637);
nand U14404 (N_14404,N_14293,N_14230);
nand U14405 (N_14405,N_13587,N_13837);
nor U14406 (N_14406,N_13275,N_14070);
or U14407 (N_14407,N_14077,N_13211);
nor U14408 (N_14408,N_13464,N_13460);
xor U14409 (N_14409,N_13853,N_13733);
xnor U14410 (N_14410,N_14008,N_14387);
xor U14411 (N_14411,N_14085,N_14378);
nand U14412 (N_14412,N_13279,N_13295);
nand U14413 (N_14413,N_13442,N_14129);
nor U14414 (N_14414,N_13476,N_13795);
nand U14415 (N_14415,N_13394,N_14116);
nor U14416 (N_14416,N_14241,N_13721);
or U14417 (N_14417,N_13423,N_13754);
xnor U14418 (N_14418,N_14282,N_13767);
nand U14419 (N_14419,N_14287,N_14171);
and U14420 (N_14420,N_13550,N_13420);
and U14421 (N_14421,N_13312,N_14096);
and U14422 (N_14422,N_14039,N_13366);
nand U14423 (N_14423,N_13504,N_14323);
nor U14424 (N_14424,N_13239,N_13957);
and U14425 (N_14425,N_14149,N_13337);
nand U14426 (N_14426,N_14027,N_13919);
xor U14427 (N_14427,N_14299,N_13936);
xor U14428 (N_14428,N_14367,N_13856);
and U14429 (N_14429,N_13758,N_13991);
nor U14430 (N_14430,N_13562,N_14217);
and U14431 (N_14431,N_13411,N_14001);
and U14432 (N_14432,N_13307,N_13415);
nor U14433 (N_14433,N_14121,N_13792);
and U14434 (N_14434,N_13854,N_13468);
nand U14435 (N_14435,N_13780,N_14144);
nand U14436 (N_14436,N_14140,N_13256);
xor U14437 (N_14437,N_13593,N_13855);
or U14438 (N_14438,N_13812,N_14091);
and U14439 (N_14439,N_13392,N_13513);
xor U14440 (N_14440,N_13743,N_14320);
xnor U14441 (N_14441,N_13974,N_13799);
or U14442 (N_14442,N_13379,N_14119);
nor U14443 (N_14443,N_13893,N_13909);
nor U14444 (N_14444,N_14256,N_14086);
nand U14445 (N_14445,N_14127,N_13454);
xnor U14446 (N_14446,N_13475,N_14097);
nand U14447 (N_14447,N_13611,N_14393);
and U14448 (N_14448,N_13290,N_13787);
and U14449 (N_14449,N_13528,N_13869);
nand U14450 (N_14450,N_13745,N_13848);
nor U14451 (N_14451,N_13655,N_14161);
or U14452 (N_14452,N_13708,N_14392);
nor U14453 (N_14453,N_13929,N_13933);
nand U14454 (N_14454,N_13425,N_13542);
and U14455 (N_14455,N_13598,N_13961);
and U14456 (N_14456,N_13693,N_13453);
nor U14457 (N_14457,N_14229,N_14196);
or U14458 (N_14458,N_13206,N_13447);
and U14459 (N_14459,N_14390,N_14107);
xor U14460 (N_14460,N_14002,N_13236);
nand U14461 (N_14461,N_13253,N_13386);
nand U14462 (N_14462,N_13959,N_13289);
or U14463 (N_14463,N_14397,N_13228);
and U14464 (N_14464,N_13649,N_13638);
nand U14465 (N_14465,N_13840,N_14347);
or U14466 (N_14466,N_13716,N_13742);
and U14467 (N_14467,N_13251,N_14351);
and U14468 (N_14468,N_13535,N_13620);
xor U14469 (N_14469,N_13766,N_13696);
or U14470 (N_14470,N_13278,N_14012);
nor U14471 (N_14471,N_13597,N_13391);
and U14472 (N_14472,N_13934,N_13369);
nor U14473 (N_14473,N_14179,N_13465);
nand U14474 (N_14474,N_13280,N_13321);
or U14475 (N_14475,N_13789,N_13700);
nor U14476 (N_14476,N_14263,N_13564);
xor U14477 (N_14477,N_14058,N_13352);
nand U14478 (N_14478,N_13822,N_13348);
and U14479 (N_14479,N_13904,N_13688);
nand U14480 (N_14480,N_14246,N_13694);
and U14481 (N_14481,N_13451,N_13891);
or U14482 (N_14482,N_13783,N_13346);
and U14483 (N_14483,N_14132,N_13622);
nand U14484 (N_14484,N_13488,N_14301);
nor U14485 (N_14485,N_14218,N_13342);
nand U14486 (N_14486,N_13586,N_13599);
xor U14487 (N_14487,N_14136,N_14377);
nand U14488 (N_14488,N_13569,N_13543);
nand U14489 (N_14489,N_14098,N_13486);
nor U14490 (N_14490,N_14051,N_13452);
nor U14491 (N_14491,N_14059,N_13724);
nand U14492 (N_14492,N_13507,N_14183);
nor U14493 (N_14493,N_13613,N_14178);
nor U14494 (N_14494,N_14037,N_14208);
or U14495 (N_14495,N_13242,N_14376);
or U14496 (N_14496,N_13470,N_14385);
nand U14497 (N_14497,N_13566,N_13482);
and U14498 (N_14498,N_14381,N_14386);
and U14499 (N_14499,N_13387,N_13798);
or U14500 (N_14500,N_13894,N_13753);
nor U14501 (N_14501,N_14063,N_14092);
or U14502 (N_14502,N_14222,N_13666);
nand U14503 (N_14503,N_14305,N_14007);
xnor U14504 (N_14504,N_13466,N_14334);
nor U14505 (N_14505,N_13523,N_13714);
nand U14506 (N_14506,N_13847,N_13719);
or U14507 (N_14507,N_14360,N_13711);
or U14508 (N_14508,N_13722,N_13519);
or U14509 (N_14509,N_13305,N_13912);
xor U14510 (N_14510,N_13435,N_13725);
and U14511 (N_14511,N_13605,N_14163);
and U14512 (N_14512,N_14286,N_13201);
nor U14513 (N_14513,N_14047,N_13986);
and U14514 (N_14514,N_13262,N_13359);
and U14515 (N_14515,N_13833,N_13330);
xnor U14516 (N_14516,N_13825,N_13553);
nand U14517 (N_14517,N_13502,N_14370);
and U14518 (N_14518,N_13831,N_14266);
nand U14519 (N_14519,N_13816,N_13508);
nand U14520 (N_14520,N_14170,N_13208);
nor U14521 (N_14521,N_13281,N_13960);
or U14522 (N_14522,N_13375,N_13418);
and U14523 (N_14523,N_13492,N_14232);
or U14524 (N_14524,N_13973,N_13480);
nor U14525 (N_14525,N_14244,N_14004);
xor U14526 (N_14526,N_14214,N_13217);
and U14527 (N_14527,N_14265,N_13252);
nand U14528 (N_14528,N_14021,N_14375);
and U14529 (N_14529,N_13802,N_14368);
nor U14530 (N_14530,N_14223,N_13405);
nand U14531 (N_14531,N_13723,N_13571);
or U14532 (N_14532,N_13607,N_14036);
xor U14533 (N_14533,N_14339,N_14396);
or U14534 (N_14534,N_13695,N_13969);
or U14535 (N_14535,N_13667,N_13344);
xnor U14536 (N_14536,N_13538,N_14204);
nand U14537 (N_14537,N_13777,N_13215);
nand U14538 (N_14538,N_13669,N_14044);
or U14539 (N_14539,N_14046,N_14173);
nand U14540 (N_14540,N_13365,N_13474);
nor U14541 (N_14541,N_13608,N_14146);
or U14542 (N_14542,N_13489,N_14324);
nand U14543 (N_14543,N_13881,N_13741);
nor U14544 (N_14544,N_13601,N_14210);
nor U14545 (N_14545,N_13509,N_14193);
xor U14546 (N_14546,N_13984,N_13472);
and U14547 (N_14547,N_13690,N_13676);
nand U14548 (N_14548,N_14154,N_13210);
xnor U14549 (N_14549,N_13319,N_13925);
or U14550 (N_14550,N_13653,N_13671);
nor U14551 (N_14551,N_13589,N_13422);
nand U14552 (N_14552,N_13877,N_13529);
xnor U14553 (N_14553,N_13626,N_13632);
nor U14554 (N_14554,N_13554,N_14143);
nand U14555 (N_14555,N_14348,N_13703);
nand U14556 (N_14556,N_14174,N_13791);
nand U14557 (N_14557,N_13552,N_13225);
and U14558 (N_14558,N_13491,N_13623);
and U14559 (N_14559,N_13624,N_13769);
nand U14560 (N_14560,N_14283,N_14157);
xnor U14561 (N_14561,N_13618,N_13205);
and U14562 (N_14562,N_13786,N_14080);
or U14563 (N_14563,N_13966,N_13467);
or U14564 (N_14564,N_14043,N_14134);
and U14565 (N_14565,N_13218,N_13362);
xor U14566 (N_14566,N_14101,N_13235);
and U14567 (N_14567,N_13495,N_14245);
nor U14568 (N_14568,N_13588,N_13230);
xnor U14569 (N_14569,N_13770,N_13374);
and U14570 (N_14570,N_13709,N_14066);
xor U14571 (N_14571,N_13325,N_13682);
or U14572 (N_14572,N_14342,N_13570);
nand U14573 (N_14573,N_13292,N_13397);
or U14574 (N_14574,N_14164,N_13246);
nand U14575 (N_14575,N_13712,N_13609);
nand U14576 (N_14576,N_13287,N_14292);
nand U14577 (N_14577,N_14354,N_13885);
nand U14578 (N_14578,N_14095,N_13445);
nor U14579 (N_14579,N_13883,N_14328);
or U14580 (N_14580,N_13594,N_13313);
nand U14581 (N_14581,N_14148,N_14090);
and U14582 (N_14582,N_14177,N_13760);
or U14583 (N_14583,N_14030,N_14382);
or U14584 (N_14584,N_14309,N_14361);
xor U14585 (N_14585,N_14062,N_14306);
and U14586 (N_14586,N_13872,N_13617);
nand U14587 (N_14587,N_13240,N_14182);
nor U14588 (N_14588,N_14373,N_13970);
xnor U14589 (N_14589,N_13510,N_13430);
or U14590 (N_14590,N_14159,N_14310);
xnor U14591 (N_14591,N_13270,N_13994);
nand U14592 (N_14592,N_14285,N_14169);
or U14593 (N_14593,N_13781,N_13746);
nand U14594 (N_14594,N_13820,N_14297);
and U14595 (N_14595,N_13980,N_13326);
or U14596 (N_14596,N_14270,N_13238);
nor U14597 (N_14597,N_14003,N_13427);
nor U14598 (N_14598,N_13540,N_14316);
nor U14599 (N_14599,N_13954,N_13497);
or U14600 (N_14600,N_13839,N_13819);
and U14601 (N_14601,N_13222,N_13784);
nor U14602 (N_14602,N_13765,N_14081);
or U14603 (N_14603,N_13274,N_14048);
and U14604 (N_14604,N_13734,N_13804);
xnor U14605 (N_14605,N_13209,N_13913);
nor U14606 (N_14606,N_14155,N_14258);
or U14607 (N_14607,N_13665,N_13384);
xor U14608 (N_14608,N_13232,N_14216);
nor U14609 (N_14609,N_13884,N_14250);
or U14610 (N_14610,N_14235,N_13923);
and U14611 (N_14611,N_14065,N_14160);
and U14612 (N_14612,N_14355,N_14124);
and U14613 (N_14613,N_13660,N_13463);
nor U14614 (N_14614,N_13450,N_14296);
nand U14615 (N_14615,N_14332,N_14076);
nand U14616 (N_14616,N_14189,N_13300);
xor U14617 (N_14617,N_13591,N_13978);
nand U14618 (N_14618,N_14053,N_14278);
or U14619 (N_14619,N_13371,N_14175);
nor U14620 (N_14620,N_14333,N_13818);
nand U14621 (N_14621,N_13559,N_13437);
and U14622 (N_14622,N_13285,N_13778);
nor U14623 (N_14623,N_13875,N_14188);
or U14624 (N_14624,N_13382,N_13698);
and U14625 (N_14625,N_14389,N_13650);
and U14626 (N_14626,N_13328,N_13927);
xor U14627 (N_14627,N_14014,N_13643);
and U14628 (N_14628,N_13311,N_13568);
nand U14629 (N_14629,N_13908,N_13866);
nand U14630 (N_14630,N_14363,N_13926);
xor U14631 (N_14631,N_14005,N_14158);
xnor U14632 (N_14632,N_14365,N_13796);
nand U14633 (N_14633,N_13651,N_14371);
nor U14634 (N_14634,N_13473,N_13843);
or U14635 (N_14635,N_13942,N_13631);
and U14636 (N_14636,N_14325,N_13383);
or U14637 (N_14637,N_14331,N_14236);
nor U14638 (N_14638,N_13229,N_13677);
xor U14639 (N_14639,N_13500,N_13248);
xor U14640 (N_14640,N_14261,N_13707);
xnor U14641 (N_14641,N_13213,N_13675);
nand U14642 (N_14642,N_13544,N_14078);
and U14643 (N_14643,N_14106,N_13360);
nor U14644 (N_14644,N_13259,N_13902);
xnor U14645 (N_14645,N_13518,N_14280);
or U14646 (N_14646,N_13768,N_14277);
xnor U14647 (N_14647,N_13512,N_13801);
nand U14648 (N_14648,N_14237,N_14364);
or U14649 (N_14649,N_13424,N_13441);
or U14650 (N_14650,N_13846,N_13870);
or U14651 (N_14651,N_13814,N_13207);
or U14652 (N_14652,N_13429,N_13868);
nor U14653 (N_14653,N_14398,N_13357);
or U14654 (N_14654,N_13214,N_13494);
nor U14655 (N_14655,N_13258,N_13662);
and U14656 (N_14656,N_14307,N_13948);
nand U14657 (N_14657,N_13731,N_13426);
nor U14658 (N_14658,N_13931,N_14259);
and U14659 (N_14659,N_13989,N_14167);
and U14660 (N_14660,N_13315,N_14304);
and U14661 (N_14661,N_13479,N_13911);
nor U14662 (N_14662,N_13499,N_13390);
nand U14663 (N_14663,N_13496,N_13490);
and U14664 (N_14664,N_14289,N_13436);
xnor U14665 (N_14665,N_14372,N_13800);
and U14666 (N_14666,N_13503,N_14340);
xor U14667 (N_14667,N_14327,N_14288);
or U14668 (N_14668,N_13979,N_13739);
and U14669 (N_14669,N_13906,N_13889);
and U14670 (N_14670,N_13581,N_13811);
or U14671 (N_14671,N_13318,N_13546);
or U14672 (N_14672,N_14290,N_13324);
nor U14673 (N_14673,N_13537,N_14011);
or U14674 (N_14674,N_13697,N_14349);
nand U14675 (N_14675,N_13575,N_13958);
xor U14676 (N_14676,N_13481,N_13341);
or U14677 (N_14677,N_13557,N_13354);
nor U14678 (N_14678,N_13203,N_13975);
xnor U14679 (N_14679,N_13938,N_14087);
or U14680 (N_14680,N_13815,N_14329);
nor U14681 (N_14681,N_14145,N_13776);
and U14682 (N_14682,N_14114,N_13773);
xor U14683 (N_14683,N_13996,N_13336);
nor U14684 (N_14684,N_14069,N_13968);
xnor U14685 (N_14685,N_13294,N_13381);
or U14686 (N_14686,N_13993,N_13668);
and U14687 (N_14687,N_13462,N_14123);
nand U14688 (N_14688,N_13433,N_13320);
xnor U14689 (N_14689,N_14399,N_14049);
and U14690 (N_14690,N_13531,N_13615);
xnor U14691 (N_14691,N_13983,N_13790);
nor U14692 (N_14692,N_13385,N_14023);
xor U14693 (N_14693,N_14060,N_14165);
nor U14694 (N_14694,N_13924,N_13556);
xor U14695 (N_14695,N_14052,N_14253);
or U14696 (N_14696,N_14317,N_13431);
xnor U14697 (N_14697,N_14084,N_14191);
nand U14698 (N_14698,N_13678,N_14100);
or U14699 (N_14699,N_13673,N_13641);
nand U14700 (N_14700,N_13689,N_13343);
and U14701 (N_14701,N_14019,N_13656);
and U14702 (N_14702,N_14168,N_13652);
nand U14703 (N_14703,N_13409,N_14029);
xnor U14704 (N_14704,N_13679,N_14279);
xor U14705 (N_14705,N_13861,N_13692);
or U14706 (N_14706,N_13304,N_14291);
xnor U14707 (N_14707,N_14026,N_13477);
or U14708 (N_14708,N_13301,N_13827);
and U14709 (N_14709,N_13558,N_14141);
nand U14710 (N_14710,N_13710,N_13751);
xor U14711 (N_14711,N_13867,N_13522);
xnor U14712 (N_14712,N_14273,N_13947);
xnor U14713 (N_14713,N_14064,N_13627);
or U14714 (N_14714,N_13396,N_14284);
xor U14715 (N_14715,N_14018,N_14135);
xor U14716 (N_14716,N_13298,N_13368);
nor U14717 (N_14717,N_13967,N_14035);
xnor U14718 (N_14718,N_13567,N_13541);
nand U14719 (N_14719,N_13525,N_13458);
or U14720 (N_14720,N_13828,N_13630);
xor U14721 (N_14721,N_13521,N_13713);
nor U14722 (N_14722,N_14198,N_13579);
or U14723 (N_14723,N_13879,N_13720);
and U14724 (N_14724,N_13842,N_14079);
xnor U14725 (N_14725,N_13511,N_13917);
nor U14726 (N_14726,N_13972,N_13204);
and U14727 (N_14727,N_13932,N_13921);
and U14728 (N_14728,N_13578,N_13705);
xnor U14729 (N_14729,N_13438,N_13681);
xor U14730 (N_14730,N_14089,N_14366);
xor U14731 (N_14731,N_13417,N_14010);
nand U14732 (N_14732,N_14192,N_14082);
and U14733 (N_14733,N_13310,N_13400);
or U14734 (N_14734,N_14269,N_14153);
xor U14735 (N_14735,N_13990,N_13226);
or U14736 (N_14736,N_13603,N_14212);
and U14737 (N_14737,N_13378,N_14335);
and U14738 (N_14738,N_14142,N_13404);
or U14739 (N_14739,N_13737,N_13347);
nand U14740 (N_14740,N_13612,N_13272);
and U14741 (N_14741,N_13871,N_13971);
or U14742 (N_14742,N_14015,N_13779);
or U14743 (N_14743,N_13728,N_14150);
nand U14744 (N_14744,N_14345,N_14383);
xor U14745 (N_14745,N_14315,N_13901);
nand U14746 (N_14746,N_13772,N_13691);
nor U14747 (N_14747,N_14394,N_13952);
and U14748 (N_14748,N_13234,N_13629);
nand U14749 (N_14749,N_13469,N_13685);
nand U14750 (N_14750,N_13551,N_13805);
nand U14751 (N_14751,N_13857,N_13530);
xor U14752 (N_14752,N_13532,N_13316);
nor U14753 (N_14753,N_13555,N_13604);
nor U14754 (N_14754,N_13271,N_13955);
or U14755 (N_14755,N_14350,N_13233);
nor U14756 (N_14756,N_13764,N_14209);
nor U14757 (N_14757,N_14352,N_13389);
or U14758 (N_14758,N_14308,N_13899);
nand U14759 (N_14759,N_13220,N_13412);
or U14760 (N_14760,N_13761,N_13880);
or U14761 (N_14761,N_14337,N_14226);
or U14762 (N_14762,N_13610,N_14126);
or U14763 (N_14763,N_13434,N_13953);
or U14764 (N_14764,N_14379,N_14017);
nor U14765 (N_14765,N_13250,N_14219);
nor U14766 (N_14766,N_13444,N_13224);
nand U14767 (N_14767,N_13351,N_13729);
nand U14768 (N_14768,N_13633,N_13327);
and U14769 (N_14769,N_13756,N_14211);
and U14770 (N_14770,N_13399,N_14055);
nand U14771 (N_14771,N_14103,N_13640);
or U14772 (N_14772,N_14302,N_14120);
nand U14773 (N_14773,N_14110,N_14061);
nand U14774 (N_14774,N_13506,N_13997);
xor U14775 (N_14775,N_13254,N_13928);
or U14776 (N_14776,N_14025,N_14067);
nand U14777 (N_14777,N_14228,N_13358);
nand U14778 (N_14778,N_13549,N_14006);
and U14779 (N_14779,N_13459,N_13355);
nor U14780 (N_14780,N_13943,N_13350);
nand U14781 (N_14781,N_13353,N_14264);
xor U14782 (N_14782,N_13393,N_13995);
or U14783 (N_14783,N_14176,N_14343);
nand U14784 (N_14784,N_13704,N_13548);
nor U14785 (N_14785,N_13657,N_14380);
or U14786 (N_14786,N_13410,N_14073);
nand U14787 (N_14787,N_14072,N_13600);
nor U14788 (N_14788,N_13858,N_13949);
xnor U14789 (N_14789,N_13247,N_13916);
xnor U14790 (N_14790,N_14321,N_14083);
or U14791 (N_14791,N_14113,N_13896);
and U14792 (N_14792,N_13363,N_13874);
or U14793 (N_14793,N_14201,N_13876);
nand U14794 (N_14794,N_13982,N_13565);
nand U14795 (N_14795,N_13408,N_13376);
xnor U14796 (N_14796,N_13628,N_14028);
xnor U14797 (N_14797,N_13976,N_13621);
nor U14798 (N_14798,N_13634,N_13699);
nand U14799 (N_14799,N_13487,N_14009);
nand U14800 (N_14800,N_13985,N_13915);
nand U14801 (N_14801,N_13664,N_14088);
and U14802 (N_14802,N_13416,N_13821);
xnor U14803 (N_14803,N_13515,N_13775);
nand U14804 (N_14804,N_13484,N_13998);
or U14805 (N_14805,N_14187,N_14233);
and U14806 (N_14806,N_13888,N_13483);
xor U14807 (N_14807,N_14068,N_13293);
nand U14808 (N_14808,N_13439,N_14369);
nand U14809 (N_14809,N_13288,N_13808);
nand U14810 (N_14810,N_14147,N_14094);
and U14811 (N_14811,N_13574,N_13702);
and U14812 (N_14812,N_13255,N_14162);
xnor U14813 (N_14813,N_13448,N_13717);
nand U14814 (N_14814,N_13810,N_14054);
nand U14815 (N_14815,N_13266,N_13331);
xnor U14816 (N_14816,N_13334,N_13738);
nor U14817 (N_14817,N_14190,N_13402);
and U14818 (N_14818,N_13388,N_13478);
xor U14819 (N_14819,N_14016,N_13432);
nor U14820 (N_14820,N_13276,N_14319);
xor U14821 (N_14821,N_13296,N_14311);
nand U14822 (N_14822,N_13687,N_13674);
nand U14823 (N_14823,N_13349,N_13735);
nand U14824 (N_14824,N_14137,N_13440);
or U14825 (N_14825,N_14013,N_14075);
or U14826 (N_14826,N_13686,N_13306);
xor U14827 (N_14827,N_13261,N_13264);
nor U14828 (N_14828,N_14194,N_14112);
nand U14829 (N_14829,N_14224,N_14131);
and U14830 (N_14830,N_14151,N_14166);
xnor U14831 (N_14831,N_13922,N_13260);
and U14832 (N_14832,N_13706,N_13299);
nor U14833 (N_14833,N_13658,N_13524);
nand U14834 (N_14834,N_14215,N_13284);
nand U14835 (N_14835,N_14243,N_13886);
and U14836 (N_14836,N_14254,N_14318);
nor U14837 (N_14837,N_13583,N_13841);
and U14838 (N_14838,N_13851,N_13606);
nor U14839 (N_14839,N_14034,N_13268);
nand U14840 (N_14840,N_13749,N_14038);
nand U14841 (N_14841,N_13788,N_14109);
or U14842 (N_14842,N_14357,N_14071);
and U14843 (N_14843,N_13887,N_13803);
or U14844 (N_14844,N_13941,N_13782);
nor U14845 (N_14845,N_14195,N_13414);
nand U14846 (N_14846,N_13635,N_14268);
nor U14847 (N_14847,N_13826,N_13560);
nand U14848 (N_14848,N_13774,N_13534);
and U14849 (N_14849,N_13263,N_13547);
xor U14850 (N_14850,N_14122,N_13838);
and U14851 (N_14851,N_13807,N_14313);
and U14852 (N_14852,N_13644,N_14181);
nor U14853 (N_14853,N_13446,N_13683);
and U14854 (N_14854,N_14041,N_13964);
and U14855 (N_14855,N_14200,N_13329);
or U14856 (N_14856,N_13536,N_13335);
or U14857 (N_14857,N_13663,N_14359);
nor U14858 (N_14858,N_13987,N_13297);
and U14859 (N_14859,N_13339,N_13977);
nand U14860 (N_14860,N_14128,N_13937);
nand U14861 (N_14861,N_13785,N_14099);
xnor U14862 (N_14862,N_13730,N_13829);
xor U14863 (N_14863,N_13830,N_13602);
nand U14864 (N_14864,N_13377,N_14274);
or U14865 (N_14865,N_13625,N_14395);
xor U14866 (N_14866,N_14248,N_13231);
xor U14867 (N_14867,N_14234,N_13905);
and U14868 (N_14868,N_13813,N_13950);
nor U14869 (N_14869,N_14353,N_13501);
and U14870 (N_14870,N_14260,N_13763);
or U14871 (N_14871,N_13865,N_14102);
xor U14872 (N_14872,N_13249,N_14262);
or U14873 (N_14873,N_13265,N_13939);
nor U14874 (N_14874,N_14257,N_13527);
or U14875 (N_14875,N_13338,N_13573);
nand U14876 (N_14876,N_14238,N_14239);
nor U14877 (N_14877,N_13380,N_13680);
nand U14878 (N_14878,N_13824,N_14186);
nor U14879 (N_14879,N_13845,N_13744);
nand U14880 (N_14880,N_13670,N_14050);
or U14881 (N_14881,N_13930,N_14115);
nor U14882 (N_14882,N_13317,N_14356);
xnor U14883 (N_14883,N_14295,N_14202);
nor U14884 (N_14884,N_13514,N_14111);
nand U14885 (N_14885,N_13449,N_14133);
or U14886 (N_14886,N_14251,N_13903);
xnor U14887 (N_14887,N_13455,N_14125);
xnor U14888 (N_14888,N_13291,N_13636);
nand U14889 (N_14889,N_14197,N_14104);
xnor U14890 (N_14890,N_13457,N_13956);
nand U14891 (N_14891,N_13793,N_13561);
nor U14892 (N_14892,N_13322,N_13576);
nor U14893 (N_14893,N_13648,N_13834);
or U14894 (N_14894,N_13309,N_14031);
nand U14895 (N_14895,N_13572,N_14185);
or U14896 (N_14896,N_13373,N_13963);
nor U14897 (N_14897,N_13493,N_14118);
or U14898 (N_14898,N_13332,N_14252);
and U14899 (N_14899,N_14108,N_14093);
nand U14900 (N_14900,N_13372,N_13944);
xor U14901 (N_14901,N_14242,N_13835);
and U14902 (N_14902,N_13740,N_13282);
nor U14903 (N_14903,N_14000,N_13461);
or U14904 (N_14904,N_13223,N_14040);
or U14905 (N_14905,N_14391,N_14213);
and U14906 (N_14906,N_14303,N_13485);
nor U14907 (N_14907,N_13962,N_13750);
or U14908 (N_14908,N_13752,N_14152);
and U14909 (N_14909,N_13992,N_14255);
or U14910 (N_14910,N_14227,N_14074);
and U14911 (N_14911,N_13595,N_14024);
xnor U14912 (N_14912,N_14184,N_13882);
and U14913 (N_14913,N_13809,N_13584);
nor U14914 (N_14914,N_14384,N_14220);
nand U14915 (N_14915,N_13257,N_14346);
nand U14916 (N_14916,N_13619,N_14336);
and U14917 (N_14917,N_13726,N_14022);
xor U14918 (N_14918,N_13273,N_13277);
and U14919 (N_14919,N_13935,N_13237);
xnor U14920 (N_14920,N_13406,N_13403);
xor U14921 (N_14921,N_13940,N_13227);
and U14922 (N_14922,N_13202,N_14203);
nand U14923 (N_14923,N_14206,N_14330);
xnor U14924 (N_14924,N_13859,N_14199);
and U14925 (N_14925,N_13577,N_13897);
and U14926 (N_14926,N_13900,N_13592);
or U14927 (N_14927,N_13946,N_13401);
nor U14928 (N_14928,N_13647,N_13614);
or U14929 (N_14929,N_13907,N_13757);
nand U14930 (N_14930,N_13890,N_13988);
xnor U14931 (N_14931,N_13302,N_13898);
nor U14932 (N_14932,N_13684,N_14341);
or U14933 (N_14933,N_13267,N_13981);
nand U14934 (N_14934,N_13863,N_13732);
nand U14935 (N_14935,N_14267,N_13616);
nor U14936 (N_14936,N_13243,N_14300);
xnor U14937 (N_14937,N_13823,N_13516);
nor U14938 (N_14938,N_14344,N_13832);
xor U14939 (N_14939,N_13836,N_13794);
xnor U14940 (N_14940,N_14042,N_13755);
or U14941 (N_14941,N_13639,N_13413);
nand U14942 (N_14942,N_13520,N_14271);
and U14943 (N_14943,N_13771,N_14275);
or U14944 (N_14944,N_14056,N_13759);
or U14945 (N_14945,N_13672,N_13718);
and U14946 (N_14946,N_13286,N_14130);
and U14947 (N_14947,N_13920,N_13545);
and U14948 (N_14948,N_13862,N_14388);
xnor U14949 (N_14949,N_13428,N_13241);
xor U14950 (N_14950,N_14247,N_14249);
xor U14951 (N_14951,N_13443,N_13701);
nand U14952 (N_14952,N_14033,N_13303);
nor U14953 (N_14953,N_14281,N_14057);
nor U14954 (N_14954,N_13999,N_13918);
and U14955 (N_14955,N_13367,N_13539);
or U14956 (N_14956,N_13817,N_13421);
nor U14957 (N_14957,N_14362,N_13736);
nand U14958 (N_14958,N_13216,N_13762);
xor U14959 (N_14959,N_13844,N_13456);
xor U14960 (N_14960,N_14225,N_13364);
nand U14961 (N_14961,N_13398,N_14221);
xnor U14962 (N_14962,N_13333,N_13370);
nand U14963 (N_14963,N_13806,N_13244);
nor U14964 (N_14964,N_13659,N_13526);
and U14965 (N_14965,N_13878,N_13715);
nor U14966 (N_14966,N_13590,N_14240);
or U14967 (N_14967,N_14358,N_14105);
nor U14968 (N_14968,N_14138,N_13727);
nand U14969 (N_14969,N_13895,N_13748);
nand U14970 (N_14970,N_13849,N_13361);
nand U14971 (N_14971,N_13395,N_14326);
and U14972 (N_14972,N_13797,N_14272);
nand U14973 (N_14973,N_14322,N_13219);
nand U14974 (N_14974,N_13407,N_14172);
and U14975 (N_14975,N_13645,N_13245);
nand U14976 (N_14976,N_13951,N_14020);
or U14977 (N_14977,N_14139,N_13585);
nor U14978 (N_14978,N_13283,N_13646);
and U14979 (N_14979,N_13945,N_13860);
or U14980 (N_14980,N_13323,N_14298);
nor U14981 (N_14981,N_13580,N_13314);
or U14982 (N_14982,N_13212,N_13654);
nor U14983 (N_14983,N_13356,N_13517);
xnor U14984 (N_14984,N_13850,N_13747);
and U14985 (N_14985,N_13892,N_13873);
and U14986 (N_14986,N_14314,N_14294);
xnor U14987 (N_14987,N_13340,N_13914);
nand U14988 (N_14988,N_14045,N_13563);
and U14989 (N_14989,N_14205,N_13642);
or U14990 (N_14990,N_13910,N_14312);
nor U14991 (N_14991,N_14231,N_13864);
xnor U14992 (N_14992,N_13308,N_14032);
nand U14993 (N_14993,N_13221,N_13582);
nor U14994 (N_14994,N_13533,N_13498);
or U14995 (N_14995,N_14276,N_14374);
nor U14996 (N_14996,N_13965,N_13269);
nor U14997 (N_14997,N_14180,N_13200);
or U14998 (N_14998,N_13471,N_13505);
nor U14999 (N_14999,N_14117,N_13852);
or U15000 (N_15000,N_14095,N_14252);
or U15001 (N_15001,N_14294,N_14269);
and U15002 (N_15002,N_13332,N_13934);
or U15003 (N_15003,N_14248,N_14273);
nand U15004 (N_15004,N_13271,N_13962);
xnor U15005 (N_15005,N_13301,N_14091);
nand U15006 (N_15006,N_13595,N_13503);
and U15007 (N_15007,N_14382,N_13871);
or U15008 (N_15008,N_14371,N_13270);
xnor U15009 (N_15009,N_13563,N_14191);
or U15010 (N_15010,N_13809,N_14347);
and U15011 (N_15011,N_14384,N_13691);
nand U15012 (N_15012,N_13625,N_13494);
nand U15013 (N_15013,N_13887,N_14293);
and U15014 (N_15014,N_13377,N_14159);
xnor U15015 (N_15015,N_13659,N_13820);
xnor U15016 (N_15016,N_14262,N_14023);
nand U15017 (N_15017,N_14299,N_13286);
nand U15018 (N_15018,N_13339,N_13600);
and U15019 (N_15019,N_14192,N_13333);
nand U15020 (N_15020,N_13778,N_14266);
nor U15021 (N_15021,N_14320,N_13645);
nor U15022 (N_15022,N_13873,N_14119);
xor U15023 (N_15023,N_13549,N_14051);
nand U15024 (N_15024,N_14238,N_13583);
or U15025 (N_15025,N_13453,N_13330);
or U15026 (N_15026,N_13903,N_13360);
xor U15027 (N_15027,N_14300,N_13402);
or U15028 (N_15028,N_14252,N_13700);
and U15029 (N_15029,N_13985,N_13391);
xnor U15030 (N_15030,N_14299,N_13505);
nand U15031 (N_15031,N_14050,N_13416);
xnor U15032 (N_15032,N_13643,N_14069);
or U15033 (N_15033,N_13456,N_14037);
nor U15034 (N_15034,N_13210,N_14132);
and U15035 (N_15035,N_14104,N_13979);
xor U15036 (N_15036,N_13374,N_13293);
nand U15037 (N_15037,N_13561,N_14019);
or U15038 (N_15038,N_13896,N_14230);
and U15039 (N_15039,N_14305,N_14271);
and U15040 (N_15040,N_13901,N_13635);
nor U15041 (N_15041,N_13695,N_14349);
nand U15042 (N_15042,N_14083,N_14034);
xnor U15043 (N_15043,N_13596,N_13932);
or U15044 (N_15044,N_14196,N_13517);
nand U15045 (N_15045,N_14181,N_13619);
and U15046 (N_15046,N_13792,N_14029);
nor U15047 (N_15047,N_14281,N_14225);
xor U15048 (N_15048,N_13376,N_14172);
or U15049 (N_15049,N_13393,N_13272);
and U15050 (N_15050,N_14319,N_14237);
or U15051 (N_15051,N_14351,N_13400);
xnor U15052 (N_15052,N_13806,N_14088);
xnor U15053 (N_15053,N_13348,N_13337);
xnor U15054 (N_15054,N_14325,N_14349);
xor U15055 (N_15055,N_13437,N_14227);
nand U15056 (N_15056,N_13571,N_13945);
and U15057 (N_15057,N_13436,N_14357);
nor U15058 (N_15058,N_14359,N_14249);
and U15059 (N_15059,N_13752,N_14084);
or U15060 (N_15060,N_13497,N_13715);
or U15061 (N_15061,N_14032,N_13549);
nand U15062 (N_15062,N_13469,N_14064);
nand U15063 (N_15063,N_14063,N_13377);
xor U15064 (N_15064,N_13470,N_13914);
xor U15065 (N_15065,N_13442,N_13943);
or U15066 (N_15066,N_14328,N_13328);
and U15067 (N_15067,N_13857,N_13827);
and U15068 (N_15068,N_13385,N_13572);
nor U15069 (N_15069,N_14011,N_13554);
xnor U15070 (N_15070,N_13706,N_13694);
nor U15071 (N_15071,N_14011,N_13557);
or U15072 (N_15072,N_14250,N_13607);
nor U15073 (N_15073,N_13205,N_13224);
nor U15074 (N_15074,N_13232,N_13688);
nor U15075 (N_15075,N_14262,N_14386);
and U15076 (N_15076,N_14361,N_13258);
nor U15077 (N_15077,N_14316,N_13480);
nand U15078 (N_15078,N_13400,N_13982);
xnor U15079 (N_15079,N_13268,N_14214);
nor U15080 (N_15080,N_13573,N_13717);
or U15081 (N_15081,N_13702,N_14101);
xor U15082 (N_15082,N_14154,N_13725);
and U15083 (N_15083,N_14038,N_13745);
and U15084 (N_15084,N_13297,N_14181);
xnor U15085 (N_15085,N_14313,N_14315);
nor U15086 (N_15086,N_13326,N_13345);
or U15087 (N_15087,N_13841,N_13628);
nand U15088 (N_15088,N_14393,N_13533);
or U15089 (N_15089,N_13228,N_13586);
nand U15090 (N_15090,N_13245,N_13348);
nor U15091 (N_15091,N_14220,N_13825);
nor U15092 (N_15092,N_13725,N_13245);
and U15093 (N_15093,N_14293,N_13905);
or U15094 (N_15094,N_13921,N_13275);
xor U15095 (N_15095,N_13597,N_14351);
or U15096 (N_15096,N_13955,N_14249);
and U15097 (N_15097,N_13903,N_14177);
and U15098 (N_15098,N_13848,N_13702);
xnor U15099 (N_15099,N_13686,N_13697);
nand U15100 (N_15100,N_14018,N_14300);
xor U15101 (N_15101,N_13327,N_13780);
xor U15102 (N_15102,N_13727,N_14145);
or U15103 (N_15103,N_13521,N_14318);
xor U15104 (N_15104,N_13576,N_14000);
nor U15105 (N_15105,N_13972,N_13862);
or U15106 (N_15106,N_14227,N_13859);
and U15107 (N_15107,N_13264,N_14394);
and U15108 (N_15108,N_13216,N_14165);
or U15109 (N_15109,N_14290,N_13310);
xnor U15110 (N_15110,N_13707,N_13338);
nand U15111 (N_15111,N_13987,N_14014);
nor U15112 (N_15112,N_13583,N_13737);
and U15113 (N_15113,N_13933,N_13510);
nor U15114 (N_15114,N_13908,N_13423);
and U15115 (N_15115,N_14394,N_14185);
nand U15116 (N_15116,N_13455,N_13772);
or U15117 (N_15117,N_13221,N_14276);
nand U15118 (N_15118,N_13696,N_14034);
or U15119 (N_15119,N_14152,N_13579);
nand U15120 (N_15120,N_13923,N_13920);
nand U15121 (N_15121,N_13650,N_14180);
nand U15122 (N_15122,N_14380,N_13613);
nor U15123 (N_15123,N_13800,N_13568);
nand U15124 (N_15124,N_14255,N_13812);
nor U15125 (N_15125,N_13897,N_13418);
nor U15126 (N_15126,N_13216,N_14042);
or U15127 (N_15127,N_13940,N_14239);
xor U15128 (N_15128,N_13450,N_14045);
and U15129 (N_15129,N_13972,N_13304);
xnor U15130 (N_15130,N_14310,N_14379);
xnor U15131 (N_15131,N_14350,N_13753);
and U15132 (N_15132,N_13674,N_14024);
and U15133 (N_15133,N_14258,N_13820);
and U15134 (N_15134,N_14233,N_13278);
and U15135 (N_15135,N_14238,N_14200);
xor U15136 (N_15136,N_14241,N_13977);
nor U15137 (N_15137,N_13599,N_13584);
and U15138 (N_15138,N_14042,N_14077);
and U15139 (N_15139,N_14194,N_14207);
nor U15140 (N_15140,N_14151,N_13402);
or U15141 (N_15141,N_13352,N_13787);
xor U15142 (N_15142,N_13499,N_14398);
and U15143 (N_15143,N_13501,N_13982);
nand U15144 (N_15144,N_13322,N_13249);
nand U15145 (N_15145,N_13615,N_13666);
xnor U15146 (N_15146,N_13370,N_13783);
nand U15147 (N_15147,N_13273,N_14001);
and U15148 (N_15148,N_14317,N_14152);
nor U15149 (N_15149,N_13376,N_14220);
nor U15150 (N_15150,N_13387,N_14085);
nor U15151 (N_15151,N_13349,N_14373);
nand U15152 (N_15152,N_14308,N_14265);
xor U15153 (N_15153,N_14312,N_13642);
nor U15154 (N_15154,N_13507,N_14055);
xnor U15155 (N_15155,N_13672,N_13756);
or U15156 (N_15156,N_13902,N_14112);
nand U15157 (N_15157,N_13798,N_13701);
and U15158 (N_15158,N_13436,N_13751);
nand U15159 (N_15159,N_14266,N_14113);
or U15160 (N_15160,N_13339,N_13586);
xor U15161 (N_15161,N_14269,N_14086);
nor U15162 (N_15162,N_14310,N_13496);
nor U15163 (N_15163,N_14073,N_13539);
xor U15164 (N_15164,N_14121,N_13260);
or U15165 (N_15165,N_14203,N_13750);
xnor U15166 (N_15166,N_13364,N_14389);
nor U15167 (N_15167,N_13805,N_13349);
or U15168 (N_15168,N_13427,N_13865);
xnor U15169 (N_15169,N_13890,N_14250);
nand U15170 (N_15170,N_13698,N_13644);
nand U15171 (N_15171,N_13284,N_13671);
or U15172 (N_15172,N_13218,N_14393);
nor U15173 (N_15173,N_14393,N_13481);
nand U15174 (N_15174,N_13961,N_13584);
or U15175 (N_15175,N_13259,N_13248);
xor U15176 (N_15176,N_13732,N_14028);
xnor U15177 (N_15177,N_14370,N_13233);
or U15178 (N_15178,N_13909,N_13654);
or U15179 (N_15179,N_13948,N_13653);
or U15180 (N_15180,N_14080,N_13586);
or U15181 (N_15181,N_14068,N_13711);
and U15182 (N_15182,N_13457,N_13410);
nand U15183 (N_15183,N_13637,N_13981);
and U15184 (N_15184,N_13263,N_13337);
xnor U15185 (N_15185,N_14037,N_13281);
and U15186 (N_15186,N_13581,N_14263);
and U15187 (N_15187,N_13378,N_14304);
or U15188 (N_15188,N_13396,N_13951);
nor U15189 (N_15189,N_13989,N_13268);
and U15190 (N_15190,N_13780,N_14130);
nor U15191 (N_15191,N_13382,N_14092);
xnor U15192 (N_15192,N_13347,N_13904);
and U15193 (N_15193,N_13223,N_13336);
nand U15194 (N_15194,N_13817,N_13507);
xnor U15195 (N_15195,N_14160,N_13518);
and U15196 (N_15196,N_14208,N_13685);
or U15197 (N_15197,N_13768,N_13910);
xnor U15198 (N_15198,N_13756,N_13799);
nor U15199 (N_15199,N_13340,N_13236);
and U15200 (N_15200,N_14007,N_13885);
and U15201 (N_15201,N_14195,N_14010);
and U15202 (N_15202,N_13964,N_14069);
nand U15203 (N_15203,N_14188,N_13631);
and U15204 (N_15204,N_14206,N_13690);
and U15205 (N_15205,N_13226,N_13920);
and U15206 (N_15206,N_14151,N_13318);
nand U15207 (N_15207,N_13880,N_13804);
nand U15208 (N_15208,N_13581,N_13288);
nor U15209 (N_15209,N_13567,N_13308);
and U15210 (N_15210,N_13233,N_14355);
xnor U15211 (N_15211,N_14097,N_13745);
xnor U15212 (N_15212,N_14076,N_13988);
and U15213 (N_15213,N_13773,N_13392);
or U15214 (N_15214,N_14338,N_14161);
nor U15215 (N_15215,N_14070,N_13994);
or U15216 (N_15216,N_13441,N_14068);
nand U15217 (N_15217,N_14146,N_13786);
nand U15218 (N_15218,N_13734,N_13234);
and U15219 (N_15219,N_14396,N_13798);
nor U15220 (N_15220,N_13705,N_14349);
nand U15221 (N_15221,N_13224,N_13308);
xnor U15222 (N_15222,N_13941,N_13733);
and U15223 (N_15223,N_13922,N_14327);
xnor U15224 (N_15224,N_13914,N_14231);
or U15225 (N_15225,N_14313,N_14231);
and U15226 (N_15226,N_13549,N_13416);
nor U15227 (N_15227,N_13589,N_13720);
xnor U15228 (N_15228,N_13998,N_13873);
xor U15229 (N_15229,N_13526,N_14279);
and U15230 (N_15230,N_13883,N_13669);
xor U15231 (N_15231,N_13261,N_14332);
or U15232 (N_15232,N_13871,N_14082);
and U15233 (N_15233,N_14363,N_13980);
or U15234 (N_15234,N_14232,N_14366);
nand U15235 (N_15235,N_13500,N_13494);
nor U15236 (N_15236,N_14056,N_13758);
nand U15237 (N_15237,N_13338,N_13200);
nor U15238 (N_15238,N_13292,N_14137);
nor U15239 (N_15239,N_13978,N_13263);
xor U15240 (N_15240,N_13783,N_13902);
nand U15241 (N_15241,N_14278,N_13920);
nor U15242 (N_15242,N_14328,N_13886);
or U15243 (N_15243,N_13870,N_13284);
nor U15244 (N_15244,N_13324,N_13645);
nor U15245 (N_15245,N_13772,N_13204);
and U15246 (N_15246,N_13785,N_13544);
nor U15247 (N_15247,N_13581,N_13424);
xnor U15248 (N_15248,N_13882,N_14282);
xnor U15249 (N_15249,N_13453,N_13402);
xnor U15250 (N_15250,N_13727,N_13599);
nor U15251 (N_15251,N_13435,N_13613);
xnor U15252 (N_15252,N_14248,N_13417);
xor U15253 (N_15253,N_13988,N_13951);
nor U15254 (N_15254,N_13744,N_13436);
nor U15255 (N_15255,N_14287,N_13785);
and U15256 (N_15256,N_13596,N_13926);
xor U15257 (N_15257,N_13290,N_13874);
nor U15258 (N_15258,N_14178,N_13684);
nor U15259 (N_15259,N_13249,N_13508);
xor U15260 (N_15260,N_14359,N_13749);
or U15261 (N_15261,N_13515,N_13267);
nor U15262 (N_15262,N_13449,N_14345);
and U15263 (N_15263,N_13767,N_13812);
and U15264 (N_15264,N_13885,N_13360);
nand U15265 (N_15265,N_13966,N_14170);
xor U15266 (N_15266,N_13301,N_13450);
nor U15267 (N_15267,N_13633,N_13333);
nor U15268 (N_15268,N_14196,N_13953);
nor U15269 (N_15269,N_13326,N_13583);
xnor U15270 (N_15270,N_14226,N_14370);
and U15271 (N_15271,N_14006,N_14152);
or U15272 (N_15272,N_14167,N_14193);
xor U15273 (N_15273,N_13341,N_14005);
nand U15274 (N_15274,N_13317,N_14248);
and U15275 (N_15275,N_13848,N_14354);
and U15276 (N_15276,N_13478,N_14201);
xor U15277 (N_15277,N_13359,N_13544);
or U15278 (N_15278,N_13279,N_14178);
or U15279 (N_15279,N_13997,N_13938);
nor U15280 (N_15280,N_14223,N_14043);
or U15281 (N_15281,N_13896,N_14364);
nand U15282 (N_15282,N_13610,N_13835);
nor U15283 (N_15283,N_13426,N_14370);
nand U15284 (N_15284,N_14009,N_13624);
nand U15285 (N_15285,N_13954,N_13993);
nand U15286 (N_15286,N_13888,N_13880);
nor U15287 (N_15287,N_13256,N_14094);
nand U15288 (N_15288,N_13630,N_14043);
xnor U15289 (N_15289,N_13945,N_14091);
nand U15290 (N_15290,N_14083,N_14345);
xor U15291 (N_15291,N_14312,N_14244);
nand U15292 (N_15292,N_13939,N_13470);
nor U15293 (N_15293,N_13915,N_14228);
nand U15294 (N_15294,N_13982,N_13349);
xor U15295 (N_15295,N_13730,N_13366);
xor U15296 (N_15296,N_14002,N_13461);
nor U15297 (N_15297,N_13441,N_14344);
nand U15298 (N_15298,N_13664,N_14325);
or U15299 (N_15299,N_14063,N_14046);
nand U15300 (N_15300,N_13717,N_14190);
or U15301 (N_15301,N_14350,N_13640);
or U15302 (N_15302,N_13528,N_13445);
nor U15303 (N_15303,N_13432,N_14299);
or U15304 (N_15304,N_13712,N_13312);
xor U15305 (N_15305,N_13850,N_13504);
nor U15306 (N_15306,N_13571,N_13736);
or U15307 (N_15307,N_13971,N_14258);
xnor U15308 (N_15308,N_13265,N_14328);
xnor U15309 (N_15309,N_13668,N_13597);
or U15310 (N_15310,N_13597,N_13459);
and U15311 (N_15311,N_13689,N_14369);
and U15312 (N_15312,N_14277,N_13542);
or U15313 (N_15313,N_14207,N_13238);
and U15314 (N_15314,N_13707,N_13804);
nand U15315 (N_15315,N_13474,N_13592);
nand U15316 (N_15316,N_13390,N_14185);
or U15317 (N_15317,N_13414,N_13442);
nor U15318 (N_15318,N_13302,N_13258);
nand U15319 (N_15319,N_14089,N_13582);
or U15320 (N_15320,N_14157,N_13781);
and U15321 (N_15321,N_13267,N_13317);
nor U15322 (N_15322,N_13703,N_13850);
nand U15323 (N_15323,N_13942,N_13441);
or U15324 (N_15324,N_13395,N_13243);
and U15325 (N_15325,N_13972,N_13268);
or U15326 (N_15326,N_14308,N_13773);
xor U15327 (N_15327,N_13969,N_13603);
nor U15328 (N_15328,N_13837,N_14179);
nor U15329 (N_15329,N_13944,N_14321);
and U15330 (N_15330,N_13874,N_14378);
nand U15331 (N_15331,N_14151,N_13690);
nand U15332 (N_15332,N_13699,N_13705);
or U15333 (N_15333,N_13251,N_13786);
and U15334 (N_15334,N_13363,N_14390);
or U15335 (N_15335,N_13819,N_13758);
xnor U15336 (N_15336,N_13344,N_13321);
nand U15337 (N_15337,N_14040,N_13301);
and U15338 (N_15338,N_13925,N_14255);
nor U15339 (N_15339,N_13876,N_13210);
and U15340 (N_15340,N_13790,N_14060);
and U15341 (N_15341,N_13465,N_13468);
xor U15342 (N_15342,N_13896,N_14301);
nor U15343 (N_15343,N_13261,N_13303);
and U15344 (N_15344,N_14093,N_14387);
or U15345 (N_15345,N_13361,N_13478);
or U15346 (N_15346,N_13897,N_14049);
nand U15347 (N_15347,N_13750,N_13615);
and U15348 (N_15348,N_14019,N_14143);
xnor U15349 (N_15349,N_13765,N_14231);
and U15350 (N_15350,N_13431,N_14346);
and U15351 (N_15351,N_13676,N_13300);
xor U15352 (N_15352,N_13997,N_14323);
or U15353 (N_15353,N_13308,N_13382);
xor U15354 (N_15354,N_13696,N_13257);
nand U15355 (N_15355,N_13241,N_13509);
and U15356 (N_15356,N_13993,N_13547);
nand U15357 (N_15357,N_14122,N_13551);
or U15358 (N_15358,N_13814,N_14227);
and U15359 (N_15359,N_13639,N_13914);
or U15360 (N_15360,N_14171,N_13756);
or U15361 (N_15361,N_13220,N_13431);
xor U15362 (N_15362,N_13827,N_13951);
nor U15363 (N_15363,N_13302,N_14294);
or U15364 (N_15364,N_13776,N_14025);
or U15365 (N_15365,N_13983,N_13222);
xnor U15366 (N_15366,N_13999,N_13978);
xor U15367 (N_15367,N_13765,N_13423);
nand U15368 (N_15368,N_13402,N_14138);
or U15369 (N_15369,N_13339,N_13366);
and U15370 (N_15370,N_13696,N_13403);
or U15371 (N_15371,N_14224,N_13320);
nand U15372 (N_15372,N_13808,N_13812);
nand U15373 (N_15373,N_13548,N_13398);
or U15374 (N_15374,N_13892,N_13657);
nor U15375 (N_15375,N_13947,N_13704);
xnor U15376 (N_15376,N_13215,N_13881);
nor U15377 (N_15377,N_13608,N_14355);
or U15378 (N_15378,N_13423,N_14238);
or U15379 (N_15379,N_14117,N_13342);
and U15380 (N_15380,N_13890,N_13824);
nor U15381 (N_15381,N_14350,N_13569);
nor U15382 (N_15382,N_13440,N_13966);
nor U15383 (N_15383,N_13590,N_13783);
nor U15384 (N_15384,N_14291,N_14262);
nor U15385 (N_15385,N_13304,N_13581);
nor U15386 (N_15386,N_13855,N_14324);
or U15387 (N_15387,N_13730,N_14323);
and U15388 (N_15388,N_13331,N_14171);
nand U15389 (N_15389,N_13393,N_13736);
nor U15390 (N_15390,N_14233,N_13898);
or U15391 (N_15391,N_13626,N_14270);
xnor U15392 (N_15392,N_14249,N_13429);
xor U15393 (N_15393,N_13561,N_13247);
nor U15394 (N_15394,N_13905,N_14366);
nor U15395 (N_15395,N_13353,N_13956);
nor U15396 (N_15396,N_13441,N_13752);
or U15397 (N_15397,N_13685,N_13294);
or U15398 (N_15398,N_13687,N_14388);
or U15399 (N_15399,N_13819,N_13845);
or U15400 (N_15400,N_14237,N_13854);
nor U15401 (N_15401,N_13750,N_13506);
and U15402 (N_15402,N_13713,N_13665);
nor U15403 (N_15403,N_13663,N_14003);
or U15404 (N_15404,N_14397,N_14240);
or U15405 (N_15405,N_14346,N_14383);
nor U15406 (N_15406,N_14095,N_13408);
nor U15407 (N_15407,N_14249,N_14168);
or U15408 (N_15408,N_13384,N_13485);
nand U15409 (N_15409,N_13713,N_13510);
xnor U15410 (N_15410,N_13572,N_13760);
xnor U15411 (N_15411,N_14006,N_13334);
or U15412 (N_15412,N_14045,N_13942);
xnor U15413 (N_15413,N_14068,N_14074);
nor U15414 (N_15414,N_13618,N_13447);
or U15415 (N_15415,N_14289,N_13805);
nor U15416 (N_15416,N_13793,N_13202);
xor U15417 (N_15417,N_13266,N_14025);
and U15418 (N_15418,N_13847,N_13297);
xnor U15419 (N_15419,N_14320,N_13360);
or U15420 (N_15420,N_14259,N_13573);
xnor U15421 (N_15421,N_13427,N_14007);
nand U15422 (N_15422,N_13617,N_13997);
xor U15423 (N_15423,N_13681,N_13465);
and U15424 (N_15424,N_13671,N_14058);
or U15425 (N_15425,N_13919,N_13532);
nand U15426 (N_15426,N_13395,N_14334);
nand U15427 (N_15427,N_13536,N_14163);
and U15428 (N_15428,N_13495,N_13406);
nand U15429 (N_15429,N_13912,N_14258);
or U15430 (N_15430,N_14323,N_14344);
and U15431 (N_15431,N_13573,N_14316);
nand U15432 (N_15432,N_13944,N_13625);
nand U15433 (N_15433,N_13341,N_13365);
or U15434 (N_15434,N_13763,N_14278);
xor U15435 (N_15435,N_14268,N_14301);
or U15436 (N_15436,N_13337,N_13396);
nand U15437 (N_15437,N_14140,N_14398);
and U15438 (N_15438,N_14368,N_13271);
or U15439 (N_15439,N_13447,N_13295);
or U15440 (N_15440,N_13345,N_14171);
or U15441 (N_15441,N_13639,N_13718);
nand U15442 (N_15442,N_14170,N_13561);
or U15443 (N_15443,N_14265,N_14054);
nor U15444 (N_15444,N_13208,N_13527);
and U15445 (N_15445,N_13731,N_13660);
and U15446 (N_15446,N_13612,N_13253);
xnor U15447 (N_15447,N_13585,N_14055);
or U15448 (N_15448,N_14380,N_13426);
or U15449 (N_15449,N_14289,N_13464);
or U15450 (N_15450,N_13681,N_14019);
nand U15451 (N_15451,N_13859,N_14107);
nand U15452 (N_15452,N_14141,N_13846);
and U15453 (N_15453,N_13489,N_13782);
nor U15454 (N_15454,N_13552,N_13610);
nand U15455 (N_15455,N_14205,N_13934);
or U15456 (N_15456,N_13601,N_13284);
nor U15457 (N_15457,N_13321,N_13304);
nor U15458 (N_15458,N_13363,N_13251);
or U15459 (N_15459,N_13752,N_13452);
or U15460 (N_15460,N_13505,N_13994);
or U15461 (N_15461,N_13233,N_13303);
xnor U15462 (N_15462,N_13472,N_13992);
nand U15463 (N_15463,N_14033,N_13620);
nor U15464 (N_15464,N_14125,N_14394);
nand U15465 (N_15465,N_14131,N_13972);
and U15466 (N_15466,N_14244,N_14252);
nand U15467 (N_15467,N_14052,N_13299);
xnor U15468 (N_15468,N_13907,N_13933);
nand U15469 (N_15469,N_13584,N_14040);
xor U15470 (N_15470,N_13387,N_13820);
nor U15471 (N_15471,N_13449,N_13648);
and U15472 (N_15472,N_13313,N_13880);
nor U15473 (N_15473,N_13250,N_13660);
nor U15474 (N_15474,N_13885,N_13778);
nand U15475 (N_15475,N_13321,N_13394);
nor U15476 (N_15476,N_13831,N_14316);
xnor U15477 (N_15477,N_13936,N_14380);
or U15478 (N_15478,N_13771,N_13630);
xor U15479 (N_15479,N_13513,N_13742);
nand U15480 (N_15480,N_13614,N_13621);
nor U15481 (N_15481,N_13610,N_13794);
xor U15482 (N_15482,N_13608,N_13491);
nand U15483 (N_15483,N_13662,N_13855);
or U15484 (N_15484,N_13512,N_14260);
and U15485 (N_15485,N_13895,N_13975);
and U15486 (N_15486,N_13677,N_13621);
nand U15487 (N_15487,N_13929,N_14284);
xnor U15488 (N_15488,N_14175,N_13657);
nand U15489 (N_15489,N_13517,N_14126);
xnor U15490 (N_15490,N_13879,N_14289);
or U15491 (N_15491,N_14233,N_13218);
or U15492 (N_15492,N_14178,N_13652);
and U15493 (N_15493,N_14233,N_13988);
xor U15494 (N_15494,N_13792,N_13269);
and U15495 (N_15495,N_13888,N_13728);
nand U15496 (N_15496,N_14351,N_14045);
nand U15497 (N_15497,N_13701,N_14290);
xor U15498 (N_15498,N_13300,N_13563);
nor U15499 (N_15499,N_14333,N_13744);
nor U15500 (N_15500,N_14357,N_13598);
nand U15501 (N_15501,N_14149,N_13502);
and U15502 (N_15502,N_14018,N_13279);
nor U15503 (N_15503,N_13769,N_13337);
xnor U15504 (N_15504,N_13952,N_13711);
nand U15505 (N_15505,N_13522,N_14009);
or U15506 (N_15506,N_14306,N_13908);
xor U15507 (N_15507,N_14309,N_13822);
nand U15508 (N_15508,N_14315,N_13442);
nand U15509 (N_15509,N_13241,N_13658);
and U15510 (N_15510,N_14062,N_13246);
nor U15511 (N_15511,N_13687,N_13610);
and U15512 (N_15512,N_14372,N_14356);
xor U15513 (N_15513,N_14336,N_13576);
and U15514 (N_15514,N_14035,N_13642);
nand U15515 (N_15515,N_14290,N_13367);
or U15516 (N_15516,N_14374,N_13325);
xnor U15517 (N_15517,N_14055,N_14007);
xor U15518 (N_15518,N_13241,N_13710);
xor U15519 (N_15519,N_14070,N_13636);
and U15520 (N_15520,N_13683,N_13868);
nand U15521 (N_15521,N_14257,N_14362);
nand U15522 (N_15522,N_13645,N_13341);
xor U15523 (N_15523,N_13448,N_14156);
xnor U15524 (N_15524,N_13314,N_14107);
or U15525 (N_15525,N_13998,N_13741);
nand U15526 (N_15526,N_14382,N_14044);
nand U15527 (N_15527,N_14240,N_13233);
or U15528 (N_15528,N_14066,N_13705);
or U15529 (N_15529,N_13406,N_13422);
or U15530 (N_15530,N_13251,N_13672);
and U15531 (N_15531,N_14231,N_13406);
or U15532 (N_15532,N_14280,N_14320);
and U15533 (N_15533,N_14198,N_14185);
or U15534 (N_15534,N_13573,N_13682);
nand U15535 (N_15535,N_14064,N_13421);
nor U15536 (N_15536,N_13489,N_13208);
nor U15537 (N_15537,N_13722,N_13494);
and U15538 (N_15538,N_13998,N_14223);
nand U15539 (N_15539,N_13254,N_13735);
nor U15540 (N_15540,N_14375,N_13532);
xnor U15541 (N_15541,N_13634,N_14359);
nand U15542 (N_15542,N_13549,N_13781);
and U15543 (N_15543,N_13523,N_13256);
and U15544 (N_15544,N_13589,N_13585);
nand U15545 (N_15545,N_13930,N_13497);
or U15546 (N_15546,N_14066,N_13382);
nor U15547 (N_15547,N_14389,N_13302);
nor U15548 (N_15548,N_13441,N_13528);
nor U15549 (N_15549,N_13306,N_14025);
nor U15550 (N_15550,N_13840,N_13969);
or U15551 (N_15551,N_13731,N_14331);
nor U15552 (N_15552,N_13252,N_13635);
xnor U15553 (N_15553,N_13778,N_13922);
nand U15554 (N_15554,N_13371,N_13361);
and U15555 (N_15555,N_13322,N_13728);
nand U15556 (N_15556,N_13579,N_14358);
or U15557 (N_15557,N_13610,N_13867);
nor U15558 (N_15558,N_13923,N_13419);
and U15559 (N_15559,N_13879,N_13981);
nor U15560 (N_15560,N_13977,N_13624);
nand U15561 (N_15561,N_13505,N_14028);
or U15562 (N_15562,N_14012,N_13786);
nor U15563 (N_15563,N_13891,N_14010);
xnor U15564 (N_15564,N_14336,N_13590);
nand U15565 (N_15565,N_14306,N_13920);
or U15566 (N_15566,N_14352,N_13268);
xnor U15567 (N_15567,N_13779,N_14250);
xor U15568 (N_15568,N_13754,N_14321);
nor U15569 (N_15569,N_13948,N_14062);
nor U15570 (N_15570,N_13225,N_13868);
nand U15571 (N_15571,N_14129,N_13530);
nor U15572 (N_15572,N_14044,N_14338);
nor U15573 (N_15573,N_13208,N_13989);
nor U15574 (N_15574,N_14140,N_13988);
nand U15575 (N_15575,N_13779,N_14219);
nor U15576 (N_15576,N_13263,N_14312);
nand U15577 (N_15577,N_13538,N_14185);
xor U15578 (N_15578,N_13372,N_14352);
xor U15579 (N_15579,N_14033,N_14290);
nor U15580 (N_15580,N_14317,N_14033);
nand U15581 (N_15581,N_14044,N_14074);
nor U15582 (N_15582,N_14154,N_13719);
or U15583 (N_15583,N_13707,N_13357);
nor U15584 (N_15584,N_13298,N_14141);
xnor U15585 (N_15585,N_13320,N_13777);
and U15586 (N_15586,N_14125,N_14031);
nand U15587 (N_15587,N_13244,N_13979);
nor U15588 (N_15588,N_14261,N_13771);
or U15589 (N_15589,N_13262,N_13728);
or U15590 (N_15590,N_14288,N_13826);
or U15591 (N_15591,N_13909,N_14269);
or U15592 (N_15592,N_13798,N_13595);
nand U15593 (N_15593,N_13220,N_13633);
xor U15594 (N_15594,N_13474,N_14256);
nand U15595 (N_15595,N_14191,N_14141);
or U15596 (N_15596,N_13956,N_14260);
and U15597 (N_15597,N_13266,N_13983);
nand U15598 (N_15598,N_13280,N_13339);
nor U15599 (N_15599,N_14307,N_13576);
or U15600 (N_15600,N_15373,N_14468);
or U15601 (N_15601,N_15176,N_15211);
and U15602 (N_15602,N_14875,N_15432);
or U15603 (N_15603,N_14976,N_15465);
nor U15604 (N_15604,N_14434,N_14848);
or U15605 (N_15605,N_14703,N_15345);
nand U15606 (N_15606,N_15040,N_14896);
or U15607 (N_15607,N_15573,N_14749);
xor U15608 (N_15608,N_15242,N_14564);
nand U15609 (N_15609,N_15082,N_15541);
or U15610 (N_15610,N_14442,N_14610);
nand U15611 (N_15611,N_14474,N_15291);
nor U15612 (N_15612,N_15116,N_15477);
nand U15613 (N_15613,N_14825,N_15275);
and U15614 (N_15614,N_14486,N_14781);
and U15615 (N_15615,N_15320,N_14722);
or U15616 (N_15616,N_15285,N_14518);
nand U15617 (N_15617,N_14786,N_14764);
nand U15618 (N_15618,N_14899,N_14915);
or U15619 (N_15619,N_14414,N_14601);
nand U15620 (N_15620,N_14403,N_15463);
or U15621 (N_15621,N_15129,N_15058);
xor U15622 (N_15622,N_14615,N_14517);
and U15623 (N_15623,N_15008,N_15219);
nand U15624 (N_15624,N_14579,N_15462);
or U15625 (N_15625,N_14589,N_15315);
xnor U15626 (N_15626,N_15046,N_15241);
and U15627 (N_15627,N_14478,N_15516);
xor U15628 (N_15628,N_14855,N_15073);
or U15629 (N_15629,N_15335,N_15287);
nand U15630 (N_15630,N_14943,N_14535);
nor U15631 (N_15631,N_15350,N_14646);
and U15632 (N_15632,N_14496,N_15153);
and U15633 (N_15633,N_14763,N_15507);
nand U15634 (N_15634,N_14778,N_15406);
nor U15635 (N_15635,N_14963,N_14955);
nand U15636 (N_15636,N_15221,N_15417);
or U15637 (N_15637,N_14485,N_14762);
xnor U15638 (N_15638,N_14631,N_15217);
xor U15639 (N_15639,N_14536,N_15007);
xnor U15640 (N_15640,N_15321,N_15124);
or U15641 (N_15641,N_14634,N_15513);
nand U15642 (N_15642,N_14920,N_14639);
or U15643 (N_15643,N_14682,N_14583);
xor U15644 (N_15644,N_14552,N_14887);
and U15645 (N_15645,N_14898,N_15254);
nor U15646 (N_15646,N_15182,N_15358);
or U15647 (N_15647,N_15147,N_15444);
nor U15648 (N_15648,N_15453,N_14572);
and U15649 (N_15649,N_14498,N_14569);
and U15650 (N_15650,N_14418,N_14904);
xnor U15651 (N_15651,N_14750,N_15024);
nor U15652 (N_15652,N_15202,N_14741);
nand U15653 (N_15653,N_14553,N_15538);
xnor U15654 (N_15654,N_14713,N_15426);
nor U15655 (N_15655,N_14939,N_14984);
xnor U15656 (N_15656,N_14982,N_14698);
and U15657 (N_15657,N_14416,N_15197);
nand U15658 (N_15658,N_14941,N_14542);
or U15659 (N_15659,N_15412,N_14958);
xnor U15660 (N_15660,N_15341,N_15314);
and U15661 (N_15661,N_15096,N_15488);
nand U15662 (N_15662,N_15000,N_15048);
nand U15663 (N_15663,N_15578,N_15105);
nor U15664 (N_15664,N_14765,N_15517);
nor U15665 (N_15665,N_14806,N_14754);
or U15666 (N_15666,N_14873,N_15244);
xor U15667 (N_15667,N_15141,N_14882);
nand U15668 (N_15668,N_14844,N_15092);
and U15669 (N_15669,N_15185,N_14706);
or U15670 (N_15670,N_14469,N_14566);
or U15671 (N_15671,N_15510,N_15121);
nand U15672 (N_15672,N_14475,N_15177);
or U15673 (N_15673,N_14483,N_15081);
and U15674 (N_15674,N_14895,N_15547);
or U15675 (N_15675,N_14885,N_14585);
or U15676 (N_15676,N_14949,N_15392);
xnor U15677 (N_15677,N_15187,N_14742);
nand U15678 (N_15678,N_14588,N_15130);
nand U15679 (N_15679,N_15173,N_14746);
and U15680 (N_15680,N_15554,N_15467);
xor U15681 (N_15681,N_14839,N_15257);
or U15682 (N_15682,N_14823,N_15296);
xor U15683 (N_15683,N_14555,N_14826);
or U15684 (N_15684,N_15284,N_14637);
or U15685 (N_15685,N_15163,N_15443);
and U15686 (N_15686,N_15482,N_14662);
nand U15687 (N_15687,N_14669,N_14780);
and U15688 (N_15688,N_14599,N_15190);
xnor U15689 (N_15689,N_14576,N_14803);
and U15690 (N_15690,N_14420,N_15133);
nor U15691 (N_15691,N_14423,N_15286);
and U15692 (N_15692,N_15340,N_15596);
or U15693 (N_15693,N_15001,N_14951);
and U15694 (N_15694,N_15599,N_14489);
nor U15695 (N_15695,N_15203,N_14507);
or U15696 (N_15696,N_15065,N_15037);
and U15697 (N_15697,N_14635,N_14683);
and U15698 (N_15698,N_15521,N_14602);
nand U15699 (N_15699,N_14559,N_14783);
nand U15700 (N_15700,N_14543,N_14604);
nand U15701 (N_15701,N_15260,N_15150);
nor U15702 (N_15702,N_15391,N_14511);
xor U15703 (N_15703,N_14852,N_14539);
nor U15704 (N_15704,N_15466,N_15589);
nor U15705 (N_15705,N_14573,N_15561);
nor U15706 (N_15706,N_14640,N_15272);
or U15707 (N_15707,N_15094,N_15123);
xnor U15708 (N_15708,N_15050,N_14522);
and U15709 (N_15709,N_14404,N_14849);
nand U15710 (N_15710,N_15175,N_14865);
nand U15711 (N_15711,N_14591,N_14837);
xor U15712 (N_15712,N_14642,N_14794);
nand U15713 (N_15713,N_15167,N_14932);
xnor U15714 (N_15714,N_15503,N_14651);
nor U15715 (N_15715,N_14558,N_15155);
xnor U15716 (N_15716,N_15414,N_15550);
nor U15717 (N_15717,N_15278,N_15383);
or U15718 (N_15718,N_15523,N_15290);
nand U15719 (N_15719,N_15549,N_14596);
or U15720 (N_15720,N_15586,N_15357);
xor U15721 (N_15721,N_14820,N_15354);
xor U15722 (N_15722,N_15128,N_14956);
and U15723 (N_15723,N_15394,N_14453);
nand U15724 (N_15724,N_15327,N_14436);
and U15725 (N_15725,N_14931,N_14718);
or U15726 (N_15726,N_15195,N_14748);
or U15727 (N_15727,N_15261,N_15558);
nand U15728 (N_15728,N_15498,N_14804);
nor U15729 (N_15729,N_15419,N_14678);
nor U15730 (N_15730,N_15085,N_14993);
nor U15731 (N_15731,N_14644,N_15434);
nor U15732 (N_15732,N_15119,N_14506);
and U15733 (N_15733,N_15288,N_15228);
and U15734 (N_15734,N_15399,N_14700);
and U15735 (N_15735,N_15071,N_15401);
xnor U15736 (N_15736,N_14648,N_14838);
nor U15737 (N_15737,N_15209,N_14740);
xor U15738 (N_15738,N_14992,N_14696);
nand U15739 (N_15739,N_14903,N_15583);
xor U15740 (N_15740,N_15464,N_15234);
nand U15741 (N_15741,N_14994,N_15424);
or U15742 (N_15742,N_14580,N_15371);
and U15743 (N_15743,N_14624,N_15556);
or U15744 (N_15744,N_15039,N_14711);
and U15745 (N_15745,N_15183,N_15049);
nor U15746 (N_15746,N_14789,N_14724);
nand U15747 (N_15747,N_14922,N_14461);
xnor U15748 (N_15748,N_14944,N_14505);
and U15749 (N_15749,N_15168,N_15070);
xor U15750 (N_15750,N_15405,N_15479);
nand U15751 (N_15751,N_14933,N_14617);
nand U15752 (N_15752,N_14728,N_15515);
and U15753 (N_15753,N_15415,N_15375);
nor U15754 (N_15754,N_15423,N_14488);
nor U15755 (N_15755,N_15529,N_15527);
or U15756 (N_15756,N_14704,N_14534);
or U15757 (N_15757,N_15107,N_15029);
or U15758 (N_15758,N_14457,N_14888);
and U15759 (N_15759,N_14914,N_14614);
nand U15760 (N_15760,N_15109,N_14495);
nand U15761 (N_15761,N_15362,N_15470);
xor U15762 (N_15762,N_15156,N_14638);
nand U15763 (N_15763,N_15233,N_14772);
nor U15764 (N_15764,N_15098,N_15279);
nand U15765 (N_15765,N_14695,N_14738);
nand U15766 (N_15766,N_15273,N_15252);
nand U15767 (N_15767,N_15258,N_15575);
or U15768 (N_15768,N_14435,N_15369);
nor U15769 (N_15769,N_15186,N_15553);
xor U15770 (N_15770,N_15250,N_14426);
nand U15771 (N_15771,N_14877,N_14481);
xnor U15772 (N_15772,N_14432,N_15179);
xor U15773 (N_15773,N_15522,N_14867);
nor U15774 (N_15774,N_14890,N_15367);
xnor U15775 (N_15775,N_15011,N_14857);
nor U15776 (N_15776,N_14608,N_14680);
nor U15777 (N_15777,N_14894,N_14541);
nand U15778 (N_15778,N_14981,N_14611);
nor U15779 (N_15779,N_15565,N_15091);
nor U15780 (N_15780,N_15162,N_14758);
and U15781 (N_15781,N_14815,N_15161);
nand U15782 (N_15782,N_14940,N_15044);
or U15783 (N_15783,N_15034,N_14902);
nor U15784 (N_15784,N_15454,N_14729);
or U15785 (N_15785,N_15594,N_15068);
and U15786 (N_15786,N_14814,N_15393);
or U15787 (N_15787,N_14441,N_15243);
xnor U15788 (N_15788,N_14942,N_15389);
or U15789 (N_15789,N_14986,N_15120);
or U15790 (N_15790,N_14437,N_15269);
nand U15791 (N_15791,N_14630,N_15416);
xnor U15792 (N_15792,N_14716,N_15570);
nand U15793 (N_15793,N_15265,N_15206);
nand U15794 (N_15794,N_14925,N_15230);
or U15795 (N_15795,N_15118,N_14664);
or U15796 (N_15796,N_15385,N_14900);
and U15797 (N_15797,N_14968,N_15598);
nand U15798 (N_15798,N_14514,N_15022);
and U15799 (N_15799,N_14901,N_15200);
nor U15800 (N_15800,N_15543,N_14653);
or U15801 (N_15801,N_15418,N_14633);
and U15802 (N_15802,N_15563,N_15164);
and U15803 (N_15803,N_15125,N_15095);
nor U15804 (N_15804,N_14590,N_14733);
and U15805 (N_15805,N_15440,N_14979);
and U15806 (N_15806,N_14800,N_14528);
nand U15807 (N_15807,N_14473,N_15456);
and U15808 (N_15808,N_14603,N_15475);
nor U15809 (N_15809,N_14419,N_15528);
xnor U15810 (N_15810,N_15409,N_15351);
nand U15811 (N_15811,N_14626,N_15555);
nand U15812 (N_15812,N_14813,N_15216);
xnor U15813 (N_15813,N_14476,N_15152);
nand U15814 (N_15814,N_14757,N_15113);
or U15815 (N_15815,N_15264,N_15582);
or U15816 (N_15816,N_15500,N_14516);
and U15817 (N_15817,N_15572,N_15038);
nand U15818 (N_15818,N_15458,N_15525);
or U15819 (N_15819,N_15237,N_14582);
xor U15820 (N_15820,N_14752,N_15526);
nor U15821 (N_15821,N_14797,N_15436);
and U15822 (N_15822,N_15455,N_15592);
or U15823 (N_15823,N_14801,N_15222);
and U15824 (N_15824,N_15089,N_14714);
or U15825 (N_15825,N_14685,N_15126);
xor U15826 (N_15826,N_15192,N_14874);
or U15827 (N_15827,N_14946,N_14934);
nand U15828 (N_15828,N_15518,N_14592);
and U15829 (N_15829,N_14753,N_14410);
xnor U15830 (N_15830,N_15535,N_14451);
xnor U15831 (N_15831,N_15043,N_15097);
xor U15832 (N_15832,N_14684,N_14759);
xnor U15833 (N_15833,N_15398,N_14532);
nand U15834 (N_15834,N_15430,N_15238);
or U15835 (N_15835,N_14405,N_15472);
xnor U15836 (N_15836,N_14647,N_15122);
nand U15837 (N_15837,N_14866,N_15359);
xor U15838 (N_15838,N_14798,N_14551);
nor U15839 (N_15839,N_15569,N_15093);
or U15840 (N_15840,N_14828,N_15353);
or U15841 (N_15841,N_15019,N_14889);
or U15842 (N_15842,N_14812,N_15157);
nand U15843 (N_15843,N_14808,N_15449);
or U15844 (N_15844,N_14538,N_15086);
nand U15845 (N_15845,N_14973,N_14492);
nor U15846 (N_15846,N_14509,N_15337);
or U15847 (N_15847,N_14502,N_15016);
nand U15848 (N_15848,N_15380,N_15326);
xnor U15849 (N_15849,N_14690,N_14650);
or U15850 (N_15850,N_14621,N_14479);
or U15851 (N_15851,N_15407,N_15002);
or U15852 (N_15852,N_15087,N_15356);
xor U15853 (N_15853,N_15307,N_15208);
xnor U15854 (N_15854,N_15239,N_15344);
nand U15855 (N_15855,N_14594,N_15442);
nor U15856 (N_15856,N_15052,N_15493);
xnor U15857 (N_15857,N_15413,N_15194);
nand U15858 (N_15858,N_15319,N_15481);
nor U15859 (N_15859,N_15331,N_14428);
xnor U15860 (N_15860,N_14667,N_14744);
nand U15861 (N_15861,N_14760,N_14666);
nor U15862 (N_15862,N_15127,N_15559);
or U15863 (N_15863,N_15274,N_14770);
and U15864 (N_15864,N_14671,N_15342);
xor U15865 (N_15865,N_14484,N_15310);
and U15866 (N_15866,N_14447,N_14600);
nor U15867 (N_15867,N_14872,N_15114);
nand U15868 (N_15868,N_15251,N_14842);
or U15869 (N_15869,N_14605,N_15499);
nand U15870 (N_15870,N_15303,N_15139);
and U15871 (N_15871,N_14415,N_15312);
nor U15872 (N_15872,N_15247,N_14980);
nor U15873 (N_15873,N_14512,N_15577);
nor U15874 (N_15874,N_14997,N_15336);
and U15875 (N_15875,N_14701,N_15159);
xor U15876 (N_15876,N_14878,N_14493);
or U15877 (N_15877,N_14454,N_15178);
xnor U15878 (N_15878,N_14715,N_15504);
and U15879 (N_15879,N_15408,N_14673);
nor U15880 (N_15880,N_14577,N_15020);
xor U15881 (N_15881,N_15519,N_14990);
nand U15882 (N_15882,N_15390,N_14452);
and U15883 (N_15883,N_14412,N_15451);
or U15884 (N_15884,N_14989,N_14521);
xor U15885 (N_15885,N_15104,N_14830);
xnor U15886 (N_15886,N_14988,N_15361);
nor U15887 (N_15887,N_15143,N_14991);
nor U15888 (N_15888,N_15474,N_14726);
and U15889 (N_15889,N_15520,N_14999);
xnor U15890 (N_15890,N_14995,N_15539);
or U15891 (N_15891,N_15425,N_15402);
nand U15892 (N_15892,N_14723,N_14679);
nor U15893 (N_15893,N_15196,N_15584);
xor U15894 (N_15894,N_14871,N_15154);
nand U15895 (N_15895,N_14969,N_15255);
or U15896 (N_15896,N_14730,N_15064);
and U15897 (N_15897,N_14840,N_14560);
and U15898 (N_15898,N_15138,N_14709);
nand U15899 (N_15899,N_15289,N_14627);
and U15900 (N_15900,N_14431,N_14775);
nor U15901 (N_15901,N_14549,N_14455);
xnor U15902 (N_15902,N_15485,N_15591);
nor U15903 (N_15903,N_15329,N_15439);
or U15904 (N_15904,N_15339,N_14965);
xnor U15905 (N_15905,N_15566,N_14921);
nand U15906 (N_15906,N_15226,N_14776);
nand U15907 (N_15907,N_14503,N_14408);
or U15908 (N_15908,N_15075,N_14557);
nor U15909 (N_15909,N_14571,N_14854);
nand U15910 (N_15910,N_14439,N_14523);
nand U15911 (N_15911,N_14876,N_14919);
nor U15912 (N_15912,N_15428,N_15056);
nand U15913 (N_15913,N_14927,N_15484);
or U15914 (N_15914,N_14743,N_15099);
nand U15915 (N_15915,N_14520,N_14905);
nand U15916 (N_15916,N_14501,N_14923);
xor U15917 (N_15917,N_14649,N_14924);
and U15918 (N_15918,N_14846,N_14545);
or U15919 (N_15919,N_15033,N_15171);
and U15920 (N_15920,N_14659,N_15397);
xnor U15921 (N_15921,N_14612,N_15343);
or U15922 (N_15922,N_15077,N_14425);
nand U15923 (N_15923,N_14427,N_15386);
nand U15924 (N_15924,N_15188,N_15246);
nand U15925 (N_15925,N_15292,N_14938);
or U15926 (N_15926,N_15452,N_14712);
and U15927 (N_15927,N_14401,N_14850);
nand U15928 (N_15928,N_14891,N_15079);
nand U15929 (N_15929,N_15060,N_15268);
nor U15930 (N_15930,N_15459,N_15468);
nand U15931 (N_15931,N_14836,N_14529);
and U15932 (N_15932,N_15142,N_15372);
or U15933 (N_15933,N_15595,N_14777);
xnor U15934 (N_15934,N_14450,N_15324);
and U15935 (N_15935,N_14856,N_14767);
and U15936 (N_15936,N_14544,N_15382);
and U15937 (N_15937,N_14864,N_15169);
xor U15938 (N_15938,N_14471,N_14996);
xnor U15939 (N_15939,N_14827,N_15030);
nand U15940 (N_15940,N_15445,N_15384);
nor U15941 (N_15941,N_14953,N_14761);
and U15942 (N_15942,N_15325,N_15478);
nor U15943 (N_15943,N_14459,N_14411);
and U15944 (N_15944,N_15067,N_15266);
or U15945 (N_15945,N_15593,N_14935);
nor U15946 (N_15946,N_15562,N_15213);
xor U15947 (N_15947,N_14625,N_15524);
nand U15948 (N_15948,N_15387,N_14952);
nand U15949 (N_15949,N_15009,N_15042);
xor U15950 (N_15950,N_15542,N_14717);
xnor U15951 (N_15951,N_15035,N_14655);
nand U15952 (N_15952,N_15259,N_15302);
and U15953 (N_15953,N_14769,N_15021);
and U15954 (N_15954,N_14689,N_14834);
nand U15955 (N_15955,N_15587,N_15015);
nor U15956 (N_15956,N_15552,N_14472);
and U15957 (N_15957,N_14672,N_14540);
nand U15958 (N_15958,N_15207,N_14790);
xor U15959 (N_15959,N_15568,N_14402);
and U15960 (N_15960,N_15437,N_14818);
or U15961 (N_15961,N_14929,N_14570);
nand U15962 (N_15962,N_14816,N_14508);
nand U15963 (N_15963,N_14609,N_15347);
and U15964 (N_15964,N_15400,N_15501);
or U15965 (N_15965,N_14597,N_15533);
or U15966 (N_15966,N_15505,N_14500);
and U15967 (N_15967,N_14692,N_15306);
and U15968 (N_15968,N_15537,N_15311);
nand U15969 (N_15969,N_14641,N_14430);
xor U15970 (N_15970,N_15318,N_15263);
xnor U15971 (N_15971,N_15532,N_14708);
nor U15972 (N_15972,N_14616,N_14499);
and U15973 (N_15973,N_14623,N_15294);
and U15974 (N_15974,N_15111,N_14413);
xor U15975 (N_15975,N_15088,N_15365);
xor U15976 (N_15976,N_14598,N_15486);
xnor U15977 (N_15977,N_14490,N_14406);
nand U15978 (N_15978,N_15205,N_15483);
and U15979 (N_15979,N_14792,N_15055);
nand U15980 (N_15980,N_14530,N_15395);
and U15981 (N_15981,N_15476,N_15283);
and U15982 (N_15982,N_15134,N_15232);
xnor U15983 (N_15983,N_15313,N_15349);
and U15984 (N_15984,N_15193,N_15054);
or U15985 (N_15985,N_15223,N_14661);
xor U15986 (N_15986,N_14527,N_15026);
nor U15987 (N_15987,N_14721,N_14697);
nor U15988 (N_15988,N_15023,N_14556);
xnor U15989 (N_15989,N_14421,N_14853);
nand U15990 (N_15990,N_15166,N_15487);
or U15991 (N_15991,N_14799,N_15041);
xnor U15992 (N_15992,N_14835,N_14586);
or U15993 (N_15993,N_14652,N_14510);
nand U15994 (N_15994,N_15446,N_15191);
nand U15995 (N_15995,N_15429,N_14702);
nand U15996 (N_15996,N_15297,N_15551);
nand U15997 (N_15997,N_15366,N_14862);
or U15998 (N_15998,N_15253,N_14824);
and U15999 (N_15999,N_14467,N_14491);
nand U16000 (N_16000,N_14618,N_15227);
or U16001 (N_16001,N_15374,N_14936);
xor U16002 (N_16002,N_15597,N_15579);
nand U16003 (N_16003,N_14851,N_15069);
nand U16004 (N_16004,N_14613,N_14732);
nand U16005 (N_16005,N_15571,N_14802);
and U16006 (N_16006,N_14668,N_14676);
xor U16007 (N_16007,N_14705,N_15180);
nor U16008 (N_16008,N_15005,N_14575);
nand U16009 (N_16009,N_15108,N_14884);
nand U16010 (N_16010,N_14462,N_14443);
nand U16011 (N_16011,N_15045,N_15184);
and U16012 (N_16012,N_14805,N_15028);
nand U16013 (N_16013,N_15492,N_15495);
nand U16014 (N_16014,N_14694,N_14911);
or U16015 (N_16015,N_14962,N_15115);
or U16016 (N_16016,N_14907,N_15376);
xnor U16017 (N_16017,N_14526,N_15170);
or U16018 (N_16018,N_14636,N_14918);
or U16019 (N_16019,N_14464,N_15461);
and U16020 (N_16020,N_14998,N_14561);
nor U16021 (N_16021,N_14987,N_15160);
xnor U16022 (N_16022,N_15047,N_14847);
xor U16023 (N_16023,N_14893,N_15144);
nand U16024 (N_16024,N_14807,N_15214);
or U16025 (N_16025,N_15172,N_14975);
nand U16026 (N_16026,N_15131,N_14658);
xnor U16027 (N_16027,N_14913,N_15072);
and U16028 (N_16028,N_15305,N_14819);
and U16029 (N_16029,N_14565,N_14587);
nand U16030 (N_16030,N_14784,N_15427);
or U16031 (N_16031,N_15420,N_15013);
nand U16032 (N_16032,N_14886,N_14463);
and U16033 (N_16033,N_15006,N_14691);
and U16034 (N_16034,N_15236,N_14710);
nand U16035 (N_16035,N_15564,N_15078);
nand U16036 (N_16036,N_15003,N_14881);
nand U16037 (N_16037,N_14967,N_15531);
or U16038 (N_16038,N_15480,N_14945);
xor U16039 (N_16039,N_14869,N_14497);
xnor U16040 (N_16040,N_14880,N_15514);
and U16041 (N_16041,N_15363,N_15580);
and U16042 (N_16042,N_14548,N_14438);
nor U16043 (N_16043,N_14859,N_14458);
nor U16044 (N_16044,N_14964,N_15585);
xor U16045 (N_16045,N_14957,N_15063);
xnor U16046 (N_16046,N_14688,N_15433);
xnor U16047 (N_16047,N_14832,N_15212);
nor U16048 (N_16048,N_15100,N_14916);
nor U16049 (N_16049,N_14687,N_15330);
xor U16050 (N_16050,N_15025,N_14845);
or U16051 (N_16051,N_15074,N_15112);
nand U16052 (N_16052,N_14657,N_14550);
or U16053 (N_16053,N_15328,N_15377);
xor U16054 (N_16054,N_15332,N_15083);
xnor U16055 (N_16055,N_14947,N_14959);
nor U16056 (N_16056,N_14567,N_14595);
nand U16057 (N_16057,N_14897,N_15145);
or U16058 (N_16058,N_14407,N_15323);
nor U16059 (N_16059,N_14656,N_15084);
xnor U16060 (N_16060,N_14966,N_15027);
xnor U16061 (N_16061,N_14654,N_15061);
nor U16062 (N_16062,N_15422,N_15245);
and U16063 (N_16063,N_14670,N_15352);
nand U16064 (N_16064,N_14515,N_15136);
xnor U16065 (N_16065,N_15370,N_14863);
or U16066 (N_16066,N_14831,N_15224);
or U16067 (N_16067,N_14645,N_14779);
nor U16068 (N_16068,N_14793,N_14768);
nand U16069 (N_16069,N_15189,N_14525);
nor U16070 (N_16070,N_14906,N_14477);
xor U16071 (N_16071,N_15544,N_14970);
and U16072 (N_16072,N_14628,N_15066);
or U16073 (N_16073,N_14465,N_14607);
nor U16074 (N_16074,N_14568,N_14796);
or U16075 (N_16075,N_15299,N_15548);
nor U16076 (N_16076,N_14547,N_15014);
nand U16077 (N_16077,N_15322,N_14504);
xnor U16078 (N_16078,N_14909,N_14449);
and U16079 (N_16079,N_14821,N_14974);
and U16080 (N_16080,N_15431,N_14870);
xnor U16081 (N_16081,N_14751,N_15102);
nand U16082 (N_16082,N_15421,N_15057);
xnor U16083 (N_16083,N_14699,N_15298);
nor U16084 (N_16084,N_14487,N_14785);
and U16085 (N_16085,N_15018,N_15300);
nor U16086 (N_16086,N_14937,N_15103);
and U16087 (N_16087,N_14861,N_15502);
nand U16088 (N_16088,N_15262,N_15010);
and U16089 (N_16089,N_14677,N_14731);
xnor U16090 (N_16090,N_15165,N_15101);
and U16091 (N_16091,N_14409,N_15174);
xor U16092 (N_16092,N_14480,N_15140);
nand U16093 (N_16093,N_14822,N_15457);
nand U16094 (N_16094,N_14727,N_15581);
or U16095 (N_16095,N_14737,N_15218);
nand U16096 (N_16096,N_15270,N_14892);
and U16097 (N_16097,N_15447,N_15545);
and U16098 (N_16098,N_14795,N_15567);
xnor U16099 (N_16099,N_14440,N_15295);
xor U16100 (N_16100,N_14494,N_15316);
nand U16101 (N_16101,N_15388,N_14766);
nand U16102 (N_16102,N_15355,N_14810);
nand U16103 (N_16103,N_15309,N_14554);
nor U16104 (N_16104,N_15198,N_14574);
and U16105 (N_16105,N_14843,N_15496);
xor U16106 (N_16106,N_14971,N_15508);
or U16107 (N_16107,N_14643,N_15364);
and U16108 (N_16108,N_15036,N_14928);
nor U16109 (N_16109,N_15546,N_14466);
nor U16110 (N_16110,N_14524,N_15151);
xor U16111 (N_16111,N_14581,N_15450);
xnor U16112 (N_16112,N_15225,N_15530);
or U16113 (N_16113,N_14665,N_14829);
nand U16114 (N_16114,N_15158,N_15491);
xor U16115 (N_16115,N_15490,N_15338);
nor U16116 (N_16116,N_14429,N_14620);
and U16117 (N_16117,N_15333,N_15090);
or U16118 (N_16118,N_15199,N_15053);
nor U16119 (N_16119,N_15281,N_15012);
and U16120 (N_16120,N_15110,N_15137);
nor U16121 (N_16121,N_15215,N_15201);
and U16122 (N_16122,N_14584,N_15249);
or U16123 (N_16123,N_14433,N_15004);
xnor U16124 (N_16124,N_15438,N_15511);
and U16125 (N_16125,N_15560,N_14860);
or U16126 (N_16126,N_15441,N_14448);
and U16127 (N_16127,N_14629,N_14622);
and U16128 (N_16128,N_15435,N_15379);
or U16129 (N_16129,N_14456,N_14739);
or U16130 (N_16130,N_14417,N_14563);
and U16131 (N_16131,N_15210,N_14446);
and U16132 (N_16132,N_14735,N_14632);
and U16133 (N_16133,N_15235,N_14858);
nor U16134 (N_16134,N_14562,N_14424);
and U16135 (N_16135,N_15017,N_15059);
or U16136 (N_16136,N_15080,N_15277);
nand U16137 (N_16137,N_14791,N_15360);
and U16138 (N_16138,N_15146,N_15106);
and U16139 (N_16139,N_15301,N_15031);
or U16140 (N_16140,N_14720,N_14745);
nor U16141 (N_16141,N_15509,N_15368);
or U16142 (N_16142,N_14736,N_15132);
nor U16143 (N_16143,N_15381,N_15220);
xor U16144 (N_16144,N_14908,N_14978);
nor U16145 (N_16145,N_15334,N_14985);
and U16146 (N_16146,N_15256,N_14771);
and U16147 (N_16147,N_14930,N_15181);
nor U16148 (N_16148,N_14533,N_15473);
and U16149 (N_16149,N_14725,N_15494);
xor U16150 (N_16150,N_14681,N_14948);
and U16151 (N_16151,N_15231,N_15346);
nor U16152 (N_16152,N_15512,N_14674);
or U16153 (N_16153,N_15348,N_15506);
or U16154 (N_16154,N_14833,N_14531);
nor U16155 (N_16155,N_15588,N_15135);
nand U16156 (N_16156,N_14841,N_14606);
nor U16157 (N_16157,N_14954,N_14513);
nand U16158 (N_16158,N_14593,N_14912);
or U16159 (N_16159,N_15317,N_15471);
xor U16160 (N_16160,N_15149,N_15276);
nand U16161 (N_16161,N_14546,N_15148);
nor U16162 (N_16162,N_15576,N_14755);
or U16163 (N_16163,N_15117,N_14950);
or U16164 (N_16164,N_15469,N_15076);
nand U16165 (N_16165,N_15304,N_14961);
nand U16166 (N_16166,N_14707,N_14926);
or U16167 (N_16167,N_15411,N_15557);
xnor U16168 (N_16168,N_14868,N_15204);
nand U16169 (N_16169,N_14460,N_15540);
or U16170 (N_16170,N_14811,N_15534);
and U16171 (N_16171,N_15403,N_15051);
and U16172 (N_16172,N_14444,N_14470);
nor U16173 (N_16173,N_15590,N_15448);
xor U16174 (N_16174,N_14660,N_14519);
nand U16175 (N_16175,N_14482,N_14972);
xor U16176 (N_16176,N_14537,N_15280);
nand U16177 (N_16177,N_14809,N_14663);
nand U16178 (N_16178,N_14787,N_15282);
xor U16179 (N_16179,N_15267,N_15308);
nor U16180 (N_16180,N_14422,N_15062);
xor U16181 (N_16181,N_15410,N_15396);
nand U16182 (N_16182,N_15404,N_14578);
nand U16183 (N_16183,N_14719,N_15229);
nor U16184 (N_16184,N_15271,N_14734);
xnor U16185 (N_16185,N_14756,N_15378);
or U16186 (N_16186,N_15240,N_14774);
nand U16187 (N_16187,N_15536,N_14445);
xor U16188 (N_16188,N_14910,N_15032);
and U16189 (N_16189,N_14400,N_15497);
and U16190 (N_16190,N_14619,N_14693);
xnor U16191 (N_16191,N_14883,N_14675);
and U16192 (N_16192,N_15460,N_14788);
xnor U16193 (N_16193,N_14817,N_15293);
and U16194 (N_16194,N_14782,N_14917);
and U16195 (N_16195,N_15248,N_15489);
nor U16196 (N_16196,N_14879,N_15574);
or U16197 (N_16197,N_14977,N_14747);
nand U16198 (N_16198,N_14983,N_14960);
or U16199 (N_16199,N_14773,N_14686);
or U16200 (N_16200,N_15145,N_14438);
nand U16201 (N_16201,N_15153,N_14909);
xnor U16202 (N_16202,N_14871,N_14446);
or U16203 (N_16203,N_15291,N_14530);
xnor U16204 (N_16204,N_15364,N_14695);
xnor U16205 (N_16205,N_15162,N_14797);
nand U16206 (N_16206,N_14677,N_14711);
xor U16207 (N_16207,N_14433,N_15081);
and U16208 (N_16208,N_15200,N_15550);
nand U16209 (N_16209,N_15046,N_15544);
and U16210 (N_16210,N_15355,N_14443);
nand U16211 (N_16211,N_15574,N_14977);
nor U16212 (N_16212,N_15206,N_15091);
and U16213 (N_16213,N_15031,N_14590);
and U16214 (N_16214,N_14894,N_14846);
nor U16215 (N_16215,N_15286,N_15143);
xnor U16216 (N_16216,N_14887,N_14845);
nand U16217 (N_16217,N_15441,N_14695);
xor U16218 (N_16218,N_14522,N_14438);
xor U16219 (N_16219,N_15287,N_15518);
nand U16220 (N_16220,N_14955,N_15493);
xnor U16221 (N_16221,N_14709,N_14644);
nor U16222 (N_16222,N_14967,N_15314);
xor U16223 (N_16223,N_15417,N_14845);
or U16224 (N_16224,N_15519,N_14418);
xor U16225 (N_16225,N_15552,N_15427);
xor U16226 (N_16226,N_15104,N_14875);
xnor U16227 (N_16227,N_15218,N_15485);
or U16228 (N_16228,N_15053,N_14516);
nand U16229 (N_16229,N_14655,N_14960);
or U16230 (N_16230,N_14450,N_15022);
nand U16231 (N_16231,N_14452,N_15554);
and U16232 (N_16232,N_14576,N_15260);
or U16233 (N_16233,N_15506,N_14784);
xor U16234 (N_16234,N_15147,N_15457);
or U16235 (N_16235,N_14862,N_14478);
nand U16236 (N_16236,N_15253,N_15053);
or U16237 (N_16237,N_15248,N_14497);
and U16238 (N_16238,N_15053,N_14850);
nand U16239 (N_16239,N_15117,N_15095);
nor U16240 (N_16240,N_15271,N_15462);
xnor U16241 (N_16241,N_15349,N_15529);
xnor U16242 (N_16242,N_14853,N_15223);
nor U16243 (N_16243,N_14918,N_15202);
and U16244 (N_16244,N_15476,N_15237);
nand U16245 (N_16245,N_14553,N_14712);
or U16246 (N_16246,N_15025,N_14796);
and U16247 (N_16247,N_15142,N_14773);
nand U16248 (N_16248,N_15268,N_15037);
nor U16249 (N_16249,N_15509,N_15128);
xor U16250 (N_16250,N_15264,N_14921);
nand U16251 (N_16251,N_15433,N_14772);
nand U16252 (N_16252,N_14946,N_14414);
and U16253 (N_16253,N_15289,N_14691);
xor U16254 (N_16254,N_15274,N_15081);
nand U16255 (N_16255,N_15330,N_15498);
and U16256 (N_16256,N_15199,N_15465);
nor U16257 (N_16257,N_15067,N_14799);
xor U16258 (N_16258,N_15373,N_15390);
xor U16259 (N_16259,N_15453,N_15429);
or U16260 (N_16260,N_14557,N_15164);
or U16261 (N_16261,N_14581,N_14663);
nor U16262 (N_16262,N_15205,N_14758);
or U16263 (N_16263,N_14455,N_14786);
and U16264 (N_16264,N_14478,N_14709);
and U16265 (N_16265,N_15201,N_14411);
and U16266 (N_16266,N_14994,N_14959);
nand U16267 (N_16267,N_15484,N_14549);
or U16268 (N_16268,N_15192,N_14568);
xor U16269 (N_16269,N_14922,N_15386);
or U16270 (N_16270,N_14616,N_14454);
and U16271 (N_16271,N_14908,N_15277);
or U16272 (N_16272,N_15252,N_14895);
nor U16273 (N_16273,N_15206,N_15038);
nor U16274 (N_16274,N_15181,N_14796);
nor U16275 (N_16275,N_15592,N_14800);
nand U16276 (N_16276,N_15562,N_14782);
nand U16277 (N_16277,N_14583,N_15336);
and U16278 (N_16278,N_15352,N_15520);
or U16279 (N_16279,N_15019,N_15163);
nor U16280 (N_16280,N_15578,N_14602);
or U16281 (N_16281,N_15415,N_14825);
and U16282 (N_16282,N_15282,N_15215);
nand U16283 (N_16283,N_14522,N_15374);
nand U16284 (N_16284,N_15591,N_14974);
nor U16285 (N_16285,N_15493,N_15072);
or U16286 (N_16286,N_15258,N_14484);
nand U16287 (N_16287,N_14992,N_14408);
nor U16288 (N_16288,N_14768,N_15197);
xor U16289 (N_16289,N_15432,N_15429);
xnor U16290 (N_16290,N_15366,N_15191);
xnor U16291 (N_16291,N_14760,N_14813);
and U16292 (N_16292,N_14743,N_15361);
xnor U16293 (N_16293,N_14996,N_14549);
and U16294 (N_16294,N_15040,N_15224);
and U16295 (N_16295,N_14990,N_14772);
nor U16296 (N_16296,N_15435,N_15522);
or U16297 (N_16297,N_15519,N_14712);
nor U16298 (N_16298,N_15522,N_14996);
or U16299 (N_16299,N_15053,N_14678);
nand U16300 (N_16300,N_14568,N_14755);
and U16301 (N_16301,N_14908,N_15189);
or U16302 (N_16302,N_14940,N_15331);
nand U16303 (N_16303,N_15260,N_15563);
or U16304 (N_16304,N_15050,N_14610);
nor U16305 (N_16305,N_14428,N_15069);
nand U16306 (N_16306,N_15228,N_14958);
xor U16307 (N_16307,N_15359,N_14638);
nor U16308 (N_16308,N_15385,N_14520);
or U16309 (N_16309,N_15484,N_14922);
or U16310 (N_16310,N_15496,N_14726);
and U16311 (N_16311,N_14483,N_15464);
and U16312 (N_16312,N_15206,N_14607);
nand U16313 (N_16313,N_15281,N_15259);
nand U16314 (N_16314,N_15072,N_14946);
and U16315 (N_16315,N_14671,N_15229);
nand U16316 (N_16316,N_14984,N_14757);
or U16317 (N_16317,N_15468,N_15023);
xor U16318 (N_16318,N_14751,N_15495);
and U16319 (N_16319,N_15557,N_14472);
nor U16320 (N_16320,N_15391,N_14859);
or U16321 (N_16321,N_15047,N_15109);
xnor U16322 (N_16322,N_14441,N_15100);
nor U16323 (N_16323,N_14819,N_15564);
nor U16324 (N_16324,N_15449,N_14463);
xor U16325 (N_16325,N_14550,N_14684);
nor U16326 (N_16326,N_14699,N_15282);
or U16327 (N_16327,N_15007,N_15184);
nand U16328 (N_16328,N_14410,N_14669);
and U16329 (N_16329,N_15140,N_15424);
nor U16330 (N_16330,N_15168,N_14741);
nor U16331 (N_16331,N_14641,N_14927);
nand U16332 (N_16332,N_15576,N_14516);
nor U16333 (N_16333,N_15508,N_14726);
and U16334 (N_16334,N_15491,N_15311);
nand U16335 (N_16335,N_14915,N_15535);
nor U16336 (N_16336,N_15024,N_14916);
nand U16337 (N_16337,N_15457,N_15383);
and U16338 (N_16338,N_14400,N_15213);
or U16339 (N_16339,N_15596,N_14490);
and U16340 (N_16340,N_15470,N_14718);
xor U16341 (N_16341,N_14488,N_15335);
xnor U16342 (N_16342,N_14522,N_14747);
and U16343 (N_16343,N_14452,N_14868);
nand U16344 (N_16344,N_14982,N_15319);
and U16345 (N_16345,N_15486,N_15561);
xnor U16346 (N_16346,N_15084,N_14511);
and U16347 (N_16347,N_15334,N_15584);
and U16348 (N_16348,N_15080,N_14597);
nor U16349 (N_16349,N_14401,N_15070);
xor U16350 (N_16350,N_14941,N_14643);
xor U16351 (N_16351,N_15540,N_15393);
xnor U16352 (N_16352,N_15484,N_14997);
and U16353 (N_16353,N_15085,N_14845);
xnor U16354 (N_16354,N_15054,N_14499);
and U16355 (N_16355,N_15380,N_15323);
nand U16356 (N_16356,N_15110,N_14846);
and U16357 (N_16357,N_14435,N_14407);
or U16358 (N_16358,N_15010,N_15376);
nand U16359 (N_16359,N_15393,N_14657);
or U16360 (N_16360,N_14669,N_15074);
nor U16361 (N_16361,N_14814,N_15160);
nor U16362 (N_16362,N_15141,N_15265);
or U16363 (N_16363,N_14945,N_14730);
or U16364 (N_16364,N_15345,N_15330);
and U16365 (N_16365,N_15533,N_15397);
xnor U16366 (N_16366,N_14985,N_14473);
nor U16367 (N_16367,N_14606,N_15486);
or U16368 (N_16368,N_15329,N_15204);
nor U16369 (N_16369,N_15520,N_15228);
or U16370 (N_16370,N_15277,N_15461);
nand U16371 (N_16371,N_15431,N_15013);
xor U16372 (N_16372,N_15329,N_15582);
or U16373 (N_16373,N_15448,N_15221);
nand U16374 (N_16374,N_14644,N_15265);
nor U16375 (N_16375,N_15234,N_14783);
nor U16376 (N_16376,N_14576,N_14504);
nor U16377 (N_16377,N_15272,N_14722);
and U16378 (N_16378,N_15467,N_14528);
or U16379 (N_16379,N_15127,N_14738);
or U16380 (N_16380,N_14793,N_14912);
or U16381 (N_16381,N_14459,N_14728);
nand U16382 (N_16382,N_14825,N_15394);
xnor U16383 (N_16383,N_15534,N_15078);
nand U16384 (N_16384,N_15554,N_15302);
or U16385 (N_16385,N_15556,N_14543);
nand U16386 (N_16386,N_14552,N_14406);
and U16387 (N_16387,N_14815,N_14589);
or U16388 (N_16388,N_14991,N_15431);
and U16389 (N_16389,N_15395,N_14528);
xor U16390 (N_16390,N_14737,N_14856);
nand U16391 (N_16391,N_15450,N_14697);
or U16392 (N_16392,N_15500,N_15136);
nand U16393 (N_16393,N_15285,N_14637);
nor U16394 (N_16394,N_14896,N_14961);
nand U16395 (N_16395,N_15174,N_15320);
nor U16396 (N_16396,N_14447,N_15038);
or U16397 (N_16397,N_14635,N_14414);
nand U16398 (N_16398,N_15042,N_15082);
xnor U16399 (N_16399,N_14487,N_14556);
xor U16400 (N_16400,N_15156,N_14788);
xor U16401 (N_16401,N_14554,N_14582);
and U16402 (N_16402,N_15594,N_14580);
nand U16403 (N_16403,N_15328,N_14467);
or U16404 (N_16404,N_14639,N_15205);
nor U16405 (N_16405,N_15010,N_14573);
xnor U16406 (N_16406,N_14929,N_14519);
nand U16407 (N_16407,N_14484,N_15075);
nand U16408 (N_16408,N_15341,N_14833);
and U16409 (N_16409,N_15305,N_14571);
xnor U16410 (N_16410,N_15541,N_15117);
nand U16411 (N_16411,N_14984,N_15303);
xnor U16412 (N_16412,N_15502,N_14671);
xnor U16413 (N_16413,N_15036,N_15026);
nand U16414 (N_16414,N_15178,N_15279);
nor U16415 (N_16415,N_15194,N_15158);
nor U16416 (N_16416,N_15168,N_15400);
and U16417 (N_16417,N_15327,N_14581);
nor U16418 (N_16418,N_15408,N_15479);
nor U16419 (N_16419,N_15225,N_14644);
nor U16420 (N_16420,N_15559,N_15010);
and U16421 (N_16421,N_15120,N_14418);
or U16422 (N_16422,N_15067,N_14695);
xnor U16423 (N_16423,N_15495,N_14813);
and U16424 (N_16424,N_15113,N_14434);
xnor U16425 (N_16425,N_14856,N_14676);
or U16426 (N_16426,N_15001,N_15032);
xnor U16427 (N_16427,N_15447,N_15403);
nor U16428 (N_16428,N_14775,N_14914);
and U16429 (N_16429,N_15445,N_15013);
nor U16430 (N_16430,N_15369,N_14501);
nand U16431 (N_16431,N_15305,N_14504);
and U16432 (N_16432,N_15088,N_15397);
or U16433 (N_16433,N_14539,N_15281);
xnor U16434 (N_16434,N_14974,N_15228);
nor U16435 (N_16435,N_15575,N_14992);
nor U16436 (N_16436,N_15350,N_15471);
or U16437 (N_16437,N_15535,N_15241);
or U16438 (N_16438,N_15379,N_14432);
or U16439 (N_16439,N_15029,N_15174);
nor U16440 (N_16440,N_14995,N_14921);
nand U16441 (N_16441,N_14854,N_14911);
xor U16442 (N_16442,N_14687,N_14628);
and U16443 (N_16443,N_15057,N_15563);
nor U16444 (N_16444,N_14788,N_15247);
nand U16445 (N_16445,N_15329,N_15093);
nor U16446 (N_16446,N_15129,N_14815);
and U16447 (N_16447,N_14929,N_14799);
nor U16448 (N_16448,N_14417,N_15513);
nand U16449 (N_16449,N_14768,N_15062);
and U16450 (N_16450,N_15042,N_14634);
nand U16451 (N_16451,N_14479,N_15019);
and U16452 (N_16452,N_14633,N_14607);
xnor U16453 (N_16453,N_14474,N_15458);
nor U16454 (N_16454,N_15485,N_15197);
xnor U16455 (N_16455,N_15237,N_15398);
and U16456 (N_16456,N_14824,N_15118);
xor U16457 (N_16457,N_15168,N_14768);
nor U16458 (N_16458,N_14876,N_14550);
and U16459 (N_16459,N_15269,N_14685);
xor U16460 (N_16460,N_15212,N_14689);
nand U16461 (N_16461,N_15037,N_15325);
nand U16462 (N_16462,N_14662,N_14796);
and U16463 (N_16463,N_15579,N_15397);
xnor U16464 (N_16464,N_14520,N_14937);
xor U16465 (N_16465,N_14859,N_15109);
nand U16466 (N_16466,N_15419,N_14537);
nor U16467 (N_16467,N_15487,N_14795);
nor U16468 (N_16468,N_14642,N_15010);
and U16469 (N_16469,N_15348,N_14664);
and U16470 (N_16470,N_14548,N_14763);
nand U16471 (N_16471,N_15506,N_15259);
xnor U16472 (N_16472,N_15573,N_14536);
and U16473 (N_16473,N_15329,N_15044);
xor U16474 (N_16474,N_15442,N_14509);
nand U16475 (N_16475,N_14612,N_15135);
or U16476 (N_16476,N_14947,N_14885);
nor U16477 (N_16477,N_15547,N_15545);
nor U16478 (N_16478,N_14447,N_14566);
and U16479 (N_16479,N_15049,N_15422);
or U16480 (N_16480,N_15374,N_15150);
or U16481 (N_16481,N_14814,N_15431);
or U16482 (N_16482,N_15198,N_14975);
or U16483 (N_16483,N_14499,N_14487);
and U16484 (N_16484,N_14604,N_15009);
nand U16485 (N_16485,N_15279,N_15327);
nand U16486 (N_16486,N_15119,N_15161);
nand U16487 (N_16487,N_15348,N_14477);
and U16488 (N_16488,N_15180,N_15381);
nor U16489 (N_16489,N_14404,N_15341);
nor U16490 (N_16490,N_14598,N_15189);
xnor U16491 (N_16491,N_15546,N_15250);
xnor U16492 (N_16492,N_15455,N_14960);
xnor U16493 (N_16493,N_15470,N_14693);
and U16494 (N_16494,N_14949,N_15569);
nand U16495 (N_16495,N_15225,N_14771);
nor U16496 (N_16496,N_15539,N_14948);
xor U16497 (N_16497,N_15540,N_15221);
and U16498 (N_16498,N_14804,N_15197);
nor U16499 (N_16499,N_14831,N_14686);
and U16500 (N_16500,N_15196,N_14570);
and U16501 (N_16501,N_15450,N_14536);
and U16502 (N_16502,N_14581,N_14950);
and U16503 (N_16503,N_15486,N_14464);
xor U16504 (N_16504,N_15276,N_15335);
or U16505 (N_16505,N_14523,N_14935);
nor U16506 (N_16506,N_15039,N_14705);
xnor U16507 (N_16507,N_15337,N_15462);
nor U16508 (N_16508,N_14649,N_15295);
or U16509 (N_16509,N_14955,N_15538);
or U16510 (N_16510,N_15136,N_15211);
nand U16511 (N_16511,N_15431,N_14718);
or U16512 (N_16512,N_14614,N_15431);
nand U16513 (N_16513,N_15523,N_14506);
or U16514 (N_16514,N_15121,N_15508);
nand U16515 (N_16515,N_15041,N_15568);
and U16516 (N_16516,N_14879,N_15176);
and U16517 (N_16517,N_14474,N_14888);
and U16518 (N_16518,N_14768,N_14774);
nor U16519 (N_16519,N_15140,N_15157);
and U16520 (N_16520,N_14977,N_15210);
and U16521 (N_16521,N_14566,N_15002);
or U16522 (N_16522,N_14735,N_15117);
nor U16523 (N_16523,N_15473,N_15324);
and U16524 (N_16524,N_15356,N_15264);
nand U16525 (N_16525,N_15242,N_15353);
nand U16526 (N_16526,N_15103,N_14694);
nor U16527 (N_16527,N_15239,N_14477);
nand U16528 (N_16528,N_14970,N_15381);
nor U16529 (N_16529,N_14878,N_14815);
and U16530 (N_16530,N_14725,N_15333);
xnor U16531 (N_16531,N_15538,N_14644);
nor U16532 (N_16532,N_14850,N_15443);
or U16533 (N_16533,N_15165,N_15397);
xnor U16534 (N_16534,N_14971,N_14798);
nand U16535 (N_16535,N_15120,N_15019);
nand U16536 (N_16536,N_15054,N_14687);
and U16537 (N_16537,N_14686,N_15359);
nand U16538 (N_16538,N_15400,N_14420);
or U16539 (N_16539,N_14804,N_14482);
nor U16540 (N_16540,N_15127,N_15221);
nand U16541 (N_16541,N_15308,N_15551);
and U16542 (N_16542,N_15053,N_14978);
and U16543 (N_16543,N_15243,N_14926);
xor U16544 (N_16544,N_15572,N_15578);
nand U16545 (N_16545,N_14733,N_14462);
xor U16546 (N_16546,N_15006,N_14762);
nand U16547 (N_16547,N_14939,N_14612);
nand U16548 (N_16548,N_14496,N_15194);
nand U16549 (N_16549,N_15496,N_15110);
and U16550 (N_16550,N_14984,N_15469);
and U16551 (N_16551,N_15421,N_15541);
or U16552 (N_16552,N_14689,N_14535);
xnor U16553 (N_16553,N_14534,N_15473);
nor U16554 (N_16554,N_14835,N_15182);
nor U16555 (N_16555,N_15296,N_15207);
nor U16556 (N_16556,N_15283,N_14997);
xor U16557 (N_16557,N_14624,N_15290);
nor U16558 (N_16558,N_15403,N_15594);
nand U16559 (N_16559,N_15324,N_15219);
xnor U16560 (N_16560,N_14429,N_14486);
nand U16561 (N_16561,N_14582,N_15377);
nor U16562 (N_16562,N_15295,N_15003);
nand U16563 (N_16563,N_15242,N_15194);
nand U16564 (N_16564,N_15565,N_15545);
nand U16565 (N_16565,N_15077,N_14642);
xnor U16566 (N_16566,N_14491,N_14569);
xnor U16567 (N_16567,N_14567,N_14858);
or U16568 (N_16568,N_15187,N_14947);
nor U16569 (N_16569,N_14930,N_15376);
or U16570 (N_16570,N_14707,N_15258);
nor U16571 (N_16571,N_15148,N_14794);
or U16572 (N_16572,N_14859,N_14908);
nor U16573 (N_16573,N_14803,N_15470);
nor U16574 (N_16574,N_15526,N_15013);
nor U16575 (N_16575,N_14709,N_14518);
and U16576 (N_16576,N_15390,N_15450);
nor U16577 (N_16577,N_14495,N_14667);
xor U16578 (N_16578,N_15437,N_15179);
nor U16579 (N_16579,N_15595,N_15315);
nand U16580 (N_16580,N_14543,N_15080);
and U16581 (N_16581,N_15384,N_14834);
nand U16582 (N_16582,N_15529,N_14655);
xor U16583 (N_16583,N_15272,N_15072);
and U16584 (N_16584,N_14564,N_15214);
or U16585 (N_16585,N_15177,N_15508);
xnor U16586 (N_16586,N_14818,N_14602);
and U16587 (N_16587,N_14857,N_14970);
or U16588 (N_16588,N_15469,N_14684);
xnor U16589 (N_16589,N_14851,N_14423);
nand U16590 (N_16590,N_15110,N_15494);
xor U16591 (N_16591,N_15059,N_14839);
xnor U16592 (N_16592,N_15098,N_15391);
nor U16593 (N_16593,N_15536,N_15301);
nor U16594 (N_16594,N_14703,N_15181);
xor U16595 (N_16595,N_14649,N_14542);
or U16596 (N_16596,N_14644,N_15214);
and U16597 (N_16597,N_14603,N_14636);
xnor U16598 (N_16598,N_15424,N_15193);
nor U16599 (N_16599,N_15327,N_15309);
nand U16600 (N_16600,N_15220,N_14686);
or U16601 (N_16601,N_14883,N_15259);
nand U16602 (N_16602,N_15069,N_15404);
nor U16603 (N_16603,N_15419,N_15405);
or U16604 (N_16604,N_14892,N_14666);
xnor U16605 (N_16605,N_15269,N_15241);
nor U16606 (N_16606,N_15421,N_14497);
xnor U16607 (N_16607,N_15565,N_14933);
nor U16608 (N_16608,N_14821,N_15592);
and U16609 (N_16609,N_15457,N_14581);
nor U16610 (N_16610,N_15180,N_15116);
nor U16611 (N_16611,N_14471,N_15241);
and U16612 (N_16612,N_14962,N_14591);
nand U16613 (N_16613,N_14641,N_15512);
nand U16614 (N_16614,N_15128,N_15030);
or U16615 (N_16615,N_14832,N_15409);
nor U16616 (N_16616,N_15200,N_15181);
and U16617 (N_16617,N_14988,N_14843);
nor U16618 (N_16618,N_15323,N_15522);
or U16619 (N_16619,N_15219,N_14995);
xnor U16620 (N_16620,N_15084,N_15505);
nor U16621 (N_16621,N_14691,N_14462);
nand U16622 (N_16622,N_14899,N_14736);
nand U16623 (N_16623,N_14438,N_15166);
or U16624 (N_16624,N_14516,N_15532);
nand U16625 (N_16625,N_15137,N_15470);
nor U16626 (N_16626,N_14460,N_14949);
nand U16627 (N_16627,N_15229,N_14581);
nor U16628 (N_16628,N_15492,N_15476);
or U16629 (N_16629,N_14543,N_14511);
nand U16630 (N_16630,N_15076,N_14914);
nor U16631 (N_16631,N_14497,N_15477);
or U16632 (N_16632,N_15283,N_15189);
xor U16633 (N_16633,N_15237,N_14850);
or U16634 (N_16634,N_15120,N_14537);
nand U16635 (N_16635,N_14443,N_15158);
or U16636 (N_16636,N_14539,N_14565);
xnor U16637 (N_16637,N_15462,N_15229);
xor U16638 (N_16638,N_15444,N_15000);
and U16639 (N_16639,N_14491,N_15257);
nand U16640 (N_16640,N_14576,N_15144);
or U16641 (N_16641,N_14537,N_14442);
nand U16642 (N_16642,N_14518,N_15433);
nand U16643 (N_16643,N_15256,N_15518);
or U16644 (N_16644,N_14988,N_15449);
or U16645 (N_16645,N_15485,N_15388);
xor U16646 (N_16646,N_15152,N_15406);
nor U16647 (N_16647,N_15477,N_15494);
nor U16648 (N_16648,N_14716,N_14513);
or U16649 (N_16649,N_14479,N_15035);
and U16650 (N_16650,N_14839,N_15295);
nand U16651 (N_16651,N_14505,N_14948);
nor U16652 (N_16652,N_15552,N_15474);
nand U16653 (N_16653,N_15562,N_15404);
nand U16654 (N_16654,N_15203,N_14603);
or U16655 (N_16655,N_14976,N_14465);
xor U16656 (N_16656,N_15224,N_14660);
nor U16657 (N_16657,N_15242,N_15342);
xnor U16658 (N_16658,N_15455,N_15310);
and U16659 (N_16659,N_15202,N_14494);
and U16660 (N_16660,N_15209,N_15064);
nor U16661 (N_16661,N_15499,N_15598);
nand U16662 (N_16662,N_15257,N_15559);
nand U16663 (N_16663,N_14514,N_15406);
nand U16664 (N_16664,N_15519,N_15561);
or U16665 (N_16665,N_14776,N_15098);
and U16666 (N_16666,N_15539,N_15255);
xnor U16667 (N_16667,N_15037,N_15486);
nor U16668 (N_16668,N_14636,N_15208);
or U16669 (N_16669,N_15010,N_14675);
or U16670 (N_16670,N_15273,N_15258);
and U16671 (N_16671,N_15345,N_14567);
xnor U16672 (N_16672,N_14673,N_15393);
and U16673 (N_16673,N_15573,N_15243);
nand U16674 (N_16674,N_14930,N_14419);
nand U16675 (N_16675,N_15507,N_15505);
xor U16676 (N_16676,N_15448,N_14647);
nor U16677 (N_16677,N_14533,N_15116);
nor U16678 (N_16678,N_14787,N_14989);
and U16679 (N_16679,N_14701,N_14697);
nor U16680 (N_16680,N_15534,N_14455);
nor U16681 (N_16681,N_14649,N_14788);
or U16682 (N_16682,N_15263,N_14833);
nand U16683 (N_16683,N_15570,N_14957);
xor U16684 (N_16684,N_15489,N_14456);
nand U16685 (N_16685,N_15351,N_14567);
nand U16686 (N_16686,N_14534,N_14552);
or U16687 (N_16687,N_15024,N_15384);
xor U16688 (N_16688,N_15489,N_15261);
xnor U16689 (N_16689,N_15330,N_14411);
xor U16690 (N_16690,N_15451,N_14525);
xnor U16691 (N_16691,N_14534,N_14603);
and U16692 (N_16692,N_14780,N_15436);
and U16693 (N_16693,N_14838,N_14535);
and U16694 (N_16694,N_14692,N_15404);
or U16695 (N_16695,N_15330,N_14614);
xnor U16696 (N_16696,N_15180,N_15427);
or U16697 (N_16697,N_14862,N_14699);
and U16698 (N_16698,N_15315,N_14672);
or U16699 (N_16699,N_15530,N_14852);
nor U16700 (N_16700,N_15233,N_15439);
and U16701 (N_16701,N_15268,N_14886);
and U16702 (N_16702,N_14722,N_14509);
xor U16703 (N_16703,N_14566,N_14948);
nor U16704 (N_16704,N_15536,N_14639);
or U16705 (N_16705,N_14861,N_14890);
or U16706 (N_16706,N_14832,N_14551);
nand U16707 (N_16707,N_14651,N_14954);
nor U16708 (N_16708,N_14659,N_15265);
and U16709 (N_16709,N_14601,N_14791);
xor U16710 (N_16710,N_14752,N_15396);
xor U16711 (N_16711,N_14427,N_14726);
nand U16712 (N_16712,N_15512,N_15058);
or U16713 (N_16713,N_15122,N_15011);
or U16714 (N_16714,N_15265,N_14581);
and U16715 (N_16715,N_14685,N_15362);
nand U16716 (N_16716,N_15464,N_14522);
and U16717 (N_16717,N_15431,N_15219);
or U16718 (N_16718,N_15322,N_14546);
nand U16719 (N_16719,N_15514,N_14724);
and U16720 (N_16720,N_15227,N_14715);
and U16721 (N_16721,N_14569,N_14689);
nor U16722 (N_16722,N_15008,N_14659);
and U16723 (N_16723,N_14434,N_14704);
and U16724 (N_16724,N_14925,N_14989);
nand U16725 (N_16725,N_14804,N_14594);
nand U16726 (N_16726,N_15556,N_15263);
nand U16727 (N_16727,N_14625,N_14897);
nand U16728 (N_16728,N_15286,N_14682);
nand U16729 (N_16729,N_14647,N_15489);
or U16730 (N_16730,N_15131,N_14549);
or U16731 (N_16731,N_15536,N_14459);
and U16732 (N_16732,N_15590,N_14528);
and U16733 (N_16733,N_15450,N_14588);
and U16734 (N_16734,N_14711,N_14637);
or U16735 (N_16735,N_14724,N_14433);
or U16736 (N_16736,N_15466,N_15170);
xor U16737 (N_16737,N_14711,N_14659);
or U16738 (N_16738,N_15525,N_15101);
and U16739 (N_16739,N_14453,N_14528);
and U16740 (N_16740,N_14870,N_15550);
or U16741 (N_16741,N_14776,N_14642);
nand U16742 (N_16742,N_14578,N_15207);
xor U16743 (N_16743,N_15504,N_15544);
nand U16744 (N_16744,N_15537,N_15568);
and U16745 (N_16745,N_14970,N_15425);
or U16746 (N_16746,N_15239,N_15096);
or U16747 (N_16747,N_15105,N_14927);
nor U16748 (N_16748,N_14803,N_14907);
and U16749 (N_16749,N_14865,N_15372);
or U16750 (N_16750,N_15532,N_14527);
nor U16751 (N_16751,N_15111,N_15203);
or U16752 (N_16752,N_14862,N_15074);
xor U16753 (N_16753,N_15557,N_14822);
and U16754 (N_16754,N_14673,N_15095);
nand U16755 (N_16755,N_15305,N_14869);
or U16756 (N_16756,N_14461,N_15463);
nor U16757 (N_16757,N_14430,N_14484);
or U16758 (N_16758,N_15203,N_14649);
nand U16759 (N_16759,N_14747,N_15368);
nand U16760 (N_16760,N_14522,N_14622);
nor U16761 (N_16761,N_14468,N_14506);
or U16762 (N_16762,N_14519,N_14569);
nand U16763 (N_16763,N_14491,N_14909);
or U16764 (N_16764,N_15574,N_15255);
xnor U16765 (N_16765,N_14882,N_15411);
xor U16766 (N_16766,N_15248,N_15491);
xor U16767 (N_16767,N_14915,N_14579);
xor U16768 (N_16768,N_14790,N_14915);
or U16769 (N_16769,N_14956,N_15518);
and U16770 (N_16770,N_14566,N_14997);
and U16771 (N_16771,N_15171,N_15310);
nand U16772 (N_16772,N_15001,N_14584);
and U16773 (N_16773,N_15131,N_15243);
nand U16774 (N_16774,N_15380,N_14632);
xnor U16775 (N_16775,N_14619,N_14812);
nand U16776 (N_16776,N_15497,N_15026);
nand U16777 (N_16777,N_14960,N_14712);
or U16778 (N_16778,N_15027,N_14885);
or U16779 (N_16779,N_15242,N_15201);
and U16780 (N_16780,N_14577,N_15247);
or U16781 (N_16781,N_14692,N_15295);
and U16782 (N_16782,N_15166,N_14461);
xor U16783 (N_16783,N_15085,N_15494);
xnor U16784 (N_16784,N_14731,N_15466);
nand U16785 (N_16785,N_15275,N_15051);
or U16786 (N_16786,N_15519,N_15469);
nand U16787 (N_16787,N_14735,N_14612);
nor U16788 (N_16788,N_15187,N_14936);
and U16789 (N_16789,N_14413,N_15573);
or U16790 (N_16790,N_14447,N_14455);
xor U16791 (N_16791,N_14702,N_15293);
xnor U16792 (N_16792,N_14650,N_14994);
or U16793 (N_16793,N_15423,N_15550);
nand U16794 (N_16794,N_14515,N_15463);
nor U16795 (N_16795,N_15201,N_14657);
and U16796 (N_16796,N_14491,N_15412);
xor U16797 (N_16797,N_14592,N_14790);
nor U16798 (N_16798,N_15489,N_15530);
or U16799 (N_16799,N_14445,N_15201);
and U16800 (N_16800,N_15792,N_16741);
and U16801 (N_16801,N_16241,N_15973);
nor U16802 (N_16802,N_16256,N_16073);
and U16803 (N_16803,N_15931,N_16394);
and U16804 (N_16804,N_16680,N_16711);
and U16805 (N_16805,N_16062,N_16556);
nand U16806 (N_16806,N_16548,N_16716);
and U16807 (N_16807,N_15847,N_15905);
and U16808 (N_16808,N_16725,N_15799);
and U16809 (N_16809,N_16583,N_16077);
xor U16810 (N_16810,N_15972,N_16646);
nand U16811 (N_16811,N_16166,N_16459);
and U16812 (N_16812,N_16371,N_15889);
and U16813 (N_16813,N_16032,N_15734);
nand U16814 (N_16814,N_16316,N_16214);
xnor U16815 (N_16815,N_15895,N_15774);
nor U16816 (N_16816,N_16497,N_15967);
xor U16817 (N_16817,N_15713,N_16204);
nand U16818 (N_16818,N_16427,N_16696);
nor U16819 (N_16819,N_16217,N_16253);
or U16820 (N_16820,N_16639,N_16345);
nand U16821 (N_16821,N_15773,N_15764);
and U16822 (N_16822,N_16428,N_15939);
and U16823 (N_16823,N_15633,N_16463);
nor U16824 (N_16824,N_16335,N_15703);
xor U16825 (N_16825,N_15708,N_16719);
xnor U16826 (N_16826,N_15927,N_16582);
and U16827 (N_16827,N_16642,N_16495);
or U16828 (N_16828,N_16012,N_16617);
and U16829 (N_16829,N_15894,N_16657);
nor U16830 (N_16830,N_16175,N_16420);
and U16831 (N_16831,N_15750,N_15740);
nor U16832 (N_16832,N_15920,N_15828);
nand U16833 (N_16833,N_16740,N_16407);
or U16834 (N_16834,N_16515,N_15963);
nand U16835 (N_16835,N_16588,N_15798);
xor U16836 (N_16836,N_16191,N_16036);
xor U16837 (N_16837,N_16195,N_16436);
nand U16838 (N_16838,N_15641,N_16013);
and U16839 (N_16839,N_16550,N_15690);
xor U16840 (N_16840,N_16792,N_16322);
or U16841 (N_16841,N_15675,N_16708);
xnor U16842 (N_16842,N_16659,N_15659);
nor U16843 (N_16843,N_16772,N_16343);
or U16844 (N_16844,N_16167,N_15677);
nand U16845 (N_16845,N_15639,N_16360);
nor U16846 (N_16846,N_16555,N_16328);
nor U16847 (N_16847,N_16462,N_15819);
nand U16848 (N_16848,N_16076,N_16765);
xnor U16849 (N_16849,N_15715,N_16121);
nor U16850 (N_16850,N_15691,N_15787);
xnor U16851 (N_16851,N_16728,N_16212);
and U16852 (N_16852,N_16361,N_16211);
xnor U16853 (N_16853,N_15755,N_16612);
xor U16854 (N_16854,N_15689,N_16049);
and U16855 (N_16855,N_16457,N_15692);
nand U16856 (N_16856,N_15849,N_16567);
or U16857 (N_16857,N_16501,N_15609);
and U16858 (N_16858,N_16664,N_16291);
xor U16859 (N_16859,N_16504,N_16480);
nand U16860 (N_16860,N_15606,N_16187);
xor U16861 (N_16861,N_16178,N_16730);
nor U16862 (N_16862,N_16472,N_16652);
and U16863 (N_16863,N_16488,N_16275);
nor U16864 (N_16864,N_16602,N_16786);
nor U16865 (N_16865,N_16162,N_16438);
or U16866 (N_16866,N_16110,N_15942);
or U16867 (N_16867,N_16372,N_16458);
and U16868 (N_16868,N_15970,N_16237);
xor U16869 (N_16869,N_16601,N_16282);
or U16870 (N_16870,N_16311,N_16240);
nor U16871 (N_16871,N_16344,N_16577);
nor U16872 (N_16872,N_16055,N_16337);
or U16873 (N_16873,N_16125,N_15861);
nor U16874 (N_16874,N_15762,N_16009);
xnor U16875 (N_16875,N_15800,N_16593);
nand U16876 (N_16876,N_16114,N_16748);
xnor U16877 (N_16877,N_15845,N_16494);
or U16878 (N_16878,N_15682,N_16339);
nand U16879 (N_16879,N_16757,N_15673);
xnor U16880 (N_16880,N_15701,N_16419);
and U16881 (N_16881,N_16262,N_16367);
nand U16882 (N_16882,N_15637,N_16284);
and U16883 (N_16883,N_16305,N_16723);
and U16884 (N_16884,N_15936,N_16425);
or U16885 (N_16885,N_16393,N_16053);
nand U16886 (N_16886,N_16455,N_15718);
nor U16887 (N_16887,N_16151,N_16700);
or U16888 (N_16888,N_15749,N_16201);
or U16889 (N_16889,N_16105,N_16699);
nand U16890 (N_16890,N_16243,N_16205);
xor U16891 (N_16891,N_16521,N_16742);
and U16892 (N_16892,N_15918,N_16492);
and U16893 (N_16893,N_15891,N_15932);
nor U16894 (N_16894,N_16308,N_15900);
nor U16895 (N_16895,N_15661,N_16138);
xor U16896 (N_16896,N_15765,N_16570);
or U16897 (N_16897,N_15980,N_16043);
xnor U16898 (N_16898,N_16010,N_16259);
and U16899 (N_16899,N_16014,N_15934);
nand U16900 (N_16900,N_16537,N_16683);
xnor U16901 (N_16901,N_16440,N_15699);
xnor U16902 (N_16902,N_16724,N_15611);
and U16903 (N_16903,N_15922,N_15618);
nand U16904 (N_16904,N_16535,N_16510);
nor U16905 (N_16905,N_16784,N_15992);
xnor U16906 (N_16906,N_16695,N_15822);
nor U16907 (N_16907,N_16296,N_16611);
nor U16908 (N_16908,N_16314,N_16518);
and U16909 (N_16909,N_15753,N_15614);
nand U16910 (N_16910,N_16264,N_16600);
nor U16911 (N_16911,N_16271,N_16397);
or U16912 (N_16912,N_16368,N_16775);
xnor U16913 (N_16913,N_15712,N_16605);
and U16914 (N_16914,N_16244,N_16760);
or U16915 (N_16915,N_15671,N_16727);
or U16916 (N_16916,N_16127,N_16050);
and U16917 (N_16917,N_15707,N_16587);
and U16918 (N_16918,N_16456,N_16622);
or U16919 (N_16919,N_16126,N_16489);
xnor U16920 (N_16920,N_16059,N_16513);
xnor U16921 (N_16921,N_16464,N_15770);
nand U16922 (N_16922,N_16029,N_16758);
xnor U16923 (N_16923,N_15772,N_16446);
xor U16924 (N_16924,N_15870,N_15860);
nor U16925 (N_16925,N_16392,N_16242);
or U16926 (N_16926,N_16576,N_15930);
and U16927 (N_16927,N_16762,N_16453);
or U16928 (N_16928,N_16402,N_15721);
nor U16929 (N_16929,N_16528,N_16389);
xnor U16930 (N_16930,N_16219,N_15783);
nand U16931 (N_16931,N_16635,N_16767);
nand U16932 (N_16932,N_15743,N_15610);
nor U16933 (N_16933,N_16268,N_15741);
xnor U16934 (N_16934,N_15790,N_16325);
and U16935 (N_16935,N_16682,N_15812);
and U16936 (N_16936,N_15758,N_16194);
xor U16937 (N_16937,N_15959,N_16406);
nor U16938 (N_16938,N_16418,N_16273);
or U16939 (N_16939,N_15766,N_15984);
nor U16940 (N_16940,N_16746,N_16040);
xor U16941 (N_16941,N_15802,N_16750);
and U16942 (N_16942,N_15638,N_16159);
nand U16943 (N_16943,N_16156,N_16118);
xnor U16944 (N_16944,N_16293,N_16207);
or U16945 (N_16945,N_15886,N_15841);
or U16946 (N_16946,N_16661,N_15901);
nand U16947 (N_16947,N_16452,N_16147);
nor U16948 (N_16948,N_15817,N_16355);
nand U16949 (N_16949,N_16479,N_15823);
xor U16950 (N_16950,N_16058,N_16737);
or U16951 (N_16951,N_16434,N_15838);
or U16952 (N_16952,N_16670,N_15757);
or U16953 (N_16953,N_15612,N_16552);
and U16954 (N_16954,N_16396,N_16713);
and U16955 (N_16955,N_16752,N_16060);
nor U16956 (N_16956,N_16277,N_16512);
or U16957 (N_16957,N_16477,N_16668);
nor U16958 (N_16958,N_16304,N_16093);
nor U16959 (N_16959,N_16132,N_15852);
or U16960 (N_16960,N_16496,N_16421);
and U16961 (N_16961,N_16616,N_15917);
xnor U16962 (N_16962,N_15977,N_16177);
nor U16963 (N_16963,N_16729,N_15957);
and U16964 (N_16964,N_15872,N_16743);
or U16965 (N_16965,N_16306,N_16689);
xor U16966 (N_16966,N_16329,N_16761);
or U16967 (N_16967,N_16584,N_15884);
nand U16968 (N_16968,N_15668,N_15897);
or U16969 (N_16969,N_15751,N_15719);
nand U16970 (N_16970,N_15794,N_16566);
xnor U16971 (N_16971,N_16365,N_16416);
nand U16972 (N_16972,N_16065,N_16313);
and U16973 (N_16973,N_16033,N_16019);
nand U16974 (N_16974,N_16056,N_16377);
xnor U16975 (N_16975,N_15694,N_16395);
nand U16976 (N_16976,N_16095,N_16349);
nand U16977 (N_16977,N_16011,N_16503);
xnor U16978 (N_16978,N_16063,N_15769);
and U16979 (N_16979,N_16348,N_16660);
nand U16980 (N_16980,N_15864,N_16034);
or U16981 (N_16981,N_15634,N_16112);
nor U16982 (N_16982,N_16514,N_16644);
xor U16983 (N_16983,N_16254,N_16720);
nand U16984 (N_16984,N_16651,N_16274);
xnor U16985 (N_16985,N_16190,N_16285);
nor U16986 (N_16986,N_15815,N_15960);
nor U16987 (N_16987,N_16656,N_16119);
xor U16988 (N_16988,N_16776,N_16078);
nor U16989 (N_16989,N_16783,N_16523);
or U16990 (N_16990,N_15966,N_16409);
nor U16991 (N_16991,N_16563,N_16744);
or U16992 (N_16992,N_16002,N_15684);
nor U16993 (N_16993,N_16267,N_16069);
xnor U16994 (N_16994,N_16183,N_16405);
and U16995 (N_16995,N_16039,N_15605);
xor U16996 (N_16996,N_16297,N_16082);
nand U16997 (N_16997,N_16735,N_16520);
and U16998 (N_16998,N_16384,N_16326);
or U16999 (N_16999,N_16613,N_16486);
xnor U17000 (N_17000,N_15602,N_16290);
nand U17001 (N_17001,N_15655,N_16410);
nand U17002 (N_17002,N_16522,N_16667);
xnor U17003 (N_17003,N_16142,N_16097);
nand U17004 (N_17004,N_16353,N_15991);
or U17005 (N_17005,N_16079,N_15746);
nor U17006 (N_17006,N_15874,N_16272);
nor U17007 (N_17007,N_15848,N_15625);
xor U17008 (N_17008,N_16454,N_16359);
xor U17009 (N_17009,N_16255,N_16764);
nor U17010 (N_17010,N_16221,N_16694);
nor U17011 (N_17011,N_15859,N_15667);
or U17012 (N_17012,N_16592,N_16681);
nor U17013 (N_17013,N_16197,N_16035);
and U17014 (N_17014,N_15644,N_16712);
xnor U17015 (N_17015,N_15883,N_15627);
nor U17016 (N_17016,N_16442,N_16531);
nor U17017 (N_17017,N_16176,N_16422);
or U17018 (N_17018,N_15670,N_16228);
and U17019 (N_17019,N_15801,N_16474);
xnor U17020 (N_17020,N_15925,N_16084);
and U17021 (N_17021,N_16623,N_16071);
or U17022 (N_17022,N_16491,N_16412);
or U17023 (N_17023,N_15808,N_15958);
xor U17024 (N_17024,N_16334,N_16092);
or U17025 (N_17025,N_16785,N_16157);
and U17026 (N_17026,N_16122,N_16266);
xor U17027 (N_17027,N_16301,N_16350);
nand U17028 (N_17028,N_15723,N_16146);
nor U17029 (N_17029,N_16323,N_15730);
nand U17030 (N_17030,N_16778,N_16276);
or U17031 (N_17031,N_16202,N_16370);
nor U17032 (N_17032,N_16170,N_15896);
nand U17033 (N_17033,N_16770,N_16490);
xnor U17034 (N_17034,N_15865,N_16100);
or U17035 (N_17035,N_16249,N_15748);
and U17036 (N_17036,N_16717,N_16051);
or U17037 (N_17037,N_16286,N_16527);
nor U17038 (N_17038,N_16650,N_16378);
or U17039 (N_17039,N_16229,N_16089);
nor U17040 (N_17040,N_16572,N_16192);
and U17041 (N_17041,N_15990,N_15926);
xor U17042 (N_17042,N_16684,N_16731);
and U17043 (N_17043,N_15988,N_16715);
and U17044 (N_17044,N_16478,N_16469);
nand U17045 (N_17045,N_15676,N_16774);
nor U17046 (N_17046,N_15853,N_16709);
nand U17047 (N_17047,N_16099,N_16338);
xnor U17048 (N_17048,N_16231,N_16686);
and U17049 (N_17049,N_15956,N_15752);
nor U17050 (N_17050,N_16104,N_15747);
nor U17051 (N_17051,N_16626,N_16358);
and U17052 (N_17052,N_15771,N_16096);
nor U17053 (N_17053,N_16248,N_15854);
and U17054 (N_17054,N_16634,N_16632);
xnor U17055 (N_17055,N_16075,N_15731);
or U17056 (N_17056,N_16590,N_16468);
xor U17057 (N_17057,N_16585,N_16356);
or U17058 (N_17058,N_16484,N_16714);
xnor U17059 (N_17059,N_15726,N_15754);
nand U17060 (N_17060,N_16481,N_16706);
xor U17061 (N_17061,N_15805,N_15919);
nand U17062 (N_17062,N_16648,N_16074);
or U17063 (N_17063,N_16134,N_15867);
and U17064 (N_17064,N_16354,N_15706);
and U17065 (N_17065,N_16210,N_16173);
and U17066 (N_17066,N_16400,N_15873);
nand U17067 (N_17067,N_16150,N_16287);
and U17068 (N_17068,N_16791,N_15698);
and U17069 (N_17069,N_15724,N_16120);
xnor U17070 (N_17070,N_15680,N_15658);
or U17071 (N_17071,N_16128,N_16441);
and U17072 (N_17072,N_15825,N_16558);
nand U17073 (N_17073,N_15842,N_16280);
xor U17074 (N_17074,N_15732,N_15810);
and U17075 (N_17075,N_16318,N_15603);
nor U17076 (N_17076,N_16732,N_16645);
nand U17077 (N_17077,N_16546,N_15780);
nand U17078 (N_17078,N_16139,N_15647);
and U17079 (N_17079,N_15814,N_15964);
xnor U17080 (N_17080,N_16090,N_16519);
xor U17081 (N_17081,N_15782,N_16363);
nor U17082 (N_17082,N_16466,N_16580);
nand U17083 (N_17083,N_16790,N_15785);
nand U17084 (N_17084,N_16754,N_16663);
and U17085 (N_17085,N_16545,N_15735);
nand U17086 (N_17086,N_15950,N_15649);
nand U17087 (N_17087,N_16245,N_15786);
xnor U17088 (N_17088,N_16766,N_15678);
or U17089 (N_17089,N_15803,N_16470);
and U17090 (N_17090,N_16148,N_15687);
or U17091 (N_17091,N_16020,N_15613);
xnor U17092 (N_17092,N_16589,N_15722);
xnor U17093 (N_17093,N_16598,N_16007);
or U17094 (N_17094,N_16530,N_16027);
and U17095 (N_17095,N_16072,N_16431);
nor U17096 (N_17096,N_16199,N_16144);
nand U17097 (N_17097,N_16437,N_15816);
and U17098 (N_17098,N_16391,N_15804);
or U17099 (N_17099,N_16006,N_16030);
xnor U17100 (N_17100,N_15954,N_15928);
xnor U17101 (N_17101,N_16718,N_15700);
and U17102 (N_17102,N_16174,N_15788);
and U17103 (N_17103,N_16113,N_16630);
nor U17104 (N_17104,N_15789,N_16230);
nor U17105 (N_17105,N_16543,N_16239);
nand U17106 (N_17106,N_16057,N_16315);
nand U17107 (N_17107,N_16123,N_15656);
and U17108 (N_17108,N_16773,N_16251);
nor U17109 (N_17109,N_16184,N_15727);
nor U17110 (N_17110,N_16739,N_15821);
nand U17111 (N_17111,N_16444,N_15696);
nand U17112 (N_17112,N_16594,N_15946);
or U17113 (N_17113,N_15768,N_16685);
and U17114 (N_17114,N_15836,N_15796);
nand U17115 (N_17115,N_16795,N_16172);
nand U17116 (N_17116,N_15940,N_15813);
nand U17117 (N_17117,N_15921,N_16140);
and U17118 (N_17118,N_15733,N_16091);
nor U17119 (N_17119,N_16238,N_15906);
and U17120 (N_17120,N_15915,N_16398);
nor U17121 (N_17121,N_16485,N_16379);
xnor U17122 (N_17122,N_16381,N_16621);
nor U17123 (N_17123,N_16722,N_15978);
xor U17124 (N_17124,N_16688,N_16232);
xnor U17125 (N_17125,N_15650,N_16534);
and U17126 (N_17126,N_16129,N_16669);
or U17127 (N_17127,N_16373,N_15855);
nand U17128 (N_17128,N_15937,N_16575);
xor U17129 (N_17129,N_16070,N_16705);
xor U17130 (N_17130,N_16294,N_16269);
nand U17131 (N_17131,N_16016,N_15778);
and U17132 (N_17132,N_16516,N_16213);
nand U17133 (N_17133,N_15826,N_16141);
or U17134 (N_17134,N_16300,N_16022);
nand U17135 (N_17135,N_15648,N_16675);
nand U17136 (N_17136,N_16330,N_15736);
and U17137 (N_17137,N_16573,N_16265);
nand U17138 (N_17138,N_16111,N_16362);
nor U17139 (N_17139,N_16557,N_16781);
or U17140 (N_17140,N_15832,N_15965);
nor U17141 (N_17141,N_16149,N_16625);
nand U17142 (N_17142,N_16799,N_16386);
xnor U17143 (N_17143,N_16532,N_15857);
nand U17144 (N_17144,N_15929,N_15902);
nor U17145 (N_17145,N_16018,N_16413);
or U17146 (N_17146,N_16155,N_15616);
or U17147 (N_17147,N_16061,N_16346);
or U17148 (N_17148,N_16653,N_16046);
nor U17149 (N_17149,N_15737,N_15617);
nand U17150 (N_17150,N_15947,N_16672);
or U17151 (N_17151,N_15811,N_16517);
nor U17152 (N_17152,N_16771,N_15890);
or U17153 (N_17153,N_15974,N_15898);
and U17154 (N_17154,N_15907,N_15744);
nor U17155 (N_17155,N_16603,N_16364);
or U17156 (N_17156,N_16483,N_16751);
nor U17157 (N_17157,N_16562,N_16636);
or U17158 (N_17158,N_16226,N_16340);
nor U17159 (N_17159,N_16042,N_16375);
or U17160 (N_17160,N_15716,N_15624);
nand U17161 (N_17161,N_16498,N_16662);
and U17162 (N_17162,N_16618,N_16533);
xor U17163 (N_17163,N_16666,N_16257);
or U17164 (N_17164,N_16606,N_15830);
or U17165 (N_17165,N_15843,N_16258);
xnor U17166 (N_17166,N_16182,N_16703);
or U17167 (N_17167,N_15968,N_15738);
and U17168 (N_17168,N_15621,N_16263);
and U17169 (N_17169,N_16180,N_16687);
nor U17170 (N_17170,N_15685,N_16756);
and U17171 (N_17171,N_16031,N_16541);
and U17172 (N_17172,N_16445,N_15835);
or U17173 (N_17173,N_16143,N_16628);
nor U17174 (N_17174,N_15831,N_16136);
nand U17175 (N_17175,N_15871,N_16317);
nand U17176 (N_17176,N_16502,N_15756);
nor U17177 (N_17177,N_15953,N_16278);
nand U17178 (N_17178,N_16094,N_15885);
and U17179 (N_17179,N_16461,N_15941);
nor U17180 (N_17180,N_15989,N_16004);
xor U17181 (N_17181,N_15600,N_15664);
or U17182 (N_17182,N_15704,N_16450);
xor U17183 (N_17183,N_15666,N_16782);
nor U17184 (N_17184,N_15739,N_16508);
nor U17185 (N_17185,N_16408,N_16295);
and U17186 (N_17186,N_15879,N_16676);
nand U17187 (N_17187,N_16203,N_16261);
xnor U17188 (N_17188,N_16574,N_16279);
and U17189 (N_17189,N_15662,N_16564);
nand U17190 (N_17190,N_16702,N_15681);
nand U17191 (N_17191,N_16052,N_16789);
nand U17192 (N_17192,N_15729,N_15914);
xnor U17193 (N_17193,N_16005,N_16482);
or U17194 (N_17194,N_16430,N_16038);
xnor U17195 (N_17195,N_16116,N_16677);
nand U17196 (N_17196,N_15912,N_16475);
and U17197 (N_17197,N_15961,N_15640);
nand U17198 (N_17198,N_15986,N_16447);
nand U17199 (N_17199,N_16347,N_16250);
nor U17200 (N_17200,N_16044,N_15702);
xnor U17201 (N_17201,N_16499,N_16235);
nand U17202 (N_17202,N_16223,N_16793);
or U17203 (N_17203,N_16327,N_16607);
xnor U17204 (N_17204,N_15952,N_16568);
xnor U17205 (N_17205,N_16423,N_15809);
or U17206 (N_17206,N_16559,N_16544);
nor U17207 (N_17207,N_15630,N_16164);
xor U17208 (N_17208,N_15777,N_16200);
nor U17209 (N_17209,N_16135,N_15863);
nor U17210 (N_17210,N_16745,N_15651);
nand U17211 (N_17211,N_16342,N_16161);
nand U17212 (N_17212,N_16595,N_16388);
or U17213 (N_17213,N_15846,N_15615);
or U17214 (N_17214,N_16218,N_16401);
or U17215 (N_17215,N_15623,N_16753);
nand U17216 (N_17216,N_16193,N_16047);
and U17217 (N_17217,N_16234,N_15892);
nor U17218 (N_17218,N_16749,N_15910);
nor U17219 (N_17219,N_16168,N_15820);
or U17220 (N_17220,N_16467,N_16565);
or U17221 (N_17221,N_15626,N_15607);
nor U17222 (N_17222,N_16578,N_15629);
or U17223 (N_17223,N_16707,N_15784);
or U17224 (N_17224,N_16198,N_16387);
or U17225 (N_17225,N_16115,N_16015);
nor U17226 (N_17226,N_16797,N_16404);
nand U17227 (N_17227,N_16500,N_15653);
nor U17228 (N_17228,N_16614,N_16341);
nor U17229 (N_17229,N_15709,N_16698);
and U17230 (N_17230,N_16619,N_16476);
or U17231 (N_17231,N_15742,N_15829);
or U17232 (N_17232,N_15909,N_16179);
or U17233 (N_17233,N_15717,N_16299);
xnor U17234 (N_17234,N_15679,N_16154);
nand U17235 (N_17235,N_16374,N_15652);
xor U17236 (N_17236,N_16003,N_16638);
xor U17237 (N_17237,N_16041,N_16553);
nand U17238 (N_17238,N_16448,N_16206);
and U17239 (N_17239,N_15714,N_15996);
xnor U17240 (N_17240,N_16734,N_15979);
nand U17241 (N_17241,N_16390,N_16509);
xnor U17242 (N_17242,N_15948,N_16270);
xnor U17243 (N_17243,N_16560,N_15725);
xor U17244 (N_17244,N_15995,N_16281);
xnor U17245 (N_17245,N_16465,N_15697);
or U17246 (N_17246,N_15985,N_16721);
nand U17247 (N_17247,N_15993,N_16678);
or U17248 (N_17248,N_16321,N_16163);
nor U17249 (N_17249,N_16380,N_16227);
nand U17250 (N_17250,N_15844,N_16539);
and U17251 (N_17251,N_16586,N_16627);
or U17252 (N_17252,N_16117,N_15881);
or U17253 (N_17253,N_16169,N_16424);
nor U17254 (N_17254,N_16647,N_16252);
nand U17255 (N_17255,N_16629,N_16021);
xnor U17256 (N_17256,N_15660,N_15645);
nor U17257 (N_17257,N_16153,N_15944);
xnor U17258 (N_17258,N_16103,N_16704);
and U17259 (N_17259,N_16086,N_16763);
or U17260 (N_17260,N_16088,N_15999);
nand U17261 (N_17261,N_16188,N_16726);
nor U17262 (N_17262,N_15663,N_15969);
and U17263 (N_17263,N_15866,N_16411);
nand U17264 (N_17264,N_16109,N_15631);
and U17265 (N_17265,N_15665,N_16087);
and U17266 (N_17266,N_15851,N_16649);
nor U17267 (N_17267,N_16507,N_16637);
nand U17268 (N_17268,N_16222,N_16597);
xnor U17269 (N_17269,N_16697,N_16124);
or U17270 (N_17270,N_16383,N_16787);
xnor U17271 (N_17271,N_16549,N_16025);
and U17272 (N_17272,N_15779,N_16604);
xor U17273 (N_17273,N_16524,N_15837);
or U17274 (N_17274,N_16596,N_15862);
or U17275 (N_17275,N_16288,N_16561);
nor U17276 (N_17276,N_15833,N_16665);
or U17277 (N_17277,N_15899,N_16493);
nor U17278 (N_17278,N_16693,N_16691);
or U17279 (N_17279,N_16196,N_15806);
nor U17280 (N_17280,N_15850,N_16145);
and U17281 (N_17281,N_15827,N_16024);
xor U17282 (N_17282,N_16152,N_16220);
and U17283 (N_17283,N_15840,N_15643);
or U17284 (N_17284,N_16292,N_16026);
nand U17285 (N_17285,N_16298,N_15818);
nand U17286 (N_17286,N_15728,N_16654);
nor U17287 (N_17287,N_16054,N_15781);
xor U17288 (N_17288,N_16671,N_16303);
nand U17289 (N_17289,N_15935,N_16439);
nor U17290 (N_17290,N_15646,N_15880);
and U17291 (N_17291,N_15683,N_16609);
xor U17292 (N_17292,N_16529,N_16777);
or U17293 (N_17293,N_15998,N_16417);
and U17294 (N_17294,N_16131,N_15877);
or U17295 (N_17295,N_15976,N_15908);
nand U17296 (N_17296,N_16160,N_15686);
and U17297 (N_17297,N_16023,N_16643);
nor U17298 (N_17298,N_16000,N_16165);
nand U17299 (N_17299,N_16747,N_15949);
or U17300 (N_17300,N_15858,N_16351);
xor U17301 (N_17301,N_16620,N_16215);
xnor U17302 (N_17302,N_15695,N_16449);
or U17303 (N_17303,N_16526,N_16569);
nor U17304 (N_17304,N_15893,N_15654);
and U17305 (N_17305,N_16171,N_16008);
and U17306 (N_17306,N_15951,N_16547);
xor U17307 (N_17307,N_16208,N_15943);
nor U17308 (N_17308,N_16506,N_15760);
xnor U17309 (N_17309,N_16357,N_16336);
or U17310 (N_17310,N_16064,N_16352);
nor U17311 (N_17311,N_15657,N_15913);
and U17312 (N_17312,N_15776,N_16460);
nand U17313 (N_17313,N_16525,N_16102);
or U17314 (N_17314,N_16571,N_16692);
xnor U17315 (N_17315,N_16068,N_16673);
and U17316 (N_17316,N_16107,N_16302);
nor U17317 (N_17317,N_16615,N_16435);
or U17318 (N_17318,N_15795,N_15962);
or U17319 (N_17319,N_16511,N_16710);
nor U17320 (N_17320,N_15938,N_16246);
and U17321 (N_17321,N_16310,N_16554);
and U17322 (N_17322,N_16471,N_16538);
xor U17323 (N_17323,N_15688,N_15672);
nor U17324 (N_17324,N_16376,N_15911);
nor U17325 (N_17325,N_16759,N_15705);
xor U17326 (N_17326,N_15710,N_16505);
or U17327 (N_17327,N_16382,N_15882);
or U17328 (N_17328,N_16542,N_15628);
xnor U17329 (N_17329,N_15903,N_15642);
or U17330 (N_17330,N_15608,N_16332);
xnor U17331 (N_17331,N_16101,N_15669);
nor U17332 (N_17332,N_16098,N_15981);
xnor U17333 (N_17333,N_16130,N_15636);
or U17334 (N_17334,N_15601,N_16599);
nand U17335 (N_17335,N_15904,N_16066);
nand U17336 (N_17336,N_16283,N_15869);
or U17337 (N_17337,N_16289,N_16236);
xnor U17338 (N_17338,N_15745,N_16794);
and U17339 (N_17339,N_16798,N_15674);
xnor U17340 (N_17340,N_16048,N_16769);
nand U17341 (N_17341,N_15876,N_16083);
and U17342 (N_17342,N_16366,N_16414);
nor U17343 (N_17343,N_15983,N_16701);
and U17344 (N_17344,N_15797,N_16780);
or U17345 (N_17345,N_16185,N_15711);
nor U17346 (N_17346,N_16433,N_16001);
or U17347 (N_17347,N_16028,N_15916);
nand U17348 (N_17348,N_15619,N_15824);
nand U17349 (N_17349,N_15620,N_15632);
nor U17350 (N_17350,N_15987,N_15923);
or U17351 (N_17351,N_16540,N_16426);
and U17352 (N_17352,N_16655,N_15693);
xnor U17353 (N_17353,N_15994,N_16319);
xor U17354 (N_17354,N_16133,N_15856);
or U17355 (N_17355,N_16443,N_15875);
nand U17356 (N_17356,N_16312,N_15971);
xnor U17357 (N_17357,N_15635,N_15868);
xnor U17358 (N_17358,N_16608,N_16674);
nor U17359 (N_17359,N_16037,N_16081);
or U17360 (N_17360,N_16331,N_16641);
xor U17361 (N_17361,N_16631,N_16736);
nor U17362 (N_17362,N_15955,N_16536);
and U17363 (N_17363,N_16679,N_16624);
nand U17364 (N_17364,N_16633,N_16658);
nor U17365 (N_17365,N_16137,N_15759);
or U17366 (N_17366,N_16189,N_16779);
xor U17367 (N_17367,N_15834,N_16333);
xor U17368 (N_17368,N_16106,N_15997);
xnor U17369 (N_17369,N_16415,N_16309);
and U17370 (N_17370,N_15888,N_16788);
and U17371 (N_17371,N_16755,N_16385);
and U17372 (N_17372,N_16551,N_16733);
or U17373 (N_17373,N_15839,N_16610);
or U17374 (N_17374,N_16085,N_16186);
or U17375 (N_17375,N_15982,N_16216);
xor U17376 (N_17376,N_15720,N_15933);
or U17377 (N_17377,N_15878,N_16209);
nor U17378 (N_17378,N_16158,N_16320);
and U17379 (N_17379,N_16399,N_15945);
or U17380 (N_17380,N_15763,N_16224);
xor U17381 (N_17381,N_15887,N_16768);
and U17382 (N_17382,N_15791,N_16233);
nand U17383 (N_17383,N_16017,N_16796);
or U17384 (N_17384,N_16225,N_16451);
xnor U17385 (N_17385,N_16579,N_16324);
nand U17386 (N_17386,N_16738,N_16080);
nand U17387 (N_17387,N_16690,N_15767);
nor U17388 (N_17388,N_16581,N_16640);
nor U17389 (N_17389,N_16260,N_15975);
or U17390 (N_17390,N_16429,N_16181);
nand U17391 (N_17391,N_16591,N_15793);
and U17392 (N_17392,N_15622,N_16473);
xnor U17393 (N_17393,N_16067,N_15807);
and U17394 (N_17394,N_16307,N_15604);
nor U17395 (N_17395,N_16369,N_16487);
nor U17396 (N_17396,N_15924,N_16045);
or U17397 (N_17397,N_15775,N_16108);
and U17398 (N_17398,N_16247,N_16403);
and U17399 (N_17399,N_15761,N_16432);
xnor U17400 (N_17400,N_16747,N_16555);
or U17401 (N_17401,N_16006,N_15646);
xor U17402 (N_17402,N_16149,N_15963);
nor U17403 (N_17403,N_15609,N_15908);
xor U17404 (N_17404,N_15699,N_15681);
nor U17405 (N_17405,N_15619,N_16246);
nor U17406 (N_17406,N_16431,N_16550);
xor U17407 (N_17407,N_15893,N_16241);
and U17408 (N_17408,N_15812,N_16338);
and U17409 (N_17409,N_16437,N_16451);
or U17410 (N_17410,N_16691,N_16327);
nand U17411 (N_17411,N_16655,N_16772);
nand U17412 (N_17412,N_16028,N_16754);
or U17413 (N_17413,N_16634,N_15955);
xnor U17414 (N_17414,N_15835,N_15815);
and U17415 (N_17415,N_15778,N_16625);
xor U17416 (N_17416,N_16338,N_16448);
xor U17417 (N_17417,N_16712,N_16062);
nand U17418 (N_17418,N_15714,N_16504);
xor U17419 (N_17419,N_16140,N_15626);
nor U17420 (N_17420,N_15660,N_16506);
nor U17421 (N_17421,N_16448,N_15645);
nand U17422 (N_17422,N_15613,N_15751);
nor U17423 (N_17423,N_16081,N_15677);
nand U17424 (N_17424,N_15756,N_16325);
or U17425 (N_17425,N_16148,N_16330);
xnor U17426 (N_17426,N_16106,N_16322);
or U17427 (N_17427,N_16570,N_16673);
nor U17428 (N_17428,N_16652,N_16119);
xor U17429 (N_17429,N_16744,N_16221);
nand U17430 (N_17430,N_16274,N_16501);
or U17431 (N_17431,N_16334,N_16413);
and U17432 (N_17432,N_15688,N_16158);
nor U17433 (N_17433,N_15769,N_16313);
or U17434 (N_17434,N_16656,N_15866);
and U17435 (N_17435,N_16056,N_16686);
or U17436 (N_17436,N_15920,N_15726);
nor U17437 (N_17437,N_16298,N_16129);
nor U17438 (N_17438,N_16029,N_15997);
nor U17439 (N_17439,N_15750,N_16437);
nand U17440 (N_17440,N_16225,N_15965);
nor U17441 (N_17441,N_16410,N_15900);
or U17442 (N_17442,N_16453,N_16682);
or U17443 (N_17443,N_16418,N_16002);
xor U17444 (N_17444,N_15835,N_16166);
nand U17445 (N_17445,N_15811,N_15601);
or U17446 (N_17446,N_15967,N_16244);
nor U17447 (N_17447,N_16089,N_15964);
xor U17448 (N_17448,N_16405,N_16366);
xor U17449 (N_17449,N_16727,N_15944);
nand U17450 (N_17450,N_15743,N_15847);
and U17451 (N_17451,N_16209,N_16432);
nor U17452 (N_17452,N_15820,N_16515);
nor U17453 (N_17453,N_16635,N_15851);
nor U17454 (N_17454,N_15774,N_15713);
nor U17455 (N_17455,N_15625,N_16153);
or U17456 (N_17456,N_15752,N_15687);
or U17457 (N_17457,N_16410,N_15940);
nand U17458 (N_17458,N_16746,N_15735);
and U17459 (N_17459,N_16212,N_15834);
nor U17460 (N_17460,N_16004,N_16171);
nand U17461 (N_17461,N_16685,N_16478);
nor U17462 (N_17462,N_16542,N_16525);
or U17463 (N_17463,N_15645,N_16062);
or U17464 (N_17464,N_16741,N_16191);
xor U17465 (N_17465,N_16046,N_16357);
xnor U17466 (N_17466,N_16573,N_16094);
xor U17467 (N_17467,N_15679,N_16038);
nand U17468 (N_17468,N_16697,N_16086);
nand U17469 (N_17469,N_16508,N_16289);
xor U17470 (N_17470,N_15761,N_15877);
and U17471 (N_17471,N_16210,N_15734);
or U17472 (N_17472,N_16564,N_15936);
nor U17473 (N_17473,N_16224,N_16512);
xnor U17474 (N_17474,N_16253,N_16044);
nor U17475 (N_17475,N_16325,N_16333);
xnor U17476 (N_17476,N_16771,N_15779);
nor U17477 (N_17477,N_16646,N_15701);
nor U17478 (N_17478,N_16528,N_16078);
or U17479 (N_17479,N_15750,N_16670);
nand U17480 (N_17480,N_15976,N_15951);
nand U17481 (N_17481,N_16251,N_16084);
or U17482 (N_17482,N_15830,N_16088);
nor U17483 (N_17483,N_15656,N_15763);
and U17484 (N_17484,N_16247,N_16569);
or U17485 (N_17485,N_15933,N_16323);
nand U17486 (N_17486,N_16197,N_16015);
xnor U17487 (N_17487,N_16514,N_16268);
nand U17488 (N_17488,N_16184,N_16636);
nor U17489 (N_17489,N_16530,N_16343);
nor U17490 (N_17490,N_15773,N_15663);
nor U17491 (N_17491,N_15869,N_16290);
and U17492 (N_17492,N_16749,N_16744);
nand U17493 (N_17493,N_15791,N_15684);
xnor U17494 (N_17494,N_16581,N_16023);
nand U17495 (N_17495,N_15997,N_16136);
nand U17496 (N_17496,N_15631,N_16363);
and U17497 (N_17497,N_16758,N_16393);
xor U17498 (N_17498,N_15938,N_16043);
xnor U17499 (N_17499,N_16024,N_16429);
nor U17500 (N_17500,N_16556,N_16095);
or U17501 (N_17501,N_16660,N_15757);
nand U17502 (N_17502,N_16438,N_15842);
xor U17503 (N_17503,N_16758,N_15693);
xnor U17504 (N_17504,N_16607,N_15878);
and U17505 (N_17505,N_15930,N_16442);
nand U17506 (N_17506,N_16310,N_15693);
nor U17507 (N_17507,N_16757,N_16117);
xor U17508 (N_17508,N_16644,N_16677);
nor U17509 (N_17509,N_16030,N_16394);
nand U17510 (N_17510,N_16332,N_16768);
nand U17511 (N_17511,N_16785,N_15697);
nand U17512 (N_17512,N_16128,N_15738);
nor U17513 (N_17513,N_16534,N_16196);
nor U17514 (N_17514,N_16668,N_16122);
xnor U17515 (N_17515,N_16052,N_15859);
xor U17516 (N_17516,N_16750,N_15656);
and U17517 (N_17517,N_16141,N_16379);
or U17518 (N_17518,N_15657,N_15608);
or U17519 (N_17519,N_16244,N_16170);
nor U17520 (N_17520,N_16273,N_15755);
or U17521 (N_17521,N_16781,N_16397);
xor U17522 (N_17522,N_16122,N_16578);
xnor U17523 (N_17523,N_15772,N_16095);
nor U17524 (N_17524,N_16331,N_15966);
nor U17525 (N_17525,N_15646,N_16317);
nand U17526 (N_17526,N_16558,N_16337);
and U17527 (N_17527,N_16756,N_16395);
nand U17528 (N_17528,N_15665,N_15740);
and U17529 (N_17529,N_15985,N_15918);
xor U17530 (N_17530,N_16016,N_15991);
nor U17531 (N_17531,N_16186,N_16178);
xnor U17532 (N_17532,N_15810,N_15907);
nor U17533 (N_17533,N_16320,N_16535);
nand U17534 (N_17534,N_16772,N_16273);
xor U17535 (N_17535,N_16363,N_16409);
xor U17536 (N_17536,N_15769,N_16110);
or U17537 (N_17537,N_16520,N_15887);
nand U17538 (N_17538,N_16754,N_15857);
or U17539 (N_17539,N_16002,N_16746);
nor U17540 (N_17540,N_16195,N_15762);
nand U17541 (N_17541,N_16063,N_16675);
nor U17542 (N_17542,N_16585,N_16152);
and U17543 (N_17543,N_16030,N_16331);
nand U17544 (N_17544,N_16051,N_16083);
nand U17545 (N_17545,N_16265,N_16216);
nand U17546 (N_17546,N_15623,N_16020);
nor U17547 (N_17547,N_16220,N_16767);
nand U17548 (N_17548,N_16658,N_15949);
and U17549 (N_17549,N_15995,N_16214);
xor U17550 (N_17550,N_15933,N_16705);
nand U17551 (N_17551,N_16376,N_16760);
nand U17552 (N_17552,N_15992,N_16643);
or U17553 (N_17553,N_16108,N_16329);
and U17554 (N_17554,N_15702,N_16547);
or U17555 (N_17555,N_16521,N_16786);
xor U17556 (N_17556,N_16502,N_16727);
nand U17557 (N_17557,N_16264,N_15789);
or U17558 (N_17558,N_16407,N_16050);
xnor U17559 (N_17559,N_16283,N_16342);
and U17560 (N_17560,N_16299,N_15828);
and U17561 (N_17561,N_16629,N_16336);
and U17562 (N_17562,N_16337,N_16054);
or U17563 (N_17563,N_16425,N_15724);
and U17564 (N_17564,N_15643,N_15950);
or U17565 (N_17565,N_16423,N_16142);
and U17566 (N_17566,N_15924,N_15980);
nor U17567 (N_17567,N_16572,N_16160);
or U17568 (N_17568,N_16205,N_16308);
and U17569 (N_17569,N_16423,N_16282);
nor U17570 (N_17570,N_15680,N_16514);
or U17571 (N_17571,N_16767,N_16063);
nor U17572 (N_17572,N_15969,N_16178);
nand U17573 (N_17573,N_15801,N_16376);
xor U17574 (N_17574,N_15671,N_16735);
and U17575 (N_17575,N_16586,N_15629);
xnor U17576 (N_17576,N_16055,N_16398);
or U17577 (N_17577,N_15902,N_15710);
xnor U17578 (N_17578,N_16366,N_15937);
nor U17579 (N_17579,N_15628,N_15774);
nand U17580 (N_17580,N_15907,N_15735);
nor U17581 (N_17581,N_16312,N_16692);
xor U17582 (N_17582,N_16405,N_16657);
xor U17583 (N_17583,N_15661,N_16679);
nand U17584 (N_17584,N_15634,N_16093);
nand U17585 (N_17585,N_16214,N_16086);
xnor U17586 (N_17586,N_16075,N_16344);
nand U17587 (N_17587,N_16476,N_16439);
nand U17588 (N_17588,N_16067,N_16769);
nand U17589 (N_17589,N_15737,N_16072);
nand U17590 (N_17590,N_15728,N_16558);
or U17591 (N_17591,N_16592,N_16653);
and U17592 (N_17592,N_15929,N_16294);
and U17593 (N_17593,N_15642,N_16237);
or U17594 (N_17594,N_16574,N_16668);
and U17595 (N_17595,N_16507,N_15733);
nor U17596 (N_17596,N_15891,N_16375);
or U17597 (N_17597,N_15651,N_16741);
and U17598 (N_17598,N_15761,N_15735);
or U17599 (N_17599,N_16523,N_16233);
and U17600 (N_17600,N_16395,N_16102);
or U17601 (N_17601,N_15652,N_16380);
or U17602 (N_17602,N_16687,N_16392);
xnor U17603 (N_17603,N_15623,N_16452);
nand U17604 (N_17604,N_16611,N_16358);
nor U17605 (N_17605,N_15808,N_16605);
xnor U17606 (N_17606,N_15837,N_16525);
xor U17607 (N_17607,N_15848,N_15911);
nand U17608 (N_17608,N_16762,N_16792);
or U17609 (N_17609,N_15726,N_16266);
nor U17610 (N_17610,N_16200,N_15816);
and U17611 (N_17611,N_16124,N_16500);
and U17612 (N_17612,N_16646,N_16661);
and U17613 (N_17613,N_16352,N_16054);
xnor U17614 (N_17614,N_16242,N_16614);
xor U17615 (N_17615,N_15901,N_16129);
or U17616 (N_17616,N_16506,N_16050);
or U17617 (N_17617,N_16371,N_16076);
nand U17618 (N_17618,N_15909,N_15642);
and U17619 (N_17619,N_16555,N_16630);
and U17620 (N_17620,N_16485,N_16087);
and U17621 (N_17621,N_15658,N_15928);
xnor U17622 (N_17622,N_16650,N_16198);
and U17623 (N_17623,N_16775,N_16067);
or U17624 (N_17624,N_15951,N_15743);
and U17625 (N_17625,N_15868,N_15840);
nor U17626 (N_17626,N_16354,N_16550);
xnor U17627 (N_17627,N_16631,N_16129);
xor U17628 (N_17628,N_15646,N_16415);
and U17629 (N_17629,N_16721,N_15750);
or U17630 (N_17630,N_16351,N_15824);
nand U17631 (N_17631,N_15920,N_16575);
and U17632 (N_17632,N_16480,N_16576);
nor U17633 (N_17633,N_16511,N_16613);
or U17634 (N_17634,N_16342,N_15606);
and U17635 (N_17635,N_16366,N_16766);
and U17636 (N_17636,N_15649,N_16293);
xor U17637 (N_17637,N_16296,N_15750);
nand U17638 (N_17638,N_15617,N_16526);
nand U17639 (N_17639,N_15903,N_16345);
nor U17640 (N_17640,N_15941,N_16335);
xnor U17641 (N_17641,N_15914,N_15894);
xnor U17642 (N_17642,N_16018,N_16797);
or U17643 (N_17643,N_15707,N_16322);
xnor U17644 (N_17644,N_15741,N_16431);
and U17645 (N_17645,N_16158,N_15763);
xor U17646 (N_17646,N_16058,N_16507);
and U17647 (N_17647,N_16473,N_16547);
nor U17648 (N_17648,N_16226,N_16791);
or U17649 (N_17649,N_16509,N_15725);
and U17650 (N_17650,N_16516,N_16284);
or U17651 (N_17651,N_16667,N_16410);
or U17652 (N_17652,N_15671,N_16157);
and U17653 (N_17653,N_16503,N_16284);
and U17654 (N_17654,N_16609,N_16724);
or U17655 (N_17655,N_16488,N_16645);
xnor U17656 (N_17656,N_16276,N_16028);
xnor U17657 (N_17657,N_16738,N_16559);
nand U17658 (N_17658,N_16782,N_15939);
nor U17659 (N_17659,N_15864,N_16478);
xnor U17660 (N_17660,N_16410,N_16794);
xor U17661 (N_17661,N_15660,N_16676);
nor U17662 (N_17662,N_16377,N_15999);
nor U17663 (N_17663,N_16282,N_16327);
nor U17664 (N_17664,N_16161,N_15718);
nand U17665 (N_17665,N_15723,N_16541);
xor U17666 (N_17666,N_15819,N_16275);
or U17667 (N_17667,N_16629,N_15696);
xnor U17668 (N_17668,N_16360,N_16753);
nor U17669 (N_17669,N_16543,N_16271);
nand U17670 (N_17670,N_15879,N_16437);
xnor U17671 (N_17671,N_16239,N_16721);
nand U17672 (N_17672,N_16322,N_15777);
nand U17673 (N_17673,N_16778,N_16308);
and U17674 (N_17674,N_16620,N_16305);
and U17675 (N_17675,N_16277,N_16378);
xor U17676 (N_17676,N_16127,N_15635);
and U17677 (N_17677,N_16299,N_16013);
nor U17678 (N_17678,N_16412,N_16465);
or U17679 (N_17679,N_15625,N_16327);
xor U17680 (N_17680,N_16590,N_16248);
xnor U17681 (N_17681,N_16683,N_15712);
xnor U17682 (N_17682,N_16492,N_16003);
xor U17683 (N_17683,N_15833,N_16348);
nor U17684 (N_17684,N_16074,N_16523);
nor U17685 (N_17685,N_15627,N_16346);
xnor U17686 (N_17686,N_15890,N_16409);
nand U17687 (N_17687,N_16322,N_16051);
xnor U17688 (N_17688,N_16138,N_16537);
nor U17689 (N_17689,N_15615,N_15836);
nand U17690 (N_17690,N_16155,N_15998);
and U17691 (N_17691,N_16036,N_16295);
nor U17692 (N_17692,N_15650,N_16186);
or U17693 (N_17693,N_15752,N_16734);
nor U17694 (N_17694,N_16089,N_16332);
xnor U17695 (N_17695,N_16242,N_15703);
or U17696 (N_17696,N_16382,N_16579);
or U17697 (N_17697,N_15730,N_15965);
nand U17698 (N_17698,N_15654,N_16175);
xor U17699 (N_17699,N_16528,N_15996);
or U17700 (N_17700,N_16406,N_16041);
and U17701 (N_17701,N_16409,N_15613);
nor U17702 (N_17702,N_16550,N_16242);
or U17703 (N_17703,N_15643,N_15936);
nand U17704 (N_17704,N_16471,N_16294);
nor U17705 (N_17705,N_16674,N_16214);
nor U17706 (N_17706,N_16481,N_16342);
nor U17707 (N_17707,N_15663,N_16514);
xor U17708 (N_17708,N_16198,N_15716);
nor U17709 (N_17709,N_16774,N_16672);
nand U17710 (N_17710,N_16742,N_15641);
and U17711 (N_17711,N_16508,N_15657);
nand U17712 (N_17712,N_16260,N_16077);
nor U17713 (N_17713,N_15831,N_16651);
xor U17714 (N_17714,N_16044,N_16335);
or U17715 (N_17715,N_16640,N_15634);
or U17716 (N_17716,N_16439,N_16521);
xnor U17717 (N_17717,N_16242,N_16202);
and U17718 (N_17718,N_16153,N_15737);
and U17719 (N_17719,N_15841,N_16134);
and U17720 (N_17720,N_15637,N_16646);
xor U17721 (N_17721,N_15716,N_16373);
xnor U17722 (N_17722,N_16143,N_15866);
and U17723 (N_17723,N_16395,N_15802);
or U17724 (N_17724,N_15712,N_16421);
or U17725 (N_17725,N_16150,N_16578);
nand U17726 (N_17726,N_16255,N_15951);
or U17727 (N_17727,N_15615,N_15843);
or U17728 (N_17728,N_16246,N_16668);
or U17729 (N_17729,N_16313,N_15759);
or U17730 (N_17730,N_16085,N_16090);
or U17731 (N_17731,N_16530,N_16433);
xnor U17732 (N_17732,N_16607,N_16113);
and U17733 (N_17733,N_16262,N_15746);
nor U17734 (N_17734,N_16509,N_15743);
and U17735 (N_17735,N_16742,N_16717);
nor U17736 (N_17736,N_16583,N_15683);
nor U17737 (N_17737,N_16383,N_15839);
xnor U17738 (N_17738,N_16765,N_15904);
nand U17739 (N_17739,N_16051,N_15724);
and U17740 (N_17740,N_16098,N_15787);
and U17741 (N_17741,N_15632,N_16733);
nand U17742 (N_17742,N_16275,N_16026);
or U17743 (N_17743,N_16430,N_16772);
xor U17744 (N_17744,N_15672,N_15943);
nor U17745 (N_17745,N_16474,N_16262);
or U17746 (N_17746,N_16044,N_16635);
nor U17747 (N_17747,N_16568,N_16135);
and U17748 (N_17748,N_16269,N_16407);
nor U17749 (N_17749,N_16226,N_16587);
or U17750 (N_17750,N_15934,N_16156);
or U17751 (N_17751,N_16682,N_16721);
xor U17752 (N_17752,N_16174,N_16248);
nor U17753 (N_17753,N_16439,N_16430);
or U17754 (N_17754,N_15737,N_16365);
and U17755 (N_17755,N_15658,N_15629);
nor U17756 (N_17756,N_15758,N_16139);
xor U17757 (N_17757,N_16057,N_15610);
or U17758 (N_17758,N_15622,N_16009);
or U17759 (N_17759,N_16134,N_15737);
nor U17760 (N_17760,N_15925,N_16716);
or U17761 (N_17761,N_16470,N_15766);
nand U17762 (N_17762,N_16446,N_16018);
xnor U17763 (N_17763,N_16757,N_15958);
nand U17764 (N_17764,N_16430,N_16149);
nor U17765 (N_17765,N_16146,N_15932);
or U17766 (N_17766,N_15926,N_16521);
or U17767 (N_17767,N_16291,N_16602);
or U17768 (N_17768,N_15885,N_15820);
or U17769 (N_17769,N_16029,N_15933);
nor U17770 (N_17770,N_15669,N_16276);
or U17771 (N_17771,N_16778,N_15624);
or U17772 (N_17772,N_16268,N_15614);
nor U17773 (N_17773,N_16370,N_16364);
or U17774 (N_17774,N_16655,N_15785);
or U17775 (N_17775,N_16608,N_16556);
and U17776 (N_17776,N_16208,N_16569);
or U17777 (N_17777,N_16592,N_16233);
or U17778 (N_17778,N_16625,N_16671);
and U17779 (N_17779,N_15968,N_16158);
or U17780 (N_17780,N_16653,N_15911);
and U17781 (N_17781,N_16643,N_16040);
or U17782 (N_17782,N_15600,N_16340);
or U17783 (N_17783,N_15852,N_15671);
nand U17784 (N_17784,N_16708,N_15699);
xnor U17785 (N_17785,N_15698,N_15900);
nor U17786 (N_17786,N_15676,N_16545);
nand U17787 (N_17787,N_16546,N_16563);
nor U17788 (N_17788,N_15933,N_16338);
or U17789 (N_17789,N_16020,N_16705);
nand U17790 (N_17790,N_16063,N_15842);
or U17791 (N_17791,N_15968,N_15894);
and U17792 (N_17792,N_16082,N_16425);
or U17793 (N_17793,N_16000,N_16777);
or U17794 (N_17794,N_16380,N_16044);
and U17795 (N_17795,N_15909,N_15942);
nor U17796 (N_17796,N_15686,N_16514);
nand U17797 (N_17797,N_16668,N_16630);
nand U17798 (N_17798,N_15747,N_16017);
nor U17799 (N_17799,N_15817,N_15934);
nor U17800 (N_17800,N_16044,N_15975);
or U17801 (N_17801,N_16045,N_16032);
xor U17802 (N_17802,N_16348,N_15984);
or U17803 (N_17803,N_16144,N_16602);
or U17804 (N_17804,N_16166,N_16456);
nand U17805 (N_17805,N_16618,N_16000);
or U17806 (N_17806,N_16769,N_16603);
or U17807 (N_17807,N_15946,N_16142);
nand U17808 (N_17808,N_16322,N_16779);
or U17809 (N_17809,N_15886,N_15788);
nor U17810 (N_17810,N_16196,N_16059);
xnor U17811 (N_17811,N_15675,N_15774);
or U17812 (N_17812,N_16342,N_16282);
and U17813 (N_17813,N_16751,N_16573);
and U17814 (N_17814,N_16792,N_15967);
xor U17815 (N_17815,N_16635,N_15747);
and U17816 (N_17816,N_16334,N_16381);
xnor U17817 (N_17817,N_16312,N_16759);
nor U17818 (N_17818,N_16213,N_15732);
and U17819 (N_17819,N_16666,N_16340);
or U17820 (N_17820,N_16549,N_15836);
nor U17821 (N_17821,N_16043,N_16482);
xor U17822 (N_17822,N_16078,N_16331);
xnor U17823 (N_17823,N_16153,N_16598);
nor U17824 (N_17824,N_16472,N_16164);
xnor U17825 (N_17825,N_15644,N_15779);
nand U17826 (N_17826,N_16667,N_15689);
xnor U17827 (N_17827,N_16777,N_16068);
nand U17828 (N_17828,N_16605,N_16614);
or U17829 (N_17829,N_16164,N_15962);
xor U17830 (N_17830,N_16467,N_15740);
nor U17831 (N_17831,N_16628,N_16380);
and U17832 (N_17832,N_16328,N_16207);
or U17833 (N_17833,N_16129,N_16127);
nand U17834 (N_17834,N_15766,N_16488);
xnor U17835 (N_17835,N_16363,N_15690);
xor U17836 (N_17836,N_16681,N_16160);
nand U17837 (N_17837,N_16629,N_16774);
xnor U17838 (N_17838,N_16112,N_16199);
xor U17839 (N_17839,N_16749,N_15936);
and U17840 (N_17840,N_16737,N_15955);
and U17841 (N_17841,N_16511,N_16344);
and U17842 (N_17842,N_16004,N_15894);
xor U17843 (N_17843,N_15825,N_15784);
or U17844 (N_17844,N_15824,N_16225);
nor U17845 (N_17845,N_16287,N_15683);
nor U17846 (N_17846,N_16381,N_16152);
and U17847 (N_17847,N_15685,N_15952);
nand U17848 (N_17848,N_16161,N_16560);
xnor U17849 (N_17849,N_16571,N_16007);
nor U17850 (N_17850,N_16212,N_16036);
nor U17851 (N_17851,N_16101,N_15849);
and U17852 (N_17852,N_16518,N_16298);
xnor U17853 (N_17853,N_16683,N_16789);
and U17854 (N_17854,N_15708,N_16790);
nand U17855 (N_17855,N_16307,N_15764);
or U17856 (N_17856,N_16591,N_15944);
nand U17857 (N_17857,N_15637,N_16701);
and U17858 (N_17858,N_16369,N_16242);
nor U17859 (N_17859,N_16338,N_16247);
nand U17860 (N_17860,N_16403,N_16576);
nor U17861 (N_17861,N_15603,N_16325);
nor U17862 (N_17862,N_16594,N_16265);
nor U17863 (N_17863,N_15908,N_16342);
xnor U17864 (N_17864,N_16476,N_15684);
or U17865 (N_17865,N_16792,N_15758);
nor U17866 (N_17866,N_15778,N_16478);
nand U17867 (N_17867,N_16502,N_15781);
or U17868 (N_17868,N_16701,N_16731);
nand U17869 (N_17869,N_15845,N_16536);
nand U17870 (N_17870,N_16537,N_15925);
and U17871 (N_17871,N_15604,N_15672);
and U17872 (N_17872,N_16431,N_16751);
nand U17873 (N_17873,N_16168,N_16418);
or U17874 (N_17874,N_16522,N_15695);
xnor U17875 (N_17875,N_16732,N_16629);
and U17876 (N_17876,N_15823,N_15751);
and U17877 (N_17877,N_15885,N_15663);
xnor U17878 (N_17878,N_16775,N_15668);
nor U17879 (N_17879,N_16770,N_16679);
or U17880 (N_17880,N_15864,N_16208);
nand U17881 (N_17881,N_16605,N_16405);
or U17882 (N_17882,N_15965,N_16070);
nand U17883 (N_17883,N_16303,N_16506);
and U17884 (N_17884,N_16053,N_15950);
xnor U17885 (N_17885,N_15636,N_16098);
nand U17886 (N_17886,N_16003,N_16369);
and U17887 (N_17887,N_15769,N_16410);
xnor U17888 (N_17888,N_16789,N_16390);
and U17889 (N_17889,N_16067,N_15648);
and U17890 (N_17890,N_16540,N_16706);
xnor U17891 (N_17891,N_15898,N_16664);
xor U17892 (N_17892,N_16009,N_15793);
and U17893 (N_17893,N_16273,N_16458);
nor U17894 (N_17894,N_15618,N_15936);
and U17895 (N_17895,N_16029,N_16631);
xnor U17896 (N_17896,N_16681,N_15874);
nand U17897 (N_17897,N_16315,N_16129);
nor U17898 (N_17898,N_16653,N_15611);
nand U17899 (N_17899,N_15670,N_16643);
and U17900 (N_17900,N_16398,N_16376);
xor U17901 (N_17901,N_15696,N_15662);
xnor U17902 (N_17902,N_15684,N_16575);
or U17903 (N_17903,N_16680,N_15826);
xnor U17904 (N_17904,N_15829,N_15777);
nand U17905 (N_17905,N_15821,N_15865);
nand U17906 (N_17906,N_16230,N_16189);
xor U17907 (N_17907,N_15823,N_15613);
or U17908 (N_17908,N_16677,N_16580);
and U17909 (N_17909,N_15896,N_15636);
xor U17910 (N_17910,N_15626,N_16056);
xnor U17911 (N_17911,N_16697,N_16282);
nor U17912 (N_17912,N_16564,N_16505);
xor U17913 (N_17913,N_15965,N_16093);
xor U17914 (N_17914,N_16731,N_15836);
or U17915 (N_17915,N_15677,N_16790);
nor U17916 (N_17916,N_16068,N_16066);
and U17917 (N_17917,N_16775,N_15664);
nor U17918 (N_17918,N_16405,N_16571);
or U17919 (N_17919,N_16193,N_15872);
or U17920 (N_17920,N_16311,N_15672);
nor U17921 (N_17921,N_15702,N_16037);
or U17922 (N_17922,N_16676,N_16004);
and U17923 (N_17923,N_16546,N_16220);
nor U17924 (N_17924,N_16047,N_16247);
nand U17925 (N_17925,N_15977,N_16321);
and U17926 (N_17926,N_16776,N_15878);
nor U17927 (N_17927,N_15981,N_16489);
and U17928 (N_17928,N_16603,N_16616);
nor U17929 (N_17929,N_16046,N_16380);
and U17930 (N_17930,N_16571,N_16520);
nor U17931 (N_17931,N_16312,N_15661);
or U17932 (N_17932,N_15663,N_15840);
nor U17933 (N_17933,N_16449,N_16632);
or U17934 (N_17934,N_16344,N_16473);
nand U17935 (N_17935,N_16426,N_15803);
nor U17936 (N_17936,N_16660,N_15822);
xnor U17937 (N_17937,N_16093,N_16191);
nor U17938 (N_17938,N_16380,N_15858);
nor U17939 (N_17939,N_15979,N_16271);
or U17940 (N_17940,N_16433,N_16417);
and U17941 (N_17941,N_16501,N_16515);
nand U17942 (N_17942,N_16056,N_16110);
nand U17943 (N_17943,N_16404,N_15860);
nand U17944 (N_17944,N_16614,N_16458);
and U17945 (N_17945,N_16339,N_16276);
nor U17946 (N_17946,N_15935,N_15904);
nor U17947 (N_17947,N_16425,N_15742);
nor U17948 (N_17948,N_16703,N_16699);
xor U17949 (N_17949,N_16369,N_16776);
or U17950 (N_17950,N_15880,N_15732);
xnor U17951 (N_17951,N_15788,N_16254);
nor U17952 (N_17952,N_16198,N_16392);
nor U17953 (N_17953,N_16062,N_16432);
or U17954 (N_17954,N_16176,N_16702);
nor U17955 (N_17955,N_16123,N_15710);
and U17956 (N_17956,N_16622,N_16667);
nand U17957 (N_17957,N_16121,N_16482);
xor U17958 (N_17958,N_16125,N_16482);
nand U17959 (N_17959,N_16227,N_16695);
nor U17960 (N_17960,N_16767,N_15781);
nand U17961 (N_17961,N_16481,N_15696);
nor U17962 (N_17962,N_15664,N_16356);
or U17963 (N_17963,N_16034,N_16613);
or U17964 (N_17964,N_16039,N_15903);
nand U17965 (N_17965,N_15685,N_15679);
and U17966 (N_17966,N_16412,N_16322);
nand U17967 (N_17967,N_16650,N_16148);
xnor U17968 (N_17968,N_16566,N_16036);
nor U17969 (N_17969,N_15805,N_15756);
xor U17970 (N_17970,N_16731,N_16687);
nor U17971 (N_17971,N_15766,N_15813);
nand U17972 (N_17972,N_16346,N_16398);
nor U17973 (N_17973,N_15989,N_16489);
or U17974 (N_17974,N_16089,N_16693);
and U17975 (N_17975,N_16192,N_16527);
nor U17976 (N_17976,N_16770,N_16080);
or U17977 (N_17977,N_15850,N_16337);
and U17978 (N_17978,N_16035,N_16442);
nand U17979 (N_17979,N_15985,N_16232);
xnor U17980 (N_17980,N_15603,N_16009);
nor U17981 (N_17981,N_16009,N_15600);
nand U17982 (N_17982,N_16374,N_15799);
nand U17983 (N_17983,N_16502,N_15961);
nand U17984 (N_17984,N_16392,N_15632);
nand U17985 (N_17985,N_16476,N_16230);
or U17986 (N_17986,N_16517,N_16635);
or U17987 (N_17987,N_16701,N_15922);
xor U17988 (N_17988,N_16730,N_16657);
nand U17989 (N_17989,N_15785,N_16437);
or U17990 (N_17990,N_16480,N_16219);
and U17991 (N_17991,N_16473,N_16282);
xnor U17992 (N_17992,N_15886,N_16262);
or U17993 (N_17993,N_15680,N_16605);
nand U17994 (N_17994,N_16628,N_15769);
xnor U17995 (N_17995,N_16631,N_15995);
or U17996 (N_17996,N_15693,N_16666);
xnor U17997 (N_17997,N_15830,N_16115);
nor U17998 (N_17998,N_15807,N_15875);
xnor U17999 (N_17999,N_16286,N_16639);
nor U18000 (N_18000,N_17446,N_16998);
or U18001 (N_18001,N_17602,N_17284);
nand U18002 (N_18002,N_17965,N_17175);
nand U18003 (N_18003,N_17991,N_17226);
or U18004 (N_18004,N_17621,N_17527);
nand U18005 (N_18005,N_17056,N_17263);
and U18006 (N_18006,N_17940,N_17320);
and U18007 (N_18007,N_17456,N_17638);
or U18008 (N_18008,N_17964,N_17029);
or U18009 (N_18009,N_17630,N_16867);
and U18010 (N_18010,N_17726,N_17240);
and U18011 (N_18011,N_17406,N_17619);
xnor U18012 (N_18012,N_17594,N_17058);
nand U18013 (N_18013,N_17738,N_17506);
and U18014 (N_18014,N_16871,N_17332);
nand U18015 (N_18015,N_17064,N_16877);
and U18016 (N_18016,N_17422,N_17835);
or U18017 (N_18017,N_17612,N_17842);
or U18018 (N_18018,N_16814,N_17901);
nor U18019 (N_18019,N_17626,N_17909);
and U18020 (N_18020,N_16819,N_17458);
nor U18021 (N_18021,N_17079,N_16833);
xor U18022 (N_18022,N_17720,N_17063);
xor U18023 (N_18023,N_17545,N_17611);
and U18024 (N_18024,N_16806,N_16995);
nor U18025 (N_18025,N_17822,N_17762);
and U18026 (N_18026,N_17742,N_17454);
xnor U18027 (N_18027,N_17334,N_17518);
nand U18028 (N_18028,N_17059,N_16807);
or U18029 (N_18029,N_17546,N_17248);
or U18030 (N_18030,N_17255,N_17864);
and U18031 (N_18031,N_17461,N_17607);
and U18032 (N_18032,N_17870,N_17409);
xor U18033 (N_18033,N_17010,N_17717);
or U18034 (N_18034,N_17593,N_17968);
and U18035 (N_18035,N_16878,N_17729);
or U18036 (N_18036,N_17140,N_17862);
nor U18037 (N_18037,N_17733,N_17889);
and U18038 (N_18038,N_17953,N_17865);
nand U18039 (N_18039,N_16853,N_17283);
nor U18040 (N_18040,N_17447,N_17294);
or U18041 (N_18041,N_16977,N_17844);
and U18042 (N_18042,N_16868,N_17723);
or U18043 (N_18043,N_17500,N_17754);
and U18044 (N_18044,N_17774,N_17945);
and U18045 (N_18045,N_17755,N_17061);
and U18046 (N_18046,N_17904,N_17526);
nor U18047 (N_18047,N_17082,N_17736);
and U18048 (N_18048,N_17978,N_17162);
or U18049 (N_18049,N_17948,N_17974);
and U18050 (N_18050,N_17687,N_17540);
nand U18051 (N_18051,N_17715,N_17967);
nand U18052 (N_18052,N_17150,N_17507);
or U18053 (N_18053,N_17353,N_17396);
xor U18054 (N_18054,N_17917,N_17452);
xor U18055 (N_18055,N_17615,N_17371);
or U18056 (N_18056,N_17293,N_16930);
or U18057 (N_18057,N_17884,N_17695);
nor U18058 (N_18058,N_16834,N_17759);
and U18059 (N_18059,N_16820,N_17138);
nand U18060 (N_18060,N_17793,N_17823);
or U18061 (N_18061,N_17208,N_16932);
or U18062 (N_18062,N_17743,N_17647);
nor U18063 (N_18063,N_17342,N_17051);
nor U18064 (N_18064,N_17840,N_17516);
nand U18065 (N_18065,N_17004,N_17400);
nand U18066 (N_18066,N_17741,N_17510);
nor U18067 (N_18067,N_17876,N_17142);
nor U18068 (N_18068,N_16831,N_17337);
and U18069 (N_18069,N_17942,N_17700);
and U18070 (N_18070,N_17411,N_17556);
and U18071 (N_18071,N_17165,N_16966);
and U18072 (N_18072,N_17013,N_16881);
or U18073 (N_18073,N_17766,N_16911);
xnor U18074 (N_18074,N_17369,N_17827);
and U18075 (N_18075,N_17895,N_17387);
nand U18076 (N_18076,N_17368,N_17662);
or U18077 (N_18077,N_17075,N_17984);
nor U18078 (N_18078,N_17437,N_16988);
xnor U18079 (N_18079,N_17911,N_17218);
nor U18080 (N_18080,N_17882,N_17204);
or U18081 (N_18081,N_17781,N_17443);
and U18082 (N_18082,N_17684,N_17280);
nand U18083 (N_18083,N_17405,N_16989);
and U18084 (N_18084,N_17017,N_17250);
xnor U18085 (N_18085,N_17644,N_17583);
nand U18086 (N_18086,N_16990,N_17114);
and U18087 (N_18087,N_17584,N_17777);
xor U18088 (N_18088,N_17314,N_17886);
or U18089 (N_18089,N_16943,N_16953);
and U18090 (N_18090,N_17676,N_17980);
and U18091 (N_18091,N_17273,N_17853);
and U18092 (N_18092,N_17893,N_17734);
xnor U18093 (N_18093,N_17773,N_17892);
nor U18094 (N_18094,N_17600,N_17290);
and U18095 (N_18095,N_17905,N_17989);
or U18096 (N_18096,N_17983,N_17450);
or U18097 (N_18097,N_17277,N_16817);
or U18098 (N_18098,N_17748,N_17832);
or U18099 (N_18099,N_17377,N_17955);
xor U18100 (N_18100,N_17499,N_16969);
and U18101 (N_18101,N_17995,N_16958);
xnor U18102 (N_18102,N_17223,N_17249);
xor U18103 (N_18103,N_17836,N_16981);
or U18104 (N_18104,N_17306,N_17419);
or U18105 (N_18105,N_17330,N_17264);
nor U18106 (N_18106,N_17515,N_17310);
nor U18107 (N_18107,N_17372,N_17744);
and U18108 (N_18108,N_17303,N_17811);
nor U18109 (N_18109,N_17451,N_16937);
or U18110 (N_18110,N_16909,N_17993);
xor U18111 (N_18111,N_17694,N_17603);
xnor U18112 (N_18112,N_16948,N_17153);
xnor U18113 (N_18113,N_17821,N_17923);
and U18114 (N_18114,N_16964,N_16876);
nor U18115 (N_18115,N_17408,N_17573);
nor U18116 (N_18116,N_17708,N_17160);
or U18117 (N_18117,N_17768,N_16847);
or U18118 (N_18118,N_17636,N_17598);
xnor U18119 (N_18119,N_17522,N_17957);
nor U18120 (N_18120,N_16912,N_17164);
xor U18121 (N_18121,N_17077,N_17872);
nand U18122 (N_18122,N_17008,N_17107);
and U18123 (N_18123,N_17686,N_17365);
nor U18124 (N_18124,N_17815,N_16846);
nand U18125 (N_18125,N_17501,N_17691);
or U18126 (N_18126,N_16974,N_17286);
nor U18127 (N_18127,N_17156,N_17807);
and U18128 (N_18128,N_17632,N_17792);
nand U18129 (N_18129,N_16890,N_17509);
or U18130 (N_18130,N_17351,N_17331);
nor U18131 (N_18131,N_17413,N_17109);
or U18132 (N_18132,N_17641,N_17355);
xor U18133 (N_18133,N_17426,N_16946);
or U18134 (N_18134,N_16852,N_17261);
and U18135 (N_18135,N_17015,N_17994);
xor U18136 (N_18136,N_17401,N_16918);
and U18137 (N_18137,N_17790,N_17505);
or U18138 (N_18138,N_17267,N_17613);
xnor U18139 (N_18139,N_17112,N_17639);
nand U18140 (N_18140,N_17242,N_17958);
or U18141 (N_18141,N_17854,N_16900);
nand U18142 (N_18142,N_16844,N_17855);
nand U18143 (N_18143,N_17992,N_17770);
nor U18144 (N_18144,N_17460,N_17683);
nor U18145 (N_18145,N_17572,N_17867);
and U18146 (N_18146,N_17378,N_17000);
or U18147 (N_18147,N_17243,N_17701);
nand U18148 (N_18148,N_16997,N_17473);
and U18149 (N_18149,N_17122,N_17035);
xor U18150 (N_18150,N_17234,N_17099);
nand U18151 (N_18151,N_17169,N_17541);
xor U18152 (N_18152,N_17783,N_16804);
nand U18153 (N_18153,N_17589,N_17352);
and U18154 (N_18154,N_17534,N_17433);
or U18155 (N_18155,N_17563,N_17794);
or U18156 (N_18156,N_17788,N_17495);
and U18157 (N_18157,N_17824,N_17588);
or U18158 (N_18158,N_17217,N_17431);
nand U18159 (N_18159,N_17739,N_17336);
xor U18160 (N_18160,N_17459,N_17067);
or U18161 (N_18161,N_17610,N_17969);
or U18162 (N_18162,N_17578,N_16872);
or U18163 (N_18163,N_17279,N_16942);
nor U18164 (N_18164,N_17721,N_16805);
and U18165 (N_18165,N_16848,N_17629);
nand U18166 (N_18166,N_17007,N_17073);
and U18167 (N_18167,N_16869,N_17281);
or U18168 (N_18168,N_17906,N_17846);
or U18169 (N_18169,N_16983,N_17430);
xnor U18170 (N_18170,N_17599,N_17653);
nor U18171 (N_18171,N_17129,N_17078);
nor U18172 (N_18172,N_17260,N_17211);
nor U18173 (N_18173,N_17549,N_17758);
nand U18174 (N_18174,N_17564,N_17577);
and U18175 (N_18175,N_17554,N_16827);
or U18176 (N_18176,N_16984,N_17222);
and U18177 (N_18177,N_17699,N_17069);
nor U18178 (N_18178,N_17338,N_17944);
xnor U18179 (N_18179,N_16919,N_17055);
xor U18180 (N_18180,N_17436,N_17977);
and U18181 (N_18181,N_16813,N_17309);
and U18182 (N_18182,N_16886,N_16945);
xor U18183 (N_18183,N_16841,N_16873);
and U18184 (N_18184,N_17535,N_17085);
nor U18185 (N_18185,N_16825,N_17354);
nand U18186 (N_18186,N_17490,N_17463);
nand U18187 (N_18187,N_17786,N_17671);
and U18188 (N_18188,N_16901,N_16856);
or U18189 (N_18189,N_17110,N_17558);
and U18190 (N_18190,N_17252,N_17998);
or U18191 (N_18191,N_17557,N_16824);
and U18192 (N_18192,N_16896,N_17825);
nor U18193 (N_18193,N_17296,N_16957);
xnor U18194 (N_18194,N_17388,N_17435);
nor U18195 (N_18195,N_17609,N_17206);
nand U18196 (N_18196,N_17019,N_17220);
xnor U18197 (N_18197,N_17034,N_17343);
or U18198 (N_18198,N_16888,N_16987);
and U18199 (N_18199,N_16811,N_17951);
or U18200 (N_18200,N_16816,N_16913);
xor U18201 (N_18201,N_17943,N_17254);
and U18202 (N_18202,N_17302,N_17414);
and U18203 (N_18203,N_17919,N_17348);
and U18204 (N_18204,N_17601,N_17221);
xor U18205 (N_18205,N_17032,N_17869);
nor U18206 (N_18206,N_17767,N_17914);
nand U18207 (N_18207,N_17925,N_17665);
xor U18208 (N_18208,N_17763,N_17673);
and U18209 (N_18209,N_17272,N_17213);
nand U18210 (N_18210,N_17997,N_16991);
and U18211 (N_18211,N_17520,N_17776);
and U18212 (N_18212,N_17384,N_17125);
and U18213 (N_18213,N_17706,N_17861);
or U18214 (N_18214,N_16933,N_17933);
and U18215 (N_18215,N_16916,N_16972);
nor U18216 (N_18216,N_17265,N_17299);
and U18217 (N_18217,N_17488,N_17144);
xnor U18218 (N_18218,N_17480,N_17782);
xnor U18219 (N_18219,N_17804,N_16879);
xor U18220 (N_18220,N_17567,N_17448);
or U18221 (N_18221,N_17237,N_16979);
or U18222 (N_18222,N_17143,N_17319);
xnor U18223 (N_18223,N_17778,N_17429);
xnor U18224 (N_18224,N_17858,N_17643);
nor U18225 (N_18225,N_17166,N_17875);
nor U18226 (N_18226,N_17379,N_17816);
nand U18227 (N_18227,N_16949,N_17373);
nor U18228 (N_18228,N_17819,N_17714);
xnor U18229 (N_18229,N_17561,N_17271);
nor U18230 (N_18230,N_16838,N_17952);
nor U18231 (N_18231,N_17344,N_16928);
nor U18232 (N_18232,N_17145,N_16892);
nand U18233 (N_18233,N_16818,N_17115);
nand U18234 (N_18234,N_17954,N_17120);
and U18235 (N_18235,N_17591,N_17266);
nor U18236 (N_18236,N_16927,N_17938);
nor U18237 (N_18237,N_17627,N_17618);
xnor U18238 (N_18238,N_17324,N_17771);
or U18239 (N_18239,N_16994,N_17322);
nand U18240 (N_18240,N_17246,N_17434);
nor U18241 (N_18241,N_17809,N_17597);
nand U18242 (N_18242,N_17972,N_17859);
nor U18243 (N_18243,N_17961,N_17048);
or U18244 (N_18244,N_17152,N_17474);
nor U18245 (N_18245,N_17190,N_17530);
and U18246 (N_18246,N_16940,N_17722);
nand U18247 (N_18247,N_17275,N_17679);
nand U18248 (N_18248,N_17642,N_17011);
or U18249 (N_18249,N_16875,N_17174);
nor U18250 (N_18250,N_17335,N_17678);
or U18251 (N_18251,N_17987,N_17806);
nor U18252 (N_18252,N_17385,N_17383);
or U18253 (N_18253,N_17956,N_16952);
xor U18254 (N_18254,N_17382,N_16963);
and U18255 (N_18255,N_17640,N_17514);
nor U18256 (N_18256,N_17851,N_16889);
xnor U18257 (N_18257,N_17394,N_17031);
nor U18258 (N_18258,N_17102,N_17635);
nand U18259 (N_18259,N_17233,N_16985);
nand U18260 (N_18260,N_17151,N_17651);
nor U18261 (N_18261,N_16800,N_17481);
nand U18262 (N_18262,N_17745,N_17848);
nor U18263 (N_18263,N_17449,N_16859);
and U18264 (N_18264,N_17521,N_17198);
or U18265 (N_18265,N_17442,N_16971);
xnor U18266 (N_18266,N_16986,N_17975);
nand U18267 (N_18267,N_17571,N_17581);
nand U18268 (N_18268,N_17149,N_17664);
xor U18269 (N_18269,N_17386,N_17608);
xor U18270 (N_18270,N_16854,N_17127);
nand U18271 (N_18271,N_16904,N_17311);
and U18272 (N_18272,N_16924,N_17698);
xnor U18273 (N_18273,N_17634,N_17622);
or U18274 (N_18274,N_17423,N_17962);
nand U18275 (N_18275,N_17941,N_17705);
xor U18276 (N_18276,N_17470,N_17569);
nand U18277 (N_18277,N_17485,N_17493);
nor U18278 (N_18278,N_16923,N_17988);
and U18279 (N_18279,N_17658,N_17345);
xor U18280 (N_18280,N_17650,N_17269);
xor U18281 (N_18281,N_16962,N_17410);
nand U18282 (N_18282,N_17543,N_17985);
nand U18283 (N_18283,N_17464,N_17071);
nand U18284 (N_18284,N_17030,N_17797);
and U18285 (N_18285,N_17259,N_17910);
and U18286 (N_18286,N_17932,N_17256);
or U18287 (N_18287,N_17391,N_17113);
xor U18288 (N_18288,N_17496,N_17046);
nor U18289 (N_18289,N_17098,N_17253);
nand U18290 (N_18290,N_17230,N_17137);
or U18291 (N_18291,N_17236,N_17922);
or U18292 (N_18292,N_16823,N_17095);
or U18293 (N_18293,N_17494,N_17913);
nand U18294 (N_18294,N_17586,N_17487);
nand U18295 (N_18295,N_16903,N_17831);
and U18296 (N_18296,N_17959,N_17022);
nand U18297 (N_18297,N_17856,N_17703);
and U18298 (N_18298,N_17347,N_17238);
or U18299 (N_18299,N_17747,N_17645);
nor U18300 (N_18300,N_17663,N_17888);
nor U18301 (N_18301,N_17565,N_17301);
and U18302 (N_18302,N_17305,N_17087);
xor U18303 (N_18303,N_17830,N_17725);
nor U18304 (N_18304,N_17136,N_17323);
nand U18305 (N_18305,N_17536,N_16835);
xnor U18306 (N_18306,N_17116,N_17927);
or U18307 (N_18307,N_17245,N_17489);
nand U18308 (N_18308,N_17130,N_17838);
nand U18309 (N_18309,N_17654,N_17042);
xor U18310 (N_18310,N_17397,N_17900);
nand U18311 (N_18311,N_17177,N_17043);
nor U18312 (N_18312,N_17214,N_17847);
and U18313 (N_18313,N_17760,N_16836);
nor U18314 (N_18314,N_17592,N_16850);
or U18315 (N_18315,N_17192,N_17887);
and U18316 (N_18316,N_17399,N_17216);
nor U18317 (N_18317,N_16845,N_17696);
nor U18318 (N_18318,N_16951,N_17229);
or U18319 (N_18319,N_16874,N_17258);
and U18320 (N_18320,N_16936,N_17356);
xnor U18321 (N_18321,N_16894,N_17878);
xor U18322 (N_18322,N_17981,N_17316);
xor U18323 (N_18323,N_17001,N_17091);
nor U18324 (N_18324,N_16934,N_17339);
nor U18325 (N_18325,N_17176,N_17963);
xnor U18326 (N_18326,N_17605,N_17502);
or U18327 (N_18327,N_16973,N_16887);
xnor U18328 (N_18328,N_17800,N_16939);
nor U18329 (N_18329,N_17812,N_16978);
nor U18330 (N_18330,N_17307,N_17935);
nand U18331 (N_18331,N_17719,N_17873);
xor U18332 (N_18332,N_17693,N_16862);
nand U18333 (N_18333,N_17879,N_17357);
nor U18334 (N_18334,N_17550,N_17682);
or U18335 (N_18335,N_17124,N_17877);
or U18336 (N_18336,N_17829,N_17239);
nor U18337 (N_18337,N_16965,N_17947);
xnor U18338 (N_18338,N_17524,N_17479);
and U18339 (N_18339,N_17054,N_17050);
nor U18340 (N_18340,N_17477,N_17003);
or U18341 (N_18341,N_17834,N_17472);
xnor U18342 (N_18342,N_16866,N_17002);
or U18343 (N_18343,N_17753,N_17133);
or U18344 (N_18344,N_17180,N_17282);
and U18345 (N_18345,N_17789,N_17866);
nor U18346 (N_18346,N_17652,N_17096);
or U18347 (N_18347,N_17202,N_17381);
and U18348 (N_18348,N_17205,N_17478);
and U18349 (N_18349,N_17841,N_16905);
or U18350 (N_18350,N_17195,N_17457);
or U18351 (N_18351,N_17045,N_17193);
nor U18352 (N_18352,N_17052,N_17750);
and U18353 (N_18353,N_17497,N_17587);
xnor U18354 (N_18354,N_16812,N_17704);
nand U18355 (N_18355,N_17668,N_17677);
or U18356 (N_18356,N_17966,N_17780);
and U18357 (N_18357,N_17020,N_17990);
or U18358 (N_18358,N_17403,N_16821);
nand U18359 (N_18359,N_17513,N_17455);
and U18360 (N_18360,N_17062,N_17146);
or U18361 (N_18361,N_17134,N_17350);
nor U18362 (N_18362,N_16906,N_17390);
and U18363 (N_18363,N_17128,N_17531);
and U18364 (N_18364,N_16822,N_17950);
nand U18365 (N_18365,N_17231,N_17200);
or U18366 (N_18366,N_17325,N_17918);
nor U18367 (N_18367,N_17089,N_17971);
xnor U18368 (N_18368,N_16893,N_17364);
and U18369 (N_18369,N_16815,N_17649);
nor U18370 (N_18370,N_17580,N_17924);
xor U18371 (N_18371,N_17276,N_17805);
nand U18372 (N_18372,N_17810,N_17775);
or U18373 (N_18373,N_17025,N_17897);
nand U18374 (N_18374,N_16902,N_17009);
xor U18375 (N_18375,N_16947,N_17596);
or U18376 (N_18376,N_17936,N_17047);
nand U18377 (N_18377,N_17718,N_17155);
nand U18378 (N_18378,N_17590,N_17675);
and U18379 (N_18379,N_17712,N_17111);
or U18380 (N_18380,N_16801,N_17105);
and U18381 (N_18381,N_17103,N_16860);
or U18382 (N_18382,N_17730,N_17986);
and U18383 (N_18383,N_17139,N_17707);
nor U18384 (N_18384,N_17081,N_17756);
nor U18385 (N_18385,N_17097,N_16857);
and U18386 (N_18386,N_16955,N_16830);
nor U18387 (N_18387,N_17716,N_17934);
or U18388 (N_18388,N_17158,N_17845);
or U18389 (N_18389,N_17210,N_17979);
or U18390 (N_18390,N_17425,N_16915);
xnor U18391 (N_18391,N_17201,N_17359);
and U18392 (N_18392,N_17582,N_17367);
and U18393 (N_18393,N_16922,N_17049);
or U18394 (N_18394,N_17287,N_17033);
nor U18395 (N_18395,N_16839,N_17224);
nand U18396 (N_18396,N_17424,N_17053);
nor U18397 (N_18397,N_17931,N_17902);
and U18398 (N_18398,N_16950,N_17746);
xor U18399 (N_18399,N_17633,N_17393);
nor U18400 (N_18400,N_17799,N_17670);
nor U18401 (N_18401,N_17949,N_17183);
and U18402 (N_18402,N_17172,N_16929);
and U18403 (N_18403,N_17570,N_17006);
and U18404 (N_18404,N_17088,N_17890);
and U18405 (N_18405,N_17814,N_17808);
and U18406 (N_18406,N_17791,N_16858);
nor U18407 (N_18407,N_17826,N_16885);
nand U18408 (N_18408,N_16842,N_17333);
or U18409 (N_18409,N_17765,N_17637);
or U18410 (N_18410,N_17674,N_17274);
xor U18411 (N_18411,N_17370,N_17508);
nand U18412 (N_18412,N_17212,N_17764);
xnor U18413 (N_18413,N_17751,N_17398);
and U18414 (N_18414,N_17044,N_17024);
nor U18415 (N_18415,N_17108,N_17432);
nor U18416 (N_18416,N_16809,N_17065);
nand U18417 (N_18417,N_17552,N_17445);
and U18418 (N_18418,N_17860,N_17187);
and U18419 (N_18419,N_17118,N_17412);
and U18420 (N_18420,N_17291,N_17476);
xnor U18421 (N_18421,N_17646,N_16959);
nand U18422 (N_18422,N_16999,N_17620);
or U18423 (N_18423,N_17757,N_17326);
and U18424 (N_18424,N_17648,N_16944);
nor U18425 (N_18425,N_17692,N_17404);
nor U18426 (N_18426,N_17121,N_17257);
nand U18427 (N_18427,N_17551,N_17363);
nor U18428 (N_18428,N_17395,N_17666);
nor U18429 (N_18429,N_17713,N_17471);
and U18430 (N_18430,N_17084,N_16920);
xnor U18431 (N_18431,N_17562,N_17227);
or U18432 (N_18432,N_17523,N_17186);
nor U18433 (N_18433,N_17376,N_17667);
xor U18434 (N_18434,N_17203,N_17681);
nand U18435 (N_18435,N_17225,N_17321);
xnor U18436 (N_18436,N_17300,N_17014);
or U18437 (N_18437,N_17937,N_16976);
nor U18438 (N_18438,N_17568,N_16837);
xor U18439 (N_18439,N_17163,N_17784);
or U18440 (N_18440,N_16870,N_17548);
xnor U18441 (N_18441,N_17247,N_16826);
nor U18442 (N_18442,N_17318,N_17288);
or U18443 (N_18443,N_17358,N_17724);
xnor U18444 (N_18444,N_17813,N_17857);
and U18445 (N_18445,N_17749,N_17148);
or U18446 (N_18446,N_17547,N_17100);
or U18447 (N_18447,N_17285,N_16914);
and U18448 (N_18448,N_17041,N_17182);
xnor U18449 (N_18449,N_17417,N_16938);
or U18450 (N_18450,N_17453,N_17057);
or U18451 (N_18451,N_17416,N_17483);
xnor U18452 (N_18452,N_17916,N_16863);
nor U18453 (N_18453,N_17772,N_17690);
and U18454 (N_18454,N_17469,N_17880);
nor U18455 (N_18455,N_16895,N_17907);
or U18456 (N_18456,N_17327,N_16855);
xor U18457 (N_18457,N_17038,N_17617);
nor U18458 (N_18458,N_17023,N_17779);
nor U18459 (N_18459,N_17818,N_16832);
or U18460 (N_18460,N_17850,N_17209);
xor U18461 (N_18461,N_17576,N_17389);
nand U18462 (N_18462,N_16908,N_17740);
and U18463 (N_18463,N_17999,N_17761);
nand U18464 (N_18464,N_17131,N_17727);
nand U18465 (N_18465,N_17094,N_17360);
nor U18466 (N_18466,N_17539,N_17921);
nor U18467 (N_18467,N_17308,N_17181);
and U18468 (N_18468,N_16861,N_17157);
or U18469 (N_18469,N_17883,N_17304);
and U18470 (N_18470,N_17555,N_17604);
nor U18471 (N_18471,N_17315,N_16993);
nand U18472 (N_18472,N_17407,N_17785);
and U18473 (N_18473,N_17802,N_17575);
nor U18474 (N_18474,N_17021,N_16961);
xnor U18475 (N_18475,N_17135,N_17538);
and U18476 (N_18476,N_17511,N_17735);
xnor U18477 (N_18477,N_17016,N_17544);
or U18478 (N_18478,N_17317,N_16960);
and U18479 (N_18479,N_17072,N_17298);
nor U18480 (N_18480,N_17891,N_16810);
nor U18481 (N_18481,N_16865,N_17475);
nand U18482 (N_18482,N_17026,N_17170);
or U18483 (N_18483,N_17533,N_17996);
or U18484 (N_18484,N_16941,N_17559);
nor U18485 (N_18485,N_16907,N_16849);
nand U18486 (N_18486,N_17616,N_17189);
xnor U18487 (N_18487,N_17930,N_16917);
nor U18488 (N_18488,N_16975,N_17728);
xor U18489 (N_18489,N_17268,N_17939);
or U18490 (N_18490,N_17005,N_17492);
nor U18491 (N_18491,N_17843,N_17068);
nand U18492 (N_18492,N_17849,N_17661);
and U18493 (N_18493,N_17894,N_16925);
and U18494 (N_18494,N_16808,N_17289);
and U18495 (N_18495,N_16803,N_17817);
nand U18496 (N_18496,N_17970,N_17215);
or U18497 (N_18497,N_17313,N_17185);
or U18498 (N_18498,N_17519,N_17585);
nand U18499 (N_18499,N_16970,N_17123);
nand U18500 (N_18500,N_17093,N_16954);
nor U18501 (N_18501,N_17484,N_17278);
nand U18502 (N_18502,N_17083,N_17486);
xor U18503 (N_18503,N_17191,N_16992);
nand U18504 (N_18504,N_17161,N_17439);
or U18505 (N_18505,N_17655,N_17090);
or U18506 (N_18506,N_17529,N_16910);
xor U18507 (N_18507,N_16851,N_17828);
nor U18508 (N_18508,N_17498,N_17184);
and U18509 (N_18509,N_17037,N_17566);
or U18510 (N_18510,N_17839,N_17798);
and U18511 (N_18511,N_17392,N_17946);
or U18512 (N_18512,N_17167,N_17117);
xor U18513 (N_18513,N_17349,N_17614);
nor U18514 (N_18514,N_17312,N_17709);
and U18515 (N_18515,N_17702,N_17973);
xor U18516 (N_18516,N_17874,N_17297);
and U18517 (N_18517,N_17868,N_17512);
nand U18518 (N_18518,N_17428,N_17074);
nand U18519 (N_18519,N_17482,N_17018);
nor U18520 (N_18520,N_17438,N_17915);
and U18521 (N_18521,N_17542,N_17669);
xnor U18522 (N_18522,N_17467,N_17219);
or U18523 (N_18523,N_17560,N_17228);
nor U18524 (N_18524,N_17270,N_16968);
nand U18525 (N_18525,N_17631,N_17863);
nand U18526 (N_18526,N_17171,N_17528);
xor U18527 (N_18527,N_16843,N_17159);
nor U18528 (N_18528,N_17262,N_17787);
nor U18529 (N_18529,N_17241,N_17251);
and U18530 (N_18530,N_17039,N_17415);
and U18531 (N_18531,N_16829,N_17375);
nor U18532 (N_18532,N_17374,N_17532);
nor U18533 (N_18533,N_17820,N_17525);
and U18534 (N_18534,N_17885,N_17132);
nand U18535 (N_18535,N_17418,N_17341);
and U18536 (N_18536,N_17711,N_17737);
nand U18537 (N_18537,N_16883,N_17689);
nor U18538 (N_18538,N_17976,N_17504);
and U18539 (N_18539,N_17732,N_17194);
and U18540 (N_18540,N_17628,N_17168);
and U18541 (N_18541,N_17926,N_17657);
xor U18542 (N_18542,N_17060,N_17752);
and U18543 (N_18543,N_17080,N_17660);
or U18544 (N_18544,N_17147,N_17465);
or U18545 (N_18545,N_16891,N_17329);
nand U18546 (N_18546,N_16967,N_17898);
nand U18547 (N_18547,N_17871,N_17106);
and U18548 (N_18548,N_17982,N_17179);
nor U18549 (N_18549,N_17623,N_17076);
or U18550 (N_18550,N_16884,N_17440);
or U18551 (N_18551,N_17769,N_17672);
xnor U18552 (N_18552,N_17908,N_17685);
nor U18553 (N_18553,N_17207,N_17154);
nor U18554 (N_18554,N_17803,N_17366);
or U18555 (N_18555,N_17899,N_17796);
nor U18556 (N_18556,N_16897,N_17896);
nor U18557 (N_18557,N_17444,N_17697);
and U18558 (N_18558,N_17517,N_17595);
or U18559 (N_18559,N_17624,N_17688);
or U18560 (N_18560,N_17466,N_17188);
or U18561 (N_18561,N_17197,N_16802);
xnor U18562 (N_18562,N_16956,N_17362);
nand U18563 (N_18563,N_17468,N_16898);
or U18564 (N_18564,N_16935,N_17199);
or U18565 (N_18565,N_17292,N_16840);
xnor U18566 (N_18566,N_17173,N_17346);
or U18567 (N_18567,N_17903,N_17579);
nand U18568 (N_18568,N_17656,N_17881);
nor U18569 (N_18569,N_17141,N_17625);
xor U18570 (N_18570,N_17086,N_16982);
nand U18571 (N_18571,N_16980,N_17126);
nand U18572 (N_18572,N_17402,N_17680);
and U18573 (N_18573,N_17340,N_17441);
nand U18574 (N_18574,N_17244,N_17027);
and U18575 (N_18575,N_17420,N_17040);
or U18576 (N_18576,N_17731,N_17104);
or U18577 (N_18577,N_17295,N_17929);
nand U18578 (N_18578,N_17101,N_17427);
nor U18579 (N_18579,N_17928,N_17491);
or U18580 (N_18580,N_17361,N_17710);
nand U18581 (N_18581,N_16931,N_17960);
or U18582 (N_18582,N_17012,N_16880);
xnor U18583 (N_18583,N_16899,N_16828);
nor U18584 (N_18584,N_17837,N_17920);
and U18585 (N_18585,N_17178,N_17070);
xor U18586 (N_18586,N_17833,N_17232);
or U18587 (N_18587,N_17092,N_17066);
nand U18588 (N_18588,N_17801,N_17553);
and U18589 (N_18589,N_17503,N_16996);
nand U18590 (N_18590,N_16921,N_16864);
nor U18591 (N_18591,N_17380,N_17119);
xor U18592 (N_18592,N_16882,N_17036);
nor U18593 (N_18593,N_17659,N_17462);
nand U18594 (N_18594,N_17421,N_17196);
or U18595 (N_18595,N_17328,N_17795);
and U18596 (N_18596,N_16926,N_17235);
nand U18597 (N_18597,N_17912,N_17852);
or U18598 (N_18598,N_17606,N_17537);
xor U18599 (N_18599,N_17574,N_17028);
nand U18600 (N_18600,N_17847,N_17227);
and U18601 (N_18601,N_17461,N_17812);
nand U18602 (N_18602,N_17267,N_17247);
nand U18603 (N_18603,N_17402,N_17327);
or U18604 (N_18604,N_17097,N_17815);
or U18605 (N_18605,N_16982,N_17533);
nor U18606 (N_18606,N_17140,N_16978);
and U18607 (N_18607,N_16956,N_16966);
or U18608 (N_18608,N_17521,N_17558);
and U18609 (N_18609,N_17479,N_17213);
nor U18610 (N_18610,N_17514,N_17313);
or U18611 (N_18611,N_17776,N_17025);
nand U18612 (N_18612,N_17356,N_17857);
nand U18613 (N_18613,N_17926,N_16966);
nor U18614 (N_18614,N_17764,N_17506);
xor U18615 (N_18615,N_17818,N_16889);
or U18616 (N_18616,N_17852,N_17772);
nand U18617 (N_18617,N_16807,N_17262);
nand U18618 (N_18618,N_17599,N_17737);
nor U18619 (N_18619,N_17412,N_17150);
nand U18620 (N_18620,N_17934,N_17380);
xnor U18621 (N_18621,N_17424,N_17951);
nand U18622 (N_18622,N_17305,N_17118);
xor U18623 (N_18623,N_17944,N_17597);
and U18624 (N_18624,N_16932,N_17865);
nand U18625 (N_18625,N_17554,N_17228);
nand U18626 (N_18626,N_17058,N_17090);
xnor U18627 (N_18627,N_17020,N_17458);
or U18628 (N_18628,N_17597,N_16972);
nand U18629 (N_18629,N_17748,N_17103);
nand U18630 (N_18630,N_17343,N_17988);
or U18631 (N_18631,N_17253,N_17278);
and U18632 (N_18632,N_17392,N_17060);
nand U18633 (N_18633,N_16851,N_17439);
and U18634 (N_18634,N_17647,N_17255);
nand U18635 (N_18635,N_17015,N_17448);
nor U18636 (N_18636,N_17184,N_17881);
nand U18637 (N_18637,N_17250,N_17451);
nand U18638 (N_18638,N_17595,N_17578);
nor U18639 (N_18639,N_17498,N_17864);
nand U18640 (N_18640,N_17508,N_16990);
nor U18641 (N_18641,N_17352,N_17314);
or U18642 (N_18642,N_17484,N_17520);
xnor U18643 (N_18643,N_17104,N_17756);
and U18644 (N_18644,N_17979,N_17305);
nand U18645 (N_18645,N_17429,N_17090);
xor U18646 (N_18646,N_17269,N_17937);
or U18647 (N_18647,N_17385,N_17124);
nand U18648 (N_18648,N_17114,N_17869);
and U18649 (N_18649,N_17234,N_17509);
or U18650 (N_18650,N_17000,N_17879);
xor U18651 (N_18651,N_17468,N_17592);
nor U18652 (N_18652,N_16961,N_17262);
nand U18653 (N_18653,N_16989,N_17437);
nor U18654 (N_18654,N_16875,N_16843);
nor U18655 (N_18655,N_17609,N_17835);
nand U18656 (N_18656,N_17320,N_17999);
xor U18657 (N_18657,N_17995,N_17506);
nor U18658 (N_18658,N_17332,N_17776);
nand U18659 (N_18659,N_17955,N_16853);
nand U18660 (N_18660,N_17732,N_17231);
or U18661 (N_18661,N_17265,N_17031);
nand U18662 (N_18662,N_17468,N_17694);
xor U18663 (N_18663,N_17648,N_17638);
nand U18664 (N_18664,N_17106,N_17188);
xnor U18665 (N_18665,N_17386,N_17571);
xnor U18666 (N_18666,N_17832,N_17211);
nand U18667 (N_18667,N_17056,N_16857);
and U18668 (N_18668,N_17101,N_17333);
or U18669 (N_18669,N_17604,N_16838);
xnor U18670 (N_18670,N_17283,N_17641);
and U18671 (N_18671,N_17266,N_17990);
and U18672 (N_18672,N_17915,N_17543);
nor U18673 (N_18673,N_17372,N_16847);
nor U18674 (N_18674,N_16811,N_17130);
xor U18675 (N_18675,N_17894,N_17775);
nor U18676 (N_18676,N_17278,N_17678);
or U18677 (N_18677,N_17383,N_17647);
xor U18678 (N_18678,N_16894,N_17870);
nor U18679 (N_18679,N_17217,N_17493);
nor U18680 (N_18680,N_16851,N_17064);
xor U18681 (N_18681,N_16940,N_17011);
nor U18682 (N_18682,N_17756,N_17096);
nor U18683 (N_18683,N_17504,N_17498);
nor U18684 (N_18684,N_17716,N_17535);
nand U18685 (N_18685,N_17076,N_17960);
or U18686 (N_18686,N_17082,N_17380);
nor U18687 (N_18687,N_17683,N_17895);
or U18688 (N_18688,N_17691,N_17843);
or U18689 (N_18689,N_17640,N_17252);
or U18690 (N_18690,N_17943,N_17870);
nand U18691 (N_18691,N_17818,N_17684);
nand U18692 (N_18692,N_17707,N_17834);
or U18693 (N_18693,N_17180,N_17718);
xnor U18694 (N_18694,N_17667,N_17507);
or U18695 (N_18695,N_17746,N_17495);
nand U18696 (N_18696,N_17164,N_17288);
and U18697 (N_18697,N_17803,N_17676);
or U18698 (N_18698,N_17188,N_17051);
xnor U18699 (N_18699,N_17959,N_16903);
xnor U18700 (N_18700,N_17704,N_17616);
nand U18701 (N_18701,N_17364,N_17839);
nor U18702 (N_18702,N_17689,N_17778);
nand U18703 (N_18703,N_17592,N_16953);
xnor U18704 (N_18704,N_17904,N_16897);
nor U18705 (N_18705,N_17367,N_17258);
and U18706 (N_18706,N_16859,N_17900);
nor U18707 (N_18707,N_17777,N_17267);
or U18708 (N_18708,N_16959,N_17206);
and U18709 (N_18709,N_17271,N_17859);
and U18710 (N_18710,N_17185,N_17283);
and U18711 (N_18711,N_17063,N_17716);
and U18712 (N_18712,N_17911,N_17376);
or U18713 (N_18713,N_17770,N_16951);
nand U18714 (N_18714,N_17194,N_17013);
and U18715 (N_18715,N_17945,N_17785);
nor U18716 (N_18716,N_16930,N_16815);
and U18717 (N_18717,N_16891,N_17691);
nor U18718 (N_18718,N_17030,N_16995);
xnor U18719 (N_18719,N_17675,N_17849);
nor U18720 (N_18720,N_17743,N_17527);
or U18721 (N_18721,N_17048,N_17806);
nand U18722 (N_18722,N_17632,N_17429);
nand U18723 (N_18723,N_16871,N_17053);
and U18724 (N_18724,N_17366,N_17778);
and U18725 (N_18725,N_16968,N_17739);
xnor U18726 (N_18726,N_17526,N_17944);
and U18727 (N_18727,N_17720,N_17801);
nand U18728 (N_18728,N_17076,N_17714);
xor U18729 (N_18729,N_17688,N_17722);
xnor U18730 (N_18730,N_17324,N_17972);
or U18731 (N_18731,N_16868,N_17064);
nor U18732 (N_18732,N_17974,N_16978);
or U18733 (N_18733,N_17101,N_17657);
or U18734 (N_18734,N_17452,N_17114);
or U18735 (N_18735,N_17153,N_17525);
nor U18736 (N_18736,N_17532,N_17670);
nand U18737 (N_18737,N_16928,N_17442);
nand U18738 (N_18738,N_17746,N_17737);
and U18739 (N_18739,N_17086,N_17112);
or U18740 (N_18740,N_16985,N_16856);
or U18741 (N_18741,N_17866,N_17761);
nand U18742 (N_18742,N_17660,N_17180);
nand U18743 (N_18743,N_17476,N_17237);
nor U18744 (N_18744,N_17413,N_17533);
nor U18745 (N_18745,N_17383,N_17289);
or U18746 (N_18746,N_17849,N_17855);
or U18747 (N_18747,N_17343,N_17740);
nor U18748 (N_18748,N_17286,N_17851);
nor U18749 (N_18749,N_16959,N_17616);
xnor U18750 (N_18750,N_17693,N_17422);
nand U18751 (N_18751,N_17085,N_17220);
or U18752 (N_18752,N_16815,N_17850);
nor U18753 (N_18753,N_16906,N_17090);
nor U18754 (N_18754,N_17765,N_17219);
and U18755 (N_18755,N_17447,N_17283);
and U18756 (N_18756,N_17535,N_17436);
and U18757 (N_18757,N_17332,N_17188);
and U18758 (N_18758,N_17262,N_17058);
nor U18759 (N_18759,N_17184,N_17957);
or U18760 (N_18760,N_17442,N_17592);
and U18761 (N_18761,N_17745,N_17235);
or U18762 (N_18762,N_17488,N_17849);
nand U18763 (N_18763,N_17353,N_17455);
xnor U18764 (N_18764,N_17099,N_17840);
or U18765 (N_18765,N_17696,N_17328);
and U18766 (N_18766,N_17955,N_16984);
or U18767 (N_18767,N_17830,N_17738);
and U18768 (N_18768,N_17958,N_17821);
xnor U18769 (N_18769,N_17975,N_17635);
xnor U18770 (N_18770,N_17776,N_16908);
and U18771 (N_18771,N_17437,N_17971);
nand U18772 (N_18772,N_17257,N_17993);
xor U18773 (N_18773,N_17894,N_16878);
nand U18774 (N_18774,N_17249,N_16809);
nand U18775 (N_18775,N_17203,N_17862);
xnor U18776 (N_18776,N_17780,N_17127);
nor U18777 (N_18777,N_17634,N_17431);
or U18778 (N_18778,N_17488,N_17942);
nand U18779 (N_18779,N_16813,N_16858);
nor U18780 (N_18780,N_17076,N_17148);
and U18781 (N_18781,N_17587,N_17582);
nor U18782 (N_18782,N_16846,N_17119);
or U18783 (N_18783,N_17335,N_17926);
xnor U18784 (N_18784,N_17023,N_17025);
and U18785 (N_18785,N_17737,N_17121);
xnor U18786 (N_18786,N_17035,N_17321);
nor U18787 (N_18787,N_17122,N_17017);
xor U18788 (N_18788,N_17774,N_17375);
nand U18789 (N_18789,N_17997,N_17113);
and U18790 (N_18790,N_17705,N_17229);
xor U18791 (N_18791,N_16813,N_16950);
xnor U18792 (N_18792,N_17769,N_17810);
nand U18793 (N_18793,N_17268,N_17455);
nand U18794 (N_18794,N_16838,N_17764);
nand U18795 (N_18795,N_17909,N_16988);
nand U18796 (N_18796,N_16890,N_17075);
xnor U18797 (N_18797,N_17979,N_17624);
nand U18798 (N_18798,N_17129,N_17789);
or U18799 (N_18799,N_17465,N_17592);
xnor U18800 (N_18800,N_17727,N_17419);
and U18801 (N_18801,N_16843,N_17120);
xor U18802 (N_18802,N_17535,N_17226);
or U18803 (N_18803,N_16904,N_17701);
xor U18804 (N_18804,N_17009,N_17978);
xnor U18805 (N_18805,N_17058,N_17139);
and U18806 (N_18806,N_16871,N_16979);
and U18807 (N_18807,N_17113,N_17137);
and U18808 (N_18808,N_16971,N_17121);
or U18809 (N_18809,N_16950,N_17029);
nor U18810 (N_18810,N_17300,N_17113);
or U18811 (N_18811,N_17106,N_17127);
nor U18812 (N_18812,N_17095,N_17706);
xor U18813 (N_18813,N_16999,N_17271);
or U18814 (N_18814,N_17210,N_17097);
nor U18815 (N_18815,N_17359,N_16820);
nand U18816 (N_18816,N_17788,N_17325);
nor U18817 (N_18817,N_17417,N_17986);
nand U18818 (N_18818,N_16929,N_16846);
nand U18819 (N_18819,N_17878,N_17374);
xnor U18820 (N_18820,N_17487,N_17268);
xor U18821 (N_18821,N_17837,N_16835);
nor U18822 (N_18822,N_17497,N_17651);
nand U18823 (N_18823,N_16832,N_16951);
nand U18824 (N_18824,N_17051,N_17416);
and U18825 (N_18825,N_17482,N_17041);
or U18826 (N_18826,N_17298,N_17222);
nor U18827 (N_18827,N_17821,N_16836);
nor U18828 (N_18828,N_17802,N_17611);
nor U18829 (N_18829,N_17746,N_17297);
or U18830 (N_18830,N_16857,N_17836);
nor U18831 (N_18831,N_17793,N_17455);
nand U18832 (N_18832,N_16832,N_17969);
nor U18833 (N_18833,N_17413,N_17618);
or U18834 (N_18834,N_17819,N_17642);
nor U18835 (N_18835,N_17605,N_17819);
or U18836 (N_18836,N_16832,N_17427);
nand U18837 (N_18837,N_17686,N_16869);
and U18838 (N_18838,N_17550,N_17828);
xor U18839 (N_18839,N_17303,N_16854);
nand U18840 (N_18840,N_17409,N_17361);
or U18841 (N_18841,N_16802,N_16993);
and U18842 (N_18842,N_17882,N_17078);
and U18843 (N_18843,N_17129,N_17965);
nand U18844 (N_18844,N_17848,N_17115);
nand U18845 (N_18845,N_17523,N_17000);
or U18846 (N_18846,N_16978,N_17951);
nand U18847 (N_18847,N_16974,N_17383);
or U18848 (N_18848,N_16861,N_17459);
xor U18849 (N_18849,N_17226,N_17231);
xor U18850 (N_18850,N_17235,N_17779);
nand U18851 (N_18851,N_16853,N_17721);
or U18852 (N_18852,N_17932,N_16982);
nand U18853 (N_18853,N_17135,N_17978);
xnor U18854 (N_18854,N_16988,N_17451);
nor U18855 (N_18855,N_17011,N_17610);
nand U18856 (N_18856,N_17409,N_17578);
nor U18857 (N_18857,N_17223,N_17264);
nor U18858 (N_18858,N_17654,N_17635);
and U18859 (N_18859,N_16805,N_17522);
nand U18860 (N_18860,N_17817,N_17921);
and U18861 (N_18861,N_17772,N_16954);
and U18862 (N_18862,N_17346,N_17272);
and U18863 (N_18863,N_17859,N_17973);
xnor U18864 (N_18864,N_17213,N_17791);
nand U18865 (N_18865,N_16833,N_16835);
xnor U18866 (N_18866,N_17781,N_17598);
nand U18867 (N_18867,N_17134,N_16818);
or U18868 (N_18868,N_16920,N_17508);
nand U18869 (N_18869,N_17275,N_16977);
nand U18870 (N_18870,N_17545,N_17464);
nand U18871 (N_18871,N_17109,N_17534);
nor U18872 (N_18872,N_17383,N_16859);
or U18873 (N_18873,N_17312,N_17593);
nand U18874 (N_18874,N_17929,N_17160);
nand U18875 (N_18875,N_17134,N_16896);
or U18876 (N_18876,N_16845,N_17903);
or U18877 (N_18877,N_17550,N_17796);
and U18878 (N_18878,N_17509,N_16824);
or U18879 (N_18879,N_17918,N_17393);
nand U18880 (N_18880,N_17205,N_16880);
xor U18881 (N_18881,N_17832,N_17169);
xnor U18882 (N_18882,N_17412,N_17091);
and U18883 (N_18883,N_16875,N_16824);
xor U18884 (N_18884,N_17975,N_17421);
nand U18885 (N_18885,N_16848,N_17372);
xor U18886 (N_18886,N_17362,N_17822);
nand U18887 (N_18887,N_17538,N_16920);
xnor U18888 (N_18888,N_17740,N_17030);
nand U18889 (N_18889,N_16940,N_16804);
nand U18890 (N_18890,N_17675,N_17098);
and U18891 (N_18891,N_17944,N_16979);
or U18892 (N_18892,N_17881,N_17875);
xnor U18893 (N_18893,N_17959,N_17752);
and U18894 (N_18894,N_17171,N_17033);
nand U18895 (N_18895,N_17459,N_17411);
nor U18896 (N_18896,N_17602,N_17304);
nor U18897 (N_18897,N_16957,N_17834);
nand U18898 (N_18898,N_17393,N_17545);
nor U18899 (N_18899,N_17720,N_17930);
nor U18900 (N_18900,N_17588,N_17725);
nand U18901 (N_18901,N_17486,N_17785);
and U18902 (N_18902,N_17687,N_17582);
or U18903 (N_18903,N_17851,N_17103);
xnor U18904 (N_18904,N_17713,N_17321);
nand U18905 (N_18905,N_17957,N_16982);
or U18906 (N_18906,N_17072,N_17138);
or U18907 (N_18907,N_16868,N_17950);
or U18908 (N_18908,N_17868,N_17978);
nand U18909 (N_18909,N_17607,N_17086);
or U18910 (N_18910,N_17913,N_16865);
nor U18911 (N_18911,N_17318,N_17195);
nor U18912 (N_18912,N_17800,N_17146);
nor U18913 (N_18913,N_17544,N_17808);
or U18914 (N_18914,N_17541,N_17516);
or U18915 (N_18915,N_17116,N_17846);
nor U18916 (N_18916,N_17112,N_17825);
xor U18917 (N_18917,N_17718,N_17372);
or U18918 (N_18918,N_16986,N_17913);
nor U18919 (N_18919,N_17220,N_17831);
nand U18920 (N_18920,N_17499,N_17068);
xnor U18921 (N_18921,N_17768,N_17626);
xnor U18922 (N_18922,N_17372,N_17408);
nor U18923 (N_18923,N_17116,N_17382);
nor U18924 (N_18924,N_17281,N_17909);
nand U18925 (N_18925,N_17672,N_17345);
or U18926 (N_18926,N_17442,N_17260);
nor U18927 (N_18927,N_17962,N_17770);
xnor U18928 (N_18928,N_17525,N_17566);
nand U18929 (N_18929,N_17590,N_17880);
and U18930 (N_18930,N_16967,N_17376);
nor U18931 (N_18931,N_17388,N_17027);
or U18932 (N_18932,N_17432,N_17385);
nor U18933 (N_18933,N_17243,N_17897);
nand U18934 (N_18934,N_17897,N_17015);
or U18935 (N_18935,N_17005,N_17310);
or U18936 (N_18936,N_17443,N_17074);
nand U18937 (N_18937,N_17531,N_16943);
xnor U18938 (N_18938,N_17945,N_17093);
and U18939 (N_18939,N_17381,N_17847);
nand U18940 (N_18940,N_17852,N_17983);
or U18941 (N_18941,N_16836,N_17914);
or U18942 (N_18942,N_17703,N_17392);
nor U18943 (N_18943,N_16848,N_16999);
xnor U18944 (N_18944,N_17789,N_17820);
or U18945 (N_18945,N_17102,N_17611);
and U18946 (N_18946,N_17452,N_17823);
nor U18947 (N_18947,N_17382,N_17441);
nand U18948 (N_18948,N_17800,N_17284);
nand U18949 (N_18949,N_17463,N_17529);
or U18950 (N_18950,N_17610,N_16959);
nand U18951 (N_18951,N_17707,N_17425);
or U18952 (N_18952,N_17068,N_17577);
xor U18953 (N_18953,N_17493,N_17356);
and U18954 (N_18954,N_17763,N_17461);
nor U18955 (N_18955,N_17513,N_17408);
and U18956 (N_18956,N_17579,N_16970);
nand U18957 (N_18957,N_16862,N_17505);
and U18958 (N_18958,N_17278,N_17651);
or U18959 (N_18959,N_17002,N_16910);
nor U18960 (N_18960,N_17282,N_17608);
nand U18961 (N_18961,N_17470,N_16898);
nor U18962 (N_18962,N_16932,N_17374);
nand U18963 (N_18963,N_17364,N_16849);
xnor U18964 (N_18964,N_17356,N_17422);
nand U18965 (N_18965,N_17136,N_17436);
or U18966 (N_18966,N_17604,N_17803);
xnor U18967 (N_18967,N_17177,N_17668);
nor U18968 (N_18968,N_17191,N_17259);
and U18969 (N_18969,N_17824,N_17648);
and U18970 (N_18970,N_17046,N_17472);
nand U18971 (N_18971,N_17775,N_17054);
and U18972 (N_18972,N_17002,N_17564);
xor U18973 (N_18973,N_17334,N_17526);
nand U18974 (N_18974,N_17753,N_17338);
or U18975 (N_18975,N_17285,N_17698);
nand U18976 (N_18976,N_16999,N_16896);
nor U18977 (N_18977,N_17096,N_17635);
xnor U18978 (N_18978,N_17549,N_17767);
xor U18979 (N_18979,N_17910,N_17737);
and U18980 (N_18980,N_17359,N_17335);
xnor U18981 (N_18981,N_17330,N_17879);
and U18982 (N_18982,N_17795,N_17132);
nand U18983 (N_18983,N_16930,N_16835);
and U18984 (N_18984,N_17225,N_17880);
or U18985 (N_18985,N_17489,N_17133);
or U18986 (N_18986,N_17835,N_17826);
nor U18987 (N_18987,N_17527,N_17099);
or U18988 (N_18988,N_17283,N_17195);
and U18989 (N_18989,N_17836,N_17965);
and U18990 (N_18990,N_17049,N_16852);
or U18991 (N_18991,N_17767,N_17633);
or U18992 (N_18992,N_17343,N_16863);
nor U18993 (N_18993,N_16948,N_17876);
nor U18994 (N_18994,N_17869,N_17889);
xor U18995 (N_18995,N_17994,N_17463);
or U18996 (N_18996,N_17963,N_17454);
nor U18997 (N_18997,N_16980,N_17985);
or U18998 (N_18998,N_17013,N_17736);
and U18999 (N_18999,N_17891,N_17075);
nand U19000 (N_19000,N_17425,N_17445);
nor U19001 (N_19001,N_17530,N_17984);
or U19002 (N_19002,N_17813,N_16817);
and U19003 (N_19003,N_16964,N_17777);
or U19004 (N_19004,N_17465,N_17662);
and U19005 (N_19005,N_17328,N_17069);
nor U19006 (N_19006,N_17801,N_17852);
and U19007 (N_19007,N_17065,N_17536);
nor U19008 (N_19008,N_17484,N_17047);
xor U19009 (N_19009,N_17817,N_17471);
and U19010 (N_19010,N_17071,N_17621);
and U19011 (N_19011,N_17829,N_17613);
and U19012 (N_19012,N_16803,N_17355);
nand U19013 (N_19013,N_16827,N_17779);
nor U19014 (N_19014,N_16862,N_17292);
nand U19015 (N_19015,N_17850,N_17483);
xnor U19016 (N_19016,N_17955,N_16880);
nand U19017 (N_19017,N_17232,N_17415);
nor U19018 (N_19018,N_17845,N_17805);
or U19019 (N_19019,N_17946,N_17224);
nor U19020 (N_19020,N_17547,N_16982);
xor U19021 (N_19021,N_17696,N_17117);
and U19022 (N_19022,N_16932,N_17787);
and U19023 (N_19023,N_17838,N_17986);
or U19024 (N_19024,N_17169,N_17540);
nor U19025 (N_19025,N_17314,N_17020);
xnor U19026 (N_19026,N_17783,N_17650);
nor U19027 (N_19027,N_17110,N_17080);
and U19028 (N_19028,N_17044,N_17966);
nand U19029 (N_19029,N_17072,N_17524);
and U19030 (N_19030,N_17817,N_17805);
nand U19031 (N_19031,N_16812,N_17234);
or U19032 (N_19032,N_17581,N_17232);
and U19033 (N_19033,N_17109,N_17766);
xnor U19034 (N_19034,N_17666,N_17331);
nor U19035 (N_19035,N_17947,N_17687);
and U19036 (N_19036,N_17230,N_17127);
nor U19037 (N_19037,N_17942,N_16803);
nor U19038 (N_19038,N_17809,N_17290);
and U19039 (N_19039,N_17053,N_17205);
nand U19040 (N_19040,N_17177,N_17126);
nand U19041 (N_19041,N_17356,N_17932);
nand U19042 (N_19042,N_17778,N_16916);
nand U19043 (N_19043,N_17052,N_17982);
or U19044 (N_19044,N_17594,N_16838);
and U19045 (N_19045,N_17234,N_17702);
xnor U19046 (N_19046,N_16811,N_17845);
nor U19047 (N_19047,N_16986,N_17712);
and U19048 (N_19048,N_17589,N_17165);
nor U19049 (N_19049,N_17852,N_17358);
or U19050 (N_19050,N_17904,N_17444);
or U19051 (N_19051,N_17265,N_17084);
nor U19052 (N_19052,N_17814,N_17117);
nor U19053 (N_19053,N_17779,N_17875);
nor U19054 (N_19054,N_17017,N_17614);
nor U19055 (N_19055,N_17647,N_17091);
nand U19056 (N_19056,N_17082,N_17915);
and U19057 (N_19057,N_17017,N_17699);
nand U19058 (N_19058,N_17791,N_17772);
nor U19059 (N_19059,N_17736,N_17780);
nor U19060 (N_19060,N_17917,N_17280);
or U19061 (N_19061,N_17252,N_16989);
nand U19062 (N_19062,N_17099,N_17540);
nand U19063 (N_19063,N_17503,N_17741);
nand U19064 (N_19064,N_17721,N_17381);
nor U19065 (N_19065,N_17376,N_17292);
xor U19066 (N_19066,N_17063,N_16819);
or U19067 (N_19067,N_17878,N_17364);
and U19068 (N_19068,N_17392,N_17307);
or U19069 (N_19069,N_17622,N_17830);
nand U19070 (N_19070,N_17920,N_17157);
or U19071 (N_19071,N_17809,N_17569);
or U19072 (N_19072,N_17820,N_17411);
and U19073 (N_19073,N_17507,N_17472);
and U19074 (N_19074,N_17433,N_16823);
and U19075 (N_19075,N_16861,N_17527);
or U19076 (N_19076,N_17608,N_17982);
xnor U19077 (N_19077,N_17566,N_17110);
nand U19078 (N_19078,N_17960,N_17743);
or U19079 (N_19079,N_17757,N_16903);
and U19080 (N_19080,N_16822,N_17266);
xnor U19081 (N_19081,N_17815,N_17693);
and U19082 (N_19082,N_17566,N_17426);
nor U19083 (N_19083,N_16862,N_17614);
or U19084 (N_19084,N_17859,N_17251);
and U19085 (N_19085,N_17214,N_17058);
or U19086 (N_19086,N_17474,N_17688);
nand U19087 (N_19087,N_16927,N_16981);
and U19088 (N_19088,N_17122,N_16850);
nand U19089 (N_19089,N_17056,N_17405);
nand U19090 (N_19090,N_17188,N_17517);
nor U19091 (N_19091,N_17782,N_17424);
xor U19092 (N_19092,N_17046,N_16979);
or U19093 (N_19093,N_17697,N_17386);
nor U19094 (N_19094,N_17272,N_17698);
or U19095 (N_19095,N_17759,N_17854);
or U19096 (N_19096,N_16937,N_17726);
nand U19097 (N_19097,N_17674,N_17445);
and U19098 (N_19098,N_17040,N_17098);
nand U19099 (N_19099,N_17910,N_17649);
nand U19100 (N_19100,N_17606,N_17271);
xor U19101 (N_19101,N_17415,N_17157);
nand U19102 (N_19102,N_17834,N_17787);
nor U19103 (N_19103,N_17374,N_17678);
and U19104 (N_19104,N_17177,N_17689);
nor U19105 (N_19105,N_17785,N_17755);
nand U19106 (N_19106,N_17282,N_17756);
or U19107 (N_19107,N_16803,N_17900);
or U19108 (N_19108,N_17439,N_16827);
and U19109 (N_19109,N_17943,N_17836);
nand U19110 (N_19110,N_17009,N_17876);
and U19111 (N_19111,N_17763,N_17291);
or U19112 (N_19112,N_16818,N_17775);
or U19113 (N_19113,N_17742,N_17693);
nand U19114 (N_19114,N_17843,N_17257);
or U19115 (N_19115,N_17978,N_16971);
nand U19116 (N_19116,N_17383,N_17258);
xor U19117 (N_19117,N_17216,N_17207);
and U19118 (N_19118,N_17203,N_17906);
nor U19119 (N_19119,N_17187,N_17466);
xor U19120 (N_19120,N_17422,N_17583);
or U19121 (N_19121,N_17467,N_17367);
xor U19122 (N_19122,N_17718,N_17528);
xnor U19123 (N_19123,N_17090,N_17226);
nor U19124 (N_19124,N_17659,N_17688);
and U19125 (N_19125,N_17916,N_17607);
nor U19126 (N_19126,N_16812,N_17458);
and U19127 (N_19127,N_16807,N_17201);
nor U19128 (N_19128,N_17378,N_17526);
xnor U19129 (N_19129,N_17682,N_17070);
nand U19130 (N_19130,N_17162,N_17674);
and U19131 (N_19131,N_16952,N_17621);
and U19132 (N_19132,N_16926,N_17273);
and U19133 (N_19133,N_17600,N_16957);
nand U19134 (N_19134,N_16930,N_17562);
and U19135 (N_19135,N_17291,N_17439);
and U19136 (N_19136,N_17563,N_17080);
or U19137 (N_19137,N_17001,N_17159);
and U19138 (N_19138,N_17772,N_17479);
or U19139 (N_19139,N_17022,N_16980);
nand U19140 (N_19140,N_17572,N_17620);
nand U19141 (N_19141,N_17406,N_17146);
or U19142 (N_19142,N_16828,N_17147);
xor U19143 (N_19143,N_17493,N_17398);
and U19144 (N_19144,N_17528,N_17204);
nor U19145 (N_19145,N_17614,N_17853);
xnor U19146 (N_19146,N_17059,N_16967);
xnor U19147 (N_19147,N_17227,N_17825);
nor U19148 (N_19148,N_17234,N_17466);
nor U19149 (N_19149,N_17072,N_17698);
xnor U19150 (N_19150,N_17278,N_17898);
xnor U19151 (N_19151,N_17016,N_17934);
or U19152 (N_19152,N_17079,N_17918);
and U19153 (N_19153,N_17506,N_17710);
nor U19154 (N_19154,N_16853,N_17343);
or U19155 (N_19155,N_17915,N_17857);
nand U19156 (N_19156,N_16882,N_17763);
xor U19157 (N_19157,N_17872,N_17430);
xnor U19158 (N_19158,N_17705,N_17486);
and U19159 (N_19159,N_17748,N_17425);
xnor U19160 (N_19160,N_17647,N_17199);
nand U19161 (N_19161,N_17229,N_16882);
xor U19162 (N_19162,N_17369,N_16964);
nand U19163 (N_19163,N_16867,N_17429);
nand U19164 (N_19164,N_17855,N_17600);
and U19165 (N_19165,N_17690,N_17217);
xnor U19166 (N_19166,N_17816,N_17831);
nor U19167 (N_19167,N_17943,N_17046);
or U19168 (N_19168,N_17118,N_17403);
nand U19169 (N_19169,N_16814,N_17647);
or U19170 (N_19170,N_17859,N_17982);
nand U19171 (N_19171,N_17050,N_16983);
xnor U19172 (N_19172,N_17868,N_17838);
and U19173 (N_19173,N_17416,N_17937);
nand U19174 (N_19174,N_16864,N_17765);
and U19175 (N_19175,N_17301,N_17905);
xor U19176 (N_19176,N_17549,N_17159);
xnor U19177 (N_19177,N_17851,N_17684);
or U19178 (N_19178,N_17554,N_17733);
xnor U19179 (N_19179,N_16956,N_17228);
xor U19180 (N_19180,N_17824,N_17674);
xnor U19181 (N_19181,N_17422,N_17947);
nor U19182 (N_19182,N_17005,N_17806);
nand U19183 (N_19183,N_17168,N_17494);
xnor U19184 (N_19184,N_17545,N_17445);
nor U19185 (N_19185,N_17510,N_17872);
or U19186 (N_19186,N_17841,N_17528);
nor U19187 (N_19187,N_17327,N_17976);
and U19188 (N_19188,N_17574,N_17479);
or U19189 (N_19189,N_17797,N_17301);
xnor U19190 (N_19190,N_17303,N_17940);
or U19191 (N_19191,N_17703,N_17276);
nand U19192 (N_19192,N_17395,N_17449);
nand U19193 (N_19193,N_17876,N_17077);
or U19194 (N_19194,N_16921,N_17617);
or U19195 (N_19195,N_17413,N_17934);
nand U19196 (N_19196,N_17802,N_16833);
xnor U19197 (N_19197,N_16875,N_17427);
or U19198 (N_19198,N_16957,N_16803);
or U19199 (N_19199,N_17499,N_17450);
or U19200 (N_19200,N_18451,N_18628);
or U19201 (N_19201,N_18692,N_18087);
or U19202 (N_19202,N_18686,N_19140);
xor U19203 (N_19203,N_18066,N_19011);
or U19204 (N_19204,N_18007,N_18926);
nand U19205 (N_19205,N_18356,N_18953);
xor U19206 (N_19206,N_18924,N_18191);
and U19207 (N_19207,N_18691,N_18154);
nand U19208 (N_19208,N_18837,N_18798);
xnor U19209 (N_19209,N_18971,N_18580);
and U19210 (N_19210,N_19006,N_19136);
or U19211 (N_19211,N_18123,N_18872);
nor U19212 (N_19212,N_18062,N_19150);
xnor U19213 (N_19213,N_18721,N_18519);
and U19214 (N_19214,N_18940,N_18917);
nand U19215 (N_19215,N_18586,N_18326);
or U19216 (N_19216,N_18044,N_18311);
and U19217 (N_19217,N_18243,N_18282);
or U19218 (N_19218,N_18323,N_18011);
nand U19219 (N_19219,N_18800,N_18269);
or U19220 (N_19220,N_18575,N_18220);
nand U19221 (N_19221,N_18083,N_18690);
nand U19222 (N_19222,N_18002,N_18255);
or U19223 (N_19223,N_18277,N_18228);
or U19224 (N_19224,N_18383,N_18640);
or U19225 (N_19225,N_18367,N_18652);
nand U19226 (N_19226,N_18649,N_18179);
nor U19227 (N_19227,N_18873,N_18127);
xnor U19228 (N_19228,N_19049,N_18241);
nand U19229 (N_19229,N_18295,N_19198);
xnor U19230 (N_19230,N_18620,N_18854);
or U19231 (N_19231,N_18942,N_18380);
nand U19232 (N_19232,N_18831,N_19099);
nand U19233 (N_19233,N_19118,N_19183);
and U19234 (N_19234,N_18515,N_18650);
nor U19235 (N_19235,N_18256,N_18545);
nand U19236 (N_19236,N_18101,N_18895);
or U19237 (N_19237,N_18463,N_18314);
and U19238 (N_19238,N_18198,N_18107);
and U19239 (N_19239,N_18009,N_18625);
nand U19240 (N_19240,N_18750,N_18542);
xor U19241 (N_19241,N_18883,N_18422);
xnor U19242 (N_19242,N_18700,N_18151);
xnor U19243 (N_19243,N_18597,N_18526);
and U19244 (N_19244,N_18371,N_18125);
nor U19245 (N_19245,N_18997,N_18109);
nand U19246 (N_19246,N_18962,N_18038);
nand U19247 (N_19247,N_18240,N_18784);
xnor U19248 (N_19248,N_18075,N_18478);
and U19249 (N_19249,N_19074,N_18560);
xor U19250 (N_19250,N_18772,N_18785);
nand U19251 (N_19251,N_18466,N_19031);
nand U19252 (N_19252,N_18826,N_18175);
xnor U19253 (N_19253,N_18681,N_18850);
xor U19254 (N_19254,N_19126,N_18008);
or U19255 (N_19255,N_18822,N_18386);
and U19256 (N_19256,N_18814,N_18782);
nand U19257 (N_19257,N_18443,N_18554);
and U19258 (N_19258,N_18131,N_18032);
nand U19259 (N_19259,N_19025,N_18048);
or U19260 (N_19260,N_18280,N_19055);
and U19261 (N_19261,N_18186,N_18161);
nand U19262 (N_19262,N_19192,N_19163);
or U19263 (N_19263,N_18321,N_18874);
or U19264 (N_19264,N_18737,N_18056);
nor U19265 (N_19265,N_18727,N_18844);
nor U19266 (N_19266,N_19159,N_18433);
nor U19267 (N_19267,N_18794,N_18548);
and U19268 (N_19268,N_18345,N_18003);
nand U19269 (N_19269,N_18055,N_18041);
nand U19270 (N_19270,N_18956,N_18808);
and U19271 (N_19271,N_18384,N_18049);
nor U19272 (N_19272,N_18335,N_19182);
and U19273 (N_19273,N_18912,N_18669);
or U19274 (N_19274,N_19103,N_18194);
nand U19275 (N_19275,N_18106,N_19082);
nor U19276 (N_19276,N_19147,N_19190);
nand U19277 (N_19277,N_18936,N_18818);
and U19278 (N_19278,N_18638,N_19153);
nor U19279 (N_19279,N_18306,N_18405);
nand U19280 (N_19280,N_18500,N_18347);
nand U19281 (N_19281,N_18033,N_18039);
nand U19282 (N_19282,N_18922,N_18525);
xnor U19283 (N_19283,N_19177,N_19085);
nand U19284 (N_19284,N_18090,N_18014);
or U19285 (N_19285,N_18735,N_18996);
nor U19286 (N_19286,N_18570,N_18390);
nand U19287 (N_19287,N_18215,N_18973);
nand U19288 (N_19288,N_18627,N_18265);
and U19289 (N_19289,N_18694,N_18455);
nor U19290 (N_19290,N_18828,N_18904);
nand U19291 (N_19291,N_18675,N_18070);
and U19292 (N_19292,N_18459,N_19073);
nand U19293 (N_19293,N_19127,N_18394);
xor U19294 (N_19294,N_18855,N_18745);
and U19295 (N_19295,N_18930,N_19187);
or U19296 (N_19296,N_18111,N_18078);
or U19297 (N_19297,N_19157,N_18832);
or U19298 (N_19298,N_18689,N_18980);
xnor U19299 (N_19299,N_18188,N_18751);
nor U19300 (N_19300,N_18209,N_18104);
nand U19301 (N_19301,N_18724,N_18567);
xor U19302 (N_19302,N_19078,N_18102);
or U19303 (N_19303,N_18440,N_18299);
nor U19304 (N_19304,N_18085,N_18250);
and U19305 (N_19305,N_18779,N_18130);
nor U19306 (N_19306,N_18132,N_18103);
nor U19307 (N_19307,N_19068,N_18609);
and U19308 (N_19308,N_18637,N_18608);
xor U19309 (N_19309,N_18088,N_18457);
and U19310 (N_19310,N_18774,N_18170);
and U19311 (N_19311,N_18113,N_18998);
nand U19312 (N_19312,N_19046,N_18482);
nor U19313 (N_19313,N_18664,N_18589);
nor U19314 (N_19314,N_18114,N_18404);
nor U19315 (N_19315,N_18835,N_19165);
xnor U19316 (N_19316,N_18484,N_18067);
and U19317 (N_19317,N_19086,N_18678);
and U19318 (N_19318,N_18730,N_18807);
xnor U19319 (N_19319,N_18577,N_18937);
nor U19320 (N_19320,N_18984,N_18925);
nor U19321 (N_19321,N_18171,N_19023);
xor U19322 (N_19322,N_18355,N_18246);
nand U19323 (N_19323,N_18605,N_18660);
and U19324 (N_19324,N_18290,N_18398);
nand U19325 (N_19325,N_19133,N_18441);
nor U19326 (N_19326,N_18214,N_18324);
nor U19327 (N_19327,N_18712,N_18871);
nor U19328 (N_19328,N_18334,N_19195);
xor U19329 (N_19329,N_19032,N_18665);
nor U19330 (N_19330,N_18923,N_18911);
nand U19331 (N_19331,N_18251,N_18167);
nand U19332 (N_19332,N_18746,N_19186);
xor U19333 (N_19333,N_18770,N_18516);
or U19334 (N_19334,N_18225,N_18933);
xor U19335 (N_19335,N_19035,N_18229);
and U19336 (N_19336,N_18447,N_18363);
and U19337 (N_19337,N_18733,N_18034);
and U19338 (N_19338,N_18181,N_19178);
and U19339 (N_19339,N_18732,N_18285);
nor U19340 (N_19340,N_19056,N_18739);
nor U19341 (N_19341,N_18564,N_18415);
nand U19342 (N_19342,N_18322,N_18557);
nand U19343 (N_19343,N_18659,N_18763);
or U19344 (N_19344,N_18811,N_18474);
nor U19345 (N_19345,N_18117,N_18619);
and U19346 (N_19346,N_18706,N_18645);
nor U19347 (N_19347,N_18533,N_18616);
nor U19348 (N_19348,N_18201,N_19061);
nor U19349 (N_19349,N_18312,N_18445);
nand U19350 (N_19350,N_18037,N_18025);
nand U19351 (N_19351,N_18110,N_18431);
or U19352 (N_19352,N_18452,N_18756);
nor U19353 (N_19353,N_18614,N_19128);
xor U19354 (N_19354,N_18054,N_18591);
nand U19355 (N_19355,N_18339,N_18695);
nand U19356 (N_19356,N_18530,N_18001);
xor U19357 (N_19357,N_18498,N_19119);
xor U19358 (N_19358,N_18658,N_18421);
and U19359 (N_19359,N_18200,N_19123);
nand U19360 (N_19360,N_18095,N_19114);
nand U19361 (N_19361,N_18680,N_18511);
nor U19362 (N_19362,N_18699,N_18333);
nand U19363 (N_19363,N_18332,N_19041);
or U19364 (N_19364,N_18419,N_18899);
and U19365 (N_19365,N_19048,N_18468);
nand U19366 (N_19366,N_18975,N_19088);
or U19367 (N_19367,N_18726,N_18178);
nand U19368 (N_19368,N_18100,N_19110);
and U19369 (N_19369,N_18242,N_18787);
xnor U19370 (N_19370,N_19017,N_18298);
xor U19371 (N_19371,N_19194,N_19059);
nor U19372 (N_19372,N_18990,N_18847);
nor U19373 (N_19373,N_18051,N_18366);
nand U19374 (N_19374,N_18610,N_18909);
or U19375 (N_19375,N_18187,N_18592);
nor U19376 (N_19376,N_18288,N_19174);
nor U19377 (N_19377,N_18042,N_18802);
nor U19378 (N_19378,N_18920,N_18579);
nor U19379 (N_19379,N_18865,N_18071);
or U19380 (N_19380,N_18999,N_18584);
nor U19381 (N_19381,N_18825,N_19009);
or U19382 (N_19382,N_18226,N_18778);
or U19383 (N_19383,N_19001,N_18024);
nand U19384 (N_19384,N_18230,N_18857);
xor U19385 (N_19385,N_18632,N_18408);
nand U19386 (N_19386,N_18365,N_18454);
nor U19387 (N_19387,N_18183,N_18821);
and U19388 (N_19388,N_18891,N_18718);
and U19389 (N_19389,N_18771,N_18646);
and U19390 (N_19390,N_18738,N_18657);
nand U19391 (N_19391,N_19018,N_18611);
and U19392 (N_19392,N_18860,N_18065);
and U19393 (N_19393,N_19148,N_18830);
and U19394 (N_19394,N_18862,N_18544);
nor U19395 (N_19395,N_18613,N_18257);
xor U19396 (N_19396,N_18254,N_18728);
xor U19397 (N_19397,N_18340,N_19138);
or U19398 (N_19398,N_19132,N_18052);
nand U19399 (N_19399,N_18907,N_18966);
nand U19400 (N_19400,N_19037,N_19051);
or U19401 (N_19401,N_18098,N_18057);
and U19402 (N_19402,N_18674,N_18166);
nand U19403 (N_19403,N_18710,N_18320);
xor U19404 (N_19404,N_18086,N_18489);
or U19405 (N_19405,N_18900,N_18399);
and U19406 (N_19406,N_18602,N_18969);
nand U19407 (N_19407,N_18853,N_18302);
and U19408 (N_19408,N_19151,N_18473);
xnor U19409 (N_19409,N_18174,N_18769);
xnor U19410 (N_19410,N_18867,N_18708);
or U19411 (N_19411,N_18604,N_18654);
or U19412 (N_19412,N_18858,N_18908);
nor U19413 (N_19413,N_18145,N_18029);
nor U19414 (N_19414,N_18734,N_18842);
or U19415 (N_19415,N_18353,N_18972);
nor U19416 (N_19416,N_18805,N_18801);
or U19417 (N_19417,N_18546,N_18758);
or U19418 (N_19418,N_18283,N_18262);
nor U19419 (N_19419,N_18995,N_18676);
nor U19420 (N_19420,N_19131,N_18133);
nor U19421 (N_19421,N_19158,N_19058);
xnor U19422 (N_19422,N_18709,N_18134);
or U19423 (N_19423,N_19089,N_18931);
or U19424 (N_19424,N_18521,N_18069);
and U19425 (N_19425,N_18596,N_18081);
nor U19426 (N_19426,N_18509,N_18437);
nor U19427 (N_19427,N_18305,N_18409);
or U19428 (N_19428,N_18742,N_18144);
nor U19429 (N_19429,N_19175,N_18590);
or U19430 (N_19430,N_18679,N_18747);
nand U19431 (N_19431,N_18612,N_18812);
or U19432 (N_19432,N_18744,N_18607);
xnor U19433 (N_19433,N_18434,N_18713);
or U19434 (N_19434,N_19117,N_19092);
xnor U19435 (N_19435,N_18291,N_18767);
xor U19436 (N_19436,N_18958,N_18886);
nor U19437 (N_19437,N_18651,N_18252);
or U19438 (N_19438,N_18279,N_18562);
or U19439 (N_19439,N_18276,N_18006);
nand U19440 (N_19440,N_18878,N_18470);
or U19441 (N_19441,N_19162,N_19002);
and U19442 (N_19442,N_18983,N_18328);
nor U19443 (N_19443,N_18236,N_18947);
and U19444 (N_19444,N_18359,N_18278);
or U19445 (N_19445,N_19076,N_18094);
xor U19446 (N_19446,N_19067,N_18864);
nor U19447 (N_19447,N_18158,N_18879);
nand U19448 (N_19448,N_18082,N_18688);
xor U19449 (N_19449,N_18450,N_18776);
nand U19450 (N_19450,N_18076,N_18631);
or U19451 (N_19451,N_18268,N_18720);
or U19452 (N_19452,N_18722,N_18513);
nor U19453 (N_19453,N_18939,N_19063);
and U19454 (N_19454,N_18211,N_18817);
nand U19455 (N_19455,N_18424,N_19169);
xor U19456 (N_19456,N_18547,N_18403);
xor U19457 (N_19457,N_18216,N_18361);
nor U19458 (N_19458,N_18633,N_18479);
nand U19459 (N_19459,N_18137,N_18881);
xor U19460 (N_19460,N_19122,N_18869);
nor U19461 (N_19461,N_19028,N_18696);
nor U19462 (N_19462,N_18022,N_18795);
nor U19463 (N_19463,N_18430,N_18296);
and U19464 (N_19464,N_18261,N_18019);
and U19465 (N_19465,N_18838,N_18761);
xor U19466 (N_19466,N_18868,N_18495);
or U19467 (N_19467,N_18558,N_18385);
nor U19468 (N_19468,N_19197,N_18193);
xnor U19469 (N_19469,N_19042,N_18264);
or U19470 (N_19470,N_18266,N_18494);
or U19471 (N_19471,N_19021,N_18496);
and U19472 (N_19472,N_18205,N_18781);
nor U19473 (N_19473,N_18587,N_18938);
xnor U19474 (N_19474,N_19171,N_18374);
and U19475 (N_19475,N_18396,N_18987);
and U19476 (N_19476,N_18594,N_18413);
and U19477 (N_19477,N_19013,N_18816);
or U19478 (N_19478,N_18461,N_18824);
and U19479 (N_19479,N_18458,N_18898);
or U19480 (N_19480,N_18989,N_18372);
nand U19481 (N_19481,N_19047,N_18128);
and U19482 (N_19482,N_18543,N_18848);
xor U19483 (N_19483,N_18523,N_18316);
nor U19484 (N_19484,N_18307,N_18199);
nor U19485 (N_19485,N_18275,N_18227);
nand U19486 (N_19486,N_19105,N_18017);
nand U19487 (N_19487,N_18503,N_19125);
nor U19488 (N_19488,N_19145,N_18204);
xnor U19489 (N_19489,N_18373,N_18121);
xor U19490 (N_19490,N_19189,N_18155);
nand U19491 (N_19491,N_18951,N_18239);
xnor U19492 (N_19492,N_18978,N_18018);
nand U19493 (N_19493,N_18714,N_19152);
and U19494 (N_19494,N_19109,N_18540);
nand U19495 (N_19495,N_18985,N_19015);
and U19496 (N_19496,N_18464,N_18013);
nand U19497 (N_19497,N_18472,N_18043);
nand U19498 (N_19498,N_18177,N_18232);
nor U19499 (N_19499,N_19053,N_18977);
and U19500 (N_19500,N_18749,N_18325);
xor U19501 (N_19501,N_18301,N_18976);
nand U19502 (N_19502,N_18249,N_18118);
nor U19503 (N_19503,N_19079,N_18428);
nor U19504 (N_19504,N_19083,N_18337);
or U19505 (N_19505,N_19154,N_18666);
nor U19506 (N_19506,N_18162,N_19000);
nand U19507 (N_19507,N_18849,N_18852);
nor U19508 (N_19508,N_18348,N_18764);
nor U19509 (N_19509,N_18753,N_18606);
or U19510 (N_19510,N_18000,N_18773);
or U19511 (N_19511,N_18124,N_18851);
and U19512 (N_19512,N_18635,N_18084);
and U19513 (N_19513,N_18202,N_18303);
nor U19514 (N_19514,N_18715,N_19100);
nand U19515 (N_19515,N_19196,N_18027);
nor U19516 (N_19516,N_18297,N_18994);
nor U19517 (N_19517,N_18642,N_18578);
xor U19518 (N_19518,N_18190,N_18598);
nor U19519 (N_19519,N_18139,N_19077);
nor U19520 (N_19520,N_18964,N_18775);
or U19521 (N_19521,N_18195,N_18023);
nand U19522 (N_19522,N_18846,N_18168);
and U19523 (N_19523,N_18510,N_18449);
and U19524 (N_19524,N_18762,N_18471);
or U19525 (N_19525,N_19167,N_18643);
nor U19526 (N_19526,N_18150,N_18378);
or U19527 (N_19527,N_19022,N_18105);
nand U19528 (N_19528,N_18395,N_18988);
and U19529 (N_19529,N_18663,N_18501);
nand U19530 (N_19530,N_18234,N_19137);
or U19531 (N_19531,N_18668,N_18512);
xnor U19532 (N_19532,N_18317,N_18360);
xnor U19533 (N_19533,N_18524,N_19071);
xor U19534 (N_19534,N_19130,N_18729);
nand U19535 (N_19535,N_18016,N_18960);
and U19536 (N_19536,N_18550,N_18407);
or U19537 (N_19537,N_18736,N_18945);
and U19538 (N_19538,N_19176,N_18423);
and U19539 (N_19539,N_19033,N_18159);
xnor U19540 (N_19540,N_18950,N_18116);
xnor U19541 (N_19541,N_19030,N_18810);
xor U19542 (N_19542,N_18556,N_18093);
or U19543 (N_19543,N_18237,N_19144);
xnor U19544 (N_19544,N_19064,N_18535);
or U19545 (N_19545,N_18740,N_18418);
and U19546 (N_19546,N_18563,N_19014);
and U19547 (N_19547,N_18901,N_18453);
or U19548 (N_19548,N_19116,N_18221);
or U19549 (N_19549,N_18803,N_18504);
and U19550 (N_19550,N_18146,N_18566);
xnor U19551 (N_19551,N_18163,N_18425);
and U19552 (N_19552,N_18683,N_18397);
and U19553 (N_19553,N_18157,N_18362);
nand U19554 (N_19554,N_18522,N_18986);
xor U19555 (N_19555,N_18112,N_19052);
xnor U19556 (N_19556,N_18702,N_18271);
or U19557 (N_19557,N_18701,N_18141);
nor U19558 (N_19558,N_18788,N_18414);
nor U19559 (N_19559,N_18446,N_18601);
nor U19560 (N_19560,N_18890,N_18968);
nor U19561 (N_19561,N_19135,N_18827);
xor U19562 (N_19562,N_18889,N_18574);
nand U19563 (N_19563,N_18823,N_19087);
nor U19564 (N_19564,N_18352,N_18491);
xor U19565 (N_19565,N_18231,N_18514);
or U19566 (N_19566,N_18477,N_18603);
nor U19567 (N_19567,N_18529,N_18402);
nand U19568 (N_19568,N_18786,N_18318);
xnor U19569 (N_19569,N_18063,N_18653);
or U19570 (N_19570,N_18080,N_18748);
or U19571 (N_19571,N_18551,N_18927);
and U19572 (N_19572,N_18725,N_18059);
or U19573 (N_19573,N_19010,N_18212);
or U19574 (N_19574,N_18126,N_18892);
and U19575 (N_19575,N_18284,N_18096);
and U19576 (N_19576,N_18329,N_18136);
nand U19577 (N_19577,N_18581,N_18272);
nand U19578 (N_19578,N_18427,N_18319);
nand U19579 (N_19579,N_19007,N_18045);
nor U19580 (N_19580,N_19199,N_19084);
nor U19581 (N_19581,N_19139,N_18308);
xnor U19582 (N_19582,N_18074,N_18010);
xor U19583 (N_19583,N_18991,N_18813);
nand U19584 (N_19584,N_19129,N_18180);
nand U19585 (N_19585,N_18527,N_18757);
xor U19586 (N_19586,N_18287,N_19040);
or U19587 (N_19587,N_18460,N_18026);
and U19588 (N_19588,N_19093,N_18583);
nor U19589 (N_19589,N_18806,N_18981);
nor U19590 (N_19590,N_18184,N_18357);
xnor U19591 (N_19591,N_18752,N_18506);
nor U19592 (N_19592,N_18887,N_18439);
nand U19593 (N_19593,N_18456,N_19160);
nand U19594 (N_19594,N_18531,N_18768);
xnor U19595 (N_19595,N_18685,N_18932);
nor U19596 (N_19596,N_18792,N_18376);
xor U19597 (N_19597,N_18364,N_18021);
nor U19598 (N_19598,N_18636,N_18576);
nand U19599 (N_19599,N_19065,N_18870);
and U19600 (N_19600,N_19090,N_19166);
or U19601 (N_19601,N_18292,N_18244);
nand U19602 (N_19602,N_18142,N_18207);
or U19603 (N_19603,N_18621,N_18442);
and U19604 (N_19604,N_18819,N_18310);
or U19605 (N_19605,N_18961,N_18091);
or U19606 (N_19606,N_18859,N_19012);
nor U19607 (N_19607,N_19168,N_18164);
xor U19608 (N_19608,N_18667,N_18875);
nor U19609 (N_19609,N_18444,N_18634);
nor U19610 (N_19610,N_18435,N_18537);
nand U19611 (N_19611,N_18882,N_18349);
and U19612 (N_19612,N_18233,N_18944);
nor U19613 (N_19613,N_18799,N_19107);
nor U19614 (N_19614,N_18916,N_19091);
xor U19615 (N_19615,N_18502,N_18189);
xnor U19616 (N_19616,N_18149,N_18182);
nor U19617 (N_19617,N_19113,N_18705);
and U19618 (N_19618,N_18330,N_18833);
or U19619 (N_19619,N_18341,N_18588);
xor U19620 (N_19620,N_19062,N_19179);
or U19621 (N_19621,N_19081,N_18222);
nor U19622 (N_19622,N_18391,N_18934);
xor U19623 (N_19623,N_18704,N_18493);
xnor U19624 (N_19624,N_18829,N_18671);
and U19625 (N_19625,N_19104,N_18684);
xnor U19626 (N_19626,N_19072,N_18248);
nor U19627 (N_19627,N_18759,N_18327);
nor U19628 (N_19628,N_18377,N_18354);
xor U19629 (N_19629,N_19066,N_19101);
xnor U19630 (N_19630,N_18336,N_18173);
nor U19631 (N_19631,N_19026,N_18893);
and U19632 (N_19632,N_18210,N_18046);
nand U19633 (N_19633,N_18959,N_18979);
or U19634 (N_19634,N_18097,N_18172);
xnor U19635 (N_19635,N_18238,N_19102);
or U19636 (N_19636,N_18982,N_18030);
and U19637 (N_19637,N_18553,N_18350);
or U19638 (N_19638,N_18913,N_18677);
nand U19639 (N_19639,N_18313,N_18368);
xnor U19640 (N_19640,N_18876,N_18490);
nand U19641 (N_19641,N_18921,N_18392);
and U19642 (N_19642,N_18682,N_18508);
or U19643 (N_19643,N_18618,N_19184);
xnor U19644 (N_19644,N_18152,N_18790);
or U19645 (N_19645,N_18487,N_18741);
nand U19646 (N_19646,N_18036,N_18541);
or U19647 (N_19647,N_18165,N_18914);
or U19648 (N_19648,N_19024,N_18375);
xnor U19649 (N_19649,N_18593,N_19060);
xor U19650 (N_19650,N_18793,N_18595);
nand U19651 (N_19651,N_19156,N_18723);
nor U19652 (N_19652,N_18861,N_18260);
or U19653 (N_19653,N_18903,N_18648);
and U19654 (N_19654,N_18197,N_19149);
nor U19655 (N_19655,N_18426,N_18885);
and U19656 (N_19656,N_18765,N_18358);
and U19657 (N_19657,N_18573,N_19180);
nand U19658 (N_19658,N_18206,N_18815);
and U19659 (N_19659,N_19038,N_19045);
or U19660 (N_19660,N_19016,N_19069);
or U19661 (N_19661,N_18119,N_19094);
or U19662 (N_19662,N_19111,N_18293);
nand U19663 (N_19663,N_18217,N_18623);
and U19664 (N_19664,N_19112,N_18532);
nand U19665 (N_19665,N_18655,N_19155);
xor U19666 (N_19666,N_19004,N_18820);
nand U19667 (N_19667,N_18286,N_18263);
nand U19668 (N_19668,N_18015,N_18615);
and U19669 (N_19669,N_18993,N_18505);
nor U19670 (N_19670,N_19170,N_18585);
nor U19671 (N_19671,N_18060,N_18219);
or U19672 (N_19672,N_18058,N_18517);
xor U19673 (N_19673,N_18662,N_19027);
nor U19674 (N_19674,N_18641,N_18549);
nand U19675 (N_19675,N_18089,N_18224);
nand U19676 (N_19676,N_18448,N_18963);
or U19677 (N_19677,N_18247,N_19142);
nand U19678 (N_19678,N_18943,N_18147);
and U19679 (N_19679,N_18534,N_18497);
and U19680 (N_19680,N_19044,N_18077);
nand U19681 (N_19681,N_18949,N_18294);
and U19682 (N_19682,N_18004,N_18518);
nor U19683 (N_19683,N_18429,N_18035);
xor U19684 (N_19684,N_19172,N_18693);
or U19685 (N_19685,N_18948,N_18401);
nor U19686 (N_19686,N_18064,N_18866);
xnor U19687 (N_19687,N_18783,N_18267);
nand U19688 (N_19688,N_18185,N_18420);
nor U19689 (N_19689,N_18381,N_19120);
and U19690 (N_19690,N_18370,N_18970);
or U19691 (N_19691,N_18079,N_18897);
and U19692 (N_19692,N_18955,N_18839);
or U19693 (N_19693,N_19173,N_19096);
or U19694 (N_19694,N_19164,N_18841);
or U19695 (N_19695,N_18346,N_18160);
and U19696 (N_19696,N_18809,N_18176);
nand U19697 (N_19697,N_18707,N_18992);
or U19698 (N_19698,N_18129,N_18946);
and U19699 (N_19699,N_19191,N_18672);
and U19700 (N_19700,N_18289,N_18974);
nand U19701 (N_19701,N_18731,N_18836);
nand U19702 (N_19702,N_18156,N_18135);
or U19703 (N_19703,N_18309,N_18040);
or U19704 (N_19704,N_18896,N_18259);
or U19705 (N_19705,N_18716,N_18203);
nand U19706 (N_19706,N_18910,N_18755);
or U19707 (N_19707,N_19185,N_19075);
nor U19708 (N_19708,N_18417,N_18952);
nand U19709 (N_19709,N_18270,N_18389);
nand U19710 (N_19710,N_18520,N_18698);
xnor U19711 (N_19711,N_18400,N_18888);
xnor U19712 (N_19712,N_18047,N_18343);
nand U19713 (N_19713,N_18143,N_18600);
and U19714 (N_19714,N_18711,N_18624);
nand U19715 (N_19715,N_18072,N_18918);
xor U19716 (N_19716,N_18393,N_19193);
or U19717 (N_19717,N_19003,N_18791);
nand U19718 (N_19718,N_18796,N_18834);
xnor U19719 (N_19719,N_18338,N_18843);
and U19720 (N_19720,N_19050,N_18050);
nand U19721 (N_19721,N_18552,N_18485);
or U19722 (N_19722,N_19141,N_19106);
and U19723 (N_19723,N_18499,N_18957);
xnor U19724 (N_19724,N_18169,N_18780);
nor U19725 (N_19725,N_19098,N_18697);
nor U19726 (N_19726,N_19124,N_18687);
nand U19727 (N_19727,N_18273,N_18572);
nand U19728 (N_19728,N_18626,N_19188);
or U19729 (N_19729,N_18416,N_18331);
nand U19730 (N_19730,N_18877,N_18192);
or U19731 (N_19731,N_18902,N_19146);
or U19732 (N_19732,N_18919,N_19020);
nand U19733 (N_19733,N_18387,N_18218);
or U19734 (N_19734,N_18777,N_18469);
and U19735 (N_19735,N_18717,N_18840);
and U19736 (N_19736,N_18630,N_18411);
nor U19737 (N_19737,N_18412,N_18342);
nand U19738 (N_19738,N_18941,N_18536);
xor U19739 (N_19739,N_18344,N_18068);
or U19740 (N_19740,N_18845,N_18138);
and U19741 (N_19741,N_18379,N_19095);
xnor U19742 (N_19742,N_18153,N_18351);
or U19743 (N_19743,N_19097,N_18223);
or U19744 (N_19744,N_18031,N_18622);
xnor U19745 (N_19745,N_18528,N_18196);
nand U19746 (N_19746,N_18492,N_18915);
or U19747 (N_19747,N_19080,N_18743);
and U19748 (N_19748,N_18789,N_18804);
nor U19749 (N_19749,N_18005,N_19161);
nand U19750 (N_19750,N_18905,N_18719);
nand U19751 (N_19751,N_18967,N_18073);
nand U19752 (N_19752,N_18928,N_18555);
nand U19753 (N_19753,N_18486,N_18954);
or U19754 (N_19754,N_19005,N_18582);
and U19755 (N_19755,N_18571,N_19008);
nand U19756 (N_19756,N_18028,N_18148);
or U19757 (N_19757,N_18476,N_18300);
or U19758 (N_19758,N_18894,N_18382);
nor U19759 (N_19759,N_18856,N_18599);
and U19760 (N_19760,N_18754,N_18304);
or U19761 (N_19761,N_19043,N_19034);
nand U19762 (N_19762,N_18245,N_18388);
and U19763 (N_19763,N_19070,N_18507);
xor U19764 (N_19764,N_18760,N_18906);
or U19765 (N_19765,N_19019,N_18436);
nand U19766 (N_19766,N_18315,N_18012);
nor U19767 (N_19767,N_18661,N_18703);
nor U19768 (N_19768,N_18880,N_18438);
nand U19769 (N_19769,N_18140,N_18258);
and U19770 (N_19770,N_18481,N_18465);
or U19771 (N_19771,N_18483,N_18929);
and U19772 (N_19772,N_18797,N_18462);
nor U19773 (N_19773,N_18092,N_18629);
xor U19774 (N_19774,N_18061,N_18480);
and U19775 (N_19775,N_18670,N_18053);
nand U19776 (N_19776,N_19036,N_18208);
nand U19777 (N_19777,N_18410,N_18213);
or U19778 (N_19778,N_18644,N_18559);
nor U19779 (N_19779,N_18432,N_18281);
or U19780 (N_19780,N_18235,N_19057);
and U19781 (N_19781,N_18766,N_18475);
xor U19782 (N_19782,N_18020,N_18656);
xor U19783 (N_19783,N_18561,N_19054);
nor U19784 (N_19784,N_19121,N_18935);
nand U19785 (N_19785,N_19181,N_18639);
nor U19786 (N_19786,N_19115,N_18467);
nand U19787 (N_19787,N_18538,N_18647);
nand U19788 (N_19788,N_18120,N_18099);
or U19789 (N_19789,N_18569,N_18488);
xor U19790 (N_19790,N_18965,N_18568);
and U19791 (N_19791,N_18115,N_18274);
or U19792 (N_19792,N_19039,N_18565);
and U19793 (N_19793,N_19143,N_19134);
nand U19794 (N_19794,N_18673,N_18369);
or U19795 (N_19795,N_18406,N_18617);
nor U19796 (N_19796,N_18253,N_19108);
and U19797 (N_19797,N_18863,N_18539);
or U19798 (N_19798,N_18108,N_18122);
nand U19799 (N_19799,N_19029,N_18884);
nor U19800 (N_19800,N_18875,N_18798);
nor U19801 (N_19801,N_18288,N_18863);
and U19802 (N_19802,N_18262,N_18729);
and U19803 (N_19803,N_18389,N_18779);
nand U19804 (N_19804,N_18675,N_18727);
nand U19805 (N_19805,N_18985,N_18338);
nand U19806 (N_19806,N_18315,N_18728);
nor U19807 (N_19807,N_18014,N_18350);
xor U19808 (N_19808,N_18208,N_19026);
nor U19809 (N_19809,N_18972,N_18815);
and U19810 (N_19810,N_18623,N_18978);
and U19811 (N_19811,N_18478,N_18102);
or U19812 (N_19812,N_18243,N_18257);
xor U19813 (N_19813,N_18039,N_18857);
and U19814 (N_19814,N_18758,N_18638);
nand U19815 (N_19815,N_18682,N_18864);
nor U19816 (N_19816,N_18295,N_18730);
nor U19817 (N_19817,N_18042,N_18538);
and U19818 (N_19818,N_18589,N_18375);
nor U19819 (N_19819,N_18281,N_18649);
nand U19820 (N_19820,N_18933,N_18217);
nand U19821 (N_19821,N_18858,N_19061);
xor U19822 (N_19822,N_18865,N_18877);
or U19823 (N_19823,N_18706,N_18431);
and U19824 (N_19824,N_18218,N_18992);
nor U19825 (N_19825,N_18819,N_18220);
nor U19826 (N_19826,N_18524,N_18837);
and U19827 (N_19827,N_18136,N_18414);
nor U19828 (N_19828,N_18769,N_18731);
xor U19829 (N_19829,N_18668,N_18662);
nor U19830 (N_19830,N_18509,N_18728);
nor U19831 (N_19831,N_18926,N_18526);
or U19832 (N_19832,N_18471,N_19139);
nor U19833 (N_19833,N_18952,N_18889);
xor U19834 (N_19834,N_18723,N_18477);
nand U19835 (N_19835,N_18401,N_18157);
nor U19836 (N_19836,N_18215,N_18760);
xor U19837 (N_19837,N_18833,N_18640);
nor U19838 (N_19838,N_18582,N_18017);
and U19839 (N_19839,N_18283,N_18627);
nor U19840 (N_19840,N_18629,N_19098);
nor U19841 (N_19841,N_18810,N_18669);
nor U19842 (N_19842,N_18280,N_19117);
or U19843 (N_19843,N_18404,N_18705);
or U19844 (N_19844,N_18642,N_18234);
xor U19845 (N_19845,N_18318,N_18385);
or U19846 (N_19846,N_18502,N_18335);
nand U19847 (N_19847,N_18190,N_18030);
nor U19848 (N_19848,N_18086,N_19068);
or U19849 (N_19849,N_18706,N_18028);
or U19850 (N_19850,N_19037,N_18728);
nand U19851 (N_19851,N_18153,N_18534);
xnor U19852 (N_19852,N_18737,N_18456);
xor U19853 (N_19853,N_18498,N_18084);
or U19854 (N_19854,N_18404,N_18044);
and U19855 (N_19855,N_19123,N_19114);
nor U19856 (N_19856,N_18045,N_18789);
nor U19857 (N_19857,N_18999,N_18990);
or U19858 (N_19858,N_18596,N_18163);
or U19859 (N_19859,N_18375,N_18571);
and U19860 (N_19860,N_19018,N_18810);
nand U19861 (N_19861,N_18772,N_18671);
or U19862 (N_19862,N_18995,N_18582);
and U19863 (N_19863,N_18248,N_18203);
and U19864 (N_19864,N_18636,N_18870);
xnor U19865 (N_19865,N_18475,N_18212);
nor U19866 (N_19866,N_18196,N_18509);
nor U19867 (N_19867,N_18370,N_18277);
and U19868 (N_19868,N_18939,N_18176);
or U19869 (N_19869,N_18428,N_18221);
nand U19870 (N_19870,N_18561,N_18385);
nor U19871 (N_19871,N_18440,N_18261);
xor U19872 (N_19872,N_18532,N_18075);
and U19873 (N_19873,N_18127,N_18449);
or U19874 (N_19874,N_18069,N_19093);
xor U19875 (N_19875,N_18896,N_18616);
and U19876 (N_19876,N_18066,N_18777);
xnor U19877 (N_19877,N_18999,N_18515);
xnor U19878 (N_19878,N_18544,N_18430);
and U19879 (N_19879,N_18542,N_19122);
and U19880 (N_19880,N_18808,N_18595);
nor U19881 (N_19881,N_18749,N_18878);
or U19882 (N_19882,N_18149,N_18337);
xor U19883 (N_19883,N_18688,N_19052);
nand U19884 (N_19884,N_19090,N_18933);
or U19885 (N_19885,N_18548,N_18524);
and U19886 (N_19886,N_18250,N_18683);
nand U19887 (N_19887,N_18565,N_18270);
or U19888 (N_19888,N_18986,N_18316);
nor U19889 (N_19889,N_18032,N_18409);
xor U19890 (N_19890,N_18903,N_18752);
nand U19891 (N_19891,N_18765,N_18471);
nor U19892 (N_19892,N_18287,N_18030);
nand U19893 (N_19893,N_18139,N_18416);
nand U19894 (N_19894,N_18763,N_18287);
nor U19895 (N_19895,N_18360,N_18845);
and U19896 (N_19896,N_18995,N_18344);
and U19897 (N_19897,N_18836,N_18022);
and U19898 (N_19898,N_18153,N_18337);
and U19899 (N_19899,N_18364,N_19144);
and U19900 (N_19900,N_18542,N_18173);
or U19901 (N_19901,N_19108,N_18218);
xnor U19902 (N_19902,N_18417,N_19188);
xnor U19903 (N_19903,N_18343,N_18211);
nand U19904 (N_19904,N_18120,N_18407);
and U19905 (N_19905,N_18309,N_18575);
xnor U19906 (N_19906,N_18222,N_18422);
or U19907 (N_19907,N_18909,N_19001);
or U19908 (N_19908,N_18035,N_18424);
or U19909 (N_19909,N_18694,N_18310);
xnor U19910 (N_19910,N_18263,N_18219);
and U19911 (N_19911,N_18606,N_18619);
xor U19912 (N_19912,N_18376,N_18720);
and U19913 (N_19913,N_18049,N_18586);
and U19914 (N_19914,N_19114,N_18928);
and U19915 (N_19915,N_18533,N_18305);
nor U19916 (N_19916,N_19064,N_18977);
and U19917 (N_19917,N_18078,N_19033);
nor U19918 (N_19918,N_18963,N_18471);
nand U19919 (N_19919,N_18303,N_18819);
or U19920 (N_19920,N_19031,N_18219);
and U19921 (N_19921,N_18633,N_18672);
and U19922 (N_19922,N_18016,N_19179);
nor U19923 (N_19923,N_19129,N_18741);
xnor U19924 (N_19924,N_18421,N_18799);
or U19925 (N_19925,N_18743,N_19175);
and U19926 (N_19926,N_18900,N_18842);
nor U19927 (N_19927,N_18750,N_18025);
xor U19928 (N_19928,N_18699,N_18380);
or U19929 (N_19929,N_18111,N_19045);
xor U19930 (N_19930,N_18106,N_18443);
and U19931 (N_19931,N_18901,N_18144);
and U19932 (N_19932,N_19125,N_18721);
and U19933 (N_19933,N_18937,N_18408);
nor U19934 (N_19934,N_19135,N_19187);
and U19935 (N_19935,N_18377,N_18337);
and U19936 (N_19936,N_18100,N_18915);
nand U19937 (N_19937,N_18111,N_18497);
nand U19938 (N_19938,N_18385,N_19128);
and U19939 (N_19939,N_18122,N_18283);
xor U19940 (N_19940,N_18600,N_18697);
xor U19941 (N_19941,N_18904,N_18143);
nor U19942 (N_19942,N_18155,N_18062);
xor U19943 (N_19943,N_18315,N_18253);
xnor U19944 (N_19944,N_18309,N_18151);
nand U19945 (N_19945,N_18910,N_18160);
or U19946 (N_19946,N_18701,N_18065);
nor U19947 (N_19947,N_18096,N_18398);
nand U19948 (N_19948,N_18376,N_18815);
or U19949 (N_19949,N_18749,N_18558);
nor U19950 (N_19950,N_18447,N_18712);
or U19951 (N_19951,N_18756,N_18890);
xnor U19952 (N_19952,N_19081,N_18185);
nor U19953 (N_19953,N_19088,N_18578);
nor U19954 (N_19954,N_18772,N_18533);
xor U19955 (N_19955,N_19081,N_18991);
and U19956 (N_19956,N_18222,N_18252);
xnor U19957 (N_19957,N_18303,N_19039);
nor U19958 (N_19958,N_18873,N_18611);
or U19959 (N_19959,N_18589,N_18826);
nand U19960 (N_19960,N_18508,N_18963);
xnor U19961 (N_19961,N_18504,N_18908);
and U19962 (N_19962,N_18169,N_18659);
nor U19963 (N_19963,N_18706,N_18561);
or U19964 (N_19964,N_18447,N_18558);
nand U19965 (N_19965,N_19151,N_18742);
nor U19966 (N_19966,N_18300,N_18861);
xor U19967 (N_19967,N_18441,N_18043);
or U19968 (N_19968,N_19179,N_18989);
nand U19969 (N_19969,N_18084,N_18510);
nand U19970 (N_19970,N_18506,N_18846);
or U19971 (N_19971,N_19144,N_18386);
or U19972 (N_19972,N_18256,N_18078);
and U19973 (N_19973,N_18541,N_18952);
nor U19974 (N_19974,N_18879,N_18028);
nand U19975 (N_19975,N_18405,N_18175);
or U19976 (N_19976,N_18822,N_18347);
xnor U19977 (N_19977,N_18878,N_18691);
nand U19978 (N_19978,N_18587,N_18044);
or U19979 (N_19979,N_18558,N_18500);
nand U19980 (N_19980,N_18751,N_18628);
xnor U19981 (N_19981,N_18425,N_18110);
xnor U19982 (N_19982,N_18167,N_18189);
nand U19983 (N_19983,N_18204,N_18295);
or U19984 (N_19984,N_19002,N_18964);
or U19985 (N_19985,N_18963,N_19000);
xor U19986 (N_19986,N_18169,N_18338);
and U19987 (N_19987,N_18195,N_18381);
xnor U19988 (N_19988,N_19001,N_18763);
nand U19989 (N_19989,N_18513,N_18460);
xor U19990 (N_19990,N_19117,N_18824);
xor U19991 (N_19991,N_18036,N_18835);
and U19992 (N_19992,N_18180,N_18798);
or U19993 (N_19993,N_18583,N_18569);
or U19994 (N_19994,N_18289,N_18801);
or U19995 (N_19995,N_18425,N_18893);
and U19996 (N_19996,N_18623,N_18710);
or U19997 (N_19997,N_18089,N_18678);
and U19998 (N_19998,N_18182,N_19064);
nor U19999 (N_19999,N_18344,N_18674);
and U20000 (N_20000,N_18456,N_19190);
xor U20001 (N_20001,N_18174,N_18343);
xnor U20002 (N_20002,N_18742,N_18600);
or U20003 (N_20003,N_18951,N_18291);
nand U20004 (N_20004,N_19038,N_18137);
nand U20005 (N_20005,N_18906,N_18860);
nor U20006 (N_20006,N_18464,N_19051);
xor U20007 (N_20007,N_18839,N_18185);
xnor U20008 (N_20008,N_19088,N_18300);
nand U20009 (N_20009,N_18696,N_18673);
nand U20010 (N_20010,N_19065,N_18220);
and U20011 (N_20011,N_19152,N_18055);
and U20012 (N_20012,N_18357,N_19049);
and U20013 (N_20013,N_18188,N_18602);
nor U20014 (N_20014,N_18255,N_18525);
or U20015 (N_20015,N_19092,N_18086);
nor U20016 (N_20016,N_18295,N_18102);
nor U20017 (N_20017,N_18085,N_18798);
nand U20018 (N_20018,N_19125,N_18304);
and U20019 (N_20019,N_19192,N_18461);
nor U20020 (N_20020,N_19021,N_18602);
xor U20021 (N_20021,N_19130,N_18802);
xnor U20022 (N_20022,N_18108,N_18582);
and U20023 (N_20023,N_19182,N_19170);
and U20024 (N_20024,N_18746,N_18933);
nor U20025 (N_20025,N_18388,N_18168);
or U20026 (N_20026,N_18737,N_18409);
nand U20027 (N_20027,N_18399,N_18869);
or U20028 (N_20028,N_18481,N_18255);
and U20029 (N_20029,N_18419,N_18504);
and U20030 (N_20030,N_19100,N_18052);
or U20031 (N_20031,N_18861,N_19144);
or U20032 (N_20032,N_18405,N_18196);
or U20033 (N_20033,N_18297,N_18746);
nand U20034 (N_20034,N_18574,N_18636);
xnor U20035 (N_20035,N_18951,N_18938);
nor U20036 (N_20036,N_18091,N_18099);
nor U20037 (N_20037,N_18579,N_18092);
nor U20038 (N_20038,N_18919,N_18188);
xnor U20039 (N_20039,N_18720,N_18918);
nor U20040 (N_20040,N_18055,N_18591);
nand U20041 (N_20041,N_18038,N_18831);
and U20042 (N_20042,N_18418,N_18733);
nand U20043 (N_20043,N_19147,N_18995);
or U20044 (N_20044,N_18717,N_18360);
nand U20045 (N_20045,N_19133,N_18271);
xor U20046 (N_20046,N_18788,N_18685);
nor U20047 (N_20047,N_18766,N_18025);
xnor U20048 (N_20048,N_18565,N_18274);
or U20049 (N_20049,N_18927,N_18825);
or U20050 (N_20050,N_18513,N_18139);
or U20051 (N_20051,N_18175,N_19033);
and U20052 (N_20052,N_18066,N_18006);
nand U20053 (N_20053,N_18005,N_18997);
or U20054 (N_20054,N_18104,N_19076);
xnor U20055 (N_20055,N_18112,N_18235);
nor U20056 (N_20056,N_18407,N_18714);
or U20057 (N_20057,N_18890,N_18545);
and U20058 (N_20058,N_19114,N_18213);
nand U20059 (N_20059,N_18225,N_18807);
nor U20060 (N_20060,N_18881,N_18192);
and U20061 (N_20061,N_18595,N_18272);
and U20062 (N_20062,N_19158,N_18968);
or U20063 (N_20063,N_18839,N_18040);
nand U20064 (N_20064,N_18155,N_18793);
nand U20065 (N_20065,N_18483,N_18984);
nor U20066 (N_20066,N_18820,N_18309);
and U20067 (N_20067,N_19090,N_19174);
or U20068 (N_20068,N_18289,N_18757);
and U20069 (N_20069,N_18915,N_18907);
xor U20070 (N_20070,N_18265,N_18461);
or U20071 (N_20071,N_18687,N_19155);
or U20072 (N_20072,N_18238,N_18977);
nor U20073 (N_20073,N_18702,N_18692);
nand U20074 (N_20074,N_18193,N_18127);
nand U20075 (N_20075,N_18385,N_18311);
nor U20076 (N_20076,N_19182,N_19096);
or U20077 (N_20077,N_18800,N_18124);
xor U20078 (N_20078,N_18822,N_19018);
or U20079 (N_20079,N_18596,N_18117);
xnor U20080 (N_20080,N_18263,N_18410);
and U20081 (N_20081,N_18412,N_18263);
nor U20082 (N_20082,N_18877,N_18001);
and U20083 (N_20083,N_18258,N_18469);
xnor U20084 (N_20084,N_18422,N_18754);
and U20085 (N_20085,N_19104,N_19044);
nor U20086 (N_20086,N_19117,N_18750);
nand U20087 (N_20087,N_18522,N_18000);
nor U20088 (N_20088,N_18252,N_19138);
and U20089 (N_20089,N_18966,N_18112);
xnor U20090 (N_20090,N_18928,N_18265);
xnor U20091 (N_20091,N_18863,N_18019);
nand U20092 (N_20092,N_18260,N_18755);
nor U20093 (N_20093,N_18492,N_19031);
nor U20094 (N_20094,N_18612,N_18432);
or U20095 (N_20095,N_18538,N_19161);
or U20096 (N_20096,N_18999,N_18612);
or U20097 (N_20097,N_18837,N_18931);
nor U20098 (N_20098,N_18841,N_19174);
or U20099 (N_20099,N_18949,N_18095);
and U20100 (N_20100,N_19176,N_18139);
or U20101 (N_20101,N_18487,N_18210);
xnor U20102 (N_20102,N_18345,N_18916);
or U20103 (N_20103,N_18980,N_18578);
xor U20104 (N_20104,N_18788,N_18881);
and U20105 (N_20105,N_18963,N_18411);
nor U20106 (N_20106,N_18111,N_19024);
nand U20107 (N_20107,N_18774,N_18216);
nand U20108 (N_20108,N_18479,N_18766);
nand U20109 (N_20109,N_19136,N_18263);
nand U20110 (N_20110,N_18479,N_18800);
or U20111 (N_20111,N_18128,N_19117);
nand U20112 (N_20112,N_18621,N_19040);
nand U20113 (N_20113,N_18886,N_19107);
xnor U20114 (N_20114,N_18294,N_18391);
or U20115 (N_20115,N_19047,N_19154);
nand U20116 (N_20116,N_18605,N_18507);
nand U20117 (N_20117,N_18538,N_18724);
nor U20118 (N_20118,N_18129,N_18516);
and U20119 (N_20119,N_18398,N_18159);
xnor U20120 (N_20120,N_18351,N_18837);
nor U20121 (N_20121,N_18654,N_18704);
nor U20122 (N_20122,N_18852,N_19127);
xnor U20123 (N_20123,N_19162,N_18729);
or U20124 (N_20124,N_18825,N_18200);
nand U20125 (N_20125,N_18620,N_18216);
xnor U20126 (N_20126,N_18161,N_19067);
xnor U20127 (N_20127,N_19179,N_18764);
xnor U20128 (N_20128,N_19198,N_19034);
nor U20129 (N_20129,N_18985,N_18747);
nor U20130 (N_20130,N_18104,N_18474);
or U20131 (N_20131,N_18963,N_18396);
nand U20132 (N_20132,N_18097,N_18404);
xor U20133 (N_20133,N_18113,N_19083);
or U20134 (N_20134,N_19041,N_18912);
or U20135 (N_20135,N_18641,N_18157);
or U20136 (N_20136,N_18875,N_19114);
and U20137 (N_20137,N_18946,N_19055);
nor U20138 (N_20138,N_18027,N_18697);
nor U20139 (N_20139,N_18569,N_18955);
nand U20140 (N_20140,N_18612,N_19068);
nand U20141 (N_20141,N_18902,N_18108);
or U20142 (N_20142,N_18300,N_18659);
or U20143 (N_20143,N_18592,N_19122);
nor U20144 (N_20144,N_18496,N_18017);
nand U20145 (N_20145,N_18967,N_18002);
nand U20146 (N_20146,N_18039,N_19139);
xnor U20147 (N_20147,N_18572,N_18410);
and U20148 (N_20148,N_19131,N_19054);
nor U20149 (N_20149,N_18408,N_18852);
and U20150 (N_20150,N_18819,N_18739);
and U20151 (N_20151,N_19021,N_18134);
xor U20152 (N_20152,N_18149,N_19020);
and U20153 (N_20153,N_18223,N_18431);
nand U20154 (N_20154,N_18566,N_18631);
nor U20155 (N_20155,N_18646,N_18418);
and U20156 (N_20156,N_18920,N_18717);
nor U20157 (N_20157,N_18918,N_18293);
nor U20158 (N_20158,N_18650,N_18008);
xor U20159 (N_20159,N_18408,N_18452);
nand U20160 (N_20160,N_18513,N_18196);
xnor U20161 (N_20161,N_18941,N_18322);
nand U20162 (N_20162,N_19075,N_18245);
or U20163 (N_20163,N_18494,N_18997);
and U20164 (N_20164,N_18681,N_18021);
or U20165 (N_20165,N_18051,N_18481);
nand U20166 (N_20166,N_18280,N_18516);
or U20167 (N_20167,N_18694,N_18007);
xor U20168 (N_20168,N_19112,N_18681);
nor U20169 (N_20169,N_18008,N_18335);
nor U20170 (N_20170,N_18509,N_18566);
xor U20171 (N_20171,N_18620,N_18125);
nand U20172 (N_20172,N_19061,N_18267);
nand U20173 (N_20173,N_19061,N_18239);
xor U20174 (N_20174,N_18179,N_18048);
nand U20175 (N_20175,N_18323,N_18920);
xor U20176 (N_20176,N_18772,N_18739);
and U20177 (N_20177,N_18797,N_18832);
and U20178 (N_20178,N_19081,N_18111);
xnor U20179 (N_20179,N_18366,N_18766);
xor U20180 (N_20180,N_18825,N_18494);
nor U20181 (N_20181,N_18138,N_18438);
or U20182 (N_20182,N_19106,N_18383);
and U20183 (N_20183,N_18095,N_18866);
and U20184 (N_20184,N_19053,N_18100);
xor U20185 (N_20185,N_18802,N_18063);
nor U20186 (N_20186,N_18668,N_18131);
nand U20187 (N_20187,N_18511,N_19176);
and U20188 (N_20188,N_18994,N_18004);
and U20189 (N_20189,N_18066,N_18243);
or U20190 (N_20190,N_19107,N_18984);
nor U20191 (N_20191,N_19134,N_19107);
nor U20192 (N_20192,N_19106,N_18949);
nor U20193 (N_20193,N_19012,N_18521);
and U20194 (N_20194,N_18166,N_19094);
nand U20195 (N_20195,N_18280,N_18261);
nor U20196 (N_20196,N_18626,N_19056);
and U20197 (N_20197,N_18664,N_18518);
nor U20198 (N_20198,N_18793,N_18097);
nand U20199 (N_20199,N_18965,N_18653);
and U20200 (N_20200,N_18237,N_19186);
and U20201 (N_20201,N_18278,N_18756);
or U20202 (N_20202,N_18206,N_19120);
xor U20203 (N_20203,N_19092,N_18455);
and U20204 (N_20204,N_18293,N_18832);
xor U20205 (N_20205,N_18079,N_18103);
nor U20206 (N_20206,N_19120,N_18395);
and U20207 (N_20207,N_18220,N_19170);
or U20208 (N_20208,N_18763,N_18530);
or U20209 (N_20209,N_18225,N_18153);
or U20210 (N_20210,N_18295,N_19015);
nor U20211 (N_20211,N_18569,N_19190);
and U20212 (N_20212,N_18928,N_19151);
and U20213 (N_20213,N_18846,N_18187);
or U20214 (N_20214,N_18811,N_19007);
xnor U20215 (N_20215,N_18057,N_18959);
xnor U20216 (N_20216,N_18445,N_18983);
and U20217 (N_20217,N_18297,N_18142);
nor U20218 (N_20218,N_19128,N_18066);
nand U20219 (N_20219,N_18621,N_18510);
or U20220 (N_20220,N_18940,N_18814);
nand U20221 (N_20221,N_19104,N_18918);
or U20222 (N_20222,N_19074,N_18288);
or U20223 (N_20223,N_18176,N_18303);
and U20224 (N_20224,N_18062,N_19051);
nand U20225 (N_20225,N_18927,N_18989);
xor U20226 (N_20226,N_19015,N_18924);
nor U20227 (N_20227,N_18086,N_19058);
nor U20228 (N_20228,N_18559,N_19145);
xnor U20229 (N_20229,N_19066,N_19022);
nand U20230 (N_20230,N_18258,N_18788);
or U20231 (N_20231,N_18332,N_19190);
or U20232 (N_20232,N_18592,N_18448);
and U20233 (N_20233,N_18441,N_18458);
or U20234 (N_20234,N_18681,N_18523);
or U20235 (N_20235,N_18463,N_18373);
xor U20236 (N_20236,N_18725,N_18741);
or U20237 (N_20237,N_18275,N_19075);
nor U20238 (N_20238,N_18942,N_18921);
xnor U20239 (N_20239,N_18920,N_18301);
and U20240 (N_20240,N_18347,N_18915);
nand U20241 (N_20241,N_18400,N_18663);
and U20242 (N_20242,N_19086,N_19190);
nor U20243 (N_20243,N_18046,N_18172);
nand U20244 (N_20244,N_18981,N_18992);
or U20245 (N_20245,N_18179,N_19140);
nand U20246 (N_20246,N_18093,N_19121);
and U20247 (N_20247,N_18908,N_19021);
xnor U20248 (N_20248,N_18822,N_19176);
nor U20249 (N_20249,N_18831,N_18729);
and U20250 (N_20250,N_18486,N_18979);
xnor U20251 (N_20251,N_18165,N_18316);
or U20252 (N_20252,N_18214,N_18105);
nand U20253 (N_20253,N_18741,N_18426);
nand U20254 (N_20254,N_18724,N_18673);
nand U20255 (N_20255,N_18031,N_18629);
nor U20256 (N_20256,N_18183,N_18002);
nor U20257 (N_20257,N_18050,N_18601);
or U20258 (N_20258,N_18170,N_18853);
nor U20259 (N_20259,N_18505,N_18094);
xor U20260 (N_20260,N_18045,N_19085);
nor U20261 (N_20261,N_18425,N_18571);
or U20262 (N_20262,N_18655,N_18990);
xnor U20263 (N_20263,N_18247,N_18352);
nor U20264 (N_20264,N_18941,N_18525);
nor U20265 (N_20265,N_18729,N_18823);
xor U20266 (N_20266,N_18336,N_18752);
xnor U20267 (N_20267,N_18257,N_18116);
or U20268 (N_20268,N_18021,N_18057);
xor U20269 (N_20269,N_19136,N_18672);
nand U20270 (N_20270,N_18863,N_18405);
nor U20271 (N_20271,N_18136,N_18536);
or U20272 (N_20272,N_19188,N_19001);
and U20273 (N_20273,N_18954,N_18514);
and U20274 (N_20274,N_18036,N_19008);
or U20275 (N_20275,N_18886,N_18666);
nand U20276 (N_20276,N_18719,N_18380);
and U20277 (N_20277,N_18569,N_18308);
nand U20278 (N_20278,N_18028,N_18898);
or U20279 (N_20279,N_19193,N_19041);
nor U20280 (N_20280,N_18970,N_19189);
xor U20281 (N_20281,N_18472,N_18623);
xnor U20282 (N_20282,N_19003,N_18540);
nand U20283 (N_20283,N_18601,N_18114);
nor U20284 (N_20284,N_19075,N_18775);
nand U20285 (N_20285,N_18679,N_18925);
xnor U20286 (N_20286,N_18578,N_18842);
nand U20287 (N_20287,N_18519,N_18829);
xor U20288 (N_20288,N_18741,N_18207);
xor U20289 (N_20289,N_19089,N_18174);
xor U20290 (N_20290,N_18342,N_18583);
xor U20291 (N_20291,N_18393,N_18849);
nand U20292 (N_20292,N_18556,N_18153);
nor U20293 (N_20293,N_18973,N_18558);
nor U20294 (N_20294,N_19110,N_18798);
nand U20295 (N_20295,N_18789,N_18518);
nand U20296 (N_20296,N_18270,N_18377);
nand U20297 (N_20297,N_18880,N_18209);
or U20298 (N_20298,N_18746,N_18575);
nand U20299 (N_20299,N_18259,N_18270);
or U20300 (N_20300,N_18805,N_18260);
or U20301 (N_20301,N_18505,N_18797);
xnor U20302 (N_20302,N_18242,N_18582);
and U20303 (N_20303,N_18815,N_18391);
or U20304 (N_20304,N_19108,N_18994);
and U20305 (N_20305,N_18777,N_18177);
xor U20306 (N_20306,N_19144,N_18635);
xor U20307 (N_20307,N_18935,N_18783);
nand U20308 (N_20308,N_18279,N_18707);
or U20309 (N_20309,N_18617,N_18978);
nor U20310 (N_20310,N_18798,N_18684);
nor U20311 (N_20311,N_18522,N_18157);
nor U20312 (N_20312,N_18645,N_18782);
nor U20313 (N_20313,N_18784,N_18604);
nand U20314 (N_20314,N_18851,N_19009);
xor U20315 (N_20315,N_18755,N_18461);
nor U20316 (N_20316,N_19095,N_18150);
nand U20317 (N_20317,N_18010,N_18143);
xor U20318 (N_20318,N_18372,N_18282);
nor U20319 (N_20319,N_19060,N_18072);
and U20320 (N_20320,N_19058,N_18560);
and U20321 (N_20321,N_19181,N_18873);
nor U20322 (N_20322,N_18754,N_18268);
and U20323 (N_20323,N_18946,N_18538);
xor U20324 (N_20324,N_19159,N_18786);
xnor U20325 (N_20325,N_18667,N_18020);
or U20326 (N_20326,N_18309,N_18972);
or U20327 (N_20327,N_18765,N_18145);
or U20328 (N_20328,N_19152,N_19017);
nor U20329 (N_20329,N_18036,N_18589);
xor U20330 (N_20330,N_18730,N_18403);
nor U20331 (N_20331,N_18968,N_18228);
and U20332 (N_20332,N_18365,N_18673);
xnor U20333 (N_20333,N_18813,N_18244);
xnor U20334 (N_20334,N_18346,N_18536);
nor U20335 (N_20335,N_18522,N_18173);
and U20336 (N_20336,N_18242,N_18412);
or U20337 (N_20337,N_18290,N_18407);
and U20338 (N_20338,N_18806,N_18757);
nand U20339 (N_20339,N_18440,N_18539);
xnor U20340 (N_20340,N_19093,N_18952);
nor U20341 (N_20341,N_18623,N_19120);
and U20342 (N_20342,N_19110,N_18633);
and U20343 (N_20343,N_18907,N_18679);
nand U20344 (N_20344,N_18358,N_18859);
nor U20345 (N_20345,N_18982,N_18628);
or U20346 (N_20346,N_18056,N_18434);
nand U20347 (N_20347,N_19072,N_18603);
nand U20348 (N_20348,N_18495,N_18077);
xnor U20349 (N_20349,N_18530,N_19191);
or U20350 (N_20350,N_18877,N_18595);
and U20351 (N_20351,N_18901,N_18661);
or U20352 (N_20352,N_18426,N_18764);
xnor U20353 (N_20353,N_18957,N_19100);
or U20354 (N_20354,N_18515,N_18660);
and U20355 (N_20355,N_18018,N_19136);
or U20356 (N_20356,N_19162,N_18658);
nand U20357 (N_20357,N_18543,N_18999);
and U20358 (N_20358,N_19087,N_18278);
or U20359 (N_20359,N_18904,N_18115);
and U20360 (N_20360,N_18225,N_18589);
nor U20361 (N_20361,N_18758,N_19167);
and U20362 (N_20362,N_18664,N_18912);
and U20363 (N_20363,N_18986,N_18448);
nand U20364 (N_20364,N_18594,N_19180);
xnor U20365 (N_20365,N_18218,N_19136);
xnor U20366 (N_20366,N_18158,N_18725);
and U20367 (N_20367,N_18634,N_18051);
or U20368 (N_20368,N_18616,N_19005);
xor U20369 (N_20369,N_18814,N_18320);
nand U20370 (N_20370,N_18243,N_18496);
or U20371 (N_20371,N_18585,N_18175);
nand U20372 (N_20372,N_18958,N_18459);
nand U20373 (N_20373,N_18568,N_19004);
nand U20374 (N_20374,N_18610,N_18640);
or U20375 (N_20375,N_18163,N_18762);
xnor U20376 (N_20376,N_18323,N_18038);
or U20377 (N_20377,N_18414,N_18597);
and U20378 (N_20378,N_18371,N_18056);
or U20379 (N_20379,N_18224,N_18772);
or U20380 (N_20380,N_18537,N_18555);
nand U20381 (N_20381,N_18563,N_19059);
or U20382 (N_20382,N_18041,N_18007);
or U20383 (N_20383,N_18110,N_18208);
nor U20384 (N_20384,N_18409,N_18920);
nand U20385 (N_20385,N_18883,N_18587);
nand U20386 (N_20386,N_18122,N_18073);
and U20387 (N_20387,N_18126,N_18595);
and U20388 (N_20388,N_18624,N_18749);
and U20389 (N_20389,N_19169,N_18652);
and U20390 (N_20390,N_19051,N_19015);
nor U20391 (N_20391,N_18782,N_19044);
nand U20392 (N_20392,N_18634,N_19158);
nand U20393 (N_20393,N_18214,N_18309);
nand U20394 (N_20394,N_18203,N_18834);
nor U20395 (N_20395,N_19179,N_19025);
nor U20396 (N_20396,N_18136,N_19184);
nor U20397 (N_20397,N_18733,N_18225);
or U20398 (N_20398,N_18402,N_19132);
or U20399 (N_20399,N_18950,N_18602);
nor U20400 (N_20400,N_19565,N_20246);
and U20401 (N_20401,N_19920,N_19921);
xor U20402 (N_20402,N_20017,N_19884);
and U20403 (N_20403,N_19350,N_19213);
and U20404 (N_20404,N_19958,N_19239);
or U20405 (N_20405,N_19789,N_19811);
xor U20406 (N_20406,N_19232,N_19806);
xor U20407 (N_20407,N_19522,N_19781);
nand U20408 (N_20408,N_20025,N_19535);
nor U20409 (N_20409,N_19221,N_19798);
nor U20410 (N_20410,N_20126,N_19562);
nor U20411 (N_20411,N_20092,N_20322);
nor U20412 (N_20412,N_19340,N_19455);
and U20413 (N_20413,N_19477,N_19763);
nor U20414 (N_20414,N_19402,N_20082);
nor U20415 (N_20415,N_19331,N_19722);
and U20416 (N_20416,N_19587,N_20319);
nor U20417 (N_20417,N_19312,N_19447);
and U20418 (N_20418,N_19534,N_19652);
xor U20419 (N_20419,N_19995,N_19757);
and U20420 (N_20420,N_19924,N_20139);
and U20421 (N_20421,N_20137,N_20200);
nor U20422 (N_20422,N_19512,N_20250);
xnor U20423 (N_20423,N_19809,N_20018);
nand U20424 (N_20424,N_19904,N_19459);
or U20425 (N_20425,N_20163,N_19976);
nand U20426 (N_20426,N_20312,N_19880);
or U20427 (N_20427,N_20247,N_20243);
xnor U20428 (N_20428,N_20181,N_19807);
or U20429 (N_20429,N_20278,N_20012);
nor U20430 (N_20430,N_19753,N_19342);
and U20431 (N_20431,N_19698,N_19495);
and U20432 (N_20432,N_19865,N_19220);
nand U20433 (N_20433,N_19760,N_20081);
or U20434 (N_20434,N_19313,N_20015);
or U20435 (N_20435,N_19877,N_20021);
xnor U20436 (N_20436,N_19917,N_19665);
nor U20437 (N_20437,N_19623,N_20316);
and U20438 (N_20438,N_19317,N_20147);
and U20439 (N_20439,N_19887,N_19948);
nor U20440 (N_20440,N_19773,N_19597);
or U20441 (N_20441,N_19429,N_19386);
xnor U20442 (N_20442,N_19749,N_20135);
or U20443 (N_20443,N_19382,N_19970);
or U20444 (N_20444,N_19225,N_19859);
or U20445 (N_20445,N_19874,N_20372);
nand U20446 (N_20446,N_20209,N_19355);
nand U20447 (N_20447,N_20130,N_19266);
and U20448 (N_20448,N_19541,N_20220);
or U20449 (N_20449,N_19236,N_19554);
xor U20450 (N_20450,N_20393,N_19633);
nor U20451 (N_20451,N_19476,N_19369);
or U20452 (N_20452,N_19205,N_20396);
xor U20453 (N_20453,N_19854,N_19758);
nand U20454 (N_20454,N_20370,N_20381);
nor U20455 (N_20455,N_19460,N_20368);
and U20456 (N_20456,N_19523,N_19850);
nor U20457 (N_20457,N_19638,N_20167);
nor U20458 (N_20458,N_19822,N_20338);
nand U20459 (N_20459,N_19670,N_19234);
xor U20460 (N_20460,N_20383,N_19388);
and U20461 (N_20461,N_19546,N_19463);
xor U20462 (N_20462,N_20307,N_19249);
nor U20463 (N_20463,N_20310,N_20212);
nand U20464 (N_20464,N_19991,N_20028);
nor U20465 (N_20465,N_19242,N_19932);
xor U20466 (N_20466,N_20303,N_19935);
nand U20467 (N_20467,N_19951,N_20240);
nand U20468 (N_20468,N_20121,N_19536);
and U20469 (N_20469,N_19748,N_19592);
xnor U20470 (N_20470,N_19503,N_19397);
nor U20471 (N_20471,N_20073,N_20297);
nand U20472 (N_20472,N_20323,N_19492);
or U20473 (N_20473,N_19409,N_19410);
nand U20474 (N_20474,N_20279,N_19867);
xor U20475 (N_20475,N_19559,N_20046);
or U20476 (N_20476,N_19391,N_19267);
or U20477 (N_20477,N_20317,N_19898);
and U20478 (N_20478,N_19516,N_20245);
nor U20479 (N_20479,N_19641,N_19444);
nor U20480 (N_20480,N_19833,N_19374);
xnor U20481 (N_20481,N_19601,N_19928);
xor U20482 (N_20482,N_20115,N_20213);
and U20483 (N_20483,N_19323,N_20127);
or U20484 (N_20484,N_20251,N_19479);
xor U20485 (N_20485,N_19680,N_20005);
nor U20486 (N_20486,N_20391,N_19414);
nor U20487 (N_20487,N_19593,N_20295);
or U20488 (N_20488,N_20238,N_19956);
xor U20489 (N_20489,N_19241,N_19849);
xor U20490 (N_20490,N_19487,N_19642);
and U20491 (N_20491,N_20131,N_20079);
and U20492 (N_20492,N_20176,N_19478);
nor U20493 (N_20493,N_19330,N_20399);
xor U20494 (N_20494,N_19706,N_19715);
nand U20495 (N_20495,N_19440,N_19343);
or U20496 (N_20496,N_20222,N_20093);
nor U20497 (N_20497,N_20029,N_19383);
or U20498 (N_20498,N_19311,N_19278);
and U20499 (N_20499,N_19978,N_20202);
nor U20500 (N_20500,N_19863,N_19513);
nand U20501 (N_20501,N_20282,N_19344);
nor U20502 (N_20502,N_19967,N_19254);
nor U20503 (N_20503,N_19654,N_20358);
or U20504 (N_20504,N_19905,N_19422);
nand U20505 (N_20505,N_19845,N_20272);
or U20506 (N_20506,N_19259,N_19988);
xor U20507 (N_20507,N_19285,N_19392);
nand U20508 (N_20508,N_19345,N_20075);
and U20509 (N_20509,N_20033,N_20002);
xor U20510 (N_20510,N_19412,N_19666);
nor U20511 (N_20511,N_19304,N_20034);
or U20512 (N_20512,N_19655,N_19589);
nand U20513 (N_20513,N_19858,N_19844);
xnor U20514 (N_20514,N_19608,N_20040);
nor U20515 (N_20515,N_19827,N_19326);
xor U20516 (N_20516,N_20366,N_20292);
or U20517 (N_20517,N_19631,N_20161);
or U20518 (N_20518,N_20004,N_19812);
or U20519 (N_20519,N_19295,N_19226);
and U20520 (N_20520,N_19333,N_19723);
and U20521 (N_20521,N_19585,N_19810);
and U20522 (N_20522,N_20165,N_20277);
xor U20523 (N_20523,N_19329,N_20225);
or U20524 (N_20524,N_19566,N_19334);
or U20525 (N_20525,N_19900,N_19711);
or U20526 (N_20526,N_19404,N_19302);
xnor U20527 (N_20527,N_19544,N_20132);
xor U20528 (N_20528,N_19338,N_19450);
nor U20529 (N_20529,N_19651,N_19971);
nand U20530 (N_20530,N_20061,N_19870);
and U20531 (N_20531,N_20268,N_19673);
and U20532 (N_20532,N_19387,N_19700);
and U20533 (N_20533,N_20120,N_19568);
xor U20534 (N_20534,N_19411,N_19914);
and U20535 (N_20535,N_20101,N_19483);
xnor U20536 (N_20536,N_20084,N_19742);
xor U20537 (N_20537,N_19699,N_20283);
or U20538 (N_20538,N_19848,N_20339);
nand U20539 (N_20539,N_20000,N_19462);
nand U20540 (N_20540,N_19674,N_20293);
or U20541 (N_20541,N_19678,N_19712);
nor U20542 (N_20542,N_19736,N_19485);
and U20543 (N_20543,N_19515,N_20068);
xor U20544 (N_20544,N_19842,N_20373);
xnor U20545 (N_20545,N_19688,N_19526);
nand U20546 (N_20546,N_19299,N_19913);
nor U20547 (N_20547,N_19964,N_20010);
xor U20548 (N_20548,N_19361,N_20374);
or U20549 (N_20549,N_19888,N_19771);
and U20550 (N_20550,N_19415,N_20327);
and U20551 (N_20551,N_20192,N_20218);
nand U20552 (N_20552,N_19290,N_19318);
nand U20553 (N_20553,N_19449,N_20355);
nand U20554 (N_20554,N_20043,N_19704);
nor U20555 (N_20555,N_19283,N_19274);
nand U20556 (N_20556,N_19755,N_20110);
or U20557 (N_20557,N_20332,N_20001);
xnor U20558 (N_20558,N_20356,N_19271);
xor U20559 (N_20559,N_19997,N_19626);
and U20560 (N_20560,N_19684,N_20064);
and U20561 (N_20561,N_20349,N_19740);
or U20562 (N_20562,N_19791,N_19737);
nand U20563 (N_20563,N_20095,N_20168);
nor U20564 (N_20564,N_20148,N_20387);
xnor U20565 (N_20565,N_20269,N_20122);
xor U20566 (N_20566,N_19857,N_19960);
or U20567 (N_20567,N_19769,N_19705);
nor U20568 (N_20568,N_19583,N_20230);
xnor U20569 (N_20569,N_19256,N_19669);
xnor U20570 (N_20570,N_19886,N_19881);
or U20571 (N_20571,N_19525,N_19795);
or U20572 (N_20572,N_19488,N_19604);
or U20573 (N_20573,N_20157,N_19765);
or U20574 (N_20574,N_19407,N_20343);
and U20575 (N_20575,N_19621,N_20186);
and U20576 (N_20576,N_19883,N_19528);
and U20577 (N_20577,N_20128,N_19839);
xor U20578 (N_20578,N_19918,N_20049);
and U20579 (N_20579,N_19393,N_19339);
or U20580 (N_20580,N_19720,N_19385);
and U20581 (N_20581,N_19911,N_20164);
nand U20582 (N_20582,N_19640,N_19425);
and U20583 (N_20583,N_19661,N_20299);
xnor U20584 (N_20584,N_20051,N_19441);
nand U20585 (N_20585,N_19486,N_19524);
or U20586 (N_20586,N_20304,N_19701);
xnor U20587 (N_20587,N_19380,N_19686);
or U20588 (N_20588,N_20175,N_19829);
and U20589 (N_20589,N_19983,N_19451);
nor U20590 (N_20590,N_19327,N_19588);
nor U20591 (N_20591,N_20233,N_19709);
and U20592 (N_20592,N_19298,N_19657);
and U20593 (N_20593,N_20057,N_20309);
nand U20594 (N_20594,N_19501,N_19885);
nor U20595 (N_20595,N_20007,N_19576);
nor U20596 (N_20596,N_19434,N_20203);
or U20597 (N_20597,N_20294,N_19797);
nor U20598 (N_20598,N_19581,N_20071);
xnor U20599 (N_20599,N_19252,N_19416);
nor U20600 (N_20600,N_19580,N_20146);
nor U20601 (N_20601,N_20050,N_19300);
and U20602 (N_20602,N_20156,N_19873);
nand U20603 (N_20603,N_20276,N_20273);
and U20604 (N_20604,N_20386,N_19465);
nor U20605 (N_20605,N_19838,N_20184);
nand U20606 (N_20606,N_19619,N_19371);
or U20607 (N_20607,N_19616,N_20172);
and U20608 (N_20608,N_19780,N_20085);
xnor U20609 (N_20609,N_19468,N_20094);
xnor U20610 (N_20610,N_20060,N_19445);
nand U20611 (N_20611,N_19985,N_19325);
and U20612 (N_20612,N_19575,N_20394);
xor U20613 (N_20613,N_19622,N_20280);
nand U20614 (N_20614,N_19752,N_19799);
xnor U20615 (N_20615,N_20378,N_20341);
or U20616 (N_20616,N_19716,N_19442);
nand U20617 (N_20617,N_20285,N_19896);
or U20618 (N_20618,N_19332,N_19211);
and U20619 (N_20619,N_20392,N_19813);
xnor U20620 (N_20620,N_20258,N_20182);
nor U20621 (N_20621,N_19618,N_19980);
and U20622 (N_20622,N_20228,N_19498);
and U20623 (N_20623,N_19933,N_19237);
and U20624 (N_20624,N_19825,N_20211);
and U20625 (N_20625,N_20194,N_20016);
nand U20626 (N_20626,N_20144,N_19824);
nand U20627 (N_20627,N_19890,N_19428);
or U20628 (N_20628,N_19993,N_19724);
nor U20629 (N_20629,N_19246,N_19987);
nor U20630 (N_20630,N_20369,N_19861);
and U20631 (N_20631,N_19969,N_19400);
or U20632 (N_20632,N_20263,N_20133);
or U20633 (N_20633,N_20106,N_19770);
or U20634 (N_20634,N_20188,N_19574);
xnor U20635 (N_20635,N_20344,N_19805);
nor U20636 (N_20636,N_19243,N_20325);
and U20637 (N_20637,N_19656,N_19820);
nand U20638 (N_20638,N_20284,N_19731);
xnor U20639 (N_20639,N_20003,N_20027);
nand U20640 (N_20640,N_19745,N_19864);
and U20641 (N_20641,N_19281,N_19836);
or U20642 (N_20642,N_19965,N_20367);
nor U20643 (N_20643,N_20191,N_20045);
or U20644 (N_20644,N_19926,N_19860);
or U20645 (N_20645,N_19250,N_19433);
nor U20646 (N_20646,N_19419,N_19275);
or U20647 (N_20647,N_19767,N_19981);
or U20648 (N_20648,N_19892,N_19600);
xnor U20649 (N_20649,N_19373,N_19787);
nor U20650 (N_20650,N_20154,N_19207);
xnor U20651 (N_20651,N_19837,N_19282);
or U20652 (N_20652,N_19693,N_19895);
xnor U20653 (N_20653,N_19718,N_19349);
nor U20654 (N_20654,N_19801,N_20150);
xnor U20655 (N_20655,N_19201,N_20056);
or U20656 (N_20656,N_19263,N_20178);
xnor U20657 (N_20657,N_20236,N_19530);
or U20658 (N_20658,N_20055,N_20052);
or U20659 (N_20659,N_19365,N_19248);
or U20660 (N_20660,N_19871,N_20187);
nand U20661 (N_20661,N_19453,N_19903);
and U20662 (N_20662,N_19491,N_19710);
nand U20663 (N_20663,N_20090,N_19303);
and U20664 (N_20664,N_19473,N_19310);
nand U20665 (N_20665,N_19443,N_20103);
nor U20666 (N_20666,N_19800,N_20171);
xor U20667 (N_20667,N_19814,N_20063);
xnor U20668 (N_20668,N_19775,N_19719);
nor U20669 (N_20669,N_20153,N_20205);
nor U20670 (N_20670,N_19308,N_19937);
nor U20671 (N_20671,N_20239,N_19542);
nand U20672 (N_20672,N_19675,N_20313);
and U20673 (N_20673,N_20062,N_19999);
nor U20674 (N_20674,N_20318,N_19435);
nand U20675 (N_20675,N_19596,N_20340);
nor U20676 (N_20676,N_20006,N_19691);
nand U20677 (N_20677,N_20143,N_19766);
nand U20678 (N_20678,N_20360,N_19552);
nand U20679 (N_20679,N_20179,N_20217);
nand U20680 (N_20680,N_20174,N_20013);
nor U20681 (N_20681,N_19816,N_19307);
nand U20682 (N_20682,N_19603,N_19645);
nand U20683 (N_20683,N_19776,N_19590);
nor U20684 (N_20684,N_19729,N_20296);
nand U20685 (N_20685,N_20350,N_19511);
nand U20686 (N_20686,N_19240,N_20031);
nor U20687 (N_20687,N_19222,N_19851);
nor U20688 (N_20688,N_19901,N_19502);
nor U20689 (N_20689,N_19354,N_20253);
xor U20690 (N_20690,N_19471,N_20232);
and U20691 (N_20691,N_19551,N_19741);
xnor U20692 (N_20692,N_20030,N_19208);
nor U20693 (N_20693,N_19467,N_20382);
xnor U20694 (N_20694,N_19634,N_19247);
nor U20695 (N_20695,N_19624,N_20346);
nor U20696 (N_20696,N_20116,N_19322);
or U20697 (N_20697,N_19555,N_19689);
xnor U20698 (N_20698,N_19907,N_20066);
nor U20699 (N_20699,N_19782,N_20199);
nand U20700 (N_20700,N_20302,N_19714);
nor U20701 (N_20701,N_19341,N_19629);
nor U20702 (N_20702,N_19792,N_19878);
or U20703 (N_20703,N_19620,N_19309);
xor U20704 (N_20704,N_20300,N_19696);
nor U20705 (N_20705,N_20330,N_19431);
nor U20706 (N_20706,N_20397,N_20237);
or U20707 (N_20707,N_19586,N_20196);
nor U20708 (N_20708,N_19943,N_19337);
xor U20709 (N_20709,N_20022,N_19916);
nand U20710 (N_20710,N_19335,N_20097);
nand U20711 (N_20711,N_19963,N_20091);
nand U20712 (N_20712,N_19959,N_19582);
nand U20713 (N_20713,N_20089,N_19457);
and U20714 (N_20714,N_19947,N_20114);
or U20715 (N_20715,N_19768,N_19268);
or U20716 (N_20716,N_20320,N_19667);
xnor U20717 (N_20717,N_19520,N_19938);
xor U20718 (N_20718,N_19632,N_19594);
and U20719 (N_20719,N_19286,N_19474);
or U20720 (N_20720,N_19977,N_20190);
xnor U20721 (N_20721,N_19612,N_19784);
nand U20722 (N_20722,N_19876,N_19521);
or U20723 (N_20723,N_20047,N_19508);
or U20724 (N_20724,N_19637,N_20076);
or U20725 (N_20725,N_19868,N_19966);
nand U20726 (N_20726,N_19872,N_19973);
nand U20727 (N_20727,N_19908,N_19683);
nand U20728 (N_20728,N_19227,N_19230);
or U20729 (N_20729,N_20201,N_19390);
xor U20730 (N_20730,N_19454,N_19989);
and U20731 (N_20731,N_19972,N_19257);
or U20732 (N_20732,N_19996,N_19889);
xnor U20733 (N_20733,N_19360,N_20117);
nor U20734 (N_20734,N_19615,N_19950);
or U20735 (N_20735,N_19423,N_20275);
nand U20736 (N_20736,N_20363,N_19613);
nor U20737 (N_20737,N_19238,N_20324);
nand U20738 (N_20738,N_19984,N_19426);
xor U20739 (N_20739,N_19672,N_19954);
xor U20740 (N_20740,N_20138,N_20384);
nor U20741 (N_20741,N_20107,N_20331);
and U20742 (N_20742,N_20354,N_19370);
or U20743 (N_20743,N_19377,N_19224);
nand U20744 (N_20744,N_20151,N_19461);
xor U20745 (N_20745,N_20096,N_19319);
or U20746 (N_20746,N_19527,N_19902);
nand U20747 (N_20747,N_19785,N_19293);
or U20748 (N_20748,N_20347,N_19569);
nor U20749 (N_20749,N_20170,N_20026);
and U20750 (N_20750,N_19563,N_20019);
and U20751 (N_20751,N_20044,N_20376);
or U20752 (N_20752,N_19315,N_20353);
nand U20753 (N_20753,N_20177,N_19272);
and U20754 (N_20754,N_19579,N_19728);
nand U20755 (N_20755,N_20267,N_19200);
nand U20756 (N_20756,N_19291,N_19940);
nand U20757 (N_20757,N_20388,N_19424);
nand U20758 (N_20758,N_19212,N_20305);
or U20759 (N_20759,N_20053,N_19694);
xor U20760 (N_20760,N_20359,N_19475);
nand U20761 (N_20761,N_20080,N_19269);
or U20762 (N_20762,N_19430,N_20334);
nor U20763 (N_20763,N_19570,N_19504);
nand U20764 (N_20764,N_19549,N_20223);
nand U20765 (N_20765,N_20104,N_19231);
nand U20766 (N_20766,N_19577,N_19650);
or U20767 (N_20767,N_19413,N_19942);
xor U20768 (N_20768,N_19764,N_20287);
nand U20769 (N_20769,N_19595,N_19671);
nand U20770 (N_20770,N_19297,N_20259);
nand U20771 (N_20771,N_19519,N_20333);
nor U20772 (N_20772,N_19636,N_19841);
nor U20773 (N_20773,N_19685,N_19677);
and U20774 (N_20774,N_19261,N_20242);
or U20775 (N_20775,N_19662,N_20159);
and U20776 (N_20776,N_19879,N_19292);
or U20777 (N_20777,N_19558,N_19472);
or U20778 (N_20778,N_20204,N_19301);
or U20779 (N_20779,N_19437,N_19253);
nor U20780 (N_20780,N_20385,N_19762);
and U20781 (N_20781,N_19692,N_19834);
nor U20782 (N_20782,N_19952,N_19264);
xor U20783 (N_20783,N_19774,N_19815);
xnor U20784 (N_20784,N_19893,N_19314);
nor U20785 (N_20785,N_19346,N_19783);
and U20786 (N_20786,N_19244,N_19277);
and U20787 (N_20787,N_20009,N_20262);
xnor U20788 (N_20788,N_19713,N_19490);
and U20789 (N_20789,N_19539,N_20244);
nor U20790 (N_20790,N_20113,N_19548);
nand U20791 (N_20791,N_19643,N_19934);
or U20792 (N_20792,N_19353,N_19817);
nand U20793 (N_20793,N_19609,N_19245);
or U20794 (N_20794,N_20070,N_19818);
or U20795 (N_20795,N_19979,N_19853);
nand U20796 (N_20796,N_19939,N_19702);
and U20797 (N_20797,N_19658,N_19202);
nor U20798 (N_20798,N_19732,N_19217);
nand U20799 (N_20799,N_20198,N_19545);
and U20800 (N_20800,N_19777,N_19955);
xnor U20801 (N_20801,N_19584,N_20083);
nor U20802 (N_20802,N_20357,N_19289);
nand U20803 (N_20803,N_19739,N_20059);
xor U20804 (N_20804,N_20099,N_20207);
or U20805 (N_20805,N_19668,N_19529);
nor U20806 (N_20806,N_20288,N_19352);
or U20807 (N_20807,N_19986,N_19210);
xor U20808 (N_20808,N_19320,N_19543);
or U20809 (N_20809,N_19925,N_19929);
xor U20810 (N_20810,N_20037,N_20261);
nand U20811 (N_20811,N_19533,N_20185);
nor U20812 (N_20812,N_19229,N_19363);
xor U20813 (N_20813,N_19953,N_20125);
or U20814 (N_20814,N_20286,N_20112);
nand U20815 (N_20815,N_19627,N_20224);
and U20816 (N_20816,N_19750,N_19945);
xnor U20817 (N_20817,N_19875,N_20119);
nand U20818 (N_20818,N_20379,N_19793);
nand U20819 (N_20819,N_20169,N_19681);
and U20820 (N_20820,N_20124,N_19846);
nor U20821 (N_20821,N_20345,N_20337);
and U20822 (N_20822,N_20260,N_20227);
nand U20823 (N_20823,N_19233,N_20072);
nor U20824 (N_20824,N_20241,N_19910);
and U20825 (N_20825,N_20235,N_19518);
xor U20826 (N_20826,N_19206,N_19540);
nand U20827 (N_20827,N_19439,N_20152);
and U20828 (N_20828,N_20291,N_19663);
or U20829 (N_20829,N_19831,N_19223);
xor U20830 (N_20830,N_19994,N_20377);
and U20831 (N_20831,N_19819,N_20321);
nor U20832 (N_20832,N_19381,N_19804);
and U20833 (N_20833,N_20221,N_19553);
nor U20834 (N_20834,N_19990,N_20197);
nand U20835 (N_20835,N_19664,N_20271);
xor U20836 (N_20836,N_19847,N_19567);
nand U20837 (N_20837,N_19305,N_19556);
or U20838 (N_20838,N_20342,N_19941);
or U20839 (N_20839,N_20234,N_19510);
nor U20840 (N_20840,N_19294,N_20248);
nand U20841 (N_20841,N_19427,N_19982);
or U20842 (N_20842,N_19496,N_19830);
or U20843 (N_20843,N_20256,N_20351);
nand U20844 (N_20844,N_20088,N_20336);
and U20845 (N_20845,N_19564,N_19296);
xor U20846 (N_20846,N_19708,N_19855);
or U20847 (N_20847,N_19276,N_19366);
nand U20848 (N_20848,N_19707,N_19362);
and U20849 (N_20849,N_19946,N_19265);
nor U20850 (N_20850,N_19808,N_20067);
xor U20851 (N_20851,N_19359,N_19690);
nor U20852 (N_20852,N_19280,N_19561);
nor U20853 (N_20853,N_19573,N_19219);
xor U20854 (N_20854,N_19284,N_20231);
or U20855 (N_20855,N_19610,N_20390);
xor U20856 (N_20856,N_19931,N_19288);
nand U20857 (N_20857,N_19336,N_19866);
and U20858 (N_20858,N_19930,N_19456);
xor U20859 (N_20859,N_19218,N_20329);
xor U20860 (N_20860,N_20118,N_19957);
nor U20861 (N_20861,N_19697,N_19406);
or U20862 (N_20862,N_19968,N_19497);
nor U20863 (N_20863,N_19214,N_20326);
xnor U20864 (N_20864,N_20335,N_19324);
xor U20865 (N_20865,N_19372,N_19398);
and U20866 (N_20866,N_19646,N_19408);
and U20867 (N_20867,N_19375,N_19507);
nand U20868 (N_20868,N_19260,N_20298);
nor U20869 (N_20869,N_19499,N_20361);
or U20870 (N_20870,N_19578,N_20158);
nand U20871 (N_20871,N_20042,N_19287);
and U20872 (N_20872,N_20041,N_19682);
and U20873 (N_20873,N_19856,N_20348);
nand U20874 (N_20874,N_20140,N_20229);
or U20875 (N_20875,N_19379,N_19727);
nand U20876 (N_20876,N_19348,N_19448);
nor U20877 (N_20877,N_20311,N_19840);
or U20878 (N_20878,N_19466,N_20077);
and U20879 (N_20879,N_20254,N_19607);
nor U20880 (N_20880,N_19828,N_20108);
or U20881 (N_20881,N_20039,N_19446);
or U20882 (N_20882,N_19403,N_19721);
nand U20883 (N_20883,N_19687,N_20036);
xnor U20884 (N_20884,N_20389,N_19639);
or U20885 (N_20885,N_19962,N_20074);
xnor U20886 (N_20886,N_20365,N_19617);
or U20887 (N_20887,N_20257,N_19321);
nor U20888 (N_20888,N_20193,N_19882);
nor U20889 (N_20889,N_19730,N_19949);
xor U20890 (N_20890,N_19306,N_20180);
nor U20891 (N_20891,N_20102,N_19751);
xor U20892 (N_20892,N_20100,N_20032);
and U20893 (N_20893,N_19399,N_19602);
nor U20894 (N_20894,N_20065,N_20210);
and U20895 (N_20895,N_19482,N_19347);
or U20896 (N_20896,N_19251,N_19452);
or U20897 (N_20897,N_19823,N_20206);
and U20898 (N_20898,N_19635,N_20214);
and U20899 (N_20899,N_19358,N_19517);
xor U20900 (N_20900,N_20281,N_19733);
nand U20901 (N_20901,N_19625,N_19376);
nor U20902 (N_20902,N_20142,N_20301);
and U20903 (N_20903,N_19746,N_19912);
xnor U20904 (N_20904,N_19328,N_19384);
xor U20905 (N_20905,N_19364,N_19395);
nand U20906 (N_20906,N_19779,N_19228);
xor U20907 (N_20907,N_20069,N_19630);
nand U20908 (N_20908,N_19899,N_19547);
nor U20909 (N_20909,N_19923,N_20011);
or U20910 (N_20910,N_19262,N_19778);
nand U20911 (N_20911,N_19803,N_20398);
nand U20912 (N_20912,N_20145,N_19919);
xor U20913 (N_20913,N_19484,N_20105);
xor U20914 (N_20914,N_19464,N_19235);
nand U20915 (N_20915,N_19599,N_19494);
nor U20916 (N_20916,N_19481,N_19915);
nand U20917 (N_20917,N_19405,N_19796);
xor U20918 (N_20918,N_20149,N_19255);
and U20919 (N_20919,N_19606,N_20078);
nor U20920 (N_20920,N_20173,N_19725);
nand U20921 (N_20921,N_20364,N_19644);
nand U20922 (N_20922,N_20264,N_20058);
and U20923 (N_20923,N_20136,N_20189);
and U20924 (N_20924,N_20266,N_19532);
nand U20925 (N_20925,N_19649,N_19557);
and U20926 (N_20926,N_19506,N_19204);
and U20927 (N_20927,N_19747,N_19922);
nand U20928 (N_20928,N_19897,N_19550);
nor U20929 (N_20929,N_19743,N_19659);
or U20930 (N_20930,N_19653,N_19537);
or U20931 (N_20931,N_19500,N_19754);
nand U20932 (N_20932,N_19489,N_19974);
or U20933 (N_20933,N_20134,N_19401);
and U20934 (N_20934,N_19611,N_20289);
and U20935 (N_20935,N_19572,N_19772);
nand U20936 (N_20936,N_19676,N_20038);
nor U20937 (N_20937,N_19538,N_19480);
nor U20938 (N_20938,N_20371,N_19614);
and U20939 (N_20939,N_19469,N_20109);
nand U20940 (N_20940,N_20308,N_20352);
xor U20941 (N_20941,N_19215,N_19421);
xnor U20942 (N_20942,N_20290,N_19531);
and U20943 (N_20943,N_20048,N_19927);
xor U20944 (N_20944,N_20315,N_19470);
and U20945 (N_20945,N_19961,N_20166);
and U20946 (N_20946,N_19598,N_19509);
nand U20947 (N_20947,N_19975,N_20020);
xor U20948 (N_20948,N_19936,N_20274);
xnor U20949 (N_20949,N_19591,N_20265);
nand U20950 (N_20950,N_19852,N_20123);
xnor U20951 (N_20951,N_20160,N_20183);
nor U20952 (N_20952,N_19992,N_20023);
nor U20953 (N_20953,N_20380,N_19906);
xor U20954 (N_20954,N_19909,N_20215);
nor U20955 (N_20955,N_19270,N_20155);
and U20956 (N_20956,N_19821,N_19571);
or U20957 (N_20957,N_20054,N_19316);
and U20958 (N_20958,N_19648,N_20208);
and U20959 (N_20959,N_19862,N_19832);
nor U20960 (N_20960,N_20111,N_20314);
xor U20961 (N_20961,N_19826,N_19209);
and U20962 (N_20962,N_19735,N_19396);
nor U20963 (N_20963,N_20086,N_19647);
and U20964 (N_20964,N_20216,N_19802);
xnor U20965 (N_20965,N_19438,N_19759);
nand U20966 (N_20966,N_19891,N_19695);
and U20967 (N_20967,N_19660,N_20219);
xor U20968 (N_20968,N_20226,N_20255);
nand U20969 (N_20969,N_19258,N_19894);
and U20970 (N_20970,N_20249,N_19744);
nor U20971 (N_20971,N_19717,N_20328);
or U20972 (N_20972,N_20024,N_19417);
nor U20973 (N_20973,N_19726,N_20087);
and U20974 (N_20974,N_19843,N_19944);
and U20975 (N_20975,N_19628,N_20035);
nand U20976 (N_20976,N_19394,N_19605);
nand U20977 (N_20977,N_19734,N_19368);
nand U20978 (N_20978,N_19378,N_20008);
xnor U20979 (N_20979,N_19505,N_19761);
xor U20980 (N_20980,N_19679,N_19203);
nor U20981 (N_20981,N_20270,N_19216);
and U20982 (N_20982,N_19514,N_19998);
or U20983 (N_20983,N_19493,N_19458);
xor U20984 (N_20984,N_19420,N_19794);
or U20985 (N_20985,N_20395,N_19788);
nor U20986 (N_20986,N_20129,N_19357);
xnor U20987 (N_20987,N_20306,N_19367);
nor U20988 (N_20988,N_19703,N_19418);
and U20989 (N_20989,N_19560,N_20098);
nand U20990 (N_20990,N_19738,N_19869);
and U20991 (N_20991,N_19279,N_19356);
or U20992 (N_20992,N_19786,N_20141);
or U20993 (N_20993,N_20252,N_19436);
or U20994 (N_20994,N_20362,N_20195);
and U20995 (N_20995,N_20162,N_20014);
and U20996 (N_20996,N_19273,N_19835);
xnor U20997 (N_20997,N_19790,N_19432);
or U20998 (N_20998,N_19756,N_19389);
or U20999 (N_20999,N_20375,N_19351);
nor U21000 (N_21000,N_19931,N_20135);
nor U21001 (N_21001,N_19317,N_19725);
or U21002 (N_21002,N_19739,N_19634);
nand U21003 (N_21003,N_20131,N_19915);
nor U21004 (N_21004,N_20239,N_19525);
or U21005 (N_21005,N_19910,N_20185);
and U21006 (N_21006,N_19217,N_19370);
or U21007 (N_21007,N_19326,N_19513);
nand U21008 (N_21008,N_19574,N_19644);
nand U21009 (N_21009,N_19308,N_20374);
xor U21010 (N_21010,N_20027,N_20356);
or U21011 (N_21011,N_20082,N_19376);
nor U21012 (N_21012,N_19664,N_19588);
or U21013 (N_21013,N_19744,N_20255);
and U21014 (N_21014,N_19910,N_20079);
or U21015 (N_21015,N_20038,N_20113);
nand U21016 (N_21016,N_19270,N_19951);
nand U21017 (N_21017,N_19352,N_20150);
nor U21018 (N_21018,N_19425,N_19775);
xnor U21019 (N_21019,N_19761,N_20036);
or U21020 (N_21020,N_19583,N_20014);
and U21021 (N_21021,N_20315,N_20010);
xor U21022 (N_21022,N_20078,N_19471);
nand U21023 (N_21023,N_20229,N_19872);
nor U21024 (N_21024,N_20116,N_20031);
or U21025 (N_21025,N_20015,N_19211);
nor U21026 (N_21026,N_20387,N_19707);
xnor U21027 (N_21027,N_19327,N_19420);
or U21028 (N_21028,N_20375,N_20041);
nand U21029 (N_21029,N_20070,N_19495);
and U21030 (N_21030,N_20048,N_19716);
xor U21031 (N_21031,N_20059,N_19425);
nor U21032 (N_21032,N_19716,N_19295);
or U21033 (N_21033,N_19288,N_19334);
nand U21034 (N_21034,N_19609,N_19983);
nand U21035 (N_21035,N_19227,N_19941);
or U21036 (N_21036,N_19313,N_20092);
nor U21037 (N_21037,N_19602,N_19766);
or U21038 (N_21038,N_19969,N_20323);
nand U21039 (N_21039,N_20394,N_20296);
or U21040 (N_21040,N_19682,N_19701);
or U21041 (N_21041,N_19864,N_19292);
nor U21042 (N_21042,N_19465,N_19572);
or U21043 (N_21043,N_20084,N_20305);
or U21044 (N_21044,N_20061,N_19827);
or U21045 (N_21045,N_19575,N_20312);
or U21046 (N_21046,N_20330,N_20050);
nand U21047 (N_21047,N_20344,N_19208);
and U21048 (N_21048,N_19367,N_19691);
nand U21049 (N_21049,N_19351,N_19620);
xor U21050 (N_21050,N_19545,N_20323);
or U21051 (N_21051,N_19431,N_20257);
or U21052 (N_21052,N_20323,N_19857);
and U21053 (N_21053,N_19675,N_19907);
nor U21054 (N_21054,N_20333,N_20366);
xor U21055 (N_21055,N_19294,N_19224);
and U21056 (N_21056,N_19826,N_19726);
xnor U21057 (N_21057,N_20027,N_19523);
and U21058 (N_21058,N_20333,N_19812);
xor U21059 (N_21059,N_19770,N_20274);
or U21060 (N_21060,N_19651,N_19594);
nor U21061 (N_21061,N_20059,N_19429);
xor U21062 (N_21062,N_19489,N_20364);
nor U21063 (N_21063,N_19977,N_19772);
nor U21064 (N_21064,N_19282,N_19343);
or U21065 (N_21065,N_20337,N_20301);
nand U21066 (N_21066,N_19639,N_20123);
nor U21067 (N_21067,N_20338,N_19317);
nor U21068 (N_21068,N_19702,N_19309);
nor U21069 (N_21069,N_19445,N_20350);
nand U21070 (N_21070,N_19880,N_19512);
xor U21071 (N_21071,N_20338,N_19766);
nor U21072 (N_21072,N_20017,N_19341);
or U21073 (N_21073,N_19538,N_19481);
nand U21074 (N_21074,N_19510,N_19839);
nand U21075 (N_21075,N_19374,N_20233);
xor U21076 (N_21076,N_19411,N_19587);
and U21077 (N_21077,N_19400,N_19915);
nor U21078 (N_21078,N_20029,N_20392);
or U21079 (N_21079,N_19961,N_19744);
xor U21080 (N_21080,N_20039,N_20321);
or U21081 (N_21081,N_19304,N_19350);
and U21082 (N_21082,N_19305,N_20014);
nor U21083 (N_21083,N_19476,N_20030);
nor U21084 (N_21084,N_19915,N_19991);
xnor U21085 (N_21085,N_19326,N_19366);
and U21086 (N_21086,N_20212,N_19485);
nor U21087 (N_21087,N_19770,N_19569);
nor U21088 (N_21088,N_20080,N_20055);
xnor U21089 (N_21089,N_20213,N_19592);
xnor U21090 (N_21090,N_19319,N_19984);
xor U21091 (N_21091,N_19640,N_20381);
or U21092 (N_21092,N_19892,N_19507);
or U21093 (N_21093,N_19418,N_20127);
nand U21094 (N_21094,N_19617,N_19680);
xor U21095 (N_21095,N_19434,N_19465);
or U21096 (N_21096,N_19615,N_20366);
or U21097 (N_21097,N_20375,N_20063);
xnor U21098 (N_21098,N_20128,N_19410);
nand U21099 (N_21099,N_19876,N_20174);
xor U21100 (N_21100,N_19772,N_20006);
nor U21101 (N_21101,N_20015,N_19658);
xor U21102 (N_21102,N_19871,N_20334);
nand U21103 (N_21103,N_19326,N_19761);
xor U21104 (N_21104,N_19356,N_20272);
or U21105 (N_21105,N_19267,N_19883);
xor U21106 (N_21106,N_19533,N_19402);
or U21107 (N_21107,N_19496,N_19224);
nor U21108 (N_21108,N_20348,N_19928);
nor U21109 (N_21109,N_20065,N_19940);
nor U21110 (N_21110,N_19515,N_20308);
nand U21111 (N_21111,N_20380,N_19943);
nor U21112 (N_21112,N_19371,N_19848);
or U21113 (N_21113,N_20375,N_19202);
and U21114 (N_21114,N_19690,N_20065);
and U21115 (N_21115,N_19747,N_19425);
and U21116 (N_21116,N_20051,N_19512);
nor U21117 (N_21117,N_19350,N_20059);
nand U21118 (N_21118,N_19700,N_19686);
nand U21119 (N_21119,N_20198,N_20338);
and U21120 (N_21120,N_19514,N_20296);
nor U21121 (N_21121,N_20361,N_20023);
and U21122 (N_21122,N_19917,N_19961);
nand U21123 (N_21123,N_19640,N_20240);
xnor U21124 (N_21124,N_20063,N_19953);
nand U21125 (N_21125,N_19242,N_19698);
and U21126 (N_21126,N_19409,N_19764);
nor U21127 (N_21127,N_19924,N_19551);
and U21128 (N_21128,N_20043,N_20297);
nand U21129 (N_21129,N_19401,N_20098);
xnor U21130 (N_21130,N_19357,N_19886);
or U21131 (N_21131,N_19617,N_19368);
xor U21132 (N_21132,N_19777,N_20151);
or U21133 (N_21133,N_19845,N_20336);
nand U21134 (N_21134,N_20215,N_19379);
nor U21135 (N_21135,N_19846,N_19558);
nand U21136 (N_21136,N_20057,N_19775);
and U21137 (N_21137,N_19265,N_19969);
nand U21138 (N_21138,N_19351,N_20310);
and U21139 (N_21139,N_20249,N_19748);
xor U21140 (N_21140,N_20149,N_19534);
nand U21141 (N_21141,N_20223,N_19760);
xnor U21142 (N_21142,N_19226,N_20100);
xor U21143 (N_21143,N_19403,N_19916);
nor U21144 (N_21144,N_19471,N_19547);
nor U21145 (N_21145,N_19785,N_19724);
or U21146 (N_21146,N_19640,N_19242);
xor U21147 (N_21147,N_19595,N_20105);
xnor U21148 (N_21148,N_19782,N_19722);
and U21149 (N_21149,N_19762,N_19350);
and U21150 (N_21150,N_19747,N_19262);
nand U21151 (N_21151,N_19549,N_19823);
nand U21152 (N_21152,N_19411,N_20394);
and U21153 (N_21153,N_20054,N_19307);
xnor U21154 (N_21154,N_19699,N_20010);
nand U21155 (N_21155,N_20395,N_19955);
or U21156 (N_21156,N_19405,N_19294);
and U21157 (N_21157,N_19736,N_19438);
nor U21158 (N_21158,N_19634,N_19415);
or U21159 (N_21159,N_20178,N_19858);
and U21160 (N_21160,N_20328,N_19370);
xor U21161 (N_21161,N_19883,N_20129);
xor U21162 (N_21162,N_19964,N_19989);
nor U21163 (N_21163,N_19228,N_19516);
nand U21164 (N_21164,N_19942,N_20116);
or U21165 (N_21165,N_19568,N_19655);
or U21166 (N_21166,N_19701,N_19977);
nand U21167 (N_21167,N_19853,N_19239);
and U21168 (N_21168,N_19250,N_19598);
or U21169 (N_21169,N_19483,N_19811);
xnor U21170 (N_21170,N_19311,N_20199);
xor U21171 (N_21171,N_19420,N_19413);
xnor U21172 (N_21172,N_20243,N_20022);
xor U21173 (N_21173,N_19855,N_19787);
nor U21174 (N_21174,N_19381,N_20171);
nand U21175 (N_21175,N_19231,N_19358);
xnor U21176 (N_21176,N_19900,N_20352);
or U21177 (N_21177,N_19480,N_20057);
nand U21178 (N_21178,N_19947,N_19486);
and U21179 (N_21179,N_19510,N_19454);
nand U21180 (N_21180,N_19596,N_19310);
or U21181 (N_21181,N_19554,N_19251);
xor U21182 (N_21182,N_19253,N_20161);
xor U21183 (N_21183,N_19633,N_19797);
xor U21184 (N_21184,N_19307,N_19780);
xnor U21185 (N_21185,N_19462,N_19696);
or U21186 (N_21186,N_19946,N_19378);
or U21187 (N_21187,N_19825,N_19203);
and U21188 (N_21188,N_20379,N_19794);
nor U21189 (N_21189,N_20079,N_19485);
or U21190 (N_21190,N_19256,N_19763);
and U21191 (N_21191,N_19696,N_19400);
and U21192 (N_21192,N_19298,N_19339);
nand U21193 (N_21193,N_19703,N_19599);
xnor U21194 (N_21194,N_19327,N_20225);
xnor U21195 (N_21195,N_19708,N_19375);
and U21196 (N_21196,N_20321,N_19744);
and U21197 (N_21197,N_19800,N_19360);
nand U21198 (N_21198,N_19840,N_19306);
or U21199 (N_21199,N_20361,N_20293);
or U21200 (N_21200,N_19726,N_19912);
xor U21201 (N_21201,N_19633,N_19925);
nand U21202 (N_21202,N_20130,N_20017);
nand U21203 (N_21203,N_20291,N_20302);
xnor U21204 (N_21204,N_19212,N_19348);
nand U21205 (N_21205,N_20281,N_19750);
xor U21206 (N_21206,N_20083,N_20065);
nand U21207 (N_21207,N_20174,N_20240);
nor U21208 (N_21208,N_19929,N_20089);
or U21209 (N_21209,N_19624,N_20295);
nand U21210 (N_21210,N_19594,N_20023);
nor U21211 (N_21211,N_20069,N_19493);
nand U21212 (N_21212,N_19374,N_19210);
nor U21213 (N_21213,N_19880,N_19722);
nand U21214 (N_21214,N_20245,N_19305);
and U21215 (N_21215,N_20367,N_19822);
and U21216 (N_21216,N_19730,N_19686);
xnor U21217 (N_21217,N_19775,N_19773);
and U21218 (N_21218,N_19410,N_19219);
xor U21219 (N_21219,N_19932,N_20258);
nor U21220 (N_21220,N_20104,N_19714);
and U21221 (N_21221,N_20240,N_20305);
and U21222 (N_21222,N_19532,N_19702);
or U21223 (N_21223,N_19450,N_19679);
xnor U21224 (N_21224,N_20197,N_19770);
xnor U21225 (N_21225,N_19786,N_19769);
or U21226 (N_21226,N_20208,N_19676);
and U21227 (N_21227,N_19790,N_19504);
nor U21228 (N_21228,N_20229,N_19915);
nand U21229 (N_21229,N_19489,N_20132);
nor U21230 (N_21230,N_19721,N_19720);
and U21231 (N_21231,N_19422,N_20396);
nand U21232 (N_21232,N_19993,N_19488);
xor U21233 (N_21233,N_19662,N_19516);
nor U21234 (N_21234,N_19811,N_19916);
xor U21235 (N_21235,N_19723,N_19446);
xor U21236 (N_21236,N_20244,N_20145);
nand U21237 (N_21237,N_19356,N_19237);
or U21238 (N_21238,N_19236,N_19585);
or U21239 (N_21239,N_20252,N_19848);
xor U21240 (N_21240,N_20032,N_19459);
nor U21241 (N_21241,N_20326,N_19606);
xor U21242 (N_21242,N_19453,N_20386);
nor U21243 (N_21243,N_19839,N_19278);
nand U21244 (N_21244,N_19621,N_20246);
nand U21245 (N_21245,N_19383,N_19748);
or U21246 (N_21246,N_20259,N_19636);
xnor U21247 (N_21247,N_19213,N_19532);
or U21248 (N_21248,N_20132,N_19944);
xor U21249 (N_21249,N_19726,N_19452);
xor U21250 (N_21250,N_19823,N_19746);
nor U21251 (N_21251,N_20151,N_19552);
or U21252 (N_21252,N_20145,N_19507);
or U21253 (N_21253,N_19531,N_20270);
nand U21254 (N_21254,N_19659,N_19481);
nor U21255 (N_21255,N_19848,N_19377);
xor U21256 (N_21256,N_19469,N_19735);
nor U21257 (N_21257,N_19841,N_19439);
nand U21258 (N_21258,N_20387,N_20383);
nor U21259 (N_21259,N_19698,N_19904);
xor U21260 (N_21260,N_20120,N_19415);
and U21261 (N_21261,N_19842,N_19201);
xor U21262 (N_21262,N_19508,N_19725);
nor U21263 (N_21263,N_19707,N_20231);
and U21264 (N_21264,N_19912,N_19236);
or U21265 (N_21265,N_19858,N_19768);
or U21266 (N_21266,N_19784,N_20012);
and U21267 (N_21267,N_20072,N_20370);
or U21268 (N_21268,N_19528,N_19533);
xnor U21269 (N_21269,N_20097,N_20243);
xor U21270 (N_21270,N_19977,N_19976);
xnor U21271 (N_21271,N_19646,N_20175);
xnor U21272 (N_21272,N_20121,N_20315);
nor U21273 (N_21273,N_19586,N_20067);
nand U21274 (N_21274,N_19526,N_19865);
xnor U21275 (N_21275,N_20125,N_19983);
nor U21276 (N_21276,N_19876,N_19789);
xnor U21277 (N_21277,N_19636,N_19572);
nor U21278 (N_21278,N_19976,N_20365);
nor U21279 (N_21279,N_19858,N_19583);
or U21280 (N_21280,N_20308,N_19554);
nor U21281 (N_21281,N_19211,N_19231);
xor U21282 (N_21282,N_19853,N_19710);
or U21283 (N_21283,N_20107,N_19487);
and U21284 (N_21284,N_19743,N_19720);
and U21285 (N_21285,N_20365,N_19631);
and U21286 (N_21286,N_19642,N_19634);
nor U21287 (N_21287,N_19579,N_19635);
nor U21288 (N_21288,N_19660,N_19577);
or U21289 (N_21289,N_19975,N_19428);
xor U21290 (N_21290,N_19292,N_19996);
nor U21291 (N_21291,N_20370,N_19965);
nor U21292 (N_21292,N_19772,N_19945);
and U21293 (N_21293,N_20343,N_19630);
or U21294 (N_21294,N_20054,N_19407);
or U21295 (N_21295,N_20233,N_19807);
and U21296 (N_21296,N_19611,N_19862);
or U21297 (N_21297,N_19755,N_19907);
and U21298 (N_21298,N_19823,N_19410);
nand U21299 (N_21299,N_19204,N_19606);
and U21300 (N_21300,N_20252,N_19415);
and U21301 (N_21301,N_19504,N_19430);
and U21302 (N_21302,N_19491,N_20184);
and U21303 (N_21303,N_19237,N_19403);
nor U21304 (N_21304,N_20011,N_19353);
nor U21305 (N_21305,N_19378,N_19448);
xnor U21306 (N_21306,N_19981,N_20198);
nor U21307 (N_21307,N_20324,N_19226);
or U21308 (N_21308,N_19696,N_19763);
nor U21309 (N_21309,N_19937,N_20074);
nand U21310 (N_21310,N_19585,N_19436);
nor U21311 (N_21311,N_20101,N_19302);
or U21312 (N_21312,N_19796,N_19960);
nor U21313 (N_21313,N_19495,N_20392);
and U21314 (N_21314,N_19304,N_20101);
nand U21315 (N_21315,N_20206,N_19287);
and U21316 (N_21316,N_20269,N_20169);
xnor U21317 (N_21317,N_19662,N_19587);
xnor U21318 (N_21318,N_19714,N_20289);
xor U21319 (N_21319,N_19640,N_19766);
and U21320 (N_21320,N_19824,N_19410);
xnor U21321 (N_21321,N_19352,N_19703);
or U21322 (N_21322,N_20221,N_20139);
nand U21323 (N_21323,N_20222,N_19775);
and U21324 (N_21324,N_19460,N_19837);
xor U21325 (N_21325,N_20130,N_19676);
xor U21326 (N_21326,N_19325,N_20143);
xnor U21327 (N_21327,N_19965,N_19482);
nand U21328 (N_21328,N_19233,N_19384);
or U21329 (N_21329,N_19378,N_19932);
nand U21330 (N_21330,N_19576,N_20157);
or U21331 (N_21331,N_20068,N_19879);
xor U21332 (N_21332,N_19295,N_19951);
nor U21333 (N_21333,N_19393,N_19719);
nor U21334 (N_21334,N_19714,N_19863);
or U21335 (N_21335,N_19645,N_19809);
nor U21336 (N_21336,N_19645,N_19210);
nand U21337 (N_21337,N_20260,N_20146);
and U21338 (N_21338,N_19755,N_19242);
xnor U21339 (N_21339,N_19733,N_19255);
nor U21340 (N_21340,N_20092,N_19490);
xor U21341 (N_21341,N_19812,N_19584);
xnor U21342 (N_21342,N_19380,N_19819);
or U21343 (N_21343,N_19907,N_20261);
and U21344 (N_21344,N_20281,N_19816);
nor U21345 (N_21345,N_19996,N_20035);
and U21346 (N_21346,N_19924,N_20150);
nor U21347 (N_21347,N_20138,N_19437);
nor U21348 (N_21348,N_20366,N_20194);
or U21349 (N_21349,N_19818,N_19888);
nor U21350 (N_21350,N_19639,N_20335);
nand U21351 (N_21351,N_19637,N_19772);
nand U21352 (N_21352,N_19970,N_19504);
and U21353 (N_21353,N_20156,N_19214);
nand U21354 (N_21354,N_19713,N_19985);
xor U21355 (N_21355,N_19906,N_19986);
nor U21356 (N_21356,N_20392,N_19606);
and U21357 (N_21357,N_19632,N_19912);
nand U21358 (N_21358,N_19578,N_20240);
and U21359 (N_21359,N_19459,N_19421);
nand U21360 (N_21360,N_19960,N_20292);
or U21361 (N_21361,N_19906,N_20092);
xnor U21362 (N_21362,N_19201,N_19602);
or U21363 (N_21363,N_20002,N_19573);
nand U21364 (N_21364,N_19294,N_19241);
nand U21365 (N_21365,N_19995,N_20312);
and U21366 (N_21366,N_19981,N_20113);
or U21367 (N_21367,N_19782,N_19584);
or U21368 (N_21368,N_19772,N_19549);
and U21369 (N_21369,N_19884,N_20327);
nor U21370 (N_21370,N_20390,N_19484);
nor U21371 (N_21371,N_20319,N_19796);
and U21372 (N_21372,N_19657,N_19546);
or U21373 (N_21373,N_19668,N_20190);
nor U21374 (N_21374,N_20214,N_19650);
nand U21375 (N_21375,N_19413,N_20108);
or U21376 (N_21376,N_19669,N_19514);
xor U21377 (N_21377,N_19965,N_19894);
nand U21378 (N_21378,N_19568,N_19595);
nand U21379 (N_21379,N_19510,N_19341);
or U21380 (N_21380,N_19732,N_20158);
or U21381 (N_21381,N_19294,N_19708);
and U21382 (N_21382,N_20290,N_19418);
or U21383 (N_21383,N_19792,N_19666);
or U21384 (N_21384,N_20371,N_19600);
nor U21385 (N_21385,N_19433,N_19971);
nand U21386 (N_21386,N_20081,N_19882);
xor U21387 (N_21387,N_19204,N_19812);
and U21388 (N_21388,N_19714,N_19470);
nor U21389 (N_21389,N_19514,N_19684);
nand U21390 (N_21390,N_19224,N_20292);
nor U21391 (N_21391,N_19227,N_19322);
or U21392 (N_21392,N_19939,N_20335);
or U21393 (N_21393,N_20121,N_19854);
nor U21394 (N_21394,N_19827,N_19370);
nand U21395 (N_21395,N_19831,N_20308);
xor U21396 (N_21396,N_19492,N_19622);
xor U21397 (N_21397,N_20317,N_19847);
nor U21398 (N_21398,N_19933,N_19234);
and U21399 (N_21399,N_20222,N_20286);
nor U21400 (N_21400,N_19856,N_19549);
nor U21401 (N_21401,N_20373,N_19686);
nand U21402 (N_21402,N_19490,N_19347);
or U21403 (N_21403,N_19451,N_19411);
and U21404 (N_21404,N_20143,N_19234);
nor U21405 (N_21405,N_19687,N_19977);
nand U21406 (N_21406,N_19370,N_19962);
xnor U21407 (N_21407,N_20241,N_19931);
nor U21408 (N_21408,N_20195,N_19816);
nand U21409 (N_21409,N_20084,N_19323);
xor U21410 (N_21410,N_20279,N_19281);
and U21411 (N_21411,N_19455,N_20124);
or U21412 (N_21412,N_19213,N_19875);
nor U21413 (N_21413,N_20185,N_19767);
and U21414 (N_21414,N_19298,N_20147);
xor U21415 (N_21415,N_19283,N_20338);
nor U21416 (N_21416,N_20009,N_20256);
nand U21417 (N_21417,N_19934,N_19247);
nand U21418 (N_21418,N_19652,N_19221);
xor U21419 (N_21419,N_19297,N_19467);
or U21420 (N_21420,N_20170,N_20308);
or U21421 (N_21421,N_19876,N_19747);
nor U21422 (N_21422,N_20226,N_19325);
and U21423 (N_21423,N_19587,N_20140);
nand U21424 (N_21424,N_20002,N_19804);
and U21425 (N_21425,N_20365,N_20167);
nand U21426 (N_21426,N_20146,N_19335);
nor U21427 (N_21427,N_19895,N_20125);
xor U21428 (N_21428,N_20163,N_19501);
nand U21429 (N_21429,N_20193,N_19693);
nand U21430 (N_21430,N_19222,N_20186);
and U21431 (N_21431,N_19337,N_19544);
nor U21432 (N_21432,N_19936,N_19244);
nor U21433 (N_21433,N_19597,N_19856);
nand U21434 (N_21434,N_19663,N_19834);
and U21435 (N_21435,N_19417,N_20036);
and U21436 (N_21436,N_19741,N_19677);
or U21437 (N_21437,N_19460,N_20118);
xnor U21438 (N_21438,N_20358,N_19690);
nor U21439 (N_21439,N_19552,N_19678);
nand U21440 (N_21440,N_19338,N_20003);
and U21441 (N_21441,N_19706,N_19653);
nand U21442 (N_21442,N_19920,N_19760);
nand U21443 (N_21443,N_19723,N_20061);
xor U21444 (N_21444,N_19887,N_20350);
or U21445 (N_21445,N_19514,N_19239);
nor U21446 (N_21446,N_19297,N_20013);
nand U21447 (N_21447,N_19970,N_19734);
xnor U21448 (N_21448,N_19317,N_19749);
or U21449 (N_21449,N_19321,N_19527);
xnor U21450 (N_21450,N_19682,N_19753);
and U21451 (N_21451,N_19239,N_19803);
nand U21452 (N_21452,N_20227,N_19717);
nor U21453 (N_21453,N_20222,N_19663);
nor U21454 (N_21454,N_19803,N_19632);
nand U21455 (N_21455,N_19241,N_20121);
and U21456 (N_21456,N_20101,N_19911);
or U21457 (N_21457,N_20262,N_19663);
nor U21458 (N_21458,N_19630,N_20002);
nor U21459 (N_21459,N_20233,N_20141);
or U21460 (N_21460,N_20221,N_19476);
nand U21461 (N_21461,N_19348,N_19833);
nor U21462 (N_21462,N_19364,N_19557);
nand U21463 (N_21463,N_19313,N_19565);
xnor U21464 (N_21464,N_19792,N_20071);
nand U21465 (N_21465,N_19790,N_19799);
nand U21466 (N_21466,N_19498,N_20017);
and U21467 (N_21467,N_20335,N_19780);
nand U21468 (N_21468,N_19888,N_19828);
or U21469 (N_21469,N_19234,N_20270);
and U21470 (N_21470,N_20131,N_19657);
and U21471 (N_21471,N_20032,N_19421);
xor U21472 (N_21472,N_19514,N_20379);
or U21473 (N_21473,N_19760,N_19545);
nand U21474 (N_21474,N_20179,N_19238);
nand U21475 (N_21475,N_20307,N_20230);
xnor U21476 (N_21476,N_19739,N_20390);
nand U21477 (N_21477,N_19261,N_19626);
xnor U21478 (N_21478,N_20091,N_19408);
nor U21479 (N_21479,N_19922,N_19334);
and U21480 (N_21480,N_20325,N_20222);
xnor U21481 (N_21481,N_19361,N_19288);
and U21482 (N_21482,N_19316,N_19420);
nor U21483 (N_21483,N_20043,N_20084);
and U21484 (N_21484,N_19731,N_20087);
xnor U21485 (N_21485,N_20046,N_19912);
or U21486 (N_21486,N_19831,N_20396);
nor U21487 (N_21487,N_20247,N_19552);
xnor U21488 (N_21488,N_19263,N_19307);
nor U21489 (N_21489,N_19228,N_19446);
xnor U21490 (N_21490,N_20368,N_20195);
or U21491 (N_21491,N_20042,N_20166);
nand U21492 (N_21492,N_20364,N_20202);
nor U21493 (N_21493,N_20062,N_19380);
xnor U21494 (N_21494,N_20196,N_19302);
and U21495 (N_21495,N_20188,N_20359);
nor U21496 (N_21496,N_19857,N_19965);
xnor U21497 (N_21497,N_19792,N_19560);
nor U21498 (N_21498,N_19522,N_20214);
nor U21499 (N_21499,N_20320,N_19947);
or U21500 (N_21500,N_19639,N_19444);
and U21501 (N_21501,N_19316,N_20085);
nand U21502 (N_21502,N_20041,N_19559);
xor U21503 (N_21503,N_20363,N_20371);
xnor U21504 (N_21504,N_20171,N_20250);
xor U21505 (N_21505,N_20215,N_19753);
xnor U21506 (N_21506,N_20228,N_20202);
and U21507 (N_21507,N_20308,N_19801);
and U21508 (N_21508,N_20353,N_19723);
and U21509 (N_21509,N_19641,N_19908);
nor U21510 (N_21510,N_20260,N_19220);
nor U21511 (N_21511,N_20111,N_20196);
or U21512 (N_21512,N_19400,N_19248);
or U21513 (N_21513,N_20203,N_19686);
or U21514 (N_21514,N_19842,N_20363);
xnor U21515 (N_21515,N_20368,N_19404);
and U21516 (N_21516,N_20379,N_19431);
xnor U21517 (N_21517,N_19664,N_20348);
and U21518 (N_21518,N_19626,N_19871);
nand U21519 (N_21519,N_19305,N_19577);
nor U21520 (N_21520,N_19439,N_19263);
nor U21521 (N_21521,N_19937,N_20315);
nand U21522 (N_21522,N_19274,N_19527);
xnor U21523 (N_21523,N_19910,N_19407);
and U21524 (N_21524,N_20146,N_20333);
and U21525 (N_21525,N_19674,N_20189);
and U21526 (N_21526,N_19798,N_20143);
nand U21527 (N_21527,N_20394,N_20155);
xnor U21528 (N_21528,N_19318,N_19424);
and U21529 (N_21529,N_20063,N_20066);
and U21530 (N_21530,N_19367,N_19244);
nand U21531 (N_21531,N_20023,N_20286);
or U21532 (N_21532,N_19541,N_20098);
or U21533 (N_21533,N_19268,N_19229);
nor U21534 (N_21534,N_20183,N_19602);
and U21535 (N_21535,N_19232,N_19341);
xor U21536 (N_21536,N_19779,N_20365);
nor U21537 (N_21537,N_19718,N_19959);
or U21538 (N_21538,N_19789,N_19584);
and U21539 (N_21539,N_19871,N_20358);
nor U21540 (N_21540,N_20328,N_20076);
xor U21541 (N_21541,N_20054,N_19736);
xor U21542 (N_21542,N_19777,N_19776);
and U21543 (N_21543,N_19342,N_19751);
nand U21544 (N_21544,N_19289,N_19529);
or U21545 (N_21545,N_20282,N_20077);
nor U21546 (N_21546,N_19611,N_19972);
xor U21547 (N_21547,N_19649,N_19808);
xor U21548 (N_21548,N_19210,N_19962);
nand U21549 (N_21549,N_19355,N_19979);
nor U21550 (N_21550,N_20245,N_19732);
and U21551 (N_21551,N_19222,N_19268);
nand U21552 (N_21552,N_19682,N_19588);
nand U21553 (N_21553,N_20087,N_20085);
or U21554 (N_21554,N_19254,N_19256);
xnor U21555 (N_21555,N_20306,N_19869);
nor U21556 (N_21556,N_20009,N_20263);
and U21557 (N_21557,N_19267,N_20294);
xor U21558 (N_21558,N_19573,N_20326);
nor U21559 (N_21559,N_20009,N_19538);
nor U21560 (N_21560,N_19557,N_20194);
nor U21561 (N_21561,N_20192,N_19282);
nor U21562 (N_21562,N_20351,N_20138);
and U21563 (N_21563,N_19339,N_19942);
or U21564 (N_21564,N_20019,N_19910);
xor U21565 (N_21565,N_19573,N_20358);
nand U21566 (N_21566,N_19388,N_20300);
or U21567 (N_21567,N_19427,N_19951);
xor U21568 (N_21568,N_19959,N_19307);
or U21569 (N_21569,N_19634,N_19660);
and U21570 (N_21570,N_19847,N_19257);
nand U21571 (N_21571,N_19258,N_19912);
nor U21572 (N_21572,N_20011,N_19347);
nand U21573 (N_21573,N_19555,N_19892);
xor U21574 (N_21574,N_19791,N_20375);
nand U21575 (N_21575,N_19579,N_20074);
or U21576 (N_21576,N_20156,N_19227);
and U21577 (N_21577,N_20311,N_19535);
nor U21578 (N_21578,N_19305,N_19788);
nor U21579 (N_21579,N_19755,N_19716);
and U21580 (N_21580,N_19867,N_19436);
xnor U21581 (N_21581,N_19398,N_19539);
and U21582 (N_21582,N_19738,N_19567);
nor U21583 (N_21583,N_19685,N_20268);
nor U21584 (N_21584,N_20328,N_19301);
xnor U21585 (N_21585,N_19408,N_19351);
or U21586 (N_21586,N_20324,N_19901);
nor U21587 (N_21587,N_19528,N_20126);
or U21588 (N_21588,N_19634,N_19245);
nand U21589 (N_21589,N_20018,N_20064);
and U21590 (N_21590,N_19498,N_20312);
nor U21591 (N_21591,N_19493,N_19931);
nor U21592 (N_21592,N_19811,N_19303);
and U21593 (N_21593,N_19749,N_19740);
or U21594 (N_21594,N_19208,N_20016);
nand U21595 (N_21595,N_20105,N_20126);
xor U21596 (N_21596,N_19509,N_20182);
or U21597 (N_21597,N_19967,N_19398);
and U21598 (N_21598,N_20271,N_20051);
xor U21599 (N_21599,N_20310,N_20291);
xor U21600 (N_21600,N_21468,N_20551);
and U21601 (N_21601,N_20737,N_20959);
nand U21602 (N_21602,N_21004,N_20542);
and U21603 (N_21603,N_20515,N_20576);
xnor U21604 (N_21604,N_20885,N_21342);
xor U21605 (N_21605,N_21106,N_20827);
and U21606 (N_21606,N_21139,N_21421);
or U21607 (N_21607,N_20539,N_20916);
or U21608 (N_21608,N_20441,N_20455);
xnor U21609 (N_21609,N_20621,N_20584);
xnor U21610 (N_21610,N_21596,N_20465);
xnor U21611 (N_21611,N_21314,N_20945);
nand U21612 (N_21612,N_21360,N_20967);
or U21613 (N_21613,N_20847,N_21080);
nand U21614 (N_21614,N_20603,N_20487);
or U21615 (N_21615,N_20588,N_20419);
nor U21616 (N_21616,N_21059,N_20920);
nand U21617 (N_21617,N_21144,N_20891);
nor U21618 (N_21618,N_21481,N_20851);
or U21619 (N_21619,N_21420,N_21132);
nor U21620 (N_21620,N_20793,N_20919);
xor U21621 (N_21621,N_20813,N_20437);
or U21622 (N_21622,N_21480,N_20569);
xor U21623 (N_21623,N_20833,N_21138);
and U21624 (N_21624,N_20453,N_21150);
xnor U21625 (N_21625,N_20805,N_21504);
and U21626 (N_21626,N_20798,N_21275);
or U21627 (N_21627,N_21437,N_21198);
xor U21628 (N_21628,N_20922,N_20877);
nor U21629 (N_21629,N_20616,N_20953);
and U21630 (N_21630,N_21436,N_20864);
xnor U21631 (N_21631,N_21321,N_21370);
nor U21632 (N_21632,N_20881,N_20933);
nor U21633 (N_21633,N_20804,N_20684);
or U21634 (N_21634,N_20510,N_21135);
xor U21635 (N_21635,N_21500,N_20788);
xor U21636 (N_21636,N_21580,N_20770);
nand U21637 (N_21637,N_21359,N_20894);
and U21638 (N_21638,N_20963,N_20928);
or U21639 (N_21639,N_21247,N_21367);
or U21640 (N_21640,N_21079,N_21007);
nand U21641 (N_21641,N_20996,N_21153);
xnor U21642 (N_21642,N_20690,N_20811);
nand U21643 (N_21643,N_21264,N_20674);
nand U21644 (N_21644,N_21239,N_21048);
xnor U21645 (N_21645,N_21305,N_20452);
and U21646 (N_21646,N_20949,N_20796);
xnor U21647 (N_21647,N_21592,N_21438);
xor U21648 (N_21648,N_20818,N_21570);
or U21649 (N_21649,N_20748,N_20589);
nand U21650 (N_21650,N_21200,N_21245);
or U21651 (N_21651,N_21373,N_21148);
xor U21652 (N_21652,N_21558,N_21161);
xor U21653 (N_21653,N_20725,N_21565);
nand U21654 (N_21654,N_20826,N_20743);
nand U21655 (N_21655,N_21113,N_20718);
nor U21656 (N_21656,N_20794,N_21499);
nand U21657 (N_21657,N_21516,N_20713);
xor U21658 (N_21658,N_21304,N_21385);
or U21659 (N_21659,N_20628,N_20611);
or U21660 (N_21660,N_21316,N_20548);
or U21661 (N_21661,N_21224,N_20578);
xor U21662 (N_21662,N_21221,N_21186);
nor U21663 (N_21663,N_21515,N_20937);
xnor U21664 (N_21664,N_20809,N_21018);
nor U21665 (N_21665,N_21082,N_20846);
xnor U21666 (N_21666,N_21534,N_20618);
and U21667 (N_21667,N_20839,N_20635);
and U21668 (N_21668,N_20544,N_21085);
nand U21669 (N_21669,N_20697,N_21593);
and U21670 (N_21670,N_20650,N_21584);
xor U21671 (N_21671,N_20552,N_20471);
xnor U21672 (N_21672,N_21492,N_20520);
or U21673 (N_21673,N_20500,N_21390);
or U21674 (N_21674,N_21361,N_21526);
or U21675 (N_21675,N_21117,N_20422);
or U21676 (N_21676,N_21181,N_20879);
and U21677 (N_21677,N_21167,N_21552);
nand U21678 (N_21678,N_21425,N_20853);
and U21679 (N_21679,N_20609,N_21339);
nand U21680 (N_21680,N_21043,N_20705);
and U21681 (N_21681,N_21017,N_20873);
nor U21682 (N_21682,N_21511,N_20456);
nor U21683 (N_21683,N_21062,N_20900);
nor U21684 (N_21684,N_21072,N_20810);
nand U21685 (N_21685,N_21077,N_21130);
nor U21686 (N_21686,N_21065,N_20675);
xor U21687 (N_21687,N_20991,N_20480);
nand U21688 (N_21688,N_21573,N_20720);
nor U21689 (N_21689,N_21013,N_21459);
and U21690 (N_21690,N_20987,N_20492);
nor U21691 (N_21691,N_20936,N_21328);
xor U21692 (N_21692,N_20403,N_21280);
nor U21693 (N_21693,N_20753,N_21574);
nand U21694 (N_21694,N_21154,N_20474);
xnor U21695 (N_21695,N_20962,N_20773);
or U21696 (N_21696,N_20482,N_21112);
or U21697 (N_21697,N_21118,N_21016);
or U21698 (N_21698,N_20964,N_20424);
nor U21699 (N_21699,N_20447,N_21332);
nand U21700 (N_21700,N_21021,N_21472);
nand U21701 (N_21701,N_21039,N_21012);
and U21702 (N_21702,N_20974,N_21075);
or U21703 (N_21703,N_21233,N_21238);
nor U21704 (N_21704,N_21493,N_21288);
nand U21705 (N_21705,N_20736,N_20844);
nor U21706 (N_21706,N_20493,N_21356);
nor U21707 (N_21707,N_20440,N_20625);
xor U21708 (N_21708,N_21488,N_20498);
or U21709 (N_21709,N_20477,N_21097);
and U21710 (N_21710,N_21454,N_21538);
nor U21711 (N_21711,N_21351,N_21358);
nor U21712 (N_21712,N_20665,N_21341);
nand U21713 (N_21713,N_20802,N_21163);
or U21714 (N_21714,N_21450,N_20405);
or U21715 (N_21715,N_20613,N_20408);
xnor U21716 (N_21716,N_20789,N_21562);
nand U21717 (N_21717,N_20745,N_21445);
or U21718 (N_21718,N_21164,N_20768);
xnor U21719 (N_21719,N_21255,N_21599);
xnor U21720 (N_21720,N_20411,N_20428);
xnor U21721 (N_21721,N_20526,N_20418);
xnor U21722 (N_21722,N_20639,N_21069);
xor U21723 (N_21723,N_20727,N_20895);
nor U21724 (N_21724,N_20950,N_21095);
xnor U21725 (N_21725,N_21152,N_20828);
or U21726 (N_21726,N_21416,N_21467);
xor U21727 (N_21727,N_21060,N_20763);
or U21728 (N_21728,N_20470,N_20606);
or U21729 (N_21729,N_21276,N_20409);
nor U21730 (N_21730,N_21386,N_21058);
xor U21731 (N_21731,N_20558,N_21108);
xor U21732 (N_21732,N_21290,N_21340);
or U21733 (N_21733,N_20443,N_21478);
xor U21734 (N_21734,N_21178,N_21347);
and U21735 (N_21735,N_21453,N_20728);
nand U21736 (N_21736,N_20931,N_21409);
nand U21737 (N_21737,N_21482,N_21536);
nor U21738 (N_21738,N_20645,N_21399);
nor U21739 (N_21739,N_20497,N_21303);
nand U21740 (N_21740,N_21365,N_20467);
and U21741 (N_21741,N_20774,N_21327);
nand U21742 (N_21742,N_21406,N_20537);
xor U21743 (N_21743,N_21171,N_20593);
nor U21744 (N_21744,N_21187,N_20730);
or U21745 (N_21745,N_20610,N_21291);
or U21746 (N_21746,N_21388,N_20733);
xor U21747 (N_21747,N_20561,N_21136);
nand U21748 (N_21748,N_21109,N_21597);
and U21749 (N_21749,N_20619,N_21297);
or U21750 (N_21750,N_20800,N_21479);
or U21751 (N_21751,N_21429,N_20431);
or U21752 (N_21752,N_20943,N_20653);
or U21753 (N_21753,N_21506,N_20444);
nand U21754 (N_21754,N_20660,N_21522);
nand U21755 (N_21755,N_20824,N_21011);
or U21756 (N_21756,N_21268,N_21334);
and U21757 (N_21757,N_21146,N_21545);
nand U21758 (N_21758,N_21142,N_20948);
xor U21759 (N_21759,N_21124,N_21322);
nand U21760 (N_21760,N_20764,N_21009);
or U21761 (N_21761,N_20785,N_21513);
nand U21762 (N_21762,N_21432,N_20981);
nand U21763 (N_21763,N_21363,N_20449);
and U21764 (N_21764,N_21527,N_20801);
nor U21765 (N_21765,N_20508,N_20631);
nand U21766 (N_21766,N_20755,N_21444);
and U21767 (N_21767,N_21179,N_21369);
nor U21768 (N_21768,N_21403,N_21311);
and U21769 (N_21769,N_20915,N_21242);
nand U21770 (N_21770,N_21234,N_21222);
and U21771 (N_21771,N_20486,N_21248);
xor U21772 (N_21772,N_21343,N_21448);
xor U21773 (N_21773,N_20462,N_20531);
or U21774 (N_21774,N_20909,N_21578);
nand U21775 (N_21775,N_21038,N_21315);
xor U21776 (N_21776,N_20630,N_20546);
nor U21777 (N_21777,N_21495,N_21357);
nor U21778 (N_21778,N_20874,N_20516);
nand U21779 (N_21779,N_21405,N_20892);
and U21780 (N_21780,N_20901,N_20756);
nor U21781 (N_21781,N_20685,N_20412);
nand U21782 (N_21782,N_20686,N_20912);
nand U21783 (N_21783,N_20760,N_20511);
nand U21784 (N_21784,N_21175,N_20734);
and U21785 (N_21785,N_21458,N_21204);
xor U21786 (N_21786,N_21494,N_21557);
or U21787 (N_21787,N_20825,N_20829);
xor U21788 (N_21788,N_21465,N_21063);
nand U21789 (N_21789,N_20681,N_21176);
or U21790 (N_21790,N_21030,N_21211);
xor U21791 (N_21791,N_20955,N_20893);
nor U21792 (N_21792,N_21031,N_21073);
and U21793 (N_21793,N_20530,N_21093);
or U21794 (N_21794,N_20680,N_21090);
or U21795 (N_21795,N_21123,N_21168);
nand U21796 (N_21796,N_21089,N_21270);
and U21797 (N_21797,N_21254,N_20598);
nor U21798 (N_21798,N_20747,N_20401);
or U21799 (N_21799,N_21419,N_20795);
nand U21800 (N_21800,N_20757,N_21035);
and U21801 (N_21801,N_21267,N_21391);
nor U21802 (N_21802,N_21446,N_20975);
nand U21803 (N_21803,N_20778,N_21330);
xnor U21804 (N_21804,N_20568,N_21217);
nor U21805 (N_21805,N_20769,N_20535);
or U21806 (N_21806,N_20518,N_21491);
nand U21807 (N_21807,N_20481,N_21568);
or U21808 (N_21808,N_20522,N_20654);
and U21809 (N_21809,N_20643,N_20523);
or U21810 (N_21810,N_20458,N_21382);
xnor U21811 (N_21811,N_20559,N_21577);
nand U21812 (N_21812,N_21583,N_21366);
and U21813 (N_21813,N_21216,N_20608);
or U21814 (N_21814,N_21532,N_20514);
and U21815 (N_21815,N_20495,N_20624);
nand U21816 (N_21816,N_20432,N_20923);
nand U21817 (N_21817,N_21046,N_20957);
nor U21818 (N_21818,N_21227,N_21244);
xnor U21819 (N_21819,N_20404,N_20865);
xor U21820 (N_21820,N_21548,N_21331);
or U21821 (N_21821,N_20636,N_21126);
xnor U21822 (N_21822,N_20792,N_20536);
or U21823 (N_21823,N_20840,N_21189);
xnor U21824 (N_21824,N_20944,N_21251);
and U21825 (N_21825,N_21026,N_20573);
nor U21826 (N_21826,N_21040,N_21354);
nor U21827 (N_21827,N_20821,N_20704);
nand U21828 (N_21828,N_20956,N_20656);
nand U21829 (N_21829,N_20822,N_20862);
or U21830 (N_21830,N_21309,N_20940);
and U21831 (N_21831,N_21439,N_21197);
and U21832 (N_21832,N_20433,N_21434);
or U21833 (N_21833,N_21215,N_20410);
and U21834 (N_21834,N_20448,N_20600);
xnor U21835 (N_21835,N_21487,N_21071);
xnor U21836 (N_21836,N_21044,N_21508);
nand U21837 (N_21837,N_20938,N_21301);
or U21838 (N_21838,N_21414,N_20958);
or U21839 (N_21839,N_21023,N_21456);
or U21840 (N_21840,N_20927,N_21166);
xor U21841 (N_21841,N_20596,N_21306);
nor U21842 (N_21842,N_20429,N_20952);
or U21843 (N_21843,N_21585,N_20466);
nand U21844 (N_21844,N_20906,N_20560);
xor U21845 (N_21845,N_21287,N_20632);
and U21846 (N_21846,N_21094,N_20907);
nor U21847 (N_21847,N_20807,N_20642);
or U21848 (N_21848,N_21129,N_21477);
nor U21849 (N_21849,N_21269,N_21134);
nor U21850 (N_21850,N_20423,N_21034);
xnor U21851 (N_21851,N_20622,N_20668);
and U21852 (N_21852,N_21127,N_20972);
nand U21853 (N_21853,N_20838,N_21353);
or U21854 (N_21854,N_20849,N_20716);
or U21855 (N_21855,N_21214,N_21283);
xor U21856 (N_21856,N_21225,N_20905);
or U21857 (N_21857,N_21313,N_20436);
nor U21858 (N_21858,N_20776,N_20977);
xor U21859 (N_21859,N_20832,N_21338);
xnor U21860 (N_21860,N_20871,N_21005);
and U21861 (N_21861,N_21451,N_21258);
or U21862 (N_21862,N_21027,N_20939);
xnor U21863 (N_21863,N_20579,N_21293);
nand U21864 (N_21864,N_21470,N_21555);
nand U21865 (N_21865,N_21520,N_20714);
nand U21866 (N_21866,N_21539,N_20563);
and U21867 (N_21867,N_20925,N_20960);
and U21868 (N_21868,N_20759,N_20499);
nand U21869 (N_21869,N_20484,N_20911);
xnor U21870 (N_21870,N_21279,N_21423);
xnor U21871 (N_21871,N_21202,N_20689);
and U21872 (N_21872,N_20994,N_21307);
and U21873 (N_21873,N_21010,N_20935);
xnor U21874 (N_21874,N_20875,N_21252);
nor U21875 (N_21875,N_21115,N_20547);
or U21876 (N_21876,N_21551,N_20751);
xnor U21877 (N_21877,N_20854,N_21497);
nand U21878 (N_21878,N_21260,N_21404);
nor U21879 (N_21879,N_21282,N_21485);
nand U21880 (N_21880,N_21246,N_21169);
nand U21881 (N_21881,N_21447,N_20472);
nand U21882 (N_21882,N_20904,N_20857);
nor U21883 (N_21883,N_21512,N_20494);
or U21884 (N_21884,N_20886,N_21469);
nor U21885 (N_21885,N_21483,N_21165);
or U21886 (N_21886,N_20671,N_20657);
nor U21887 (N_21887,N_21368,N_20435);
and U21888 (N_21888,N_21586,N_21542);
nand U21889 (N_21889,N_21022,N_21582);
nand U21890 (N_21890,N_21078,N_20662);
nand U21891 (N_21891,N_21519,N_21336);
or U21892 (N_21892,N_20664,N_20717);
or U21893 (N_21893,N_21442,N_21412);
and U21894 (N_21894,N_20669,N_21559);
xor U21895 (N_21895,N_21571,N_21070);
or U21896 (N_21896,N_21277,N_20791);
and U21897 (N_21897,N_20746,N_21033);
and U21898 (N_21898,N_21104,N_20597);
nand U21899 (N_21899,N_21317,N_21424);
xor U21900 (N_21900,N_21145,N_21474);
and U21901 (N_21901,N_21119,N_21333);
or U21902 (N_21902,N_20426,N_20623);
nor U21903 (N_21903,N_21231,N_20852);
nand U21904 (N_21904,N_21084,N_20702);
nand U21905 (N_21905,N_20999,N_21100);
and U21906 (N_21906,N_21344,N_21426);
and U21907 (N_21907,N_20682,N_21524);
or U21908 (N_21908,N_20965,N_21281);
nand U21909 (N_21909,N_20688,N_20858);
and U21910 (N_21910,N_21335,N_21476);
or U21911 (N_21911,N_20430,N_20869);
xnor U21912 (N_21912,N_20476,N_21208);
nor U21913 (N_21913,N_21230,N_20451);
and U21914 (N_21914,N_20841,N_20533);
nor U21915 (N_21915,N_20557,N_20509);
xnor U21916 (N_21916,N_21387,N_20941);
and U21917 (N_21917,N_21151,N_20979);
xor U21918 (N_21918,N_20951,N_20903);
xnor U21919 (N_21919,N_21261,N_20843);
nand U21920 (N_21920,N_20607,N_21392);
or U21921 (N_21921,N_20438,N_20407);
and U21922 (N_21922,N_21249,N_20910);
nand U21923 (N_21923,N_21308,N_20421);
or U21924 (N_21924,N_20729,N_20652);
nor U21925 (N_21925,N_20525,N_20504);
nand U21926 (N_21926,N_20961,N_21041);
xor U21927 (N_21927,N_21226,N_21503);
and U21928 (N_21928,N_20651,N_20666);
and U21929 (N_21929,N_21285,N_20779);
nor U21930 (N_21930,N_21173,N_20888);
nand U21931 (N_21931,N_21296,N_21320);
nand U21932 (N_21932,N_21433,N_21220);
xnor U21933 (N_21933,N_21210,N_20954);
or U21934 (N_21934,N_21116,N_21489);
and U21935 (N_21935,N_20890,N_20781);
and U21936 (N_21936,N_21273,N_21380);
and U21937 (N_21937,N_20703,N_21182);
xor U21938 (N_21938,N_21449,N_21008);
and U21939 (N_21939,N_20914,N_20541);
nand U21940 (N_21940,N_21457,N_20816);
xnor U21941 (N_21941,N_21535,N_21372);
or U21942 (N_21942,N_20540,N_21203);
xnor U21943 (N_21943,N_21411,N_21521);
or U21944 (N_21944,N_20633,N_20501);
or U21945 (N_21945,N_20754,N_20599);
nand U21946 (N_21946,N_20868,N_20580);
xor U21947 (N_21947,N_21143,N_21323);
or U21948 (N_21948,N_20677,N_20947);
and U21949 (N_21949,N_21422,N_20724);
nand U21950 (N_21950,N_21529,N_20762);
nand U21951 (N_21951,N_21378,N_20420);
nor U21952 (N_21952,N_21110,N_21196);
or U21953 (N_21953,N_21137,N_20679);
or U21954 (N_21954,N_20620,N_20924);
or U21955 (N_21955,N_21128,N_20988);
nor U21956 (N_21956,N_21371,N_21199);
and U21957 (N_21957,N_21505,N_20878);
xor U21958 (N_21958,N_21501,N_20581);
xnor U21959 (N_21959,N_20591,N_20836);
nor U21960 (N_21960,N_20750,N_20771);
or U21961 (N_21961,N_20659,N_20842);
nand U21962 (N_21962,N_21241,N_21598);
and U21963 (N_21963,N_21096,N_21190);
or U21964 (N_21964,N_21289,N_21443);
nor U21965 (N_21965,N_20766,N_21410);
xnor U21966 (N_21966,N_21595,N_21006);
xnor U21967 (N_21967,N_20461,N_21431);
and U21968 (N_21968,N_21484,N_21417);
nand U21969 (N_21969,N_21384,N_20637);
nand U21970 (N_21970,N_21355,N_20738);
nand U21971 (N_21971,N_21594,N_20899);
nor U21972 (N_21972,N_20932,N_20698);
xnor U21973 (N_21973,N_20434,N_21374);
nor U21974 (N_21974,N_20855,N_21083);
nor U21975 (N_21975,N_20880,N_21122);
nand U21976 (N_21976,N_21101,N_21028);
nand U21977 (N_21977,N_20982,N_20752);
xnor U21978 (N_21978,N_21274,N_20971);
xnor U21979 (N_21979,N_20913,N_21589);
xor U21980 (N_21980,N_21286,N_20627);
and U21981 (N_21981,N_20612,N_20983);
nor U21982 (N_21982,N_21345,N_20966);
nor U21983 (N_21983,N_20695,N_20896);
nand U21984 (N_21984,N_21057,N_20799);
and U21985 (N_21985,N_21235,N_20882);
nor U21986 (N_21986,N_20427,N_21473);
and U21987 (N_21987,N_21440,N_20532);
nand U21988 (N_21988,N_20787,N_20739);
nor U21989 (N_21989,N_21061,N_20694);
nor U21990 (N_21990,N_20594,N_21540);
xor U21991 (N_21991,N_21180,N_21563);
nand U21992 (N_21992,N_20845,N_21103);
nor U21993 (N_21993,N_21206,N_21502);
xor U21994 (N_21994,N_21088,N_20574);
nand U21995 (N_21995,N_20969,N_20700);
nor U21996 (N_21996,N_20506,N_21407);
nand U21997 (N_21997,N_21319,N_20555);
and U21998 (N_21998,N_21398,N_20808);
and U21999 (N_21999,N_20978,N_21195);
and U22000 (N_22000,N_20595,N_21158);
xnor U22001 (N_22001,N_20819,N_21350);
xnor U22002 (N_22002,N_21091,N_21174);
xor U22003 (N_22003,N_20726,N_20583);
and U22004 (N_22004,N_20735,N_20450);
xor U22005 (N_22005,N_21566,N_21262);
xor U22006 (N_22006,N_21408,N_20614);
or U22007 (N_22007,N_21564,N_21185);
and U22008 (N_22008,N_20732,N_20775);
or U22009 (N_22009,N_21299,N_20538);
or U22010 (N_22010,N_20908,N_20439);
and U22011 (N_22011,N_20806,N_21256);
nor U22012 (N_22012,N_21149,N_20721);
nor U22013 (N_22013,N_21510,N_21157);
xnor U22014 (N_22014,N_20565,N_20459);
and U22015 (N_22015,N_20490,N_20850);
or U22016 (N_22016,N_20970,N_21554);
or U22017 (N_22017,N_20820,N_21086);
xnor U22018 (N_22018,N_20691,N_21184);
nor U22019 (N_22019,N_21223,N_20817);
and U22020 (N_22020,N_21383,N_21509);
or U22021 (N_22021,N_20711,N_20496);
xor U22022 (N_22022,N_20780,N_20758);
nand U22023 (N_22023,N_20921,N_21415);
and U22024 (N_22024,N_21105,N_21219);
xor U22025 (N_22025,N_21427,N_21212);
xnor U22026 (N_22026,N_21015,N_20777);
nor U22027 (N_22027,N_21049,N_21402);
or U22028 (N_22028,N_20926,N_20634);
and U22029 (N_22029,N_20709,N_20989);
or U22030 (N_22030,N_21528,N_20658);
nand U22031 (N_22031,N_21537,N_21576);
nand U22032 (N_22032,N_21092,N_21243);
nand U22033 (N_22033,N_20861,N_20812);
and U22034 (N_22034,N_21324,N_21591);
nand U22035 (N_22035,N_21462,N_21236);
and U22036 (N_22036,N_20867,N_20837);
nor U22037 (N_22037,N_21302,N_20876);
nand U22038 (N_22038,N_20414,N_21561);
nand U22039 (N_22039,N_21120,N_21588);
and U22040 (N_22040,N_20898,N_21194);
and U22041 (N_22041,N_21032,N_20749);
and U22042 (N_22042,N_21053,N_21569);
xnor U22043 (N_22043,N_20934,N_20930);
nand U22044 (N_22044,N_20998,N_21162);
nor U22045 (N_22045,N_20507,N_21172);
and U22046 (N_22046,N_20483,N_20446);
nor U22047 (N_22047,N_21253,N_20503);
and U22048 (N_22048,N_20997,N_20670);
nand U22049 (N_22049,N_21364,N_20765);
and U22050 (N_22050,N_20577,N_20712);
or U22051 (N_22051,N_21192,N_20566);
nand U22052 (N_22052,N_21329,N_21461);
xor U22053 (N_22053,N_20457,N_21400);
and U22054 (N_22054,N_21544,N_21518);
xor U22055 (N_22055,N_21418,N_21001);
nor U22056 (N_22056,N_20460,N_21074);
xnor U22057 (N_22057,N_21201,N_20673);
nand U22058 (N_22058,N_20491,N_20887);
or U22059 (N_22059,N_20556,N_20767);
or U22060 (N_22060,N_20863,N_21155);
and U22061 (N_22061,N_20406,N_21466);
xor U22062 (N_22062,N_20469,N_20782);
nor U22063 (N_22063,N_21209,N_20866);
nor U22064 (N_22064,N_20860,N_21218);
nand U22065 (N_22065,N_20502,N_20870);
nor U22066 (N_22066,N_21292,N_21579);
nor U22067 (N_22067,N_20413,N_20917);
nand U22068 (N_22068,N_21525,N_20835);
xnor U22069 (N_22069,N_21054,N_21193);
or U22070 (N_22070,N_20696,N_21547);
nor U22071 (N_22071,N_21401,N_20701);
xor U22072 (N_22072,N_21055,N_20731);
xor U22073 (N_22073,N_20995,N_21250);
or U22074 (N_22074,N_21575,N_20534);
nand U22075 (N_22075,N_21232,N_20601);
or U22076 (N_22076,N_20485,N_21298);
nor U22077 (N_22077,N_21435,N_21295);
and U22078 (N_22078,N_20602,N_20571);
nand U22079 (N_22079,N_21000,N_21228);
or U22080 (N_22080,N_21377,N_21428);
and U22081 (N_22081,N_20647,N_20990);
nor U22082 (N_22082,N_21496,N_20676);
xor U22083 (N_22083,N_20872,N_20463);
nor U22084 (N_22084,N_20562,N_21348);
xor U22085 (N_22085,N_21272,N_21349);
and U22086 (N_22086,N_21523,N_21533);
nand U22087 (N_22087,N_20572,N_21133);
and U22088 (N_22088,N_21362,N_21068);
and U22089 (N_22089,N_21237,N_21486);
nand U22090 (N_22090,N_20445,N_20968);
and U22091 (N_22091,N_21213,N_21376);
nand U22092 (N_22092,N_21460,N_20442);
xnor U22093 (N_22093,N_21278,N_21550);
nor U22094 (N_22094,N_21590,N_21531);
nand U22095 (N_22095,N_21003,N_21543);
and U22096 (N_22096,N_20786,N_21455);
or U22097 (N_22097,N_21140,N_20464);
and U22098 (N_22098,N_21310,N_21463);
nor U22099 (N_22099,N_20587,N_21546);
nor U22100 (N_22100,N_20946,N_21259);
or U22101 (N_22101,N_21240,N_21475);
xor U22102 (N_22102,N_20488,N_21081);
xor U22103 (N_22103,N_20549,N_21318);
xnor U22104 (N_22104,N_20723,N_20706);
nand U22105 (N_22105,N_21107,N_20672);
nand U22106 (N_22106,N_20683,N_21025);
nor U22107 (N_22107,N_21325,N_20513);
xor U22108 (N_22108,N_21397,N_20626);
or U22109 (N_22109,N_20992,N_20400);
xor U22110 (N_22110,N_21067,N_21036);
nand U22111 (N_22111,N_21393,N_21587);
nand U22112 (N_22112,N_20929,N_20942);
and U22113 (N_22113,N_21160,N_20784);
nor U22114 (N_22114,N_21389,N_21326);
and U22115 (N_22115,N_21170,N_21430);
xnor U22116 (N_22116,N_21066,N_20667);
xnor U22117 (N_22117,N_20889,N_20814);
nand U22118 (N_22118,N_21553,N_21572);
xor U22119 (N_22119,N_20976,N_20761);
nor U22120 (N_22120,N_20521,N_20823);
or U22121 (N_22121,N_21188,N_20454);
nor U22122 (N_22122,N_20803,N_20902);
nand U22123 (N_22123,N_20719,N_21037);
and U22124 (N_22124,N_20517,N_20638);
xnor U22125 (N_22125,N_21045,N_20710);
nand U22126 (N_22126,N_20744,N_20986);
nand U22127 (N_22127,N_20797,N_21517);
nor U22128 (N_22128,N_21294,N_20848);
nand U22129 (N_22129,N_20692,N_20475);
and U22130 (N_22130,N_20856,N_21265);
nor U22131 (N_22131,N_21050,N_21056);
nor U22132 (N_22132,N_21159,N_21087);
or U22133 (N_22133,N_21125,N_20699);
or U22134 (N_22134,N_21271,N_20550);
xor U22135 (N_22135,N_21002,N_20742);
xor U22136 (N_22136,N_20604,N_20505);
nand U22137 (N_22137,N_21121,N_21395);
and U22138 (N_22138,N_20663,N_20582);
and U22139 (N_22139,N_20783,N_21099);
nand U22140 (N_22140,N_21284,N_20815);
or U22141 (N_22141,N_20567,N_20708);
and U22142 (N_22142,N_21337,N_20479);
and U22143 (N_22143,N_20512,N_21498);
or U22144 (N_22144,N_21490,N_20646);
and U22145 (N_22145,N_20478,N_21464);
xnor U22146 (N_22146,N_20524,N_20985);
nor U22147 (N_22147,N_21042,N_20772);
nand U22148 (N_22148,N_20830,N_21352);
xor U22149 (N_22149,N_20592,N_21300);
nand U22150 (N_22150,N_20543,N_20707);
nand U22151 (N_22151,N_20605,N_21312);
and U22152 (N_22152,N_20740,N_21560);
nor U22153 (N_22153,N_21514,N_20554);
xor U22154 (N_22154,N_21266,N_21207);
and U22155 (N_22155,N_20468,N_20831);
and U22156 (N_22156,N_21441,N_20590);
or U22157 (N_22157,N_21029,N_21379);
or U22158 (N_22158,N_20678,N_21263);
nor U22159 (N_22159,N_21375,N_20586);
xor U22160 (N_22160,N_20741,N_20417);
nand U22161 (N_22161,N_21396,N_21541);
or U22162 (N_22162,N_21381,N_20897);
and U22163 (N_22163,N_20489,N_21076);
nor U22164 (N_22164,N_21452,N_20884);
xor U22165 (N_22165,N_20722,N_21567);
or U22166 (N_22166,N_20649,N_21205);
or U22167 (N_22167,N_21111,N_20980);
and U22168 (N_22168,N_20655,N_20790);
nor U22169 (N_22169,N_21530,N_21413);
or U22170 (N_22170,N_21020,N_20641);
nor U22171 (N_22171,N_21156,N_21191);
nand U22172 (N_22172,N_20883,N_20687);
and U22173 (N_22173,N_20644,N_20918);
or U22174 (N_22174,N_21141,N_21051);
nand U22175 (N_22175,N_20425,N_20629);
xor U22176 (N_22176,N_20529,N_21098);
and U22177 (N_22177,N_21549,N_21394);
or U22178 (N_22178,N_20617,N_21047);
and U22179 (N_22179,N_20973,N_21131);
or U22180 (N_22180,N_20993,N_20615);
nand U22181 (N_22181,N_20693,N_20984);
or U22182 (N_22182,N_21229,N_21581);
nor U22183 (N_22183,N_21024,N_20570);
and U22184 (N_22184,N_20859,N_21507);
nand U22185 (N_22185,N_20834,N_21177);
nand U22186 (N_22186,N_20575,N_20545);
and U22187 (N_22187,N_21257,N_21014);
xor U22188 (N_22188,N_20648,N_21147);
nor U22189 (N_22189,N_20715,N_20564);
nand U22190 (N_22190,N_20640,N_20416);
xor U22191 (N_22191,N_21346,N_21102);
nand U22192 (N_22192,N_20585,N_21019);
xnor U22193 (N_22193,N_20661,N_20528);
or U22194 (N_22194,N_21052,N_20415);
nor U22195 (N_22195,N_21114,N_21556);
nand U22196 (N_22196,N_21183,N_21471);
nand U22197 (N_22197,N_20527,N_20519);
nor U22198 (N_22198,N_20402,N_21064);
nor U22199 (N_22199,N_20473,N_20553);
and U22200 (N_22200,N_21526,N_21294);
and U22201 (N_22201,N_20529,N_20630);
or U22202 (N_22202,N_21096,N_21014);
xor U22203 (N_22203,N_20686,N_21041);
and U22204 (N_22204,N_20959,N_20630);
and U22205 (N_22205,N_20990,N_21107);
xnor U22206 (N_22206,N_20642,N_21169);
or U22207 (N_22207,N_20434,N_20400);
nand U22208 (N_22208,N_20846,N_21391);
or U22209 (N_22209,N_21594,N_21307);
nor U22210 (N_22210,N_20921,N_20664);
nand U22211 (N_22211,N_20643,N_21218);
nand U22212 (N_22212,N_21462,N_20738);
nor U22213 (N_22213,N_21026,N_21226);
xor U22214 (N_22214,N_21304,N_20836);
nand U22215 (N_22215,N_21577,N_21387);
nand U22216 (N_22216,N_20689,N_21123);
and U22217 (N_22217,N_20529,N_20721);
xnor U22218 (N_22218,N_20701,N_20456);
and U22219 (N_22219,N_20936,N_21074);
or U22220 (N_22220,N_20436,N_20497);
and U22221 (N_22221,N_20447,N_20712);
nand U22222 (N_22222,N_21580,N_21573);
nand U22223 (N_22223,N_20905,N_20965);
nor U22224 (N_22224,N_20788,N_21594);
nand U22225 (N_22225,N_21527,N_21009);
nand U22226 (N_22226,N_21186,N_20787);
xor U22227 (N_22227,N_21121,N_21066);
or U22228 (N_22228,N_20917,N_20408);
and U22229 (N_22229,N_21298,N_21241);
nand U22230 (N_22230,N_20765,N_21029);
or U22231 (N_22231,N_20824,N_20871);
or U22232 (N_22232,N_21561,N_20819);
and U22233 (N_22233,N_21496,N_21127);
or U22234 (N_22234,N_20727,N_20754);
or U22235 (N_22235,N_20692,N_21562);
nand U22236 (N_22236,N_20465,N_21568);
nor U22237 (N_22237,N_21528,N_20922);
and U22238 (N_22238,N_21483,N_20736);
xor U22239 (N_22239,N_20885,N_20766);
or U22240 (N_22240,N_21081,N_21452);
and U22241 (N_22241,N_21578,N_20679);
nand U22242 (N_22242,N_21042,N_20821);
nor U22243 (N_22243,N_20867,N_20674);
xor U22244 (N_22244,N_20603,N_21312);
nor U22245 (N_22245,N_21312,N_20630);
or U22246 (N_22246,N_20977,N_20662);
nor U22247 (N_22247,N_21006,N_21090);
nand U22248 (N_22248,N_20648,N_21375);
and U22249 (N_22249,N_20805,N_21365);
nor U22250 (N_22250,N_20633,N_20651);
or U22251 (N_22251,N_21146,N_21369);
and U22252 (N_22252,N_20417,N_20634);
nor U22253 (N_22253,N_21415,N_20914);
nand U22254 (N_22254,N_20993,N_20918);
and U22255 (N_22255,N_20927,N_20748);
xnor U22256 (N_22256,N_20970,N_21278);
or U22257 (N_22257,N_20434,N_20736);
and U22258 (N_22258,N_20663,N_21413);
nand U22259 (N_22259,N_20810,N_20628);
nand U22260 (N_22260,N_21391,N_21594);
and U22261 (N_22261,N_21066,N_20668);
nand U22262 (N_22262,N_20542,N_21584);
nand U22263 (N_22263,N_21242,N_20635);
nor U22264 (N_22264,N_20752,N_21422);
or U22265 (N_22265,N_20811,N_21344);
and U22266 (N_22266,N_21285,N_20491);
or U22267 (N_22267,N_20728,N_21042);
and U22268 (N_22268,N_20417,N_20971);
and U22269 (N_22269,N_20446,N_21242);
xor U22270 (N_22270,N_21493,N_21222);
or U22271 (N_22271,N_21508,N_20478);
nor U22272 (N_22272,N_20983,N_21161);
xor U22273 (N_22273,N_20422,N_21266);
or U22274 (N_22274,N_20813,N_20841);
or U22275 (N_22275,N_20419,N_21055);
xnor U22276 (N_22276,N_20443,N_20804);
xor U22277 (N_22277,N_20936,N_20920);
and U22278 (N_22278,N_21594,N_21411);
nand U22279 (N_22279,N_21215,N_21257);
and U22280 (N_22280,N_21335,N_20621);
nor U22281 (N_22281,N_21056,N_21136);
nor U22282 (N_22282,N_20490,N_20910);
xnor U22283 (N_22283,N_21248,N_21212);
xnor U22284 (N_22284,N_21302,N_21041);
and U22285 (N_22285,N_21538,N_20848);
nor U22286 (N_22286,N_21406,N_21033);
or U22287 (N_22287,N_21294,N_20904);
and U22288 (N_22288,N_20493,N_21088);
xor U22289 (N_22289,N_21525,N_20770);
or U22290 (N_22290,N_21222,N_20625);
nand U22291 (N_22291,N_21292,N_21059);
nand U22292 (N_22292,N_21403,N_21188);
or U22293 (N_22293,N_21588,N_21304);
nand U22294 (N_22294,N_21045,N_21048);
or U22295 (N_22295,N_20507,N_21346);
and U22296 (N_22296,N_21341,N_21195);
xor U22297 (N_22297,N_20733,N_20512);
nor U22298 (N_22298,N_21492,N_20569);
nand U22299 (N_22299,N_20549,N_20495);
and U22300 (N_22300,N_21519,N_20499);
xor U22301 (N_22301,N_21553,N_20921);
xnor U22302 (N_22302,N_21211,N_20921);
nand U22303 (N_22303,N_20477,N_20715);
nor U22304 (N_22304,N_21082,N_21536);
and U22305 (N_22305,N_20745,N_21038);
nand U22306 (N_22306,N_20568,N_20646);
nor U22307 (N_22307,N_20712,N_21177);
nand U22308 (N_22308,N_21388,N_21135);
xor U22309 (N_22309,N_20406,N_20809);
nand U22310 (N_22310,N_20443,N_20727);
or U22311 (N_22311,N_21017,N_21505);
nor U22312 (N_22312,N_21294,N_20783);
nand U22313 (N_22313,N_21193,N_21355);
and U22314 (N_22314,N_21276,N_21375);
and U22315 (N_22315,N_20841,N_21141);
nor U22316 (N_22316,N_21160,N_20906);
nand U22317 (N_22317,N_20556,N_20543);
xnor U22318 (N_22318,N_21352,N_20590);
nor U22319 (N_22319,N_21122,N_21121);
xnor U22320 (N_22320,N_20913,N_21055);
or U22321 (N_22321,N_21562,N_21550);
nand U22322 (N_22322,N_20928,N_20898);
nor U22323 (N_22323,N_21124,N_20811);
or U22324 (N_22324,N_20975,N_20678);
nor U22325 (N_22325,N_20867,N_21316);
or U22326 (N_22326,N_21487,N_21200);
or U22327 (N_22327,N_21309,N_20698);
nand U22328 (N_22328,N_20986,N_20965);
xnor U22329 (N_22329,N_20519,N_21594);
nand U22330 (N_22330,N_20875,N_20702);
and U22331 (N_22331,N_20693,N_20704);
nand U22332 (N_22332,N_21336,N_21259);
nor U22333 (N_22333,N_20735,N_21256);
nor U22334 (N_22334,N_21006,N_21150);
and U22335 (N_22335,N_20733,N_20612);
nand U22336 (N_22336,N_20921,N_20814);
nand U22337 (N_22337,N_21502,N_21531);
or U22338 (N_22338,N_20820,N_21208);
xor U22339 (N_22339,N_20752,N_20573);
and U22340 (N_22340,N_20956,N_21354);
nand U22341 (N_22341,N_20459,N_20876);
xor U22342 (N_22342,N_21351,N_20453);
xnor U22343 (N_22343,N_21310,N_20649);
nor U22344 (N_22344,N_20643,N_20884);
nor U22345 (N_22345,N_20493,N_20480);
nor U22346 (N_22346,N_21309,N_20946);
nor U22347 (N_22347,N_21230,N_20674);
nor U22348 (N_22348,N_21262,N_20751);
and U22349 (N_22349,N_21278,N_20653);
and U22350 (N_22350,N_21516,N_20679);
xnor U22351 (N_22351,N_21381,N_21520);
xnor U22352 (N_22352,N_21106,N_20756);
or U22353 (N_22353,N_20454,N_20966);
xor U22354 (N_22354,N_20543,N_21118);
xor U22355 (N_22355,N_21592,N_21362);
nor U22356 (N_22356,N_20769,N_20566);
nand U22357 (N_22357,N_21358,N_21365);
nand U22358 (N_22358,N_21472,N_20741);
xnor U22359 (N_22359,N_20741,N_20627);
or U22360 (N_22360,N_21435,N_20617);
or U22361 (N_22361,N_20418,N_21236);
xnor U22362 (N_22362,N_21517,N_20538);
or U22363 (N_22363,N_21305,N_20855);
xnor U22364 (N_22364,N_21118,N_20884);
and U22365 (N_22365,N_21535,N_20528);
or U22366 (N_22366,N_20443,N_20731);
xor U22367 (N_22367,N_20999,N_20805);
and U22368 (N_22368,N_21137,N_20745);
nor U22369 (N_22369,N_21223,N_20868);
and U22370 (N_22370,N_21000,N_20564);
nand U22371 (N_22371,N_20623,N_20832);
or U22372 (N_22372,N_20951,N_20501);
and U22373 (N_22373,N_20718,N_20803);
or U22374 (N_22374,N_21427,N_21431);
xor U22375 (N_22375,N_20843,N_20593);
xnor U22376 (N_22376,N_20737,N_21257);
xor U22377 (N_22377,N_20497,N_21438);
nand U22378 (N_22378,N_21569,N_21462);
xor U22379 (N_22379,N_20423,N_20975);
nor U22380 (N_22380,N_21534,N_21126);
nand U22381 (N_22381,N_21219,N_20988);
nand U22382 (N_22382,N_21027,N_21203);
xnor U22383 (N_22383,N_20638,N_20760);
or U22384 (N_22384,N_21336,N_20579);
xnor U22385 (N_22385,N_21238,N_20954);
nor U22386 (N_22386,N_21557,N_20931);
nand U22387 (N_22387,N_21460,N_21131);
or U22388 (N_22388,N_20534,N_20577);
xnor U22389 (N_22389,N_20485,N_21284);
nor U22390 (N_22390,N_20820,N_21343);
nand U22391 (N_22391,N_21292,N_20420);
and U22392 (N_22392,N_21232,N_21110);
nor U22393 (N_22393,N_20410,N_21522);
xor U22394 (N_22394,N_20685,N_21410);
nand U22395 (N_22395,N_21183,N_20569);
nor U22396 (N_22396,N_20462,N_20525);
xor U22397 (N_22397,N_20836,N_20633);
xor U22398 (N_22398,N_21444,N_21297);
nand U22399 (N_22399,N_21508,N_20425);
and U22400 (N_22400,N_20792,N_20952);
xor U22401 (N_22401,N_20660,N_20677);
nand U22402 (N_22402,N_21094,N_21472);
nor U22403 (N_22403,N_20599,N_21066);
or U22404 (N_22404,N_20881,N_21586);
or U22405 (N_22405,N_20463,N_20972);
xor U22406 (N_22406,N_21073,N_20520);
and U22407 (N_22407,N_20567,N_20947);
nand U22408 (N_22408,N_21567,N_20427);
and U22409 (N_22409,N_21570,N_21155);
nor U22410 (N_22410,N_21418,N_21353);
nand U22411 (N_22411,N_20880,N_21410);
or U22412 (N_22412,N_20941,N_21417);
nand U22413 (N_22413,N_20439,N_20713);
nor U22414 (N_22414,N_20912,N_20763);
or U22415 (N_22415,N_20733,N_20759);
nor U22416 (N_22416,N_21240,N_21597);
xor U22417 (N_22417,N_20767,N_21440);
nor U22418 (N_22418,N_20634,N_20759);
nor U22419 (N_22419,N_21132,N_21505);
xnor U22420 (N_22420,N_21071,N_21191);
nor U22421 (N_22421,N_21158,N_20416);
nor U22422 (N_22422,N_20562,N_20698);
or U22423 (N_22423,N_20949,N_21027);
nor U22424 (N_22424,N_20587,N_21394);
or U22425 (N_22425,N_21039,N_20882);
nor U22426 (N_22426,N_20829,N_21082);
xnor U22427 (N_22427,N_20784,N_20629);
or U22428 (N_22428,N_21135,N_20752);
nor U22429 (N_22429,N_20785,N_21099);
xor U22430 (N_22430,N_21566,N_21382);
and U22431 (N_22431,N_21406,N_21064);
nand U22432 (N_22432,N_21110,N_20684);
nor U22433 (N_22433,N_20615,N_20753);
or U22434 (N_22434,N_21042,N_21067);
or U22435 (N_22435,N_20790,N_20868);
nand U22436 (N_22436,N_21067,N_21397);
or U22437 (N_22437,N_21343,N_20972);
nand U22438 (N_22438,N_20814,N_21069);
nor U22439 (N_22439,N_21234,N_21172);
or U22440 (N_22440,N_21223,N_20756);
or U22441 (N_22441,N_21307,N_20784);
xnor U22442 (N_22442,N_21060,N_20519);
and U22443 (N_22443,N_21410,N_20456);
nor U22444 (N_22444,N_20701,N_21292);
nor U22445 (N_22445,N_20906,N_20885);
nand U22446 (N_22446,N_20990,N_21501);
or U22447 (N_22447,N_21182,N_21458);
and U22448 (N_22448,N_21091,N_21311);
nor U22449 (N_22449,N_21578,N_21206);
and U22450 (N_22450,N_21554,N_21031);
or U22451 (N_22451,N_21094,N_21004);
xor U22452 (N_22452,N_21462,N_21094);
or U22453 (N_22453,N_20607,N_21044);
or U22454 (N_22454,N_20930,N_21252);
nand U22455 (N_22455,N_20555,N_21494);
nand U22456 (N_22456,N_21433,N_21359);
xnor U22457 (N_22457,N_21344,N_20445);
nand U22458 (N_22458,N_20975,N_20920);
or U22459 (N_22459,N_20777,N_20833);
and U22460 (N_22460,N_21348,N_20738);
nor U22461 (N_22461,N_21551,N_20813);
and U22462 (N_22462,N_21183,N_21447);
nor U22463 (N_22463,N_20783,N_21085);
and U22464 (N_22464,N_20456,N_21389);
nand U22465 (N_22465,N_20769,N_20804);
and U22466 (N_22466,N_21392,N_20489);
xnor U22467 (N_22467,N_20486,N_20835);
nor U22468 (N_22468,N_21292,N_20555);
xor U22469 (N_22469,N_21569,N_21359);
nor U22470 (N_22470,N_21180,N_20839);
nor U22471 (N_22471,N_20631,N_20957);
nor U22472 (N_22472,N_21512,N_20685);
nor U22473 (N_22473,N_20912,N_21154);
xor U22474 (N_22474,N_21217,N_20670);
nor U22475 (N_22475,N_20810,N_20552);
and U22476 (N_22476,N_20791,N_21310);
nor U22477 (N_22477,N_21036,N_21336);
or U22478 (N_22478,N_21306,N_21212);
or U22479 (N_22479,N_21187,N_20455);
nor U22480 (N_22480,N_21369,N_20421);
xnor U22481 (N_22481,N_21116,N_21167);
nor U22482 (N_22482,N_21591,N_20403);
nor U22483 (N_22483,N_20885,N_20560);
xnor U22484 (N_22484,N_21171,N_20617);
nand U22485 (N_22485,N_20547,N_20701);
and U22486 (N_22486,N_20575,N_21459);
nand U22487 (N_22487,N_20407,N_21511);
xnor U22488 (N_22488,N_21516,N_21223);
nor U22489 (N_22489,N_20772,N_20870);
nor U22490 (N_22490,N_20478,N_20518);
nand U22491 (N_22491,N_21160,N_21029);
or U22492 (N_22492,N_20722,N_20451);
nand U22493 (N_22493,N_21299,N_20694);
nor U22494 (N_22494,N_20714,N_20475);
or U22495 (N_22495,N_21535,N_21404);
nand U22496 (N_22496,N_20630,N_21571);
and U22497 (N_22497,N_20967,N_21213);
nor U22498 (N_22498,N_20797,N_21534);
nor U22499 (N_22499,N_20705,N_21562);
nor U22500 (N_22500,N_21207,N_20766);
and U22501 (N_22501,N_20853,N_20577);
nand U22502 (N_22502,N_20414,N_20942);
nor U22503 (N_22503,N_20871,N_21394);
and U22504 (N_22504,N_21326,N_21134);
nand U22505 (N_22505,N_20617,N_20808);
nand U22506 (N_22506,N_20565,N_20647);
and U22507 (N_22507,N_20623,N_21545);
xor U22508 (N_22508,N_21582,N_21521);
xnor U22509 (N_22509,N_21012,N_21065);
nand U22510 (N_22510,N_20711,N_21507);
xnor U22511 (N_22511,N_21588,N_21042);
xor U22512 (N_22512,N_21112,N_21030);
nand U22513 (N_22513,N_21577,N_20521);
nor U22514 (N_22514,N_21133,N_21311);
and U22515 (N_22515,N_21025,N_20553);
nand U22516 (N_22516,N_20807,N_21048);
or U22517 (N_22517,N_21521,N_20582);
and U22518 (N_22518,N_21275,N_20525);
nor U22519 (N_22519,N_21020,N_21214);
and U22520 (N_22520,N_21503,N_21048);
nand U22521 (N_22521,N_21519,N_20697);
and U22522 (N_22522,N_20636,N_21071);
or U22523 (N_22523,N_20594,N_21566);
nor U22524 (N_22524,N_20832,N_20478);
nor U22525 (N_22525,N_21156,N_21571);
or U22526 (N_22526,N_20642,N_20427);
or U22527 (N_22527,N_20463,N_21260);
nand U22528 (N_22528,N_20899,N_21375);
nand U22529 (N_22529,N_21091,N_20505);
or U22530 (N_22530,N_21325,N_21518);
and U22531 (N_22531,N_21200,N_20976);
nor U22532 (N_22532,N_21096,N_20400);
xor U22533 (N_22533,N_20910,N_21538);
xnor U22534 (N_22534,N_20744,N_20854);
xor U22535 (N_22535,N_21314,N_20881);
and U22536 (N_22536,N_20537,N_20697);
nor U22537 (N_22537,N_21233,N_21047);
or U22538 (N_22538,N_21167,N_20464);
nor U22539 (N_22539,N_21240,N_20584);
xor U22540 (N_22540,N_20649,N_20765);
nor U22541 (N_22541,N_20510,N_21383);
and U22542 (N_22542,N_21038,N_20817);
nand U22543 (N_22543,N_20977,N_20705);
nand U22544 (N_22544,N_20411,N_20739);
nand U22545 (N_22545,N_20684,N_20614);
nand U22546 (N_22546,N_20415,N_20998);
and U22547 (N_22547,N_20456,N_21509);
xnor U22548 (N_22548,N_20898,N_21202);
and U22549 (N_22549,N_21055,N_21301);
and U22550 (N_22550,N_20851,N_20470);
xnor U22551 (N_22551,N_21148,N_20401);
or U22552 (N_22552,N_20750,N_21546);
nor U22553 (N_22553,N_21587,N_21516);
or U22554 (N_22554,N_21158,N_21326);
or U22555 (N_22555,N_21032,N_20478);
nor U22556 (N_22556,N_20851,N_20471);
xnor U22557 (N_22557,N_20674,N_21273);
nand U22558 (N_22558,N_21332,N_21202);
nand U22559 (N_22559,N_20927,N_20779);
nor U22560 (N_22560,N_20825,N_21220);
nor U22561 (N_22561,N_20714,N_20986);
and U22562 (N_22562,N_21590,N_20905);
nor U22563 (N_22563,N_21059,N_20504);
and U22564 (N_22564,N_20994,N_21450);
nand U22565 (N_22565,N_21143,N_21338);
xor U22566 (N_22566,N_20543,N_21076);
xnor U22567 (N_22567,N_20993,N_20422);
nand U22568 (N_22568,N_20755,N_21358);
nand U22569 (N_22569,N_21575,N_20824);
nand U22570 (N_22570,N_21302,N_21165);
nor U22571 (N_22571,N_20837,N_21576);
nor U22572 (N_22572,N_20777,N_20951);
or U22573 (N_22573,N_21250,N_20704);
or U22574 (N_22574,N_21387,N_21217);
xor U22575 (N_22575,N_21205,N_20402);
nand U22576 (N_22576,N_21066,N_20698);
and U22577 (N_22577,N_20747,N_21125);
and U22578 (N_22578,N_21171,N_21403);
nand U22579 (N_22579,N_20807,N_21517);
and U22580 (N_22580,N_20553,N_21391);
nor U22581 (N_22581,N_21113,N_21215);
or U22582 (N_22582,N_20681,N_21437);
or U22583 (N_22583,N_21185,N_20944);
and U22584 (N_22584,N_20888,N_21323);
nor U22585 (N_22585,N_20861,N_21409);
nor U22586 (N_22586,N_20894,N_20521);
xnor U22587 (N_22587,N_20916,N_21326);
nor U22588 (N_22588,N_21166,N_21153);
and U22589 (N_22589,N_20779,N_21490);
and U22590 (N_22590,N_21353,N_20407);
nand U22591 (N_22591,N_20854,N_20717);
or U22592 (N_22592,N_20717,N_20583);
or U22593 (N_22593,N_21590,N_20585);
and U22594 (N_22594,N_21473,N_20645);
and U22595 (N_22595,N_20909,N_20627);
nand U22596 (N_22596,N_20432,N_20463);
and U22597 (N_22597,N_20873,N_20905);
xnor U22598 (N_22598,N_20908,N_21573);
xnor U22599 (N_22599,N_20820,N_20429);
or U22600 (N_22600,N_21321,N_21535);
nor U22601 (N_22601,N_20865,N_21290);
and U22602 (N_22602,N_21201,N_21062);
and U22603 (N_22603,N_20585,N_21320);
nand U22604 (N_22604,N_21100,N_21144);
xnor U22605 (N_22605,N_21196,N_20817);
xor U22606 (N_22606,N_20837,N_20987);
nand U22607 (N_22607,N_21139,N_21195);
and U22608 (N_22608,N_21332,N_21492);
and U22609 (N_22609,N_20511,N_20433);
or U22610 (N_22610,N_21067,N_21491);
xnor U22611 (N_22611,N_21215,N_20761);
or U22612 (N_22612,N_21254,N_21058);
or U22613 (N_22613,N_20460,N_20774);
nor U22614 (N_22614,N_20945,N_21296);
nor U22615 (N_22615,N_21347,N_21130);
xnor U22616 (N_22616,N_20547,N_20551);
nand U22617 (N_22617,N_21481,N_20652);
nand U22618 (N_22618,N_20722,N_20736);
xor U22619 (N_22619,N_21064,N_21132);
nand U22620 (N_22620,N_20587,N_21462);
or U22621 (N_22621,N_20973,N_20746);
or U22622 (N_22622,N_21207,N_20932);
or U22623 (N_22623,N_20427,N_21219);
nor U22624 (N_22624,N_20936,N_21350);
nand U22625 (N_22625,N_20705,N_20653);
nand U22626 (N_22626,N_20452,N_20898);
or U22627 (N_22627,N_20433,N_21527);
nand U22628 (N_22628,N_20885,N_21059);
or U22629 (N_22629,N_21188,N_20760);
and U22630 (N_22630,N_21320,N_20928);
nand U22631 (N_22631,N_20845,N_21215);
nand U22632 (N_22632,N_21220,N_21569);
nor U22633 (N_22633,N_20647,N_21563);
or U22634 (N_22634,N_20557,N_21063);
and U22635 (N_22635,N_21340,N_20589);
and U22636 (N_22636,N_21187,N_20874);
nor U22637 (N_22637,N_20574,N_21212);
and U22638 (N_22638,N_20885,N_21107);
and U22639 (N_22639,N_20634,N_21550);
xor U22640 (N_22640,N_21238,N_21440);
or U22641 (N_22641,N_20801,N_21427);
and U22642 (N_22642,N_21566,N_21544);
or U22643 (N_22643,N_20847,N_20621);
xor U22644 (N_22644,N_20835,N_21397);
and U22645 (N_22645,N_21330,N_20443);
nor U22646 (N_22646,N_21292,N_20971);
nand U22647 (N_22647,N_20893,N_20411);
or U22648 (N_22648,N_20854,N_21360);
xor U22649 (N_22649,N_21561,N_20958);
and U22650 (N_22650,N_20549,N_21384);
and U22651 (N_22651,N_21261,N_20692);
nor U22652 (N_22652,N_21456,N_21495);
nor U22653 (N_22653,N_21094,N_21282);
xnor U22654 (N_22654,N_21310,N_21231);
nand U22655 (N_22655,N_21595,N_21213);
and U22656 (N_22656,N_21165,N_21213);
or U22657 (N_22657,N_21087,N_20916);
xnor U22658 (N_22658,N_20432,N_21032);
or U22659 (N_22659,N_20459,N_20410);
xor U22660 (N_22660,N_21037,N_21218);
or U22661 (N_22661,N_21180,N_21264);
xor U22662 (N_22662,N_20824,N_21540);
and U22663 (N_22663,N_21289,N_20479);
or U22664 (N_22664,N_21400,N_21352);
nand U22665 (N_22665,N_21045,N_21070);
xnor U22666 (N_22666,N_21110,N_21295);
or U22667 (N_22667,N_21434,N_21121);
and U22668 (N_22668,N_20752,N_20851);
xor U22669 (N_22669,N_21187,N_21521);
xnor U22670 (N_22670,N_20902,N_20591);
and U22671 (N_22671,N_21377,N_20508);
nand U22672 (N_22672,N_21489,N_21334);
xor U22673 (N_22673,N_20476,N_21066);
nor U22674 (N_22674,N_21373,N_21183);
or U22675 (N_22675,N_21013,N_21433);
xnor U22676 (N_22676,N_20690,N_20797);
or U22677 (N_22677,N_21058,N_20740);
and U22678 (N_22678,N_21354,N_21404);
xor U22679 (N_22679,N_20975,N_20924);
xnor U22680 (N_22680,N_20960,N_21074);
and U22681 (N_22681,N_21058,N_21180);
nor U22682 (N_22682,N_21394,N_20531);
nand U22683 (N_22683,N_20839,N_20841);
or U22684 (N_22684,N_20615,N_21512);
and U22685 (N_22685,N_21545,N_21445);
and U22686 (N_22686,N_21193,N_20734);
and U22687 (N_22687,N_21387,N_20528);
and U22688 (N_22688,N_21344,N_20810);
nand U22689 (N_22689,N_20685,N_20752);
xor U22690 (N_22690,N_20995,N_20771);
nand U22691 (N_22691,N_21130,N_20693);
nand U22692 (N_22692,N_20608,N_21081);
nand U22693 (N_22693,N_21400,N_20656);
xnor U22694 (N_22694,N_20886,N_21463);
or U22695 (N_22695,N_21141,N_20706);
or U22696 (N_22696,N_20864,N_20881);
and U22697 (N_22697,N_20547,N_20852);
or U22698 (N_22698,N_21449,N_21218);
or U22699 (N_22699,N_20826,N_21238);
xor U22700 (N_22700,N_20405,N_20594);
xor U22701 (N_22701,N_21342,N_21539);
nand U22702 (N_22702,N_21061,N_21478);
xor U22703 (N_22703,N_20806,N_21183);
or U22704 (N_22704,N_20498,N_21258);
nor U22705 (N_22705,N_21138,N_21333);
nand U22706 (N_22706,N_20409,N_20661);
xor U22707 (N_22707,N_20748,N_20953);
and U22708 (N_22708,N_20716,N_20456);
nor U22709 (N_22709,N_20904,N_21452);
or U22710 (N_22710,N_21478,N_21593);
nand U22711 (N_22711,N_21135,N_20455);
nand U22712 (N_22712,N_20653,N_20947);
or U22713 (N_22713,N_20743,N_20829);
nand U22714 (N_22714,N_21089,N_21452);
or U22715 (N_22715,N_21536,N_20775);
and U22716 (N_22716,N_21481,N_20662);
xor U22717 (N_22717,N_20956,N_21593);
nand U22718 (N_22718,N_20734,N_20465);
xor U22719 (N_22719,N_20970,N_20553);
and U22720 (N_22720,N_21520,N_20607);
nand U22721 (N_22721,N_20955,N_21533);
nand U22722 (N_22722,N_20587,N_20952);
or U22723 (N_22723,N_21262,N_20948);
or U22724 (N_22724,N_21260,N_20862);
nand U22725 (N_22725,N_20886,N_20670);
and U22726 (N_22726,N_21546,N_20882);
or U22727 (N_22727,N_20419,N_21266);
and U22728 (N_22728,N_20682,N_21009);
nor U22729 (N_22729,N_20862,N_21444);
nor U22730 (N_22730,N_20992,N_20984);
xor U22731 (N_22731,N_20584,N_21281);
and U22732 (N_22732,N_21493,N_20477);
and U22733 (N_22733,N_20411,N_21115);
or U22734 (N_22734,N_20670,N_20917);
nor U22735 (N_22735,N_20495,N_20579);
nor U22736 (N_22736,N_20993,N_20806);
nand U22737 (N_22737,N_21520,N_20749);
and U22738 (N_22738,N_21416,N_21057);
nor U22739 (N_22739,N_20777,N_20802);
nand U22740 (N_22740,N_20816,N_21596);
nor U22741 (N_22741,N_21498,N_20918);
or U22742 (N_22742,N_21336,N_21086);
or U22743 (N_22743,N_21043,N_21137);
xor U22744 (N_22744,N_20505,N_21075);
nand U22745 (N_22745,N_20540,N_20756);
nor U22746 (N_22746,N_20773,N_20924);
nand U22747 (N_22747,N_21034,N_21406);
or U22748 (N_22748,N_21538,N_20922);
nand U22749 (N_22749,N_20566,N_21571);
or U22750 (N_22750,N_20560,N_21571);
nand U22751 (N_22751,N_20632,N_21531);
nand U22752 (N_22752,N_20841,N_21190);
nand U22753 (N_22753,N_20822,N_20531);
xnor U22754 (N_22754,N_20551,N_21599);
xor U22755 (N_22755,N_20697,N_20938);
nand U22756 (N_22756,N_21490,N_20419);
nor U22757 (N_22757,N_20990,N_21291);
nor U22758 (N_22758,N_20980,N_20929);
and U22759 (N_22759,N_20739,N_21153);
nor U22760 (N_22760,N_21251,N_21127);
xor U22761 (N_22761,N_20964,N_20453);
and U22762 (N_22762,N_21073,N_21056);
nand U22763 (N_22763,N_21095,N_21504);
nor U22764 (N_22764,N_21424,N_21453);
and U22765 (N_22765,N_21042,N_21188);
nor U22766 (N_22766,N_21450,N_20621);
nand U22767 (N_22767,N_21148,N_21031);
xor U22768 (N_22768,N_21425,N_20663);
nand U22769 (N_22769,N_21436,N_20769);
xor U22770 (N_22770,N_21293,N_20705);
or U22771 (N_22771,N_21231,N_20638);
xor U22772 (N_22772,N_21578,N_20930);
nor U22773 (N_22773,N_21468,N_21031);
or U22774 (N_22774,N_20515,N_20997);
and U22775 (N_22775,N_20641,N_20423);
and U22776 (N_22776,N_21203,N_21060);
nand U22777 (N_22777,N_21199,N_21219);
xor U22778 (N_22778,N_20562,N_21332);
nor U22779 (N_22779,N_20604,N_21406);
nor U22780 (N_22780,N_20976,N_20604);
xor U22781 (N_22781,N_20764,N_20740);
nor U22782 (N_22782,N_21379,N_20912);
or U22783 (N_22783,N_21446,N_21297);
xnor U22784 (N_22784,N_20718,N_21202);
nand U22785 (N_22785,N_20676,N_20859);
nor U22786 (N_22786,N_20776,N_20411);
and U22787 (N_22787,N_20803,N_20795);
or U22788 (N_22788,N_20773,N_21240);
nand U22789 (N_22789,N_20742,N_20980);
nor U22790 (N_22790,N_21137,N_21543);
nor U22791 (N_22791,N_21546,N_20898);
and U22792 (N_22792,N_21508,N_20957);
nor U22793 (N_22793,N_20446,N_21250);
xor U22794 (N_22794,N_21134,N_20482);
nand U22795 (N_22795,N_21141,N_20897);
nand U22796 (N_22796,N_20945,N_20693);
or U22797 (N_22797,N_20593,N_20518);
or U22798 (N_22798,N_21399,N_20974);
or U22799 (N_22799,N_20845,N_20664);
or U22800 (N_22800,N_22253,N_21754);
nand U22801 (N_22801,N_22069,N_22372);
or U22802 (N_22802,N_21888,N_22721);
nor U22803 (N_22803,N_22529,N_22118);
and U22804 (N_22804,N_21820,N_22186);
xnor U22805 (N_22805,N_21833,N_21895);
nand U22806 (N_22806,N_22342,N_22267);
xnor U22807 (N_22807,N_21899,N_22676);
nand U22808 (N_22808,N_21817,N_22214);
nand U22809 (N_22809,N_22475,N_22123);
and U22810 (N_22810,N_22140,N_22446);
nor U22811 (N_22811,N_22579,N_22737);
nor U22812 (N_22812,N_22039,N_22428);
nor U22813 (N_22813,N_22405,N_22463);
nand U22814 (N_22814,N_22127,N_21733);
nand U22815 (N_22815,N_22569,N_22301);
xor U22816 (N_22816,N_21887,N_22340);
nand U22817 (N_22817,N_22431,N_22504);
nand U22818 (N_22818,N_21779,N_21898);
nor U22819 (N_22819,N_22448,N_22541);
nand U22820 (N_22820,N_22568,N_22600);
and U22821 (N_22821,N_21753,N_21613);
nand U22822 (N_22822,N_22153,N_22499);
or U22823 (N_22823,N_21800,N_21974);
or U22824 (N_22824,N_22205,N_22731);
nand U22825 (N_22825,N_21710,N_22485);
xnor U22826 (N_22826,N_21855,N_22400);
nor U22827 (N_22827,N_22430,N_21691);
and U22828 (N_22828,N_22029,N_22723);
and U22829 (N_22829,N_22699,N_22018);
or U22830 (N_22830,N_21614,N_21845);
nand U22831 (N_22831,N_22521,N_22285);
nor U22832 (N_22832,N_22654,N_22658);
or U22833 (N_22833,N_22193,N_22451);
nand U22834 (N_22834,N_22596,N_22407);
nand U22835 (N_22835,N_22549,N_22108);
and U22836 (N_22836,N_22173,N_21826);
or U22837 (N_22837,N_22082,N_22065);
nand U22838 (N_22838,N_21901,N_21958);
nand U22839 (N_22839,N_22727,N_21952);
nor U22840 (N_22840,N_21813,N_22129);
xnor U22841 (N_22841,N_22365,N_22518);
and U22842 (N_22842,N_22696,N_21853);
nor U22843 (N_22843,N_22093,N_22537);
nor U22844 (N_22844,N_22413,N_22182);
nor U22845 (N_22845,N_22197,N_22750);
xnor U22846 (N_22846,N_22777,N_22782);
nor U22847 (N_22847,N_22177,N_21795);
xor U22848 (N_22848,N_22701,N_22606);
nor U22849 (N_22849,N_22771,N_22590);
and U22850 (N_22850,N_22617,N_22289);
or U22851 (N_22851,N_22785,N_22345);
xnor U22852 (N_22852,N_21724,N_22509);
or U22853 (N_22853,N_21831,N_22300);
nand U22854 (N_22854,N_21949,N_21842);
and U22855 (N_22855,N_22211,N_22359);
or U22856 (N_22856,N_22415,N_21657);
nand U22857 (N_22857,N_22057,N_22049);
and U22858 (N_22858,N_22068,N_22061);
nand U22859 (N_22859,N_21970,N_22382);
or U22860 (N_22860,N_21784,N_22574);
and U22861 (N_22861,N_22735,N_22126);
nand U22862 (N_22862,N_22483,N_22510);
and U22863 (N_22863,N_21967,N_22674);
nor U22864 (N_22864,N_22292,N_22507);
xor U22865 (N_22865,N_22150,N_22634);
xnor U22866 (N_22866,N_22328,N_22505);
nand U22867 (N_22867,N_21619,N_22387);
xor U22868 (N_22868,N_22531,N_22477);
xor U22869 (N_22869,N_21882,N_22604);
nor U22870 (N_22870,N_21607,N_21893);
xnor U22871 (N_22871,N_22054,N_22511);
or U22872 (N_22872,N_21803,N_22402);
or U22873 (N_22873,N_22255,N_22031);
or U22874 (N_22874,N_22035,N_21760);
nand U22875 (N_22875,N_22670,N_21656);
or U22876 (N_22876,N_21781,N_22225);
xor U22877 (N_22877,N_21715,N_21945);
nand U22878 (N_22878,N_22200,N_21675);
nand U22879 (N_22879,N_22074,N_22168);
nand U22880 (N_22880,N_22545,N_22616);
nand U22881 (N_22881,N_21641,N_22046);
nor U22882 (N_22882,N_22482,N_22624);
and U22883 (N_22883,N_22156,N_21862);
or U22884 (N_22884,N_22138,N_22673);
or U22885 (N_22885,N_22661,N_22429);
xnor U22886 (N_22886,N_22189,N_21809);
nand U22887 (N_22887,N_21909,N_21615);
nor U22888 (N_22888,N_22135,N_22277);
or U22889 (N_22889,N_21763,N_22154);
nor U22890 (N_22890,N_22730,N_22075);
nor U22891 (N_22891,N_22651,N_22744);
or U22892 (N_22892,N_22041,N_22611);
xnor U22893 (N_22893,N_21667,N_22274);
or U22894 (N_22894,N_22199,N_22646);
nand U22895 (N_22895,N_22757,N_22103);
or U22896 (N_22896,N_22139,N_21964);
or U22897 (N_22897,N_22224,N_22412);
nor U22898 (N_22898,N_21943,N_22663);
nor U22899 (N_22899,N_21627,N_21937);
xnor U22900 (N_22900,N_22178,N_21783);
xnor U22901 (N_22901,N_22265,N_21962);
and U22902 (N_22902,N_21906,N_21929);
xor U22903 (N_22903,N_22618,N_22249);
and U22904 (N_22904,N_22597,N_22439);
nor U22905 (N_22905,N_21912,N_22733);
nand U22906 (N_22906,N_22263,N_22652);
nand U22907 (N_22907,N_21734,N_21677);
nor U22908 (N_22908,N_22572,N_21844);
nand U22909 (N_22909,N_21985,N_22761);
or U22910 (N_22910,N_22272,N_21757);
or U22911 (N_22911,N_22621,N_21666);
nand U22912 (N_22912,N_22738,N_22036);
and U22913 (N_22913,N_22498,N_22546);
xnor U22914 (N_22914,N_22554,N_22517);
xor U22915 (N_22915,N_22566,N_22467);
xor U22916 (N_22916,N_22079,N_22377);
or U22917 (N_22917,N_21915,N_22134);
xnor U22918 (N_22918,N_21850,N_22087);
xor U22919 (N_22919,N_22598,N_22608);
xor U22920 (N_22920,N_22005,N_21664);
or U22921 (N_22921,N_22076,N_22337);
nand U22922 (N_22922,N_21731,N_21746);
xnor U22923 (N_22923,N_21730,N_22719);
or U22924 (N_22924,N_22141,N_22742);
nor U22925 (N_22925,N_21684,N_22729);
nor U22926 (N_22926,N_22014,N_22097);
or U22927 (N_22927,N_22112,N_21606);
nand U22928 (N_22928,N_22081,N_22148);
or U22929 (N_22929,N_21859,N_21794);
nor U22930 (N_22930,N_22725,N_21647);
nor U22931 (N_22931,N_21665,N_22464);
and U22932 (N_22932,N_22688,N_22707);
nand U22933 (N_22933,N_21628,N_22749);
nand U22934 (N_22934,N_21774,N_22760);
nand U22935 (N_22935,N_22424,N_22739);
or U22936 (N_22936,N_22789,N_22091);
nand U22937 (N_22937,N_21861,N_21840);
xnor U22938 (N_22938,N_22408,N_21884);
nand U22939 (N_22939,N_22680,N_21714);
nor U22940 (N_22940,N_22346,N_22060);
xnor U22941 (N_22941,N_21905,N_22470);
nand U22942 (N_22942,N_22171,N_22686);
nand U22943 (N_22943,N_22349,N_21732);
and U22944 (N_22944,N_22512,N_22716);
xor U22945 (N_22945,N_22032,N_22694);
nor U22946 (N_22946,N_21998,N_22333);
xor U22947 (N_22947,N_21834,N_22548);
nand U22948 (N_22948,N_21908,N_22573);
or U22949 (N_22949,N_22151,N_22648);
nor U22950 (N_22950,N_21877,N_21860);
nor U22951 (N_22951,N_21863,N_22383);
xor U22952 (N_22952,N_22350,N_22145);
nand U22953 (N_22953,N_22086,N_22288);
xor U22954 (N_22954,N_22105,N_22790);
nor U22955 (N_22955,N_21631,N_21719);
nand U22956 (N_22956,N_21776,N_22259);
or U22957 (N_22957,N_21810,N_21749);
and U22958 (N_22958,N_21913,N_22244);
or U22959 (N_22959,N_22258,N_22612);
xor U22960 (N_22960,N_22672,N_22276);
nand U22961 (N_22961,N_22660,N_22453);
and U22962 (N_22962,N_22714,N_22264);
xnor U22963 (N_22963,N_22266,N_22275);
and U22964 (N_22964,N_22011,N_21917);
nor U22965 (N_22965,N_22454,N_21701);
and U22966 (N_22966,N_21990,N_22309);
or U22967 (N_22967,N_21727,N_22639);
and U22968 (N_22968,N_21683,N_21654);
nor U22969 (N_22969,N_22117,N_22291);
xnor U22970 (N_22970,N_22325,N_21920);
xnor U22971 (N_22971,N_21679,N_22500);
nor U22972 (N_22972,N_22360,N_22229);
and U22973 (N_22973,N_21758,N_22513);
nand U22974 (N_22974,N_22551,N_22395);
xor U22975 (N_22975,N_22305,N_22284);
and U22976 (N_22976,N_22491,N_22710);
xor U22977 (N_22977,N_22709,N_21982);
and U22978 (N_22978,N_22717,N_22004);
nand U22979 (N_22979,N_22157,N_22756);
nor U22980 (N_22980,N_22779,N_22653);
and U22981 (N_22981,N_22316,N_22198);
nand U22982 (N_22982,N_21708,N_22533);
and U22983 (N_22983,N_22209,N_21989);
xor U22984 (N_22984,N_22434,N_21938);
nor U22985 (N_22985,N_21707,N_22559);
nand U22986 (N_22986,N_21942,N_21827);
or U22987 (N_22987,N_22002,N_21694);
nor U22988 (N_22988,N_21873,N_21875);
nor U22989 (N_22989,N_22250,N_21680);
nor U22990 (N_22990,N_22798,N_22550);
nor U22991 (N_22991,N_22524,N_21856);
nand U22992 (N_22992,N_22218,N_22636);
nand U22993 (N_22993,N_22702,N_21668);
and U22994 (N_22994,N_22480,N_21977);
xor U22995 (N_22995,N_22191,N_21788);
nor U22996 (N_22996,N_22233,N_22013);
and U22997 (N_22997,N_22746,N_21816);
and U22998 (N_22998,N_22104,N_21866);
nand U22999 (N_22999,N_22064,N_22167);
xor U23000 (N_23000,N_21698,N_22073);
nand U23001 (N_23001,N_22147,N_21818);
nor U23002 (N_23002,N_21921,N_22166);
nor U23003 (N_23003,N_22599,N_22242);
nand U23004 (N_23004,N_21897,N_22023);
and U23005 (N_23005,N_22689,N_22063);
xnor U23006 (N_23006,N_22748,N_22366);
nand U23007 (N_23007,N_22114,N_21980);
xor U23008 (N_23008,N_22764,N_22762);
and U23009 (N_23009,N_21644,N_22208);
nand U23010 (N_23010,N_22247,N_22560);
nand U23011 (N_23011,N_22149,N_22356);
nor U23012 (N_23012,N_22071,N_21930);
nor U23013 (N_23013,N_22037,N_22235);
and U23014 (N_23014,N_21926,N_22295);
or U23015 (N_23015,N_22206,N_22799);
nand U23016 (N_23016,N_21965,N_22184);
xnor U23017 (N_23017,N_22256,N_22718);
and U23018 (N_23018,N_21717,N_21704);
and U23019 (N_23019,N_22027,N_22028);
or U23020 (N_23020,N_22313,N_22327);
or U23021 (N_23021,N_22332,N_22787);
or U23022 (N_23022,N_22297,N_22195);
or U23023 (N_23023,N_22704,N_22090);
nor U23024 (N_23024,N_22558,N_22122);
or U23025 (N_23025,N_22298,N_21690);
nand U23026 (N_23026,N_22115,N_22170);
and U23027 (N_23027,N_22099,N_22347);
nor U23028 (N_23028,N_22666,N_21904);
nor U23029 (N_23029,N_21652,N_21601);
nand U23030 (N_23030,N_22240,N_21934);
nand U23031 (N_23031,N_22210,N_22338);
nor U23032 (N_23032,N_22113,N_21892);
nand U23033 (N_23033,N_22238,N_22752);
nand U23034 (N_23034,N_22444,N_21723);
nand U23035 (N_23035,N_22629,N_21655);
nand U23036 (N_23036,N_22774,N_22472);
nand U23037 (N_23037,N_22784,N_21973);
nand U23038 (N_23038,N_21660,N_21700);
and U23039 (N_23039,N_21610,N_22675);
xor U23040 (N_23040,N_22271,N_22755);
and U23041 (N_23041,N_22581,N_22404);
and U23042 (N_23042,N_21725,N_21736);
and U23043 (N_23043,N_21849,N_21716);
xnor U23044 (N_23044,N_22589,N_22681);
nor U23045 (N_23045,N_22192,N_22237);
xor U23046 (N_23046,N_22506,N_21622);
or U23047 (N_23047,N_22445,N_22136);
nand U23048 (N_23048,N_22098,N_22243);
or U23049 (N_23049,N_21630,N_21750);
xor U23050 (N_23050,N_22286,N_22695);
nand U23051 (N_23051,N_22715,N_21857);
or U23052 (N_23052,N_22066,N_21771);
and U23053 (N_23053,N_21948,N_21832);
or U23054 (N_23054,N_22732,N_22522);
or U23055 (N_23055,N_21720,N_22106);
and U23056 (N_23056,N_22741,N_22133);
and U23057 (N_23057,N_21772,N_21624);
xor U23058 (N_23058,N_21739,N_22768);
xnor U23059 (N_23059,N_21959,N_21709);
nor U23060 (N_23060,N_21991,N_22318);
nor U23061 (N_23061,N_22204,N_21659);
or U23062 (N_23062,N_21748,N_22364);
nand U23063 (N_23063,N_22311,N_22792);
xor U23064 (N_23064,N_22003,N_22547);
xnor U23065 (N_23065,N_21648,N_22435);
and U23066 (N_23066,N_22664,N_22322);
and U23067 (N_23067,N_21636,N_22223);
xor U23068 (N_23068,N_22495,N_22623);
nor U23069 (N_23069,N_22376,N_22519);
and U23070 (N_23070,N_21954,N_22146);
and U23071 (N_23071,N_22261,N_21759);
nand U23072 (N_23072,N_22423,N_22362);
xnor U23073 (N_23073,N_22226,N_22765);
nor U23074 (N_23074,N_21940,N_22283);
nand U23075 (N_23075,N_22001,N_22232);
nand U23076 (N_23076,N_22780,N_21986);
or U23077 (N_23077,N_22268,N_22181);
nand U23078 (N_23078,N_21812,N_22307);
nor U23079 (N_23079,N_22503,N_22588);
and U23080 (N_23080,N_21824,N_21806);
nor U23081 (N_23081,N_22024,N_22484);
nor U23082 (N_23082,N_21927,N_22698);
or U23083 (N_23083,N_22645,N_21638);
xor U23084 (N_23084,N_22317,N_22578);
xnor U23085 (N_23085,N_22239,N_22532);
nand U23086 (N_23086,N_22058,N_21852);
or U23087 (N_23087,N_22033,N_22647);
nor U23088 (N_23088,N_22137,N_21916);
or U23089 (N_23089,N_22438,N_22143);
xor U23090 (N_23090,N_22441,N_21928);
nor U23091 (N_23091,N_21941,N_22713);
nand U23092 (N_23092,N_21799,N_22794);
or U23093 (N_23093,N_22062,N_22523);
and U23094 (N_23094,N_22493,N_22330);
nand U23095 (N_23095,N_22034,N_21639);
and U23096 (N_23096,N_21947,N_22452);
nor U23097 (N_23097,N_22323,N_21765);
nor U23098 (N_23098,N_21987,N_21747);
or U23099 (N_23099,N_21984,N_22326);
and U23100 (N_23100,N_21600,N_22474);
xor U23101 (N_23101,N_21874,N_22685);
xor U23102 (N_23102,N_21713,N_22396);
nor U23103 (N_23103,N_21837,N_22577);
xor U23104 (N_23104,N_22657,N_21769);
and U23105 (N_23105,N_21787,N_21919);
nor U23106 (N_23106,N_21718,N_21871);
or U23107 (N_23107,N_21963,N_21983);
nand U23108 (N_23108,N_22655,N_22466);
nor U23109 (N_23109,N_22190,N_22254);
xnor U23110 (N_23110,N_22697,N_22659);
nand U23111 (N_23111,N_22595,N_22691);
xor U23112 (N_23112,N_22007,N_21914);
nand U23113 (N_23113,N_21918,N_22460);
xnor U23114 (N_23114,N_22385,N_22393);
or U23115 (N_23115,N_22165,N_22469);
nor U23116 (N_23116,N_22273,N_22626);
nand U23117 (N_23117,N_21711,N_22743);
nand U23118 (N_23118,N_21629,N_21618);
and U23119 (N_23119,N_21876,N_22684);
and U23120 (N_23120,N_21706,N_22020);
nand U23121 (N_23121,N_22067,N_22745);
nor U23122 (N_23122,N_22754,N_22770);
and U23123 (N_23123,N_21865,N_22488);
and U23124 (N_23124,N_21752,N_22728);
and U23125 (N_23125,N_21858,N_22095);
and U23126 (N_23126,N_22048,N_21685);
and U23127 (N_23127,N_22227,N_22433);
and U23128 (N_23128,N_21658,N_22586);
xnor U23129 (N_23129,N_22776,N_22038);
nor U23130 (N_23130,N_21702,N_22582);
and U23131 (N_23131,N_21995,N_22487);
nand U23132 (N_23132,N_21886,N_22563);
nor U23133 (N_23133,N_22241,N_22219);
and U23134 (N_23134,N_22072,N_22107);
and U23135 (N_23135,N_21835,N_22462);
nand U23136 (N_23136,N_22363,N_22530);
and U23137 (N_23137,N_22257,N_21968);
nand U23138 (N_23138,N_22607,N_22443);
xnor U23139 (N_23139,N_22544,N_22683);
nand U23140 (N_23140,N_22269,N_22580);
nand U23141 (N_23141,N_22516,N_22236);
xor U23142 (N_23142,N_21923,N_21872);
or U23143 (N_23143,N_22747,N_21742);
nor U23144 (N_23144,N_21688,N_22391);
nor U23145 (N_23145,N_21696,N_21672);
nand U23146 (N_23146,N_22180,N_21822);
or U23147 (N_23147,N_22162,N_22172);
nand U23148 (N_23148,N_21740,N_22203);
nor U23149 (N_23149,N_22315,N_21796);
nand U23150 (N_23150,N_21762,N_22693);
nor U23151 (N_23151,N_22628,N_22409);
nor U23152 (N_23152,N_22527,N_22319);
xor U23153 (N_23153,N_21646,N_21999);
nor U23154 (N_23154,N_22406,N_22632);
xnor U23155 (N_23155,N_22354,N_22245);
nor U23156 (N_23156,N_21620,N_21682);
nand U23157 (N_23157,N_21957,N_22175);
or U23158 (N_23158,N_22006,N_21789);
xor U23159 (N_23159,N_22656,N_22160);
nor U23160 (N_23160,N_22690,N_22720);
and U23161 (N_23161,N_21738,N_22478);
nand U23162 (N_23162,N_22388,N_21900);
nor U23163 (N_23163,N_21773,N_22092);
xor U23164 (N_23164,N_22142,N_21880);
or U23165 (N_23165,N_22128,N_21891);
nor U23166 (N_23166,N_21878,N_21766);
or U23167 (N_23167,N_21939,N_21770);
and U23168 (N_23168,N_21663,N_22047);
and U23169 (N_23169,N_21961,N_22427);
or U23170 (N_23170,N_22212,N_21604);
nand U23171 (N_23171,N_22392,N_22335);
and U23172 (N_23172,N_22692,N_21829);
or U23173 (N_23173,N_22389,N_22051);
nand U23174 (N_23174,N_21775,N_22793);
nand U23175 (N_23175,N_22078,N_22030);
nor U23176 (N_23176,N_22411,N_21802);
nor U23177 (N_23177,N_22185,N_22471);
or U23178 (N_23178,N_21782,N_22216);
and U23179 (N_23179,N_22759,N_22116);
or U23180 (N_23180,N_22341,N_22593);
nor U23181 (N_23181,N_22009,N_22610);
xnor U23182 (N_23182,N_22535,N_22329);
nand U23183 (N_23183,N_22538,N_22763);
xnor U23184 (N_23184,N_21889,N_21642);
xor U23185 (N_23185,N_22620,N_22525);
or U23186 (N_23186,N_22124,N_22450);
nand U23187 (N_23187,N_22279,N_22421);
xor U23188 (N_23188,N_21616,N_22201);
xnor U23189 (N_23189,N_22459,N_22419);
or U23190 (N_23190,N_21879,N_22370);
or U23191 (N_23191,N_22246,N_22627);
nor U23192 (N_23192,N_21744,N_21910);
and U23193 (N_23193,N_21662,N_22635);
or U23194 (N_23194,N_22213,N_21819);
and U23195 (N_23195,N_21681,N_22637);
nand U23196 (N_23196,N_21645,N_22120);
nand U23197 (N_23197,N_22567,N_22615);
and U23198 (N_23198,N_22640,N_21791);
and U23199 (N_23199,N_21793,N_21761);
nor U23200 (N_23200,N_22642,N_22287);
nand U23201 (N_23201,N_21670,N_22486);
nand U23202 (N_23202,N_21976,N_22025);
nand U23203 (N_23203,N_22781,N_22294);
nand U23204 (N_23204,N_22222,N_22775);
or U23205 (N_23205,N_22679,N_21903);
or U23206 (N_23206,N_21617,N_21686);
nand U23207 (N_23207,N_22552,N_22678);
and U23208 (N_23208,N_22102,N_22625);
nand U23209 (N_23209,N_22740,N_22473);
and U23210 (N_23210,N_22085,N_21946);
xnor U23211 (N_23211,N_21843,N_22280);
nor U23212 (N_23212,N_21605,N_22314);
and U23213 (N_23213,N_22706,N_21621);
and U23214 (N_23214,N_22476,N_22501);
nor U23215 (N_23215,N_22378,N_21851);
nor U23216 (N_23216,N_22682,N_22155);
and U23217 (N_23217,N_21890,N_21634);
and U23218 (N_23218,N_22416,N_22797);
nor U23219 (N_23219,N_21728,N_21797);
nor U23220 (N_23220,N_21695,N_22125);
or U23221 (N_23221,N_22215,N_22161);
nor U23222 (N_23222,N_21956,N_22619);
xnor U23223 (N_23223,N_21881,N_21678);
or U23224 (N_23224,N_21721,N_22368);
xnor U23225 (N_23225,N_22278,N_22119);
nand U23226 (N_23226,N_22643,N_21815);
and U23227 (N_23227,N_22230,N_21981);
nand U23228 (N_23228,N_21780,N_21801);
or U23229 (N_23229,N_22668,N_22587);
and U23230 (N_23230,N_22361,N_22447);
and U23231 (N_23231,N_22687,N_22571);
nor U23232 (N_23232,N_21935,N_22352);
nor U23233 (N_23233,N_22708,N_22260);
nand U23234 (N_23234,N_22758,N_22344);
xnor U23235 (N_23235,N_22055,N_22602);
nor U23236 (N_23236,N_22576,N_22353);
nand U23237 (N_23237,N_22613,N_22302);
or U23238 (N_23238,N_22724,N_21931);
or U23239 (N_23239,N_21830,N_22017);
nor U23240 (N_23240,N_21971,N_22788);
or U23241 (N_23241,N_22592,N_21612);
or U23242 (N_23242,N_22183,N_22021);
or U23243 (N_23243,N_22508,N_22158);
or U23244 (N_23244,N_22252,N_22420);
nor U23245 (N_23245,N_22380,N_22012);
and U23246 (N_23246,N_21996,N_21811);
nor U23247 (N_23247,N_22543,N_21689);
and U23248 (N_23248,N_21902,N_21944);
and U23249 (N_23249,N_21997,N_22561);
nor U23250 (N_23250,N_22514,N_22109);
nor U23251 (N_23251,N_21687,N_21883);
or U23252 (N_23252,N_22649,N_22080);
nand U23253 (N_23253,N_21741,N_21839);
and U23254 (N_23254,N_22520,N_22070);
nor U23255 (N_23255,N_22016,N_21697);
and U23256 (N_23256,N_22026,N_21825);
nor U23257 (N_23257,N_21790,N_22583);
or U23258 (N_23258,N_22791,N_22334);
and U23259 (N_23259,N_21867,N_22008);
nor U23260 (N_23260,N_21777,N_22783);
and U23261 (N_23261,N_21969,N_22772);
xor U23262 (N_23262,N_22575,N_21699);
nand U23263 (N_23263,N_21609,N_21870);
nand U23264 (N_23264,N_22536,N_22282);
and U23265 (N_23265,N_22767,N_22426);
and U23266 (N_23266,N_21854,N_21756);
and U23267 (N_23267,N_22553,N_22490);
nor U23268 (N_23268,N_22019,N_22010);
xor U23269 (N_23269,N_22373,N_21848);
nor U23270 (N_23270,N_22705,N_22605);
or U23271 (N_23271,N_22769,N_22456);
and U23272 (N_23272,N_22458,N_21661);
or U23273 (N_23273,N_22440,N_21804);
and U23274 (N_23274,N_22374,N_22712);
xnor U23275 (N_23275,N_22465,N_22089);
and U23276 (N_23276,N_22594,N_22662);
or U23277 (N_23277,N_22565,N_22320);
xnor U23278 (N_23278,N_22132,N_22773);
or U23279 (N_23279,N_22641,N_22357);
and U23280 (N_23280,N_22375,N_21608);
xor U23281 (N_23281,N_22355,N_21705);
xor U23282 (N_23282,N_21611,N_21922);
or U23283 (N_23283,N_22700,N_22432);
or U23284 (N_23284,N_22515,N_22540);
or U23285 (N_23285,N_22348,N_22384);
or U23286 (N_23286,N_22677,N_22321);
nand U23287 (N_23287,N_22394,N_22410);
nor U23288 (N_23288,N_22358,N_21836);
nor U23289 (N_23289,N_22176,N_22449);
and U23290 (N_23290,N_22293,N_21847);
nor U23291 (N_23291,N_22056,N_22194);
or U23292 (N_23292,N_22050,N_21925);
nor U23293 (N_23293,N_22202,N_22736);
xor U23294 (N_23294,N_22481,N_22425);
and U23295 (N_23295,N_22401,N_22665);
nor U23296 (N_23296,N_21894,N_22262);
nor U23297 (N_23297,N_22131,N_21798);
or U23298 (N_23298,N_22022,N_21896);
xor U23299 (N_23299,N_22526,N_22669);
or U23300 (N_23300,N_21643,N_22187);
or U23301 (N_23301,N_21729,N_22207);
and U23302 (N_23302,N_22630,N_22778);
nor U23303 (N_23303,N_21924,N_22455);
or U23304 (N_23304,N_22528,N_21823);
xnor U23305 (N_23305,N_22343,N_22367);
nand U23306 (N_23306,N_22570,N_21755);
nor U23307 (N_23307,N_21933,N_22303);
nand U23308 (N_23308,N_22234,N_22795);
nand U23309 (N_23309,N_21737,N_21735);
xnor U23310 (N_23310,N_22457,N_21692);
nor U23311 (N_23311,N_21768,N_22094);
and U23312 (N_23312,N_22304,N_22753);
xor U23313 (N_23313,N_21653,N_22703);
nor U23314 (N_23314,N_22556,N_21864);
nand U23315 (N_23315,N_21693,N_22751);
xnor U23316 (N_23316,N_22000,N_22591);
nor U23317 (N_23317,N_22043,N_22100);
nand U23318 (N_23318,N_22174,N_21869);
nor U23319 (N_23319,N_22164,N_22614);
and U23320 (N_23320,N_22667,N_22088);
nand U23321 (N_23321,N_22417,N_22494);
and U23322 (N_23322,N_21623,N_22422);
nand U23323 (N_23323,N_22766,N_22281);
nor U23324 (N_23324,N_22052,N_22096);
nor U23325 (N_23325,N_22418,N_22163);
or U23326 (N_23326,N_21805,N_22601);
or U23327 (N_23327,N_21778,N_21745);
or U23328 (N_23328,N_22381,N_21978);
nor U23329 (N_23329,N_22083,N_21603);
xor U23330 (N_23330,N_22248,N_22339);
xnor U23331 (N_23331,N_22290,N_22040);
and U23332 (N_23332,N_21650,N_22324);
nand U23333 (N_23333,N_22251,N_21637);
nand U23334 (N_23334,N_21785,N_22179);
or U23335 (N_23335,N_21602,N_21993);
and U23336 (N_23336,N_21972,N_21676);
and U23337 (N_23337,N_22734,N_22603);
xnor U23338 (N_23338,N_22015,N_22042);
nor U23339 (N_23339,N_22414,N_21633);
xor U23340 (N_23340,N_22390,N_21932);
nor U23341 (N_23341,N_21885,N_22169);
and U23342 (N_23342,N_22111,N_22196);
or U23343 (N_23343,N_22351,N_22542);
or U23344 (N_23344,N_22492,N_21649);
and U23345 (N_23345,N_22461,N_21828);
nor U23346 (N_23346,N_21953,N_21751);
nand U23347 (N_23347,N_21703,N_21988);
and U23348 (N_23348,N_22650,N_21951);
nor U23349 (N_23349,N_21764,N_22121);
and U23350 (N_23350,N_22221,N_21808);
xnor U23351 (N_23351,N_22564,N_22371);
xnor U23352 (N_23352,N_22609,N_21807);
or U23353 (N_23353,N_22622,N_21950);
xnor U23354 (N_23354,N_22584,N_22306);
xnor U23355 (N_23355,N_22633,N_22059);
or U23356 (N_23356,N_22644,N_22044);
and U23357 (N_23357,N_22228,N_21767);
and U23358 (N_23358,N_22671,N_22436);
nand U23359 (N_23359,N_22379,N_21640);
or U23360 (N_23360,N_22296,N_21841);
nor U23361 (N_23361,N_22722,N_21960);
nor U23362 (N_23362,N_22152,N_21792);
nand U23363 (N_23363,N_21994,N_22786);
and U23364 (N_23364,N_22631,N_22397);
and U23365 (N_23365,N_22638,N_21992);
and U23366 (N_23366,N_22101,N_21626);
nand U23367 (N_23367,N_22502,N_22489);
nor U23368 (N_23368,N_22369,N_21868);
nand U23369 (N_23369,N_22403,N_22497);
and U23370 (N_23370,N_22270,N_21673);
nor U23371 (N_23371,N_22220,N_22217);
xor U23372 (N_23372,N_21979,N_21671);
xor U23373 (N_23373,N_21669,N_21821);
xor U23374 (N_23374,N_21966,N_22562);
xnor U23375 (N_23375,N_22557,N_21712);
and U23376 (N_23376,N_21625,N_22534);
xnor U23377 (N_23377,N_21743,N_22299);
nor U23378 (N_23378,N_21722,N_22398);
xor U23379 (N_23379,N_21814,N_22555);
and U23380 (N_23380,N_22159,N_21726);
nor U23381 (N_23381,N_22539,N_22045);
nand U23382 (N_23382,N_22468,N_22496);
xnor U23383 (N_23383,N_22386,N_22399);
nor U23384 (N_23384,N_22331,N_22437);
nand U23385 (N_23385,N_22231,N_22310);
and U23386 (N_23386,N_22336,N_22585);
and U23387 (N_23387,N_21632,N_22144);
nand U23388 (N_23388,N_22084,N_21955);
and U23389 (N_23389,N_22726,N_22711);
or U23390 (N_23390,N_22077,N_22312);
and U23391 (N_23391,N_22110,N_22796);
nor U23392 (N_23392,N_21907,N_22442);
nand U23393 (N_23393,N_21846,N_21838);
nand U23394 (N_23394,N_21911,N_22479);
nand U23395 (N_23395,N_21635,N_21975);
and U23396 (N_23396,N_22053,N_22308);
and U23397 (N_23397,N_21936,N_21674);
nor U23398 (N_23398,N_21786,N_22188);
or U23399 (N_23399,N_22130,N_21651);
nand U23400 (N_23400,N_22120,N_22236);
and U23401 (N_23401,N_22723,N_22742);
nand U23402 (N_23402,N_21816,N_22439);
xor U23403 (N_23403,N_22491,N_22121);
xor U23404 (N_23404,N_21869,N_22521);
xnor U23405 (N_23405,N_21953,N_22299);
or U23406 (N_23406,N_22137,N_22482);
or U23407 (N_23407,N_21872,N_22352);
xor U23408 (N_23408,N_21976,N_22440);
nand U23409 (N_23409,N_22692,N_22605);
and U23410 (N_23410,N_21744,N_22565);
and U23411 (N_23411,N_21741,N_22221);
nor U23412 (N_23412,N_22181,N_22793);
xor U23413 (N_23413,N_22751,N_21787);
or U23414 (N_23414,N_22179,N_22227);
or U23415 (N_23415,N_22709,N_21772);
nor U23416 (N_23416,N_21812,N_21813);
or U23417 (N_23417,N_22460,N_22117);
or U23418 (N_23418,N_22101,N_22135);
xnor U23419 (N_23419,N_21692,N_21936);
or U23420 (N_23420,N_22158,N_22749);
or U23421 (N_23421,N_22035,N_21744);
nand U23422 (N_23422,N_22123,N_22116);
nand U23423 (N_23423,N_22449,N_22706);
nor U23424 (N_23424,N_22773,N_22370);
or U23425 (N_23425,N_21828,N_21836);
or U23426 (N_23426,N_21765,N_22239);
nor U23427 (N_23427,N_21952,N_21675);
or U23428 (N_23428,N_22237,N_22701);
xnor U23429 (N_23429,N_22242,N_22622);
nor U23430 (N_23430,N_22126,N_22766);
or U23431 (N_23431,N_22006,N_22727);
or U23432 (N_23432,N_22231,N_21718);
nand U23433 (N_23433,N_22661,N_21845);
xor U23434 (N_23434,N_22727,N_22180);
or U23435 (N_23435,N_22340,N_21615);
xor U23436 (N_23436,N_22058,N_22301);
and U23437 (N_23437,N_22793,N_22534);
nor U23438 (N_23438,N_22576,N_22021);
nand U23439 (N_23439,N_21605,N_21791);
and U23440 (N_23440,N_21860,N_22467);
nor U23441 (N_23441,N_22784,N_21867);
nor U23442 (N_23442,N_22012,N_21814);
or U23443 (N_23443,N_22344,N_22112);
nor U23444 (N_23444,N_22298,N_22290);
or U23445 (N_23445,N_22491,N_21893);
and U23446 (N_23446,N_22033,N_21787);
xnor U23447 (N_23447,N_22366,N_22681);
xnor U23448 (N_23448,N_22738,N_21800);
or U23449 (N_23449,N_22138,N_22126);
or U23450 (N_23450,N_21981,N_22771);
and U23451 (N_23451,N_22408,N_21680);
nor U23452 (N_23452,N_22579,N_22115);
or U23453 (N_23453,N_22595,N_21757);
nor U23454 (N_23454,N_22796,N_21973);
nor U23455 (N_23455,N_22771,N_21877);
xnor U23456 (N_23456,N_21782,N_22217);
xor U23457 (N_23457,N_21973,N_22722);
xnor U23458 (N_23458,N_21820,N_22422);
nand U23459 (N_23459,N_21978,N_22794);
and U23460 (N_23460,N_22377,N_21946);
nand U23461 (N_23461,N_22594,N_21857);
and U23462 (N_23462,N_21694,N_22259);
and U23463 (N_23463,N_21986,N_22712);
or U23464 (N_23464,N_22364,N_22083);
xnor U23465 (N_23465,N_22703,N_22498);
nand U23466 (N_23466,N_21677,N_22098);
xnor U23467 (N_23467,N_21874,N_21987);
nor U23468 (N_23468,N_22181,N_21794);
nand U23469 (N_23469,N_22413,N_21611);
and U23470 (N_23470,N_22173,N_22188);
and U23471 (N_23471,N_21786,N_22738);
nand U23472 (N_23472,N_21661,N_22656);
nand U23473 (N_23473,N_22296,N_21877);
and U23474 (N_23474,N_21668,N_22525);
and U23475 (N_23475,N_22720,N_21629);
xor U23476 (N_23476,N_22367,N_22019);
xnor U23477 (N_23477,N_22497,N_21683);
nand U23478 (N_23478,N_21830,N_22194);
nor U23479 (N_23479,N_22177,N_22737);
nor U23480 (N_23480,N_21676,N_22626);
or U23481 (N_23481,N_21691,N_22271);
or U23482 (N_23482,N_22781,N_22024);
and U23483 (N_23483,N_22441,N_22524);
nand U23484 (N_23484,N_22694,N_22179);
or U23485 (N_23485,N_22592,N_22479);
and U23486 (N_23486,N_21973,N_22744);
nand U23487 (N_23487,N_21799,N_22608);
nand U23488 (N_23488,N_22558,N_22337);
nor U23489 (N_23489,N_22361,N_22555);
xor U23490 (N_23490,N_22356,N_21647);
nand U23491 (N_23491,N_21873,N_22385);
nand U23492 (N_23492,N_22300,N_22240);
xor U23493 (N_23493,N_22677,N_21849);
nor U23494 (N_23494,N_21830,N_22032);
nand U23495 (N_23495,N_22323,N_21969);
and U23496 (N_23496,N_22640,N_22616);
nor U23497 (N_23497,N_21789,N_22088);
nand U23498 (N_23498,N_22002,N_21763);
nand U23499 (N_23499,N_22164,N_22194);
nand U23500 (N_23500,N_22589,N_22269);
xor U23501 (N_23501,N_22659,N_21910);
or U23502 (N_23502,N_22573,N_22282);
nor U23503 (N_23503,N_22579,N_22533);
or U23504 (N_23504,N_21936,N_22734);
nand U23505 (N_23505,N_21779,N_21613);
or U23506 (N_23506,N_22475,N_22186);
or U23507 (N_23507,N_21954,N_22015);
nand U23508 (N_23508,N_21975,N_22224);
xor U23509 (N_23509,N_22183,N_22712);
nand U23510 (N_23510,N_22692,N_22296);
and U23511 (N_23511,N_22593,N_22722);
xor U23512 (N_23512,N_21980,N_22058);
xor U23513 (N_23513,N_22380,N_21651);
xor U23514 (N_23514,N_22089,N_21816);
nor U23515 (N_23515,N_21630,N_22080);
xor U23516 (N_23516,N_22700,N_21970);
nand U23517 (N_23517,N_22200,N_22664);
and U23518 (N_23518,N_21725,N_21880);
and U23519 (N_23519,N_21991,N_22556);
nor U23520 (N_23520,N_22243,N_21658);
or U23521 (N_23521,N_21757,N_21655);
nand U23522 (N_23522,N_22729,N_22176);
and U23523 (N_23523,N_21693,N_22184);
nand U23524 (N_23524,N_21647,N_21640);
and U23525 (N_23525,N_22748,N_21761);
and U23526 (N_23526,N_22594,N_22611);
and U23527 (N_23527,N_22321,N_22443);
nor U23528 (N_23528,N_22786,N_21749);
xor U23529 (N_23529,N_22623,N_22110);
nor U23530 (N_23530,N_21906,N_21616);
nand U23531 (N_23531,N_21627,N_22679);
or U23532 (N_23532,N_22382,N_21950);
and U23533 (N_23533,N_22614,N_22371);
or U23534 (N_23534,N_22272,N_22486);
xor U23535 (N_23535,N_22758,N_21912);
and U23536 (N_23536,N_22625,N_22128);
nand U23537 (N_23537,N_22634,N_22465);
nand U23538 (N_23538,N_22033,N_21973);
xor U23539 (N_23539,N_21957,N_22629);
nor U23540 (N_23540,N_22417,N_22466);
nand U23541 (N_23541,N_21672,N_22038);
nand U23542 (N_23542,N_21991,N_22751);
and U23543 (N_23543,N_22390,N_22330);
nor U23544 (N_23544,N_21820,N_22063);
xor U23545 (N_23545,N_22314,N_22012);
nand U23546 (N_23546,N_21875,N_22136);
or U23547 (N_23547,N_21943,N_22677);
and U23548 (N_23548,N_22338,N_21815);
or U23549 (N_23549,N_22765,N_21982);
or U23550 (N_23550,N_22327,N_22584);
nor U23551 (N_23551,N_21955,N_22772);
or U23552 (N_23552,N_22557,N_22442);
or U23553 (N_23553,N_22462,N_22024);
nand U23554 (N_23554,N_21854,N_22693);
xor U23555 (N_23555,N_22610,N_22437);
nand U23556 (N_23556,N_22792,N_22520);
or U23557 (N_23557,N_21637,N_21609);
nand U23558 (N_23558,N_21664,N_22696);
or U23559 (N_23559,N_21630,N_22139);
nand U23560 (N_23560,N_22256,N_21883);
and U23561 (N_23561,N_22754,N_22140);
nor U23562 (N_23562,N_22297,N_22240);
or U23563 (N_23563,N_22783,N_22107);
or U23564 (N_23564,N_22375,N_22612);
nand U23565 (N_23565,N_21877,N_21683);
xnor U23566 (N_23566,N_22102,N_21734);
or U23567 (N_23567,N_22362,N_21668);
nand U23568 (N_23568,N_21685,N_22292);
or U23569 (N_23569,N_22467,N_22276);
or U23570 (N_23570,N_22573,N_22499);
and U23571 (N_23571,N_21969,N_21915);
nor U23572 (N_23572,N_22341,N_21768);
nand U23573 (N_23573,N_22741,N_21832);
nor U23574 (N_23574,N_22769,N_22239);
nor U23575 (N_23575,N_22316,N_22486);
xor U23576 (N_23576,N_22666,N_22167);
or U23577 (N_23577,N_21914,N_22023);
xor U23578 (N_23578,N_21763,N_21805);
nor U23579 (N_23579,N_22008,N_22693);
nor U23580 (N_23580,N_22547,N_22127);
xor U23581 (N_23581,N_21613,N_22076);
and U23582 (N_23582,N_22306,N_22265);
or U23583 (N_23583,N_22594,N_22370);
and U23584 (N_23584,N_22485,N_21935);
and U23585 (N_23585,N_21981,N_22453);
xnor U23586 (N_23586,N_21883,N_22237);
nor U23587 (N_23587,N_22353,N_21854);
xor U23588 (N_23588,N_21859,N_22526);
nand U23589 (N_23589,N_22312,N_21600);
and U23590 (N_23590,N_22604,N_22488);
or U23591 (N_23591,N_22755,N_22217);
nor U23592 (N_23592,N_21872,N_21645);
xor U23593 (N_23593,N_22479,N_22648);
xnor U23594 (N_23594,N_21761,N_21664);
and U23595 (N_23595,N_21793,N_22446);
nand U23596 (N_23596,N_21727,N_21957);
and U23597 (N_23597,N_22453,N_22287);
nand U23598 (N_23598,N_21954,N_22282);
xnor U23599 (N_23599,N_22675,N_21600);
nand U23600 (N_23600,N_21718,N_21840);
or U23601 (N_23601,N_22523,N_22234);
nand U23602 (N_23602,N_22399,N_21787);
nor U23603 (N_23603,N_21891,N_21790);
nor U23604 (N_23604,N_22218,N_21759);
nand U23605 (N_23605,N_22384,N_22534);
or U23606 (N_23606,N_21876,N_22056);
or U23607 (N_23607,N_21789,N_22339);
xnor U23608 (N_23608,N_21737,N_22676);
nor U23609 (N_23609,N_22035,N_21899);
nand U23610 (N_23610,N_21758,N_22785);
and U23611 (N_23611,N_22635,N_21605);
nor U23612 (N_23612,N_22262,N_22762);
and U23613 (N_23613,N_21736,N_22296);
nor U23614 (N_23614,N_22489,N_22143);
or U23615 (N_23615,N_21838,N_21623);
and U23616 (N_23616,N_21938,N_22209);
or U23617 (N_23617,N_22169,N_22456);
xnor U23618 (N_23618,N_21606,N_22721);
xor U23619 (N_23619,N_22098,N_21771);
and U23620 (N_23620,N_21714,N_21923);
or U23621 (N_23621,N_21970,N_22465);
nand U23622 (N_23622,N_22011,N_22265);
or U23623 (N_23623,N_22191,N_22406);
nor U23624 (N_23624,N_22414,N_21859);
nor U23625 (N_23625,N_21839,N_22346);
nand U23626 (N_23626,N_21950,N_22291);
and U23627 (N_23627,N_22727,N_22053);
nand U23628 (N_23628,N_22027,N_21683);
nand U23629 (N_23629,N_21953,N_21817);
xnor U23630 (N_23630,N_22293,N_21862);
or U23631 (N_23631,N_22206,N_22462);
nor U23632 (N_23632,N_22298,N_22388);
nand U23633 (N_23633,N_22266,N_21968);
nand U23634 (N_23634,N_22451,N_21709);
and U23635 (N_23635,N_22683,N_21681);
and U23636 (N_23636,N_22129,N_21898);
nor U23637 (N_23637,N_21673,N_21998);
nor U23638 (N_23638,N_22061,N_21876);
or U23639 (N_23639,N_22785,N_22050);
nand U23640 (N_23640,N_21631,N_22296);
or U23641 (N_23641,N_21645,N_21857);
xnor U23642 (N_23642,N_22085,N_22408);
nor U23643 (N_23643,N_22341,N_21637);
nor U23644 (N_23644,N_22759,N_21739);
xor U23645 (N_23645,N_22645,N_22259);
nand U23646 (N_23646,N_21931,N_22383);
nor U23647 (N_23647,N_21947,N_22646);
or U23648 (N_23648,N_21933,N_22579);
nand U23649 (N_23649,N_22790,N_22252);
and U23650 (N_23650,N_22324,N_22521);
or U23651 (N_23651,N_22388,N_22030);
or U23652 (N_23652,N_21690,N_22311);
nor U23653 (N_23653,N_22331,N_21636);
or U23654 (N_23654,N_22723,N_21754);
xnor U23655 (N_23655,N_22753,N_22489);
nor U23656 (N_23656,N_22126,N_21987);
xor U23657 (N_23657,N_22204,N_22702);
xor U23658 (N_23658,N_22732,N_22351);
nand U23659 (N_23659,N_22175,N_22682);
nand U23660 (N_23660,N_22325,N_22401);
xnor U23661 (N_23661,N_22438,N_22388);
and U23662 (N_23662,N_22604,N_22491);
nand U23663 (N_23663,N_21996,N_22386);
nand U23664 (N_23664,N_21999,N_22240);
nand U23665 (N_23665,N_21786,N_22171);
or U23666 (N_23666,N_22188,N_22285);
nand U23667 (N_23667,N_22487,N_22774);
nor U23668 (N_23668,N_21784,N_22639);
nand U23669 (N_23669,N_22221,N_22467);
or U23670 (N_23670,N_21618,N_22259);
and U23671 (N_23671,N_22184,N_22249);
or U23672 (N_23672,N_22238,N_21894);
xor U23673 (N_23673,N_21677,N_22731);
nand U23674 (N_23674,N_22455,N_22378);
nor U23675 (N_23675,N_22757,N_22027);
and U23676 (N_23676,N_21869,N_22432);
and U23677 (N_23677,N_22492,N_22293);
or U23678 (N_23678,N_22455,N_22213);
or U23679 (N_23679,N_22347,N_22675);
nand U23680 (N_23680,N_21911,N_22184);
nor U23681 (N_23681,N_21895,N_22677);
and U23682 (N_23682,N_21892,N_21966);
and U23683 (N_23683,N_21648,N_21851);
or U23684 (N_23684,N_21997,N_22632);
nor U23685 (N_23685,N_22336,N_22314);
or U23686 (N_23686,N_22742,N_21656);
nand U23687 (N_23687,N_22670,N_21698);
xor U23688 (N_23688,N_22624,N_21850);
xnor U23689 (N_23689,N_22518,N_22798);
xnor U23690 (N_23690,N_22154,N_22707);
nand U23691 (N_23691,N_21990,N_22415);
nor U23692 (N_23692,N_22377,N_22396);
nand U23693 (N_23693,N_21951,N_22588);
or U23694 (N_23694,N_22538,N_21985);
nand U23695 (N_23695,N_22196,N_22297);
or U23696 (N_23696,N_21639,N_22751);
nor U23697 (N_23697,N_22374,N_22263);
and U23698 (N_23698,N_22240,N_22418);
nor U23699 (N_23699,N_22377,N_22608);
or U23700 (N_23700,N_22182,N_22218);
or U23701 (N_23701,N_21772,N_22573);
nand U23702 (N_23702,N_22110,N_22626);
nor U23703 (N_23703,N_21606,N_21943);
and U23704 (N_23704,N_22606,N_22663);
xor U23705 (N_23705,N_22507,N_21931);
nor U23706 (N_23706,N_22574,N_22457);
nand U23707 (N_23707,N_22106,N_22186);
nor U23708 (N_23708,N_22005,N_22155);
nor U23709 (N_23709,N_21970,N_22562);
nand U23710 (N_23710,N_21860,N_22339);
nand U23711 (N_23711,N_22507,N_22171);
xor U23712 (N_23712,N_22064,N_22315);
and U23713 (N_23713,N_22221,N_22063);
and U23714 (N_23714,N_22283,N_22453);
nand U23715 (N_23715,N_22799,N_22597);
nor U23716 (N_23716,N_22556,N_21833);
and U23717 (N_23717,N_22327,N_21934);
xnor U23718 (N_23718,N_22566,N_22613);
nor U23719 (N_23719,N_22510,N_21752);
xor U23720 (N_23720,N_22759,N_22271);
nor U23721 (N_23721,N_22328,N_22313);
and U23722 (N_23722,N_22456,N_21772);
nor U23723 (N_23723,N_22702,N_22403);
and U23724 (N_23724,N_22690,N_21938);
xor U23725 (N_23725,N_22519,N_21868);
xor U23726 (N_23726,N_21827,N_22734);
and U23727 (N_23727,N_22679,N_21671);
or U23728 (N_23728,N_22226,N_22697);
or U23729 (N_23729,N_21813,N_22599);
and U23730 (N_23730,N_21721,N_22606);
and U23731 (N_23731,N_22080,N_21820);
xnor U23732 (N_23732,N_21946,N_22120);
nand U23733 (N_23733,N_21959,N_22556);
and U23734 (N_23734,N_22231,N_21723);
nor U23735 (N_23735,N_21755,N_22113);
xnor U23736 (N_23736,N_21626,N_22185);
nor U23737 (N_23737,N_22195,N_21842);
nor U23738 (N_23738,N_21626,N_21931);
or U23739 (N_23739,N_22038,N_22003);
and U23740 (N_23740,N_22637,N_22405);
or U23741 (N_23741,N_21951,N_21791);
xor U23742 (N_23742,N_22770,N_21671);
nand U23743 (N_23743,N_22081,N_21999);
xnor U23744 (N_23744,N_22666,N_22761);
and U23745 (N_23745,N_22022,N_21912);
xnor U23746 (N_23746,N_22584,N_22393);
or U23747 (N_23747,N_21663,N_22020);
or U23748 (N_23748,N_21614,N_21728);
and U23749 (N_23749,N_21639,N_21714);
nor U23750 (N_23750,N_21805,N_21603);
or U23751 (N_23751,N_22517,N_22158);
and U23752 (N_23752,N_21917,N_22199);
nand U23753 (N_23753,N_21698,N_22599);
nor U23754 (N_23754,N_22176,N_22787);
and U23755 (N_23755,N_22563,N_21675);
nand U23756 (N_23756,N_22196,N_21869);
xnor U23757 (N_23757,N_22199,N_22016);
xnor U23758 (N_23758,N_21753,N_21754);
nand U23759 (N_23759,N_22215,N_22341);
and U23760 (N_23760,N_21919,N_22169);
nand U23761 (N_23761,N_21712,N_21817);
and U23762 (N_23762,N_21995,N_22500);
or U23763 (N_23763,N_22291,N_22534);
nand U23764 (N_23764,N_21714,N_22036);
xnor U23765 (N_23765,N_21945,N_21837);
nand U23766 (N_23766,N_22130,N_22714);
xnor U23767 (N_23767,N_21967,N_22500);
or U23768 (N_23768,N_22482,N_21781);
nand U23769 (N_23769,N_22515,N_21999);
or U23770 (N_23770,N_21667,N_21755);
xor U23771 (N_23771,N_22010,N_21852);
nor U23772 (N_23772,N_22648,N_21716);
xor U23773 (N_23773,N_22448,N_22096);
nand U23774 (N_23774,N_22590,N_21773);
xnor U23775 (N_23775,N_22101,N_22729);
or U23776 (N_23776,N_22644,N_21654);
and U23777 (N_23777,N_22182,N_21946);
nor U23778 (N_23778,N_21678,N_22789);
xnor U23779 (N_23779,N_22768,N_22756);
and U23780 (N_23780,N_22013,N_21721);
or U23781 (N_23781,N_22114,N_21977);
nor U23782 (N_23782,N_22301,N_22712);
nor U23783 (N_23783,N_22297,N_22049);
nor U23784 (N_23784,N_22091,N_21908);
nand U23785 (N_23785,N_22001,N_22550);
nor U23786 (N_23786,N_22015,N_22280);
or U23787 (N_23787,N_21674,N_22766);
nor U23788 (N_23788,N_21703,N_22514);
xnor U23789 (N_23789,N_22796,N_21949);
xor U23790 (N_23790,N_22130,N_21871);
xnor U23791 (N_23791,N_22067,N_22215);
nor U23792 (N_23792,N_22040,N_21878);
nor U23793 (N_23793,N_21960,N_22328);
nand U23794 (N_23794,N_21923,N_22415);
nand U23795 (N_23795,N_22124,N_22070);
nor U23796 (N_23796,N_22409,N_22492);
or U23797 (N_23797,N_22503,N_22734);
and U23798 (N_23798,N_21636,N_21859);
nor U23799 (N_23799,N_22372,N_22152);
or U23800 (N_23800,N_22596,N_21793);
nor U23801 (N_23801,N_22519,N_22172);
nor U23802 (N_23802,N_22080,N_21700);
nand U23803 (N_23803,N_22777,N_21945);
nor U23804 (N_23804,N_22380,N_22325);
or U23805 (N_23805,N_22650,N_22015);
and U23806 (N_23806,N_21813,N_22211);
or U23807 (N_23807,N_22737,N_21622);
nor U23808 (N_23808,N_22120,N_22615);
xnor U23809 (N_23809,N_22740,N_22386);
nor U23810 (N_23810,N_22662,N_22544);
xnor U23811 (N_23811,N_22424,N_22506);
nand U23812 (N_23812,N_21633,N_22687);
or U23813 (N_23813,N_22362,N_21880);
nor U23814 (N_23814,N_22574,N_21713);
nand U23815 (N_23815,N_22639,N_22439);
nand U23816 (N_23816,N_22243,N_21652);
nor U23817 (N_23817,N_22433,N_22799);
xnor U23818 (N_23818,N_21820,N_22150);
and U23819 (N_23819,N_21801,N_22699);
nand U23820 (N_23820,N_22601,N_22502);
xnor U23821 (N_23821,N_22529,N_22388);
or U23822 (N_23822,N_21966,N_22409);
xnor U23823 (N_23823,N_22360,N_21626);
nor U23824 (N_23824,N_21989,N_21869);
xnor U23825 (N_23825,N_22200,N_21831);
or U23826 (N_23826,N_22694,N_21914);
or U23827 (N_23827,N_22155,N_22520);
or U23828 (N_23828,N_21668,N_22298);
or U23829 (N_23829,N_22786,N_22332);
xnor U23830 (N_23830,N_21832,N_22160);
xnor U23831 (N_23831,N_22590,N_22614);
xor U23832 (N_23832,N_22649,N_22003);
nor U23833 (N_23833,N_22688,N_22779);
nor U23834 (N_23834,N_22524,N_22269);
nand U23835 (N_23835,N_22528,N_22718);
nand U23836 (N_23836,N_22549,N_22052);
and U23837 (N_23837,N_22587,N_22767);
xnor U23838 (N_23838,N_22561,N_22543);
xor U23839 (N_23839,N_21605,N_22179);
xnor U23840 (N_23840,N_22032,N_21871);
nor U23841 (N_23841,N_22371,N_21733);
xor U23842 (N_23842,N_22333,N_22007);
nand U23843 (N_23843,N_22560,N_21615);
and U23844 (N_23844,N_21792,N_21909);
and U23845 (N_23845,N_21947,N_21635);
xnor U23846 (N_23846,N_21788,N_21620);
or U23847 (N_23847,N_22537,N_22115);
or U23848 (N_23848,N_21816,N_21717);
xor U23849 (N_23849,N_22230,N_22399);
xor U23850 (N_23850,N_21859,N_22648);
and U23851 (N_23851,N_22478,N_22398);
and U23852 (N_23852,N_21877,N_22707);
nand U23853 (N_23853,N_22404,N_22661);
or U23854 (N_23854,N_21732,N_22541);
and U23855 (N_23855,N_21677,N_21691);
and U23856 (N_23856,N_22743,N_22135);
xnor U23857 (N_23857,N_21807,N_21917);
nor U23858 (N_23858,N_22478,N_21943);
nand U23859 (N_23859,N_22790,N_22266);
nand U23860 (N_23860,N_22439,N_21621);
nand U23861 (N_23861,N_22557,N_21665);
nor U23862 (N_23862,N_21754,N_22107);
nand U23863 (N_23863,N_22531,N_22435);
and U23864 (N_23864,N_22000,N_22625);
or U23865 (N_23865,N_22061,N_22417);
or U23866 (N_23866,N_21960,N_22600);
nor U23867 (N_23867,N_22296,N_22471);
or U23868 (N_23868,N_21902,N_21971);
or U23869 (N_23869,N_22094,N_21614);
nor U23870 (N_23870,N_21666,N_21680);
nand U23871 (N_23871,N_21865,N_21831);
or U23872 (N_23872,N_21861,N_22056);
and U23873 (N_23873,N_22318,N_22774);
nor U23874 (N_23874,N_22632,N_21669);
nor U23875 (N_23875,N_22728,N_22149);
nor U23876 (N_23876,N_21680,N_21645);
nor U23877 (N_23877,N_22633,N_21614);
nand U23878 (N_23878,N_22070,N_22148);
nor U23879 (N_23879,N_21760,N_21737);
and U23880 (N_23880,N_21634,N_22019);
xnor U23881 (N_23881,N_22530,N_22477);
and U23882 (N_23882,N_22242,N_21834);
or U23883 (N_23883,N_22316,N_22290);
nor U23884 (N_23884,N_22107,N_21864);
xor U23885 (N_23885,N_22197,N_21820);
nor U23886 (N_23886,N_22736,N_22501);
and U23887 (N_23887,N_22090,N_22435);
nand U23888 (N_23888,N_21923,N_21645);
nor U23889 (N_23889,N_22768,N_21889);
nor U23890 (N_23890,N_22485,N_22141);
xor U23891 (N_23891,N_22371,N_22711);
and U23892 (N_23892,N_22655,N_22765);
or U23893 (N_23893,N_22136,N_21626);
and U23894 (N_23894,N_22797,N_22026);
xnor U23895 (N_23895,N_22119,N_22630);
or U23896 (N_23896,N_21968,N_22228);
nor U23897 (N_23897,N_21691,N_22171);
xor U23898 (N_23898,N_22238,N_22329);
nor U23899 (N_23899,N_21651,N_22379);
nand U23900 (N_23900,N_21980,N_22015);
and U23901 (N_23901,N_22342,N_21840);
or U23902 (N_23902,N_22255,N_21633);
or U23903 (N_23903,N_21736,N_22578);
or U23904 (N_23904,N_21849,N_22181);
or U23905 (N_23905,N_21854,N_21822);
xor U23906 (N_23906,N_22646,N_22735);
xnor U23907 (N_23907,N_22746,N_22252);
or U23908 (N_23908,N_22087,N_22770);
and U23909 (N_23909,N_22307,N_22419);
xnor U23910 (N_23910,N_22397,N_21739);
nor U23911 (N_23911,N_21979,N_21770);
or U23912 (N_23912,N_22190,N_22096);
and U23913 (N_23913,N_21930,N_22127);
xnor U23914 (N_23914,N_22128,N_22705);
nand U23915 (N_23915,N_22030,N_22205);
nand U23916 (N_23916,N_22512,N_22692);
nor U23917 (N_23917,N_22149,N_21935);
nor U23918 (N_23918,N_22341,N_21702);
nor U23919 (N_23919,N_21846,N_22531);
xnor U23920 (N_23920,N_22670,N_21717);
xor U23921 (N_23921,N_22603,N_21610);
nor U23922 (N_23922,N_21631,N_21746);
and U23923 (N_23923,N_21718,N_21731);
nand U23924 (N_23924,N_21841,N_22263);
and U23925 (N_23925,N_22298,N_21794);
or U23926 (N_23926,N_21917,N_22541);
xnor U23927 (N_23927,N_22068,N_22163);
xnor U23928 (N_23928,N_22537,N_21726);
nand U23929 (N_23929,N_22617,N_21981);
xnor U23930 (N_23930,N_22394,N_22191);
and U23931 (N_23931,N_21695,N_22277);
nor U23932 (N_23932,N_21804,N_21788);
or U23933 (N_23933,N_22640,N_21808);
xnor U23934 (N_23934,N_22110,N_22551);
or U23935 (N_23935,N_22067,N_21658);
xnor U23936 (N_23936,N_22182,N_21690);
nand U23937 (N_23937,N_22187,N_22127);
xnor U23938 (N_23938,N_21879,N_22097);
nand U23939 (N_23939,N_22701,N_22646);
or U23940 (N_23940,N_22276,N_22583);
xnor U23941 (N_23941,N_22064,N_21709);
and U23942 (N_23942,N_21853,N_21690);
xor U23943 (N_23943,N_21783,N_22625);
or U23944 (N_23944,N_22672,N_21754);
xor U23945 (N_23945,N_22579,N_22628);
nor U23946 (N_23946,N_21997,N_22670);
or U23947 (N_23947,N_22475,N_22187);
and U23948 (N_23948,N_21872,N_22331);
nand U23949 (N_23949,N_21683,N_21849);
nand U23950 (N_23950,N_21976,N_21910);
or U23951 (N_23951,N_22770,N_22461);
nor U23952 (N_23952,N_22197,N_21872);
nor U23953 (N_23953,N_22633,N_21757);
nor U23954 (N_23954,N_21737,N_22451);
or U23955 (N_23955,N_22519,N_22292);
xnor U23956 (N_23956,N_22558,N_22371);
or U23957 (N_23957,N_22522,N_22422);
or U23958 (N_23958,N_22662,N_22677);
xor U23959 (N_23959,N_22742,N_22777);
and U23960 (N_23960,N_22657,N_22512);
nor U23961 (N_23961,N_21768,N_21654);
nor U23962 (N_23962,N_22276,N_21974);
and U23963 (N_23963,N_22077,N_22675);
nand U23964 (N_23964,N_21609,N_22081);
or U23965 (N_23965,N_22003,N_22675);
xor U23966 (N_23966,N_21925,N_22255);
nand U23967 (N_23967,N_21664,N_22022);
and U23968 (N_23968,N_21723,N_22253);
or U23969 (N_23969,N_22444,N_22188);
or U23970 (N_23970,N_22313,N_21794);
xnor U23971 (N_23971,N_21894,N_22557);
nand U23972 (N_23972,N_22554,N_21725);
xnor U23973 (N_23973,N_21951,N_21684);
nor U23974 (N_23974,N_22389,N_21772);
and U23975 (N_23975,N_22788,N_22621);
and U23976 (N_23976,N_21739,N_21666);
nand U23977 (N_23977,N_21634,N_22737);
nand U23978 (N_23978,N_22424,N_21698);
or U23979 (N_23979,N_22664,N_22006);
nor U23980 (N_23980,N_22562,N_22060);
nand U23981 (N_23981,N_22335,N_22035);
nand U23982 (N_23982,N_21875,N_22042);
or U23983 (N_23983,N_22350,N_22728);
nand U23984 (N_23984,N_22398,N_21610);
nor U23985 (N_23985,N_22028,N_21750);
or U23986 (N_23986,N_22322,N_21889);
xnor U23987 (N_23987,N_21960,N_22105);
nand U23988 (N_23988,N_21601,N_22650);
or U23989 (N_23989,N_21980,N_22626);
or U23990 (N_23990,N_21665,N_21861);
nor U23991 (N_23991,N_21997,N_21748);
or U23992 (N_23992,N_22343,N_22539);
xor U23993 (N_23993,N_22706,N_22769);
and U23994 (N_23994,N_22581,N_21837);
nor U23995 (N_23995,N_22023,N_22706);
nand U23996 (N_23996,N_22105,N_21668);
xor U23997 (N_23997,N_21679,N_22609);
nor U23998 (N_23998,N_22673,N_22646);
nor U23999 (N_23999,N_22456,N_21802);
and U24000 (N_24000,N_23909,N_23806);
and U24001 (N_24001,N_23392,N_23800);
nor U24002 (N_24002,N_23462,N_23687);
or U24003 (N_24003,N_23463,N_23683);
nand U24004 (N_24004,N_23423,N_23070);
or U24005 (N_24005,N_23726,N_23970);
and U24006 (N_24006,N_23551,N_23669);
nand U24007 (N_24007,N_23252,N_22821);
nand U24008 (N_24008,N_23224,N_23881);
xor U24009 (N_24009,N_22894,N_23426);
and U24010 (N_24010,N_23651,N_23022);
nand U24011 (N_24011,N_23573,N_23418);
and U24012 (N_24012,N_23405,N_23384);
and U24013 (N_24013,N_23615,N_23364);
xor U24014 (N_24014,N_22925,N_23213);
nor U24015 (N_24015,N_23483,N_23212);
or U24016 (N_24016,N_23717,N_23904);
and U24017 (N_24017,N_23265,N_23744);
nor U24018 (N_24018,N_22830,N_23964);
and U24019 (N_24019,N_23903,N_23398);
or U24020 (N_24020,N_23182,N_23766);
xor U24021 (N_24021,N_23201,N_23568);
nor U24022 (N_24022,N_23007,N_23288);
nand U24023 (N_24023,N_23145,N_23066);
nor U24024 (N_24024,N_23893,N_23016);
or U24025 (N_24025,N_23880,N_23550);
xnor U24026 (N_24026,N_23902,N_23057);
nand U24027 (N_24027,N_23994,N_23046);
nand U24028 (N_24028,N_23808,N_23660);
nand U24029 (N_24029,N_23014,N_23792);
and U24030 (N_24030,N_23432,N_23622);
or U24031 (N_24031,N_23699,N_23887);
nor U24032 (N_24032,N_23328,N_23067);
xnor U24033 (N_24033,N_23225,N_23873);
and U24034 (N_24034,N_23498,N_23454);
nor U24035 (N_24035,N_23018,N_23960);
and U24036 (N_24036,N_23223,N_22924);
or U24037 (N_24037,N_23092,N_23291);
nor U24038 (N_24038,N_22928,N_23209);
or U24039 (N_24039,N_23511,N_22882);
or U24040 (N_24040,N_22845,N_23048);
xnor U24041 (N_24041,N_23495,N_23528);
nor U24042 (N_24042,N_23434,N_23440);
and U24043 (N_24043,N_22805,N_23202);
and U24044 (N_24044,N_22919,N_22858);
nor U24045 (N_24045,N_23343,N_23389);
and U24046 (N_24046,N_23447,N_23085);
nand U24047 (N_24047,N_23408,N_23886);
and U24048 (N_24048,N_22914,N_23136);
nand U24049 (N_24049,N_23997,N_23376);
nor U24050 (N_24050,N_23159,N_23080);
xnor U24051 (N_24051,N_23190,N_23117);
or U24052 (N_24052,N_23888,N_23137);
xor U24053 (N_24053,N_23712,N_23298);
or U24054 (N_24054,N_23630,N_23931);
nor U24055 (N_24055,N_23126,N_23461);
and U24056 (N_24056,N_23756,N_23788);
xor U24057 (N_24057,N_23820,N_23193);
and U24058 (N_24058,N_23277,N_23656);
or U24059 (N_24059,N_23335,N_23465);
nor U24060 (N_24060,N_23588,N_22897);
and U24061 (N_24061,N_23394,N_23877);
and U24062 (N_24062,N_23305,N_23684);
or U24063 (N_24063,N_23499,N_23316);
nor U24064 (N_24064,N_22840,N_23179);
nand U24065 (N_24065,N_23946,N_22950);
nor U24066 (N_24066,N_23555,N_23494);
nand U24067 (N_24067,N_23192,N_23149);
nor U24068 (N_24068,N_23696,N_23093);
or U24069 (N_24069,N_23090,N_23890);
nor U24070 (N_24070,N_23488,N_23464);
nor U24071 (N_24071,N_23337,N_23832);
nor U24072 (N_24072,N_23530,N_22901);
or U24073 (N_24073,N_23670,N_22905);
and U24074 (N_24074,N_23134,N_23311);
and U24075 (N_24075,N_23409,N_23532);
nor U24076 (N_24076,N_22896,N_22910);
nor U24077 (N_24077,N_23099,N_22942);
and U24078 (N_24078,N_23767,N_23563);
xor U24079 (N_24079,N_23241,N_22999);
or U24080 (N_24080,N_23130,N_23375);
nand U24081 (N_24081,N_23798,N_23724);
xnor U24082 (N_24082,N_22956,N_23242);
xor U24083 (N_24083,N_23781,N_23680);
or U24084 (N_24084,N_23072,N_23613);
xnor U24085 (N_24085,N_23005,N_23834);
xnor U24086 (N_24086,N_23089,N_23616);
nor U24087 (N_24087,N_23172,N_23361);
or U24088 (N_24088,N_23108,N_23574);
or U24089 (N_24089,N_23966,N_23611);
nand U24090 (N_24090,N_23791,N_23111);
and U24091 (N_24091,N_23129,N_23849);
xor U24092 (N_24092,N_23292,N_23632);
nor U24093 (N_24093,N_22957,N_23497);
nand U24094 (N_24094,N_23865,N_23100);
and U24095 (N_24095,N_23743,N_22889);
nor U24096 (N_24096,N_23539,N_23989);
nand U24097 (N_24097,N_23101,N_23704);
or U24098 (N_24098,N_23502,N_23779);
nor U24099 (N_24099,N_22826,N_22979);
nand U24100 (N_24100,N_23233,N_22932);
and U24101 (N_24101,N_22902,N_23326);
nor U24102 (N_24102,N_23173,N_23648);
xnor U24103 (N_24103,N_23591,N_23942);
and U24104 (N_24104,N_23203,N_23937);
and U24105 (N_24105,N_23621,N_22884);
and U24106 (N_24106,N_22809,N_23855);
and U24107 (N_24107,N_22920,N_23629);
nand U24108 (N_24108,N_23810,N_23360);
nand U24109 (N_24109,N_22982,N_23689);
or U24110 (N_24110,N_23737,N_23762);
and U24111 (N_24111,N_22996,N_23439);
and U24112 (N_24112,N_23554,N_23122);
or U24113 (N_24113,N_22991,N_23986);
xnor U24114 (N_24114,N_23191,N_23441);
xor U24115 (N_24115,N_23627,N_23165);
xnor U24116 (N_24116,N_22968,N_23535);
and U24117 (N_24117,N_23900,N_23525);
nor U24118 (N_24118,N_23027,N_23754);
and U24119 (N_24119,N_22817,N_22945);
nor U24120 (N_24120,N_23701,N_23026);
xor U24121 (N_24121,N_23578,N_23515);
nor U24122 (N_24122,N_23895,N_23777);
xnor U24123 (N_24123,N_23036,N_23056);
xnor U24124 (N_24124,N_23366,N_23114);
xor U24125 (N_24125,N_23208,N_22974);
xnor U24126 (N_24126,N_23590,N_23536);
and U24127 (N_24127,N_23968,N_23200);
or U24128 (N_24128,N_23459,N_23761);
and U24129 (N_24129,N_22931,N_23716);
nand U24130 (N_24130,N_22997,N_22983);
xor U24131 (N_24131,N_23647,N_23526);
nand U24132 (N_24132,N_22908,N_23857);
nand U24133 (N_24133,N_23572,N_22955);
and U24134 (N_24134,N_22855,N_23169);
or U24135 (N_24135,N_23091,N_23393);
and U24136 (N_24136,N_22978,N_23512);
xnor U24137 (N_24137,N_23469,N_23379);
and U24138 (N_24138,N_22958,N_23848);
and U24139 (N_24139,N_23851,N_23310);
nand U24140 (N_24140,N_23234,N_23853);
xor U24141 (N_24141,N_23164,N_23665);
xor U24142 (N_24142,N_23320,N_23050);
xor U24143 (N_24143,N_23839,N_23858);
xor U24144 (N_24144,N_23715,N_23713);
nor U24145 (N_24145,N_23667,N_23823);
xor U24146 (N_24146,N_23745,N_23885);
nor U24147 (N_24147,N_23596,N_23150);
xnor U24148 (N_24148,N_22811,N_23017);
or U24149 (N_24149,N_22904,N_23321);
xnor U24150 (N_24150,N_23044,N_22933);
and U24151 (N_24151,N_22869,N_22984);
xnor U24152 (N_24152,N_22895,N_22870);
nand U24153 (N_24153,N_23939,N_23482);
nand U24154 (N_24154,N_23421,N_23474);
and U24155 (N_24155,N_23269,N_22954);
nand U24156 (N_24156,N_23308,N_23034);
nor U24157 (N_24157,N_23345,N_22867);
nor U24158 (N_24158,N_22841,N_23544);
or U24159 (N_24159,N_23442,N_23843);
nor U24160 (N_24160,N_23312,N_22969);
xor U24161 (N_24161,N_23628,N_23987);
or U24162 (N_24162,N_22916,N_22857);
and U24163 (N_24163,N_22806,N_23958);
nand U24164 (N_24164,N_23491,N_23437);
or U24165 (N_24165,N_23760,N_23993);
or U24166 (N_24166,N_23362,N_23861);
xnor U24167 (N_24167,N_23496,N_22887);
nor U24168 (N_24168,N_23677,N_23260);
or U24169 (N_24169,N_23157,N_23471);
xor U24170 (N_24170,N_23232,N_23062);
nand U24171 (N_24171,N_23840,N_23445);
nand U24172 (N_24172,N_23370,N_23905);
or U24173 (N_24173,N_23266,N_23207);
and U24174 (N_24174,N_23693,N_23750);
or U24175 (N_24175,N_23247,N_23322);
nand U24176 (N_24176,N_23317,N_22804);
and U24177 (N_24177,N_22898,N_23028);
nor U24178 (N_24178,N_23729,N_23147);
xor U24179 (N_24179,N_23639,N_23151);
and U24180 (N_24180,N_23776,N_23246);
and U24181 (N_24181,N_22812,N_23927);
xnor U24182 (N_24182,N_23112,N_23035);
nor U24183 (N_24183,N_23372,N_23924);
and U24184 (N_24184,N_23119,N_23864);
xnor U24185 (N_24185,N_23076,N_23486);
xnor U24186 (N_24186,N_23603,N_23801);
nor U24187 (N_24187,N_23949,N_22906);
or U24188 (N_24188,N_23505,N_23118);
nor U24189 (N_24189,N_23448,N_23926);
nand U24190 (N_24190,N_22814,N_23371);
xnor U24191 (N_24191,N_23581,N_22847);
and U24192 (N_24192,N_23153,N_22948);
nand U24193 (N_24193,N_23912,N_23047);
nor U24194 (N_24194,N_23218,N_23354);
xor U24195 (N_24195,N_23884,N_23868);
or U24196 (N_24196,N_22810,N_23506);
xor U24197 (N_24197,N_23794,N_23334);
nand U24198 (N_24198,N_23679,N_23614);
nor U24199 (N_24199,N_23065,N_23274);
xor U24200 (N_24200,N_23721,N_23079);
or U24201 (N_24201,N_23774,N_23470);
nand U24202 (N_24202,N_23413,N_23636);
and U24203 (N_24203,N_23981,N_23514);
and U24204 (N_24204,N_23074,N_23874);
nand U24205 (N_24205,N_22886,N_22967);
xnor U24206 (N_24206,N_23131,N_23082);
nand U24207 (N_24207,N_22856,N_22940);
and U24208 (N_24208,N_23640,N_23429);
nor U24209 (N_24209,N_23500,N_23175);
nand U24210 (N_24210,N_23040,N_23492);
or U24211 (N_24211,N_23913,N_23870);
or U24212 (N_24212,N_23195,N_22813);
nand U24213 (N_24213,N_23543,N_23263);
or U24214 (N_24214,N_23720,N_22871);
nand U24215 (N_24215,N_23746,N_23533);
xnor U24216 (N_24216,N_23597,N_22923);
nor U24217 (N_24217,N_23625,N_23013);
nand U24218 (N_24218,N_23400,N_23301);
nand U24219 (N_24219,N_23347,N_23280);
nand U24220 (N_24220,N_23475,N_23285);
and U24221 (N_24221,N_23414,N_22952);
nor U24222 (N_24222,N_23249,N_23768);
xnor U24223 (N_24223,N_23623,N_23407);
and U24224 (N_24224,N_23974,N_23898);
nand U24225 (N_24225,N_23654,N_23318);
or U24226 (N_24226,N_23055,N_23239);
xor U24227 (N_24227,N_22818,N_23527);
and U24228 (N_24228,N_23152,N_23410);
nand U24229 (N_24229,N_23455,N_23243);
and U24230 (N_24230,N_22820,N_23163);
xnor U24231 (N_24231,N_23124,N_23951);
nand U24232 (N_24232,N_23547,N_23261);
and U24233 (N_24233,N_23183,N_23350);
nor U24234 (N_24234,N_23446,N_23943);
and U24235 (N_24235,N_23338,N_23795);
or U24236 (N_24236,N_23197,N_23382);
or U24237 (N_24237,N_23765,N_23336);
and U24238 (N_24238,N_23708,N_23549);
or U24239 (N_24239,N_23256,N_23235);
nand U24240 (N_24240,N_23566,N_23211);
nand U24241 (N_24241,N_22977,N_23349);
and U24242 (N_24242,N_23189,N_23919);
nand U24243 (N_24243,N_23564,N_23930);
xnor U24244 (N_24244,N_23732,N_22962);
xnor U24245 (N_24245,N_22922,N_23524);
or U24246 (N_24246,N_23967,N_23087);
xor U24247 (N_24247,N_23682,N_23793);
nand U24248 (N_24248,N_23999,N_23599);
nor U24249 (N_24249,N_23748,N_23678);
or U24250 (N_24250,N_22947,N_23039);
xor U24251 (N_24251,N_22943,N_23782);
nand U24252 (N_24252,N_22877,N_23819);
xor U24253 (N_24253,N_23841,N_23828);
or U24254 (N_24254,N_23978,N_22935);
or U24255 (N_24255,N_23457,N_23472);
or U24256 (N_24256,N_23620,N_23979);
nand U24257 (N_24257,N_23922,N_23609);
and U24258 (N_24258,N_22842,N_23267);
nor U24259 (N_24259,N_23307,N_23811);
or U24260 (N_24260,N_23341,N_22851);
nor U24261 (N_24261,N_23452,N_23545);
or U24262 (N_24262,N_23977,N_23866);
xor U24263 (N_24263,N_23741,N_23757);
nor U24264 (N_24264,N_23854,N_23646);
nand U24265 (N_24265,N_23068,N_23420);
nor U24266 (N_24266,N_23763,N_23042);
or U24267 (N_24267,N_22854,N_23313);
and U24268 (N_24268,N_23214,N_23148);
nor U24269 (N_24269,N_23863,N_23259);
and U24270 (N_24270,N_23797,N_23161);
xor U24271 (N_24271,N_22998,N_23438);
nand U24272 (N_24272,N_23064,N_23155);
nand U24273 (N_24273,N_23228,N_23641);
and U24274 (N_24274,N_23695,N_23378);
nand U24275 (N_24275,N_23711,N_23916);
nor U24276 (N_24276,N_23758,N_23894);
xnor U24277 (N_24277,N_22832,N_23710);
or U24278 (N_24278,N_23879,N_23883);
and U24279 (N_24279,N_22946,N_23254);
nand U24280 (N_24280,N_22866,N_23504);
or U24281 (N_24281,N_23860,N_22964);
xor U24282 (N_24282,N_23030,N_23755);
xor U24283 (N_24283,N_23236,N_22828);
nor U24284 (N_24284,N_22900,N_23602);
xor U24285 (N_24285,N_23272,N_23178);
xnor U24286 (N_24286,N_23891,N_23899);
and U24287 (N_24287,N_22899,N_23466);
or U24288 (N_24288,N_23580,N_23397);
or U24289 (N_24289,N_23479,N_23552);
and U24290 (N_24290,N_23809,N_23098);
or U24291 (N_24291,N_23953,N_23156);
or U24292 (N_24292,N_23634,N_23339);
and U24293 (N_24293,N_23817,N_23135);
and U24294 (N_24294,N_23402,N_22937);
xnor U24295 (N_24295,N_22836,N_23358);
nor U24296 (N_24296,N_22918,N_23619);
nor U24297 (N_24297,N_22903,N_22863);
nor U24298 (N_24298,N_23830,N_23216);
nor U24299 (N_24299,N_23643,N_23045);
nor U24300 (N_24300,N_23577,N_23009);
nand U24301 (N_24301,N_23273,N_22800);
xnor U24302 (N_24302,N_23676,N_23692);
and U24303 (N_24303,N_22913,N_23271);
or U24304 (N_24304,N_23296,N_23920);
or U24305 (N_24305,N_23411,N_23657);
or U24306 (N_24306,N_23231,N_23896);
nor U24307 (N_24307,N_23003,N_23807);
nand U24308 (N_24308,N_23723,N_22864);
nand U24309 (N_24309,N_22874,N_23770);
nor U24310 (N_24310,N_23008,N_23673);
xor U24311 (N_24311,N_23585,N_23139);
and U24312 (N_24312,N_23262,N_23104);
or U24313 (N_24313,N_23295,N_22850);
and U24314 (N_24314,N_23698,N_23584);
xor U24315 (N_24315,N_23033,N_22915);
xor U24316 (N_24316,N_23029,N_23529);
or U24317 (N_24317,N_23836,N_23735);
xor U24318 (N_24318,N_23826,N_23416);
or U24319 (N_24319,N_23473,N_22926);
and U24320 (N_24320,N_23606,N_23133);
nor U24321 (N_24321,N_23901,N_23346);
or U24322 (N_24322,N_23404,N_23401);
and U24323 (N_24323,N_23752,N_23096);
and U24324 (N_24324,N_23257,N_23290);
nor U24325 (N_24325,N_23867,N_23661);
and U24326 (N_24326,N_23390,N_23510);
and U24327 (N_24327,N_23833,N_23031);
xor U24328 (N_24328,N_23185,N_23969);
xor U24329 (N_24329,N_23303,N_22973);
and U24330 (N_24330,N_22875,N_23001);
xnor U24331 (N_24331,N_23373,N_23534);
and U24332 (N_24332,N_23635,N_23422);
xnor U24333 (N_24333,N_23785,N_23168);
or U24334 (N_24334,N_23921,N_23540);
nor U24335 (N_24335,N_23956,N_22986);
nor U24336 (N_24336,N_22815,N_23058);
nand U24337 (N_24337,N_23204,N_23694);
nor U24338 (N_24338,N_23914,N_23323);
xnor U24339 (N_24339,N_22992,N_23309);
and U24340 (N_24340,N_23998,N_23468);
nor U24341 (N_24341,N_23188,N_23976);
xnor U24342 (N_24342,N_22876,N_22824);
nor U24343 (N_24343,N_23229,N_23283);
xnor U24344 (N_24344,N_22929,N_22819);
and U24345 (N_24345,N_23831,N_23822);
or U24346 (N_24346,N_23363,N_23198);
xor U24347 (N_24347,N_23929,N_23187);
nand U24348 (N_24348,N_23075,N_23381);
nor U24349 (N_24349,N_23764,N_23561);
xnor U24350 (N_24350,N_23624,N_23444);
nand U24351 (N_24351,N_23889,N_22949);
nand U24352 (N_24352,N_23365,N_22843);
or U24353 (N_24353,N_22834,N_23541);
xor U24354 (N_24354,N_23771,N_23294);
or U24355 (N_24355,N_22823,N_23436);
nand U24356 (N_24356,N_22878,N_23049);
or U24357 (N_24357,N_23480,N_23199);
nand U24358 (N_24358,N_23355,N_23041);
or U24359 (N_24359,N_23751,N_23804);
and U24360 (N_24360,N_22885,N_23289);
xor U24361 (N_24361,N_22881,N_23796);
or U24362 (N_24362,N_22912,N_22848);
nor U24363 (N_24363,N_23778,N_23589);
xnor U24364 (N_24364,N_23424,N_23595);
or U24365 (N_24365,N_23742,N_23383);
nor U24366 (N_24366,N_23671,N_23513);
nand U24367 (N_24367,N_23556,N_23730);
xor U24368 (N_24368,N_23842,N_23054);
xor U24369 (N_24369,N_23938,N_23226);
and U24370 (N_24370,N_23024,N_23433);
nor U24371 (N_24371,N_23116,N_22941);
nand U24372 (N_24372,N_23132,N_23980);
and U24373 (N_24373,N_23351,N_22990);
or U24374 (N_24374,N_23688,N_23772);
and U24375 (N_24375,N_23507,N_23481);
xor U24376 (N_24376,N_22893,N_23668);
nand U24377 (N_24377,N_23847,N_23608);
nor U24378 (N_24378,N_23516,N_23872);
nand U24379 (N_24379,N_23982,N_23000);
xor U24380 (N_24380,N_22987,N_23988);
xnor U24381 (N_24381,N_23825,N_23374);
xor U24382 (N_24382,N_22852,N_23838);
or U24383 (N_24383,N_23348,N_22888);
nor U24384 (N_24384,N_23088,N_23061);
and U24385 (N_24385,N_23251,N_23522);
xor U24386 (N_24386,N_22963,N_23655);
nor U24387 (N_24387,N_23722,N_23220);
xnor U24388 (N_24388,N_23631,N_23509);
or U24389 (N_24389,N_23484,N_23652);
nor U24390 (N_24390,N_23955,N_23146);
nand U24391 (N_24391,N_23476,N_22822);
nor U24392 (N_24392,N_23813,N_23542);
and U24393 (N_24393,N_23971,N_23086);
xnor U24394 (N_24394,N_22988,N_23417);
and U24395 (N_24395,N_23718,N_23666);
xnor U24396 (N_24396,N_23586,N_23835);
or U24397 (N_24397,N_23799,N_22936);
xor U24398 (N_24398,N_23703,N_23435);
xor U24399 (N_24399,N_23845,N_23553);
and U24400 (N_24400,N_23642,N_23012);
nand U24401 (N_24401,N_22909,N_23177);
nor U24402 (N_24402,N_23583,N_23369);
or U24403 (N_24403,N_22816,N_23650);
nand U24404 (N_24404,N_23051,N_22859);
xor U24405 (N_24405,N_22808,N_23749);
or U24406 (N_24406,N_23010,N_23908);
or U24407 (N_24407,N_23824,N_23610);
or U24408 (N_24408,N_23945,N_23786);
nand U24409 (N_24409,N_23965,N_23734);
nand U24410 (N_24410,N_23907,N_22839);
xor U24411 (N_24411,N_23431,N_22861);
nor U24412 (N_24412,N_23059,N_23215);
nand U24413 (N_24413,N_23385,N_23477);
nand U24414 (N_24414,N_23219,N_23478);
xnor U24415 (N_24415,N_23569,N_23485);
xor U24416 (N_24416,N_23353,N_23517);
and U24417 (N_24417,N_23601,N_23052);
nand U24418 (N_24418,N_23518,N_23663);
xor U24419 (N_24419,N_22907,N_23174);
or U24420 (N_24420,N_23276,N_23783);
nor U24421 (N_24421,N_23327,N_23357);
nand U24422 (N_24422,N_22892,N_23270);
and U24423 (N_24423,N_23637,N_23690);
nor U24424 (N_24424,N_23253,N_23167);
nand U24425 (N_24425,N_22833,N_23427);
nor U24426 (N_24426,N_23456,N_23659);
and U24427 (N_24427,N_23941,N_22951);
and U24428 (N_24428,N_22801,N_23206);
xor U24429 (N_24429,N_23923,N_23015);
xor U24430 (N_24430,N_23503,N_23519);
nor U24431 (N_24431,N_23709,N_23395);
nand U24432 (N_24432,N_23892,N_22829);
nand U24433 (N_24433,N_23546,N_23275);
xnor U24434 (N_24434,N_23244,N_23560);
and U24435 (N_24435,N_23391,N_23399);
and U24436 (N_24436,N_23240,N_22853);
nand U24437 (N_24437,N_23196,N_23450);
nor U24438 (N_24438,N_23846,N_23973);
nor U24439 (N_24439,N_23377,N_23245);
or U24440 (N_24440,N_22802,N_23406);
or U24441 (N_24441,N_23430,N_22890);
and U24442 (N_24442,N_23837,N_23158);
nand U24443 (N_24443,N_22970,N_23340);
nand U24444 (N_24444,N_23645,N_23996);
xnor U24445 (N_24445,N_23658,N_23862);
and U24446 (N_24446,N_23963,N_23775);
and U24447 (N_24447,N_23284,N_23501);
xor U24448 (N_24448,N_23097,N_23180);
or U24449 (N_24449,N_23342,N_23672);
xnor U24450 (N_24450,N_23818,N_23523);
nor U24451 (N_24451,N_23412,N_23784);
nand U24452 (N_24452,N_23077,N_23802);
xnor U24453 (N_24453,N_23021,N_22981);
nor U24454 (N_24454,N_23415,N_23935);
nor U24455 (N_24455,N_23186,N_23237);
nand U24456 (N_24456,N_22993,N_22953);
xor U24457 (N_24457,N_22862,N_23006);
nor U24458 (N_24458,N_23910,N_23460);
nor U24459 (N_24459,N_23829,N_23143);
nand U24460 (N_24460,N_23449,N_23081);
nand U24461 (N_24461,N_23230,N_23282);
xnor U24462 (N_24462,N_22917,N_23990);
nor U24463 (N_24463,N_23815,N_23140);
nand U24464 (N_24464,N_23329,N_23906);
nor U24465 (N_24465,N_22846,N_23386);
nor U24466 (N_24466,N_23985,N_22807);
nor U24467 (N_24467,N_23992,N_23612);
and U24468 (N_24468,N_23875,N_22927);
and U24469 (N_24469,N_22939,N_23127);
or U24470 (N_24470,N_23940,N_22849);
nand U24471 (N_24471,N_22934,N_22965);
and U24472 (N_24472,N_23171,N_23069);
nor U24473 (N_24473,N_23706,N_23521);
nand U24474 (N_24474,N_23210,N_23936);
and U24475 (N_24475,N_23816,N_23882);
xor U24476 (N_24476,N_23011,N_23812);
nand U24477 (N_24477,N_23306,N_23733);
nor U24478 (N_24478,N_23053,N_23649);
or U24479 (N_24479,N_23859,N_22944);
nor U24480 (N_24480,N_23562,N_23821);
or U24481 (N_24481,N_22960,N_23508);
and U24482 (N_24482,N_22837,N_23110);
nor U24483 (N_24483,N_23367,N_23789);
xor U24484 (N_24484,N_22980,N_23570);
or U24485 (N_24485,N_23707,N_23925);
or U24486 (N_24486,N_23102,N_23094);
or U24487 (N_24487,N_22995,N_23221);
and U24488 (N_24488,N_23739,N_23538);
and U24489 (N_24489,N_23995,N_22835);
xor U24490 (N_24490,N_23037,N_23878);
nor U24491 (N_24491,N_23557,N_23120);
nand U24492 (N_24492,N_23268,N_22975);
or U24493 (N_24493,N_23915,N_23747);
xnor U24494 (N_24494,N_23934,N_22868);
or U24495 (N_24495,N_22966,N_23917);
nor U24496 (N_24496,N_22930,N_23107);
and U24497 (N_24497,N_22911,N_23142);
and U24498 (N_24498,N_23493,N_23113);
nand U24499 (N_24499,N_23852,N_23759);
xnor U24500 (N_24500,N_23753,N_23644);
or U24501 (N_24501,N_23453,N_23071);
xnor U24502 (N_24502,N_22921,N_23396);
and U24503 (N_24503,N_23984,N_23662);
xor U24504 (N_24504,N_23537,N_23387);
nand U24505 (N_24505,N_23356,N_23575);
nor U24506 (N_24506,N_23388,N_23983);
and U24507 (N_24507,N_23238,N_23685);
nor U24508 (N_24508,N_23918,N_23103);
and U24509 (N_24509,N_23095,N_23170);
and U24510 (N_24510,N_23731,N_23587);
and U24511 (N_24511,N_23217,N_22825);
xnor U24512 (N_24512,N_23325,N_23330);
and U24513 (N_24513,N_22989,N_23952);
or U24514 (N_24514,N_23138,N_23638);
and U24515 (N_24515,N_23869,N_22838);
nor U24516 (N_24516,N_23805,N_23176);
nand U24517 (N_24517,N_22883,N_23032);
or U24518 (N_24518,N_22831,N_23043);
nor U24519 (N_24519,N_23972,N_23331);
xnor U24520 (N_24520,N_22865,N_23576);
and U24521 (N_24521,N_23141,N_23063);
and U24522 (N_24522,N_23255,N_23736);
nor U24523 (N_24523,N_22938,N_22844);
nand U24524 (N_24524,N_23293,N_23769);
xor U24525 (N_24525,N_23876,N_23125);
nor U24526 (N_24526,N_22860,N_23975);
nand U24527 (N_24527,N_22803,N_23911);
nor U24528 (N_24528,N_23598,N_23957);
or U24529 (N_24529,N_23205,N_23959);
or U24530 (N_24530,N_23773,N_23565);
nand U24531 (N_24531,N_23954,N_23944);
xnor U24532 (N_24532,N_22994,N_23258);
xor U24533 (N_24533,N_23359,N_23109);
or U24534 (N_24534,N_23933,N_23250);
xor U24535 (N_24535,N_23002,N_23850);
or U24536 (N_24536,N_23490,N_23279);
and U24537 (N_24537,N_23023,N_23827);
and U24538 (N_24538,N_23324,N_23618);
or U24539 (N_24539,N_23700,N_23019);
nand U24540 (N_24540,N_23567,N_23674);
or U24541 (N_24541,N_23675,N_23419);
or U24542 (N_24542,N_23333,N_23314);
nor U24543 (N_24543,N_23950,N_23004);
nor U24544 (N_24544,N_23697,N_23844);
xor U24545 (N_24545,N_23559,N_23060);
and U24546 (N_24546,N_23344,N_23691);
or U24547 (N_24547,N_22985,N_23702);
or U24548 (N_24548,N_23281,N_23686);
or U24549 (N_24549,N_23304,N_23319);
and U24550 (N_24550,N_23287,N_23605);
nand U24551 (N_24551,N_23428,N_23300);
and U24552 (N_24552,N_23487,N_23548);
nor U24553 (N_24553,N_23194,N_23144);
and U24554 (N_24554,N_23264,N_23948);
or U24555 (N_24555,N_23380,N_23531);
or U24556 (N_24556,N_23425,N_23123);
xnor U24557 (N_24557,N_23991,N_23617);
and U24558 (N_24558,N_23073,N_23403);
nand U24559 (N_24559,N_23352,N_23467);
and U24560 (N_24560,N_23728,N_23947);
or U24561 (N_24561,N_23166,N_23705);
xor U24562 (N_24562,N_23626,N_23790);
nand U24563 (N_24563,N_23664,N_23787);
nand U24564 (N_24564,N_23928,N_23162);
and U24565 (N_24565,N_23443,N_22880);
nor U24566 (N_24566,N_23593,N_23128);
and U24567 (N_24567,N_23315,N_23604);
xnor U24568 (N_24568,N_23719,N_23856);
nand U24569 (N_24569,N_23653,N_23286);
nor U24570 (N_24570,N_23248,N_23814);
and U24571 (N_24571,N_23600,N_23181);
or U24572 (N_24572,N_22959,N_22873);
xnor U24573 (N_24573,N_23582,N_23160);
and U24574 (N_24574,N_23154,N_23025);
or U24575 (N_24575,N_22972,N_23714);
and U24576 (N_24576,N_23084,N_23078);
or U24577 (N_24577,N_23451,N_23932);
nor U24578 (N_24578,N_23299,N_23579);
xor U24579 (N_24579,N_23106,N_23571);
and U24580 (N_24580,N_23725,N_23962);
and U24581 (N_24581,N_23105,N_23803);
nor U24582 (N_24582,N_22976,N_23594);
xnor U24583 (N_24583,N_22872,N_23592);
and U24584 (N_24584,N_23681,N_23332);
or U24585 (N_24585,N_23302,N_23368);
nor U24586 (N_24586,N_22879,N_23558);
or U24587 (N_24587,N_22827,N_23184);
or U24588 (N_24588,N_23520,N_23038);
and U24589 (N_24589,N_23458,N_23607);
nand U24590 (N_24590,N_23633,N_23222);
nand U24591 (N_24591,N_23727,N_23278);
xnor U24592 (N_24592,N_22971,N_23083);
or U24593 (N_24593,N_23489,N_22891);
nor U24594 (N_24594,N_23227,N_23780);
nor U24595 (N_24595,N_23961,N_23897);
nor U24596 (N_24596,N_23115,N_23738);
nor U24597 (N_24597,N_23020,N_23871);
nand U24598 (N_24598,N_23740,N_22961);
nand U24599 (N_24599,N_23121,N_23297);
nand U24600 (N_24600,N_23401,N_22973);
xnor U24601 (N_24601,N_23798,N_23905);
nor U24602 (N_24602,N_23620,N_23368);
nor U24603 (N_24603,N_22912,N_23459);
nor U24604 (N_24604,N_23907,N_22882);
nand U24605 (N_24605,N_23747,N_23671);
nor U24606 (N_24606,N_23339,N_23868);
xor U24607 (N_24607,N_23633,N_22998);
or U24608 (N_24608,N_23120,N_23842);
or U24609 (N_24609,N_22939,N_23855);
nor U24610 (N_24610,N_23407,N_23655);
nor U24611 (N_24611,N_23653,N_23409);
xor U24612 (N_24612,N_23816,N_23694);
xor U24613 (N_24613,N_23139,N_23540);
or U24614 (N_24614,N_23035,N_23302);
nor U24615 (N_24615,N_23357,N_23029);
nand U24616 (N_24616,N_23450,N_23523);
xor U24617 (N_24617,N_23646,N_23636);
and U24618 (N_24618,N_23888,N_23363);
xnor U24619 (N_24619,N_23084,N_22904);
nand U24620 (N_24620,N_23000,N_23873);
nor U24621 (N_24621,N_23176,N_23445);
nand U24622 (N_24622,N_22830,N_23532);
nand U24623 (N_24623,N_23315,N_23194);
nand U24624 (N_24624,N_23105,N_22993);
nand U24625 (N_24625,N_23243,N_22811);
nor U24626 (N_24626,N_23886,N_23290);
nand U24627 (N_24627,N_22898,N_23040);
xor U24628 (N_24628,N_23957,N_23368);
and U24629 (N_24629,N_22836,N_23687);
nand U24630 (N_24630,N_23149,N_23539);
xor U24631 (N_24631,N_22956,N_23911);
xor U24632 (N_24632,N_22981,N_23847);
or U24633 (N_24633,N_22823,N_23284);
or U24634 (N_24634,N_22810,N_23752);
xnor U24635 (N_24635,N_23788,N_23905);
nand U24636 (N_24636,N_23591,N_23030);
xor U24637 (N_24637,N_22824,N_23988);
nor U24638 (N_24638,N_22960,N_23881);
nand U24639 (N_24639,N_23074,N_23879);
xnor U24640 (N_24640,N_23660,N_23666);
and U24641 (N_24641,N_23945,N_22844);
nor U24642 (N_24642,N_22801,N_23815);
xnor U24643 (N_24643,N_22800,N_23677);
xor U24644 (N_24644,N_23038,N_22878);
or U24645 (N_24645,N_23320,N_23674);
or U24646 (N_24646,N_23051,N_23614);
nand U24647 (N_24647,N_23732,N_23127);
nor U24648 (N_24648,N_22946,N_23045);
nand U24649 (N_24649,N_23016,N_23533);
xnor U24650 (N_24650,N_23555,N_23316);
xor U24651 (N_24651,N_22807,N_23832);
and U24652 (N_24652,N_23687,N_23108);
and U24653 (N_24653,N_22858,N_22938);
and U24654 (N_24654,N_23127,N_23792);
or U24655 (N_24655,N_23969,N_23005);
nand U24656 (N_24656,N_23607,N_23006);
nand U24657 (N_24657,N_23639,N_23952);
xnor U24658 (N_24658,N_23715,N_22878);
xnor U24659 (N_24659,N_23897,N_23538);
or U24660 (N_24660,N_23760,N_22868);
and U24661 (N_24661,N_23066,N_23897);
and U24662 (N_24662,N_23988,N_22940);
xor U24663 (N_24663,N_23143,N_22962);
or U24664 (N_24664,N_23290,N_23360);
nand U24665 (N_24665,N_23557,N_23815);
nand U24666 (N_24666,N_23699,N_23683);
and U24667 (N_24667,N_23418,N_23825);
xnor U24668 (N_24668,N_23930,N_23948);
or U24669 (N_24669,N_23675,N_23353);
nor U24670 (N_24670,N_22964,N_23917);
or U24671 (N_24671,N_23403,N_23721);
or U24672 (N_24672,N_23913,N_23661);
and U24673 (N_24673,N_23320,N_22880);
nand U24674 (N_24674,N_23848,N_23687);
or U24675 (N_24675,N_23954,N_22954);
and U24676 (N_24676,N_23396,N_22915);
nor U24677 (N_24677,N_23511,N_23277);
xnor U24678 (N_24678,N_23983,N_23015);
or U24679 (N_24679,N_23161,N_23152);
or U24680 (N_24680,N_22863,N_22820);
or U24681 (N_24681,N_23892,N_22905);
or U24682 (N_24682,N_23997,N_23634);
or U24683 (N_24683,N_23783,N_23611);
or U24684 (N_24684,N_23624,N_23842);
and U24685 (N_24685,N_23511,N_23115);
and U24686 (N_24686,N_23713,N_23766);
nand U24687 (N_24687,N_23542,N_23119);
or U24688 (N_24688,N_22894,N_23268);
and U24689 (N_24689,N_23648,N_23193);
nand U24690 (N_24690,N_23549,N_22904);
or U24691 (N_24691,N_22993,N_23033);
and U24692 (N_24692,N_23124,N_23729);
nor U24693 (N_24693,N_23840,N_22905);
or U24694 (N_24694,N_22942,N_22804);
or U24695 (N_24695,N_23431,N_23979);
nand U24696 (N_24696,N_22824,N_23792);
or U24697 (N_24697,N_22856,N_23566);
or U24698 (N_24698,N_23417,N_22930);
nand U24699 (N_24699,N_23035,N_23102);
or U24700 (N_24700,N_23561,N_23157);
or U24701 (N_24701,N_23783,N_23462);
nand U24702 (N_24702,N_23533,N_23321);
nand U24703 (N_24703,N_23022,N_23416);
or U24704 (N_24704,N_23967,N_23261);
or U24705 (N_24705,N_23892,N_23860);
nor U24706 (N_24706,N_23158,N_23727);
xnor U24707 (N_24707,N_22997,N_22906);
or U24708 (N_24708,N_23158,N_22802);
nand U24709 (N_24709,N_23253,N_23453);
or U24710 (N_24710,N_23633,N_23376);
and U24711 (N_24711,N_23195,N_23425);
nor U24712 (N_24712,N_22817,N_23310);
or U24713 (N_24713,N_23288,N_23538);
xnor U24714 (N_24714,N_23634,N_23201);
xnor U24715 (N_24715,N_23525,N_22821);
nor U24716 (N_24716,N_23916,N_23927);
or U24717 (N_24717,N_23846,N_23695);
nand U24718 (N_24718,N_23863,N_23323);
nor U24719 (N_24719,N_23945,N_23411);
nor U24720 (N_24720,N_23824,N_23278);
nor U24721 (N_24721,N_23111,N_23534);
nand U24722 (N_24722,N_22921,N_23414);
xnor U24723 (N_24723,N_23064,N_23329);
and U24724 (N_24724,N_22983,N_23028);
nand U24725 (N_24725,N_23123,N_23882);
xor U24726 (N_24726,N_23104,N_23218);
and U24727 (N_24727,N_23640,N_23424);
nand U24728 (N_24728,N_23975,N_23238);
and U24729 (N_24729,N_23675,N_22930);
nor U24730 (N_24730,N_23356,N_23908);
nor U24731 (N_24731,N_23157,N_23976);
and U24732 (N_24732,N_23247,N_23325);
nor U24733 (N_24733,N_23713,N_23426);
or U24734 (N_24734,N_23629,N_22892);
xnor U24735 (N_24735,N_23892,N_23611);
nor U24736 (N_24736,N_23666,N_23144);
or U24737 (N_24737,N_23522,N_23234);
or U24738 (N_24738,N_23611,N_23324);
or U24739 (N_24739,N_23524,N_23607);
nor U24740 (N_24740,N_22819,N_23247);
or U24741 (N_24741,N_23251,N_23838);
nor U24742 (N_24742,N_23363,N_23871);
and U24743 (N_24743,N_23545,N_23262);
xor U24744 (N_24744,N_23557,N_23349);
or U24745 (N_24745,N_23757,N_22885);
xor U24746 (N_24746,N_23266,N_23364);
or U24747 (N_24747,N_23890,N_23463);
and U24748 (N_24748,N_23011,N_23544);
nor U24749 (N_24749,N_23118,N_23476);
nand U24750 (N_24750,N_23163,N_23090);
and U24751 (N_24751,N_23114,N_23238);
xor U24752 (N_24752,N_23218,N_23061);
xor U24753 (N_24753,N_23028,N_23677);
xor U24754 (N_24754,N_23827,N_23547);
nand U24755 (N_24755,N_23890,N_23095);
and U24756 (N_24756,N_23008,N_23949);
xnor U24757 (N_24757,N_23193,N_23685);
nand U24758 (N_24758,N_23027,N_23714);
xor U24759 (N_24759,N_23878,N_23351);
xor U24760 (N_24760,N_22985,N_22840);
nand U24761 (N_24761,N_23063,N_23545);
nor U24762 (N_24762,N_22988,N_22879);
or U24763 (N_24763,N_23038,N_23061);
nor U24764 (N_24764,N_23219,N_23232);
xnor U24765 (N_24765,N_23817,N_23319);
nor U24766 (N_24766,N_23917,N_23903);
or U24767 (N_24767,N_23994,N_23936);
nor U24768 (N_24768,N_23002,N_23993);
and U24769 (N_24769,N_23762,N_23950);
or U24770 (N_24770,N_23565,N_23169);
nand U24771 (N_24771,N_22981,N_23767);
nand U24772 (N_24772,N_23875,N_23359);
and U24773 (N_24773,N_23251,N_23953);
nand U24774 (N_24774,N_23324,N_23098);
and U24775 (N_24775,N_23198,N_23453);
nand U24776 (N_24776,N_23847,N_23351);
nand U24777 (N_24777,N_23940,N_23832);
xor U24778 (N_24778,N_23697,N_23650);
or U24779 (N_24779,N_23755,N_23096);
or U24780 (N_24780,N_23126,N_23175);
xor U24781 (N_24781,N_23172,N_23077);
or U24782 (N_24782,N_23365,N_22964);
and U24783 (N_24783,N_22990,N_23547);
nand U24784 (N_24784,N_23060,N_22908);
nand U24785 (N_24785,N_22836,N_23904);
nor U24786 (N_24786,N_23145,N_23293);
nand U24787 (N_24787,N_23221,N_23635);
and U24788 (N_24788,N_23704,N_23361);
nor U24789 (N_24789,N_23209,N_23329);
nor U24790 (N_24790,N_22975,N_23011);
nand U24791 (N_24791,N_23083,N_23601);
and U24792 (N_24792,N_23106,N_23587);
nand U24793 (N_24793,N_23252,N_23009);
or U24794 (N_24794,N_23395,N_23659);
xor U24795 (N_24795,N_23501,N_23631);
xor U24796 (N_24796,N_23073,N_23270);
xor U24797 (N_24797,N_23819,N_23850);
nor U24798 (N_24798,N_23704,N_23784);
xnor U24799 (N_24799,N_23211,N_23573);
nor U24800 (N_24800,N_23561,N_23244);
xor U24801 (N_24801,N_23765,N_23615);
nand U24802 (N_24802,N_23048,N_23720);
nand U24803 (N_24803,N_23017,N_23469);
nand U24804 (N_24804,N_23441,N_22999);
nand U24805 (N_24805,N_23568,N_23376);
or U24806 (N_24806,N_23816,N_23264);
or U24807 (N_24807,N_23117,N_23403);
xor U24808 (N_24808,N_23575,N_23224);
and U24809 (N_24809,N_22867,N_23302);
or U24810 (N_24810,N_23875,N_22845);
nor U24811 (N_24811,N_22876,N_22875);
or U24812 (N_24812,N_23356,N_23175);
nand U24813 (N_24813,N_23702,N_22891);
nand U24814 (N_24814,N_23911,N_23445);
and U24815 (N_24815,N_22906,N_23608);
nor U24816 (N_24816,N_23597,N_23666);
nand U24817 (N_24817,N_23639,N_23766);
nand U24818 (N_24818,N_22971,N_23019);
or U24819 (N_24819,N_23305,N_22971);
and U24820 (N_24820,N_23258,N_23869);
nand U24821 (N_24821,N_23608,N_23460);
nand U24822 (N_24822,N_23122,N_23521);
xnor U24823 (N_24823,N_23160,N_23470);
and U24824 (N_24824,N_23537,N_23060);
xnor U24825 (N_24825,N_22869,N_23920);
or U24826 (N_24826,N_23101,N_23695);
or U24827 (N_24827,N_23642,N_22884);
or U24828 (N_24828,N_23842,N_23461);
xnor U24829 (N_24829,N_23385,N_22859);
nor U24830 (N_24830,N_23657,N_23649);
and U24831 (N_24831,N_22801,N_23494);
and U24832 (N_24832,N_23196,N_22844);
or U24833 (N_24833,N_23551,N_23530);
and U24834 (N_24834,N_22911,N_23799);
xor U24835 (N_24835,N_23937,N_23905);
nor U24836 (N_24836,N_22873,N_23999);
or U24837 (N_24837,N_23796,N_23722);
or U24838 (N_24838,N_23119,N_22924);
nand U24839 (N_24839,N_23270,N_23057);
nand U24840 (N_24840,N_23727,N_23751);
nor U24841 (N_24841,N_23075,N_22992);
nand U24842 (N_24842,N_23959,N_23260);
nand U24843 (N_24843,N_23480,N_23736);
xor U24844 (N_24844,N_22874,N_22908);
xnor U24845 (N_24845,N_23137,N_23394);
and U24846 (N_24846,N_23856,N_23459);
and U24847 (N_24847,N_23802,N_23550);
nor U24848 (N_24848,N_23399,N_23658);
nand U24849 (N_24849,N_23958,N_22877);
xor U24850 (N_24850,N_23238,N_23823);
and U24851 (N_24851,N_23769,N_23493);
or U24852 (N_24852,N_23589,N_23656);
nand U24853 (N_24853,N_23352,N_22932);
or U24854 (N_24854,N_23102,N_23608);
xor U24855 (N_24855,N_23527,N_23796);
xor U24856 (N_24856,N_23730,N_23459);
nor U24857 (N_24857,N_22880,N_23568);
nor U24858 (N_24858,N_23616,N_23578);
and U24859 (N_24859,N_23326,N_23685);
nand U24860 (N_24860,N_23423,N_23833);
nand U24861 (N_24861,N_22829,N_23192);
and U24862 (N_24862,N_22897,N_23181);
and U24863 (N_24863,N_23216,N_23355);
xor U24864 (N_24864,N_23029,N_23930);
and U24865 (N_24865,N_23765,N_23632);
and U24866 (N_24866,N_22954,N_23512);
nor U24867 (N_24867,N_23187,N_23665);
or U24868 (N_24868,N_23911,N_23116);
and U24869 (N_24869,N_23785,N_23937);
nand U24870 (N_24870,N_23625,N_23552);
nand U24871 (N_24871,N_23667,N_23988);
nand U24872 (N_24872,N_23439,N_22915);
or U24873 (N_24873,N_23973,N_23447);
nor U24874 (N_24874,N_22921,N_22850);
nand U24875 (N_24875,N_23792,N_23922);
or U24876 (N_24876,N_23421,N_23798);
nor U24877 (N_24877,N_23626,N_23546);
xor U24878 (N_24878,N_23782,N_23346);
xnor U24879 (N_24879,N_22862,N_23212);
nand U24880 (N_24880,N_23775,N_23193);
xor U24881 (N_24881,N_23999,N_23970);
and U24882 (N_24882,N_23305,N_23459);
xor U24883 (N_24883,N_23357,N_23541);
xor U24884 (N_24884,N_23430,N_23836);
and U24885 (N_24885,N_23405,N_23666);
and U24886 (N_24886,N_23554,N_23998);
and U24887 (N_24887,N_23264,N_23430);
or U24888 (N_24888,N_23150,N_23776);
nor U24889 (N_24889,N_23861,N_23348);
nand U24890 (N_24890,N_23419,N_23869);
nand U24891 (N_24891,N_23649,N_23553);
xnor U24892 (N_24892,N_23032,N_23555);
and U24893 (N_24893,N_23237,N_23044);
nand U24894 (N_24894,N_23230,N_22871);
nand U24895 (N_24895,N_23537,N_23853);
or U24896 (N_24896,N_23316,N_23284);
nand U24897 (N_24897,N_23780,N_23334);
and U24898 (N_24898,N_23287,N_23781);
and U24899 (N_24899,N_23362,N_23137);
nor U24900 (N_24900,N_23225,N_23028);
nand U24901 (N_24901,N_23832,N_23643);
or U24902 (N_24902,N_23861,N_23173);
nand U24903 (N_24903,N_23282,N_23943);
or U24904 (N_24904,N_23856,N_23314);
xor U24905 (N_24905,N_23039,N_23452);
or U24906 (N_24906,N_23498,N_22908);
and U24907 (N_24907,N_22853,N_23638);
or U24908 (N_24908,N_23433,N_22809);
nand U24909 (N_24909,N_23306,N_22932);
or U24910 (N_24910,N_23567,N_23288);
xor U24911 (N_24911,N_23218,N_22865);
xnor U24912 (N_24912,N_23970,N_22956);
nor U24913 (N_24913,N_23606,N_23347);
and U24914 (N_24914,N_23618,N_23174);
nand U24915 (N_24915,N_22989,N_23417);
or U24916 (N_24916,N_23715,N_23719);
and U24917 (N_24917,N_23014,N_23336);
nor U24918 (N_24918,N_22973,N_22870);
xor U24919 (N_24919,N_23345,N_23505);
nand U24920 (N_24920,N_23669,N_23138);
or U24921 (N_24921,N_23495,N_23534);
xor U24922 (N_24922,N_22954,N_23319);
nand U24923 (N_24923,N_22827,N_22943);
nor U24924 (N_24924,N_23183,N_23835);
and U24925 (N_24925,N_23531,N_23825);
or U24926 (N_24926,N_23886,N_23659);
xor U24927 (N_24927,N_23738,N_23001);
nor U24928 (N_24928,N_23415,N_22863);
xor U24929 (N_24929,N_22851,N_23469);
nor U24930 (N_24930,N_23366,N_23008);
and U24931 (N_24931,N_22800,N_22908);
nand U24932 (N_24932,N_23692,N_23145);
and U24933 (N_24933,N_23094,N_23635);
or U24934 (N_24934,N_22946,N_23773);
or U24935 (N_24935,N_23255,N_23813);
or U24936 (N_24936,N_23269,N_23355);
xor U24937 (N_24937,N_23002,N_23410);
xnor U24938 (N_24938,N_23094,N_22885);
or U24939 (N_24939,N_22831,N_23685);
nand U24940 (N_24940,N_23595,N_23937);
or U24941 (N_24941,N_22938,N_23159);
nor U24942 (N_24942,N_23000,N_23848);
nor U24943 (N_24943,N_23751,N_23889);
nand U24944 (N_24944,N_23290,N_23593);
nor U24945 (N_24945,N_23541,N_23503);
or U24946 (N_24946,N_23586,N_23058);
and U24947 (N_24947,N_22819,N_22936);
or U24948 (N_24948,N_23666,N_22850);
and U24949 (N_24949,N_23344,N_23084);
and U24950 (N_24950,N_23717,N_23126);
or U24951 (N_24951,N_23682,N_23579);
or U24952 (N_24952,N_23040,N_23695);
nand U24953 (N_24953,N_23936,N_23118);
nor U24954 (N_24954,N_23228,N_23124);
nand U24955 (N_24955,N_23958,N_23524);
xor U24956 (N_24956,N_23462,N_23048);
nor U24957 (N_24957,N_23735,N_23157);
and U24958 (N_24958,N_23878,N_23105);
xor U24959 (N_24959,N_23952,N_23814);
or U24960 (N_24960,N_23196,N_23419);
or U24961 (N_24961,N_23523,N_23706);
nor U24962 (N_24962,N_23072,N_23771);
nor U24963 (N_24963,N_23275,N_22939);
xnor U24964 (N_24964,N_23701,N_22862);
nor U24965 (N_24965,N_23311,N_22934);
or U24966 (N_24966,N_23368,N_23372);
nand U24967 (N_24967,N_23332,N_22826);
nor U24968 (N_24968,N_23139,N_23384);
xnor U24969 (N_24969,N_23113,N_22878);
or U24970 (N_24970,N_23691,N_23535);
and U24971 (N_24971,N_23376,N_22937);
xor U24972 (N_24972,N_23205,N_23364);
nand U24973 (N_24973,N_23794,N_23527);
and U24974 (N_24974,N_22909,N_23377);
nand U24975 (N_24975,N_23151,N_22971);
xnor U24976 (N_24976,N_23536,N_23252);
nor U24977 (N_24977,N_23820,N_23085);
and U24978 (N_24978,N_22842,N_22883);
nand U24979 (N_24979,N_23429,N_23040);
or U24980 (N_24980,N_23249,N_23097);
nand U24981 (N_24981,N_23021,N_23026);
nand U24982 (N_24982,N_23546,N_23111);
xnor U24983 (N_24983,N_22832,N_23744);
and U24984 (N_24984,N_23266,N_23225);
and U24985 (N_24985,N_23756,N_22938);
xnor U24986 (N_24986,N_23084,N_23080);
xnor U24987 (N_24987,N_23147,N_23262);
and U24988 (N_24988,N_23270,N_22940);
and U24989 (N_24989,N_22891,N_23804);
nand U24990 (N_24990,N_23302,N_23412);
and U24991 (N_24991,N_23855,N_23266);
nand U24992 (N_24992,N_23364,N_23460);
and U24993 (N_24993,N_23316,N_23415);
and U24994 (N_24994,N_23510,N_23122);
nor U24995 (N_24995,N_23107,N_23376);
and U24996 (N_24996,N_23343,N_23773);
and U24997 (N_24997,N_22873,N_23266);
nand U24998 (N_24998,N_22848,N_23788);
or U24999 (N_24999,N_23942,N_23206);
and U25000 (N_25000,N_23377,N_23364);
nor U25001 (N_25001,N_23158,N_23583);
or U25002 (N_25002,N_22891,N_23794);
xor U25003 (N_25003,N_23036,N_23437);
and U25004 (N_25004,N_23089,N_22806);
xnor U25005 (N_25005,N_23889,N_23094);
and U25006 (N_25006,N_23528,N_22930);
nor U25007 (N_25007,N_23310,N_23740);
nand U25008 (N_25008,N_23745,N_23837);
or U25009 (N_25009,N_23263,N_23055);
or U25010 (N_25010,N_23091,N_23093);
or U25011 (N_25011,N_23353,N_23025);
nand U25012 (N_25012,N_23547,N_23099);
nand U25013 (N_25013,N_23408,N_23484);
or U25014 (N_25014,N_23907,N_22961);
or U25015 (N_25015,N_23875,N_23692);
and U25016 (N_25016,N_23898,N_23516);
nor U25017 (N_25017,N_23593,N_23515);
xor U25018 (N_25018,N_23480,N_22871);
and U25019 (N_25019,N_23377,N_23313);
nor U25020 (N_25020,N_23738,N_23805);
or U25021 (N_25021,N_23334,N_22978);
or U25022 (N_25022,N_23317,N_23110);
nor U25023 (N_25023,N_23050,N_23137);
xor U25024 (N_25024,N_22988,N_23147);
or U25025 (N_25025,N_23470,N_23916);
or U25026 (N_25026,N_23989,N_23487);
nand U25027 (N_25027,N_23464,N_23212);
nand U25028 (N_25028,N_23086,N_23338);
nor U25029 (N_25029,N_23459,N_23620);
and U25030 (N_25030,N_22993,N_23432);
nand U25031 (N_25031,N_23180,N_22960);
nor U25032 (N_25032,N_22886,N_23959);
xnor U25033 (N_25033,N_23096,N_23445);
nand U25034 (N_25034,N_23160,N_23428);
and U25035 (N_25035,N_23341,N_23338);
xor U25036 (N_25036,N_23771,N_23064);
and U25037 (N_25037,N_23661,N_23793);
nand U25038 (N_25038,N_23295,N_23865);
nor U25039 (N_25039,N_23567,N_23287);
nor U25040 (N_25040,N_23762,N_23401);
and U25041 (N_25041,N_23560,N_23863);
and U25042 (N_25042,N_23328,N_23854);
nor U25043 (N_25043,N_23820,N_23818);
nor U25044 (N_25044,N_23738,N_23270);
or U25045 (N_25045,N_23918,N_22963);
or U25046 (N_25046,N_23868,N_23900);
nand U25047 (N_25047,N_22868,N_23746);
or U25048 (N_25048,N_23940,N_22990);
nand U25049 (N_25049,N_23332,N_23623);
nor U25050 (N_25050,N_23164,N_23793);
or U25051 (N_25051,N_23077,N_23779);
nor U25052 (N_25052,N_23469,N_23117);
or U25053 (N_25053,N_23053,N_23597);
nand U25054 (N_25054,N_23411,N_23467);
nand U25055 (N_25055,N_22846,N_23899);
and U25056 (N_25056,N_23133,N_23966);
and U25057 (N_25057,N_22921,N_23377);
and U25058 (N_25058,N_22933,N_23017);
or U25059 (N_25059,N_23943,N_22944);
xor U25060 (N_25060,N_23233,N_23867);
and U25061 (N_25061,N_22813,N_22848);
or U25062 (N_25062,N_22968,N_23339);
xnor U25063 (N_25063,N_22939,N_23319);
and U25064 (N_25064,N_22948,N_23612);
nor U25065 (N_25065,N_23798,N_23160);
nand U25066 (N_25066,N_22836,N_23626);
nor U25067 (N_25067,N_23075,N_23913);
and U25068 (N_25068,N_23090,N_23725);
nand U25069 (N_25069,N_23223,N_23489);
nand U25070 (N_25070,N_23056,N_23009);
and U25071 (N_25071,N_23167,N_23177);
xor U25072 (N_25072,N_23524,N_23447);
and U25073 (N_25073,N_23155,N_23319);
nor U25074 (N_25074,N_22969,N_23015);
xnor U25075 (N_25075,N_23148,N_23820);
or U25076 (N_25076,N_23149,N_23728);
or U25077 (N_25077,N_22972,N_23539);
nand U25078 (N_25078,N_23999,N_23725);
xor U25079 (N_25079,N_23667,N_23530);
or U25080 (N_25080,N_23517,N_22978);
nor U25081 (N_25081,N_23124,N_23564);
nand U25082 (N_25082,N_23968,N_23957);
or U25083 (N_25083,N_23006,N_23348);
nand U25084 (N_25084,N_23355,N_22970);
xor U25085 (N_25085,N_23206,N_23962);
xnor U25086 (N_25086,N_23923,N_23550);
nand U25087 (N_25087,N_23123,N_23637);
nor U25088 (N_25088,N_23207,N_22891);
xnor U25089 (N_25089,N_23150,N_23676);
xor U25090 (N_25090,N_23856,N_22809);
nand U25091 (N_25091,N_23256,N_22901);
xor U25092 (N_25092,N_23156,N_22912);
or U25093 (N_25093,N_23457,N_23922);
and U25094 (N_25094,N_23813,N_23543);
nand U25095 (N_25095,N_23223,N_23768);
or U25096 (N_25096,N_22973,N_23441);
nand U25097 (N_25097,N_23698,N_23076);
and U25098 (N_25098,N_23904,N_23455);
and U25099 (N_25099,N_23255,N_23242);
or U25100 (N_25100,N_22904,N_22930);
nor U25101 (N_25101,N_23125,N_23394);
or U25102 (N_25102,N_23694,N_23505);
and U25103 (N_25103,N_23990,N_23735);
nor U25104 (N_25104,N_23704,N_22918);
nand U25105 (N_25105,N_22814,N_22935);
nor U25106 (N_25106,N_23811,N_23951);
and U25107 (N_25107,N_23299,N_23629);
nand U25108 (N_25108,N_23322,N_23908);
and U25109 (N_25109,N_22883,N_23479);
nor U25110 (N_25110,N_23027,N_23743);
nor U25111 (N_25111,N_23701,N_23755);
and U25112 (N_25112,N_23964,N_23288);
nand U25113 (N_25113,N_23121,N_23096);
and U25114 (N_25114,N_22928,N_23062);
and U25115 (N_25115,N_23040,N_23326);
nor U25116 (N_25116,N_23360,N_23573);
nand U25117 (N_25117,N_22860,N_23428);
nor U25118 (N_25118,N_23904,N_22991);
nor U25119 (N_25119,N_23588,N_23008);
and U25120 (N_25120,N_23149,N_23378);
or U25121 (N_25121,N_22971,N_23529);
nor U25122 (N_25122,N_23088,N_23211);
nand U25123 (N_25123,N_23086,N_23491);
nand U25124 (N_25124,N_23546,N_23128);
xor U25125 (N_25125,N_23985,N_23472);
or U25126 (N_25126,N_23912,N_23967);
nand U25127 (N_25127,N_23826,N_23453);
and U25128 (N_25128,N_23465,N_23822);
or U25129 (N_25129,N_23164,N_23039);
and U25130 (N_25130,N_22919,N_23569);
and U25131 (N_25131,N_22862,N_23923);
xor U25132 (N_25132,N_23379,N_23149);
nand U25133 (N_25133,N_23732,N_23348);
nand U25134 (N_25134,N_23116,N_23325);
nor U25135 (N_25135,N_23622,N_23792);
xor U25136 (N_25136,N_22983,N_22939);
nand U25137 (N_25137,N_23822,N_22959);
xor U25138 (N_25138,N_22882,N_23393);
and U25139 (N_25139,N_23233,N_23260);
and U25140 (N_25140,N_23115,N_23352);
nor U25141 (N_25141,N_23776,N_23889);
or U25142 (N_25142,N_23933,N_22893);
xnor U25143 (N_25143,N_23441,N_23319);
xor U25144 (N_25144,N_23986,N_23646);
and U25145 (N_25145,N_23592,N_23084);
and U25146 (N_25146,N_23706,N_23003);
or U25147 (N_25147,N_22868,N_22906);
nand U25148 (N_25148,N_23396,N_23788);
or U25149 (N_25149,N_23408,N_23710);
nand U25150 (N_25150,N_23663,N_23858);
or U25151 (N_25151,N_23773,N_23594);
nand U25152 (N_25152,N_23721,N_22831);
nor U25153 (N_25153,N_23969,N_22958);
or U25154 (N_25154,N_23216,N_23869);
and U25155 (N_25155,N_23559,N_23025);
or U25156 (N_25156,N_23793,N_22854);
nand U25157 (N_25157,N_23261,N_23550);
nor U25158 (N_25158,N_23637,N_23075);
nand U25159 (N_25159,N_23863,N_23024);
and U25160 (N_25160,N_23719,N_23026);
xor U25161 (N_25161,N_23165,N_23624);
xnor U25162 (N_25162,N_23762,N_22834);
xnor U25163 (N_25163,N_23534,N_23828);
xnor U25164 (N_25164,N_23368,N_23580);
xor U25165 (N_25165,N_23037,N_23275);
xnor U25166 (N_25166,N_23386,N_23962);
and U25167 (N_25167,N_23679,N_23441);
and U25168 (N_25168,N_23527,N_23642);
or U25169 (N_25169,N_23161,N_23116);
or U25170 (N_25170,N_23405,N_23712);
xor U25171 (N_25171,N_23004,N_23594);
or U25172 (N_25172,N_23707,N_23534);
nor U25173 (N_25173,N_23142,N_23610);
nor U25174 (N_25174,N_23293,N_23260);
xnor U25175 (N_25175,N_23966,N_23523);
or U25176 (N_25176,N_23937,N_23475);
or U25177 (N_25177,N_23672,N_22894);
and U25178 (N_25178,N_23068,N_23641);
xor U25179 (N_25179,N_23232,N_23572);
xor U25180 (N_25180,N_23353,N_23727);
and U25181 (N_25181,N_23711,N_23683);
nand U25182 (N_25182,N_23184,N_23515);
nor U25183 (N_25183,N_23609,N_22971);
nand U25184 (N_25184,N_23128,N_23334);
and U25185 (N_25185,N_23673,N_23693);
xnor U25186 (N_25186,N_23520,N_23474);
and U25187 (N_25187,N_23101,N_22904);
and U25188 (N_25188,N_23386,N_23804);
nor U25189 (N_25189,N_23971,N_23173);
or U25190 (N_25190,N_23774,N_22885);
xor U25191 (N_25191,N_23001,N_23473);
and U25192 (N_25192,N_22821,N_23950);
or U25193 (N_25193,N_23595,N_22956);
nand U25194 (N_25194,N_23223,N_23509);
or U25195 (N_25195,N_22805,N_23878);
nand U25196 (N_25196,N_23619,N_23251);
and U25197 (N_25197,N_23298,N_23254);
or U25198 (N_25198,N_23463,N_23833);
xor U25199 (N_25199,N_23219,N_23812);
nand U25200 (N_25200,N_24684,N_24158);
or U25201 (N_25201,N_25044,N_24065);
or U25202 (N_25202,N_24826,N_24448);
and U25203 (N_25203,N_24904,N_24700);
and U25204 (N_25204,N_24502,N_24841);
or U25205 (N_25205,N_24405,N_24882);
xnor U25206 (N_25206,N_24265,N_25121);
nand U25207 (N_25207,N_24136,N_24352);
xnor U25208 (N_25208,N_24433,N_25034);
or U25209 (N_25209,N_24422,N_24881);
nor U25210 (N_25210,N_25071,N_24141);
xnor U25211 (N_25211,N_24244,N_24368);
xnor U25212 (N_25212,N_25186,N_24095);
and U25213 (N_25213,N_24230,N_24128);
or U25214 (N_25214,N_24913,N_24513);
nor U25215 (N_25215,N_24171,N_24457);
xnor U25216 (N_25216,N_24500,N_25015);
nand U25217 (N_25217,N_24733,N_24454);
nor U25218 (N_25218,N_24002,N_24226);
nand U25219 (N_25219,N_25178,N_24963);
nand U25220 (N_25220,N_24111,N_24617);
nor U25221 (N_25221,N_24253,N_24739);
nor U25222 (N_25222,N_25166,N_24694);
xor U25223 (N_25223,N_25100,N_24523);
xor U25224 (N_25224,N_24059,N_24940);
or U25225 (N_25225,N_24926,N_24183);
nor U25226 (N_25226,N_24706,N_24668);
xnor U25227 (N_25227,N_24315,N_24318);
nor U25228 (N_25228,N_24554,N_24228);
and U25229 (N_25229,N_24595,N_24300);
xnor U25230 (N_25230,N_25056,N_24221);
nor U25231 (N_25231,N_24395,N_24851);
and U25232 (N_25232,N_24919,N_24723);
xor U25233 (N_25233,N_24822,N_24125);
nor U25234 (N_25234,N_24623,N_24567);
xnor U25235 (N_25235,N_24387,N_24943);
and U25236 (N_25236,N_24665,N_24123);
nor U25237 (N_25237,N_24600,N_24051);
and U25238 (N_25238,N_24113,N_25170);
nor U25239 (N_25239,N_24843,N_24467);
and U25240 (N_25240,N_24752,N_24207);
nand U25241 (N_25241,N_24304,N_25079);
xor U25242 (N_25242,N_24363,N_24450);
or U25243 (N_25243,N_24197,N_24890);
nor U25244 (N_25244,N_24515,N_24129);
xnor U25245 (N_25245,N_24252,N_24028);
nand U25246 (N_25246,N_24747,N_24067);
nor U25247 (N_25247,N_24174,N_25132);
xnor U25248 (N_25248,N_25066,N_24869);
xnor U25249 (N_25249,N_24534,N_24414);
xor U25250 (N_25250,N_24885,N_24487);
xor U25251 (N_25251,N_24358,N_24219);
nor U25252 (N_25252,N_24704,N_24858);
and U25253 (N_25253,N_24536,N_25123);
xnor U25254 (N_25254,N_24316,N_24582);
nor U25255 (N_25255,N_24211,N_24026);
or U25256 (N_25256,N_25112,N_24836);
xor U25257 (N_25257,N_24268,N_24692);
xor U25258 (N_25258,N_25025,N_24222);
nand U25259 (N_25259,N_24660,N_25062);
nand U25260 (N_25260,N_24401,N_24996);
or U25261 (N_25261,N_25067,N_25190);
nor U25262 (N_25262,N_25181,N_24463);
xor U25263 (N_25263,N_25131,N_24278);
and U25264 (N_25264,N_24664,N_24772);
or U25265 (N_25265,N_24200,N_25038);
and U25266 (N_25266,N_24017,N_25001);
nor U25267 (N_25267,N_24437,N_24553);
and U25268 (N_25268,N_25115,N_24399);
or U25269 (N_25269,N_24449,N_24066);
nand U25270 (N_25270,N_24371,N_24242);
nand U25271 (N_25271,N_24774,N_24879);
xnor U25272 (N_25272,N_24193,N_24459);
nand U25273 (N_25273,N_24642,N_24055);
or U25274 (N_25274,N_25125,N_24194);
or U25275 (N_25275,N_24181,N_24037);
xor U25276 (N_25276,N_24032,N_24314);
nor U25277 (N_25277,N_24382,N_24683);
nor U25278 (N_25278,N_24864,N_24833);
xor U25279 (N_25279,N_24994,N_24925);
and U25280 (N_25280,N_24409,N_24731);
nand U25281 (N_25281,N_24447,N_24022);
and U25282 (N_25282,N_25084,N_24143);
xnor U25283 (N_25283,N_25091,N_24245);
xnor U25284 (N_25284,N_24276,N_24535);
xor U25285 (N_25285,N_24525,N_24626);
nand U25286 (N_25286,N_24488,N_24816);
or U25287 (N_25287,N_24532,N_24917);
nand U25288 (N_25288,N_24077,N_24896);
nand U25289 (N_25289,N_24991,N_24929);
and U25290 (N_25290,N_25054,N_24044);
nor U25291 (N_25291,N_25046,N_24549);
or U25292 (N_25292,N_24272,N_24894);
or U25293 (N_25293,N_24170,N_24608);
and U25294 (N_25294,N_24381,N_24821);
nand U25295 (N_25295,N_24482,N_25085);
and U25296 (N_25296,N_24884,N_24950);
or U25297 (N_25297,N_24237,N_24182);
nand U25298 (N_25298,N_24935,N_24360);
xor U25299 (N_25299,N_24832,N_24464);
and U25300 (N_25300,N_24990,N_24877);
or U25301 (N_25301,N_25198,N_24819);
or U25302 (N_25302,N_24442,N_24737);
or U25303 (N_25303,N_24485,N_24741);
or U25304 (N_25304,N_24889,N_24845);
nor U25305 (N_25305,N_24875,N_25090);
or U25306 (N_25306,N_24840,N_24186);
nor U25307 (N_25307,N_25134,N_24235);
nand U25308 (N_25308,N_24199,N_24027);
nand U25309 (N_25309,N_25024,N_24231);
or U25310 (N_25310,N_24388,N_24526);
and U25311 (N_25311,N_24472,N_25097);
nor U25312 (N_25312,N_24375,N_24019);
or U25313 (N_25313,N_24941,N_24176);
nand U25314 (N_25314,N_24351,N_24153);
and U25315 (N_25315,N_24758,N_24953);
nor U25316 (N_25316,N_24899,N_24372);
and U25317 (N_25317,N_25154,N_25078);
xnor U25318 (N_25318,N_24920,N_24512);
or U25319 (N_25319,N_24797,N_25087);
xor U25320 (N_25320,N_24520,N_24949);
or U25321 (N_25321,N_24540,N_24932);
nor U25322 (N_25322,N_24234,N_25157);
xor U25323 (N_25323,N_24976,N_24332);
and U25324 (N_25324,N_24178,N_24508);
nand U25325 (N_25325,N_24988,N_24585);
or U25326 (N_25326,N_25013,N_24249);
or U25327 (N_25327,N_24588,N_24987);
xnor U25328 (N_25328,N_24239,N_24719);
and U25329 (N_25329,N_24290,N_25148);
nand U25330 (N_25330,N_24269,N_24112);
and U25331 (N_25331,N_24154,N_24362);
and U25332 (N_25332,N_24313,N_24054);
and U25333 (N_25333,N_24616,N_24808);
xnor U25334 (N_25334,N_24257,N_24630);
nand U25335 (N_25335,N_24813,N_24394);
nand U25336 (N_25336,N_24205,N_24714);
nor U25337 (N_25337,N_24831,N_24560);
or U25338 (N_25338,N_24238,N_24267);
and U25339 (N_25339,N_25068,N_24168);
nor U25340 (N_25340,N_24246,N_24184);
nor U25341 (N_25341,N_24644,N_24411);
nand U25342 (N_25342,N_24736,N_24530);
xnor U25343 (N_25343,N_24201,N_24435);
xnor U25344 (N_25344,N_25057,N_25145);
nand U25345 (N_25345,N_25004,N_25153);
nand U25346 (N_25346,N_24477,N_25027);
and U25347 (N_25347,N_25018,N_24258);
nand U25348 (N_25348,N_24559,N_24287);
and U25349 (N_25349,N_24213,N_24794);
xnor U25350 (N_25350,N_24020,N_24126);
and U25351 (N_25351,N_24860,N_24220);
or U25352 (N_25352,N_24676,N_25088);
nor U25353 (N_25353,N_25060,N_24104);
nor U25354 (N_25354,N_24574,N_24995);
xnor U25355 (N_25355,N_24420,N_24369);
nor U25356 (N_25356,N_24521,N_25127);
nor U25357 (N_25357,N_24192,N_24336);
nor U25358 (N_25358,N_25086,N_24229);
nand U25359 (N_25359,N_25003,N_24685);
nand U25360 (N_25360,N_24357,N_25063);
nand U25361 (N_25361,N_24568,N_24460);
nand U25362 (N_25362,N_24867,N_24264);
or U25363 (N_25363,N_24479,N_24686);
xor U25364 (N_25364,N_25147,N_25017);
xor U25365 (N_25365,N_24277,N_24946);
and U25366 (N_25366,N_25105,N_24654);
or U25367 (N_25367,N_24149,N_24791);
nor U25368 (N_25368,N_24602,N_24757);
or U25369 (N_25369,N_24402,N_24601);
or U25370 (N_25370,N_24106,N_24891);
nand U25371 (N_25371,N_24349,N_24556);
or U25372 (N_25372,N_24274,N_24726);
or U25373 (N_25373,N_24625,N_24528);
or U25374 (N_25374,N_24466,N_24137);
nand U25375 (N_25375,N_25098,N_24338);
nor U25376 (N_25376,N_24783,N_25156);
xor U25377 (N_25377,N_24620,N_24799);
nor U25378 (N_25378,N_24294,N_25159);
nand U25379 (N_25379,N_24016,N_24915);
or U25380 (N_25380,N_24850,N_24591);
or U25381 (N_25381,N_24471,N_24531);
and U25382 (N_25382,N_24425,N_24416);
nand U25383 (N_25383,N_24715,N_24754);
or U25384 (N_25384,N_24190,N_24615);
nand U25385 (N_25385,N_24622,N_24140);
xnor U25386 (N_25386,N_24886,N_24820);
xnor U25387 (N_25387,N_24179,N_24883);
or U25388 (N_25388,N_24273,N_24682);
nor U25389 (N_25389,N_24551,N_25126);
or U25390 (N_25390,N_24426,N_24086);
or U25391 (N_25391,N_24959,N_24476);
and U25392 (N_25392,N_24366,N_24364);
nor U25393 (N_25393,N_24803,N_24418);
and U25394 (N_25394,N_24356,N_24519);
or U25395 (N_25395,N_24501,N_24347);
xor U25396 (N_25396,N_24827,N_24577);
and U25397 (N_25397,N_24857,N_24335);
xnor U25398 (N_25398,N_24818,N_24761);
or U25399 (N_25399,N_24039,N_24350);
nor U25400 (N_25400,N_25043,N_25174);
and U25401 (N_25401,N_24147,N_24599);
or U25402 (N_25402,N_24829,N_24048);
xor U25403 (N_25403,N_24023,N_24480);
or U25404 (N_25404,N_24047,N_24611);
xnor U25405 (N_25405,N_24473,N_24275);
nor U25406 (N_25406,N_25150,N_24470);
or U25407 (N_25407,N_24948,N_24444);
xnor U25408 (N_25408,N_24596,N_24432);
or U25409 (N_25409,N_24765,N_24367);
xor U25410 (N_25410,N_24282,N_25101);
nand U25411 (N_25411,N_24796,N_24456);
and U25412 (N_25412,N_24573,N_24853);
or U25413 (N_25413,N_24339,N_24775);
nand U25414 (N_25414,N_24874,N_24966);
nor U25415 (N_25415,N_25028,N_24308);
xnor U25416 (N_25416,N_24583,N_24795);
nand U25417 (N_25417,N_24353,N_24045);
nor U25418 (N_25418,N_24397,N_25137);
or U25419 (N_25419,N_25073,N_24924);
or U25420 (N_25420,N_25142,N_24053);
and U25421 (N_25421,N_25111,N_24021);
nand U25422 (N_25422,N_24354,N_24981);
nor U25423 (N_25423,N_24155,N_24666);
and U25424 (N_25424,N_24578,N_24090);
nor U25425 (N_25425,N_24063,N_24419);
or U25426 (N_25426,N_24605,N_24421);
nand U25427 (N_25427,N_24825,N_24541);
nand U25428 (N_25428,N_24497,N_24749);
nand U25429 (N_25429,N_24971,N_24687);
xnor U25430 (N_25430,N_25055,N_24955);
nand U25431 (N_25431,N_24546,N_24771);
and U25432 (N_25432,N_24474,N_24438);
and U25433 (N_25433,N_24114,N_24076);
nor U25434 (N_25434,N_24333,N_24289);
nand U25435 (N_25435,N_24727,N_24099);
or U25436 (N_25436,N_24407,N_24345);
nor U25437 (N_25437,N_24041,N_24740);
or U25438 (N_25438,N_24678,N_24029);
and U25439 (N_25439,N_24606,N_24322);
and U25440 (N_25440,N_25050,N_24306);
or U25441 (N_25441,N_24396,N_24744);
nor U25442 (N_25442,N_24293,N_25103);
xor U25443 (N_25443,N_25058,N_24815);
xnor U25444 (N_25444,N_24030,N_24598);
and U25445 (N_25445,N_24280,N_24310);
and U25446 (N_25446,N_24547,N_24163);
nand U25447 (N_25447,N_24580,N_24557);
nor U25448 (N_25448,N_24710,N_24057);
nor U25449 (N_25449,N_25089,N_24101);
nand U25450 (N_25450,N_24597,N_24712);
xnor U25451 (N_25451,N_24956,N_24009);
and U25452 (N_25452,N_24010,N_24074);
or U25453 (N_25453,N_24478,N_25120);
nand U25454 (N_25454,N_24961,N_24458);
nor U25455 (N_25455,N_24814,N_24681);
xnor U25456 (N_25456,N_24575,N_24716);
and U25457 (N_25457,N_24524,N_24571);
nor U25458 (N_25458,N_24812,N_24514);
xor U25459 (N_25459,N_24035,N_24916);
xnor U25460 (N_25460,N_25110,N_24902);
nand U25461 (N_25461,N_25199,N_24689);
xnor U25462 (N_25462,N_24015,N_24581);
xor U25463 (N_25463,N_24297,N_24980);
xor U25464 (N_25464,N_24007,N_24062);
nor U25465 (N_25465,N_25061,N_24124);
and U25466 (N_25466,N_25107,N_25197);
nor U25467 (N_25467,N_24905,N_24378);
nor U25468 (N_25468,N_24227,N_24589);
nor U25469 (N_25469,N_24173,N_24910);
nor U25470 (N_25470,N_24769,N_24992);
and U25471 (N_25471,N_24906,N_24337);
xor U25472 (N_25472,N_24697,N_24653);
nor U25473 (N_25473,N_24871,N_24056);
xnor U25474 (N_25474,N_24495,N_24957);
and U25475 (N_25475,N_24110,N_25032);
nor U25476 (N_25476,N_24504,N_25168);
nand U25477 (N_25477,N_24722,N_24374);
xor U25478 (N_25478,N_24156,N_24713);
nor U25479 (N_25479,N_25011,N_25118);
xor U25480 (N_25480,N_24717,N_25141);
xnor U25481 (N_25481,N_24698,N_24768);
nor U25482 (N_25482,N_25116,N_24001);
nor U25483 (N_25483,N_24105,N_24693);
or U25484 (N_25484,N_24975,N_25000);
xor U25485 (N_25485,N_24970,N_24562);
and U25486 (N_25486,N_24406,N_24983);
or U25487 (N_25487,N_24968,N_24301);
and U25488 (N_25488,N_25042,N_25081);
or U25489 (N_25489,N_25037,N_24824);
or U25490 (N_25490,N_25007,N_24281);
nor U25491 (N_25491,N_24417,N_24198);
xor U25492 (N_25492,N_24341,N_24108);
and U25493 (N_25493,N_24895,N_25104);
or U25494 (N_25494,N_24159,N_25083);
xnor U25495 (N_25495,N_24587,N_24671);
or U25496 (N_25496,N_24636,N_24511);
or U25497 (N_25497,N_24400,N_24172);
and U25498 (N_25498,N_24389,N_24392);
nand U25499 (N_25499,N_24656,N_24675);
and U25500 (N_25500,N_24638,N_24973);
nand U25501 (N_25501,N_24166,N_25039);
xnor U25502 (N_25502,N_24185,N_24552);
xor U25503 (N_25503,N_24109,N_24324);
nor U25504 (N_25504,N_24901,N_25136);
xnor U25505 (N_25505,N_25029,N_24355);
and U25506 (N_25506,N_24548,N_25144);
nand U25507 (N_25507,N_24784,N_25185);
xnor U25508 (N_25508,N_24650,N_24031);
nor U25509 (N_25509,N_24468,N_24251);
nand U25510 (N_25510,N_24586,N_24590);
nor U25511 (N_25511,N_25077,N_24933);
nand U25512 (N_25512,N_24923,N_24380);
nor U25513 (N_25513,N_24319,N_24817);
nor U25514 (N_25514,N_24967,N_24579);
xnor U25515 (N_25515,N_24255,N_24075);
nor U25516 (N_25516,N_24746,N_24061);
and U25517 (N_25517,N_24785,N_24115);
nor U25518 (N_25518,N_24455,N_24751);
nand U25519 (N_25519,N_24064,N_25019);
and U25520 (N_25520,N_24830,N_25128);
nor U25521 (N_25521,N_24927,N_24218);
xnor U25522 (N_25522,N_25026,N_24998);
or U25523 (N_25523,N_24013,N_24809);
nand U25524 (N_25524,N_24759,N_24475);
and U25525 (N_25525,N_24259,N_24699);
nor U25526 (N_25526,N_25187,N_24702);
or U25527 (N_25527,N_24262,N_24564);
xnor U25528 (N_25528,N_25059,N_25020);
xor U25529 (N_25529,N_25163,N_24974);
and U25530 (N_25530,N_24823,N_24499);
or U25531 (N_25531,N_24930,N_24555);
and U25532 (N_25532,N_24365,N_25072);
or U25533 (N_25533,N_24655,N_24707);
nor U25534 (N_25534,N_24730,N_24999);
and U25535 (N_25535,N_24295,N_24688);
or U25536 (N_25536,N_24328,N_24735);
and U25537 (N_25537,N_24142,N_24517);
xnor U25538 (N_25538,N_24073,N_24412);
nand U25539 (N_25539,N_24404,N_25096);
xnor U25540 (N_25540,N_25167,N_25053);
nand U25541 (N_25541,N_24937,N_24743);
nand U25542 (N_25542,N_24776,N_24645);
xnor U25543 (N_25543,N_24872,N_24842);
xor U25544 (N_25544,N_24321,N_24331);
nor U25545 (N_25545,N_25082,N_24806);
or U25546 (N_25546,N_24773,N_24079);
and U25547 (N_25547,N_24627,N_24088);
and U25548 (N_25548,N_24939,N_24811);
nor U25549 (N_25549,N_24903,N_24505);
and U25550 (N_25550,N_24880,N_24732);
xor U25551 (N_25551,N_24091,N_25047);
nor U25552 (N_25552,N_24834,N_24346);
and U25553 (N_25553,N_24005,N_25065);
nor U25554 (N_25554,N_24250,N_25014);
and U25555 (N_25555,N_25035,N_24592);
xnor U25556 (N_25556,N_24718,N_24648);
nand U25557 (N_25557,N_24789,N_24083);
xnor U25558 (N_25558,N_24326,N_24344);
and U25559 (N_25559,N_25064,N_24279);
and U25560 (N_25560,N_24708,N_24068);
nand U25561 (N_25561,N_24152,N_24921);
and U25562 (N_25562,N_25129,N_24240);
xnor U25563 (N_25563,N_24835,N_24084);
xor U25564 (N_25564,N_25161,N_24261);
nor U25565 (N_25565,N_24303,N_24046);
nand U25566 (N_25566,N_24492,N_24146);
nand U25567 (N_25567,N_25138,N_25182);
nand U25568 (N_25568,N_24640,N_24911);
xnor U25569 (N_25569,N_24863,N_24750);
nor U25570 (N_25570,N_24945,N_24214);
or U25571 (N_25571,N_24087,N_24805);
xor U25572 (N_25572,N_24912,N_24018);
nand U25573 (N_25573,N_25033,N_24085);
xor U25574 (N_25574,N_24434,N_24914);
or U25575 (N_25575,N_24868,N_24243);
or U25576 (N_25576,N_24728,N_24134);
nand U25577 (N_25577,N_24558,N_24725);
nor U25578 (N_25578,N_24493,N_24691);
and U25579 (N_25579,N_24217,N_24071);
and U25580 (N_25580,N_25036,N_25094);
nor U25581 (N_25581,N_25114,N_24865);
nor U25582 (N_25582,N_24878,N_24777);
and U25583 (N_25583,N_24139,N_24801);
nand U25584 (N_25584,N_25010,N_24748);
nor U25585 (N_25585,N_24483,N_24311);
and U25586 (N_25586,N_24756,N_24131);
xor U25587 (N_25587,N_24543,N_24424);
nand U25588 (N_25588,N_24340,N_24008);
and U25589 (N_25589,N_24533,N_24361);
and U25590 (N_25590,N_24379,N_24305);
xor U25591 (N_25591,N_24330,N_25099);
and U25592 (N_25592,N_24386,N_24191);
nor U25593 (N_25593,N_24802,N_24936);
xor U25594 (N_25594,N_24846,N_24373);
xor U25595 (N_25595,N_24133,N_24663);
and U25596 (N_25596,N_24167,N_24288);
nor U25597 (N_25597,N_24058,N_25069);
and U25598 (N_25598,N_24177,N_24206);
or U25599 (N_25599,N_24770,N_24078);
and U25600 (N_25600,N_24203,N_24286);
xor U25601 (N_25601,N_25183,N_24703);
xor U25602 (N_25602,N_24119,N_24720);
or U25603 (N_25603,N_24610,N_24122);
and U25604 (N_25604,N_24491,N_25149);
xor U25605 (N_25605,N_24518,N_24069);
or U25606 (N_25606,N_24189,N_25021);
or U25607 (N_25607,N_24624,N_25113);
or U25608 (N_25608,N_24673,N_24270);
nor U25609 (N_25609,N_24307,N_24667);
xnor U25610 (N_25610,N_24161,N_24006);
and U25611 (N_25611,N_24603,N_25171);
xor U25612 (N_25612,N_25108,N_25052);
and U25613 (N_25613,N_24652,N_25175);
and U25614 (N_25614,N_24538,N_24979);
nor U25615 (N_25615,N_24408,N_24393);
nand U25616 (N_25616,N_24873,N_24679);
nand U25617 (N_25617,N_25023,N_24753);
nand U25618 (N_25618,N_24978,N_25122);
nand U25619 (N_25619,N_24223,N_24888);
xor U25620 (N_25620,N_24036,N_24516);
xor U25621 (N_25621,N_24745,N_24539);
and U25622 (N_25622,N_24762,N_24484);
and U25623 (N_25623,N_25002,N_24439);
xor U25624 (N_25624,N_24096,N_25176);
and U25625 (N_25625,N_24696,N_25133);
nor U25626 (N_25626,N_24529,N_24012);
nand U25627 (N_25627,N_24612,N_24210);
nand U25628 (N_25628,N_25070,N_24132);
or U25629 (N_25629,N_25092,N_24942);
and U25630 (N_25630,N_24861,N_24343);
nor U25631 (N_25631,N_24446,N_24734);
or U25632 (N_25632,N_24897,N_24248);
nor U25633 (N_25633,N_24285,N_24537);
nor U25634 (N_25634,N_24481,N_24680);
nor U25635 (N_25635,N_24283,N_25106);
or U25636 (N_25636,N_24431,N_25095);
xnor U25637 (N_25637,N_25160,N_24320);
nor U25638 (N_25638,N_24195,N_24157);
and U25639 (N_25639,N_24103,N_24609);
nor U25640 (N_25640,N_24164,N_24342);
or U25641 (N_25641,N_25189,N_25045);
and U25642 (N_25642,N_24893,N_24145);
and U25643 (N_25643,N_25165,N_25009);
xnor U25644 (N_25644,N_24080,N_24498);
and U25645 (N_25645,N_24325,N_25031);
nand U25646 (N_25646,N_24451,N_24410);
nand U25647 (N_25647,N_25164,N_24000);
xor U25648 (N_25648,N_24993,N_24461);
xor U25649 (N_25649,N_24862,N_24024);
and U25650 (N_25650,N_24790,N_24089);
nand U25651 (N_25651,N_24180,N_24788);
nor U25652 (N_25652,N_25093,N_24507);
xor U25653 (N_25653,N_24565,N_25143);
or U25654 (N_25654,N_24093,N_24490);
nor U25655 (N_25655,N_25173,N_24954);
nor U25656 (N_25656,N_24003,N_25117);
xnor U25657 (N_25657,N_24570,N_24254);
xnor U25658 (N_25658,N_24398,N_24951);
xnor U25659 (N_25659,N_24839,N_24900);
nand U25660 (N_25660,N_24208,N_24440);
xor U25661 (N_25661,N_24317,N_24649);
or U25662 (N_25662,N_24637,N_24849);
nand U25663 (N_25663,N_25139,N_24677);
nor U25664 (N_25664,N_24989,N_25193);
or U25665 (N_25665,N_25191,N_25196);
nand U25666 (N_25666,N_24972,N_24510);
xnor U25667 (N_25667,N_24844,N_24496);
or U25668 (N_25668,N_24632,N_24204);
xor U25669 (N_25669,N_24385,N_24506);
or U25670 (N_25670,N_24327,N_24323);
and U25671 (N_25671,N_25162,N_24938);
xor U25672 (N_25672,N_25109,N_25102);
and U25673 (N_25673,N_24641,N_24070);
or U25674 (N_25674,N_24670,N_24033);
nor U25675 (N_25675,N_24838,N_24962);
nand U25676 (N_25676,N_24550,N_24052);
nor U25677 (N_25677,N_24787,N_24561);
nand U25678 (N_25678,N_24527,N_24292);
or U25679 (N_25679,N_24465,N_24705);
xor U25680 (N_25680,N_25184,N_24494);
or U25681 (N_25681,N_24120,N_24800);
or U25682 (N_25682,N_25146,N_24618);
and U25683 (N_25683,N_24629,N_24870);
and U25684 (N_25684,N_24709,N_24907);
or U25685 (N_25685,N_24828,N_24233);
or U25686 (N_25686,N_24247,N_24049);
xnor U25687 (N_25687,N_24130,N_24212);
xnor U25688 (N_25688,N_25192,N_24782);
or U25689 (N_25689,N_24441,N_24025);
or U25690 (N_25690,N_24856,N_24376);
and U25691 (N_25691,N_24760,N_24659);
xnor U25692 (N_25692,N_25006,N_24302);
nor U25693 (N_25693,N_24584,N_24763);
and U25694 (N_25694,N_24639,N_24038);
nor U25695 (N_25695,N_24377,N_24430);
and U25696 (N_25696,N_24415,N_24876);
or U25697 (N_25697,N_24072,N_24766);
and U25698 (N_25698,N_24778,N_24004);
nand U25699 (N_25699,N_24931,N_24082);
xor U25700 (N_25700,N_24651,N_24793);
nor U25701 (N_25701,N_24764,N_24162);
xnor U25702 (N_25702,N_25048,N_24138);
xnor U25703 (N_25703,N_24810,N_24423);
xor U25704 (N_25704,N_24779,N_24545);
nand U25705 (N_25705,N_24042,N_24014);
or U25706 (N_25706,N_24569,N_24701);
or U25707 (N_25707,N_24224,N_24209);
nor U25708 (N_25708,N_24271,N_25140);
and U25709 (N_25709,N_25151,N_24175);
nor U25710 (N_25710,N_24909,N_24798);
xor U25711 (N_25711,N_24117,N_24984);
nand U25712 (N_25712,N_25012,N_24135);
xor U25713 (N_25713,N_24724,N_24786);
or U25714 (N_25714,N_24804,N_24160);
xor U25715 (N_25715,N_24284,N_24594);
or U25716 (N_25716,N_24960,N_24628);
nor U25717 (N_25717,N_24661,N_24848);
xnor U25718 (N_25718,N_24118,N_24619);
or U25719 (N_25719,N_24631,N_24633);
nor U25720 (N_25720,N_24121,N_24256);
and U25721 (N_25721,N_24098,N_24621);
xor U25722 (N_25722,N_24944,N_24428);
nor U25723 (N_25723,N_24542,N_25074);
nor U25724 (N_25724,N_25179,N_24196);
nand U25725 (N_25725,N_24729,N_24662);
nor U25726 (N_25726,N_24266,N_24165);
or U25727 (N_25727,N_24509,N_24982);
and U25728 (N_25728,N_24898,N_25041);
nand U25729 (N_25729,N_24672,N_24081);
nand U25730 (N_25730,N_24225,N_24384);
nor U25731 (N_25731,N_24572,N_24593);
and U25732 (N_25732,N_24958,N_24607);
and U25733 (N_25733,N_24767,N_24859);
nand U25734 (N_25734,N_24922,N_24711);
and U25735 (N_25735,N_25040,N_24780);
nand U25736 (N_25736,N_25016,N_24383);
or U25737 (N_25737,N_24847,N_24260);
nand U25738 (N_25738,N_24427,N_24390);
nor U25739 (N_25739,N_25152,N_24965);
and U25740 (N_25740,N_25005,N_24443);
or U25741 (N_25741,N_24486,N_24034);
nand U25742 (N_25742,N_25080,N_24102);
xnor U25743 (N_25743,N_25075,N_24403);
nand U25744 (N_25744,N_24522,N_25180);
nor U25745 (N_25745,N_25130,N_25177);
nand U25746 (N_25746,N_24050,N_24148);
nor U25747 (N_25747,N_24236,N_24646);
and U25748 (N_25748,N_25188,N_24348);
and U25749 (N_25749,N_24969,N_25022);
and U25750 (N_25750,N_24908,N_24216);
nor U25751 (N_25751,N_24263,N_24738);
nand U25752 (N_25752,N_24934,N_24097);
or U25753 (N_25753,N_24312,N_24566);
nand U25754 (N_25754,N_24997,N_24635);
xnor U25755 (N_25755,N_24643,N_24309);
or U25756 (N_25756,N_24299,N_24116);
xnor U25757 (N_25757,N_25155,N_24855);
and U25758 (N_25758,N_24391,N_24429);
nand U25759 (N_25759,N_24202,N_24043);
or U25760 (N_25760,N_24469,N_24887);
nor U25761 (N_25761,N_24792,N_24452);
nand U25762 (N_25762,N_24151,N_24918);
xnor U25763 (N_25763,N_24866,N_24695);
or U25764 (N_25764,N_24755,N_24503);
xor U25765 (N_25765,N_25119,N_24674);
xnor U25766 (N_25766,N_25135,N_24604);
nor U25767 (N_25767,N_24011,N_25124);
nand U25768 (N_25768,N_25169,N_24462);
xor U25769 (N_25769,N_24144,N_24092);
xnor U25770 (N_25770,N_24544,N_25076);
nand U25771 (N_25771,N_24647,N_24169);
nand U25772 (N_25772,N_24977,N_24329);
and U25773 (N_25773,N_24947,N_24298);
nand U25774 (N_25774,N_24150,N_24964);
nor U25775 (N_25775,N_25030,N_24187);
nor U25776 (N_25776,N_24781,N_24952);
or U25777 (N_25777,N_24040,N_24614);
or U25778 (N_25778,N_24296,N_24985);
nand U25779 (N_25779,N_24232,N_24986);
xnor U25780 (N_25780,N_24854,N_24094);
xnor U25781 (N_25781,N_24489,N_24928);
nor U25782 (N_25782,N_24291,N_24436);
or U25783 (N_25783,N_24634,N_25194);
and U25784 (N_25784,N_25008,N_24188);
and U25785 (N_25785,N_25158,N_24690);
or U25786 (N_25786,N_24359,N_24892);
and U25787 (N_25787,N_25051,N_24413);
or U25788 (N_25788,N_25172,N_25195);
nor U25789 (N_25789,N_24445,N_24576);
and U25790 (N_25790,N_24241,N_24721);
xnor U25791 (N_25791,N_24334,N_24127);
nand U25792 (N_25792,N_24613,N_24742);
and U25793 (N_25793,N_24215,N_24453);
xnor U25794 (N_25794,N_24837,N_24107);
and U25795 (N_25795,N_24669,N_24100);
nor U25796 (N_25796,N_24370,N_24060);
nand U25797 (N_25797,N_25049,N_24563);
nor U25798 (N_25798,N_24657,N_24807);
and U25799 (N_25799,N_24658,N_24852);
nor U25800 (N_25800,N_24918,N_24909);
nor U25801 (N_25801,N_24808,N_24582);
xnor U25802 (N_25802,N_25117,N_24865);
or U25803 (N_25803,N_24729,N_25033);
or U25804 (N_25804,N_24992,N_24732);
nor U25805 (N_25805,N_24023,N_24012);
or U25806 (N_25806,N_24733,N_24535);
nand U25807 (N_25807,N_25156,N_24996);
or U25808 (N_25808,N_24498,N_24173);
xnor U25809 (N_25809,N_24882,N_24642);
xor U25810 (N_25810,N_24724,N_24153);
nand U25811 (N_25811,N_24552,N_24755);
or U25812 (N_25812,N_24073,N_24588);
nor U25813 (N_25813,N_25122,N_24854);
or U25814 (N_25814,N_25178,N_24780);
and U25815 (N_25815,N_24445,N_24548);
xor U25816 (N_25816,N_24569,N_24426);
or U25817 (N_25817,N_24812,N_24932);
or U25818 (N_25818,N_24319,N_24678);
xor U25819 (N_25819,N_24028,N_25051);
xnor U25820 (N_25820,N_24844,N_24734);
or U25821 (N_25821,N_24007,N_25136);
nand U25822 (N_25822,N_24887,N_24713);
or U25823 (N_25823,N_24814,N_24866);
or U25824 (N_25824,N_24589,N_24969);
and U25825 (N_25825,N_24652,N_25010);
nor U25826 (N_25826,N_25079,N_25085);
xor U25827 (N_25827,N_24134,N_25060);
xor U25828 (N_25828,N_24573,N_24791);
nor U25829 (N_25829,N_25127,N_24470);
xnor U25830 (N_25830,N_24610,N_24580);
and U25831 (N_25831,N_25137,N_24082);
and U25832 (N_25832,N_25145,N_24377);
or U25833 (N_25833,N_24589,N_24148);
nand U25834 (N_25834,N_25188,N_24615);
nand U25835 (N_25835,N_24099,N_24139);
or U25836 (N_25836,N_24730,N_24447);
nand U25837 (N_25837,N_24105,N_24088);
xor U25838 (N_25838,N_24073,N_24956);
or U25839 (N_25839,N_24422,N_24920);
xnor U25840 (N_25840,N_24149,N_24191);
nor U25841 (N_25841,N_24706,N_24563);
nor U25842 (N_25842,N_24264,N_25100);
nor U25843 (N_25843,N_24363,N_24794);
nor U25844 (N_25844,N_25161,N_24332);
xnor U25845 (N_25845,N_24848,N_24895);
nor U25846 (N_25846,N_24353,N_24441);
nand U25847 (N_25847,N_24298,N_24646);
or U25848 (N_25848,N_24470,N_24844);
nand U25849 (N_25849,N_24723,N_24077);
or U25850 (N_25850,N_24165,N_25091);
nand U25851 (N_25851,N_24383,N_24550);
nand U25852 (N_25852,N_24217,N_24390);
or U25853 (N_25853,N_24803,N_24675);
xnor U25854 (N_25854,N_24243,N_25038);
xor U25855 (N_25855,N_24475,N_24876);
or U25856 (N_25856,N_24049,N_24795);
or U25857 (N_25857,N_24433,N_25187);
nand U25858 (N_25858,N_24649,N_25182);
nor U25859 (N_25859,N_25131,N_24552);
nand U25860 (N_25860,N_24393,N_25014);
and U25861 (N_25861,N_24036,N_24271);
nor U25862 (N_25862,N_24698,N_24572);
and U25863 (N_25863,N_24007,N_25097);
or U25864 (N_25864,N_25046,N_24735);
nand U25865 (N_25865,N_24653,N_24685);
and U25866 (N_25866,N_24721,N_24874);
nor U25867 (N_25867,N_24602,N_24945);
xor U25868 (N_25868,N_24626,N_25145);
xor U25869 (N_25869,N_24793,N_24455);
and U25870 (N_25870,N_24471,N_24221);
xor U25871 (N_25871,N_24833,N_24134);
or U25872 (N_25872,N_25068,N_24178);
nor U25873 (N_25873,N_25193,N_24039);
nor U25874 (N_25874,N_24656,N_24245);
xor U25875 (N_25875,N_24529,N_24585);
xor U25876 (N_25876,N_24688,N_24518);
nand U25877 (N_25877,N_25057,N_25113);
nor U25878 (N_25878,N_24035,N_24954);
xnor U25879 (N_25879,N_24004,N_24724);
or U25880 (N_25880,N_25167,N_25060);
nand U25881 (N_25881,N_25169,N_24544);
and U25882 (N_25882,N_24033,N_24682);
nor U25883 (N_25883,N_24904,N_24793);
xor U25884 (N_25884,N_24079,N_24399);
nand U25885 (N_25885,N_24405,N_25019);
and U25886 (N_25886,N_24544,N_24791);
xnor U25887 (N_25887,N_24739,N_25056);
nor U25888 (N_25888,N_24196,N_24361);
and U25889 (N_25889,N_24729,N_24691);
nand U25890 (N_25890,N_24910,N_24792);
xor U25891 (N_25891,N_24948,N_24166);
nor U25892 (N_25892,N_24981,N_24079);
and U25893 (N_25893,N_24062,N_24999);
nor U25894 (N_25894,N_24239,N_24819);
xor U25895 (N_25895,N_24234,N_24440);
or U25896 (N_25896,N_24018,N_24100);
xor U25897 (N_25897,N_24881,N_24247);
nor U25898 (N_25898,N_24407,N_24743);
nor U25899 (N_25899,N_24543,N_24648);
nand U25900 (N_25900,N_24223,N_24597);
xor U25901 (N_25901,N_24086,N_24639);
or U25902 (N_25902,N_24706,N_24769);
or U25903 (N_25903,N_25175,N_24599);
nor U25904 (N_25904,N_24679,N_24977);
xnor U25905 (N_25905,N_24728,N_25089);
nor U25906 (N_25906,N_24542,N_24066);
or U25907 (N_25907,N_24647,N_24822);
xnor U25908 (N_25908,N_24597,N_24695);
and U25909 (N_25909,N_24371,N_24195);
nor U25910 (N_25910,N_24891,N_25099);
xnor U25911 (N_25911,N_24289,N_24856);
or U25912 (N_25912,N_24273,N_24608);
nand U25913 (N_25913,N_24566,N_24045);
and U25914 (N_25914,N_24680,N_24154);
or U25915 (N_25915,N_24075,N_24893);
or U25916 (N_25916,N_24386,N_24972);
nand U25917 (N_25917,N_24922,N_24509);
and U25918 (N_25918,N_24338,N_24508);
nand U25919 (N_25919,N_24100,N_25107);
or U25920 (N_25920,N_24441,N_24101);
nand U25921 (N_25921,N_24721,N_25126);
and U25922 (N_25922,N_24057,N_24531);
nor U25923 (N_25923,N_25142,N_24876);
or U25924 (N_25924,N_24139,N_24405);
or U25925 (N_25925,N_24476,N_24328);
and U25926 (N_25926,N_24450,N_24881);
and U25927 (N_25927,N_24458,N_24392);
nand U25928 (N_25928,N_24974,N_24510);
xor U25929 (N_25929,N_24758,N_24097);
nor U25930 (N_25930,N_24856,N_24769);
nor U25931 (N_25931,N_25173,N_25163);
nand U25932 (N_25932,N_24953,N_24423);
xor U25933 (N_25933,N_24574,N_24287);
and U25934 (N_25934,N_24129,N_24955);
and U25935 (N_25935,N_24728,N_24876);
and U25936 (N_25936,N_25012,N_24017);
and U25937 (N_25937,N_24890,N_24053);
and U25938 (N_25938,N_24101,N_25136);
or U25939 (N_25939,N_24298,N_25010);
or U25940 (N_25940,N_24160,N_24221);
nand U25941 (N_25941,N_24550,N_24610);
or U25942 (N_25942,N_24358,N_24184);
and U25943 (N_25943,N_24938,N_24192);
nor U25944 (N_25944,N_24754,N_25091);
nand U25945 (N_25945,N_25146,N_24376);
nor U25946 (N_25946,N_24274,N_24772);
nor U25947 (N_25947,N_24570,N_24346);
and U25948 (N_25948,N_24754,N_24758);
xnor U25949 (N_25949,N_24695,N_24693);
nor U25950 (N_25950,N_24389,N_24017);
nor U25951 (N_25951,N_24811,N_24406);
nand U25952 (N_25952,N_25029,N_24154);
and U25953 (N_25953,N_24452,N_24701);
nor U25954 (N_25954,N_24267,N_24717);
xnor U25955 (N_25955,N_24838,N_25120);
and U25956 (N_25956,N_24599,N_24628);
xor U25957 (N_25957,N_24735,N_25011);
xor U25958 (N_25958,N_24981,N_24836);
or U25959 (N_25959,N_24851,N_24158);
or U25960 (N_25960,N_24120,N_24294);
xor U25961 (N_25961,N_24412,N_24284);
nand U25962 (N_25962,N_24069,N_24153);
nand U25963 (N_25963,N_24458,N_24873);
or U25964 (N_25964,N_24031,N_24318);
and U25965 (N_25965,N_24133,N_24899);
nand U25966 (N_25966,N_24606,N_24991);
nand U25967 (N_25967,N_24722,N_24795);
or U25968 (N_25968,N_24348,N_24475);
and U25969 (N_25969,N_25037,N_24366);
xor U25970 (N_25970,N_25142,N_24807);
nand U25971 (N_25971,N_24904,N_25129);
or U25972 (N_25972,N_25055,N_24375);
and U25973 (N_25973,N_24537,N_25127);
xor U25974 (N_25974,N_25117,N_24661);
xnor U25975 (N_25975,N_24873,N_25138);
xor U25976 (N_25976,N_24103,N_24249);
nand U25977 (N_25977,N_24411,N_24545);
or U25978 (N_25978,N_24068,N_24829);
nor U25979 (N_25979,N_24383,N_24057);
and U25980 (N_25980,N_24874,N_24517);
and U25981 (N_25981,N_24036,N_24064);
and U25982 (N_25982,N_24701,N_24965);
and U25983 (N_25983,N_24203,N_24701);
nor U25984 (N_25984,N_24429,N_24266);
and U25985 (N_25985,N_24821,N_24908);
nand U25986 (N_25986,N_24295,N_24070);
xnor U25987 (N_25987,N_24651,N_24339);
and U25988 (N_25988,N_24588,N_24629);
nand U25989 (N_25989,N_24728,N_25076);
xor U25990 (N_25990,N_24134,N_25135);
xor U25991 (N_25991,N_24338,N_25084);
and U25992 (N_25992,N_24043,N_24094);
xor U25993 (N_25993,N_24680,N_24510);
nor U25994 (N_25994,N_24712,N_24547);
nand U25995 (N_25995,N_24128,N_24396);
xnor U25996 (N_25996,N_24829,N_24239);
nand U25997 (N_25997,N_24223,N_24623);
and U25998 (N_25998,N_24309,N_24195);
xnor U25999 (N_25999,N_24082,N_24018);
xnor U26000 (N_26000,N_24353,N_24355);
xor U26001 (N_26001,N_24864,N_24952);
nand U26002 (N_26002,N_25114,N_24635);
xnor U26003 (N_26003,N_24292,N_24609);
or U26004 (N_26004,N_24221,N_24878);
xnor U26005 (N_26005,N_24877,N_25094);
or U26006 (N_26006,N_24835,N_24984);
or U26007 (N_26007,N_24158,N_24653);
nor U26008 (N_26008,N_24795,N_24075);
or U26009 (N_26009,N_24308,N_24297);
nand U26010 (N_26010,N_25118,N_24494);
xor U26011 (N_26011,N_24549,N_24889);
nand U26012 (N_26012,N_25174,N_24233);
xnor U26013 (N_26013,N_24590,N_25088);
or U26014 (N_26014,N_25092,N_25158);
nand U26015 (N_26015,N_24988,N_24997);
and U26016 (N_26016,N_24741,N_24726);
or U26017 (N_26017,N_24642,N_24139);
or U26018 (N_26018,N_24048,N_24175);
nor U26019 (N_26019,N_24223,N_24298);
xor U26020 (N_26020,N_24065,N_24142);
nor U26021 (N_26021,N_24976,N_24225);
nand U26022 (N_26022,N_24549,N_24782);
xnor U26023 (N_26023,N_24213,N_24477);
nand U26024 (N_26024,N_24822,N_24054);
and U26025 (N_26025,N_25055,N_24305);
xor U26026 (N_26026,N_24504,N_24686);
nand U26027 (N_26027,N_24854,N_24003);
nor U26028 (N_26028,N_25053,N_24060);
xor U26029 (N_26029,N_24067,N_24302);
xnor U26030 (N_26030,N_24924,N_24316);
nor U26031 (N_26031,N_24527,N_24758);
or U26032 (N_26032,N_24227,N_25073);
xor U26033 (N_26033,N_24340,N_24880);
nand U26034 (N_26034,N_24420,N_24216);
xnor U26035 (N_26035,N_24664,N_24442);
xnor U26036 (N_26036,N_24373,N_24038);
xnor U26037 (N_26037,N_25175,N_24629);
or U26038 (N_26038,N_24382,N_24373);
nor U26039 (N_26039,N_24587,N_24254);
nand U26040 (N_26040,N_24406,N_24425);
nand U26041 (N_26041,N_24085,N_24665);
nor U26042 (N_26042,N_25197,N_25186);
nor U26043 (N_26043,N_24250,N_24053);
nor U26044 (N_26044,N_24861,N_24416);
nand U26045 (N_26045,N_24585,N_24820);
nand U26046 (N_26046,N_24476,N_24001);
xor U26047 (N_26047,N_24732,N_24224);
xor U26048 (N_26048,N_24826,N_24843);
and U26049 (N_26049,N_24352,N_25067);
nand U26050 (N_26050,N_24131,N_24494);
xor U26051 (N_26051,N_25139,N_24212);
and U26052 (N_26052,N_24403,N_24751);
or U26053 (N_26053,N_24762,N_24029);
or U26054 (N_26054,N_24225,N_24650);
and U26055 (N_26055,N_24621,N_24981);
or U26056 (N_26056,N_24763,N_25131);
or U26057 (N_26057,N_24848,N_25123);
nor U26058 (N_26058,N_24930,N_24209);
xnor U26059 (N_26059,N_24476,N_24568);
nand U26060 (N_26060,N_24138,N_24826);
nand U26061 (N_26061,N_24414,N_24309);
or U26062 (N_26062,N_24149,N_24145);
or U26063 (N_26063,N_24833,N_24012);
xnor U26064 (N_26064,N_24879,N_24315);
nand U26065 (N_26065,N_24680,N_24783);
or U26066 (N_26066,N_24537,N_24602);
nand U26067 (N_26067,N_25165,N_25113);
and U26068 (N_26068,N_24974,N_24642);
nor U26069 (N_26069,N_24671,N_24602);
or U26070 (N_26070,N_24283,N_24861);
xnor U26071 (N_26071,N_24544,N_24147);
xnor U26072 (N_26072,N_24024,N_24331);
nor U26073 (N_26073,N_24200,N_25198);
nor U26074 (N_26074,N_24576,N_25121);
xnor U26075 (N_26075,N_24487,N_25008);
nor U26076 (N_26076,N_24009,N_24709);
or U26077 (N_26077,N_24058,N_24229);
nand U26078 (N_26078,N_24452,N_24432);
nand U26079 (N_26079,N_24995,N_24749);
xor U26080 (N_26080,N_24788,N_24228);
or U26081 (N_26081,N_24344,N_24640);
or U26082 (N_26082,N_24207,N_24648);
nand U26083 (N_26083,N_25118,N_24786);
and U26084 (N_26084,N_24624,N_25174);
nor U26085 (N_26085,N_24162,N_24569);
and U26086 (N_26086,N_24213,N_24771);
or U26087 (N_26087,N_24210,N_25145);
nand U26088 (N_26088,N_24871,N_24122);
xnor U26089 (N_26089,N_24354,N_25136);
or U26090 (N_26090,N_24954,N_25102);
nand U26091 (N_26091,N_25153,N_24772);
or U26092 (N_26092,N_25022,N_24045);
or U26093 (N_26093,N_24502,N_24961);
nor U26094 (N_26094,N_24609,N_24840);
or U26095 (N_26095,N_25169,N_24279);
nand U26096 (N_26096,N_24395,N_24905);
xnor U26097 (N_26097,N_25119,N_24718);
xor U26098 (N_26098,N_24741,N_24651);
nand U26099 (N_26099,N_24258,N_24175);
or U26100 (N_26100,N_24801,N_24357);
xor U26101 (N_26101,N_24592,N_25031);
or U26102 (N_26102,N_24104,N_24511);
nand U26103 (N_26103,N_24112,N_24383);
nor U26104 (N_26104,N_24922,N_24975);
and U26105 (N_26105,N_24625,N_24896);
and U26106 (N_26106,N_25064,N_24995);
xor U26107 (N_26107,N_24433,N_24723);
and U26108 (N_26108,N_24165,N_25153);
and U26109 (N_26109,N_24848,N_24421);
and U26110 (N_26110,N_25102,N_24782);
and U26111 (N_26111,N_24424,N_24288);
nand U26112 (N_26112,N_24765,N_24802);
nor U26113 (N_26113,N_24524,N_24916);
or U26114 (N_26114,N_24220,N_24261);
nand U26115 (N_26115,N_24811,N_24415);
and U26116 (N_26116,N_24807,N_24373);
nand U26117 (N_26117,N_25068,N_24843);
nand U26118 (N_26118,N_24604,N_24821);
xor U26119 (N_26119,N_24711,N_24622);
or U26120 (N_26120,N_24315,N_24628);
xor U26121 (N_26121,N_25107,N_24231);
and U26122 (N_26122,N_24084,N_24951);
xor U26123 (N_26123,N_25151,N_24141);
nand U26124 (N_26124,N_25052,N_25013);
nand U26125 (N_26125,N_25198,N_24373);
xnor U26126 (N_26126,N_25060,N_24616);
nand U26127 (N_26127,N_24476,N_24641);
and U26128 (N_26128,N_24961,N_25182);
nand U26129 (N_26129,N_24080,N_25027);
and U26130 (N_26130,N_24472,N_24643);
or U26131 (N_26131,N_24179,N_25122);
and U26132 (N_26132,N_24056,N_24983);
xnor U26133 (N_26133,N_24718,N_24946);
and U26134 (N_26134,N_25141,N_24656);
nor U26135 (N_26135,N_24789,N_24207);
xor U26136 (N_26136,N_24043,N_24554);
and U26137 (N_26137,N_24035,N_25128);
and U26138 (N_26138,N_24590,N_24647);
nor U26139 (N_26139,N_24648,N_24267);
or U26140 (N_26140,N_25162,N_25174);
nand U26141 (N_26141,N_24464,N_24454);
nand U26142 (N_26142,N_24785,N_24467);
nor U26143 (N_26143,N_24881,N_25160);
or U26144 (N_26144,N_25073,N_24589);
nor U26145 (N_26145,N_24641,N_24326);
nor U26146 (N_26146,N_24198,N_24687);
nand U26147 (N_26147,N_24696,N_24398);
or U26148 (N_26148,N_24584,N_24423);
nand U26149 (N_26149,N_24971,N_24523);
nand U26150 (N_26150,N_25102,N_24622);
nand U26151 (N_26151,N_24110,N_24604);
and U26152 (N_26152,N_24430,N_25168);
and U26153 (N_26153,N_24437,N_24483);
or U26154 (N_26154,N_24013,N_24781);
or U26155 (N_26155,N_24392,N_25173);
nand U26156 (N_26156,N_24130,N_24702);
and U26157 (N_26157,N_24575,N_24995);
and U26158 (N_26158,N_24467,N_24524);
nand U26159 (N_26159,N_24817,N_24685);
and U26160 (N_26160,N_24392,N_24929);
nand U26161 (N_26161,N_24597,N_24856);
xnor U26162 (N_26162,N_24911,N_24200);
nor U26163 (N_26163,N_24640,N_24523);
and U26164 (N_26164,N_24216,N_25036);
and U26165 (N_26165,N_24578,N_24058);
or U26166 (N_26166,N_24215,N_24349);
xnor U26167 (N_26167,N_24047,N_24257);
or U26168 (N_26168,N_25021,N_24764);
or U26169 (N_26169,N_24825,N_24401);
nand U26170 (N_26170,N_24491,N_24953);
or U26171 (N_26171,N_24728,N_24304);
or U26172 (N_26172,N_24871,N_24079);
nor U26173 (N_26173,N_24596,N_25182);
nand U26174 (N_26174,N_24084,N_24377);
and U26175 (N_26175,N_24092,N_24942);
and U26176 (N_26176,N_24019,N_24213);
or U26177 (N_26177,N_24588,N_24317);
or U26178 (N_26178,N_24018,N_24362);
nor U26179 (N_26179,N_24125,N_24730);
xnor U26180 (N_26180,N_24619,N_24285);
xnor U26181 (N_26181,N_24455,N_24873);
and U26182 (N_26182,N_24581,N_24906);
and U26183 (N_26183,N_25159,N_24960);
and U26184 (N_26184,N_24184,N_24437);
or U26185 (N_26185,N_24069,N_24823);
or U26186 (N_26186,N_24344,N_24795);
nor U26187 (N_26187,N_24654,N_24305);
nand U26188 (N_26188,N_24013,N_24500);
and U26189 (N_26189,N_24826,N_24702);
nor U26190 (N_26190,N_24609,N_24370);
or U26191 (N_26191,N_24824,N_24645);
or U26192 (N_26192,N_24937,N_24046);
nand U26193 (N_26193,N_24683,N_24332);
xnor U26194 (N_26194,N_24726,N_25175);
and U26195 (N_26195,N_25096,N_24884);
or U26196 (N_26196,N_24531,N_24249);
or U26197 (N_26197,N_24015,N_24355);
and U26198 (N_26198,N_24780,N_24758);
or U26199 (N_26199,N_24891,N_25163);
and U26200 (N_26200,N_24205,N_24007);
nor U26201 (N_26201,N_24051,N_24123);
xor U26202 (N_26202,N_25170,N_24506);
nand U26203 (N_26203,N_24126,N_24381);
nand U26204 (N_26204,N_25077,N_25070);
nand U26205 (N_26205,N_25188,N_24750);
xnor U26206 (N_26206,N_24038,N_25013);
xnor U26207 (N_26207,N_24939,N_24968);
nand U26208 (N_26208,N_24561,N_24335);
xor U26209 (N_26209,N_24402,N_24873);
or U26210 (N_26210,N_24539,N_24654);
or U26211 (N_26211,N_24527,N_25137);
or U26212 (N_26212,N_25187,N_24251);
and U26213 (N_26213,N_24312,N_24854);
or U26214 (N_26214,N_24530,N_24625);
nand U26215 (N_26215,N_24633,N_24999);
nor U26216 (N_26216,N_24437,N_24310);
and U26217 (N_26217,N_25046,N_25181);
nor U26218 (N_26218,N_25004,N_24445);
nand U26219 (N_26219,N_24994,N_24204);
xor U26220 (N_26220,N_25048,N_24641);
nor U26221 (N_26221,N_24933,N_24080);
xnor U26222 (N_26222,N_24958,N_25005);
and U26223 (N_26223,N_24790,N_24727);
nand U26224 (N_26224,N_24827,N_24186);
xor U26225 (N_26225,N_24670,N_24040);
and U26226 (N_26226,N_24120,N_24588);
nand U26227 (N_26227,N_24800,N_24711);
xnor U26228 (N_26228,N_24697,N_24533);
or U26229 (N_26229,N_25132,N_24559);
xnor U26230 (N_26230,N_24490,N_24902);
and U26231 (N_26231,N_24675,N_25186);
or U26232 (N_26232,N_24856,N_24118);
nand U26233 (N_26233,N_24159,N_24507);
nor U26234 (N_26234,N_24628,N_24217);
xor U26235 (N_26235,N_24990,N_24884);
xor U26236 (N_26236,N_24610,N_24758);
and U26237 (N_26237,N_24371,N_24146);
and U26238 (N_26238,N_24566,N_24012);
and U26239 (N_26239,N_24755,N_25134);
nor U26240 (N_26240,N_24946,N_24320);
and U26241 (N_26241,N_24526,N_24606);
and U26242 (N_26242,N_24757,N_24991);
or U26243 (N_26243,N_24537,N_25164);
nor U26244 (N_26244,N_24127,N_24392);
xor U26245 (N_26245,N_24763,N_24157);
nor U26246 (N_26246,N_24868,N_24448);
and U26247 (N_26247,N_24198,N_25177);
nand U26248 (N_26248,N_24136,N_24594);
xor U26249 (N_26249,N_24760,N_25166);
nand U26250 (N_26250,N_24176,N_24236);
and U26251 (N_26251,N_25075,N_24334);
or U26252 (N_26252,N_24900,N_24119);
nand U26253 (N_26253,N_24558,N_24388);
or U26254 (N_26254,N_24262,N_24177);
nor U26255 (N_26255,N_24597,N_25034);
xor U26256 (N_26256,N_24330,N_25003);
nand U26257 (N_26257,N_24307,N_24444);
nor U26258 (N_26258,N_24863,N_24564);
nand U26259 (N_26259,N_24630,N_24417);
nor U26260 (N_26260,N_24535,N_24722);
xnor U26261 (N_26261,N_24270,N_25153);
xor U26262 (N_26262,N_25046,N_25089);
or U26263 (N_26263,N_24200,N_24025);
nand U26264 (N_26264,N_24038,N_25017);
or U26265 (N_26265,N_25131,N_25157);
or U26266 (N_26266,N_24457,N_25166);
xnor U26267 (N_26267,N_24425,N_24742);
nand U26268 (N_26268,N_24071,N_24925);
nand U26269 (N_26269,N_24229,N_24275);
nand U26270 (N_26270,N_25043,N_24986);
and U26271 (N_26271,N_24960,N_24934);
and U26272 (N_26272,N_24978,N_24692);
nor U26273 (N_26273,N_24206,N_24211);
and U26274 (N_26274,N_24919,N_24366);
or U26275 (N_26275,N_24185,N_24901);
nor U26276 (N_26276,N_24082,N_25123);
nand U26277 (N_26277,N_24708,N_24259);
nand U26278 (N_26278,N_24417,N_24808);
nand U26279 (N_26279,N_24087,N_24420);
xnor U26280 (N_26280,N_24037,N_24185);
xnor U26281 (N_26281,N_24530,N_24202);
and U26282 (N_26282,N_24124,N_24839);
or U26283 (N_26283,N_25090,N_24158);
nand U26284 (N_26284,N_24145,N_25038);
nor U26285 (N_26285,N_24259,N_24177);
nor U26286 (N_26286,N_24743,N_25196);
nand U26287 (N_26287,N_24468,N_24748);
nor U26288 (N_26288,N_24809,N_24837);
nand U26289 (N_26289,N_24978,N_24718);
and U26290 (N_26290,N_24330,N_24936);
and U26291 (N_26291,N_25130,N_24478);
and U26292 (N_26292,N_24076,N_24599);
and U26293 (N_26293,N_25110,N_25192);
xnor U26294 (N_26294,N_24890,N_24361);
and U26295 (N_26295,N_24518,N_24203);
nor U26296 (N_26296,N_24409,N_24334);
nand U26297 (N_26297,N_24225,N_24296);
nor U26298 (N_26298,N_24907,N_24957);
nor U26299 (N_26299,N_24585,N_24642);
or U26300 (N_26300,N_24193,N_25044);
xnor U26301 (N_26301,N_24922,N_24303);
xor U26302 (N_26302,N_25014,N_24846);
or U26303 (N_26303,N_24321,N_24057);
nand U26304 (N_26304,N_24737,N_24054);
nor U26305 (N_26305,N_24193,N_24482);
xnor U26306 (N_26306,N_25185,N_24475);
or U26307 (N_26307,N_24850,N_24630);
and U26308 (N_26308,N_24624,N_24298);
nor U26309 (N_26309,N_24522,N_24342);
and U26310 (N_26310,N_24781,N_24700);
or U26311 (N_26311,N_24048,N_24396);
nor U26312 (N_26312,N_24313,N_24178);
or U26313 (N_26313,N_24232,N_25100);
or U26314 (N_26314,N_24219,N_24339);
or U26315 (N_26315,N_24449,N_24295);
xor U26316 (N_26316,N_25046,N_24346);
xnor U26317 (N_26317,N_24714,N_24478);
nand U26318 (N_26318,N_24353,N_24098);
or U26319 (N_26319,N_24263,N_24919);
and U26320 (N_26320,N_24951,N_24595);
xor U26321 (N_26321,N_24466,N_24957);
and U26322 (N_26322,N_24530,N_25087);
xor U26323 (N_26323,N_24447,N_24804);
and U26324 (N_26324,N_24662,N_24047);
nand U26325 (N_26325,N_24156,N_24102);
and U26326 (N_26326,N_24560,N_24910);
and U26327 (N_26327,N_24472,N_24225);
and U26328 (N_26328,N_24206,N_24914);
xnor U26329 (N_26329,N_25178,N_24900);
nand U26330 (N_26330,N_24418,N_25069);
nor U26331 (N_26331,N_24696,N_24455);
xnor U26332 (N_26332,N_24881,N_24986);
or U26333 (N_26333,N_24401,N_24657);
nor U26334 (N_26334,N_24326,N_24828);
or U26335 (N_26335,N_24057,N_24886);
and U26336 (N_26336,N_24691,N_24234);
and U26337 (N_26337,N_24396,N_24434);
or U26338 (N_26338,N_24315,N_24231);
or U26339 (N_26339,N_24075,N_25007);
nand U26340 (N_26340,N_24656,N_25082);
or U26341 (N_26341,N_24619,N_24658);
or U26342 (N_26342,N_24247,N_24944);
xor U26343 (N_26343,N_25004,N_24317);
xnor U26344 (N_26344,N_24703,N_24013);
or U26345 (N_26345,N_24147,N_24468);
nor U26346 (N_26346,N_24498,N_24629);
nand U26347 (N_26347,N_25051,N_24314);
and U26348 (N_26348,N_24777,N_24368);
and U26349 (N_26349,N_25165,N_24572);
xnor U26350 (N_26350,N_24371,N_24240);
xnor U26351 (N_26351,N_24065,N_25112);
nor U26352 (N_26352,N_24275,N_24191);
nand U26353 (N_26353,N_25033,N_24267);
nand U26354 (N_26354,N_24003,N_24168);
nor U26355 (N_26355,N_24031,N_25025);
xnor U26356 (N_26356,N_24158,N_24511);
and U26357 (N_26357,N_24006,N_24357);
xor U26358 (N_26358,N_24458,N_24650);
nor U26359 (N_26359,N_24529,N_24287);
nor U26360 (N_26360,N_24903,N_24211);
or U26361 (N_26361,N_24634,N_24761);
nand U26362 (N_26362,N_24704,N_25082);
nor U26363 (N_26363,N_24929,N_24934);
xnor U26364 (N_26364,N_24371,N_24340);
nand U26365 (N_26365,N_24493,N_25105);
and U26366 (N_26366,N_24975,N_24052);
nand U26367 (N_26367,N_24330,N_25058);
nor U26368 (N_26368,N_24779,N_24106);
or U26369 (N_26369,N_24915,N_24733);
or U26370 (N_26370,N_24023,N_24350);
xor U26371 (N_26371,N_24797,N_24661);
and U26372 (N_26372,N_24113,N_24088);
nor U26373 (N_26373,N_24871,N_24738);
xor U26374 (N_26374,N_24742,N_24240);
nand U26375 (N_26375,N_24318,N_24157);
or U26376 (N_26376,N_24711,N_24930);
and U26377 (N_26377,N_24981,N_24966);
nand U26378 (N_26378,N_24080,N_25144);
nor U26379 (N_26379,N_24001,N_24022);
or U26380 (N_26380,N_24083,N_25030);
xnor U26381 (N_26381,N_24836,N_24175);
nor U26382 (N_26382,N_24029,N_24675);
xor U26383 (N_26383,N_24454,N_24256);
xnor U26384 (N_26384,N_24630,N_24681);
xnor U26385 (N_26385,N_24772,N_24457);
nand U26386 (N_26386,N_25078,N_24087);
nand U26387 (N_26387,N_24121,N_24299);
and U26388 (N_26388,N_24325,N_25078);
and U26389 (N_26389,N_24715,N_24342);
xor U26390 (N_26390,N_24344,N_25147);
and U26391 (N_26391,N_24707,N_24370);
xor U26392 (N_26392,N_24166,N_25057);
nand U26393 (N_26393,N_24537,N_24505);
nor U26394 (N_26394,N_24978,N_24629);
nor U26395 (N_26395,N_24936,N_24679);
nand U26396 (N_26396,N_24267,N_24046);
nand U26397 (N_26397,N_24579,N_24808);
and U26398 (N_26398,N_24526,N_24064);
and U26399 (N_26399,N_24163,N_24190);
and U26400 (N_26400,N_26016,N_25218);
nand U26401 (N_26401,N_26273,N_25400);
xnor U26402 (N_26402,N_25326,N_26315);
or U26403 (N_26403,N_25894,N_25712);
or U26404 (N_26404,N_25747,N_26262);
or U26405 (N_26405,N_26151,N_25691);
and U26406 (N_26406,N_25944,N_25336);
or U26407 (N_26407,N_25949,N_25500);
or U26408 (N_26408,N_25236,N_26179);
nor U26409 (N_26409,N_25437,N_26389);
and U26410 (N_26410,N_25463,N_25857);
xor U26411 (N_26411,N_25334,N_25749);
and U26412 (N_26412,N_25958,N_26268);
nand U26413 (N_26413,N_26109,N_26154);
nand U26414 (N_26414,N_26146,N_25621);
nand U26415 (N_26415,N_25455,N_26038);
nand U26416 (N_26416,N_25587,N_26275);
or U26417 (N_26417,N_26283,N_26105);
xor U26418 (N_26418,N_25456,N_26312);
xor U26419 (N_26419,N_25491,N_25699);
nor U26420 (N_26420,N_25531,N_26333);
nand U26421 (N_26421,N_26061,N_26090);
xnor U26422 (N_26422,N_25237,N_25864);
xnor U26423 (N_26423,N_25503,N_25450);
or U26424 (N_26424,N_25506,N_26013);
and U26425 (N_26425,N_25207,N_25243);
and U26426 (N_26426,N_25411,N_26040);
or U26427 (N_26427,N_25302,N_26205);
nor U26428 (N_26428,N_25341,N_25911);
xor U26429 (N_26429,N_25555,N_26354);
and U26430 (N_26430,N_25553,N_25808);
and U26431 (N_26431,N_25282,N_26189);
nor U26432 (N_26432,N_25255,N_25263);
nand U26433 (N_26433,N_25759,N_25375);
nor U26434 (N_26434,N_26102,N_25510);
nand U26435 (N_26435,N_25995,N_25443);
and U26436 (N_26436,N_25863,N_26006);
xnor U26437 (N_26437,N_25420,N_26286);
nand U26438 (N_26438,N_26106,N_25370);
or U26439 (N_26439,N_25946,N_25515);
or U26440 (N_26440,N_25608,N_26089);
and U26441 (N_26441,N_25261,N_26256);
nand U26442 (N_26442,N_25895,N_26091);
or U26443 (N_26443,N_25920,N_26015);
nor U26444 (N_26444,N_25815,N_25671);
xor U26445 (N_26445,N_25265,N_25512);
xor U26446 (N_26446,N_25554,N_26330);
nand U26447 (N_26447,N_25381,N_25602);
nor U26448 (N_26448,N_25366,N_25896);
or U26449 (N_26449,N_25718,N_25980);
nor U26450 (N_26450,N_26281,N_25720);
nor U26451 (N_26451,N_26181,N_26134);
and U26452 (N_26452,N_25917,N_25574);
nor U26453 (N_26453,N_25286,N_25357);
and U26454 (N_26454,N_26382,N_26245);
xnor U26455 (N_26455,N_26055,N_25541);
or U26456 (N_26456,N_26085,N_25490);
and U26457 (N_26457,N_25543,N_26067);
and U26458 (N_26458,N_25790,N_25998);
nor U26459 (N_26459,N_26225,N_25916);
and U26460 (N_26460,N_25414,N_25853);
nor U26461 (N_26461,N_25644,N_25557);
and U26462 (N_26462,N_25881,N_25509);
or U26463 (N_26463,N_25732,N_26374);
xnor U26464 (N_26464,N_25733,N_26168);
nor U26465 (N_26465,N_25914,N_26131);
and U26466 (N_26466,N_26327,N_25385);
or U26467 (N_26467,N_25270,N_26249);
or U26468 (N_26468,N_26296,N_26349);
and U26469 (N_26469,N_25795,N_25383);
nand U26470 (N_26470,N_26182,N_26025);
and U26471 (N_26471,N_25227,N_25902);
nor U26472 (N_26472,N_26053,N_25729);
nor U26473 (N_26473,N_26149,N_26171);
nand U26474 (N_26474,N_25724,N_25208);
and U26475 (N_26475,N_25735,N_25384);
nand U26476 (N_26476,N_26384,N_25498);
nand U26477 (N_26477,N_26282,N_26045);
nor U26478 (N_26478,N_25473,N_26071);
and U26479 (N_26479,N_25992,N_26211);
and U26480 (N_26480,N_26394,N_25812);
xnor U26481 (N_26481,N_25952,N_26231);
nor U26482 (N_26482,N_25344,N_25764);
nand U26483 (N_26483,N_25762,N_26087);
nor U26484 (N_26484,N_25530,N_26056);
xor U26485 (N_26485,N_26012,N_26223);
nor U26486 (N_26486,N_26203,N_25943);
nand U26487 (N_26487,N_25754,N_25360);
or U26488 (N_26488,N_25818,N_25628);
xnor U26489 (N_26489,N_25890,N_25390);
nor U26490 (N_26490,N_25775,N_25313);
xnor U26491 (N_26491,N_26062,N_25717);
or U26492 (N_26492,N_25904,N_26024);
or U26493 (N_26493,N_25690,N_26185);
xnor U26494 (N_26494,N_25471,N_26216);
or U26495 (N_26495,N_26356,N_25327);
and U26496 (N_26496,N_26371,N_25311);
nand U26497 (N_26497,N_25810,N_26079);
xor U26498 (N_26498,N_25955,N_25453);
nor U26499 (N_26499,N_26021,N_25329);
nand U26500 (N_26500,N_26165,N_26169);
xor U26501 (N_26501,N_25993,N_26117);
or U26502 (N_26502,N_25449,N_26298);
nor U26503 (N_26503,N_25589,N_25533);
and U26504 (N_26504,N_25353,N_25367);
or U26505 (N_26505,N_25565,N_25852);
xnor U26506 (N_26506,N_26258,N_25285);
nor U26507 (N_26507,N_25880,N_25447);
xor U26508 (N_26508,N_25734,N_26058);
xor U26509 (N_26509,N_26043,N_25428);
and U26510 (N_26510,N_25746,N_26277);
nand U26511 (N_26511,N_26167,N_25518);
and U26512 (N_26512,N_25758,N_25290);
xnor U26513 (N_26513,N_25647,N_26379);
and U26514 (N_26514,N_26158,N_25232);
or U26515 (N_26515,N_25568,N_25933);
nor U26516 (N_26516,N_25607,N_25984);
or U26517 (N_26517,N_25844,N_26338);
xnor U26518 (N_26518,N_25798,N_26299);
nand U26519 (N_26519,N_26121,N_25297);
nor U26520 (N_26520,N_25600,N_25703);
and U26521 (N_26521,N_25292,N_25362);
or U26522 (N_26522,N_25637,N_25959);
nand U26523 (N_26523,N_25882,N_25953);
and U26524 (N_26524,N_26235,N_26074);
nor U26525 (N_26525,N_25532,N_25440);
or U26526 (N_26526,N_25640,N_25427);
and U26527 (N_26527,N_25348,N_25773);
nor U26528 (N_26528,N_25900,N_25272);
and U26529 (N_26529,N_26057,N_25805);
or U26530 (N_26530,N_25422,N_26322);
xnor U26531 (N_26531,N_25763,N_26019);
nand U26532 (N_26532,N_25672,N_25639);
or U26533 (N_26533,N_25927,N_25337);
xor U26534 (N_26534,N_25251,N_26314);
nand U26535 (N_26535,N_25583,N_25433);
xor U26536 (N_26536,N_25289,N_26307);
or U26537 (N_26537,N_25250,N_25737);
nand U26538 (N_26538,N_25664,N_25591);
or U26539 (N_26539,N_25338,N_26030);
nor U26540 (N_26540,N_25392,N_25968);
and U26541 (N_26541,N_25750,N_26092);
or U26542 (N_26542,N_25741,N_25238);
xnor U26543 (N_26543,N_26157,N_25310);
or U26544 (N_26544,N_25402,N_26359);
or U26545 (N_26545,N_26065,N_26125);
nor U26546 (N_26546,N_25909,N_25800);
xor U26547 (N_26547,N_25442,N_25839);
nor U26548 (N_26548,N_25331,N_25934);
nor U26549 (N_26549,N_26034,N_25861);
nor U26550 (N_26550,N_25889,N_25778);
xor U26551 (N_26551,N_25830,N_25472);
xnor U26552 (N_26552,N_25981,N_25947);
and U26553 (N_26553,N_25298,N_26214);
nor U26554 (N_26554,N_26098,N_26237);
nor U26555 (N_26555,N_26114,N_25316);
xnor U26556 (N_26556,N_26335,N_25504);
nor U26557 (N_26557,N_25675,N_26292);
xnor U26558 (N_26558,N_25211,N_26357);
and U26559 (N_26559,N_25303,N_25976);
and U26560 (N_26560,N_26103,N_25979);
or U26561 (N_26561,N_25252,N_26267);
nor U26562 (N_26562,N_25626,N_25835);
or U26563 (N_26563,N_26007,N_26200);
or U26564 (N_26564,N_25652,N_26177);
or U26565 (N_26565,N_25828,N_26378);
nand U26566 (N_26566,N_26112,N_26093);
xor U26567 (N_26567,N_26122,N_25714);
and U26568 (N_26568,N_25833,N_25431);
and U26569 (N_26569,N_25249,N_25556);
xor U26570 (N_26570,N_25802,N_25674);
nand U26571 (N_26571,N_26035,N_26377);
nand U26572 (N_26572,N_26070,N_25725);
and U26573 (N_26573,N_26077,N_26289);
nand U26574 (N_26574,N_25831,N_25209);
or U26575 (N_26575,N_25539,N_25971);
xnor U26576 (N_26576,N_25845,N_25215);
or U26577 (N_26577,N_26241,N_25730);
and U26578 (N_26578,N_25693,N_26175);
and U26579 (N_26579,N_26138,N_26368);
or U26580 (N_26580,N_25566,N_25941);
xnor U26581 (N_26581,N_26159,N_25776);
nor U26582 (N_26582,N_25304,N_25342);
or U26583 (N_26583,N_26000,N_26284);
nor U26584 (N_26584,N_25448,N_26392);
or U26585 (N_26585,N_26005,N_26041);
nand U26586 (N_26586,N_25657,N_25634);
nand U26587 (N_26587,N_25906,N_26320);
nor U26588 (N_26588,N_26161,N_25784);
nor U26589 (N_26589,N_25929,N_25570);
xnor U26590 (N_26590,N_25796,N_25722);
nand U26591 (N_26591,N_25579,N_25616);
nand U26592 (N_26592,N_25507,N_25723);
nor U26593 (N_26593,N_26329,N_25409);
or U26594 (N_26594,N_25423,N_25288);
nor U26595 (N_26595,N_25697,N_26328);
xor U26596 (N_26596,N_25965,N_25642);
xor U26597 (N_26597,N_25840,N_25323);
xnor U26598 (N_26598,N_25974,N_25740);
xnor U26599 (N_26599,N_25494,N_25225);
nor U26600 (N_26600,N_25314,N_25551);
nor U26601 (N_26601,N_25226,N_25903);
xor U26602 (N_26602,N_25445,N_26325);
or U26603 (N_26603,N_26300,N_25223);
nor U26604 (N_26604,N_25614,N_25982);
xnor U26605 (N_26605,N_25465,N_25562);
xor U26606 (N_26606,N_25351,N_26039);
nand U26607 (N_26607,N_25827,N_26269);
and U26608 (N_26608,N_26010,N_25312);
or U26609 (N_26609,N_25849,N_25649);
nand U26610 (N_26610,N_25239,N_25511);
nand U26611 (N_26611,N_26381,N_25470);
or U26612 (N_26612,N_25493,N_25783);
nand U26613 (N_26613,N_25676,N_26048);
nor U26614 (N_26614,N_25659,N_25240);
or U26615 (N_26615,N_25374,N_26340);
or U26616 (N_26616,N_25726,N_25985);
xor U26617 (N_26617,N_25997,N_26014);
and U26618 (N_26618,N_25508,N_25571);
and U26619 (N_26619,N_25829,N_25418);
or U26620 (N_26620,N_25680,N_26032);
and U26621 (N_26621,N_26324,N_26022);
xor U26622 (N_26622,N_25459,N_25373);
nand U26623 (N_26623,N_25434,N_25273);
nor U26624 (N_26624,N_25281,N_25970);
or U26625 (N_26625,N_26336,N_25537);
or U26626 (N_26626,N_26366,N_25388);
or U26627 (N_26627,N_25661,N_25843);
and U26628 (N_26628,N_26060,N_25613);
nor U26629 (N_26629,N_25766,N_25820);
nand U26630 (N_26630,N_26194,N_25436);
nand U26631 (N_26631,N_25987,N_26209);
or U26632 (N_26632,N_26051,N_26029);
nand U26633 (N_26633,N_25709,N_26050);
and U26634 (N_26634,N_25645,N_26229);
xor U26635 (N_26635,N_25293,N_26355);
or U26636 (N_26636,N_25467,N_25529);
nor U26637 (N_26637,N_26127,N_25309);
nand U26638 (N_26638,N_25951,N_26266);
or U26639 (N_26639,N_25899,N_25922);
or U26640 (N_26640,N_25578,N_25935);
and U26641 (N_26641,N_25253,N_25678);
nand U26642 (N_26642,N_25387,N_26193);
xnor U26643 (N_26643,N_26084,N_26135);
and U26644 (N_26644,N_25221,N_25689);
xnor U26645 (N_26645,N_26238,N_25969);
and U26646 (N_26646,N_26027,N_25241);
or U26647 (N_26647,N_25753,N_25478);
nor U26648 (N_26648,N_25660,N_26246);
xor U26649 (N_26649,N_26352,N_25668);
nand U26650 (N_26650,N_25203,N_26236);
xnor U26651 (N_26651,N_25874,N_25405);
nand U26652 (N_26652,N_25622,N_25322);
nor U26653 (N_26653,N_26118,N_25266);
and U26654 (N_26654,N_25960,N_25558);
nor U26655 (N_26655,N_25742,N_26173);
nor U26656 (N_26656,N_26222,N_26001);
xnor U26657 (N_26657,N_26063,N_25915);
nand U26658 (N_26658,N_26270,N_25938);
xor U26659 (N_26659,N_26153,N_26008);
xor U26660 (N_26660,N_25877,N_25786);
or U26661 (N_26661,N_26124,N_26028);
nor U26662 (N_26662,N_25777,N_26257);
xor U26663 (N_26663,N_25205,N_26278);
and U26664 (N_26664,N_26059,N_26380);
nand U26665 (N_26665,N_25686,N_25569);
or U26666 (N_26666,N_25536,N_25325);
or U26667 (N_26667,N_26309,N_25978);
and U26668 (N_26668,N_25495,N_26248);
xor U26669 (N_26669,N_25561,N_25332);
or U26670 (N_26670,N_25278,N_25564);
or U26671 (N_26671,N_26254,N_25983);
xnor U26672 (N_26672,N_25658,N_25576);
nor U26673 (N_26673,N_26166,N_26215);
or U26674 (N_26674,N_25785,N_25458);
nor U26675 (N_26675,N_25867,N_25596);
or U26676 (N_26676,N_25279,N_25716);
nor U26677 (N_26677,N_26397,N_25771);
nor U26678 (N_26678,N_25986,N_25772);
nand U26679 (N_26679,N_25931,N_25866);
nand U26680 (N_26680,N_26361,N_25841);
nor U26681 (N_26681,N_25228,N_25248);
nor U26682 (N_26682,N_25345,N_25213);
and U26683 (N_26683,N_25299,N_25319);
or U26684 (N_26684,N_26064,N_26375);
and U26685 (N_26685,N_25277,N_26126);
xor U26686 (N_26686,N_25363,N_25468);
xnor U26687 (N_26687,N_25954,N_25807);
and U26688 (N_26688,N_26319,N_25797);
nand U26689 (N_26689,N_25372,N_25590);
xor U26690 (N_26690,N_26207,N_25623);
xnor U26691 (N_26691,N_25328,N_26210);
xor U26692 (N_26692,N_25646,N_25609);
and U26693 (N_26693,N_26178,N_26142);
nand U26694 (N_26694,N_26233,N_25519);
nand U26695 (N_26695,N_25575,N_25430);
nor U26696 (N_26696,N_25296,N_25701);
and U26697 (N_26697,N_25999,N_26387);
and U26698 (N_26698,N_26206,N_25306);
and U26699 (N_26699,N_26107,N_25694);
or U26700 (N_26700,N_26137,N_25760);
and U26701 (N_26701,N_25582,N_25665);
xor U26702 (N_26702,N_25315,N_26049);
and U26703 (N_26703,N_25869,N_25897);
and U26704 (N_26704,N_25271,N_26306);
or U26705 (N_26705,N_25625,N_25663);
and U26706 (N_26706,N_25408,N_25403);
nor U26707 (N_26707,N_25682,N_25876);
and U26708 (N_26708,N_26372,N_25966);
and U26709 (N_26709,N_26195,N_25435);
xnor U26710 (N_26710,N_26099,N_25755);
and U26711 (N_26711,N_25545,N_25603);
nand U26712 (N_26712,N_25346,N_25688);
and U26713 (N_26713,N_25521,N_26075);
nor U26714 (N_26714,N_25848,N_25872);
and U26715 (N_26715,N_26297,N_26370);
nor U26716 (N_26716,N_26343,N_26365);
nand U26717 (N_26717,N_25748,N_25605);
and U26718 (N_26718,N_25768,N_26160);
nor U26719 (N_26719,N_26190,N_25548);
nor U26720 (N_26720,N_25617,N_25485);
or U26721 (N_26721,N_25563,N_25260);
xnor U26722 (N_26722,N_26148,N_25779);
xnor U26723 (N_26723,N_25862,N_26046);
nor U26724 (N_26724,N_26294,N_25301);
nand U26725 (N_26725,N_26100,N_26310);
nor U26726 (N_26726,N_26304,N_25814);
nand U26727 (N_26727,N_26009,N_26110);
nor U26728 (N_26728,N_25695,N_25247);
or U26729 (N_26729,N_25884,N_25859);
and U26730 (N_26730,N_26183,N_26066);
nor U26731 (N_26731,N_26260,N_26252);
xor U26732 (N_26732,N_26052,N_26076);
nand U26733 (N_26733,N_25318,N_25480);
and U26734 (N_26734,N_26080,N_26265);
nor U26735 (N_26735,N_25234,N_25534);
or U26736 (N_26736,N_26255,N_25751);
nor U26737 (N_26737,N_25501,N_25242);
nand U26738 (N_26738,N_25923,N_25404);
nor U26739 (N_26739,N_25956,N_26191);
xor U26740 (N_26740,N_25333,N_26120);
xor U26741 (N_26741,N_26342,N_25816);
nand U26742 (N_26742,N_25624,N_26344);
nor U26743 (N_26743,N_25454,N_25441);
xor U26744 (N_26744,N_25886,N_25438);
nor U26745 (N_26745,N_26155,N_25977);
nand U26746 (N_26746,N_26323,N_25481);
nor U26747 (N_26747,N_26228,N_25888);
or U26748 (N_26748,N_26002,N_25854);
nor U26749 (N_26749,N_25809,N_26170);
xor U26750 (N_26750,N_25873,N_26351);
and U26751 (N_26751,N_25222,N_25417);
or U26752 (N_26752,N_25425,N_26263);
nand U26753 (N_26753,N_26128,N_25502);
nor U26754 (N_26754,N_25516,N_25499);
xnor U26755 (N_26755,N_25567,N_25817);
and U26756 (N_26756,N_26054,N_25486);
and U26757 (N_26757,N_25662,N_26253);
and U26758 (N_26758,N_25908,N_25280);
or U26759 (N_26759,N_25517,N_26004);
and U26760 (N_26760,N_25856,N_25648);
or U26761 (N_26761,N_26201,N_25618);
xor U26762 (N_26762,N_25950,N_25787);
or U26763 (N_26763,N_25926,N_25451);
xor U26764 (N_26764,N_26243,N_25257);
nor U26765 (N_26765,N_26271,N_26391);
and U26766 (N_26766,N_25972,N_26083);
or U26767 (N_26767,N_26348,N_25898);
nand U26768 (N_26768,N_25415,N_25728);
or U26769 (N_26769,N_25667,N_25948);
or U26770 (N_26770,N_25632,N_25653);
and U26771 (N_26771,N_25719,N_25887);
and U26772 (N_26772,N_26111,N_26184);
and U26773 (N_26773,N_26279,N_25460);
nor U26774 (N_26774,N_25397,N_26156);
nor U26775 (N_26775,N_25819,N_25756);
nor U26776 (N_26776,N_25782,N_25837);
or U26777 (N_26777,N_26388,N_26383);
nand U26778 (N_26778,N_26398,N_26217);
or U26779 (N_26779,N_25713,N_25924);
and U26780 (N_26780,N_26082,N_25401);
nand U26781 (N_26781,N_25604,N_25484);
nor U26782 (N_26782,N_25912,N_25369);
xor U26783 (N_26783,N_25330,N_26318);
and U26784 (N_26784,N_25487,N_26303);
or U26785 (N_26785,N_25838,N_25631);
or U26786 (N_26786,N_26023,N_25520);
nand U26787 (N_26787,N_26287,N_26140);
nand U26788 (N_26788,N_25633,N_25523);
and U26789 (N_26789,N_25368,N_25842);
and U26790 (N_26790,N_25540,N_25457);
xor U26791 (N_26791,N_26290,N_25291);
nand U26792 (N_26792,N_25254,N_25704);
or U26793 (N_26793,N_25921,N_26176);
nor U26794 (N_26794,N_26003,N_25708);
and U26795 (N_26795,N_26162,N_25581);
or U26796 (N_26796,N_25394,N_25464);
xor U26797 (N_26797,N_25489,N_25352);
nand U26798 (N_26798,N_25477,N_25514);
nand U26799 (N_26799,N_26221,N_25721);
nor U26800 (N_26800,N_25823,N_25643);
or U26801 (N_26801,N_25988,N_25585);
xnor U26802 (N_26802,N_25560,N_25586);
or U26803 (N_26803,N_25870,N_25594);
nor U26804 (N_26804,N_26069,N_26086);
nand U26805 (N_26805,N_25738,N_25426);
or U26806 (N_26806,N_25201,N_26044);
nand U26807 (N_26807,N_26373,N_25547);
nand U26808 (N_26808,N_25317,N_25365);
or U26809 (N_26809,N_26199,N_25630);
and U26810 (N_26810,N_26152,N_25656);
nand U26811 (N_26811,N_25865,N_25268);
nand U26812 (N_26812,N_26313,N_25542);
nand U26813 (N_26813,N_25940,N_25910);
nor U26814 (N_26814,N_26396,N_26172);
and U26815 (N_26815,N_26180,N_26244);
xnor U26816 (N_26816,N_26017,N_25216);
nor U26817 (N_26817,N_26302,N_25918);
nor U26818 (N_26818,N_25466,N_25769);
xnor U26819 (N_26819,N_25687,N_25580);
and U26820 (N_26820,N_26399,N_25421);
xnor U26821 (N_26821,N_25527,N_25552);
or U26822 (N_26822,N_25380,N_25789);
xor U26823 (N_26823,N_26393,N_25476);
xor U26824 (N_26824,N_26317,N_26358);
nand U26825 (N_26825,N_25524,N_25343);
nand U26826 (N_26826,N_25892,N_25361);
xnor U26827 (N_26827,N_26291,N_25599);
and U26828 (N_26828,N_25217,N_26251);
and U26829 (N_26829,N_26141,N_25655);
xnor U26830 (N_26830,N_25505,N_25711);
nor U26831 (N_26831,N_25359,N_26326);
nor U26832 (N_26832,N_25919,N_25761);
nand U26833 (N_26833,N_25780,N_25654);
nor U26834 (N_26834,N_25707,N_25350);
nand U26835 (N_26835,N_26295,N_26031);
nand U26836 (N_26836,N_25528,N_25413);
xor U26837 (N_26837,N_26363,N_25419);
nor U26838 (N_26838,N_26196,N_25396);
nor U26839 (N_26839,N_25597,N_26250);
and U26840 (N_26840,N_26037,N_25496);
nand U26841 (N_26841,N_25650,N_25942);
and U26842 (N_26842,N_25803,N_25407);
xor U26843 (N_26843,N_26042,N_25305);
nand U26844 (N_26844,N_25791,N_25669);
and U26845 (N_26845,N_25535,N_25627);
and U26846 (N_26846,N_26345,N_26280);
nand U26847 (N_26847,N_25378,N_25846);
nor U26848 (N_26848,N_25355,N_26192);
nor U26849 (N_26849,N_25767,N_26337);
xor U26850 (N_26850,N_25264,N_26367);
or U26851 (N_26851,N_25300,N_25598);
xnor U26852 (N_26852,N_25788,N_25757);
xor U26853 (N_26853,N_25684,N_25224);
or U26854 (N_26854,N_25398,N_26198);
and U26855 (N_26855,N_25612,N_26316);
nand U26856 (N_26856,N_25479,N_26139);
nand U26857 (N_26857,N_25619,N_25439);
nor U26858 (N_26858,N_26311,N_26033);
xnor U26859 (N_26859,N_25214,N_26386);
nor U26860 (N_26860,N_26218,N_25936);
and U26861 (N_26861,N_25245,N_25573);
and U26862 (N_26862,N_25860,N_25967);
or U26863 (N_26863,N_26197,N_25677);
or U26864 (N_26864,N_25276,N_26108);
nand U26865 (N_26865,N_25259,N_26219);
nand U26866 (N_26866,N_25611,N_26187);
nand U26867 (N_26867,N_25356,N_25577);
xor U26868 (N_26868,N_25432,N_26230);
xor U26869 (N_26869,N_25868,N_25399);
nor U26870 (N_26870,N_25731,N_26259);
or U26871 (N_26871,N_26020,N_26026);
or U26872 (N_26872,N_25962,N_25262);
xnor U26873 (N_26873,N_26129,N_25593);
xnor U26874 (N_26874,N_25416,N_26301);
xnor U26875 (N_26875,N_26147,N_25636);
nand U26876 (N_26876,N_26261,N_26208);
nor U26877 (N_26877,N_26224,N_26308);
or U26878 (N_26878,N_25386,N_25744);
nand U26879 (N_26879,N_25584,N_25444);
nor U26880 (N_26880,N_25269,N_25932);
and U26881 (N_26881,N_26390,N_25233);
and U26882 (N_26882,N_25811,N_25620);
nor U26883 (N_26883,N_26240,N_25801);
nand U26884 (N_26884,N_25606,N_26285);
nor U26885 (N_26885,N_26341,N_26186);
xor U26886 (N_26886,N_26104,N_26047);
xor U26887 (N_26887,N_25821,N_26220);
nand U26888 (N_26888,N_25231,N_25412);
nor U26889 (N_26889,N_25204,N_25850);
xnor U26890 (N_26890,N_26234,N_25961);
nor U26891 (N_26891,N_26346,N_25549);
nor U26892 (N_26892,N_25794,N_26094);
and U26893 (N_26893,N_25666,N_25715);
and U26894 (N_26894,N_25964,N_25893);
or U26895 (N_26895,N_25937,N_25220);
nor U26896 (N_26896,N_25851,N_25267);
or U26897 (N_26897,N_25641,N_25804);
and U26898 (N_26898,N_25939,N_25358);
or U26899 (N_26899,N_25752,N_25525);
and U26900 (N_26900,N_25610,N_25700);
nor U26901 (N_26901,N_25354,N_26364);
nor U26902 (N_26902,N_25410,N_25364);
xor U26903 (N_26903,N_25376,N_25526);
nand U26904 (N_26904,N_26095,N_25483);
or U26905 (N_26905,N_25615,N_25320);
or U26906 (N_26906,N_25258,N_25321);
xor U26907 (N_26907,N_26144,N_25670);
xor U26908 (N_26908,N_25371,N_25774);
and U26909 (N_26909,N_25875,N_26339);
xor U26910 (N_26910,N_25274,N_25544);
nand U26911 (N_26911,N_26321,N_25871);
nand U26912 (N_26912,N_26332,N_26202);
xnor U26913 (N_26913,N_25475,N_25878);
or U26914 (N_26914,N_25806,N_26101);
and U26915 (N_26915,N_26232,N_25692);
xnor U26916 (N_26916,N_25736,N_26212);
nor U26917 (N_26917,N_25497,N_26395);
nand U26918 (N_26918,N_25284,N_26143);
nand U26919 (N_26919,N_25825,N_25382);
xor U26920 (N_26920,N_25474,N_26078);
and U26921 (N_26921,N_26119,N_25488);
or U26922 (N_26922,N_26242,N_25424);
and U26923 (N_26923,N_26204,N_26164);
nor U26924 (N_26924,N_26239,N_25990);
and U26925 (N_26925,N_26130,N_26088);
nand U26926 (N_26926,N_25377,N_25592);
xnor U26927 (N_26927,N_25492,N_25229);
nor U26928 (N_26928,N_25513,N_25957);
nand U26929 (N_26929,N_26097,N_26288);
xnor U26930 (N_26930,N_26385,N_25308);
nand U26931 (N_26931,N_26362,N_25901);
nand U26932 (N_26932,N_25781,N_25406);
xnor U26933 (N_26933,N_25696,N_25246);
nor U26934 (N_26934,N_25685,N_25393);
xnor U26935 (N_26935,N_25989,N_26227);
or U26936 (N_26936,N_25834,N_25883);
xnor U26937 (N_26937,N_26073,N_25847);
and U26938 (N_26938,N_25452,N_25638);
xnor U26939 (N_26939,N_26145,N_25244);
nand U26940 (N_26940,N_25679,N_25347);
or U26941 (N_26941,N_25210,N_25651);
xor U26942 (N_26942,N_26274,N_25212);
or U26943 (N_26943,N_25905,N_25891);
nand U26944 (N_26944,N_26136,N_25283);
and U26945 (N_26945,N_25832,N_25996);
or U26946 (N_26946,N_25702,N_25461);
xor U26947 (N_26947,N_25287,N_26174);
xnor U26948 (N_26948,N_25673,N_25885);
xor U26949 (N_26949,N_26116,N_25930);
or U26950 (N_26950,N_25522,N_25538);
nor U26951 (N_26951,N_25928,N_25855);
nor U26952 (N_26952,N_25446,N_26350);
nor U26953 (N_26953,N_25339,N_26018);
nor U26954 (N_26954,N_25705,N_25765);
nor U26955 (N_26955,N_25770,N_25635);
and U26956 (N_26956,N_26226,N_26334);
or U26957 (N_26957,N_25739,N_25743);
xor U26958 (N_26958,N_25683,N_25206);
xnor U26959 (N_26959,N_26188,N_25588);
and U26960 (N_26960,N_26331,N_25975);
nand U26961 (N_26961,N_25991,N_25295);
or U26962 (N_26962,N_26096,N_25813);
nand U26963 (N_26963,N_26133,N_26376);
and U26964 (N_26964,N_26115,N_25601);
nor U26965 (N_26965,N_25429,N_26072);
xor U26966 (N_26966,N_25793,N_25202);
or U26967 (N_26967,N_26305,N_25913);
xor U26968 (N_26968,N_25349,N_26150);
nand U26969 (N_26969,N_26011,N_26132);
nor U26970 (N_26970,N_25858,N_25826);
nand U26971 (N_26971,N_25595,N_26276);
and U26972 (N_26972,N_25230,N_25698);
xnor U26973 (N_26973,N_25324,N_26123);
or U26974 (N_26974,N_25792,N_25706);
nor U26975 (N_26975,N_25307,N_25710);
or U26976 (N_26976,N_26353,N_26272);
xor U26977 (N_26977,N_25294,N_25379);
nor U26978 (N_26978,N_25925,N_26163);
nand U26979 (N_26979,N_25335,N_26247);
nand U26980 (N_26980,N_25945,N_25462);
xnor U26981 (N_26981,N_25629,N_26113);
or U26982 (N_26982,N_25559,N_26293);
and U26983 (N_26983,N_26264,N_25550);
and U26984 (N_26984,N_25745,N_26369);
nand U26985 (N_26985,N_25200,N_25389);
and U26986 (N_26986,N_25799,N_25907);
xor U26987 (N_26987,N_25395,N_26347);
and U26988 (N_26988,N_26068,N_25482);
and U26989 (N_26989,N_25469,N_25391);
nand U26990 (N_26990,N_25824,N_26213);
nor U26991 (N_26991,N_26036,N_25256);
or U26992 (N_26992,N_25727,N_25879);
nor U26993 (N_26993,N_25275,N_25219);
or U26994 (N_26994,N_25340,N_25836);
and U26995 (N_26995,N_25546,N_25973);
nand U26996 (N_26996,N_25572,N_25822);
and U26997 (N_26997,N_25963,N_26081);
nor U26998 (N_26998,N_25994,N_25681);
and U26999 (N_26999,N_25235,N_26360);
or U27000 (N_27000,N_25491,N_25798);
and U27001 (N_27001,N_25912,N_25476);
or U27002 (N_27002,N_25808,N_25300);
nand U27003 (N_27003,N_26274,N_25787);
nor U27004 (N_27004,N_25698,N_26230);
nand U27005 (N_27005,N_25912,N_25764);
nor U27006 (N_27006,N_25394,N_25606);
and U27007 (N_27007,N_25224,N_26056);
or U27008 (N_27008,N_25981,N_25979);
nand U27009 (N_27009,N_25607,N_25788);
and U27010 (N_27010,N_26113,N_26315);
nand U27011 (N_27011,N_25905,N_25973);
xnor U27012 (N_27012,N_26214,N_25814);
and U27013 (N_27013,N_25938,N_25325);
nor U27014 (N_27014,N_25645,N_25943);
and U27015 (N_27015,N_25851,N_25817);
or U27016 (N_27016,N_25865,N_25901);
xnor U27017 (N_27017,N_26080,N_25504);
and U27018 (N_27018,N_26306,N_26103);
nand U27019 (N_27019,N_25895,N_26020);
nor U27020 (N_27020,N_25560,N_25626);
and U27021 (N_27021,N_25252,N_25749);
or U27022 (N_27022,N_26306,N_26059);
nor U27023 (N_27023,N_25265,N_25580);
and U27024 (N_27024,N_26262,N_25261);
xor U27025 (N_27025,N_25896,N_25395);
and U27026 (N_27026,N_25442,N_25264);
and U27027 (N_27027,N_25593,N_25445);
xor U27028 (N_27028,N_25714,N_25454);
xor U27029 (N_27029,N_25687,N_26076);
nor U27030 (N_27030,N_25592,N_25863);
xor U27031 (N_27031,N_25720,N_25645);
xnor U27032 (N_27032,N_26253,N_25221);
xnor U27033 (N_27033,N_26200,N_25819);
nand U27034 (N_27034,N_25774,N_26346);
nor U27035 (N_27035,N_25759,N_26316);
nor U27036 (N_27036,N_25751,N_25210);
or U27037 (N_27037,N_25668,N_25917);
xnor U27038 (N_27038,N_25739,N_25876);
and U27039 (N_27039,N_26241,N_26380);
or U27040 (N_27040,N_25483,N_25893);
and U27041 (N_27041,N_26183,N_25278);
and U27042 (N_27042,N_25687,N_25869);
and U27043 (N_27043,N_25562,N_25301);
or U27044 (N_27044,N_25759,N_25641);
nand U27045 (N_27045,N_25678,N_25852);
nor U27046 (N_27046,N_26395,N_25451);
xnor U27047 (N_27047,N_25352,N_25264);
or U27048 (N_27048,N_25613,N_25585);
nor U27049 (N_27049,N_26171,N_25743);
nand U27050 (N_27050,N_26344,N_25569);
nand U27051 (N_27051,N_25215,N_25670);
nand U27052 (N_27052,N_25826,N_25282);
nand U27053 (N_27053,N_26146,N_26133);
or U27054 (N_27054,N_25714,N_25323);
and U27055 (N_27055,N_25994,N_25890);
xor U27056 (N_27056,N_26094,N_25634);
nor U27057 (N_27057,N_25930,N_25988);
xor U27058 (N_27058,N_26241,N_25605);
and U27059 (N_27059,N_26068,N_25695);
nor U27060 (N_27060,N_25363,N_26073);
xor U27061 (N_27061,N_25957,N_25207);
nor U27062 (N_27062,N_25220,N_25284);
and U27063 (N_27063,N_25418,N_25959);
nand U27064 (N_27064,N_26073,N_26296);
and U27065 (N_27065,N_25894,N_25984);
nand U27066 (N_27066,N_25779,N_25566);
and U27067 (N_27067,N_26337,N_26136);
nor U27068 (N_27068,N_25911,N_25406);
and U27069 (N_27069,N_25554,N_25918);
xnor U27070 (N_27070,N_26397,N_25502);
xnor U27071 (N_27071,N_25366,N_25704);
xnor U27072 (N_27072,N_26178,N_26113);
or U27073 (N_27073,N_26118,N_25750);
and U27074 (N_27074,N_25273,N_25801);
or U27075 (N_27075,N_26097,N_26340);
nor U27076 (N_27076,N_25339,N_26258);
nor U27077 (N_27077,N_25666,N_26345);
nor U27078 (N_27078,N_26136,N_25267);
nor U27079 (N_27079,N_25990,N_25761);
nor U27080 (N_27080,N_25207,N_25336);
or U27081 (N_27081,N_25427,N_25272);
or U27082 (N_27082,N_25217,N_26145);
xnor U27083 (N_27083,N_25573,N_26311);
nor U27084 (N_27084,N_26071,N_26358);
or U27085 (N_27085,N_25240,N_25578);
and U27086 (N_27086,N_26271,N_26315);
and U27087 (N_27087,N_25351,N_25288);
nand U27088 (N_27088,N_26370,N_25784);
nor U27089 (N_27089,N_26266,N_25656);
and U27090 (N_27090,N_25305,N_26073);
xnor U27091 (N_27091,N_26299,N_25881);
nor U27092 (N_27092,N_26108,N_25743);
xor U27093 (N_27093,N_25785,N_25839);
xnor U27094 (N_27094,N_26338,N_25949);
nand U27095 (N_27095,N_25315,N_25861);
nor U27096 (N_27096,N_25699,N_25724);
nand U27097 (N_27097,N_25439,N_25974);
or U27098 (N_27098,N_25458,N_26086);
nand U27099 (N_27099,N_25413,N_26353);
xnor U27100 (N_27100,N_25340,N_25578);
or U27101 (N_27101,N_25429,N_25944);
nor U27102 (N_27102,N_25756,N_25369);
xor U27103 (N_27103,N_25234,N_26042);
xnor U27104 (N_27104,N_25635,N_25489);
or U27105 (N_27105,N_25644,N_26184);
nand U27106 (N_27106,N_25733,N_25207);
and U27107 (N_27107,N_26162,N_26181);
xnor U27108 (N_27108,N_26075,N_25709);
nand U27109 (N_27109,N_25270,N_25551);
nand U27110 (N_27110,N_25421,N_25474);
nor U27111 (N_27111,N_25966,N_26316);
nor U27112 (N_27112,N_25349,N_25415);
xor U27113 (N_27113,N_26399,N_25308);
nor U27114 (N_27114,N_26172,N_26077);
xor U27115 (N_27115,N_25877,N_25792);
nor U27116 (N_27116,N_25650,N_26216);
xor U27117 (N_27117,N_26394,N_25739);
nor U27118 (N_27118,N_25771,N_26071);
and U27119 (N_27119,N_26108,N_25333);
or U27120 (N_27120,N_26013,N_25765);
and U27121 (N_27121,N_25977,N_26219);
nor U27122 (N_27122,N_25363,N_26201);
nor U27123 (N_27123,N_25208,N_25784);
and U27124 (N_27124,N_25931,N_25948);
nand U27125 (N_27125,N_25606,N_26100);
nor U27126 (N_27126,N_25822,N_26236);
nand U27127 (N_27127,N_25686,N_25824);
nor U27128 (N_27128,N_25965,N_25422);
nor U27129 (N_27129,N_25786,N_26327);
nand U27130 (N_27130,N_26155,N_25215);
or U27131 (N_27131,N_26023,N_26389);
and U27132 (N_27132,N_26351,N_26211);
nand U27133 (N_27133,N_25762,N_25639);
and U27134 (N_27134,N_25305,N_25451);
and U27135 (N_27135,N_25352,N_25388);
nand U27136 (N_27136,N_26301,N_26069);
or U27137 (N_27137,N_26209,N_25579);
or U27138 (N_27138,N_25276,N_25660);
nor U27139 (N_27139,N_25909,N_25826);
nand U27140 (N_27140,N_25474,N_25212);
xor U27141 (N_27141,N_25877,N_26063);
and U27142 (N_27142,N_26304,N_25712);
xnor U27143 (N_27143,N_26223,N_25808);
nand U27144 (N_27144,N_25839,N_26111);
nand U27145 (N_27145,N_26348,N_26274);
nor U27146 (N_27146,N_25900,N_25495);
xor U27147 (N_27147,N_25708,N_26242);
or U27148 (N_27148,N_25894,N_25870);
nand U27149 (N_27149,N_26267,N_25477);
and U27150 (N_27150,N_25723,N_25484);
nor U27151 (N_27151,N_26397,N_25756);
or U27152 (N_27152,N_25908,N_25318);
and U27153 (N_27153,N_26109,N_25961);
nand U27154 (N_27154,N_25665,N_25532);
nand U27155 (N_27155,N_25610,N_25993);
nand U27156 (N_27156,N_25695,N_25383);
xnor U27157 (N_27157,N_25694,N_25836);
or U27158 (N_27158,N_25587,N_25236);
nor U27159 (N_27159,N_25414,N_25692);
or U27160 (N_27160,N_26028,N_26062);
nor U27161 (N_27161,N_26031,N_25316);
xor U27162 (N_27162,N_26141,N_25639);
and U27163 (N_27163,N_26285,N_25477);
or U27164 (N_27164,N_25714,N_26071);
or U27165 (N_27165,N_25518,N_25364);
xor U27166 (N_27166,N_25728,N_25490);
nor U27167 (N_27167,N_26390,N_25205);
nor U27168 (N_27168,N_25272,N_26124);
or U27169 (N_27169,N_25772,N_25876);
or U27170 (N_27170,N_25242,N_26140);
xor U27171 (N_27171,N_25370,N_25536);
nand U27172 (N_27172,N_26176,N_25446);
nand U27173 (N_27173,N_26000,N_25542);
and U27174 (N_27174,N_26072,N_25441);
or U27175 (N_27175,N_25717,N_25654);
and U27176 (N_27176,N_25951,N_25573);
nand U27177 (N_27177,N_26320,N_25723);
nor U27178 (N_27178,N_25237,N_25635);
nor U27179 (N_27179,N_25725,N_25773);
nor U27180 (N_27180,N_25840,N_26018);
nand U27181 (N_27181,N_25454,N_25203);
and U27182 (N_27182,N_25218,N_25260);
xnor U27183 (N_27183,N_26144,N_26000);
xor U27184 (N_27184,N_25237,N_26173);
nand U27185 (N_27185,N_25641,N_26270);
nor U27186 (N_27186,N_25315,N_25563);
nand U27187 (N_27187,N_26189,N_26210);
and U27188 (N_27188,N_26358,N_25555);
nand U27189 (N_27189,N_25429,N_25236);
and U27190 (N_27190,N_25693,N_25332);
nand U27191 (N_27191,N_25784,N_25324);
xnor U27192 (N_27192,N_26393,N_25733);
or U27193 (N_27193,N_25666,N_25725);
or U27194 (N_27194,N_25447,N_25497);
nand U27195 (N_27195,N_25909,N_26021);
xnor U27196 (N_27196,N_25804,N_25295);
nand U27197 (N_27197,N_26230,N_26002);
xor U27198 (N_27198,N_26081,N_25948);
nor U27199 (N_27199,N_25789,N_25981);
nand U27200 (N_27200,N_25434,N_26118);
nand U27201 (N_27201,N_25655,N_25577);
and U27202 (N_27202,N_25958,N_26148);
xnor U27203 (N_27203,N_26125,N_26056);
nor U27204 (N_27204,N_25890,N_25457);
nor U27205 (N_27205,N_25415,N_25218);
xnor U27206 (N_27206,N_25515,N_25857);
or U27207 (N_27207,N_25619,N_25560);
nand U27208 (N_27208,N_25971,N_26243);
xor U27209 (N_27209,N_25241,N_26353);
and U27210 (N_27210,N_26179,N_25495);
or U27211 (N_27211,N_25704,N_25757);
and U27212 (N_27212,N_25935,N_26122);
nor U27213 (N_27213,N_26198,N_25523);
nand U27214 (N_27214,N_25757,N_25332);
nand U27215 (N_27215,N_25317,N_25993);
or U27216 (N_27216,N_26213,N_25486);
nand U27217 (N_27217,N_26278,N_25321);
nand U27218 (N_27218,N_25775,N_26015);
nand U27219 (N_27219,N_26238,N_26152);
xnor U27220 (N_27220,N_25723,N_26289);
xnor U27221 (N_27221,N_25263,N_25231);
and U27222 (N_27222,N_25632,N_25864);
xnor U27223 (N_27223,N_26304,N_25242);
nor U27224 (N_27224,N_25374,N_25673);
xor U27225 (N_27225,N_25408,N_25871);
nor U27226 (N_27226,N_25335,N_26349);
nand U27227 (N_27227,N_26362,N_26266);
xnor U27228 (N_27228,N_25389,N_25540);
nand U27229 (N_27229,N_25318,N_26340);
or U27230 (N_27230,N_25612,N_25575);
or U27231 (N_27231,N_25912,N_26310);
or U27232 (N_27232,N_26102,N_25698);
nand U27233 (N_27233,N_25380,N_25855);
and U27234 (N_27234,N_25454,N_25527);
and U27235 (N_27235,N_25210,N_25302);
nand U27236 (N_27236,N_25510,N_26375);
xor U27237 (N_27237,N_25490,N_25921);
or U27238 (N_27238,N_25715,N_26383);
xnor U27239 (N_27239,N_26064,N_25545);
or U27240 (N_27240,N_26139,N_25837);
nor U27241 (N_27241,N_25986,N_26371);
nand U27242 (N_27242,N_26046,N_25218);
and U27243 (N_27243,N_25276,N_25202);
xor U27244 (N_27244,N_25670,N_25635);
or U27245 (N_27245,N_25844,N_25611);
and U27246 (N_27246,N_26184,N_25369);
nor U27247 (N_27247,N_26332,N_26301);
xnor U27248 (N_27248,N_25797,N_26345);
or U27249 (N_27249,N_25647,N_26014);
or U27250 (N_27250,N_26262,N_25520);
and U27251 (N_27251,N_25267,N_25819);
and U27252 (N_27252,N_25578,N_25606);
and U27253 (N_27253,N_26160,N_25754);
and U27254 (N_27254,N_25379,N_25879);
xor U27255 (N_27255,N_26342,N_25712);
xnor U27256 (N_27256,N_25358,N_25860);
or U27257 (N_27257,N_26013,N_25915);
or U27258 (N_27258,N_25263,N_26058);
or U27259 (N_27259,N_25679,N_25721);
and U27260 (N_27260,N_25420,N_26186);
and U27261 (N_27261,N_26229,N_25391);
xnor U27262 (N_27262,N_25673,N_26322);
or U27263 (N_27263,N_25618,N_26319);
nor U27264 (N_27264,N_25756,N_26085);
and U27265 (N_27265,N_25495,N_26383);
nand U27266 (N_27266,N_25984,N_26203);
xnor U27267 (N_27267,N_26064,N_25989);
nand U27268 (N_27268,N_25771,N_25323);
nand U27269 (N_27269,N_26117,N_26259);
or U27270 (N_27270,N_25876,N_25241);
xnor U27271 (N_27271,N_25549,N_25974);
nor U27272 (N_27272,N_25555,N_25485);
or U27273 (N_27273,N_26142,N_25496);
nand U27274 (N_27274,N_25336,N_25846);
xnor U27275 (N_27275,N_25781,N_26272);
nor U27276 (N_27276,N_26360,N_25216);
and U27277 (N_27277,N_25242,N_25820);
xor U27278 (N_27278,N_26163,N_25576);
and U27279 (N_27279,N_25827,N_26339);
nand U27280 (N_27280,N_25775,N_25955);
nand U27281 (N_27281,N_25334,N_25839);
nor U27282 (N_27282,N_25473,N_26125);
nand U27283 (N_27283,N_26003,N_25697);
nand U27284 (N_27284,N_25633,N_25205);
or U27285 (N_27285,N_25290,N_25661);
or U27286 (N_27286,N_25261,N_26337);
nand U27287 (N_27287,N_25533,N_25681);
and U27288 (N_27288,N_26176,N_25991);
xnor U27289 (N_27289,N_25435,N_26097);
and U27290 (N_27290,N_26088,N_25831);
xor U27291 (N_27291,N_26354,N_26065);
xor U27292 (N_27292,N_25817,N_25637);
or U27293 (N_27293,N_25440,N_26333);
nor U27294 (N_27294,N_25633,N_25761);
xnor U27295 (N_27295,N_25832,N_26361);
nand U27296 (N_27296,N_26021,N_26395);
nor U27297 (N_27297,N_25791,N_25672);
nand U27298 (N_27298,N_25469,N_26379);
nand U27299 (N_27299,N_25922,N_25495);
nor U27300 (N_27300,N_25712,N_25447);
nor U27301 (N_27301,N_25394,N_25402);
xnor U27302 (N_27302,N_25879,N_25700);
nor U27303 (N_27303,N_25491,N_26289);
and U27304 (N_27304,N_25681,N_25614);
and U27305 (N_27305,N_25375,N_26368);
xor U27306 (N_27306,N_25694,N_25943);
nor U27307 (N_27307,N_26179,N_26338);
xnor U27308 (N_27308,N_25513,N_25455);
and U27309 (N_27309,N_26131,N_25406);
or U27310 (N_27310,N_25891,N_26351);
or U27311 (N_27311,N_26354,N_25631);
or U27312 (N_27312,N_26261,N_25994);
xnor U27313 (N_27313,N_25770,N_25976);
and U27314 (N_27314,N_25582,N_25367);
or U27315 (N_27315,N_26101,N_25318);
nand U27316 (N_27316,N_25836,N_26253);
nand U27317 (N_27317,N_25830,N_25811);
or U27318 (N_27318,N_25931,N_25710);
nand U27319 (N_27319,N_25278,N_25475);
nand U27320 (N_27320,N_26374,N_25929);
xor U27321 (N_27321,N_25727,N_25970);
or U27322 (N_27322,N_25418,N_26014);
nand U27323 (N_27323,N_25217,N_26233);
and U27324 (N_27324,N_25281,N_25933);
nand U27325 (N_27325,N_25803,N_25547);
xor U27326 (N_27326,N_25954,N_25643);
or U27327 (N_27327,N_25646,N_26203);
or U27328 (N_27328,N_25386,N_25341);
xor U27329 (N_27329,N_25521,N_25301);
nand U27330 (N_27330,N_25239,N_25305);
xnor U27331 (N_27331,N_25812,N_25542);
nand U27332 (N_27332,N_25935,N_25773);
nand U27333 (N_27333,N_26291,N_25957);
nor U27334 (N_27334,N_26327,N_25638);
xor U27335 (N_27335,N_25403,N_25535);
and U27336 (N_27336,N_25945,N_26135);
and U27337 (N_27337,N_26367,N_25682);
nand U27338 (N_27338,N_25898,N_25344);
xnor U27339 (N_27339,N_25938,N_26102);
and U27340 (N_27340,N_26165,N_25522);
and U27341 (N_27341,N_25397,N_25374);
nor U27342 (N_27342,N_26372,N_25260);
nor U27343 (N_27343,N_25265,N_25567);
or U27344 (N_27344,N_25569,N_26079);
nor U27345 (N_27345,N_26049,N_26119);
and U27346 (N_27346,N_25523,N_26306);
nand U27347 (N_27347,N_25512,N_25734);
nor U27348 (N_27348,N_25703,N_25882);
or U27349 (N_27349,N_26137,N_25569);
xor U27350 (N_27350,N_25541,N_25435);
nand U27351 (N_27351,N_26145,N_25219);
nor U27352 (N_27352,N_25824,N_25776);
nor U27353 (N_27353,N_25380,N_25521);
and U27354 (N_27354,N_26084,N_26359);
xnor U27355 (N_27355,N_25474,N_26300);
nand U27356 (N_27356,N_25200,N_25439);
and U27357 (N_27357,N_25649,N_25653);
xor U27358 (N_27358,N_26152,N_25687);
or U27359 (N_27359,N_25868,N_25280);
nor U27360 (N_27360,N_26344,N_26266);
and U27361 (N_27361,N_26078,N_25946);
and U27362 (N_27362,N_26223,N_26190);
nand U27363 (N_27363,N_25590,N_26128);
and U27364 (N_27364,N_25213,N_26235);
nand U27365 (N_27365,N_26073,N_26244);
xor U27366 (N_27366,N_25726,N_26248);
nor U27367 (N_27367,N_26212,N_25454);
nand U27368 (N_27368,N_25695,N_26349);
and U27369 (N_27369,N_25972,N_25948);
nand U27370 (N_27370,N_26306,N_26183);
nor U27371 (N_27371,N_25751,N_25761);
nand U27372 (N_27372,N_25268,N_25448);
or U27373 (N_27373,N_25827,N_25800);
and U27374 (N_27374,N_25318,N_26002);
xnor U27375 (N_27375,N_26017,N_25556);
nand U27376 (N_27376,N_26276,N_26211);
or U27377 (N_27377,N_26111,N_26206);
nand U27378 (N_27378,N_25346,N_26216);
nand U27379 (N_27379,N_26279,N_26308);
xnor U27380 (N_27380,N_26360,N_25602);
nor U27381 (N_27381,N_25917,N_25630);
nand U27382 (N_27382,N_25426,N_26110);
and U27383 (N_27383,N_25806,N_26177);
nor U27384 (N_27384,N_25936,N_26252);
nor U27385 (N_27385,N_26015,N_25458);
and U27386 (N_27386,N_25551,N_25767);
nor U27387 (N_27387,N_26277,N_25498);
nand U27388 (N_27388,N_26289,N_25305);
nor U27389 (N_27389,N_25383,N_25885);
or U27390 (N_27390,N_25946,N_26088);
nand U27391 (N_27391,N_25519,N_26153);
or U27392 (N_27392,N_25398,N_25995);
or U27393 (N_27393,N_25476,N_25715);
nand U27394 (N_27394,N_25678,N_25453);
nand U27395 (N_27395,N_25946,N_26001);
xor U27396 (N_27396,N_26214,N_25891);
and U27397 (N_27397,N_26141,N_26035);
and U27398 (N_27398,N_25903,N_26368);
or U27399 (N_27399,N_25559,N_25811);
and U27400 (N_27400,N_26082,N_26328);
and U27401 (N_27401,N_26103,N_26212);
or U27402 (N_27402,N_26010,N_25979);
or U27403 (N_27403,N_25743,N_25511);
xor U27404 (N_27404,N_25776,N_25639);
nor U27405 (N_27405,N_26108,N_26241);
xor U27406 (N_27406,N_25477,N_25988);
xor U27407 (N_27407,N_26351,N_25768);
and U27408 (N_27408,N_25852,N_26074);
or U27409 (N_27409,N_26267,N_25717);
xnor U27410 (N_27410,N_25255,N_26181);
nor U27411 (N_27411,N_26345,N_25223);
and U27412 (N_27412,N_25560,N_25422);
nand U27413 (N_27413,N_25664,N_26330);
nor U27414 (N_27414,N_26187,N_25411);
nor U27415 (N_27415,N_26220,N_25683);
xor U27416 (N_27416,N_25742,N_25409);
and U27417 (N_27417,N_26132,N_26274);
nor U27418 (N_27418,N_25623,N_26222);
nand U27419 (N_27419,N_25466,N_25446);
nand U27420 (N_27420,N_25685,N_26058);
xor U27421 (N_27421,N_26181,N_26008);
nand U27422 (N_27422,N_25340,N_26247);
xnor U27423 (N_27423,N_25374,N_26163);
xnor U27424 (N_27424,N_26240,N_26024);
and U27425 (N_27425,N_25777,N_26142);
nand U27426 (N_27426,N_25450,N_25491);
xnor U27427 (N_27427,N_26245,N_26021);
and U27428 (N_27428,N_25480,N_25312);
nand U27429 (N_27429,N_25650,N_25372);
nand U27430 (N_27430,N_26291,N_25334);
and U27431 (N_27431,N_25550,N_26269);
nand U27432 (N_27432,N_25806,N_25507);
and U27433 (N_27433,N_25805,N_25839);
and U27434 (N_27434,N_25380,N_26091);
nor U27435 (N_27435,N_25845,N_25341);
nand U27436 (N_27436,N_26266,N_25417);
or U27437 (N_27437,N_25778,N_25488);
nor U27438 (N_27438,N_26336,N_26047);
nand U27439 (N_27439,N_25441,N_25316);
nor U27440 (N_27440,N_26288,N_25819);
or U27441 (N_27441,N_26010,N_25549);
and U27442 (N_27442,N_25242,N_25860);
nand U27443 (N_27443,N_25381,N_25235);
and U27444 (N_27444,N_25243,N_25699);
nand U27445 (N_27445,N_25200,N_25264);
or U27446 (N_27446,N_25916,N_25600);
nand U27447 (N_27447,N_26278,N_26011);
nand U27448 (N_27448,N_25496,N_26005);
xor U27449 (N_27449,N_25655,N_25950);
nand U27450 (N_27450,N_25533,N_25639);
xor U27451 (N_27451,N_25806,N_25563);
or U27452 (N_27452,N_26054,N_26271);
nor U27453 (N_27453,N_26173,N_25929);
nor U27454 (N_27454,N_25920,N_26303);
xor U27455 (N_27455,N_26255,N_25526);
or U27456 (N_27456,N_26205,N_25560);
xor U27457 (N_27457,N_26114,N_26297);
nor U27458 (N_27458,N_25681,N_26354);
nand U27459 (N_27459,N_26301,N_25481);
xor U27460 (N_27460,N_25453,N_25312);
nor U27461 (N_27461,N_26378,N_25946);
nand U27462 (N_27462,N_26176,N_25340);
nand U27463 (N_27463,N_26380,N_26146);
xor U27464 (N_27464,N_26293,N_25580);
xor U27465 (N_27465,N_25449,N_26236);
nor U27466 (N_27466,N_26306,N_26286);
nor U27467 (N_27467,N_25522,N_25354);
nand U27468 (N_27468,N_25729,N_26188);
nor U27469 (N_27469,N_26273,N_26000);
xor U27470 (N_27470,N_25783,N_26131);
or U27471 (N_27471,N_26005,N_25473);
nand U27472 (N_27472,N_25251,N_25880);
nand U27473 (N_27473,N_26225,N_25664);
nand U27474 (N_27474,N_25301,N_25884);
nand U27475 (N_27475,N_26285,N_25470);
nand U27476 (N_27476,N_26052,N_25558);
and U27477 (N_27477,N_25304,N_25768);
or U27478 (N_27478,N_26265,N_26323);
or U27479 (N_27479,N_25573,N_25262);
nor U27480 (N_27480,N_25858,N_25805);
xnor U27481 (N_27481,N_25514,N_25679);
nor U27482 (N_27482,N_25513,N_25415);
xnor U27483 (N_27483,N_25743,N_25968);
or U27484 (N_27484,N_25773,N_25962);
and U27485 (N_27485,N_26187,N_25249);
nor U27486 (N_27486,N_26158,N_26221);
xnor U27487 (N_27487,N_25836,N_25787);
nand U27488 (N_27488,N_25980,N_25652);
xnor U27489 (N_27489,N_26302,N_25667);
or U27490 (N_27490,N_25247,N_26258);
xnor U27491 (N_27491,N_25261,N_25664);
nor U27492 (N_27492,N_26355,N_25779);
or U27493 (N_27493,N_25639,N_26118);
nand U27494 (N_27494,N_25303,N_25246);
nor U27495 (N_27495,N_26335,N_25692);
nand U27496 (N_27496,N_25337,N_25373);
xnor U27497 (N_27497,N_25919,N_25586);
and U27498 (N_27498,N_25699,N_25547);
nand U27499 (N_27499,N_25776,N_25965);
xnor U27500 (N_27500,N_25994,N_26165);
or U27501 (N_27501,N_25222,N_25954);
or U27502 (N_27502,N_26187,N_26159);
xor U27503 (N_27503,N_26146,N_26197);
xnor U27504 (N_27504,N_25678,N_25612);
nand U27505 (N_27505,N_25978,N_25697);
or U27506 (N_27506,N_26108,N_26333);
nor U27507 (N_27507,N_26122,N_25844);
and U27508 (N_27508,N_25656,N_25974);
nor U27509 (N_27509,N_25909,N_26335);
nand U27510 (N_27510,N_25410,N_26042);
and U27511 (N_27511,N_25745,N_25738);
nand U27512 (N_27512,N_25495,N_25930);
nor U27513 (N_27513,N_26104,N_25405);
xnor U27514 (N_27514,N_25298,N_26328);
or U27515 (N_27515,N_26088,N_25341);
xor U27516 (N_27516,N_26257,N_26356);
and U27517 (N_27517,N_25589,N_26179);
nand U27518 (N_27518,N_25450,N_26008);
and U27519 (N_27519,N_26249,N_25539);
or U27520 (N_27520,N_25236,N_26132);
and U27521 (N_27521,N_25691,N_25688);
nand U27522 (N_27522,N_25730,N_25358);
xor U27523 (N_27523,N_25435,N_26210);
and U27524 (N_27524,N_25513,N_25284);
nand U27525 (N_27525,N_25397,N_26178);
xor U27526 (N_27526,N_26212,N_26139);
xnor U27527 (N_27527,N_26219,N_25573);
nor U27528 (N_27528,N_25400,N_26306);
or U27529 (N_27529,N_25358,N_25612);
and U27530 (N_27530,N_26248,N_25372);
nor U27531 (N_27531,N_25920,N_25481);
nor U27532 (N_27532,N_25391,N_25452);
nand U27533 (N_27533,N_25241,N_25884);
nand U27534 (N_27534,N_25748,N_25907);
nor U27535 (N_27535,N_25391,N_25897);
and U27536 (N_27536,N_25946,N_25930);
nand U27537 (N_27537,N_25399,N_26288);
nand U27538 (N_27538,N_25736,N_25880);
nand U27539 (N_27539,N_26058,N_25252);
nand U27540 (N_27540,N_25340,N_26370);
and U27541 (N_27541,N_26009,N_26157);
nor U27542 (N_27542,N_26059,N_26046);
xnor U27543 (N_27543,N_25481,N_26302);
xnor U27544 (N_27544,N_25929,N_26276);
or U27545 (N_27545,N_26283,N_25523);
nor U27546 (N_27546,N_25902,N_25222);
or U27547 (N_27547,N_25856,N_25960);
xor U27548 (N_27548,N_25996,N_25677);
or U27549 (N_27549,N_26354,N_25939);
nor U27550 (N_27550,N_25245,N_25383);
xor U27551 (N_27551,N_25411,N_25453);
nand U27552 (N_27552,N_25774,N_25435);
nand U27553 (N_27553,N_25206,N_26107);
and U27554 (N_27554,N_25421,N_25723);
and U27555 (N_27555,N_26087,N_25584);
nand U27556 (N_27556,N_25621,N_25538);
and U27557 (N_27557,N_26042,N_26129);
and U27558 (N_27558,N_26181,N_25966);
and U27559 (N_27559,N_26236,N_25444);
xnor U27560 (N_27560,N_25850,N_25869);
xnor U27561 (N_27561,N_25991,N_25811);
xnor U27562 (N_27562,N_25593,N_25812);
nor U27563 (N_27563,N_25218,N_26354);
or U27564 (N_27564,N_25900,N_25846);
nor U27565 (N_27565,N_26199,N_25899);
or U27566 (N_27566,N_26033,N_26350);
nor U27567 (N_27567,N_26036,N_26235);
or U27568 (N_27568,N_26333,N_26285);
xnor U27569 (N_27569,N_25523,N_25522);
xor U27570 (N_27570,N_26367,N_25936);
nor U27571 (N_27571,N_25207,N_25540);
xnor U27572 (N_27572,N_25559,N_26044);
or U27573 (N_27573,N_25637,N_25416);
and U27574 (N_27574,N_25540,N_25560);
or U27575 (N_27575,N_25560,N_26025);
nor U27576 (N_27576,N_25997,N_25867);
nand U27577 (N_27577,N_25461,N_25210);
nand U27578 (N_27578,N_26100,N_25822);
or U27579 (N_27579,N_26336,N_25306);
and U27580 (N_27580,N_25432,N_26206);
or U27581 (N_27581,N_25588,N_25647);
or U27582 (N_27582,N_25696,N_25730);
xnor U27583 (N_27583,N_26022,N_25427);
and U27584 (N_27584,N_25855,N_25798);
and U27585 (N_27585,N_25230,N_25255);
xor U27586 (N_27586,N_25711,N_25861);
xnor U27587 (N_27587,N_25994,N_26036);
nor U27588 (N_27588,N_26065,N_26051);
xor U27589 (N_27589,N_25843,N_25389);
nand U27590 (N_27590,N_25296,N_25804);
nor U27591 (N_27591,N_25893,N_25413);
xnor U27592 (N_27592,N_25515,N_25626);
nand U27593 (N_27593,N_25683,N_26052);
nand U27594 (N_27594,N_26185,N_26011);
nand U27595 (N_27595,N_26171,N_25874);
nand U27596 (N_27596,N_25461,N_25933);
nand U27597 (N_27597,N_25895,N_26292);
nor U27598 (N_27598,N_26226,N_25491);
or U27599 (N_27599,N_25641,N_26359);
or U27600 (N_27600,N_26641,N_26624);
nand U27601 (N_27601,N_27393,N_26408);
xor U27602 (N_27602,N_26994,N_27136);
nor U27603 (N_27603,N_27459,N_27301);
xor U27604 (N_27604,N_26459,N_26474);
and U27605 (N_27605,N_27138,N_26855);
and U27606 (N_27606,N_27395,N_27058);
nand U27607 (N_27607,N_27519,N_27500);
and U27608 (N_27608,N_27013,N_27348);
xnor U27609 (N_27609,N_27274,N_27465);
nor U27610 (N_27610,N_27026,N_26784);
nor U27611 (N_27611,N_27344,N_26582);
nand U27612 (N_27612,N_27496,N_26669);
xor U27613 (N_27613,N_26511,N_27286);
nor U27614 (N_27614,N_26958,N_26460);
or U27615 (N_27615,N_27197,N_26527);
nor U27616 (N_27616,N_26708,N_27206);
nand U27617 (N_27617,N_26550,N_27285);
or U27618 (N_27618,N_27472,N_26545);
and U27619 (N_27619,N_26993,N_26439);
nor U27620 (N_27620,N_26814,N_26894);
nand U27621 (N_27621,N_27583,N_27124);
or U27622 (N_27622,N_27208,N_27488);
nor U27623 (N_27623,N_26653,N_27094);
xor U27624 (N_27624,N_26904,N_26940);
nand U27625 (N_27625,N_26872,N_27159);
xor U27626 (N_27626,N_26988,N_27232);
and U27627 (N_27627,N_26429,N_27375);
nor U27628 (N_27628,N_26839,N_26650);
nor U27629 (N_27629,N_26404,N_26818);
or U27630 (N_27630,N_27568,N_26926);
or U27631 (N_27631,N_26598,N_27214);
nand U27632 (N_27632,N_26645,N_26970);
nand U27633 (N_27633,N_27421,N_26754);
xor U27634 (N_27634,N_26701,N_26692);
or U27635 (N_27635,N_26447,N_27116);
nor U27636 (N_27636,N_26575,N_27100);
and U27637 (N_27637,N_27433,N_27569);
nand U27638 (N_27638,N_27384,N_27054);
or U27639 (N_27639,N_26472,N_26965);
and U27640 (N_27640,N_26841,N_26978);
and U27641 (N_27641,N_27202,N_26949);
or U27642 (N_27642,N_27552,N_27133);
or U27643 (N_27643,N_26477,N_27516);
and U27644 (N_27644,N_27430,N_27311);
and U27645 (N_27645,N_27553,N_27302);
or U27646 (N_27646,N_26987,N_27529);
nand U27647 (N_27647,N_26829,N_26751);
or U27648 (N_27648,N_26589,N_27570);
nor U27649 (N_27649,N_27059,N_27199);
xnor U27650 (N_27650,N_26743,N_27092);
nor U27651 (N_27651,N_27461,N_26611);
and U27652 (N_27652,N_27271,N_27466);
nor U27653 (N_27653,N_26897,N_27216);
nor U27654 (N_27654,N_26436,N_26485);
or U27655 (N_27655,N_27139,N_27339);
and U27656 (N_27656,N_26973,N_26509);
and U27657 (N_27657,N_26632,N_27024);
nor U27658 (N_27658,N_27134,N_26934);
xor U27659 (N_27659,N_26448,N_27071);
xor U27660 (N_27660,N_26735,N_27505);
and U27661 (N_27661,N_27336,N_27597);
xnor U27662 (N_27662,N_26562,N_26832);
and U27663 (N_27663,N_27480,N_26420);
or U27664 (N_27664,N_27450,N_26608);
or U27665 (N_27665,N_27074,N_27445);
and U27666 (N_27666,N_27317,N_27276);
nand U27667 (N_27667,N_27019,N_26648);
nor U27668 (N_27668,N_26670,N_27104);
nand U27669 (N_27669,N_26785,N_26428);
nand U27670 (N_27670,N_26826,N_26774);
or U27671 (N_27671,N_27371,N_27175);
nand U27672 (N_27672,N_27534,N_26676);
nand U27673 (N_27673,N_27492,N_27145);
nand U27674 (N_27674,N_26452,N_27356);
nor U27675 (N_27675,N_26523,N_27319);
nand U27676 (N_27676,N_27210,N_27008);
and U27677 (N_27677,N_27442,N_26488);
and U27678 (N_27678,N_26732,N_27331);
nor U27679 (N_27679,N_26954,N_26665);
or U27680 (N_27680,N_26552,N_27475);
nor U27681 (N_27681,N_27447,N_26466);
and U27682 (N_27682,N_27556,N_26974);
or U27683 (N_27683,N_26667,N_26528);
nor U27684 (N_27684,N_27086,N_27070);
and U27685 (N_27685,N_26519,N_26601);
nand U27686 (N_27686,N_26685,N_27245);
xor U27687 (N_27687,N_27293,N_26604);
or U27688 (N_27688,N_26504,N_26563);
xor U27689 (N_27689,N_26532,N_27588);
nor U27690 (N_27690,N_27332,N_26433);
and U27691 (N_27691,N_27284,N_27052);
xor U27692 (N_27692,N_26997,N_26462);
nor U27693 (N_27693,N_26757,N_26998);
xor U27694 (N_27694,N_27471,N_26556);
and U27695 (N_27695,N_27030,N_27547);
nor U27696 (N_27696,N_27185,N_26609);
or U27697 (N_27697,N_26649,N_27267);
xnor U27698 (N_27698,N_26765,N_26635);
or U27699 (N_27699,N_27045,N_27165);
xor U27700 (N_27700,N_26790,N_27292);
nor U27701 (N_27701,N_27179,N_27487);
nand U27702 (N_27702,N_26434,N_26764);
xor U27703 (N_27703,N_26400,N_26697);
and U27704 (N_27704,N_26592,N_27053);
or U27705 (N_27705,N_26600,N_27509);
and U27706 (N_27706,N_27571,N_27338);
and U27707 (N_27707,N_26857,N_27237);
and U27708 (N_27708,N_27434,N_26524);
or U27709 (N_27709,N_26664,N_27127);
xor U27710 (N_27710,N_27313,N_27454);
and U27711 (N_27711,N_27296,N_26888);
and U27712 (N_27712,N_26843,N_26744);
xnor U27713 (N_27713,N_27241,N_27040);
or U27714 (N_27714,N_27358,N_26808);
and U27715 (N_27715,N_27028,N_27372);
and U27716 (N_27716,N_26959,N_26567);
nand U27717 (N_27717,N_27464,N_26778);
nand U27718 (N_27718,N_26864,N_26963);
or U27719 (N_27719,N_26554,N_27373);
xor U27720 (N_27720,N_26558,N_26517);
or U27721 (N_27721,N_27424,N_27323);
and U27722 (N_27722,N_26686,N_27536);
xnor U27723 (N_27723,N_27405,N_27204);
nand U27724 (N_27724,N_26457,N_26865);
or U27725 (N_27725,N_27484,N_27451);
or U27726 (N_27726,N_26950,N_26727);
nor U27727 (N_27727,N_26587,N_26724);
and U27728 (N_27728,N_26642,N_27004);
nand U27729 (N_27729,N_26791,N_27361);
or U27730 (N_27730,N_26846,N_27140);
nand U27731 (N_27731,N_26662,N_27404);
and U27732 (N_27732,N_27452,N_26895);
or U27733 (N_27733,N_27119,N_27121);
xnor U27734 (N_27734,N_26631,N_27223);
nor U27735 (N_27735,N_27585,N_27343);
nand U27736 (N_27736,N_27038,N_27158);
or U27737 (N_27737,N_26691,N_26638);
or U27738 (N_27738,N_26551,N_26672);
nand U27739 (N_27739,N_27096,N_27504);
nand U27740 (N_27740,N_26972,N_27391);
nor U27741 (N_27741,N_27173,N_26902);
xnor U27742 (N_27742,N_26489,N_26435);
or U27743 (N_27743,N_26693,N_27577);
nand U27744 (N_27744,N_27221,N_26546);
nor U27745 (N_27745,N_27181,N_26518);
nor U27746 (N_27746,N_27359,N_26866);
nand U27747 (N_27747,N_27575,N_26892);
nor U27748 (N_27748,N_26515,N_26520);
xnor U27749 (N_27749,N_27089,N_27238);
or U27750 (N_27750,N_26695,N_26438);
nor U27751 (N_27751,N_26471,N_26899);
and U27752 (N_27752,N_27226,N_27506);
nor U27753 (N_27753,N_27309,N_27501);
xnor U27754 (N_27754,N_27439,N_27110);
nand U27755 (N_27755,N_27595,N_27530);
xnor U27756 (N_27756,N_27422,N_27299);
nor U27757 (N_27757,N_26753,N_27236);
nor U27758 (N_27758,N_27369,N_27322);
nand U27759 (N_27759,N_27243,N_26737);
nand U27760 (N_27760,N_26657,N_26514);
and U27761 (N_27761,N_26782,N_27493);
xor U27762 (N_27762,N_27025,N_27112);
nand U27763 (N_27763,N_26677,N_26503);
or U27764 (N_27764,N_27362,N_27537);
nor U27765 (N_27765,N_26405,N_26446);
xor U27766 (N_27766,N_27084,N_26752);
nor U27767 (N_27767,N_27360,N_26960);
nand U27768 (N_27768,N_26887,N_27346);
nand U27769 (N_27769,N_27087,N_26789);
and U27770 (N_27770,N_26516,N_27418);
nand U27771 (N_27771,N_26481,N_26507);
and U27772 (N_27772,N_26838,N_26473);
nand U27773 (N_27773,N_27021,N_27258);
nor U27774 (N_27774,N_27065,N_27168);
xnor U27775 (N_27775,N_26454,N_26956);
or U27776 (N_27776,N_27507,N_27381);
or U27777 (N_27777,N_27268,N_27508);
nor U27778 (N_27778,N_27126,N_27032);
nor U27779 (N_27779,N_26805,N_27400);
nand U27780 (N_27780,N_27080,N_26681);
and U27781 (N_27781,N_27003,N_26534);
nor U27782 (N_27782,N_26606,N_26847);
and U27783 (N_27783,N_26898,N_27176);
or U27784 (N_27784,N_26432,N_26853);
xnor U27785 (N_27785,N_26739,N_27253);
nor U27786 (N_27786,N_26756,N_27386);
and U27787 (N_27787,N_26467,N_27357);
nand U27788 (N_27788,N_26759,N_27482);
nand U27789 (N_27789,N_26618,N_27290);
nor U27790 (N_27790,N_26513,N_27446);
nand U27791 (N_27791,N_27209,N_27042);
nor U27792 (N_27792,N_27273,N_27314);
and U27793 (N_27793,N_26840,N_27177);
and U27794 (N_27794,N_26947,N_27060);
or U27795 (N_27795,N_26639,N_27211);
xnor U27796 (N_27796,N_26936,N_26871);
and U27797 (N_27797,N_27098,N_27551);
or U27798 (N_27798,N_27544,N_27022);
and U27799 (N_27799,N_27486,N_27282);
nor U27800 (N_27800,N_27172,N_26798);
or U27801 (N_27801,N_27476,N_27467);
nand U27802 (N_27802,N_27154,N_26482);
or U27803 (N_27803,N_26713,N_26538);
and U27804 (N_27804,N_27051,N_27366);
nor U27805 (N_27805,N_27184,N_27441);
nor U27806 (N_27806,N_27498,N_27540);
nor U27807 (N_27807,N_26647,N_27162);
and U27808 (N_27808,N_27415,N_26529);
xnor U27809 (N_27809,N_26869,N_26905);
nor U27810 (N_27810,N_27294,N_27079);
or U27811 (N_27811,N_27029,N_26748);
xnor U27812 (N_27812,N_26602,N_26456);
nor U27813 (N_27813,N_27122,N_27192);
nor U27814 (N_27814,N_26629,N_26819);
nand U27815 (N_27815,N_26773,N_27351);
and U27816 (N_27816,N_27037,N_26607);
or U27817 (N_27817,N_26971,N_27503);
xor U27818 (N_27818,N_27355,N_27532);
or U27819 (N_27819,N_26415,N_26679);
nand U27820 (N_27820,N_27289,N_26862);
or U27821 (N_27821,N_27423,N_27440);
or U27822 (N_27822,N_26946,N_27244);
nand U27823 (N_27823,N_26923,N_26999);
and U27824 (N_27824,N_27191,N_26644);
nand U27825 (N_27825,N_26766,N_26745);
nor U27826 (N_27826,N_27525,N_27041);
nor U27827 (N_27827,N_26623,N_27228);
or U27828 (N_27828,N_27117,N_26835);
and U27829 (N_27829,N_26579,N_26540);
nand U27830 (N_27830,N_26401,N_27520);
xor U27831 (N_27831,N_26821,N_26793);
xor U27832 (N_27832,N_27420,N_27494);
xnor U27833 (N_27833,N_26740,N_26596);
and U27834 (N_27834,N_27535,N_27269);
xor U27835 (N_27835,N_26569,N_27015);
xnor U27836 (N_27836,N_27164,N_27064);
and U27837 (N_27837,N_26705,N_26564);
nand U27838 (N_27838,N_27016,N_26718);
xor U27839 (N_27839,N_27167,N_27526);
nor U27840 (N_27840,N_27218,N_27468);
or U27841 (N_27841,N_26750,N_27152);
or U27842 (N_27842,N_27156,N_27205);
and U27843 (N_27843,N_26621,N_27304);
or U27844 (N_27844,N_27436,N_26915);
and U27845 (N_27845,N_26512,N_26711);
nor U27846 (N_27846,N_27142,N_26588);
nand U27847 (N_27847,N_27190,N_27573);
nor U27848 (N_27848,N_26730,N_26483);
xnor U27849 (N_27849,N_27334,N_26860);
and U27850 (N_27850,N_27128,N_27095);
nor U27851 (N_27851,N_27131,N_26935);
xnor U27852 (N_27852,N_26414,N_27009);
xor U27853 (N_27853,N_27598,N_26628);
nand U27854 (N_27854,N_27398,N_26694);
and U27855 (N_27855,N_26767,N_27143);
nand U27856 (N_27856,N_27272,N_26937);
and U27857 (N_27857,N_27266,N_27252);
xor U27858 (N_27858,N_26852,N_27521);
nand U27859 (N_27859,N_27246,N_27380);
xor U27860 (N_27860,N_26610,N_26844);
nand U27861 (N_27861,N_27528,N_26702);
and U27862 (N_27862,N_26968,N_27113);
nand U27863 (N_27863,N_26918,N_27248);
xnor U27864 (N_27864,N_27478,N_27264);
nand U27865 (N_27865,N_26521,N_26901);
nor U27866 (N_27866,N_26427,N_26633);
nor U27867 (N_27867,N_26827,N_27410);
nor U27868 (N_27868,N_26830,N_27186);
and U27869 (N_27869,N_27533,N_27596);
or U27870 (N_27870,N_26910,N_26728);
nor U27871 (N_27871,N_27125,N_27287);
nand U27872 (N_27872,N_27378,N_26927);
xnor U27873 (N_27873,N_26712,N_27091);
nor U27874 (N_27874,N_27543,N_27444);
xor U27875 (N_27875,N_26989,N_27189);
xor U27876 (N_27876,N_26555,N_26673);
xnor U27877 (N_27877,N_26465,N_27411);
nor U27878 (N_27878,N_26549,N_26506);
xnor U27879 (N_27879,N_27335,N_26911);
nor U27880 (N_27880,N_26557,N_27067);
xnor U27881 (N_27881,N_27427,N_27169);
and U27882 (N_27882,N_26985,N_26912);
nand U27883 (N_27883,N_26682,N_27278);
xnor U27884 (N_27884,N_26969,N_26553);
nand U27885 (N_27885,N_27036,N_26464);
nand U27886 (N_27886,N_27502,N_26416);
nand U27887 (N_27887,N_26548,N_27578);
and U27888 (N_27888,N_26565,N_27081);
or U27889 (N_27889,N_27342,N_27101);
nand U27890 (N_27890,N_26944,N_26953);
nand U27891 (N_27891,N_27239,N_26842);
or U27892 (N_27892,N_27425,N_26809);
nor U27893 (N_27893,N_27329,N_26799);
and U27894 (N_27894,N_26689,N_27102);
or U27895 (N_27895,N_27324,N_26725);
nand U27896 (N_27896,N_26879,N_26714);
xor U27897 (N_27897,N_27183,N_26812);
nand U27898 (N_27898,N_26680,N_27303);
nor U27899 (N_27899,N_27483,N_26526);
and U27900 (N_27900,N_26403,N_27367);
or U27901 (N_27901,N_26502,N_26537);
or U27902 (N_27902,N_27409,N_26803);
nand U27903 (N_27903,N_27105,N_26794);
xor U27904 (N_27904,N_26729,N_26889);
nor U27905 (N_27905,N_26720,N_27062);
nand U27906 (N_27906,N_27160,N_26499);
or U27907 (N_27907,N_26873,N_26777);
nand U27908 (N_27908,N_27187,N_26850);
nand U27909 (N_27909,N_26617,N_26413);
nand U27910 (N_27910,N_26749,N_26484);
and U27911 (N_27911,N_27230,N_27545);
nand U27912 (N_27912,N_27590,N_26948);
nor U27913 (N_27913,N_26786,N_27407);
and U27914 (N_27914,N_26591,N_26921);
or U27915 (N_27915,N_27277,N_27215);
nand U27916 (N_27916,N_27456,N_27213);
nand U27917 (N_27917,N_27146,N_27001);
nand U27918 (N_27918,N_27443,N_26813);
nand U27919 (N_27919,N_27559,N_27396);
or U27920 (N_27920,N_26619,N_26652);
nor U27921 (N_27921,N_26461,N_27118);
nand U27922 (N_27922,N_26699,N_27163);
or U27923 (N_27923,N_26599,N_27275);
nor U27924 (N_27924,N_27103,N_26731);
nand U27925 (N_27925,N_27408,N_27035);
nand U27926 (N_27926,N_27390,N_27061);
nand U27927 (N_27927,N_26900,N_27229);
nand U27928 (N_27928,N_27147,N_27349);
xnor U27929 (N_27929,N_26833,N_27083);
nand U27930 (N_27930,N_26417,N_27463);
nor U27931 (N_27931,N_27429,N_27082);
xor U27932 (N_27932,N_26468,N_26683);
nor U27933 (N_27933,N_27376,N_26469);
xor U27934 (N_27934,N_27171,N_26738);
xor U27935 (N_27935,N_26654,N_27075);
and U27936 (N_27936,N_26884,N_26792);
xor U27937 (N_27937,N_26962,N_26703);
or U27938 (N_27938,N_27281,N_26533);
and U27939 (N_27939,N_27566,N_26449);
nand U27940 (N_27940,N_27090,N_26580);
xor U27941 (N_27941,N_26834,N_26995);
xnor U27942 (N_27942,N_26836,N_26723);
nor U27943 (N_27943,N_26991,N_27320);
xnor U27944 (N_27944,N_26411,N_27044);
nand U27945 (N_27945,N_26858,N_26658);
or U27946 (N_27946,N_27524,N_27458);
nand U27947 (N_27947,N_26412,N_27259);
nand U27948 (N_27948,N_26674,N_27155);
or U27949 (N_27949,N_26746,N_26781);
or U27950 (N_27950,N_26721,N_27402);
nor U27951 (N_27951,N_27220,N_27477);
xnor U27952 (N_27952,N_27310,N_27203);
nor U27953 (N_27953,N_26547,N_26585);
xnor U27954 (N_27954,N_27288,N_27305);
nor U27955 (N_27955,N_26986,N_27593);
xnor U27956 (N_27956,N_27586,N_27308);
and U27957 (N_27957,N_27383,N_27539);
nor U27958 (N_27958,N_26407,N_27234);
and U27959 (N_27959,N_27263,N_26859);
nand U27960 (N_27960,N_26957,N_26486);
nor U27961 (N_27961,N_26885,N_26581);
xnor U27962 (N_27962,N_26663,N_27150);
nor U27963 (N_27963,N_27511,N_26666);
and U27964 (N_27964,N_27023,N_27068);
nand U27965 (N_27965,N_26525,N_27354);
or U27966 (N_27966,N_26530,N_26849);
or U27967 (N_27967,N_27129,N_26470);
or U27968 (N_27968,N_27564,N_27307);
xor U27969 (N_27969,N_26480,N_27431);
nor U27970 (N_27970,N_26716,N_27546);
or U27971 (N_27971,N_26795,N_27365);
and U27972 (N_27972,N_26583,N_26640);
nor U27973 (N_27973,N_26845,N_27379);
nand U27974 (N_27974,N_26494,N_27517);
nor U27975 (N_27975,N_27257,N_26816);
xnor U27976 (N_27976,N_26458,N_27260);
nor U27977 (N_27977,N_27579,N_27114);
nand U27978 (N_27978,N_26479,N_26425);
nor U27979 (N_27979,N_27262,N_26455);
or U27980 (N_27980,N_26535,N_27574);
and U27981 (N_27981,N_27182,N_26736);
xor U27982 (N_27982,N_26917,N_26930);
nor U27983 (N_27983,N_26430,N_27198);
nor U27984 (N_27984,N_27499,N_27018);
and U27985 (N_27985,N_27397,N_27219);
nor U27986 (N_27986,N_27194,N_26637);
and U27987 (N_27987,N_26584,N_26951);
and U27988 (N_27988,N_26976,N_26522);
nand U27989 (N_27989,N_27078,N_26938);
or U27990 (N_27990,N_26593,N_26614);
xnor U27991 (N_27991,N_27581,N_26955);
nand U27992 (N_27992,N_27170,N_27561);
nor U27993 (N_27993,N_26924,N_27161);
nor U27994 (N_27994,N_26801,N_27312);
xor U27995 (N_27995,N_27031,N_27584);
xor U27996 (N_27996,N_26559,N_26780);
nor U27997 (N_27997,N_27120,N_26800);
nand U27998 (N_27998,N_26874,N_27063);
and U27999 (N_27999,N_26913,N_26939);
and U28000 (N_28000,N_26423,N_27151);
xnor U28001 (N_28001,N_26931,N_27148);
xor U28002 (N_28002,N_27270,N_27069);
or U28003 (N_28003,N_26544,N_26861);
nor U28004 (N_28004,N_26646,N_27123);
xnor U28005 (N_28005,N_26687,N_27562);
xor U28006 (N_28006,N_27033,N_27453);
nand U28007 (N_28007,N_27563,N_26797);
nand U28008 (N_28008,N_26586,N_27006);
xor U28009 (N_28009,N_27193,N_27283);
or U28010 (N_28010,N_26651,N_27256);
xor U28011 (N_28011,N_26903,N_27377);
xor U28012 (N_28012,N_27353,N_26594);
xor U28013 (N_28013,N_27251,N_27178);
or U28014 (N_28014,N_27428,N_26990);
and U28015 (N_28015,N_27485,N_26914);
xor U28016 (N_28016,N_26541,N_26788);
or U28017 (N_28017,N_27135,N_26979);
and U28018 (N_28018,N_26487,N_27093);
and U28019 (N_28019,N_27394,N_26571);
nand U28020 (N_28020,N_27325,N_26908);
and U28021 (N_28021,N_27416,N_27412);
nor U28022 (N_28022,N_27157,N_26597);
xor U28023 (N_28023,N_26445,N_26932);
or U28024 (N_28024,N_26876,N_26984);
or U28025 (N_28025,N_27388,N_26722);
or U28026 (N_28026,N_26442,N_27300);
xnor U28027 (N_28027,N_27099,N_27457);
nor U28028 (N_28028,N_26823,N_26402);
nor U28029 (N_28029,N_26967,N_27510);
nor U28030 (N_28030,N_27531,N_27414);
and U28031 (N_28031,N_26925,N_26536);
nor U28032 (N_28032,N_26761,N_26741);
or U28033 (N_28033,N_26496,N_26568);
xor U28034 (N_28034,N_26421,N_27490);
nor U28035 (N_28035,N_27330,N_26636);
and U28036 (N_28036,N_27587,N_27523);
and U28037 (N_28037,N_27249,N_27316);
xor U28038 (N_28038,N_27491,N_26762);
nor U28039 (N_28039,N_27049,N_27557);
nor U28040 (N_28040,N_26775,N_27011);
and U28041 (N_28041,N_26877,N_27130);
xor U28042 (N_28042,N_26660,N_26776);
nand U28043 (N_28043,N_26804,N_26922);
nand U28044 (N_28044,N_27389,N_26878);
or U28045 (N_28045,N_27227,N_26709);
and U28046 (N_28046,N_27195,N_27470);
nand U28047 (N_28047,N_26802,N_26578);
or U28048 (N_28048,N_27034,N_27550);
nor U28049 (N_28049,N_26981,N_26570);
nor U28050 (N_28050,N_26495,N_27554);
xnor U28051 (N_28051,N_26612,N_26690);
nor U28052 (N_28052,N_27462,N_26431);
nor U28053 (N_28053,N_27403,N_26419);
nor U28054 (N_28054,N_26856,N_27326);
nand U28055 (N_28055,N_26625,N_27180);
and U28056 (N_28056,N_27497,N_26909);
nor U28057 (N_28057,N_26531,N_27043);
nor U28058 (N_28058,N_26719,N_26406);
and U28059 (N_28059,N_27291,N_27072);
nor U28060 (N_28060,N_26490,N_26573);
xnor U28061 (N_28061,N_27419,N_26706);
nor U28062 (N_28062,N_27374,N_26620);
nor U28063 (N_28063,N_26977,N_27406);
nor U28064 (N_28064,N_26498,N_26510);
nand U28065 (N_28065,N_27002,N_26707);
and U28066 (N_28066,N_26867,N_26811);
xor U28067 (N_28067,N_26964,N_26615);
xnor U28068 (N_28068,N_26890,N_26875);
and U28069 (N_28069,N_27242,N_26848);
nor U28070 (N_28070,N_26613,N_26671);
nor U28071 (N_28071,N_26574,N_26768);
or U28072 (N_28072,N_27153,N_27261);
and U28073 (N_28073,N_26919,N_26772);
or U28074 (N_28074,N_26975,N_26418);
and U28075 (N_28075,N_26543,N_27254);
nand U28076 (N_28076,N_27144,N_27481);
xnor U28077 (N_28077,N_27088,N_26688);
and U28078 (N_28078,N_27166,N_27318);
or U28079 (N_28079,N_26576,N_27538);
nand U28080 (N_28080,N_27141,N_26726);
nand U28081 (N_28081,N_27247,N_27435);
nand U28082 (N_28082,N_26450,N_26831);
or U28083 (N_28083,N_26920,N_27201);
nand U28084 (N_28084,N_27111,N_27265);
or U28085 (N_28085,N_26661,N_26815);
nand U28086 (N_28086,N_27306,N_27555);
and U28087 (N_28087,N_27340,N_26605);
and U28088 (N_28088,N_26755,N_27240);
or U28089 (N_28089,N_26929,N_27438);
or U28090 (N_28090,N_27315,N_27558);
and U28091 (N_28091,N_27515,N_26542);
nor U28092 (N_28092,N_27364,N_26453);
nor U28093 (N_28093,N_26655,N_27222);
or U28094 (N_28094,N_26851,N_27512);
or U28095 (N_28095,N_27235,N_27327);
nor U28096 (N_28096,N_27565,N_26476);
or U28097 (N_28097,N_27109,N_26539);
nand U28098 (N_28098,N_27077,N_26966);
and U28099 (N_28099,N_27056,N_27297);
nand U28100 (N_28100,N_27572,N_26643);
and U28101 (N_28101,N_27212,N_26616);
or U28102 (N_28102,N_26942,N_26822);
xor U28103 (N_28103,N_26668,N_27055);
or U28104 (N_28104,N_27548,N_27132);
and U28105 (N_28105,N_26992,N_27250);
or U28106 (N_28106,N_27066,N_27233);
or U28107 (N_28107,N_26881,N_27370);
xor U28108 (N_28108,N_26820,N_26742);
and U28109 (N_28109,N_27591,N_27225);
xnor U28110 (N_28110,N_26560,N_26566);
nand U28111 (N_28111,N_27000,N_27417);
nand U28112 (N_28112,N_27455,N_27017);
xor U28113 (N_28113,N_27217,N_27027);
nand U28114 (N_28114,N_27298,N_27460);
and U28115 (N_28115,N_27449,N_26996);
or U28116 (N_28116,N_26603,N_27295);
xor U28117 (N_28117,N_27200,N_26684);
xor U28118 (N_28118,N_27073,N_26817);
or U28119 (N_28119,N_27399,N_27474);
xnor U28120 (N_28120,N_26928,N_27255);
or U28121 (N_28121,N_26627,N_26696);
and U28122 (N_28122,N_27594,N_27328);
nand U28123 (N_28123,N_27580,N_27448);
nand U28124 (N_28124,N_26444,N_26441);
or U28125 (N_28125,N_27020,N_27576);
or U28126 (N_28126,N_27085,N_26678);
or U28127 (N_28127,N_27107,N_27341);
nor U28128 (N_28128,N_27392,N_26760);
nand U28129 (N_28129,N_27387,N_26493);
and U28130 (N_28130,N_27014,N_27513);
xnor U28131 (N_28131,N_26717,N_27469);
nor U28132 (N_28132,N_26983,N_27489);
and U28133 (N_28133,N_27337,N_26410);
nand U28134 (N_28134,N_26916,N_27224);
or U28135 (N_28135,N_26491,N_27350);
or U28136 (N_28136,N_26577,N_26810);
or U28137 (N_28137,N_27437,N_26733);
or U28138 (N_28138,N_27010,N_27599);
nor U28139 (N_28139,N_26828,N_26700);
nor U28140 (N_28140,N_27207,N_26945);
nand U28141 (N_28141,N_26758,N_27048);
nand U28142 (N_28142,N_27280,N_26475);
nor U28143 (N_28143,N_27368,N_26886);
nand U28144 (N_28144,N_26882,N_26837);
xnor U28145 (N_28145,N_26941,N_27321);
or U28146 (N_28146,N_26590,N_26409);
or U28147 (N_28147,N_27522,N_26492);
and U28148 (N_28148,N_27345,N_27047);
and U28149 (N_28149,N_26443,N_27231);
xnor U28150 (N_28150,N_26508,N_27057);
nand U28151 (N_28151,N_26704,N_27514);
xnor U28152 (N_28152,N_26779,N_27007);
xor U28153 (N_28153,N_26659,N_26863);
nor U28154 (N_28154,N_27149,N_26893);
and U28155 (N_28155,N_26422,N_26715);
or U28156 (N_28156,N_26501,N_26426);
nor U28157 (N_28157,N_27549,N_27115);
nor U28158 (N_28158,N_27541,N_26626);
xnor U28159 (N_28159,N_26463,N_26883);
xor U28160 (N_28160,N_27382,N_27352);
nand U28161 (N_28161,N_27012,N_26437);
xor U28162 (N_28162,N_26943,N_26933);
or U28163 (N_28163,N_27363,N_26500);
nand U28164 (N_28164,N_27542,N_26451);
xnor U28165 (N_28165,N_27196,N_27050);
nor U28166 (N_28166,N_26824,N_27560);
nand U28167 (N_28167,N_27005,N_26880);
nand U28168 (N_28168,N_27401,N_26825);
and U28169 (N_28169,N_26796,N_27188);
nor U28170 (N_28170,N_27426,N_26807);
or U28171 (N_28171,N_27518,N_26675);
xor U28172 (N_28172,N_27473,N_26440);
nor U28173 (N_28173,N_26770,N_26734);
or U28174 (N_28174,N_27567,N_26710);
or U28175 (N_28175,N_26783,N_26747);
and U28176 (N_28176,N_26854,N_26505);
nor U28177 (N_28177,N_27333,N_27174);
nand U28178 (N_28178,N_26806,N_26891);
nand U28179 (N_28179,N_26868,N_27097);
and U28180 (N_28180,N_27582,N_26982);
or U28181 (N_28181,N_26896,N_26478);
nand U28182 (N_28182,N_27106,N_27347);
xnor U28183 (N_28183,N_27279,N_26595);
or U28184 (N_28184,N_26572,N_27108);
nand U28185 (N_28185,N_26424,N_26497);
nand U28186 (N_28186,N_27039,N_26980);
and U28187 (N_28187,N_26961,N_27432);
or U28188 (N_28188,N_26763,N_27046);
or U28189 (N_28189,N_27385,N_26952);
or U28190 (N_28190,N_27413,N_26656);
nand U28191 (N_28191,N_26698,N_27592);
and U28192 (N_28192,N_27495,N_27527);
and U28193 (N_28193,N_26870,N_26787);
nand U28194 (N_28194,N_26630,N_26771);
or U28195 (N_28195,N_26769,N_26906);
xnor U28196 (N_28196,N_26561,N_26907);
and U28197 (N_28197,N_26622,N_26634);
or U28198 (N_28198,N_27076,N_27589);
or U28199 (N_28199,N_27137,N_27479);
xnor U28200 (N_28200,N_27579,N_27192);
and U28201 (N_28201,N_27270,N_26501);
and U28202 (N_28202,N_27296,N_27491);
or U28203 (N_28203,N_27120,N_27572);
and U28204 (N_28204,N_27256,N_27048);
and U28205 (N_28205,N_27457,N_26777);
nor U28206 (N_28206,N_26907,N_26745);
nand U28207 (N_28207,N_26730,N_26545);
and U28208 (N_28208,N_26913,N_27071);
and U28209 (N_28209,N_26583,N_26919);
nand U28210 (N_28210,N_27575,N_27016);
and U28211 (N_28211,N_27288,N_26768);
nor U28212 (N_28212,N_27585,N_27090);
nand U28213 (N_28213,N_26816,N_26998);
nor U28214 (N_28214,N_27356,N_27522);
or U28215 (N_28215,N_27176,N_26491);
nand U28216 (N_28216,N_27504,N_26771);
xor U28217 (N_28217,N_27530,N_27067);
or U28218 (N_28218,N_26717,N_27455);
or U28219 (N_28219,N_27143,N_26480);
xor U28220 (N_28220,N_27563,N_27032);
and U28221 (N_28221,N_27029,N_26657);
nand U28222 (N_28222,N_26684,N_27559);
nor U28223 (N_28223,N_26908,N_26512);
nand U28224 (N_28224,N_26888,N_27256);
or U28225 (N_28225,N_27111,N_27134);
nor U28226 (N_28226,N_26612,N_27117);
xor U28227 (N_28227,N_26703,N_27540);
and U28228 (N_28228,N_26420,N_26933);
nand U28229 (N_28229,N_26792,N_26800);
or U28230 (N_28230,N_26939,N_26738);
xor U28231 (N_28231,N_27313,N_26548);
nor U28232 (N_28232,N_26408,N_27083);
and U28233 (N_28233,N_27018,N_26506);
or U28234 (N_28234,N_26749,N_27594);
xnor U28235 (N_28235,N_27523,N_26649);
or U28236 (N_28236,N_27365,N_26411);
and U28237 (N_28237,N_27132,N_26481);
nand U28238 (N_28238,N_27524,N_26597);
nor U28239 (N_28239,N_27110,N_27151);
or U28240 (N_28240,N_26989,N_27258);
and U28241 (N_28241,N_27055,N_27078);
or U28242 (N_28242,N_26934,N_26745);
nor U28243 (N_28243,N_27045,N_26859);
and U28244 (N_28244,N_26426,N_27325);
or U28245 (N_28245,N_27393,N_27517);
nor U28246 (N_28246,N_26437,N_26729);
or U28247 (N_28247,N_26478,N_27245);
xor U28248 (N_28248,N_27116,N_26734);
or U28249 (N_28249,N_27553,N_26766);
or U28250 (N_28250,N_26653,N_27245);
xor U28251 (N_28251,N_27523,N_27214);
xnor U28252 (N_28252,N_26529,N_26441);
and U28253 (N_28253,N_26805,N_27515);
and U28254 (N_28254,N_26411,N_26948);
or U28255 (N_28255,N_26565,N_26625);
nand U28256 (N_28256,N_27396,N_27576);
nor U28257 (N_28257,N_27157,N_26904);
nor U28258 (N_28258,N_27536,N_27006);
or U28259 (N_28259,N_26980,N_27474);
xor U28260 (N_28260,N_27432,N_27486);
nand U28261 (N_28261,N_26471,N_27517);
or U28262 (N_28262,N_27439,N_26925);
nor U28263 (N_28263,N_26695,N_26801);
nor U28264 (N_28264,N_26783,N_26617);
xor U28265 (N_28265,N_26692,N_27535);
nand U28266 (N_28266,N_26470,N_26742);
and U28267 (N_28267,N_27397,N_27051);
or U28268 (N_28268,N_27316,N_27330);
or U28269 (N_28269,N_26888,N_26793);
xnor U28270 (N_28270,N_26568,N_27166);
and U28271 (N_28271,N_27347,N_26525);
and U28272 (N_28272,N_27441,N_27233);
nand U28273 (N_28273,N_27248,N_26540);
and U28274 (N_28274,N_27362,N_27207);
nor U28275 (N_28275,N_26701,N_26607);
nand U28276 (N_28276,N_27378,N_27486);
nor U28277 (N_28277,N_27249,N_26411);
or U28278 (N_28278,N_27264,N_26739);
xor U28279 (N_28279,N_26618,N_26407);
nand U28280 (N_28280,N_27358,N_26872);
xor U28281 (N_28281,N_26439,N_27233);
or U28282 (N_28282,N_26491,N_27085);
xor U28283 (N_28283,N_26786,N_27290);
nand U28284 (N_28284,N_27585,N_26669);
and U28285 (N_28285,N_26911,N_26404);
and U28286 (N_28286,N_26955,N_26624);
xor U28287 (N_28287,N_27476,N_26760);
nor U28288 (N_28288,N_26488,N_27320);
xnor U28289 (N_28289,N_27492,N_26882);
and U28290 (N_28290,N_26468,N_27279);
nor U28291 (N_28291,N_27120,N_27583);
and U28292 (N_28292,N_27547,N_27542);
or U28293 (N_28293,N_26533,N_27092);
xor U28294 (N_28294,N_26670,N_27470);
and U28295 (N_28295,N_27299,N_27450);
or U28296 (N_28296,N_26944,N_27288);
xor U28297 (N_28297,N_26995,N_26741);
and U28298 (N_28298,N_27355,N_26516);
and U28299 (N_28299,N_26639,N_26729);
and U28300 (N_28300,N_26550,N_26963);
or U28301 (N_28301,N_26877,N_26999);
xor U28302 (N_28302,N_26431,N_26517);
or U28303 (N_28303,N_26762,N_27563);
nand U28304 (N_28304,N_26400,N_26590);
or U28305 (N_28305,N_26584,N_26517);
nand U28306 (N_28306,N_26853,N_26869);
and U28307 (N_28307,N_26559,N_27578);
xnor U28308 (N_28308,N_27292,N_26811);
or U28309 (N_28309,N_26827,N_27043);
nor U28310 (N_28310,N_26703,N_27321);
xor U28311 (N_28311,N_26774,N_27317);
and U28312 (N_28312,N_27054,N_27030);
or U28313 (N_28313,N_26426,N_27452);
nand U28314 (N_28314,N_27300,N_27588);
and U28315 (N_28315,N_27397,N_26409);
xnor U28316 (N_28316,N_27460,N_26899);
xor U28317 (N_28317,N_27300,N_26897);
nor U28318 (N_28318,N_27268,N_27109);
and U28319 (N_28319,N_27085,N_27342);
or U28320 (N_28320,N_27184,N_27123);
nand U28321 (N_28321,N_26997,N_26805);
and U28322 (N_28322,N_27408,N_27111);
xor U28323 (N_28323,N_26512,N_26506);
nor U28324 (N_28324,N_26871,N_26776);
or U28325 (N_28325,N_26629,N_27280);
nand U28326 (N_28326,N_26693,N_27578);
xor U28327 (N_28327,N_26955,N_27343);
and U28328 (N_28328,N_27560,N_27311);
nand U28329 (N_28329,N_27374,N_27485);
nand U28330 (N_28330,N_27266,N_27082);
and U28331 (N_28331,N_26990,N_26689);
nor U28332 (N_28332,N_27198,N_27168);
xnor U28333 (N_28333,N_26788,N_26548);
nand U28334 (N_28334,N_26759,N_26634);
or U28335 (N_28335,N_26794,N_27208);
nor U28336 (N_28336,N_26683,N_26728);
xnor U28337 (N_28337,N_26907,N_27292);
xor U28338 (N_28338,N_27482,N_26488);
or U28339 (N_28339,N_26435,N_26409);
nor U28340 (N_28340,N_27206,N_26470);
and U28341 (N_28341,N_27253,N_27199);
nor U28342 (N_28342,N_27126,N_27146);
or U28343 (N_28343,N_27147,N_27493);
nor U28344 (N_28344,N_27548,N_27226);
xnor U28345 (N_28345,N_26846,N_26821);
nand U28346 (N_28346,N_27224,N_26627);
or U28347 (N_28347,N_27558,N_27360);
or U28348 (N_28348,N_27273,N_26562);
nor U28349 (N_28349,N_26529,N_26475);
and U28350 (N_28350,N_26491,N_26827);
and U28351 (N_28351,N_26570,N_27537);
nor U28352 (N_28352,N_26445,N_27206);
nand U28353 (N_28353,N_27155,N_27373);
nor U28354 (N_28354,N_27366,N_27517);
or U28355 (N_28355,N_27196,N_26750);
and U28356 (N_28356,N_26578,N_26798);
or U28357 (N_28357,N_26944,N_26594);
xor U28358 (N_28358,N_27159,N_27298);
or U28359 (N_28359,N_26793,N_27108);
xnor U28360 (N_28360,N_27573,N_26608);
or U28361 (N_28361,N_27440,N_27175);
or U28362 (N_28362,N_27235,N_26859);
nand U28363 (N_28363,N_27177,N_27286);
and U28364 (N_28364,N_26446,N_27006);
xor U28365 (N_28365,N_26771,N_27443);
nor U28366 (N_28366,N_27576,N_26806);
nand U28367 (N_28367,N_27460,N_26916);
nor U28368 (N_28368,N_27344,N_27175);
nand U28369 (N_28369,N_26754,N_26818);
or U28370 (N_28370,N_26972,N_27244);
xor U28371 (N_28371,N_26978,N_27422);
xor U28372 (N_28372,N_27201,N_26556);
xnor U28373 (N_28373,N_27530,N_27238);
and U28374 (N_28374,N_26577,N_26911);
and U28375 (N_28375,N_27122,N_27372);
nand U28376 (N_28376,N_27035,N_26498);
nor U28377 (N_28377,N_27173,N_26823);
xor U28378 (N_28378,N_27533,N_26953);
and U28379 (N_28379,N_27552,N_27297);
nand U28380 (N_28380,N_26781,N_27080);
nand U28381 (N_28381,N_27563,N_26545);
nor U28382 (N_28382,N_27585,N_26444);
nor U28383 (N_28383,N_27258,N_26550);
nor U28384 (N_28384,N_26658,N_27571);
nand U28385 (N_28385,N_27568,N_26889);
nor U28386 (N_28386,N_26642,N_26568);
and U28387 (N_28387,N_26943,N_27512);
or U28388 (N_28388,N_26553,N_27185);
nor U28389 (N_28389,N_27172,N_26975);
nand U28390 (N_28390,N_27019,N_27044);
nand U28391 (N_28391,N_27026,N_27388);
nor U28392 (N_28392,N_27258,N_27528);
nand U28393 (N_28393,N_26627,N_27011);
nor U28394 (N_28394,N_26926,N_26868);
or U28395 (N_28395,N_27076,N_27103);
xnor U28396 (N_28396,N_27268,N_26508);
or U28397 (N_28397,N_27251,N_26725);
or U28398 (N_28398,N_26691,N_26534);
and U28399 (N_28399,N_27078,N_26485);
and U28400 (N_28400,N_27124,N_27166);
or U28401 (N_28401,N_26590,N_26657);
xnor U28402 (N_28402,N_26475,N_26881);
nand U28403 (N_28403,N_27526,N_27197);
nand U28404 (N_28404,N_26808,N_27061);
nor U28405 (N_28405,N_27592,N_26756);
or U28406 (N_28406,N_27197,N_27033);
xor U28407 (N_28407,N_27513,N_26884);
and U28408 (N_28408,N_26544,N_26470);
nand U28409 (N_28409,N_27081,N_26868);
nand U28410 (N_28410,N_27417,N_27339);
nand U28411 (N_28411,N_27054,N_26760);
or U28412 (N_28412,N_26740,N_26609);
nor U28413 (N_28413,N_26757,N_27015);
xor U28414 (N_28414,N_27273,N_26610);
nand U28415 (N_28415,N_27113,N_27278);
nand U28416 (N_28416,N_26633,N_26532);
or U28417 (N_28417,N_26651,N_26626);
and U28418 (N_28418,N_27138,N_26447);
xnor U28419 (N_28419,N_26633,N_26563);
and U28420 (N_28420,N_26488,N_27305);
xnor U28421 (N_28421,N_27392,N_26619);
or U28422 (N_28422,N_26727,N_27582);
nand U28423 (N_28423,N_26691,N_27483);
xor U28424 (N_28424,N_26885,N_27541);
xnor U28425 (N_28425,N_26817,N_26738);
xnor U28426 (N_28426,N_26788,N_26749);
xor U28427 (N_28427,N_27273,N_27064);
nor U28428 (N_28428,N_27319,N_27095);
xnor U28429 (N_28429,N_26678,N_27303);
nand U28430 (N_28430,N_27049,N_26611);
or U28431 (N_28431,N_27331,N_26974);
or U28432 (N_28432,N_27123,N_26551);
xor U28433 (N_28433,N_26453,N_26698);
nand U28434 (N_28434,N_27144,N_26656);
nor U28435 (N_28435,N_27522,N_27516);
nand U28436 (N_28436,N_27208,N_27469);
nor U28437 (N_28437,N_27160,N_26696);
and U28438 (N_28438,N_27142,N_26992);
xor U28439 (N_28439,N_26864,N_26772);
nand U28440 (N_28440,N_27501,N_27526);
nand U28441 (N_28441,N_27507,N_27167);
nor U28442 (N_28442,N_26963,N_26890);
nor U28443 (N_28443,N_26726,N_26734);
nand U28444 (N_28444,N_26421,N_27176);
xor U28445 (N_28445,N_26871,N_27179);
and U28446 (N_28446,N_26984,N_26709);
or U28447 (N_28447,N_26745,N_27418);
nor U28448 (N_28448,N_27326,N_27355);
or U28449 (N_28449,N_27463,N_27362);
xor U28450 (N_28450,N_27019,N_26629);
nand U28451 (N_28451,N_26688,N_26719);
nor U28452 (N_28452,N_26540,N_27126);
xnor U28453 (N_28453,N_26583,N_26826);
nor U28454 (N_28454,N_26666,N_27096);
or U28455 (N_28455,N_27436,N_26679);
nand U28456 (N_28456,N_26986,N_26788);
or U28457 (N_28457,N_27004,N_27011);
and U28458 (N_28458,N_26775,N_27564);
and U28459 (N_28459,N_27224,N_26912);
or U28460 (N_28460,N_27230,N_26986);
or U28461 (N_28461,N_26890,N_26545);
or U28462 (N_28462,N_26668,N_27450);
nand U28463 (N_28463,N_27559,N_27430);
nor U28464 (N_28464,N_27264,N_26923);
or U28465 (N_28465,N_26792,N_26995);
nor U28466 (N_28466,N_26668,N_26567);
nor U28467 (N_28467,N_26558,N_26412);
and U28468 (N_28468,N_26986,N_27288);
and U28469 (N_28469,N_26456,N_27008);
xor U28470 (N_28470,N_27597,N_26519);
or U28471 (N_28471,N_27475,N_26504);
or U28472 (N_28472,N_27317,N_26966);
and U28473 (N_28473,N_27018,N_27523);
nand U28474 (N_28474,N_26880,N_26975);
xor U28475 (N_28475,N_27044,N_26570);
nand U28476 (N_28476,N_27365,N_26653);
or U28477 (N_28477,N_26681,N_26831);
or U28478 (N_28478,N_27545,N_27145);
and U28479 (N_28479,N_26473,N_27501);
xor U28480 (N_28480,N_26792,N_27223);
and U28481 (N_28481,N_27296,N_27421);
and U28482 (N_28482,N_27461,N_27198);
or U28483 (N_28483,N_26918,N_27042);
and U28484 (N_28484,N_26917,N_26436);
and U28485 (N_28485,N_26581,N_27456);
or U28486 (N_28486,N_26604,N_27065);
nor U28487 (N_28487,N_26677,N_26630);
xor U28488 (N_28488,N_27084,N_27509);
xnor U28489 (N_28489,N_26835,N_26785);
or U28490 (N_28490,N_27339,N_26951);
and U28491 (N_28491,N_26718,N_27599);
and U28492 (N_28492,N_27478,N_27275);
nor U28493 (N_28493,N_26677,N_27202);
or U28494 (N_28494,N_26964,N_27166);
and U28495 (N_28495,N_26413,N_27595);
and U28496 (N_28496,N_27316,N_26588);
nor U28497 (N_28497,N_27312,N_26650);
or U28498 (N_28498,N_27430,N_26996);
nand U28499 (N_28499,N_26622,N_27034);
or U28500 (N_28500,N_27421,N_26979);
and U28501 (N_28501,N_27511,N_26903);
or U28502 (N_28502,N_26564,N_26792);
nor U28503 (N_28503,N_26773,N_26986);
nor U28504 (N_28504,N_27353,N_27541);
or U28505 (N_28505,N_27317,N_26633);
nor U28506 (N_28506,N_27415,N_26842);
nand U28507 (N_28507,N_26699,N_27503);
nor U28508 (N_28508,N_26878,N_27343);
nand U28509 (N_28509,N_27178,N_26444);
or U28510 (N_28510,N_27102,N_27132);
xor U28511 (N_28511,N_26828,N_27330);
or U28512 (N_28512,N_26781,N_27139);
and U28513 (N_28513,N_27473,N_26437);
or U28514 (N_28514,N_27582,N_27309);
xor U28515 (N_28515,N_27131,N_27497);
and U28516 (N_28516,N_27593,N_26950);
nand U28517 (N_28517,N_27567,N_26647);
nor U28518 (N_28518,N_26732,N_26405);
or U28519 (N_28519,N_26540,N_26947);
nor U28520 (N_28520,N_27335,N_26568);
nand U28521 (N_28521,N_27302,N_26669);
nand U28522 (N_28522,N_27564,N_26639);
nor U28523 (N_28523,N_26822,N_26557);
xnor U28524 (N_28524,N_26952,N_26997);
xor U28525 (N_28525,N_27057,N_27193);
or U28526 (N_28526,N_27549,N_26733);
or U28527 (N_28527,N_27287,N_26461);
xnor U28528 (N_28528,N_27380,N_26565);
and U28529 (N_28529,N_27201,N_26505);
and U28530 (N_28530,N_26947,N_27035);
or U28531 (N_28531,N_26927,N_26828);
nand U28532 (N_28532,N_27305,N_27254);
nand U28533 (N_28533,N_27200,N_26765);
or U28534 (N_28534,N_26527,N_27485);
xor U28535 (N_28535,N_26668,N_26571);
or U28536 (N_28536,N_26942,N_26971);
and U28537 (N_28537,N_26471,N_26655);
nand U28538 (N_28538,N_26840,N_27560);
nor U28539 (N_28539,N_27052,N_26755);
and U28540 (N_28540,N_27118,N_26578);
or U28541 (N_28541,N_26696,N_27473);
and U28542 (N_28542,N_26576,N_27073);
or U28543 (N_28543,N_27196,N_26828);
xnor U28544 (N_28544,N_26599,N_27499);
or U28545 (N_28545,N_26412,N_27536);
or U28546 (N_28546,N_27373,N_26755);
nand U28547 (N_28547,N_27139,N_26488);
or U28548 (N_28548,N_26822,N_27510);
nand U28549 (N_28549,N_26509,N_26591);
xnor U28550 (N_28550,N_26613,N_27117);
xnor U28551 (N_28551,N_27313,N_26880);
or U28552 (N_28552,N_27096,N_26679);
xnor U28553 (N_28553,N_26974,N_27490);
and U28554 (N_28554,N_27588,N_27573);
nor U28555 (N_28555,N_26654,N_27121);
nor U28556 (N_28556,N_26601,N_26477);
or U28557 (N_28557,N_26756,N_26966);
nand U28558 (N_28558,N_26546,N_27583);
nand U28559 (N_28559,N_27515,N_27020);
or U28560 (N_28560,N_27392,N_26920);
nor U28561 (N_28561,N_27329,N_26644);
and U28562 (N_28562,N_27116,N_27129);
or U28563 (N_28563,N_26763,N_27273);
xor U28564 (N_28564,N_26798,N_26730);
nor U28565 (N_28565,N_26472,N_27555);
and U28566 (N_28566,N_26519,N_26994);
and U28567 (N_28567,N_26644,N_27268);
nand U28568 (N_28568,N_26403,N_26915);
nand U28569 (N_28569,N_27459,N_27232);
or U28570 (N_28570,N_26940,N_27330);
or U28571 (N_28571,N_26709,N_27522);
nor U28572 (N_28572,N_27272,N_27585);
nand U28573 (N_28573,N_26664,N_26544);
xnor U28574 (N_28574,N_26882,N_26674);
or U28575 (N_28575,N_27191,N_26643);
and U28576 (N_28576,N_26504,N_26985);
or U28577 (N_28577,N_27556,N_27473);
and U28578 (N_28578,N_27555,N_26947);
xor U28579 (N_28579,N_26474,N_27330);
and U28580 (N_28580,N_26525,N_27152);
or U28581 (N_28581,N_26897,N_27222);
nor U28582 (N_28582,N_26568,N_27239);
or U28583 (N_28583,N_26664,N_27260);
and U28584 (N_28584,N_27442,N_26474);
nand U28585 (N_28585,N_27343,N_27339);
or U28586 (N_28586,N_27149,N_26968);
and U28587 (N_28587,N_27122,N_27214);
nor U28588 (N_28588,N_27039,N_26914);
or U28589 (N_28589,N_27093,N_27579);
nor U28590 (N_28590,N_27272,N_27362);
nand U28591 (N_28591,N_27403,N_26556);
nor U28592 (N_28592,N_27475,N_26499);
or U28593 (N_28593,N_26878,N_27261);
xnor U28594 (N_28594,N_26429,N_27512);
or U28595 (N_28595,N_27067,N_27462);
nor U28596 (N_28596,N_27285,N_26580);
xnor U28597 (N_28597,N_26784,N_27289);
and U28598 (N_28598,N_27252,N_26539);
and U28599 (N_28599,N_26836,N_26570);
nand U28600 (N_28600,N_27116,N_26793);
and U28601 (N_28601,N_26601,N_27489);
xnor U28602 (N_28602,N_26418,N_27301);
and U28603 (N_28603,N_26463,N_27432);
or U28604 (N_28604,N_27061,N_26579);
and U28605 (N_28605,N_26901,N_26527);
xnor U28606 (N_28606,N_27223,N_26491);
and U28607 (N_28607,N_26555,N_27251);
nand U28608 (N_28608,N_27507,N_26463);
and U28609 (N_28609,N_27510,N_27524);
nor U28610 (N_28610,N_27571,N_26499);
or U28611 (N_28611,N_26607,N_26680);
or U28612 (N_28612,N_26776,N_27152);
nor U28613 (N_28613,N_27559,N_26527);
and U28614 (N_28614,N_27200,N_27374);
nand U28615 (N_28615,N_26436,N_26622);
nand U28616 (N_28616,N_26413,N_27232);
or U28617 (N_28617,N_27033,N_27567);
xor U28618 (N_28618,N_26464,N_26788);
xor U28619 (N_28619,N_27503,N_26808);
nor U28620 (N_28620,N_27419,N_27143);
nand U28621 (N_28621,N_27205,N_27541);
xnor U28622 (N_28622,N_26945,N_26961);
nor U28623 (N_28623,N_26929,N_27132);
nor U28624 (N_28624,N_26459,N_26550);
nor U28625 (N_28625,N_26883,N_26469);
or U28626 (N_28626,N_26506,N_27261);
and U28627 (N_28627,N_26926,N_27571);
nand U28628 (N_28628,N_26839,N_26465);
xor U28629 (N_28629,N_27459,N_27345);
xor U28630 (N_28630,N_26841,N_26786);
xnor U28631 (N_28631,N_26757,N_26441);
or U28632 (N_28632,N_26569,N_27077);
nor U28633 (N_28633,N_26416,N_26668);
and U28634 (N_28634,N_26441,N_27458);
nand U28635 (N_28635,N_27175,N_27128);
xor U28636 (N_28636,N_27227,N_26782);
xor U28637 (N_28637,N_27561,N_26853);
or U28638 (N_28638,N_27544,N_27126);
or U28639 (N_28639,N_27149,N_27022);
nand U28640 (N_28640,N_26961,N_27150);
nand U28641 (N_28641,N_27418,N_27128);
nor U28642 (N_28642,N_26864,N_27195);
nor U28643 (N_28643,N_26757,N_27227);
xor U28644 (N_28644,N_27479,N_27005);
xor U28645 (N_28645,N_26555,N_27454);
xnor U28646 (N_28646,N_26731,N_27494);
nor U28647 (N_28647,N_27040,N_27564);
nor U28648 (N_28648,N_27016,N_26882);
nor U28649 (N_28649,N_26843,N_26564);
and U28650 (N_28650,N_26494,N_27491);
and U28651 (N_28651,N_27145,N_26772);
and U28652 (N_28652,N_27507,N_26977);
and U28653 (N_28653,N_26541,N_27124);
nor U28654 (N_28654,N_26936,N_26501);
nor U28655 (N_28655,N_27452,N_26582);
nand U28656 (N_28656,N_27176,N_26423);
or U28657 (N_28657,N_26668,N_27014);
nand U28658 (N_28658,N_26656,N_27544);
nor U28659 (N_28659,N_26891,N_27189);
and U28660 (N_28660,N_26834,N_26749);
xnor U28661 (N_28661,N_26627,N_27283);
nand U28662 (N_28662,N_27303,N_27019);
nand U28663 (N_28663,N_27180,N_26890);
and U28664 (N_28664,N_26622,N_26959);
or U28665 (N_28665,N_26917,N_26830);
or U28666 (N_28666,N_27157,N_26662);
and U28667 (N_28667,N_26465,N_27162);
xor U28668 (N_28668,N_26476,N_27260);
nand U28669 (N_28669,N_26588,N_26517);
nand U28670 (N_28670,N_27179,N_27104);
and U28671 (N_28671,N_27220,N_27294);
nor U28672 (N_28672,N_26687,N_27044);
and U28673 (N_28673,N_26607,N_27360);
xor U28674 (N_28674,N_26840,N_26419);
xor U28675 (N_28675,N_26434,N_27058);
and U28676 (N_28676,N_27513,N_27462);
xnor U28677 (N_28677,N_26571,N_27556);
and U28678 (N_28678,N_27256,N_27550);
or U28679 (N_28679,N_26944,N_26633);
or U28680 (N_28680,N_27414,N_27520);
nor U28681 (N_28681,N_27393,N_26917);
xor U28682 (N_28682,N_26711,N_27337);
xnor U28683 (N_28683,N_26880,N_26636);
and U28684 (N_28684,N_26603,N_26988);
or U28685 (N_28685,N_27239,N_26527);
nor U28686 (N_28686,N_26601,N_26719);
nor U28687 (N_28687,N_26439,N_26913);
or U28688 (N_28688,N_27227,N_26475);
and U28689 (N_28689,N_26685,N_26939);
xnor U28690 (N_28690,N_26814,N_26989);
nor U28691 (N_28691,N_26710,N_27590);
xnor U28692 (N_28692,N_27287,N_27487);
or U28693 (N_28693,N_26444,N_27296);
or U28694 (N_28694,N_27266,N_26441);
xnor U28695 (N_28695,N_27219,N_26539);
or U28696 (N_28696,N_26910,N_27459);
xnor U28697 (N_28697,N_26812,N_26564);
nand U28698 (N_28698,N_26591,N_27495);
nand U28699 (N_28699,N_26471,N_27493);
and U28700 (N_28700,N_27270,N_27593);
nand U28701 (N_28701,N_27258,N_27283);
nand U28702 (N_28702,N_26637,N_27290);
nand U28703 (N_28703,N_27171,N_27005);
nand U28704 (N_28704,N_27495,N_27180);
and U28705 (N_28705,N_27403,N_27542);
xnor U28706 (N_28706,N_26462,N_26514);
nand U28707 (N_28707,N_26820,N_26547);
nor U28708 (N_28708,N_27511,N_26596);
and U28709 (N_28709,N_26710,N_27262);
and U28710 (N_28710,N_27297,N_26954);
xnor U28711 (N_28711,N_26676,N_26749);
xor U28712 (N_28712,N_27349,N_26831);
nor U28713 (N_28713,N_27427,N_27123);
nand U28714 (N_28714,N_26892,N_26735);
nand U28715 (N_28715,N_26904,N_26410);
or U28716 (N_28716,N_27344,N_27570);
and U28717 (N_28717,N_26896,N_27342);
nand U28718 (N_28718,N_27168,N_26897);
xnor U28719 (N_28719,N_27553,N_26560);
or U28720 (N_28720,N_26974,N_27448);
xnor U28721 (N_28721,N_26946,N_27237);
nor U28722 (N_28722,N_27417,N_26546);
nor U28723 (N_28723,N_27014,N_26725);
nand U28724 (N_28724,N_26473,N_27077);
nor U28725 (N_28725,N_26890,N_26738);
and U28726 (N_28726,N_27203,N_26948);
and U28727 (N_28727,N_27166,N_26944);
xnor U28728 (N_28728,N_27066,N_27255);
or U28729 (N_28729,N_27081,N_26532);
xnor U28730 (N_28730,N_27093,N_26651);
and U28731 (N_28731,N_26629,N_26928);
and U28732 (N_28732,N_26585,N_26675);
or U28733 (N_28733,N_27527,N_27526);
or U28734 (N_28734,N_26452,N_26866);
nand U28735 (N_28735,N_26608,N_26780);
nor U28736 (N_28736,N_26746,N_27103);
nor U28737 (N_28737,N_27109,N_26437);
nand U28738 (N_28738,N_26738,N_27345);
and U28739 (N_28739,N_27173,N_26931);
nor U28740 (N_28740,N_26716,N_26528);
nand U28741 (N_28741,N_26428,N_27288);
nand U28742 (N_28742,N_27335,N_27393);
xor U28743 (N_28743,N_26509,N_26884);
nor U28744 (N_28744,N_27068,N_27469);
nor U28745 (N_28745,N_27339,N_26472);
nor U28746 (N_28746,N_26755,N_27222);
and U28747 (N_28747,N_26487,N_26874);
xnor U28748 (N_28748,N_26947,N_27112);
xnor U28749 (N_28749,N_27382,N_27395);
xnor U28750 (N_28750,N_27450,N_26757);
or U28751 (N_28751,N_27396,N_27020);
and U28752 (N_28752,N_26825,N_27466);
nor U28753 (N_28753,N_26723,N_26708);
or U28754 (N_28754,N_26830,N_27466);
or U28755 (N_28755,N_27128,N_26623);
xor U28756 (N_28756,N_27315,N_27525);
or U28757 (N_28757,N_27239,N_26622);
or U28758 (N_28758,N_27592,N_27199);
or U28759 (N_28759,N_26662,N_27131);
nand U28760 (N_28760,N_27306,N_26860);
nand U28761 (N_28761,N_26684,N_26730);
xnor U28762 (N_28762,N_26635,N_26890);
xnor U28763 (N_28763,N_26985,N_27110);
or U28764 (N_28764,N_27548,N_26913);
nand U28765 (N_28765,N_26403,N_27145);
nand U28766 (N_28766,N_26791,N_26866);
and U28767 (N_28767,N_27068,N_27464);
nor U28768 (N_28768,N_26494,N_27089);
xor U28769 (N_28769,N_27053,N_27197);
and U28770 (N_28770,N_27177,N_26848);
or U28771 (N_28771,N_27112,N_26693);
and U28772 (N_28772,N_26429,N_27280);
and U28773 (N_28773,N_27333,N_26830);
and U28774 (N_28774,N_27217,N_27515);
nand U28775 (N_28775,N_27592,N_27512);
or U28776 (N_28776,N_26684,N_27230);
xnor U28777 (N_28777,N_27209,N_26505);
and U28778 (N_28778,N_26629,N_27494);
nand U28779 (N_28779,N_26917,N_27008);
nor U28780 (N_28780,N_27378,N_27325);
nor U28781 (N_28781,N_27366,N_26801);
and U28782 (N_28782,N_26455,N_27072);
and U28783 (N_28783,N_26861,N_27346);
or U28784 (N_28784,N_26735,N_26714);
nand U28785 (N_28785,N_26987,N_26521);
or U28786 (N_28786,N_27232,N_26587);
nor U28787 (N_28787,N_27211,N_27108);
xnor U28788 (N_28788,N_26518,N_27490);
xnor U28789 (N_28789,N_26475,N_27197);
nor U28790 (N_28790,N_26681,N_26932);
or U28791 (N_28791,N_27320,N_27125);
xor U28792 (N_28792,N_27555,N_27283);
nor U28793 (N_28793,N_26719,N_27276);
xnor U28794 (N_28794,N_27188,N_26710);
xnor U28795 (N_28795,N_27345,N_27553);
and U28796 (N_28796,N_27212,N_27382);
or U28797 (N_28797,N_27215,N_27002);
or U28798 (N_28798,N_27279,N_27552);
nor U28799 (N_28799,N_26989,N_27201);
xnor U28800 (N_28800,N_27660,N_28393);
or U28801 (N_28801,N_27811,N_28308);
xnor U28802 (N_28802,N_27852,N_28006);
or U28803 (N_28803,N_28727,N_28603);
xor U28804 (N_28804,N_28711,N_28556);
and U28805 (N_28805,N_28516,N_27642);
nor U28806 (N_28806,N_28779,N_27965);
nand U28807 (N_28807,N_28125,N_27862);
nor U28808 (N_28808,N_27768,N_27946);
nor U28809 (N_28809,N_28731,N_27955);
or U28810 (N_28810,N_28139,N_28301);
or U28811 (N_28811,N_28191,N_28661);
and U28812 (N_28812,N_28617,N_27601);
or U28813 (N_28813,N_27614,N_28734);
nor U28814 (N_28814,N_27608,N_28065);
xor U28815 (N_28815,N_28233,N_27915);
xnor U28816 (N_28816,N_28672,N_28657);
or U28817 (N_28817,N_28230,N_27931);
nor U28818 (N_28818,N_27849,N_27712);
or U28819 (N_28819,N_27684,N_28189);
xor U28820 (N_28820,N_28045,N_28532);
or U28821 (N_28821,N_28654,N_28753);
and U28822 (N_28822,N_27855,N_27966);
nand U28823 (N_28823,N_28201,N_28291);
nand U28824 (N_28824,N_28119,N_28051);
nor U28825 (N_28825,N_28417,N_27674);
or U28826 (N_28826,N_27630,N_28548);
or U28827 (N_28827,N_27845,N_28104);
and U28828 (N_28828,N_28165,N_28785);
nand U28829 (N_28829,N_27791,N_27787);
or U28830 (N_28830,N_28101,N_28052);
nand U28831 (N_28831,N_28091,N_28110);
xnor U28832 (N_28832,N_28276,N_28525);
and U28833 (N_28833,N_28684,N_27767);
xor U28834 (N_28834,N_28792,N_28690);
nor U28835 (N_28835,N_27889,N_28437);
nand U28836 (N_28836,N_28044,N_28416);
or U28837 (N_28837,N_27802,N_28318);
xnor U28838 (N_28838,N_28788,N_27603);
and U28839 (N_28839,N_28742,N_28133);
xnor U28840 (N_28840,N_28592,N_28312);
nor U28841 (N_28841,N_27902,N_28306);
nand U28842 (N_28842,N_28762,N_27675);
nor U28843 (N_28843,N_28632,N_28060);
nor U28844 (N_28844,N_27950,N_28665);
nand U28845 (N_28845,N_28170,N_28799);
nor U28846 (N_28846,N_28202,N_27779);
xor U28847 (N_28847,N_28138,N_27774);
or U28848 (N_28848,N_27804,N_28345);
and U28849 (N_28849,N_28273,N_28253);
nand U28850 (N_28850,N_28135,N_28067);
nor U28851 (N_28851,N_28623,N_28611);
nand U28852 (N_28852,N_28396,N_27998);
xor U28853 (N_28853,N_27869,N_28163);
nor U28854 (N_28854,N_28172,N_28012);
nand U28855 (N_28855,N_28086,N_27813);
nand U28856 (N_28856,N_28697,N_28484);
nand U28857 (N_28857,N_28586,N_27692);
nor U28858 (N_28858,N_28224,N_28718);
nand U28859 (N_28859,N_28288,N_28407);
and U28860 (N_28860,N_28517,N_28313);
or U28861 (N_28861,N_27724,N_27663);
nor U28862 (N_28862,N_28177,N_28155);
nor U28863 (N_28863,N_28036,N_28059);
nor U28864 (N_28864,N_28771,N_28058);
xnor U28865 (N_28865,N_28076,N_28499);
or U28866 (N_28866,N_27727,N_28021);
nand U28867 (N_28867,N_28171,N_28325);
nor U28868 (N_28868,N_27857,N_28496);
xor U28869 (N_28869,N_27866,N_27693);
and U28870 (N_28870,N_28609,N_28565);
xor U28871 (N_28871,N_28142,N_28430);
xor U28872 (N_28872,N_28551,N_28440);
nand U28873 (N_28873,N_28703,N_27820);
xnor U28874 (N_28874,N_28315,N_28053);
nand U28875 (N_28875,N_28151,N_28732);
and U28876 (N_28876,N_28213,N_27618);
xor U28877 (N_28877,N_28112,N_27864);
nand U28878 (N_28878,N_28794,N_28098);
nand U28879 (N_28879,N_28714,N_28476);
xnor U28880 (N_28880,N_27858,N_28227);
nand U28881 (N_28881,N_28716,N_28048);
or U28882 (N_28882,N_28722,N_28200);
nor U28883 (N_28883,N_28628,N_28196);
or U28884 (N_28884,N_28512,N_28748);
xor U28885 (N_28885,N_27686,N_27705);
and U28886 (N_28886,N_27985,N_28321);
xor U28887 (N_28887,N_27891,N_27934);
or U28888 (N_28888,N_28751,N_28745);
nor U28889 (N_28889,N_28185,N_28557);
nor U28890 (N_28890,N_28109,N_28298);
or U28891 (N_28891,N_27873,N_27798);
nand U28892 (N_28892,N_28005,N_27745);
nor U28893 (N_28893,N_28515,N_28578);
nand U28894 (N_28894,N_28116,N_27837);
nand U28895 (N_28895,N_27839,N_27664);
nor U28896 (N_28896,N_28131,N_28243);
nand U28897 (N_28897,N_28257,N_27631);
or U28898 (N_28898,N_27942,N_28505);
or U28899 (N_28899,N_28521,N_27754);
or U28900 (N_28900,N_28520,N_28420);
and U28901 (N_28901,N_28130,N_28602);
and U28902 (N_28902,N_28421,N_28775);
and U28903 (N_28903,N_27979,N_28625);
and U28904 (N_28904,N_27817,N_27667);
and U28905 (N_28905,N_28681,N_28134);
xnor U28906 (N_28906,N_27990,N_28295);
xnor U28907 (N_28907,N_28563,N_28282);
nor U28908 (N_28908,N_28409,N_28376);
nand U28909 (N_28909,N_28507,N_27759);
xor U28910 (N_28910,N_28346,N_28490);
xor U28911 (N_28911,N_27823,N_27854);
nor U28912 (N_28912,N_28489,N_27903);
and U28913 (N_28913,N_28141,N_28226);
and U28914 (N_28914,N_28194,N_27808);
nor U28915 (N_28915,N_27919,N_27848);
or U28916 (N_28916,N_27948,N_27769);
or U28917 (N_28917,N_28702,N_27656);
xor U28918 (N_28918,N_28685,N_28148);
nand U28919 (N_28919,N_28175,N_27909);
and U28920 (N_28920,N_28581,N_28766);
and U28921 (N_28921,N_28494,N_28608);
or U28922 (N_28922,N_27790,N_28793);
nand U28923 (N_28923,N_28206,N_27821);
nand U28924 (N_28924,N_28540,N_28388);
nand U28925 (N_28925,N_28310,N_27792);
xor U28926 (N_28926,N_28728,N_28418);
and U28927 (N_28927,N_28103,N_28402);
xnor U28928 (N_28928,N_28468,N_28649);
nand U28929 (N_28929,N_27969,N_28176);
xor U28930 (N_28930,N_28755,N_28300);
xnor U28931 (N_28931,N_27805,N_28047);
nor U28932 (N_28932,N_28641,N_28464);
xor U28933 (N_28933,N_27758,N_28050);
nor U28934 (N_28934,N_28278,N_27868);
or U28935 (N_28935,N_27635,N_27795);
nor U28936 (N_28936,N_28495,N_28616);
nor U28937 (N_28937,N_28397,N_28500);
and U28938 (N_28938,N_28216,N_28349);
and U28939 (N_28939,N_28289,N_27720);
and U28940 (N_28940,N_27905,N_27981);
or U28941 (N_28941,N_28032,N_28725);
nor U28942 (N_28942,N_27937,N_28311);
xor U28943 (N_28943,N_27682,N_28622);
or U28944 (N_28944,N_28089,N_27600);
nand U28945 (N_28945,N_28225,N_28473);
nand U28946 (N_28946,N_28128,N_28046);
xor U28947 (N_28947,N_28744,N_27789);
and U28948 (N_28948,N_28683,N_28283);
nand U28949 (N_28949,N_28575,N_27696);
xnor U28950 (N_28950,N_27606,N_27906);
and U28951 (N_28951,N_28077,N_27812);
nor U28952 (N_28952,N_28763,N_27972);
nor U28953 (N_28953,N_27890,N_28447);
nor U28954 (N_28954,N_28518,N_28092);
or U28955 (N_28955,N_28558,N_27651);
or U28956 (N_28956,N_28704,N_28188);
or U28957 (N_28957,N_28668,N_27835);
and U28958 (N_28958,N_28033,N_27671);
or U28959 (N_28959,N_28250,N_28597);
or U28960 (N_28960,N_28566,N_27910);
or U28961 (N_28961,N_28014,N_28004);
xnor U28962 (N_28962,N_27916,N_27959);
and U28963 (N_28963,N_28377,N_27755);
nand U28964 (N_28964,N_28193,N_27613);
and U28965 (N_28965,N_27681,N_28299);
nand U28966 (N_28966,N_28159,N_28035);
nand U28967 (N_28967,N_27943,N_27741);
and U28968 (N_28968,N_28259,N_27737);
or U28969 (N_28969,N_28061,N_27939);
nand U28970 (N_28970,N_28009,N_28705);
xnor U28971 (N_28971,N_28026,N_27640);
or U28972 (N_28972,N_27929,N_28737);
nor U28973 (N_28973,N_28404,N_28309);
nand U28974 (N_28974,N_27807,N_28750);
and U28975 (N_28975,N_28640,N_28229);
xnor U28976 (N_28976,N_28761,N_28013);
nor U28977 (N_28977,N_28570,N_28419);
or U28978 (N_28978,N_28514,N_27748);
and U28979 (N_28979,N_28270,N_28221);
or U28980 (N_28980,N_28337,N_28441);
nand U28981 (N_28981,N_28504,N_28503);
and U28982 (N_28982,N_27992,N_27715);
nand U28983 (N_28983,N_28352,N_28248);
nor U28984 (N_28984,N_28353,N_28773);
and U28985 (N_28985,N_28712,N_27662);
nor U28986 (N_28986,N_28261,N_28482);
xor U28987 (N_28987,N_28429,N_28215);
nand U28988 (N_28988,N_28660,N_28593);
nor U28989 (N_28989,N_28363,N_27698);
or U28990 (N_28990,N_28756,N_27747);
nor U28991 (N_28991,N_28591,N_28027);
and U28992 (N_28992,N_28509,N_27997);
or U28993 (N_28993,N_27841,N_28583);
nor U28994 (N_28994,N_28576,N_28414);
and U28995 (N_28995,N_28524,N_28222);
nor U28996 (N_28996,N_28327,N_28530);
nor U28997 (N_28997,N_28040,N_27780);
xor U28998 (N_28998,N_27924,N_28568);
nor U28999 (N_28999,N_28721,N_28472);
and U29000 (N_29000,N_28707,N_28427);
or U29001 (N_29001,N_28379,N_27994);
xor U29002 (N_29002,N_27672,N_27734);
xnor U29003 (N_29003,N_28178,N_27914);
xnor U29004 (N_29004,N_27954,N_28203);
and U29005 (N_29005,N_28358,N_28634);
xnor U29006 (N_29006,N_28117,N_27694);
nor U29007 (N_29007,N_28544,N_28535);
nand U29008 (N_29008,N_27801,N_28387);
xor U29009 (N_29009,N_28284,N_28105);
or U29010 (N_29010,N_28372,N_28160);
xor U29011 (N_29011,N_28264,N_28650);
and U29012 (N_29012,N_27649,N_27933);
nand U29013 (N_29013,N_27809,N_28236);
and U29014 (N_29014,N_28220,N_28642);
and U29015 (N_29015,N_28587,N_28635);
nor U29016 (N_29016,N_27898,N_27986);
nand U29017 (N_29017,N_28412,N_28774);
xnor U29018 (N_29018,N_28391,N_27806);
nand U29019 (N_29019,N_28735,N_28644);
nand U29020 (N_29020,N_28256,N_27655);
and U29021 (N_29021,N_28434,N_28477);
nor U29022 (N_29022,N_28538,N_28674);
and U29023 (N_29023,N_27610,N_28231);
or U29024 (N_29024,N_27927,N_27775);
and U29025 (N_29025,N_27704,N_27678);
nand U29026 (N_29026,N_28317,N_27746);
nor U29027 (N_29027,N_27615,N_27657);
xnor U29028 (N_29028,N_28174,N_28340);
or U29029 (N_29029,N_28297,N_28095);
xnor U29030 (N_29030,N_28621,N_28405);
xor U29031 (N_29031,N_27895,N_28513);
and U29032 (N_29032,N_27803,N_27627);
nand U29033 (N_29033,N_28341,N_28150);
nand U29034 (N_29034,N_28457,N_27622);
and U29035 (N_29035,N_28765,N_28329);
and U29036 (N_29036,N_28102,N_28610);
nor U29037 (N_29037,N_27968,N_28688);
nand U29038 (N_29038,N_27743,N_27762);
nand U29039 (N_29039,N_28195,N_28678);
or U29040 (N_29040,N_27900,N_28562);
xnor U29041 (N_29041,N_28533,N_28706);
or U29042 (N_29042,N_27978,N_28480);
and U29043 (N_29043,N_28199,N_27766);
nand U29044 (N_29044,N_27974,N_27763);
nand U29045 (N_29045,N_27607,N_27800);
nor U29046 (N_29046,N_28454,N_28746);
or U29047 (N_29047,N_27647,N_28435);
nor U29048 (N_29048,N_28000,N_28605);
or U29049 (N_29049,N_27888,N_28475);
nor U29050 (N_29050,N_28791,N_27928);
nand U29051 (N_29051,N_28571,N_28439);
and U29052 (N_29052,N_28646,N_27732);
xor U29053 (N_29053,N_28686,N_28274);
nor U29054 (N_29054,N_27717,N_28770);
nand U29055 (N_29055,N_28433,N_27654);
nand U29056 (N_29056,N_28483,N_28554);
and U29057 (N_29057,N_28389,N_27819);
and U29058 (N_29058,N_28332,N_27977);
xor U29059 (N_29059,N_28385,N_28280);
nand U29060 (N_29060,N_27797,N_28212);
nor U29061 (N_29061,N_28010,N_28210);
or U29062 (N_29062,N_28536,N_27865);
nand U29063 (N_29063,N_27625,N_28692);
xnor U29064 (N_29064,N_28423,N_27669);
or U29065 (N_29065,N_27788,N_28754);
nand U29066 (N_29066,N_28463,N_28449);
or U29067 (N_29067,N_28431,N_28508);
xnor U29068 (N_29068,N_28161,N_28720);
and U29069 (N_29069,N_27679,N_28118);
nand U29070 (N_29070,N_28620,N_28790);
or U29071 (N_29071,N_28369,N_28022);
nor U29072 (N_29072,N_27861,N_28739);
nand U29073 (N_29073,N_28375,N_28063);
or U29074 (N_29074,N_28445,N_27999);
nand U29075 (N_29075,N_28265,N_27621);
or U29076 (N_29076,N_27984,N_27646);
or U29077 (N_29077,N_28262,N_28465);
xnor U29078 (N_29078,N_28663,N_27620);
or U29079 (N_29079,N_28460,N_27653);
nand U29080 (N_29080,N_28572,N_28676);
nor U29081 (N_29081,N_27901,N_27751);
and U29082 (N_29082,N_28180,N_27702);
nand U29083 (N_29083,N_28054,N_28157);
nand U29084 (N_29084,N_28542,N_27783);
xor U29085 (N_29085,N_27949,N_28382);
and U29086 (N_29086,N_27636,N_27771);
nand U29087 (N_29087,N_27628,N_28740);
nor U29088 (N_29088,N_28582,N_28687);
and U29089 (N_29089,N_28541,N_28474);
nor U29090 (N_29090,N_28075,N_27668);
nand U29091 (N_29091,N_28614,N_28333);
or U29092 (N_29092,N_28258,N_27982);
nand U29093 (N_29093,N_28549,N_28410);
xnor U29094 (N_29094,N_27918,N_27879);
and U29095 (N_29095,N_27719,N_28787);
nor U29096 (N_29096,N_28316,N_28747);
xor U29097 (N_29097,N_27700,N_27947);
xor U29098 (N_29098,N_28156,N_28240);
and U29099 (N_29099,N_28539,N_28392);
nor U29100 (N_29100,N_28645,N_27665);
xnor U29101 (N_29101,N_28039,N_27673);
nand U29102 (N_29102,N_28028,N_27714);
and U29103 (N_29103,N_28008,N_27639);
nor U29104 (N_29104,N_27683,N_28506);
nor U29105 (N_29105,N_27967,N_28458);
or U29106 (N_29106,N_27709,N_28169);
nor U29107 (N_29107,N_27987,N_28730);
nor U29108 (N_29108,N_28042,N_28637);
xor U29109 (N_29109,N_28015,N_27920);
and U29110 (N_29110,N_28680,N_28374);
and U29111 (N_29111,N_27847,N_27761);
nand U29112 (N_29112,N_27739,N_27650);
nand U29113 (N_29113,N_28145,N_28772);
nor U29114 (N_29114,N_28670,N_28319);
nand U29115 (N_29115,N_28723,N_28481);
and U29116 (N_29116,N_28550,N_28588);
nand U29117 (N_29117,N_28675,N_28064);
or U29118 (N_29118,N_28235,N_27907);
xnor U29119 (N_29119,N_28424,N_28486);
or U29120 (N_29120,N_27963,N_28425);
nor U29121 (N_29121,N_27602,N_27925);
nand U29122 (N_29122,N_28164,N_28677);
and U29123 (N_29123,N_27701,N_28360);
and U29124 (N_29124,N_28294,N_28784);
and U29125 (N_29125,N_28088,N_28600);
nand U29126 (N_29126,N_28371,N_28251);
and U29127 (N_29127,N_28287,N_28669);
nand U29128 (N_29128,N_28709,N_27824);
or U29129 (N_29129,N_27731,N_28777);
nor U29130 (N_29130,N_28038,N_28380);
or U29131 (N_29131,N_28082,N_28384);
xnor U29132 (N_29132,N_27930,N_28573);
and U29133 (N_29133,N_28612,N_27624);
and U29134 (N_29134,N_28488,N_27786);
nor U29135 (N_29135,N_28127,N_28079);
nand U29136 (N_29136,N_28598,N_28303);
xor U29137 (N_29137,N_28383,N_28099);
and U29138 (N_29138,N_27899,N_28403);
or U29139 (N_29139,N_27887,N_27836);
and U29140 (N_29140,N_28795,N_27842);
nor U29141 (N_29141,N_28024,N_28255);
or U29142 (N_29142,N_27884,N_28302);
or U29143 (N_29143,N_28342,N_27964);
nor U29144 (N_29144,N_27749,N_28083);
nand U29145 (N_29145,N_27828,N_28395);
nand U29146 (N_29146,N_28528,N_28204);
and U29147 (N_29147,N_27744,N_28534);
nor U29148 (N_29148,N_28030,N_28643);
nor U29149 (N_29149,N_28461,N_28003);
nand U29150 (N_29150,N_27765,N_28693);
or U29151 (N_29151,N_28594,N_27917);
nor U29152 (N_29152,N_28595,N_28147);
nand U29153 (N_29153,N_28368,N_28252);
nand U29154 (N_29154,N_28606,N_27793);
nor U29155 (N_29155,N_27772,N_27723);
nor U29156 (N_29156,N_27711,N_28334);
and U29157 (N_29157,N_28659,N_28510);
nand U29158 (N_29158,N_28238,N_27680);
or U29159 (N_29159,N_27814,N_28658);
or U29160 (N_29160,N_28219,N_27882);
xor U29161 (N_29161,N_28630,N_27892);
and U29162 (N_29162,N_27750,N_27878);
nor U29163 (N_29163,N_28398,N_27874);
or U29164 (N_29164,N_27796,N_27952);
nand U29165 (N_29165,N_27922,N_28168);
xnor U29166 (N_29166,N_27742,N_27983);
nand U29167 (N_29167,N_27722,N_28268);
nor U29168 (N_29168,N_28760,N_28492);
nand U29169 (N_29169,N_27778,N_28260);
nor U29170 (N_29170,N_27973,N_27638);
or U29171 (N_29171,N_28149,N_27757);
and U29172 (N_29172,N_28113,N_28187);
or U29173 (N_29173,N_28631,N_27752);
or U29174 (N_29174,N_28599,N_28197);
or U29175 (N_29175,N_28162,N_27623);
nand U29176 (N_29176,N_28037,N_28624);
nand U29177 (N_29177,N_28017,N_28502);
and U29178 (N_29178,N_28023,N_27770);
and U29179 (N_29179,N_28713,N_27637);
or U29180 (N_29180,N_27913,N_27735);
nor U29181 (N_29181,N_28069,N_28182);
xor U29182 (N_29182,N_28071,N_28797);
xnor U29183 (N_29183,N_28406,N_27846);
or U29184 (N_29184,N_28184,N_28589);
xnor U29185 (N_29185,N_28639,N_28198);
or U29186 (N_29186,N_28002,N_28186);
and U29187 (N_29187,N_28526,N_28344);
nor U29188 (N_29188,N_28618,N_28081);
nor U29189 (N_29189,N_28537,N_27794);
nand U29190 (N_29190,N_28656,N_28561);
xnor U29191 (N_29191,N_28636,N_27605);
xnor U29192 (N_29192,N_28682,N_27725);
or U29193 (N_29193,N_27825,N_28090);
and U29194 (N_29194,N_28084,N_27644);
nor U29195 (N_29195,N_28529,N_28356);
xor U29196 (N_29196,N_28601,N_27945);
or U29197 (N_29197,N_28776,N_28034);
nor U29198 (N_29198,N_28237,N_27995);
nand U29199 (N_29199,N_27894,N_27877);
nor U29200 (N_29200,N_28320,N_28696);
xnor U29201 (N_29201,N_28132,N_28293);
xnor U29202 (N_29202,N_28339,N_28016);
nor U29203 (N_29203,N_28767,N_27648);
and U29204 (N_29204,N_27944,N_28183);
nand U29205 (N_29205,N_27781,N_28359);
xnor U29206 (N_29206,N_28370,N_28700);
nor U29207 (N_29207,N_28366,N_28667);
nand U29208 (N_29208,N_27687,N_28173);
nand U29209 (N_29209,N_27785,N_27632);
or U29210 (N_29210,N_27911,N_27989);
xor U29211 (N_29211,N_27832,N_28559);
or U29212 (N_29212,N_28121,N_27853);
and U29213 (N_29213,N_28780,N_28126);
nor U29214 (N_29214,N_27867,N_28564);
xnor U29215 (N_29215,N_27726,N_28154);
or U29216 (N_29216,N_28136,N_27926);
and U29217 (N_29217,N_27962,N_28577);
and U29218 (N_29218,N_28627,N_28671);
xor U29219 (N_29219,N_28519,N_27626);
nor U29220 (N_29220,N_28455,N_27896);
and U29221 (N_29221,N_27840,N_27604);
and U29222 (N_29222,N_28580,N_28323);
nor U29223 (N_29223,N_28574,N_27991);
and U29224 (N_29224,N_27729,N_28769);
nor U29225 (N_29225,N_28234,N_27876);
and U29226 (N_29226,N_27830,N_27980);
nor U29227 (N_29227,N_28267,N_28400);
or U29228 (N_29228,N_28655,N_28205);
xor U29229 (N_29229,N_27728,N_28497);
and U29230 (N_29230,N_28350,N_28122);
xor U29231 (N_29231,N_28019,N_28355);
nor U29232 (N_29232,N_27689,N_28638);
xor U29233 (N_29233,N_28426,N_28254);
nor U29234 (N_29234,N_27721,N_28511);
or U29235 (N_29235,N_28401,N_28569);
nor U29236 (N_29236,N_27953,N_27956);
nor U29237 (N_29237,N_28698,N_28242);
nand U29238 (N_29238,N_28487,N_28144);
and U29239 (N_29239,N_28218,N_28552);
or U29240 (N_29240,N_27733,N_27872);
nand U29241 (N_29241,N_28115,N_27643);
and U29242 (N_29242,N_28211,N_28373);
and U29243 (N_29243,N_28691,N_28097);
and U29244 (N_29244,N_27713,N_28448);
nand U29245 (N_29245,N_28555,N_28422);
nor U29246 (N_29246,N_27941,N_27697);
nand U29247 (N_29247,N_27730,N_28247);
nand U29248 (N_29248,N_27756,N_27661);
and U29249 (N_29249,N_28324,N_28719);
nand U29250 (N_29250,N_27976,N_28432);
xnor U29251 (N_29251,N_28633,N_28129);
nand U29252 (N_29252,N_28055,N_27951);
and U29253 (N_29253,N_28778,N_28613);
or U29254 (N_29254,N_27958,N_28666);
and U29255 (N_29255,N_28469,N_27834);
or U29256 (N_29256,N_28604,N_28114);
nor U29257 (N_29257,N_28367,N_28001);
nor U29258 (N_29258,N_28029,N_28100);
nor U29259 (N_29259,N_28152,N_28501);
nand U29260 (N_29260,N_27971,N_28232);
nor U29261 (N_29261,N_28689,N_28647);
xnor U29262 (N_29262,N_28223,N_28362);
and U29263 (N_29263,N_28462,N_28733);
and U29264 (N_29264,N_28347,N_28246);
nand U29265 (N_29265,N_27940,N_28331);
and U29266 (N_29266,N_27863,N_28007);
and U29267 (N_29267,N_27816,N_28607);
nor U29268 (N_29268,N_28498,N_28411);
or U29269 (N_29269,N_28446,N_27760);
or U29270 (N_29270,N_28143,N_28348);
nand U29271 (N_29271,N_28442,N_28543);
or U29272 (N_29272,N_27677,N_27875);
nor U29273 (N_29273,N_28020,N_27908);
xor U29274 (N_29274,N_28438,N_28768);
and U29275 (N_29275,N_27708,N_28459);
nand U29276 (N_29276,N_27753,N_27619);
nand U29277 (N_29277,N_28304,N_28279);
nor U29278 (N_29278,N_27829,N_28615);
and U29279 (N_29279,N_28249,N_28018);
xor U29280 (N_29280,N_27784,N_27961);
nand U29281 (N_29281,N_27690,N_28031);
xor U29282 (N_29282,N_28120,N_28078);
or U29283 (N_29283,N_28579,N_28789);
or U29284 (N_29284,N_28715,N_28073);
or U29285 (N_29285,N_27716,N_27691);
and U29286 (N_29286,N_28286,N_28738);
or U29287 (N_29287,N_28049,N_28123);
and U29288 (N_29288,N_28757,N_28328);
and U29289 (N_29289,N_28781,N_27659);
or U29290 (N_29290,N_27706,N_28783);
nand U29291 (N_29291,N_27764,N_27611);
or U29292 (N_29292,N_27938,N_28652);
nor U29293 (N_29293,N_28585,N_28107);
or U29294 (N_29294,N_28390,N_28093);
and U29295 (N_29295,N_28057,N_28080);
and U29296 (N_29296,N_28108,N_27886);
nand U29297 (N_29297,N_27904,N_28653);
xor U29298 (N_29298,N_27695,N_27871);
and U29299 (N_29299,N_28106,N_28782);
nor U29300 (N_29300,N_28357,N_27883);
nor U29301 (N_29301,N_27707,N_28281);
and U29302 (N_29302,N_28560,N_28749);
xnor U29303 (N_29303,N_27776,N_28664);
xnor U29304 (N_29304,N_28531,N_28330);
nor U29305 (N_29305,N_28269,N_28217);
or U29306 (N_29306,N_27617,N_28285);
nand U29307 (N_29307,N_27676,N_27718);
nor U29308 (N_29308,N_27777,N_28796);
xor U29309 (N_29309,N_27844,N_28399);
nand U29310 (N_29310,N_27641,N_28066);
and U29311 (N_29311,N_27699,N_27799);
xor U29312 (N_29312,N_27935,N_27826);
nor U29313 (N_29313,N_28124,N_27957);
nand U29314 (N_29314,N_28158,N_28451);
nor U29315 (N_29315,N_28786,N_28338);
and U29316 (N_29316,N_28444,N_28011);
or U29317 (N_29317,N_28724,N_28056);
or U29318 (N_29318,N_28190,N_28491);
or U29319 (N_29319,N_28111,N_28179);
or U29320 (N_29320,N_27818,N_28553);
xor U29321 (N_29321,N_27860,N_28074);
or U29322 (N_29322,N_28167,N_27993);
nand U29323 (N_29323,N_28743,N_27893);
xor U29324 (N_29324,N_27634,N_28336);
nand U29325 (N_29325,N_28326,N_28364);
or U29326 (N_29326,N_28322,N_28729);
and U29327 (N_29327,N_27685,N_28701);
xnor U29328 (N_29328,N_28292,N_28381);
xor U29329 (N_29329,N_28343,N_27645);
and U29330 (N_29330,N_27856,N_28296);
or U29331 (N_29331,N_28436,N_28140);
xnor U29332 (N_29332,N_28413,N_28266);
nand U29333 (N_29333,N_27782,N_28798);
nor U29334 (N_29334,N_28694,N_27740);
nand U29335 (N_29335,N_28485,N_28452);
and U29336 (N_29336,N_27859,N_27822);
nor U29337 (N_29337,N_28758,N_27710);
nor U29338 (N_29338,N_28072,N_27936);
or U29339 (N_29339,N_28277,N_28085);
and U29340 (N_29340,N_28428,N_28307);
xnor U29341 (N_29341,N_28087,N_27827);
and U29342 (N_29342,N_27666,N_28567);
xor U29343 (N_29343,N_28096,N_28479);
xor U29344 (N_29344,N_28726,N_27921);
nand U29345 (N_29345,N_28062,N_28041);
xor U29346 (N_29346,N_27996,N_28025);
nor U29347 (N_29347,N_28450,N_28662);
nand U29348 (N_29348,N_28192,N_27897);
and U29349 (N_29349,N_27932,N_28527);
or U29350 (N_29350,N_28094,N_28146);
or U29351 (N_29351,N_27703,N_28522);
nand U29352 (N_29352,N_28228,N_28365);
and U29353 (N_29353,N_28547,N_28619);
xnor U29354 (N_29354,N_27773,N_28679);
xnor U29355 (N_29355,N_27970,N_28245);
nand U29356 (N_29356,N_28351,N_27850);
nor U29357 (N_29357,N_28068,N_28736);
xnor U29358 (N_29358,N_27870,N_28546);
nor U29359 (N_29359,N_28741,N_28523);
nand U29360 (N_29360,N_28290,N_28272);
nand U29361 (N_29361,N_27880,N_28545);
xor U29362 (N_29362,N_28386,N_28478);
nor U29363 (N_29363,N_27616,N_28394);
nor U29364 (N_29364,N_28695,N_27851);
xnor U29365 (N_29365,N_28471,N_27738);
nor U29366 (N_29366,N_28456,N_28470);
nor U29367 (N_29367,N_28415,N_28717);
or U29368 (N_29368,N_28271,N_28263);
and U29369 (N_29369,N_27988,N_28314);
nor U29370 (N_29370,N_28759,N_28626);
nand U29371 (N_29371,N_28239,N_28335);
and U29372 (N_29372,N_28673,N_27960);
and U29373 (N_29373,N_27658,N_27629);
nand U29374 (N_29374,N_28354,N_28207);
or U29375 (N_29375,N_28153,N_28699);
or U29376 (N_29376,N_27815,N_27843);
nand U29377 (N_29377,N_28241,N_28651);
or U29378 (N_29378,N_27736,N_27609);
or U29379 (N_29379,N_27881,N_27612);
nor U29380 (N_29380,N_28590,N_28209);
nor U29381 (N_29381,N_28493,N_27885);
nor U29382 (N_29382,N_27652,N_28181);
or U29383 (N_29383,N_28361,N_28043);
nor U29384 (N_29384,N_27833,N_27975);
and U29385 (N_29385,N_28584,N_27838);
and U29386 (N_29386,N_27670,N_27688);
or U29387 (N_29387,N_28752,N_28467);
or U29388 (N_29388,N_28453,N_28443);
and U29389 (N_29389,N_27633,N_28137);
nor U29390 (N_29390,N_28648,N_27831);
nor U29391 (N_29391,N_28466,N_28275);
nand U29392 (N_29392,N_28305,N_28629);
xnor U29393 (N_29393,N_28244,N_28764);
and U29394 (N_29394,N_28208,N_27810);
and U29395 (N_29395,N_27912,N_28214);
or U29396 (N_29396,N_28708,N_28166);
or U29397 (N_29397,N_28710,N_27923);
or U29398 (N_29398,N_28408,N_28070);
xnor U29399 (N_29399,N_28378,N_28596);
xnor U29400 (N_29400,N_27908,N_27949);
nor U29401 (N_29401,N_27664,N_27845);
nand U29402 (N_29402,N_28778,N_28233);
and U29403 (N_29403,N_28244,N_28618);
and U29404 (N_29404,N_28668,N_28047);
xor U29405 (N_29405,N_27933,N_28730);
and U29406 (N_29406,N_28678,N_27888);
and U29407 (N_29407,N_28615,N_28527);
and U29408 (N_29408,N_28044,N_27990);
nand U29409 (N_29409,N_27999,N_28647);
nor U29410 (N_29410,N_28244,N_28077);
nand U29411 (N_29411,N_28194,N_28303);
nor U29412 (N_29412,N_28084,N_28494);
nor U29413 (N_29413,N_28551,N_28265);
and U29414 (N_29414,N_28447,N_28655);
nor U29415 (N_29415,N_27653,N_27705);
nor U29416 (N_29416,N_28786,N_28541);
or U29417 (N_29417,N_28295,N_28747);
and U29418 (N_29418,N_28442,N_28229);
nand U29419 (N_29419,N_28297,N_28593);
xnor U29420 (N_29420,N_28445,N_27786);
nor U29421 (N_29421,N_28558,N_27956);
or U29422 (N_29422,N_28302,N_28491);
nand U29423 (N_29423,N_27657,N_28514);
nand U29424 (N_29424,N_28397,N_27824);
nor U29425 (N_29425,N_28460,N_28206);
and U29426 (N_29426,N_27776,N_27833);
and U29427 (N_29427,N_28033,N_28151);
nor U29428 (N_29428,N_27944,N_27712);
and U29429 (N_29429,N_28478,N_28313);
or U29430 (N_29430,N_27644,N_28491);
or U29431 (N_29431,N_28355,N_27865);
and U29432 (N_29432,N_27949,N_28679);
xor U29433 (N_29433,N_28232,N_27717);
xor U29434 (N_29434,N_28217,N_28170);
or U29435 (N_29435,N_28466,N_27703);
nand U29436 (N_29436,N_28185,N_28453);
nor U29437 (N_29437,N_27771,N_27991);
and U29438 (N_29438,N_28546,N_28287);
xor U29439 (N_29439,N_28481,N_28484);
xnor U29440 (N_29440,N_28507,N_28315);
and U29441 (N_29441,N_27947,N_27768);
nand U29442 (N_29442,N_28037,N_27761);
nor U29443 (N_29443,N_27887,N_28277);
or U29444 (N_29444,N_28736,N_28677);
nand U29445 (N_29445,N_27843,N_28750);
nand U29446 (N_29446,N_27835,N_28447);
nand U29447 (N_29447,N_28238,N_28526);
and U29448 (N_29448,N_28687,N_28799);
and U29449 (N_29449,N_27738,N_28233);
or U29450 (N_29450,N_27764,N_28419);
nand U29451 (N_29451,N_27674,N_28595);
nand U29452 (N_29452,N_27676,N_28439);
or U29453 (N_29453,N_28066,N_27775);
nor U29454 (N_29454,N_28052,N_27950);
xor U29455 (N_29455,N_28759,N_27678);
nand U29456 (N_29456,N_27840,N_28175);
and U29457 (N_29457,N_28731,N_28681);
xor U29458 (N_29458,N_28394,N_27760);
nor U29459 (N_29459,N_28563,N_28576);
nor U29460 (N_29460,N_28563,N_28470);
nor U29461 (N_29461,N_27916,N_27889);
and U29462 (N_29462,N_27869,N_27919);
nand U29463 (N_29463,N_28516,N_27760);
nor U29464 (N_29464,N_28051,N_27992);
and U29465 (N_29465,N_28536,N_28336);
xnor U29466 (N_29466,N_28041,N_28027);
nor U29467 (N_29467,N_27751,N_27659);
nand U29468 (N_29468,N_27791,N_28137);
nand U29469 (N_29469,N_28499,N_28101);
and U29470 (N_29470,N_28544,N_28086);
and U29471 (N_29471,N_28109,N_28016);
xor U29472 (N_29472,N_27674,N_28098);
xnor U29473 (N_29473,N_27740,N_27737);
nor U29474 (N_29474,N_28694,N_28562);
nand U29475 (N_29475,N_28759,N_28308);
or U29476 (N_29476,N_27645,N_28572);
and U29477 (N_29477,N_28371,N_27620);
and U29478 (N_29478,N_28748,N_28775);
or U29479 (N_29479,N_27813,N_28170);
or U29480 (N_29480,N_28158,N_28251);
xnor U29481 (N_29481,N_28691,N_28604);
nand U29482 (N_29482,N_27801,N_27910);
xor U29483 (N_29483,N_28499,N_28279);
nand U29484 (N_29484,N_28183,N_28466);
nand U29485 (N_29485,N_28001,N_27852);
or U29486 (N_29486,N_28447,N_28716);
and U29487 (N_29487,N_27924,N_27817);
xor U29488 (N_29488,N_28546,N_27713);
nand U29489 (N_29489,N_28390,N_28761);
xor U29490 (N_29490,N_28176,N_27801);
nor U29491 (N_29491,N_27874,N_27927);
or U29492 (N_29492,N_28716,N_28666);
nand U29493 (N_29493,N_27872,N_28432);
nor U29494 (N_29494,N_27774,N_28035);
nor U29495 (N_29495,N_28590,N_28323);
nor U29496 (N_29496,N_28296,N_28232);
xor U29497 (N_29497,N_27665,N_28112);
nand U29498 (N_29498,N_28733,N_27624);
nand U29499 (N_29499,N_28162,N_28099);
and U29500 (N_29500,N_28174,N_28160);
nand U29501 (N_29501,N_27879,N_28384);
or U29502 (N_29502,N_28329,N_28797);
and U29503 (N_29503,N_28627,N_27686);
xor U29504 (N_29504,N_28764,N_28353);
xnor U29505 (N_29505,N_27694,N_28744);
xnor U29506 (N_29506,N_28481,N_28244);
xnor U29507 (N_29507,N_28338,N_28084);
and U29508 (N_29508,N_28395,N_27753);
and U29509 (N_29509,N_27977,N_28421);
xor U29510 (N_29510,N_28634,N_28703);
xor U29511 (N_29511,N_28744,N_27986);
nor U29512 (N_29512,N_27871,N_27916);
xor U29513 (N_29513,N_28624,N_27879);
nand U29514 (N_29514,N_27630,N_27699);
nor U29515 (N_29515,N_28363,N_28098);
or U29516 (N_29516,N_28690,N_28603);
xor U29517 (N_29517,N_28620,N_27748);
xnor U29518 (N_29518,N_28275,N_28024);
or U29519 (N_29519,N_27931,N_27847);
or U29520 (N_29520,N_28066,N_27651);
and U29521 (N_29521,N_28574,N_28792);
xor U29522 (N_29522,N_28366,N_28542);
and U29523 (N_29523,N_28512,N_28509);
or U29524 (N_29524,N_27956,N_28469);
nand U29525 (N_29525,N_27885,N_28186);
or U29526 (N_29526,N_28504,N_28008);
nand U29527 (N_29527,N_28652,N_28710);
or U29528 (N_29528,N_27735,N_28634);
and U29529 (N_29529,N_28281,N_27862);
and U29530 (N_29530,N_28654,N_27710);
or U29531 (N_29531,N_28371,N_28253);
nor U29532 (N_29532,N_28539,N_28306);
xnor U29533 (N_29533,N_28089,N_28008);
nand U29534 (N_29534,N_27910,N_28132);
and U29535 (N_29535,N_27785,N_27740);
or U29536 (N_29536,N_28191,N_28268);
nor U29537 (N_29537,N_28693,N_28304);
nand U29538 (N_29538,N_27935,N_28063);
nor U29539 (N_29539,N_28142,N_27850);
nor U29540 (N_29540,N_28540,N_28312);
or U29541 (N_29541,N_27721,N_27642);
and U29542 (N_29542,N_27953,N_27892);
nor U29543 (N_29543,N_27725,N_27909);
or U29544 (N_29544,N_28346,N_27610);
or U29545 (N_29545,N_28175,N_28186);
and U29546 (N_29546,N_27901,N_27799);
and U29547 (N_29547,N_28687,N_28795);
and U29548 (N_29548,N_28398,N_28195);
nand U29549 (N_29549,N_27988,N_28401);
and U29550 (N_29550,N_28322,N_28562);
xnor U29551 (N_29551,N_27619,N_27860);
and U29552 (N_29552,N_28689,N_28583);
xor U29553 (N_29553,N_27839,N_27729);
xnor U29554 (N_29554,N_27950,N_28027);
or U29555 (N_29555,N_28643,N_28495);
or U29556 (N_29556,N_28573,N_28574);
nor U29557 (N_29557,N_27685,N_28542);
or U29558 (N_29558,N_27968,N_28255);
nand U29559 (N_29559,N_27871,N_27631);
or U29560 (N_29560,N_28275,N_28405);
and U29561 (N_29561,N_28290,N_28297);
nor U29562 (N_29562,N_27740,N_28453);
nand U29563 (N_29563,N_28786,N_28254);
nand U29564 (N_29564,N_28571,N_27760);
and U29565 (N_29565,N_28295,N_28781);
xor U29566 (N_29566,N_28460,N_28694);
nor U29567 (N_29567,N_28418,N_27774);
and U29568 (N_29568,N_28108,N_28483);
xor U29569 (N_29569,N_28258,N_27855);
and U29570 (N_29570,N_28264,N_27641);
nor U29571 (N_29571,N_27631,N_28792);
xor U29572 (N_29572,N_28440,N_28387);
xor U29573 (N_29573,N_28683,N_28066);
nor U29574 (N_29574,N_27915,N_28410);
nor U29575 (N_29575,N_28616,N_28406);
xor U29576 (N_29576,N_27940,N_28180);
xnor U29577 (N_29577,N_28362,N_27757);
nand U29578 (N_29578,N_27901,N_28760);
xor U29579 (N_29579,N_28070,N_28611);
or U29580 (N_29580,N_28259,N_28248);
or U29581 (N_29581,N_28316,N_28287);
xnor U29582 (N_29582,N_27893,N_28643);
xnor U29583 (N_29583,N_28276,N_28182);
nand U29584 (N_29584,N_28249,N_27627);
nand U29585 (N_29585,N_28163,N_28234);
xnor U29586 (N_29586,N_28480,N_27810);
nand U29587 (N_29587,N_28013,N_28219);
nor U29588 (N_29588,N_28522,N_28235);
xnor U29589 (N_29589,N_27821,N_28586);
nand U29590 (N_29590,N_27870,N_27705);
nor U29591 (N_29591,N_28603,N_27662);
nor U29592 (N_29592,N_28534,N_27894);
or U29593 (N_29593,N_28707,N_27666);
xor U29594 (N_29594,N_28336,N_28497);
xor U29595 (N_29595,N_27847,N_28065);
nand U29596 (N_29596,N_28316,N_28145);
xor U29597 (N_29597,N_28799,N_28770);
xnor U29598 (N_29598,N_28240,N_28499);
or U29599 (N_29599,N_28157,N_28166);
xnor U29600 (N_29600,N_27902,N_27711);
xor U29601 (N_29601,N_28692,N_28234);
nor U29602 (N_29602,N_28415,N_27816);
and U29603 (N_29603,N_27979,N_28300);
xor U29604 (N_29604,N_27753,N_27810);
nand U29605 (N_29605,N_28118,N_28348);
or U29606 (N_29606,N_28770,N_27670);
xnor U29607 (N_29607,N_27754,N_28564);
xor U29608 (N_29608,N_27904,N_28591);
and U29609 (N_29609,N_27608,N_27816);
nand U29610 (N_29610,N_28457,N_28631);
nor U29611 (N_29611,N_28577,N_28181);
and U29612 (N_29612,N_27951,N_27609);
xnor U29613 (N_29613,N_27967,N_28798);
nand U29614 (N_29614,N_27956,N_27732);
xor U29615 (N_29615,N_28798,N_28742);
nand U29616 (N_29616,N_28506,N_28052);
nand U29617 (N_29617,N_28115,N_28604);
and U29618 (N_29618,N_27688,N_28728);
or U29619 (N_29619,N_28271,N_28689);
and U29620 (N_29620,N_27662,N_28690);
xor U29621 (N_29621,N_28527,N_28620);
and U29622 (N_29622,N_28009,N_27610);
xor U29623 (N_29623,N_28626,N_28481);
nor U29624 (N_29624,N_28489,N_28203);
and U29625 (N_29625,N_27792,N_27929);
or U29626 (N_29626,N_27614,N_27798);
nand U29627 (N_29627,N_28028,N_28314);
and U29628 (N_29628,N_28052,N_28091);
xor U29629 (N_29629,N_28036,N_28529);
nor U29630 (N_29630,N_28213,N_28128);
or U29631 (N_29631,N_28533,N_28422);
xor U29632 (N_29632,N_28355,N_28539);
xor U29633 (N_29633,N_28038,N_28326);
nand U29634 (N_29634,N_27686,N_28761);
nand U29635 (N_29635,N_27947,N_28714);
nand U29636 (N_29636,N_28585,N_28681);
and U29637 (N_29637,N_27856,N_27666);
and U29638 (N_29638,N_27908,N_27854);
nor U29639 (N_29639,N_27908,N_28198);
and U29640 (N_29640,N_28026,N_28172);
and U29641 (N_29641,N_28130,N_28774);
nand U29642 (N_29642,N_28629,N_28134);
nand U29643 (N_29643,N_28383,N_27719);
nand U29644 (N_29644,N_28535,N_28468);
and U29645 (N_29645,N_27863,N_27900);
nand U29646 (N_29646,N_28076,N_27676);
xor U29647 (N_29647,N_28401,N_28675);
and U29648 (N_29648,N_28245,N_28644);
nand U29649 (N_29649,N_27825,N_28702);
nand U29650 (N_29650,N_28762,N_28183);
xor U29651 (N_29651,N_28450,N_27694);
and U29652 (N_29652,N_28752,N_27847);
nor U29653 (N_29653,N_27852,N_27933);
xnor U29654 (N_29654,N_28150,N_28206);
xnor U29655 (N_29655,N_27708,N_28392);
nand U29656 (N_29656,N_28380,N_27641);
xor U29657 (N_29657,N_27608,N_27714);
or U29658 (N_29658,N_27940,N_28028);
nor U29659 (N_29659,N_28429,N_28483);
and U29660 (N_29660,N_28498,N_28074);
xor U29661 (N_29661,N_27661,N_27819);
nand U29662 (N_29662,N_28360,N_28758);
nor U29663 (N_29663,N_28560,N_28356);
xnor U29664 (N_29664,N_28159,N_28388);
xnor U29665 (N_29665,N_28284,N_28639);
nand U29666 (N_29666,N_28674,N_28515);
nand U29667 (N_29667,N_28315,N_28405);
and U29668 (N_29668,N_28531,N_28275);
and U29669 (N_29669,N_28574,N_27780);
nor U29670 (N_29670,N_27966,N_28489);
nor U29671 (N_29671,N_27810,N_28773);
and U29672 (N_29672,N_28503,N_28306);
nand U29673 (N_29673,N_28253,N_28534);
xor U29674 (N_29674,N_27862,N_27600);
or U29675 (N_29675,N_28006,N_28766);
and U29676 (N_29676,N_27996,N_28054);
or U29677 (N_29677,N_28643,N_28733);
xnor U29678 (N_29678,N_27758,N_28633);
and U29679 (N_29679,N_28503,N_27966);
nand U29680 (N_29680,N_28778,N_28744);
and U29681 (N_29681,N_28549,N_28133);
nand U29682 (N_29682,N_28274,N_28788);
nand U29683 (N_29683,N_28612,N_27644);
nor U29684 (N_29684,N_28314,N_28104);
nor U29685 (N_29685,N_28234,N_28720);
and U29686 (N_29686,N_28455,N_28249);
and U29687 (N_29687,N_27792,N_28142);
nor U29688 (N_29688,N_27800,N_28773);
xor U29689 (N_29689,N_28031,N_28032);
xor U29690 (N_29690,N_27703,N_27871);
xnor U29691 (N_29691,N_28466,N_28545);
and U29692 (N_29692,N_27765,N_28341);
or U29693 (N_29693,N_28366,N_28150);
xnor U29694 (N_29694,N_28576,N_27947);
and U29695 (N_29695,N_28538,N_28109);
nor U29696 (N_29696,N_28308,N_27678);
or U29697 (N_29697,N_28605,N_28068);
xnor U29698 (N_29698,N_28717,N_27849);
nor U29699 (N_29699,N_28100,N_28757);
and U29700 (N_29700,N_28515,N_28207);
nand U29701 (N_29701,N_28320,N_27724);
and U29702 (N_29702,N_28636,N_28350);
or U29703 (N_29703,N_28223,N_28263);
xnor U29704 (N_29704,N_28555,N_27609);
or U29705 (N_29705,N_28384,N_28092);
and U29706 (N_29706,N_28343,N_27759);
nand U29707 (N_29707,N_27917,N_28636);
nand U29708 (N_29708,N_28749,N_28286);
and U29709 (N_29709,N_27972,N_28579);
nor U29710 (N_29710,N_27992,N_28311);
nor U29711 (N_29711,N_27656,N_28360);
and U29712 (N_29712,N_28454,N_27876);
and U29713 (N_29713,N_28044,N_28759);
or U29714 (N_29714,N_27934,N_28625);
nand U29715 (N_29715,N_28325,N_28274);
nor U29716 (N_29716,N_27606,N_28014);
nand U29717 (N_29717,N_28465,N_27927);
nand U29718 (N_29718,N_28280,N_28080);
xnor U29719 (N_29719,N_27874,N_27778);
nand U29720 (N_29720,N_28497,N_27784);
or U29721 (N_29721,N_28527,N_27906);
and U29722 (N_29722,N_27870,N_28377);
xor U29723 (N_29723,N_28019,N_27928);
nand U29724 (N_29724,N_27676,N_27994);
and U29725 (N_29725,N_27714,N_27872);
and U29726 (N_29726,N_27690,N_28010);
and U29727 (N_29727,N_28121,N_28738);
or U29728 (N_29728,N_28718,N_28026);
and U29729 (N_29729,N_28464,N_27945);
nand U29730 (N_29730,N_28659,N_27662);
and U29731 (N_29731,N_28479,N_28011);
nand U29732 (N_29732,N_27857,N_27976);
and U29733 (N_29733,N_27852,N_28270);
nor U29734 (N_29734,N_28406,N_27727);
or U29735 (N_29735,N_28522,N_27655);
xor U29736 (N_29736,N_27692,N_28370);
or U29737 (N_29737,N_28638,N_28676);
nand U29738 (N_29738,N_28229,N_28691);
or U29739 (N_29739,N_28381,N_28678);
nand U29740 (N_29740,N_28234,N_28249);
nand U29741 (N_29741,N_28669,N_28688);
nor U29742 (N_29742,N_28665,N_28062);
xnor U29743 (N_29743,N_28156,N_28116);
and U29744 (N_29744,N_28681,N_28526);
or U29745 (N_29745,N_28655,N_28014);
or U29746 (N_29746,N_27968,N_28592);
xnor U29747 (N_29747,N_28731,N_28652);
nand U29748 (N_29748,N_27946,N_28021);
nor U29749 (N_29749,N_28494,N_28517);
nor U29750 (N_29750,N_28728,N_27852);
nor U29751 (N_29751,N_27930,N_27870);
and U29752 (N_29752,N_28146,N_28717);
and U29753 (N_29753,N_28079,N_28775);
or U29754 (N_29754,N_27704,N_28455);
and U29755 (N_29755,N_28632,N_28448);
and U29756 (N_29756,N_28660,N_28478);
or U29757 (N_29757,N_28627,N_27658);
nor U29758 (N_29758,N_28653,N_28252);
nand U29759 (N_29759,N_27655,N_28730);
and U29760 (N_29760,N_28177,N_28199);
nor U29761 (N_29761,N_28329,N_28469);
nor U29762 (N_29762,N_28778,N_28212);
nor U29763 (N_29763,N_28243,N_28697);
nand U29764 (N_29764,N_27978,N_28792);
and U29765 (N_29765,N_28228,N_28118);
xor U29766 (N_29766,N_28459,N_28249);
nand U29767 (N_29767,N_28796,N_28043);
and U29768 (N_29768,N_27837,N_27907);
nor U29769 (N_29769,N_28461,N_28777);
and U29770 (N_29770,N_27664,N_28517);
or U29771 (N_29771,N_28132,N_28074);
nand U29772 (N_29772,N_27858,N_27890);
and U29773 (N_29773,N_27800,N_28169);
xnor U29774 (N_29774,N_27918,N_28699);
or U29775 (N_29775,N_28636,N_27853);
xor U29776 (N_29776,N_27795,N_28401);
or U29777 (N_29777,N_27659,N_27733);
nand U29778 (N_29778,N_27957,N_28176);
and U29779 (N_29779,N_27965,N_28644);
or U29780 (N_29780,N_28693,N_27921);
nand U29781 (N_29781,N_28017,N_27871);
xnor U29782 (N_29782,N_28233,N_27622);
xnor U29783 (N_29783,N_28700,N_28052);
or U29784 (N_29784,N_27940,N_28761);
xnor U29785 (N_29785,N_28635,N_27673);
nand U29786 (N_29786,N_28008,N_28106);
nor U29787 (N_29787,N_28722,N_28016);
and U29788 (N_29788,N_28747,N_28478);
nand U29789 (N_29789,N_28517,N_28222);
xnor U29790 (N_29790,N_28226,N_28093);
or U29791 (N_29791,N_28237,N_28284);
nand U29792 (N_29792,N_28055,N_28656);
nor U29793 (N_29793,N_28574,N_27921);
nand U29794 (N_29794,N_27702,N_27843);
xnor U29795 (N_29795,N_28442,N_28734);
xor U29796 (N_29796,N_28519,N_27662);
nand U29797 (N_29797,N_28588,N_27967);
xnor U29798 (N_29798,N_27743,N_28012);
nor U29799 (N_29799,N_28510,N_28793);
nor U29800 (N_29800,N_28024,N_27637);
nand U29801 (N_29801,N_28019,N_28569);
and U29802 (N_29802,N_28131,N_28356);
nor U29803 (N_29803,N_27671,N_27854);
nand U29804 (N_29804,N_28343,N_28647);
xor U29805 (N_29805,N_28585,N_28410);
or U29806 (N_29806,N_28333,N_27861);
nand U29807 (N_29807,N_27765,N_28346);
xnor U29808 (N_29808,N_28478,N_28296);
xor U29809 (N_29809,N_28662,N_28143);
nor U29810 (N_29810,N_28029,N_28781);
or U29811 (N_29811,N_28545,N_28098);
or U29812 (N_29812,N_28236,N_27841);
xor U29813 (N_29813,N_28200,N_27728);
nor U29814 (N_29814,N_27600,N_27702);
nand U29815 (N_29815,N_27689,N_28032);
and U29816 (N_29816,N_28168,N_28529);
nand U29817 (N_29817,N_28777,N_28637);
and U29818 (N_29818,N_28337,N_27644);
nand U29819 (N_29819,N_28405,N_28759);
and U29820 (N_29820,N_28624,N_28605);
and U29821 (N_29821,N_27845,N_28543);
nand U29822 (N_29822,N_28715,N_28447);
and U29823 (N_29823,N_28754,N_28228);
nand U29824 (N_29824,N_27775,N_28488);
or U29825 (N_29825,N_28595,N_27886);
xor U29826 (N_29826,N_28007,N_28321);
and U29827 (N_29827,N_28082,N_28228);
and U29828 (N_29828,N_28211,N_28538);
or U29829 (N_29829,N_28436,N_27905);
nor U29830 (N_29830,N_28048,N_28159);
nor U29831 (N_29831,N_27869,N_28440);
and U29832 (N_29832,N_28396,N_27657);
nor U29833 (N_29833,N_28224,N_28664);
and U29834 (N_29834,N_27928,N_28460);
or U29835 (N_29835,N_27798,N_28003);
xor U29836 (N_29836,N_28775,N_28643);
or U29837 (N_29837,N_28648,N_28096);
and U29838 (N_29838,N_27609,N_27630);
and U29839 (N_29839,N_27642,N_28508);
and U29840 (N_29840,N_28482,N_28086);
nor U29841 (N_29841,N_28443,N_28499);
nand U29842 (N_29842,N_27628,N_28556);
and U29843 (N_29843,N_27759,N_27654);
nor U29844 (N_29844,N_27895,N_27791);
nor U29845 (N_29845,N_28047,N_27788);
or U29846 (N_29846,N_28186,N_28286);
nor U29847 (N_29847,N_28117,N_28068);
nand U29848 (N_29848,N_28791,N_28561);
xor U29849 (N_29849,N_28411,N_28432);
and U29850 (N_29850,N_28528,N_28070);
or U29851 (N_29851,N_28041,N_27801);
nand U29852 (N_29852,N_28788,N_28172);
or U29853 (N_29853,N_28708,N_28666);
and U29854 (N_29854,N_28219,N_28572);
or U29855 (N_29855,N_28259,N_27862);
nand U29856 (N_29856,N_27608,N_28396);
or U29857 (N_29857,N_27667,N_28480);
nand U29858 (N_29858,N_28715,N_27858);
nand U29859 (N_29859,N_27956,N_28548);
or U29860 (N_29860,N_27743,N_27927);
xnor U29861 (N_29861,N_27829,N_28043);
nor U29862 (N_29862,N_27813,N_28574);
nor U29863 (N_29863,N_28754,N_27950);
or U29864 (N_29864,N_27912,N_28434);
or U29865 (N_29865,N_28261,N_27948);
nand U29866 (N_29866,N_27754,N_27810);
xor U29867 (N_29867,N_27813,N_27796);
xnor U29868 (N_29868,N_27842,N_28136);
xnor U29869 (N_29869,N_28115,N_28584);
or U29870 (N_29870,N_28407,N_28764);
or U29871 (N_29871,N_27715,N_28082);
or U29872 (N_29872,N_28458,N_28100);
or U29873 (N_29873,N_28405,N_27879);
and U29874 (N_29874,N_27803,N_27960);
and U29875 (N_29875,N_27905,N_28442);
or U29876 (N_29876,N_27692,N_28052);
nor U29877 (N_29877,N_28071,N_27748);
or U29878 (N_29878,N_27979,N_28019);
nand U29879 (N_29879,N_27965,N_28793);
and U29880 (N_29880,N_28608,N_27719);
xnor U29881 (N_29881,N_27933,N_28532);
and U29882 (N_29882,N_27633,N_28534);
nand U29883 (N_29883,N_27996,N_28492);
or U29884 (N_29884,N_28747,N_27979);
xnor U29885 (N_29885,N_27895,N_27986);
xnor U29886 (N_29886,N_27706,N_27925);
nand U29887 (N_29887,N_28108,N_27716);
nand U29888 (N_29888,N_28553,N_27911);
and U29889 (N_29889,N_28497,N_27766);
nor U29890 (N_29890,N_28083,N_27887);
nor U29891 (N_29891,N_28717,N_28437);
nor U29892 (N_29892,N_28730,N_28783);
xnor U29893 (N_29893,N_27848,N_28760);
and U29894 (N_29894,N_28743,N_28467);
and U29895 (N_29895,N_28797,N_27950);
or U29896 (N_29896,N_27893,N_28435);
and U29897 (N_29897,N_28125,N_28770);
and U29898 (N_29898,N_28477,N_27617);
nand U29899 (N_29899,N_28099,N_28593);
and U29900 (N_29900,N_28211,N_28593);
and U29901 (N_29901,N_28670,N_27974);
nand U29902 (N_29902,N_28094,N_28607);
xnor U29903 (N_29903,N_27938,N_27935);
or U29904 (N_29904,N_28582,N_27813);
nand U29905 (N_29905,N_27950,N_28755);
xnor U29906 (N_29906,N_27640,N_28230);
or U29907 (N_29907,N_27968,N_27627);
and U29908 (N_29908,N_28468,N_28100);
nor U29909 (N_29909,N_27788,N_28109);
nor U29910 (N_29910,N_28304,N_28087);
xnor U29911 (N_29911,N_27689,N_27608);
nand U29912 (N_29912,N_27769,N_28694);
nand U29913 (N_29913,N_28247,N_28261);
or U29914 (N_29914,N_28158,N_27809);
nand U29915 (N_29915,N_28775,N_28335);
and U29916 (N_29916,N_28429,N_28239);
nor U29917 (N_29917,N_28273,N_28173);
nor U29918 (N_29918,N_27906,N_28129);
and U29919 (N_29919,N_27959,N_28524);
nand U29920 (N_29920,N_28573,N_28547);
and U29921 (N_29921,N_28695,N_28125);
xor U29922 (N_29922,N_28457,N_28773);
and U29923 (N_29923,N_28507,N_28401);
nand U29924 (N_29924,N_27716,N_28072);
nor U29925 (N_29925,N_28452,N_27656);
nor U29926 (N_29926,N_28273,N_27669);
nor U29927 (N_29927,N_28531,N_28589);
or U29928 (N_29928,N_28156,N_28242);
nor U29929 (N_29929,N_28105,N_28051);
and U29930 (N_29930,N_27905,N_28728);
nand U29931 (N_29931,N_28559,N_27884);
xor U29932 (N_29932,N_28785,N_28128);
xnor U29933 (N_29933,N_27904,N_27753);
nand U29934 (N_29934,N_27762,N_28007);
nor U29935 (N_29935,N_28097,N_28047);
or U29936 (N_29936,N_28104,N_28585);
and U29937 (N_29937,N_28014,N_28780);
nor U29938 (N_29938,N_27656,N_28724);
and U29939 (N_29939,N_28346,N_28760);
nor U29940 (N_29940,N_28498,N_28605);
or U29941 (N_29941,N_28456,N_27869);
nor U29942 (N_29942,N_28460,N_27602);
nor U29943 (N_29943,N_28172,N_28269);
and U29944 (N_29944,N_28118,N_27914);
nand U29945 (N_29945,N_28536,N_28603);
nor U29946 (N_29946,N_27729,N_27889);
or U29947 (N_29947,N_28027,N_28357);
nand U29948 (N_29948,N_28575,N_28522);
nand U29949 (N_29949,N_28001,N_28038);
or U29950 (N_29950,N_28620,N_28255);
and U29951 (N_29951,N_27925,N_27908);
and U29952 (N_29952,N_28048,N_28659);
xnor U29953 (N_29953,N_28574,N_28435);
and U29954 (N_29954,N_27831,N_28212);
nor U29955 (N_29955,N_27737,N_28693);
nand U29956 (N_29956,N_28486,N_27805);
nand U29957 (N_29957,N_28281,N_28226);
xor U29958 (N_29958,N_28513,N_28263);
xnor U29959 (N_29959,N_28527,N_28393);
nand U29960 (N_29960,N_28599,N_28294);
xor U29961 (N_29961,N_28251,N_27937);
nand U29962 (N_29962,N_27802,N_28516);
nor U29963 (N_29963,N_28734,N_27701);
nor U29964 (N_29964,N_27965,N_28623);
nand U29965 (N_29965,N_27603,N_28152);
nand U29966 (N_29966,N_27938,N_27625);
and U29967 (N_29967,N_27800,N_28545);
and U29968 (N_29968,N_28424,N_28422);
xor U29969 (N_29969,N_28064,N_27882);
nand U29970 (N_29970,N_28231,N_28058);
nand U29971 (N_29971,N_28000,N_27855);
xor U29972 (N_29972,N_28620,N_28289);
nand U29973 (N_29973,N_28507,N_28300);
nor U29974 (N_29974,N_27910,N_28308);
nand U29975 (N_29975,N_27608,N_28266);
or U29976 (N_29976,N_28159,N_28090);
and U29977 (N_29977,N_28591,N_27742);
xnor U29978 (N_29978,N_28270,N_28475);
nor U29979 (N_29979,N_28157,N_27743);
or U29980 (N_29980,N_27996,N_28015);
or U29981 (N_29981,N_28108,N_28472);
and U29982 (N_29982,N_27771,N_28445);
nor U29983 (N_29983,N_28603,N_28736);
nor U29984 (N_29984,N_28204,N_28659);
and U29985 (N_29985,N_27910,N_27790);
nand U29986 (N_29986,N_28431,N_27778);
nor U29987 (N_29987,N_27814,N_27887);
nor U29988 (N_29988,N_28797,N_28760);
xnor U29989 (N_29989,N_28429,N_28501);
xor U29990 (N_29990,N_28608,N_28558);
nor U29991 (N_29991,N_28636,N_28628);
nand U29992 (N_29992,N_28726,N_28035);
xnor U29993 (N_29993,N_28461,N_28061);
nor U29994 (N_29994,N_28668,N_28690);
nand U29995 (N_29995,N_28748,N_27860);
and U29996 (N_29996,N_28127,N_27879);
nor U29997 (N_29997,N_28221,N_27900);
nand U29998 (N_29998,N_27711,N_27877);
nor U29999 (N_29999,N_28330,N_28653);
nor UO_0 (O_0,N_29461,N_29601);
xor UO_1 (O_1,N_28962,N_29607);
or UO_2 (O_2,N_29546,N_29274);
or UO_3 (O_3,N_29189,N_28882);
nand UO_4 (O_4,N_29340,N_29393);
or UO_5 (O_5,N_29207,N_28911);
nor UO_6 (O_6,N_29270,N_29375);
or UO_7 (O_7,N_29067,N_29783);
nor UO_8 (O_8,N_28822,N_28832);
or UO_9 (O_9,N_29473,N_29186);
nand UO_10 (O_10,N_29451,N_29438);
xor UO_11 (O_11,N_29527,N_29622);
nand UO_12 (O_12,N_29924,N_29633);
nor UO_13 (O_13,N_29048,N_29082);
xnor UO_14 (O_14,N_29730,N_29807);
xnor UO_15 (O_15,N_29655,N_29430);
or UO_16 (O_16,N_29355,N_28864);
nand UO_17 (O_17,N_29107,N_29420);
nand UO_18 (O_18,N_29839,N_29698);
nor UO_19 (O_19,N_29648,N_28886);
xor UO_20 (O_20,N_29244,N_29614);
xor UO_21 (O_21,N_28859,N_29610);
nand UO_22 (O_22,N_29694,N_29753);
nor UO_23 (O_23,N_29594,N_29298);
xor UO_24 (O_24,N_29021,N_29977);
and UO_25 (O_25,N_29624,N_28936);
and UO_26 (O_26,N_29341,N_29014);
nor UO_27 (O_27,N_29167,N_29154);
or UO_28 (O_28,N_29141,N_29504);
xor UO_29 (O_29,N_28918,N_29321);
and UO_30 (O_30,N_29976,N_29988);
or UO_31 (O_31,N_29351,N_29705);
nand UO_32 (O_32,N_29644,N_28914);
xnor UO_33 (O_33,N_29348,N_28961);
nand UO_34 (O_34,N_29044,N_29866);
and UO_35 (O_35,N_28993,N_29671);
xnor UO_36 (O_36,N_29702,N_29758);
nor UO_37 (O_37,N_29236,N_29523);
nand UO_38 (O_38,N_29040,N_28837);
or UO_39 (O_39,N_29304,N_29996);
xor UO_40 (O_40,N_29492,N_29467);
and UO_41 (O_41,N_29910,N_29446);
and UO_42 (O_42,N_29894,N_29043);
nand UO_43 (O_43,N_29199,N_29934);
xor UO_44 (O_44,N_29445,N_29809);
nand UO_45 (O_45,N_29584,N_29363);
and UO_46 (O_46,N_29469,N_29171);
xnor UO_47 (O_47,N_29872,N_29975);
xor UO_48 (O_48,N_29468,N_29058);
nor UO_49 (O_49,N_29264,N_29091);
xor UO_50 (O_50,N_29819,N_29103);
xor UO_51 (O_51,N_29704,N_29687);
nand UO_52 (O_52,N_29350,N_28897);
nand UO_53 (O_53,N_29087,N_29638);
and UO_54 (O_54,N_29306,N_29050);
and UO_55 (O_55,N_29686,N_29347);
or UO_56 (O_56,N_29431,N_29148);
nand UO_57 (O_57,N_29441,N_29402);
xnor UO_58 (O_58,N_29057,N_29994);
xnor UO_59 (O_59,N_28969,N_29405);
or UO_60 (O_60,N_29273,N_29602);
nand UO_61 (O_61,N_29185,N_29653);
xor UO_62 (O_62,N_29121,N_29053);
xnor UO_63 (O_63,N_28998,N_29582);
nand UO_64 (O_64,N_29125,N_29980);
nand UO_65 (O_65,N_29621,N_29917);
or UO_66 (O_66,N_29826,N_29200);
nor UO_67 (O_67,N_29684,N_29964);
or UO_68 (O_68,N_29209,N_29913);
xnor UO_69 (O_69,N_29104,N_28881);
xnor UO_70 (O_70,N_29381,N_29847);
or UO_71 (O_71,N_28974,N_29318);
xor UO_72 (O_72,N_29890,N_29165);
nand UO_73 (O_73,N_29233,N_29025);
nand UO_74 (O_74,N_29898,N_29069);
and UO_75 (O_75,N_29105,N_29259);
and UO_76 (O_76,N_29282,N_29689);
nand UO_77 (O_77,N_28963,N_29499);
nand UO_78 (O_78,N_29736,N_29322);
nor UO_79 (O_79,N_29314,N_29214);
and UO_80 (O_80,N_29965,N_29804);
xnor UO_81 (O_81,N_29588,N_28863);
and UO_82 (O_82,N_29463,N_29863);
or UO_83 (O_83,N_29423,N_29138);
nor UO_84 (O_84,N_29531,N_28937);
xor UO_85 (O_85,N_29260,N_29170);
and UO_86 (O_86,N_29746,N_29083);
or UO_87 (O_87,N_29706,N_29026);
nor UO_88 (O_88,N_29658,N_29859);
nand UO_89 (O_89,N_29479,N_29424);
nor UO_90 (O_90,N_29845,N_29500);
and UO_91 (O_91,N_29299,N_29568);
nor UO_92 (O_92,N_28844,N_29246);
xor UO_93 (O_93,N_29202,N_29302);
or UO_94 (O_94,N_29751,N_29747);
nand UO_95 (O_95,N_29609,N_29665);
nor UO_96 (O_96,N_29211,N_29824);
and UO_97 (O_97,N_29635,N_29449);
or UO_98 (O_98,N_28867,N_28989);
nor UO_99 (O_99,N_29590,N_29742);
nor UO_100 (O_100,N_29313,N_28893);
and UO_101 (O_101,N_29691,N_29779);
and UO_102 (O_102,N_29963,N_28856);
xnor UO_103 (O_103,N_29902,N_28942);
xor UO_104 (O_104,N_29586,N_29720);
nor UO_105 (O_105,N_28819,N_29992);
nor UO_106 (O_106,N_28924,N_29254);
nor UO_107 (O_107,N_28892,N_29459);
xor UO_108 (O_108,N_29745,N_29339);
nand UO_109 (O_109,N_29549,N_29123);
and UO_110 (O_110,N_29851,N_29275);
nand UO_111 (O_111,N_29943,N_28906);
xor UO_112 (O_112,N_29080,N_29010);
nor UO_113 (O_113,N_29909,N_29835);
nor UO_114 (O_114,N_29404,N_29179);
or UO_115 (O_115,N_29825,N_28919);
nor UO_116 (O_116,N_28866,N_29970);
nand UO_117 (O_117,N_29657,N_29247);
nand UO_118 (O_118,N_28813,N_29364);
or UO_119 (O_119,N_29421,N_29618);
nand UO_120 (O_120,N_29036,N_29817);
xnor UO_121 (O_121,N_29379,N_29544);
xnor UO_122 (O_122,N_28811,N_29256);
nor UO_123 (O_123,N_29249,N_29700);
xnor UO_124 (O_124,N_28869,N_28991);
and UO_125 (O_125,N_28887,N_29112);
or UO_126 (O_126,N_29358,N_29354);
and UO_127 (O_127,N_29785,N_29216);
nor UO_128 (O_128,N_29109,N_29464);
or UO_129 (O_129,N_29137,N_29896);
and UO_130 (O_130,N_29049,N_29713);
nor UO_131 (O_131,N_28908,N_29161);
nor UO_132 (O_132,N_29497,N_29001);
or UO_133 (O_133,N_29636,N_28817);
and UO_134 (O_134,N_29515,N_29243);
nand UO_135 (O_135,N_29195,N_29272);
or UO_136 (O_136,N_29643,N_28909);
and UO_137 (O_137,N_29478,N_29875);
nor UO_138 (O_138,N_29009,N_29511);
and UO_139 (O_139,N_29815,N_28935);
nand UO_140 (O_140,N_28951,N_28996);
and UO_141 (O_141,N_29735,N_29608);
and UO_142 (O_142,N_29984,N_29989);
nand UO_143 (O_143,N_29038,N_29927);
and UO_144 (O_144,N_29072,N_29415);
xor UO_145 (O_145,N_29520,N_29928);
nand UO_146 (O_146,N_29570,N_29793);
or UO_147 (O_147,N_29718,N_29554);
nor UO_148 (O_148,N_29887,N_29501);
nor UO_149 (O_149,N_29990,N_28805);
xor UO_150 (O_150,N_29972,N_29215);
or UO_151 (O_151,N_29953,N_29158);
nand UO_152 (O_152,N_28923,N_29372);
nand UO_153 (O_153,N_28899,N_29032);
nand UO_154 (O_154,N_29222,N_29483);
nor UO_155 (O_155,N_29255,N_29157);
and UO_156 (O_156,N_28857,N_29294);
nand UO_157 (O_157,N_29081,N_29832);
xor UO_158 (O_158,N_29239,N_28843);
xnor UO_159 (O_159,N_29368,N_29485);
or UO_160 (O_160,N_29035,N_28938);
nor UO_161 (O_161,N_29551,N_29432);
or UO_162 (O_162,N_29100,N_29919);
nor UO_163 (O_163,N_29287,N_28978);
and UO_164 (O_164,N_29346,N_29290);
or UO_165 (O_165,N_29181,N_29951);
nor UO_166 (O_166,N_29842,N_29664);
nand UO_167 (O_167,N_29663,N_28928);
and UO_168 (O_168,N_29006,N_29818);
and UO_169 (O_169,N_29987,N_29367);
nand UO_170 (O_170,N_28971,N_28827);
or UO_171 (O_171,N_29721,N_29333);
nand UO_172 (O_172,N_29289,N_28992);
nand UO_173 (O_173,N_28939,N_29914);
nand UO_174 (O_174,N_29978,N_29791);
xor UO_175 (O_175,N_29935,N_29688);
or UO_176 (O_176,N_29886,N_29337);
nand UO_177 (O_177,N_28894,N_29144);
and UO_178 (O_178,N_29061,N_29147);
or UO_179 (O_179,N_29108,N_29427);
nand UO_180 (O_180,N_29525,N_29258);
nand UO_181 (O_181,N_29699,N_28834);
nand UO_182 (O_182,N_28806,N_29595);
or UO_183 (O_183,N_29277,N_29457);
or UO_184 (O_184,N_29417,N_29135);
nor UO_185 (O_185,N_29159,N_28812);
xor UO_186 (O_186,N_29074,N_29649);
and UO_187 (O_187,N_29345,N_29076);
nor UO_188 (O_188,N_29208,N_28841);
xnor UO_189 (O_189,N_29143,N_29606);
nand UO_190 (O_190,N_29654,N_29533);
xor UO_191 (O_191,N_29764,N_29918);
nor UO_192 (O_192,N_29979,N_29521);
or UO_193 (O_193,N_29580,N_29681);
nor UO_194 (O_194,N_29332,N_29997);
or UO_195 (O_195,N_29338,N_29008);
nor UO_196 (O_196,N_29693,N_29106);
nor UO_197 (O_197,N_29781,N_29915);
or UO_198 (O_198,N_28940,N_29117);
or UO_199 (O_199,N_29085,N_29054);
or UO_200 (O_200,N_29670,N_29099);
xor UO_201 (O_201,N_29242,N_29230);
nand UO_202 (O_202,N_29465,N_29903);
nand UO_203 (O_203,N_29548,N_29127);
nor UO_204 (O_204,N_29516,N_29944);
nand UO_205 (O_205,N_29995,N_29470);
nor UO_206 (O_206,N_29399,N_28845);
nand UO_207 (O_207,N_29950,N_29833);
nand UO_208 (O_208,N_29792,N_29068);
and UO_209 (O_209,N_29041,N_29110);
and UO_210 (O_210,N_29675,N_29496);
nor UO_211 (O_211,N_29382,N_29190);
nand UO_212 (O_212,N_29812,N_29855);
nor UO_213 (O_213,N_29889,N_29203);
xor UO_214 (O_214,N_29707,N_29301);
nand UO_215 (O_215,N_29475,N_29572);
nand UO_216 (O_216,N_29336,N_29846);
xnor UO_217 (O_217,N_29952,N_29150);
xor UO_218 (O_218,N_29201,N_28831);
or UO_219 (O_219,N_29407,N_29151);
nand UO_220 (O_220,N_29263,N_29873);
or UO_221 (O_221,N_29276,N_29756);
or UO_222 (O_222,N_28804,N_29947);
nand UO_223 (O_223,N_29071,N_28800);
and UO_224 (O_224,N_29932,N_29122);
or UO_225 (O_225,N_29578,N_29948);
xnor UO_226 (O_226,N_29581,N_28958);
and UO_227 (O_227,N_28945,N_29557);
nand UO_228 (O_228,N_29062,N_28801);
nand UO_229 (O_229,N_28915,N_29899);
and UO_230 (O_230,N_29639,N_29723);
nor UO_231 (O_231,N_29986,N_28952);
nand UO_232 (O_232,N_29860,N_28912);
xnor UO_233 (O_233,N_29234,N_29460);
or UO_234 (O_234,N_29732,N_29380);
nand UO_235 (O_235,N_29271,N_29505);
or UO_236 (O_236,N_29065,N_29840);
nor UO_237 (O_237,N_28855,N_29089);
nor UO_238 (O_238,N_29406,N_29991);
or UO_239 (O_239,N_29774,N_29418);
nor UO_240 (O_240,N_29510,N_28916);
or UO_241 (O_241,N_28946,N_29034);
and UO_242 (O_242,N_29439,N_28848);
xor UO_243 (O_243,N_29891,N_29268);
xnor UO_244 (O_244,N_28877,N_28975);
xnor UO_245 (O_245,N_29882,N_29491);
nand UO_246 (O_246,N_29710,N_29966);
xor UO_247 (O_247,N_29225,N_28926);
or UO_248 (O_248,N_29413,N_29836);
xor UO_249 (O_249,N_28947,N_29019);
and UO_250 (O_250,N_28891,N_29864);
nor UO_251 (O_251,N_28985,N_29365);
nor UO_252 (O_252,N_29949,N_29480);
nand UO_253 (O_253,N_29517,N_29507);
xor UO_254 (O_254,N_29596,N_29772);
and UO_255 (O_255,N_29388,N_29474);
nor UO_256 (O_256,N_29204,N_29174);
xor UO_257 (O_257,N_29395,N_29398);
nand UO_258 (O_258,N_29680,N_29056);
nor UO_259 (O_259,N_29798,N_29617);
xnor UO_260 (O_260,N_28904,N_29788);
nor UO_261 (O_261,N_28970,N_29059);
nand UO_262 (O_262,N_29317,N_29193);
or UO_263 (O_263,N_29003,N_29701);
and UO_264 (O_264,N_29325,N_29018);
or UO_265 (O_265,N_29033,N_29737);
and UO_266 (O_266,N_29132,N_28815);
or UO_267 (O_267,N_28862,N_29900);
nand UO_268 (O_268,N_29397,N_28954);
nand UO_269 (O_269,N_29146,N_28931);
nor UO_270 (O_270,N_29969,N_28976);
and UO_271 (O_271,N_29309,N_29725);
xor UO_272 (O_272,N_29519,N_29955);
or UO_273 (O_273,N_29906,N_29235);
or UO_274 (O_274,N_29786,N_29615);
xor UO_275 (O_275,N_29856,N_29028);
nand UO_276 (O_276,N_28983,N_29489);
or UO_277 (O_277,N_28810,N_29794);
nand UO_278 (O_278,N_28876,N_29187);
nand UO_279 (O_279,N_29210,N_29163);
nand UO_280 (O_280,N_28943,N_29946);
nor UO_281 (O_281,N_29526,N_28825);
nor UO_282 (O_282,N_28956,N_29284);
or UO_283 (O_283,N_29771,N_29153);
nor UO_284 (O_284,N_29974,N_28949);
or UO_285 (O_285,N_28955,N_29802);
xnor UO_286 (O_286,N_29385,N_29757);
xnor UO_287 (O_287,N_29376,N_29861);
and UO_288 (O_288,N_29047,N_29806);
or UO_289 (O_289,N_29542,N_29394);
and UO_290 (O_290,N_29509,N_29567);
xnor UO_291 (O_291,N_29015,N_29327);
xnor UO_292 (O_292,N_29434,N_29871);
nand UO_293 (O_293,N_29066,N_29440);
and UO_294 (O_294,N_29411,N_29005);
nand UO_295 (O_295,N_29717,N_29213);
and UO_296 (O_296,N_29937,N_28987);
or UO_297 (O_297,N_29877,N_29400);
nand UO_298 (O_298,N_29353,N_29403);
and UO_299 (O_299,N_29763,N_29682);
or UO_300 (O_300,N_29620,N_29960);
or UO_301 (O_301,N_29295,N_29878);
or UO_302 (O_302,N_29113,N_28870);
xnor UO_303 (O_303,N_29941,N_29442);
or UO_304 (O_304,N_29448,N_29383);
and UO_305 (O_305,N_29538,N_29184);
and UO_306 (O_306,N_29731,N_29770);
xnor UO_307 (O_307,N_29569,N_29821);
nand UO_308 (O_308,N_29555,N_29940);
nand UO_309 (O_309,N_29754,N_29311);
xor UO_310 (O_310,N_29727,N_29084);
nand UO_311 (O_311,N_29923,N_29556);
nor UO_312 (O_312,N_29343,N_28871);
or UO_313 (O_313,N_29429,N_29734);
xnor UO_314 (O_314,N_29114,N_29092);
and UO_315 (O_315,N_29612,N_29037);
or UO_316 (O_316,N_29422,N_29192);
and UO_317 (O_317,N_29857,N_29384);
and UO_318 (O_318,N_29326,N_28934);
and UO_319 (O_319,N_29098,N_29967);
and UO_320 (O_320,N_29073,N_29623);
or UO_321 (O_321,N_29901,N_29046);
xor UO_322 (O_322,N_29884,N_29176);
and UO_323 (O_323,N_29852,N_29583);
nand UO_324 (O_324,N_29998,N_28860);
nor UO_325 (O_325,N_29627,N_29140);
xor UO_326 (O_326,N_29816,N_29926);
nor UO_327 (O_327,N_29799,N_29733);
nand UO_328 (O_328,N_29933,N_29868);
or UO_329 (O_329,N_29392,N_29945);
and UO_330 (O_330,N_29958,N_29888);
and UO_331 (O_331,N_29739,N_29361);
and UO_332 (O_332,N_29879,N_29116);
and UO_333 (O_333,N_29371,N_29055);
nor UO_334 (O_334,N_29676,N_29016);
nand UO_335 (O_335,N_28953,N_29129);
and UO_336 (O_336,N_29592,N_29444);
or UO_337 (O_337,N_29000,N_29391);
or UO_338 (O_338,N_29064,N_29843);
xnor UO_339 (O_339,N_29637,N_29954);
nand UO_340 (O_340,N_28868,N_29814);
nor UO_341 (O_341,N_29205,N_29063);
or UO_342 (O_342,N_29892,N_28803);
xnor UO_343 (O_343,N_29973,N_29956);
xor UO_344 (O_344,N_29759,N_28972);
nor UO_345 (O_345,N_29029,N_29493);
nand UO_346 (O_346,N_29262,N_29435);
xnor UO_347 (O_347,N_29631,N_29678);
nand UO_348 (O_348,N_29591,N_29983);
nand UO_349 (O_349,N_29052,N_29690);
nor UO_350 (O_350,N_29715,N_29853);
and UO_351 (O_351,N_29450,N_29683);
nand UO_352 (O_352,N_28986,N_29738);
xor UO_353 (O_353,N_29039,N_29942);
xor UO_354 (O_354,N_29456,N_29454);
or UO_355 (O_355,N_29265,N_29514);
nor UO_356 (O_356,N_29959,N_29765);
xor UO_357 (O_357,N_29605,N_28885);
or UO_358 (O_358,N_29227,N_28917);
xor UO_359 (O_359,N_29045,N_29775);
and UO_360 (O_360,N_29708,N_29022);
nand UO_361 (O_361,N_29830,N_29562);
and UO_362 (O_362,N_29288,N_29659);
xor UO_363 (O_363,N_29752,N_29498);
nand UO_364 (O_364,N_29630,N_29593);
and UO_365 (O_365,N_28921,N_29502);
xnor UO_366 (O_366,N_29634,N_29280);
nor UO_367 (O_367,N_29575,N_29805);
nand UO_368 (O_368,N_29982,N_28941);
or UO_369 (O_369,N_29308,N_29436);
xnor UO_370 (O_370,N_29921,N_29640);
nand UO_371 (O_371,N_29503,N_29012);
or UO_372 (O_372,N_28999,N_29585);
or UO_373 (O_373,N_28836,N_29476);
xor UO_374 (O_374,N_29545,N_29632);
or UO_375 (O_375,N_29957,N_28808);
or UO_376 (O_376,N_29820,N_29748);
or UO_377 (O_377,N_28948,N_28950);
or UO_378 (O_378,N_29374,N_29342);
xnor UO_379 (O_379,N_29011,N_29360);
or UO_380 (O_380,N_29539,N_29778);
nand UO_381 (O_381,N_29389,N_29660);
and UO_382 (O_382,N_29724,N_29228);
xnor UO_383 (O_383,N_29145,N_29378);
xor UO_384 (O_384,N_29838,N_29841);
nand UO_385 (O_385,N_29075,N_28842);
nor UO_386 (O_386,N_29194,N_28979);
and UO_387 (O_387,N_28851,N_29283);
xor UO_388 (O_388,N_29261,N_29530);
and UO_389 (O_389,N_29766,N_28984);
or UO_390 (O_390,N_29359,N_29453);
or UO_391 (O_391,N_29813,N_29823);
or UO_392 (O_392,N_28907,N_29716);
and UO_393 (O_393,N_29328,N_29662);
xor UO_394 (O_394,N_29870,N_28895);
nand UO_395 (O_395,N_29668,N_29600);
nand UO_396 (O_396,N_29711,N_29124);
or UO_397 (O_397,N_28990,N_28884);
or UO_398 (O_398,N_29310,N_29552);
nand UO_399 (O_399,N_28966,N_29789);
nand UO_400 (O_400,N_29629,N_29466);
nand UO_401 (O_401,N_29938,N_29795);
xnor UO_402 (O_402,N_28933,N_28875);
nor UO_403 (O_403,N_29490,N_29850);
and UO_404 (O_404,N_29077,N_28820);
and UO_405 (O_405,N_29537,N_29532);
xor UO_406 (O_406,N_28977,N_29096);
or UO_407 (O_407,N_28826,N_29628);
nand UO_408 (O_408,N_29240,N_29981);
nor UO_409 (O_409,N_29414,N_29656);
nand UO_410 (O_410,N_29494,N_28858);
and UO_411 (O_411,N_29168,N_29292);
nand UO_412 (O_412,N_29611,N_29646);
and UO_413 (O_413,N_29241,N_29741);
and UO_414 (O_414,N_29692,N_28925);
nand UO_415 (O_415,N_29579,N_29088);
nor UO_416 (O_416,N_28865,N_29782);
nor UO_417 (O_417,N_29811,N_29709);
xnor UO_418 (O_418,N_28957,N_29251);
nor UO_419 (O_419,N_29437,N_29922);
or UO_420 (O_420,N_29279,N_29156);
and UO_421 (O_421,N_29278,N_28964);
xor UO_422 (O_422,N_29223,N_29729);
nand UO_423 (O_423,N_28967,N_29768);
and UO_424 (O_424,N_29312,N_29094);
xor UO_425 (O_425,N_29316,N_29433);
and UO_426 (O_426,N_29740,N_29206);
nand UO_427 (O_427,N_29196,N_29291);
nand UO_428 (O_428,N_29547,N_29911);
nand UO_429 (O_429,N_28913,N_29408);
nor UO_430 (O_430,N_28901,N_29931);
nor UO_431 (O_431,N_29020,N_29300);
and UO_432 (O_432,N_28905,N_28927);
or UO_433 (O_433,N_29269,N_29577);
and UO_434 (O_434,N_29603,N_28828);
xnor UO_435 (O_435,N_29142,N_29303);
nand UO_436 (O_436,N_28965,N_29673);
xnor UO_437 (O_437,N_29305,N_29182);
nor UO_438 (O_438,N_29559,N_29443);
or UO_439 (O_439,N_28839,N_29095);
xnor UO_440 (O_440,N_29220,N_28854);
and UO_441 (O_441,N_28896,N_29744);
xnor UO_442 (O_442,N_29226,N_29139);
nand UO_443 (O_443,N_29257,N_29626);
and UO_444 (O_444,N_29844,N_29152);
and UO_445 (O_445,N_28821,N_29776);
nand UO_446 (O_446,N_29352,N_29412);
nand UO_447 (O_447,N_29641,N_28988);
nand UO_448 (O_448,N_29344,N_29722);
nor UO_449 (O_449,N_29912,N_29849);
nand UO_450 (O_450,N_29876,N_29248);
or UO_451 (O_451,N_28835,N_29522);
nand UO_452 (O_452,N_29477,N_29541);
or UO_453 (O_453,N_29285,N_28861);
xor UO_454 (O_454,N_29564,N_28902);
nand UO_455 (O_455,N_29281,N_29419);
xor UO_456 (O_456,N_29885,N_28850);
nand UO_457 (O_457,N_29513,N_29128);
or UO_458 (O_458,N_29166,N_29550);
nand UO_459 (O_459,N_29481,N_29221);
or UO_460 (O_460,N_29297,N_29330);
nor UO_461 (O_461,N_29808,N_29097);
or UO_462 (O_462,N_28816,N_29471);
and UO_463 (O_463,N_28829,N_29616);
or UO_464 (O_464,N_29224,N_29452);
or UO_465 (O_465,N_29925,N_29484);
nor UO_466 (O_466,N_29331,N_29004);
and UO_467 (O_467,N_29827,N_29217);
nand UO_468 (O_468,N_29455,N_28824);
or UO_469 (O_469,N_28879,N_28982);
nand UO_470 (O_470,N_29357,N_28910);
nand UO_471 (O_471,N_29023,N_28873);
nor UO_472 (O_472,N_29252,N_29416);
nand UO_473 (O_473,N_29916,N_29130);
or UO_474 (O_474,N_29212,N_29164);
xor UO_475 (O_475,N_29695,N_29535);
xnor UO_476 (O_476,N_29796,N_29131);
and UO_477 (O_477,N_29534,N_29750);
or UO_478 (O_478,N_29232,N_29183);
nand UO_479 (O_479,N_29625,N_28922);
xnor UO_480 (O_480,N_29674,N_29560);
xnor UO_481 (O_481,N_28853,N_29697);
xor UO_482 (O_482,N_28838,N_28823);
or UO_483 (O_483,N_29822,N_29160);
xnor UO_484 (O_484,N_29895,N_29553);
xor UO_485 (O_485,N_29172,N_29854);
nand UO_486 (O_486,N_29120,N_29386);
xnor UO_487 (O_487,N_29324,N_29093);
nand UO_488 (O_488,N_29865,N_29672);
xnor UO_489 (O_489,N_29829,N_29679);
nand UO_490 (O_490,N_29307,N_29362);
xnor UO_491 (O_491,N_28847,N_29652);
nor UO_492 (O_492,N_29651,N_29512);
nand UO_493 (O_493,N_29410,N_29565);
and UO_494 (O_494,N_29862,N_29027);
xnor UO_495 (O_495,N_29013,N_29540);
or UO_496 (O_496,N_29169,N_28883);
nand UO_497 (O_497,N_29198,N_29370);
xnor UO_498 (O_498,N_28809,N_28903);
nor UO_499 (O_499,N_29667,N_29219);
or UO_500 (O_500,N_29366,N_29472);
xnor UO_501 (O_501,N_29831,N_29563);
or UO_502 (O_502,N_29930,N_29323);
and UO_503 (O_503,N_29373,N_29677);
or UO_504 (O_504,N_29936,N_28840);
and UO_505 (O_505,N_29719,N_28814);
and UO_506 (O_506,N_29007,N_29908);
or UO_507 (O_507,N_29377,N_29134);
and UO_508 (O_508,N_29573,N_29286);
nand UO_509 (O_509,N_29175,N_29002);
xnor UO_510 (O_510,N_29396,N_29426);
nand UO_511 (O_511,N_29837,N_29867);
nand UO_512 (O_512,N_29238,N_29115);
nand UO_513 (O_513,N_29961,N_29329);
nand UO_514 (O_514,N_28818,N_29409);
and UO_515 (O_515,N_29571,N_29237);
nand UO_516 (O_516,N_29803,N_29787);
nand UO_517 (O_517,N_29661,N_29760);
or UO_518 (O_518,N_29971,N_29425);
xor UO_519 (O_519,N_28802,N_28973);
nor UO_520 (O_520,N_29587,N_29090);
nand UO_521 (O_521,N_29267,N_28981);
nand UO_522 (O_522,N_28849,N_29149);
nor UO_523 (O_523,N_29762,N_29848);
nor UO_524 (O_524,N_29506,N_29030);
xnor UO_525 (O_525,N_29784,N_29387);
or UO_526 (O_526,N_29874,N_29558);
xnor UO_527 (O_527,N_28997,N_29907);
and UO_528 (O_528,N_29356,N_29599);
xor UO_529 (O_529,N_29266,N_29642);
nand UO_530 (O_530,N_29102,N_29229);
xor UO_531 (O_531,N_29250,N_29647);
xor UO_532 (O_532,N_29810,N_29920);
and UO_533 (O_533,N_29962,N_29773);
nor UO_534 (O_534,N_29666,N_28959);
xnor UO_535 (O_535,N_29458,N_28944);
nor UO_536 (O_536,N_29401,N_29119);
and UO_537 (O_537,N_29335,N_29574);
xnor UO_538 (O_538,N_29650,N_28932);
or UO_539 (O_539,N_28929,N_29968);
nor UO_540 (O_540,N_29893,N_29883);
or UO_541 (O_541,N_28874,N_29619);
xnor UO_542 (O_542,N_29031,N_29999);
xor UO_543 (O_543,N_29696,N_28920);
and UO_544 (O_544,N_29253,N_29334);
nand UO_545 (O_545,N_29767,N_29790);
xnor UO_546 (O_546,N_29155,N_29597);
nor UO_547 (O_547,N_29904,N_29669);
xor UO_548 (O_548,N_29929,N_28888);
xor UO_549 (O_549,N_28995,N_29528);
xor UO_550 (O_550,N_29133,N_29111);
nor UO_551 (O_551,N_28930,N_29869);
xnor UO_552 (O_552,N_29777,N_29749);
xor UO_553 (O_553,N_29118,N_29613);
and UO_554 (O_554,N_29126,N_29780);
and UO_555 (O_555,N_29728,N_29188);
nand UO_556 (O_556,N_28980,N_29180);
or UO_557 (O_557,N_29447,N_29101);
nor UO_558 (O_558,N_29566,N_29881);
and UO_559 (O_559,N_28852,N_29495);
nand UO_560 (O_560,N_29315,N_29518);
or UO_561 (O_561,N_29293,N_29800);
and UO_562 (O_562,N_29743,N_29051);
nand UO_563 (O_563,N_29801,N_28880);
and UO_564 (O_564,N_29858,N_29177);
nand UO_565 (O_565,N_28872,N_29524);
and UO_566 (O_566,N_28807,N_29024);
nor UO_567 (O_567,N_28833,N_28994);
nand UO_568 (O_568,N_29543,N_29017);
xnor UO_569 (O_569,N_29508,N_29761);
and UO_570 (O_570,N_29070,N_29320);
xnor UO_571 (O_571,N_29296,N_29712);
nand UO_572 (O_572,N_29486,N_29218);
nand UO_573 (O_573,N_29589,N_29319);
xnor UO_574 (O_574,N_28890,N_29834);
nor UO_575 (O_575,N_29086,N_28960);
xor UO_576 (O_576,N_29191,N_29231);
nand UO_577 (O_577,N_29797,N_29178);
or UO_578 (O_578,N_29939,N_29245);
nor UO_579 (O_579,N_29078,N_29985);
xnor UO_580 (O_580,N_29487,N_29529);
xor UO_581 (O_581,N_29905,N_29462);
nor UO_582 (O_582,N_29703,N_29536);
and UO_583 (O_583,N_29369,N_29136);
nor UO_584 (O_584,N_29726,N_29197);
nor UO_585 (O_585,N_29576,N_29042);
nand UO_586 (O_586,N_28968,N_29561);
or UO_587 (O_587,N_29993,N_29162);
nand UO_588 (O_588,N_29173,N_28878);
xnor UO_589 (O_589,N_29390,N_29755);
and UO_590 (O_590,N_29598,N_28830);
nor UO_591 (O_591,N_29060,N_29714);
nand UO_592 (O_592,N_29482,N_29604);
nand UO_593 (O_593,N_28900,N_29488);
and UO_594 (O_594,N_29828,N_29769);
or UO_595 (O_595,N_29685,N_29079);
or UO_596 (O_596,N_29645,N_28898);
or UO_597 (O_597,N_29349,N_29897);
nor UO_598 (O_598,N_29428,N_29880);
xnor UO_599 (O_599,N_28889,N_28846);
nor UO_600 (O_600,N_29851,N_29720);
or UO_601 (O_601,N_29689,N_29897);
nand UO_602 (O_602,N_29464,N_29342);
nor UO_603 (O_603,N_29817,N_29191);
and UO_604 (O_604,N_29919,N_29495);
and UO_605 (O_605,N_28922,N_29384);
xnor UO_606 (O_606,N_29931,N_29663);
nor UO_607 (O_607,N_29254,N_29556);
nor UO_608 (O_608,N_29342,N_29527);
and UO_609 (O_609,N_29337,N_29756);
or UO_610 (O_610,N_29388,N_29549);
nor UO_611 (O_611,N_29114,N_29357);
and UO_612 (O_612,N_29793,N_29821);
xor UO_613 (O_613,N_29331,N_29993);
nor UO_614 (O_614,N_29687,N_29706);
nand UO_615 (O_615,N_28936,N_29778);
nor UO_616 (O_616,N_29405,N_29093);
xnor UO_617 (O_617,N_29686,N_29323);
nor UO_618 (O_618,N_29771,N_29652);
nor UO_619 (O_619,N_29468,N_29604);
xor UO_620 (O_620,N_28921,N_29850);
nor UO_621 (O_621,N_28968,N_29949);
and UO_622 (O_622,N_29136,N_28806);
and UO_623 (O_623,N_29382,N_29028);
nor UO_624 (O_624,N_29973,N_28882);
or UO_625 (O_625,N_29864,N_29222);
nor UO_626 (O_626,N_29617,N_29388);
nor UO_627 (O_627,N_29694,N_29603);
nor UO_628 (O_628,N_29025,N_29823);
and UO_629 (O_629,N_28866,N_29102);
nor UO_630 (O_630,N_29704,N_29819);
and UO_631 (O_631,N_29315,N_29862);
and UO_632 (O_632,N_29744,N_29118);
or UO_633 (O_633,N_29381,N_29849);
nor UO_634 (O_634,N_29421,N_29696);
xnor UO_635 (O_635,N_29001,N_29950);
xor UO_636 (O_636,N_28897,N_29857);
xor UO_637 (O_637,N_29682,N_29758);
or UO_638 (O_638,N_29169,N_28977);
and UO_639 (O_639,N_29449,N_29496);
or UO_640 (O_640,N_29464,N_29450);
or UO_641 (O_641,N_29880,N_29054);
xnor UO_642 (O_642,N_29132,N_29393);
nor UO_643 (O_643,N_28966,N_29577);
nand UO_644 (O_644,N_29038,N_29389);
xor UO_645 (O_645,N_29946,N_29537);
nand UO_646 (O_646,N_29454,N_29591);
nand UO_647 (O_647,N_29903,N_29366);
nand UO_648 (O_648,N_29236,N_29814);
or UO_649 (O_649,N_29804,N_28841);
or UO_650 (O_650,N_29914,N_28809);
and UO_651 (O_651,N_29582,N_29449);
xnor UO_652 (O_652,N_29871,N_29429);
nand UO_653 (O_653,N_28888,N_29759);
nand UO_654 (O_654,N_29331,N_29585);
and UO_655 (O_655,N_29015,N_29301);
nand UO_656 (O_656,N_29533,N_29543);
nand UO_657 (O_657,N_29187,N_28909);
xor UO_658 (O_658,N_29826,N_29619);
xnor UO_659 (O_659,N_29317,N_29920);
nor UO_660 (O_660,N_29726,N_29940);
xor UO_661 (O_661,N_29170,N_29449);
and UO_662 (O_662,N_29410,N_29769);
xnor UO_663 (O_663,N_29148,N_28816);
or UO_664 (O_664,N_29479,N_29607);
or UO_665 (O_665,N_29911,N_29607);
or UO_666 (O_666,N_29232,N_29574);
or UO_667 (O_667,N_28885,N_29070);
or UO_668 (O_668,N_29222,N_29523);
and UO_669 (O_669,N_28872,N_29035);
or UO_670 (O_670,N_29940,N_29008);
or UO_671 (O_671,N_29066,N_29775);
nand UO_672 (O_672,N_28816,N_28928);
nor UO_673 (O_673,N_28844,N_29657);
nor UO_674 (O_674,N_28859,N_28972);
nand UO_675 (O_675,N_29578,N_29876);
or UO_676 (O_676,N_29117,N_29411);
nor UO_677 (O_677,N_29635,N_29378);
or UO_678 (O_678,N_29734,N_28990);
nand UO_679 (O_679,N_29604,N_29086);
nor UO_680 (O_680,N_29390,N_29435);
nand UO_681 (O_681,N_29383,N_29262);
or UO_682 (O_682,N_29366,N_29320);
nor UO_683 (O_683,N_29850,N_29776);
nand UO_684 (O_684,N_29952,N_29403);
xnor UO_685 (O_685,N_29754,N_29072);
or UO_686 (O_686,N_29434,N_29990);
and UO_687 (O_687,N_29511,N_29363);
xor UO_688 (O_688,N_29814,N_28847);
or UO_689 (O_689,N_29978,N_29787);
nor UO_690 (O_690,N_29639,N_28993);
xor UO_691 (O_691,N_29703,N_28866);
nor UO_692 (O_692,N_28955,N_29419);
and UO_693 (O_693,N_29421,N_29361);
nand UO_694 (O_694,N_29800,N_29980);
nor UO_695 (O_695,N_29207,N_29506);
nor UO_696 (O_696,N_29938,N_29800);
and UO_697 (O_697,N_29626,N_29460);
and UO_698 (O_698,N_29431,N_29185);
nand UO_699 (O_699,N_29712,N_29255);
or UO_700 (O_700,N_28950,N_28974);
nor UO_701 (O_701,N_28883,N_28895);
or UO_702 (O_702,N_28878,N_29846);
nor UO_703 (O_703,N_29508,N_29341);
xnor UO_704 (O_704,N_28850,N_28942);
nor UO_705 (O_705,N_29888,N_29800);
nor UO_706 (O_706,N_28957,N_29971);
nand UO_707 (O_707,N_29274,N_29944);
and UO_708 (O_708,N_29084,N_28853);
nor UO_709 (O_709,N_29053,N_29113);
nor UO_710 (O_710,N_29472,N_29794);
nor UO_711 (O_711,N_29059,N_29517);
nand UO_712 (O_712,N_29852,N_29076);
nand UO_713 (O_713,N_29832,N_29358);
nor UO_714 (O_714,N_29964,N_29258);
and UO_715 (O_715,N_28833,N_28812);
or UO_716 (O_716,N_29450,N_29713);
nand UO_717 (O_717,N_29124,N_29440);
xor UO_718 (O_718,N_29433,N_29162);
and UO_719 (O_719,N_29789,N_29001);
and UO_720 (O_720,N_29624,N_29710);
and UO_721 (O_721,N_29434,N_29722);
or UO_722 (O_722,N_28960,N_29116);
xor UO_723 (O_723,N_29223,N_29089);
or UO_724 (O_724,N_28946,N_29675);
nand UO_725 (O_725,N_29378,N_29787);
or UO_726 (O_726,N_29100,N_29543);
nor UO_727 (O_727,N_29314,N_29608);
nand UO_728 (O_728,N_29068,N_29870);
nand UO_729 (O_729,N_29612,N_28887);
xnor UO_730 (O_730,N_29961,N_29988);
or UO_731 (O_731,N_29035,N_29853);
or UO_732 (O_732,N_29430,N_29832);
or UO_733 (O_733,N_29944,N_29176);
nand UO_734 (O_734,N_29740,N_29598);
nand UO_735 (O_735,N_28974,N_29811);
or UO_736 (O_736,N_29138,N_29988);
nor UO_737 (O_737,N_28990,N_29341);
or UO_738 (O_738,N_29772,N_29292);
and UO_739 (O_739,N_29242,N_29009);
xnor UO_740 (O_740,N_29317,N_29879);
or UO_741 (O_741,N_28805,N_29404);
and UO_742 (O_742,N_29476,N_29286);
xnor UO_743 (O_743,N_29996,N_28922);
or UO_744 (O_744,N_29337,N_29365);
nor UO_745 (O_745,N_28973,N_28830);
or UO_746 (O_746,N_29941,N_29187);
or UO_747 (O_747,N_29979,N_29234);
nor UO_748 (O_748,N_29261,N_29604);
and UO_749 (O_749,N_29157,N_29108);
nor UO_750 (O_750,N_29169,N_29811);
and UO_751 (O_751,N_28990,N_29222);
nand UO_752 (O_752,N_29923,N_29762);
or UO_753 (O_753,N_29960,N_29148);
or UO_754 (O_754,N_29845,N_29091);
and UO_755 (O_755,N_29963,N_29461);
and UO_756 (O_756,N_29772,N_29817);
nand UO_757 (O_757,N_29334,N_29177);
nor UO_758 (O_758,N_29804,N_29179);
xor UO_759 (O_759,N_29743,N_29612);
nor UO_760 (O_760,N_29129,N_29249);
nor UO_761 (O_761,N_29376,N_29787);
nor UO_762 (O_762,N_28844,N_29619);
nor UO_763 (O_763,N_29613,N_29262);
xnor UO_764 (O_764,N_29287,N_29125);
nand UO_765 (O_765,N_29938,N_29074);
xnor UO_766 (O_766,N_28988,N_29162);
or UO_767 (O_767,N_29830,N_29931);
and UO_768 (O_768,N_28885,N_29177);
nor UO_769 (O_769,N_29716,N_29572);
nor UO_770 (O_770,N_29296,N_29941);
nor UO_771 (O_771,N_29267,N_28899);
nor UO_772 (O_772,N_29307,N_29264);
or UO_773 (O_773,N_28963,N_28938);
nor UO_774 (O_774,N_29226,N_29746);
xor UO_775 (O_775,N_29509,N_29155);
xor UO_776 (O_776,N_29873,N_29282);
and UO_777 (O_777,N_29557,N_29630);
nor UO_778 (O_778,N_29598,N_29899);
nand UO_779 (O_779,N_28902,N_29073);
and UO_780 (O_780,N_29365,N_29606);
nand UO_781 (O_781,N_29886,N_29190);
nand UO_782 (O_782,N_29881,N_28973);
nor UO_783 (O_783,N_29117,N_29401);
or UO_784 (O_784,N_29054,N_29309);
nor UO_785 (O_785,N_29464,N_29690);
or UO_786 (O_786,N_29563,N_29148);
xor UO_787 (O_787,N_29102,N_29777);
nor UO_788 (O_788,N_29108,N_29360);
or UO_789 (O_789,N_29206,N_29234);
or UO_790 (O_790,N_29817,N_29583);
and UO_791 (O_791,N_29921,N_29612);
and UO_792 (O_792,N_29530,N_29727);
xor UO_793 (O_793,N_29959,N_29287);
nand UO_794 (O_794,N_29958,N_29002);
nand UO_795 (O_795,N_29938,N_28877);
or UO_796 (O_796,N_29488,N_29400);
nand UO_797 (O_797,N_29429,N_29218);
nor UO_798 (O_798,N_28896,N_29970);
and UO_799 (O_799,N_29190,N_29556);
and UO_800 (O_800,N_29652,N_29168);
nand UO_801 (O_801,N_28864,N_29591);
nand UO_802 (O_802,N_28806,N_29687);
and UO_803 (O_803,N_28816,N_29606);
xor UO_804 (O_804,N_28976,N_29817);
and UO_805 (O_805,N_29786,N_28811);
or UO_806 (O_806,N_29341,N_29536);
or UO_807 (O_807,N_29296,N_29544);
nor UO_808 (O_808,N_29034,N_29090);
and UO_809 (O_809,N_29326,N_28832);
or UO_810 (O_810,N_29072,N_29627);
and UO_811 (O_811,N_29243,N_29223);
or UO_812 (O_812,N_29385,N_29623);
nor UO_813 (O_813,N_29784,N_29350);
nand UO_814 (O_814,N_29955,N_29724);
and UO_815 (O_815,N_29042,N_29825);
and UO_816 (O_816,N_29758,N_29360);
and UO_817 (O_817,N_29197,N_29880);
nor UO_818 (O_818,N_29658,N_29231);
and UO_819 (O_819,N_29687,N_28910);
nor UO_820 (O_820,N_29654,N_29825);
and UO_821 (O_821,N_29520,N_29916);
nand UO_822 (O_822,N_29390,N_29659);
nor UO_823 (O_823,N_29788,N_29395);
nor UO_824 (O_824,N_29639,N_29349);
and UO_825 (O_825,N_29105,N_29649);
nor UO_826 (O_826,N_28982,N_29241);
or UO_827 (O_827,N_29919,N_29926);
nand UO_828 (O_828,N_28847,N_29976);
xor UO_829 (O_829,N_29077,N_29012);
xor UO_830 (O_830,N_29282,N_28938);
and UO_831 (O_831,N_29598,N_29012);
nand UO_832 (O_832,N_28829,N_29688);
xor UO_833 (O_833,N_29331,N_29606);
and UO_834 (O_834,N_29528,N_29527);
and UO_835 (O_835,N_28975,N_29102);
nor UO_836 (O_836,N_29678,N_29365);
nand UO_837 (O_837,N_29347,N_28985);
and UO_838 (O_838,N_28917,N_28966);
or UO_839 (O_839,N_29863,N_29675);
xnor UO_840 (O_840,N_28921,N_29856);
and UO_841 (O_841,N_29522,N_29651);
nand UO_842 (O_842,N_29482,N_29047);
and UO_843 (O_843,N_29003,N_29686);
or UO_844 (O_844,N_28823,N_29509);
and UO_845 (O_845,N_29173,N_29770);
nor UO_846 (O_846,N_29705,N_28978);
xnor UO_847 (O_847,N_29485,N_29986);
nor UO_848 (O_848,N_29297,N_28997);
nand UO_849 (O_849,N_29908,N_29780);
or UO_850 (O_850,N_29953,N_28960);
nand UO_851 (O_851,N_29035,N_29965);
nor UO_852 (O_852,N_29737,N_29758);
xnor UO_853 (O_853,N_29471,N_29221);
nor UO_854 (O_854,N_29275,N_28969);
xor UO_855 (O_855,N_29325,N_29332);
and UO_856 (O_856,N_29294,N_29958);
xnor UO_857 (O_857,N_29588,N_29172);
or UO_858 (O_858,N_29143,N_29077);
nor UO_859 (O_859,N_29474,N_29717);
nor UO_860 (O_860,N_29964,N_29389);
or UO_861 (O_861,N_29265,N_29947);
and UO_862 (O_862,N_29345,N_29700);
or UO_863 (O_863,N_29150,N_29916);
nor UO_864 (O_864,N_29698,N_29520);
or UO_865 (O_865,N_29408,N_28920);
nand UO_866 (O_866,N_28804,N_29814);
xor UO_867 (O_867,N_29863,N_29805);
nand UO_868 (O_868,N_29995,N_29500);
nor UO_869 (O_869,N_28910,N_28967);
or UO_870 (O_870,N_29022,N_28805);
nand UO_871 (O_871,N_29919,N_29451);
or UO_872 (O_872,N_29999,N_29529);
and UO_873 (O_873,N_29445,N_29797);
nor UO_874 (O_874,N_29456,N_29012);
nand UO_875 (O_875,N_29180,N_29010);
and UO_876 (O_876,N_28942,N_29831);
nand UO_877 (O_877,N_29528,N_29149);
or UO_878 (O_878,N_28940,N_29873);
nor UO_879 (O_879,N_28930,N_28894);
nor UO_880 (O_880,N_29506,N_29487);
and UO_881 (O_881,N_29684,N_29521);
and UO_882 (O_882,N_29954,N_29746);
or UO_883 (O_883,N_29845,N_29251);
nor UO_884 (O_884,N_29914,N_29371);
nor UO_885 (O_885,N_29001,N_29930);
and UO_886 (O_886,N_29410,N_29316);
nand UO_887 (O_887,N_29348,N_29244);
nor UO_888 (O_888,N_29733,N_29176);
nand UO_889 (O_889,N_29504,N_29524);
nand UO_890 (O_890,N_29598,N_29858);
and UO_891 (O_891,N_29259,N_28961);
nor UO_892 (O_892,N_29717,N_29877);
nand UO_893 (O_893,N_29802,N_29109);
and UO_894 (O_894,N_29247,N_28852);
and UO_895 (O_895,N_29484,N_29191);
nand UO_896 (O_896,N_29738,N_28886);
nand UO_897 (O_897,N_29279,N_29582);
and UO_898 (O_898,N_29277,N_29147);
nor UO_899 (O_899,N_29684,N_29298);
xor UO_900 (O_900,N_29791,N_28952);
nand UO_901 (O_901,N_29219,N_29486);
or UO_902 (O_902,N_29027,N_29537);
and UO_903 (O_903,N_28800,N_29302);
or UO_904 (O_904,N_29881,N_29850);
xor UO_905 (O_905,N_29309,N_29221);
and UO_906 (O_906,N_29081,N_29944);
nor UO_907 (O_907,N_28851,N_29371);
and UO_908 (O_908,N_29738,N_29857);
xor UO_909 (O_909,N_29499,N_29123);
or UO_910 (O_910,N_29736,N_29595);
and UO_911 (O_911,N_29133,N_29476);
and UO_912 (O_912,N_29655,N_29064);
xor UO_913 (O_913,N_28895,N_29560);
nor UO_914 (O_914,N_29491,N_29358);
and UO_915 (O_915,N_29448,N_29460);
or UO_916 (O_916,N_29462,N_29142);
xnor UO_917 (O_917,N_28900,N_28967);
xnor UO_918 (O_918,N_29518,N_29076);
and UO_919 (O_919,N_29634,N_29394);
or UO_920 (O_920,N_28942,N_29683);
nand UO_921 (O_921,N_29578,N_29381);
xnor UO_922 (O_922,N_29388,N_29279);
xor UO_923 (O_923,N_29430,N_29987);
nand UO_924 (O_924,N_29902,N_29584);
nor UO_925 (O_925,N_28984,N_29259);
nor UO_926 (O_926,N_29487,N_29186);
nand UO_927 (O_927,N_29205,N_29456);
xor UO_928 (O_928,N_29311,N_29792);
nand UO_929 (O_929,N_28832,N_29256);
or UO_930 (O_930,N_29641,N_29931);
and UO_931 (O_931,N_29994,N_29443);
nand UO_932 (O_932,N_29415,N_29663);
or UO_933 (O_933,N_29930,N_29872);
xnor UO_934 (O_934,N_29961,N_29780);
nand UO_935 (O_935,N_29711,N_29594);
and UO_936 (O_936,N_29256,N_28848);
nor UO_937 (O_937,N_29798,N_29440);
xor UO_938 (O_938,N_29844,N_29551);
xor UO_939 (O_939,N_29083,N_29077);
and UO_940 (O_940,N_28895,N_29125);
xor UO_941 (O_941,N_29968,N_28941);
nand UO_942 (O_942,N_29046,N_29669);
or UO_943 (O_943,N_28948,N_29266);
nand UO_944 (O_944,N_28904,N_28802);
and UO_945 (O_945,N_29325,N_29972);
nor UO_946 (O_946,N_29232,N_29980);
nor UO_947 (O_947,N_29868,N_28858);
xor UO_948 (O_948,N_28825,N_29498);
nand UO_949 (O_949,N_29020,N_29154);
and UO_950 (O_950,N_28950,N_28803);
xnor UO_951 (O_951,N_29081,N_29907);
nor UO_952 (O_952,N_29353,N_28875);
or UO_953 (O_953,N_29760,N_29858);
or UO_954 (O_954,N_29916,N_28998);
or UO_955 (O_955,N_29981,N_29740);
nand UO_956 (O_956,N_29932,N_28884);
nand UO_957 (O_957,N_29034,N_29530);
or UO_958 (O_958,N_28860,N_28907);
nor UO_959 (O_959,N_29658,N_29269);
nand UO_960 (O_960,N_29072,N_29498);
nor UO_961 (O_961,N_29795,N_29835);
nor UO_962 (O_962,N_28916,N_29192);
or UO_963 (O_963,N_29627,N_28999);
nand UO_964 (O_964,N_29622,N_29713);
nand UO_965 (O_965,N_29881,N_29692);
and UO_966 (O_966,N_29570,N_29668);
nor UO_967 (O_967,N_29861,N_29724);
nor UO_968 (O_968,N_29712,N_29853);
and UO_969 (O_969,N_29254,N_29602);
nor UO_970 (O_970,N_28975,N_29249);
and UO_971 (O_971,N_29219,N_29504);
or UO_972 (O_972,N_28887,N_29017);
nand UO_973 (O_973,N_29660,N_29327);
xnor UO_974 (O_974,N_29482,N_29981);
xor UO_975 (O_975,N_29758,N_29450);
xor UO_976 (O_976,N_28930,N_29843);
or UO_977 (O_977,N_29229,N_29203);
and UO_978 (O_978,N_29115,N_29360);
and UO_979 (O_979,N_29335,N_29726);
nor UO_980 (O_980,N_29669,N_29526);
nor UO_981 (O_981,N_28914,N_29934);
xor UO_982 (O_982,N_29605,N_29202);
or UO_983 (O_983,N_29989,N_29226);
xnor UO_984 (O_984,N_29620,N_29856);
and UO_985 (O_985,N_29462,N_29359);
nand UO_986 (O_986,N_29498,N_29517);
nand UO_987 (O_987,N_29705,N_29960);
or UO_988 (O_988,N_29257,N_29777);
and UO_989 (O_989,N_28876,N_28996);
and UO_990 (O_990,N_29047,N_29524);
and UO_991 (O_991,N_29956,N_29721);
nand UO_992 (O_992,N_29696,N_29990);
xnor UO_993 (O_993,N_29218,N_29328);
nand UO_994 (O_994,N_29083,N_29450);
nand UO_995 (O_995,N_28995,N_29168);
xor UO_996 (O_996,N_29403,N_29387);
or UO_997 (O_997,N_29754,N_29025);
and UO_998 (O_998,N_29986,N_28907);
xnor UO_999 (O_999,N_29084,N_28928);
and UO_1000 (O_1000,N_29141,N_29905);
nor UO_1001 (O_1001,N_29458,N_29465);
or UO_1002 (O_1002,N_29767,N_29560);
nand UO_1003 (O_1003,N_28933,N_29987);
nor UO_1004 (O_1004,N_28816,N_29418);
or UO_1005 (O_1005,N_29058,N_29704);
xor UO_1006 (O_1006,N_29183,N_29816);
nor UO_1007 (O_1007,N_29105,N_28843);
nand UO_1008 (O_1008,N_29315,N_29344);
or UO_1009 (O_1009,N_29853,N_29933);
or UO_1010 (O_1010,N_29703,N_29759);
nor UO_1011 (O_1011,N_29478,N_29658);
xnor UO_1012 (O_1012,N_29093,N_29754);
or UO_1013 (O_1013,N_29160,N_29715);
xnor UO_1014 (O_1014,N_29662,N_29205);
and UO_1015 (O_1015,N_29443,N_29317);
nor UO_1016 (O_1016,N_29306,N_29720);
xnor UO_1017 (O_1017,N_29590,N_29376);
and UO_1018 (O_1018,N_29759,N_29398);
nor UO_1019 (O_1019,N_29348,N_28839);
or UO_1020 (O_1020,N_28953,N_29376);
or UO_1021 (O_1021,N_29344,N_28958);
nor UO_1022 (O_1022,N_29739,N_29924);
nand UO_1023 (O_1023,N_29149,N_28926);
and UO_1024 (O_1024,N_28865,N_29436);
nand UO_1025 (O_1025,N_29554,N_29929);
nor UO_1026 (O_1026,N_29992,N_29734);
and UO_1027 (O_1027,N_29892,N_29395);
nand UO_1028 (O_1028,N_29357,N_29626);
nand UO_1029 (O_1029,N_29085,N_29458);
or UO_1030 (O_1030,N_29878,N_29603);
xor UO_1031 (O_1031,N_29747,N_29869);
and UO_1032 (O_1032,N_29964,N_29512);
nand UO_1033 (O_1033,N_29490,N_29784);
nor UO_1034 (O_1034,N_28987,N_29088);
xor UO_1035 (O_1035,N_28931,N_29013);
and UO_1036 (O_1036,N_29473,N_28867);
xnor UO_1037 (O_1037,N_29116,N_28955);
and UO_1038 (O_1038,N_29752,N_29872);
or UO_1039 (O_1039,N_29964,N_29829);
xor UO_1040 (O_1040,N_29758,N_29384);
xnor UO_1041 (O_1041,N_29074,N_29543);
nor UO_1042 (O_1042,N_28924,N_29523);
xor UO_1043 (O_1043,N_29381,N_28898);
and UO_1044 (O_1044,N_29998,N_29105);
and UO_1045 (O_1045,N_29510,N_29564);
nand UO_1046 (O_1046,N_29267,N_29127);
and UO_1047 (O_1047,N_29300,N_29823);
nor UO_1048 (O_1048,N_29491,N_29792);
nand UO_1049 (O_1049,N_29654,N_29065);
or UO_1050 (O_1050,N_29950,N_29059);
nor UO_1051 (O_1051,N_29488,N_29287);
nor UO_1052 (O_1052,N_29197,N_29220);
and UO_1053 (O_1053,N_29822,N_29702);
nand UO_1054 (O_1054,N_29119,N_29404);
xor UO_1055 (O_1055,N_29472,N_29290);
and UO_1056 (O_1056,N_29210,N_29204);
and UO_1057 (O_1057,N_28936,N_29361);
nand UO_1058 (O_1058,N_29163,N_29565);
and UO_1059 (O_1059,N_29460,N_29754);
and UO_1060 (O_1060,N_29851,N_28850);
and UO_1061 (O_1061,N_29150,N_29878);
and UO_1062 (O_1062,N_29410,N_28958);
and UO_1063 (O_1063,N_29704,N_29820);
nand UO_1064 (O_1064,N_29288,N_29898);
and UO_1065 (O_1065,N_29661,N_29879);
nand UO_1066 (O_1066,N_29513,N_29987);
xor UO_1067 (O_1067,N_29041,N_29614);
xor UO_1068 (O_1068,N_29065,N_29018);
nand UO_1069 (O_1069,N_29634,N_29039);
and UO_1070 (O_1070,N_29728,N_29541);
nand UO_1071 (O_1071,N_29499,N_29862);
and UO_1072 (O_1072,N_29400,N_28933);
xnor UO_1073 (O_1073,N_29349,N_29310);
nand UO_1074 (O_1074,N_28917,N_28993);
or UO_1075 (O_1075,N_29909,N_29069);
and UO_1076 (O_1076,N_28994,N_29286);
nor UO_1077 (O_1077,N_29089,N_29463);
and UO_1078 (O_1078,N_29422,N_29521);
nand UO_1079 (O_1079,N_29754,N_29520);
nor UO_1080 (O_1080,N_29643,N_29634);
or UO_1081 (O_1081,N_29129,N_29879);
xor UO_1082 (O_1082,N_28929,N_29480);
or UO_1083 (O_1083,N_29003,N_29640);
or UO_1084 (O_1084,N_28850,N_29271);
nor UO_1085 (O_1085,N_29493,N_29372);
xnor UO_1086 (O_1086,N_29810,N_29012);
nand UO_1087 (O_1087,N_28808,N_29071);
or UO_1088 (O_1088,N_29140,N_29760);
or UO_1089 (O_1089,N_29117,N_28977);
nor UO_1090 (O_1090,N_29796,N_29453);
nor UO_1091 (O_1091,N_29817,N_29591);
nor UO_1092 (O_1092,N_29533,N_29992);
and UO_1093 (O_1093,N_29704,N_29290);
and UO_1094 (O_1094,N_29430,N_29405);
xnor UO_1095 (O_1095,N_29631,N_29375);
and UO_1096 (O_1096,N_28937,N_29829);
xor UO_1097 (O_1097,N_29969,N_29753);
and UO_1098 (O_1098,N_29163,N_29455);
and UO_1099 (O_1099,N_29497,N_29637);
or UO_1100 (O_1100,N_29998,N_29855);
xnor UO_1101 (O_1101,N_28825,N_29496);
nor UO_1102 (O_1102,N_29246,N_29123);
and UO_1103 (O_1103,N_29445,N_29652);
xor UO_1104 (O_1104,N_28863,N_29637);
nor UO_1105 (O_1105,N_29954,N_29639);
or UO_1106 (O_1106,N_29296,N_28988);
xnor UO_1107 (O_1107,N_29461,N_28946);
or UO_1108 (O_1108,N_28877,N_29652);
xor UO_1109 (O_1109,N_29878,N_29521);
and UO_1110 (O_1110,N_28964,N_29754);
and UO_1111 (O_1111,N_29902,N_28844);
nand UO_1112 (O_1112,N_29878,N_29103);
and UO_1113 (O_1113,N_29247,N_29154);
or UO_1114 (O_1114,N_29815,N_29115);
or UO_1115 (O_1115,N_29006,N_29462);
nand UO_1116 (O_1116,N_29874,N_29488);
nand UO_1117 (O_1117,N_28991,N_28870);
or UO_1118 (O_1118,N_28834,N_29343);
nand UO_1119 (O_1119,N_28898,N_28868);
xor UO_1120 (O_1120,N_29891,N_29934);
xnor UO_1121 (O_1121,N_29810,N_29802);
nand UO_1122 (O_1122,N_29061,N_29411);
nor UO_1123 (O_1123,N_29159,N_29729);
or UO_1124 (O_1124,N_28880,N_29861);
or UO_1125 (O_1125,N_29277,N_29630);
nor UO_1126 (O_1126,N_29448,N_29359);
and UO_1127 (O_1127,N_28940,N_29475);
xor UO_1128 (O_1128,N_29417,N_29950);
xnor UO_1129 (O_1129,N_29110,N_29286);
nor UO_1130 (O_1130,N_29606,N_29553);
or UO_1131 (O_1131,N_29106,N_28974);
or UO_1132 (O_1132,N_28924,N_29202);
nor UO_1133 (O_1133,N_29264,N_29399);
and UO_1134 (O_1134,N_28816,N_29572);
nor UO_1135 (O_1135,N_29371,N_29821);
or UO_1136 (O_1136,N_29698,N_29180);
nand UO_1137 (O_1137,N_29803,N_29134);
xnor UO_1138 (O_1138,N_28965,N_29406);
or UO_1139 (O_1139,N_28978,N_29546);
nand UO_1140 (O_1140,N_29711,N_29441);
and UO_1141 (O_1141,N_29158,N_29857);
and UO_1142 (O_1142,N_28982,N_29366);
and UO_1143 (O_1143,N_28884,N_29926);
nand UO_1144 (O_1144,N_29336,N_29448);
nand UO_1145 (O_1145,N_29678,N_29759);
xnor UO_1146 (O_1146,N_29452,N_29102);
and UO_1147 (O_1147,N_29879,N_29585);
nor UO_1148 (O_1148,N_29432,N_28915);
xor UO_1149 (O_1149,N_28954,N_29872);
nor UO_1150 (O_1150,N_29262,N_29962);
nand UO_1151 (O_1151,N_29479,N_29836);
nand UO_1152 (O_1152,N_29882,N_28877);
and UO_1153 (O_1153,N_29124,N_29183);
nand UO_1154 (O_1154,N_28997,N_28855);
nand UO_1155 (O_1155,N_28956,N_29405);
nor UO_1156 (O_1156,N_28916,N_29809);
and UO_1157 (O_1157,N_29342,N_28856);
or UO_1158 (O_1158,N_29803,N_29700);
nor UO_1159 (O_1159,N_29498,N_29618);
and UO_1160 (O_1160,N_29770,N_29782);
xnor UO_1161 (O_1161,N_29884,N_28985);
nor UO_1162 (O_1162,N_29883,N_28806);
or UO_1163 (O_1163,N_29311,N_29712);
nand UO_1164 (O_1164,N_29551,N_28886);
nand UO_1165 (O_1165,N_29219,N_29607);
xnor UO_1166 (O_1166,N_28804,N_28873);
nor UO_1167 (O_1167,N_28974,N_29222);
xnor UO_1168 (O_1168,N_28843,N_29504);
nand UO_1169 (O_1169,N_29125,N_28817);
xnor UO_1170 (O_1170,N_29818,N_29820);
and UO_1171 (O_1171,N_29174,N_29790);
nand UO_1172 (O_1172,N_29249,N_29062);
xnor UO_1173 (O_1173,N_29385,N_29422);
nand UO_1174 (O_1174,N_29209,N_29941);
nor UO_1175 (O_1175,N_29406,N_29146);
nor UO_1176 (O_1176,N_29131,N_28986);
nor UO_1177 (O_1177,N_29485,N_29139);
or UO_1178 (O_1178,N_29088,N_29621);
nand UO_1179 (O_1179,N_29514,N_29402);
xor UO_1180 (O_1180,N_28891,N_28805);
and UO_1181 (O_1181,N_29619,N_29809);
or UO_1182 (O_1182,N_29054,N_29705);
nor UO_1183 (O_1183,N_29755,N_29083);
and UO_1184 (O_1184,N_29215,N_29169);
or UO_1185 (O_1185,N_29670,N_29940);
nand UO_1186 (O_1186,N_29180,N_29920);
or UO_1187 (O_1187,N_28929,N_29198);
or UO_1188 (O_1188,N_29435,N_28845);
nand UO_1189 (O_1189,N_29081,N_29767);
nor UO_1190 (O_1190,N_29854,N_29273);
and UO_1191 (O_1191,N_29887,N_29728);
xnor UO_1192 (O_1192,N_29658,N_29934);
and UO_1193 (O_1193,N_29474,N_29438);
or UO_1194 (O_1194,N_29320,N_29601);
nor UO_1195 (O_1195,N_29755,N_29250);
nor UO_1196 (O_1196,N_29039,N_29514);
and UO_1197 (O_1197,N_29680,N_29023);
xnor UO_1198 (O_1198,N_28970,N_29269);
or UO_1199 (O_1199,N_29541,N_29789);
or UO_1200 (O_1200,N_29708,N_28899);
or UO_1201 (O_1201,N_29403,N_28843);
or UO_1202 (O_1202,N_29343,N_29387);
or UO_1203 (O_1203,N_29549,N_29424);
nor UO_1204 (O_1204,N_29288,N_29913);
and UO_1205 (O_1205,N_29145,N_28907);
or UO_1206 (O_1206,N_29709,N_28944);
nand UO_1207 (O_1207,N_29990,N_29485);
nor UO_1208 (O_1208,N_29241,N_29307);
or UO_1209 (O_1209,N_29571,N_29630);
or UO_1210 (O_1210,N_29689,N_29948);
and UO_1211 (O_1211,N_29595,N_29668);
nor UO_1212 (O_1212,N_29686,N_29688);
or UO_1213 (O_1213,N_28991,N_29458);
xnor UO_1214 (O_1214,N_29473,N_29555);
nand UO_1215 (O_1215,N_29051,N_29053);
nand UO_1216 (O_1216,N_28922,N_29553);
nor UO_1217 (O_1217,N_29891,N_29013);
and UO_1218 (O_1218,N_29748,N_29543);
xor UO_1219 (O_1219,N_29043,N_29726);
nor UO_1220 (O_1220,N_29154,N_28896);
and UO_1221 (O_1221,N_29533,N_29314);
xnor UO_1222 (O_1222,N_29458,N_29464);
or UO_1223 (O_1223,N_29183,N_29585);
or UO_1224 (O_1224,N_29570,N_29872);
nor UO_1225 (O_1225,N_29635,N_29487);
nor UO_1226 (O_1226,N_29394,N_29662);
xnor UO_1227 (O_1227,N_29240,N_29889);
nand UO_1228 (O_1228,N_29058,N_28896);
xor UO_1229 (O_1229,N_29633,N_29640);
or UO_1230 (O_1230,N_29558,N_28969);
and UO_1231 (O_1231,N_29704,N_29538);
and UO_1232 (O_1232,N_29950,N_29703);
or UO_1233 (O_1233,N_29735,N_28847);
xor UO_1234 (O_1234,N_29406,N_29134);
xor UO_1235 (O_1235,N_28956,N_28816);
nand UO_1236 (O_1236,N_29928,N_29978);
and UO_1237 (O_1237,N_29167,N_29968);
or UO_1238 (O_1238,N_29872,N_29465);
nand UO_1239 (O_1239,N_29790,N_29670);
nand UO_1240 (O_1240,N_29205,N_29355);
nor UO_1241 (O_1241,N_28973,N_29302);
and UO_1242 (O_1242,N_29019,N_29573);
or UO_1243 (O_1243,N_29606,N_29683);
or UO_1244 (O_1244,N_29877,N_29588);
or UO_1245 (O_1245,N_28809,N_29164);
xnor UO_1246 (O_1246,N_28954,N_28952);
xor UO_1247 (O_1247,N_29376,N_29607);
or UO_1248 (O_1248,N_29568,N_29015);
xor UO_1249 (O_1249,N_29016,N_29758);
xnor UO_1250 (O_1250,N_29820,N_29796);
and UO_1251 (O_1251,N_28902,N_29923);
nor UO_1252 (O_1252,N_29487,N_29926);
and UO_1253 (O_1253,N_29641,N_29332);
and UO_1254 (O_1254,N_29260,N_28918);
nor UO_1255 (O_1255,N_29933,N_29170);
nand UO_1256 (O_1256,N_28971,N_28825);
or UO_1257 (O_1257,N_29290,N_29660);
nand UO_1258 (O_1258,N_29191,N_29567);
xnor UO_1259 (O_1259,N_29330,N_29504);
xnor UO_1260 (O_1260,N_29091,N_29402);
and UO_1261 (O_1261,N_28894,N_29373);
nor UO_1262 (O_1262,N_29413,N_28856);
and UO_1263 (O_1263,N_29904,N_29487);
nor UO_1264 (O_1264,N_29587,N_29464);
nand UO_1265 (O_1265,N_29237,N_29623);
xor UO_1266 (O_1266,N_29352,N_29999);
nor UO_1267 (O_1267,N_29887,N_29983);
xor UO_1268 (O_1268,N_28954,N_29906);
and UO_1269 (O_1269,N_29975,N_29710);
and UO_1270 (O_1270,N_29918,N_28838);
nor UO_1271 (O_1271,N_29988,N_29624);
xnor UO_1272 (O_1272,N_28861,N_29413);
or UO_1273 (O_1273,N_29375,N_29166);
nor UO_1274 (O_1274,N_28994,N_29205);
xnor UO_1275 (O_1275,N_29786,N_29402);
xnor UO_1276 (O_1276,N_29615,N_29071);
nand UO_1277 (O_1277,N_29217,N_28851);
xor UO_1278 (O_1278,N_29820,N_29129);
nor UO_1279 (O_1279,N_29560,N_29410);
or UO_1280 (O_1280,N_29182,N_29829);
xor UO_1281 (O_1281,N_29079,N_29935);
nor UO_1282 (O_1282,N_28859,N_29179);
nand UO_1283 (O_1283,N_28816,N_29738);
nand UO_1284 (O_1284,N_29570,N_28899);
nand UO_1285 (O_1285,N_29093,N_29111);
xor UO_1286 (O_1286,N_29866,N_29939);
nand UO_1287 (O_1287,N_29124,N_29145);
xnor UO_1288 (O_1288,N_28909,N_29608);
nor UO_1289 (O_1289,N_29593,N_29847);
xnor UO_1290 (O_1290,N_29923,N_28894);
or UO_1291 (O_1291,N_29763,N_29610);
nor UO_1292 (O_1292,N_28840,N_28849);
and UO_1293 (O_1293,N_29490,N_29170);
nor UO_1294 (O_1294,N_29512,N_29994);
and UO_1295 (O_1295,N_29515,N_29724);
nand UO_1296 (O_1296,N_28845,N_29343);
nor UO_1297 (O_1297,N_29823,N_29227);
or UO_1298 (O_1298,N_29900,N_29040);
xor UO_1299 (O_1299,N_29857,N_29695);
or UO_1300 (O_1300,N_29870,N_29192);
xor UO_1301 (O_1301,N_29006,N_29260);
nand UO_1302 (O_1302,N_29085,N_29489);
and UO_1303 (O_1303,N_29092,N_29526);
and UO_1304 (O_1304,N_28826,N_28864);
nor UO_1305 (O_1305,N_29826,N_29274);
xor UO_1306 (O_1306,N_29218,N_29017);
or UO_1307 (O_1307,N_29548,N_28940);
xor UO_1308 (O_1308,N_29695,N_29982);
or UO_1309 (O_1309,N_29269,N_29901);
nand UO_1310 (O_1310,N_29171,N_29211);
xor UO_1311 (O_1311,N_29798,N_29148);
xor UO_1312 (O_1312,N_29576,N_29144);
xor UO_1313 (O_1313,N_29375,N_29900);
or UO_1314 (O_1314,N_28994,N_28965);
nor UO_1315 (O_1315,N_29219,N_29027);
or UO_1316 (O_1316,N_29322,N_28993);
or UO_1317 (O_1317,N_29550,N_29670);
and UO_1318 (O_1318,N_28982,N_29230);
xnor UO_1319 (O_1319,N_28974,N_29559);
or UO_1320 (O_1320,N_29087,N_29222);
and UO_1321 (O_1321,N_29351,N_29119);
and UO_1322 (O_1322,N_29369,N_29289);
nor UO_1323 (O_1323,N_29486,N_29973);
nor UO_1324 (O_1324,N_29751,N_29191);
or UO_1325 (O_1325,N_28919,N_29938);
xnor UO_1326 (O_1326,N_29144,N_29890);
nor UO_1327 (O_1327,N_29959,N_29182);
nor UO_1328 (O_1328,N_29894,N_29224);
or UO_1329 (O_1329,N_29188,N_29534);
nand UO_1330 (O_1330,N_29397,N_29957);
and UO_1331 (O_1331,N_29902,N_29534);
or UO_1332 (O_1332,N_29954,N_28847);
xor UO_1333 (O_1333,N_29637,N_28990);
and UO_1334 (O_1334,N_28985,N_29402);
nor UO_1335 (O_1335,N_29900,N_29839);
or UO_1336 (O_1336,N_28973,N_29501);
nand UO_1337 (O_1337,N_29612,N_28801);
and UO_1338 (O_1338,N_29300,N_29770);
xor UO_1339 (O_1339,N_29772,N_29069);
or UO_1340 (O_1340,N_29025,N_29399);
nor UO_1341 (O_1341,N_29904,N_29302);
nand UO_1342 (O_1342,N_29542,N_29872);
nand UO_1343 (O_1343,N_29833,N_28982);
xor UO_1344 (O_1344,N_28896,N_29924);
or UO_1345 (O_1345,N_29427,N_29551);
and UO_1346 (O_1346,N_29073,N_29933);
nand UO_1347 (O_1347,N_29541,N_29715);
nand UO_1348 (O_1348,N_29075,N_28991);
and UO_1349 (O_1349,N_29116,N_29536);
or UO_1350 (O_1350,N_29616,N_29216);
nor UO_1351 (O_1351,N_29100,N_29468);
and UO_1352 (O_1352,N_29526,N_29550);
xnor UO_1353 (O_1353,N_29867,N_29263);
nor UO_1354 (O_1354,N_29642,N_29420);
or UO_1355 (O_1355,N_29245,N_29503);
xor UO_1356 (O_1356,N_28897,N_29540);
and UO_1357 (O_1357,N_29779,N_29559);
or UO_1358 (O_1358,N_29178,N_29096);
and UO_1359 (O_1359,N_29059,N_29996);
or UO_1360 (O_1360,N_29150,N_29572);
xnor UO_1361 (O_1361,N_29488,N_28892);
or UO_1362 (O_1362,N_29087,N_29275);
nand UO_1363 (O_1363,N_29012,N_29086);
nand UO_1364 (O_1364,N_29460,N_29098);
or UO_1365 (O_1365,N_29297,N_29335);
or UO_1366 (O_1366,N_29784,N_29647);
nand UO_1367 (O_1367,N_29541,N_29786);
or UO_1368 (O_1368,N_29784,N_29177);
or UO_1369 (O_1369,N_28900,N_29690);
nand UO_1370 (O_1370,N_29553,N_29343);
xor UO_1371 (O_1371,N_29242,N_29171);
and UO_1372 (O_1372,N_29751,N_29425);
xnor UO_1373 (O_1373,N_28879,N_29193);
xor UO_1374 (O_1374,N_29667,N_29035);
xnor UO_1375 (O_1375,N_29018,N_28953);
nor UO_1376 (O_1376,N_29901,N_28941);
nand UO_1377 (O_1377,N_28946,N_28912);
xor UO_1378 (O_1378,N_29000,N_28925);
or UO_1379 (O_1379,N_29395,N_28910);
nor UO_1380 (O_1380,N_29876,N_29192);
nand UO_1381 (O_1381,N_29140,N_29928);
nand UO_1382 (O_1382,N_29805,N_29396);
xnor UO_1383 (O_1383,N_29298,N_29665);
nor UO_1384 (O_1384,N_29141,N_29037);
nand UO_1385 (O_1385,N_29368,N_29910);
or UO_1386 (O_1386,N_29786,N_29317);
nor UO_1387 (O_1387,N_28900,N_29720);
or UO_1388 (O_1388,N_29379,N_28839);
and UO_1389 (O_1389,N_29207,N_29092);
and UO_1390 (O_1390,N_29460,N_29113);
nand UO_1391 (O_1391,N_28820,N_28942);
xor UO_1392 (O_1392,N_29608,N_28931);
nor UO_1393 (O_1393,N_29283,N_29608);
xor UO_1394 (O_1394,N_29741,N_29499);
nor UO_1395 (O_1395,N_29183,N_29804);
and UO_1396 (O_1396,N_29331,N_29622);
nand UO_1397 (O_1397,N_28899,N_29926);
or UO_1398 (O_1398,N_29428,N_29009);
nor UO_1399 (O_1399,N_29054,N_29415);
xor UO_1400 (O_1400,N_28846,N_29075);
nand UO_1401 (O_1401,N_29186,N_29768);
xnor UO_1402 (O_1402,N_28815,N_29498);
nand UO_1403 (O_1403,N_29883,N_29129);
and UO_1404 (O_1404,N_29442,N_29188);
nor UO_1405 (O_1405,N_29746,N_29184);
or UO_1406 (O_1406,N_29957,N_28865);
xor UO_1407 (O_1407,N_28994,N_29861);
nand UO_1408 (O_1408,N_29446,N_29790);
nand UO_1409 (O_1409,N_29128,N_28911);
xnor UO_1410 (O_1410,N_29030,N_29296);
nand UO_1411 (O_1411,N_28940,N_28857);
nand UO_1412 (O_1412,N_28953,N_29203);
xor UO_1413 (O_1413,N_29780,N_29268);
or UO_1414 (O_1414,N_29667,N_29172);
nor UO_1415 (O_1415,N_29381,N_29582);
nor UO_1416 (O_1416,N_29360,N_29088);
and UO_1417 (O_1417,N_29468,N_29879);
xor UO_1418 (O_1418,N_29501,N_29062);
and UO_1419 (O_1419,N_29573,N_29449);
nor UO_1420 (O_1420,N_29782,N_29616);
and UO_1421 (O_1421,N_29676,N_29974);
nor UO_1422 (O_1422,N_29273,N_29317);
xnor UO_1423 (O_1423,N_29610,N_29590);
xnor UO_1424 (O_1424,N_29093,N_29488);
or UO_1425 (O_1425,N_28975,N_29622);
or UO_1426 (O_1426,N_29000,N_29072);
xor UO_1427 (O_1427,N_29315,N_29566);
or UO_1428 (O_1428,N_29518,N_29392);
and UO_1429 (O_1429,N_29423,N_29330);
xor UO_1430 (O_1430,N_28880,N_29627);
xor UO_1431 (O_1431,N_29845,N_29062);
nand UO_1432 (O_1432,N_29193,N_29868);
xnor UO_1433 (O_1433,N_29371,N_29237);
nor UO_1434 (O_1434,N_29981,N_28992);
and UO_1435 (O_1435,N_29401,N_28814);
nand UO_1436 (O_1436,N_29276,N_29103);
xor UO_1437 (O_1437,N_29627,N_28944);
or UO_1438 (O_1438,N_28949,N_28942);
nor UO_1439 (O_1439,N_29904,N_29419);
nor UO_1440 (O_1440,N_29672,N_29933);
or UO_1441 (O_1441,N_29043,N_29727);
nand UO_1442 (O_1442,N_29873,N_29917);
and UO_1443 (O_1443,N_29495,N_28819);
or UO_1444 (O_1444,N_28827,N_29586);
xor UO_1445 (O_1445,N_29382,N_29689);
nor UO_1446 (O_1446,N_29474,N_29669);
xor UO_1447 (O_1447,N_29450,N_29939);
nor UO_1448 (O_1448,N_29908,N_29282);
or UO_1449 (O_1449,N_29595,N_29827);
xnor UO_1450 (O_1450,N_29248,N_29244);
or UO_1451 (O_1451,N_29943,N_29774);
nand UO_1452 (O_1452,N_29877,N_29035);
and UO_1453 (O_1453,N_28888,N_29087);
and UO_1454 (O_1454,N_29568,N_28865);
and UO_1455 (O_1455,N_29422,N_29088);
nor UO_1456 (O_1456,N_29091,N_29408);
nor UO_1457 (O_1457,N_29714,N_28930);
or UO_1458 (O_1458,N_29890,N_29187);
or UO_1459 (O_1459,N_29698,N_29528);
xnor UO_1460 (O_1460,N_29270,N_29506);
nor UO_1461 (O_1461,N_29392,N_29550);
xnor UO_1462 (O_1462,N_29690,N_29324);
or UO_1463 (O_1463,N_29238,N_28926);
xor UO_1464 (O_1464,N_29994,N_29374);
nor UO_1465 (O_1465,N_29793,N_29167);
or UO_1466 (O_1466,N_28944,N_29429);
or UO_1467 (O_1467,N_29173,N_29101);
and UO_1468 (O_1468,N_29816,N_29509);
and UO_1469 (O_1469,N_29564,N_28999);
nor UO_1470 (O_1470,N_29862,N_29611);
and UO_1471 (O_1471,N_29526,N_29189);
nand UO_1472 (O_1472,N_29335,N_29277);
and UO_1473 (O_1473,N_29090,N_29693);
and UO_1474 (O_1474,N_29023,N_29569);
nand UO_1475 (O_1475,N_28927,N_29853);
xnor UO_1476 (O_1476,N_29869,N_29667);
xnor UO_1477 (O_1477,N_28909,N_29165);
nor UO_1478 (O_1478,N_29772,N_28882);
xnor UO_1479 (O_1479,N_29546,N_29523);
xnor UO_1480 (O_1480,N_29838,N_29925);
xor UO_1481 (O_1481,N_29228,N_28832);
or UO_1482 (O_1482,N_29688,N_29619);
or UO_1483 (O_1483,N_29347,N_29438);
and UO_1484 (O_1484,N_28946,N_29704);
nand UO_1485 (O_1485,N_29346,N_29819);
nand UO_1486 (O_1486,N_29114,N_29389);
nor UO_1487 (O_1487,N_29204,N_28839);
xor UO_1488 (O_1488,N_29350,N_29349);
xnor UO_1489 (O_1489,N_28991,N_29364);
nor UO_1490 (O_1490,N_29139,N_29613);
xnor UO_1491 (O_1491,N_29180,N_29896);
and UO_1492 (O_1492,N_29603,N_29747);
xor UO_1493 (O_1493,N_28827,N_29434);
xnor UO_1494 (O_1494,N_29982,N_29387);
or UO_1495 (O_1495,N_29329,N_29785);
and UO_1496 (O_1496,N_29829,N_29499);
or UO_1497 (O_1497,N_28893,N_29571);
nand UO_1498 (O_1498,N_29428,N_29823);
and UO_1499 (O_1499,N_29786,N_28912);
nand UO_1500 (O_1500,N_29826,N_29222);
and UO_1501 (O_1501,N_29013,N_29154);
or UO_1502 (O_1502,N_28825,N_28883);
nor UO_1503 (O_1503,N_29647,N_29324);
nor UO_1504 (O_1504,N_29124,N_29505);
nand UO_1505 (O_1505,N_29453,N_28915);
and UO_1506 (O_1506,N_29885,N_29028);
nand UO_1507 (O_1507,N_29583,N_29690);
or UO_1508 (O_1508,N_29781,N_29995);
or UO_1509 (O_1509,N_29338,N_29229);
nand UO_1510 (O_1510,N_29676,N_29108);
xnor UO_1511 (O_1511,N_28826,N_28982);
and UO_1512 (O_1512,N_29959,N_29528);
nor UO_1513 (O_1513,N_29085,N_29601);
nor UO_1514 (O_1514,N_29584,N_29659);
or UO_1515 (O_1515,N_29705,N_29707);
nand UO_1516 (O_1516,N_29937,N_29343);
nand UO_1517 (O_1517,N_29974,N_29336);
nor UO_1518 (O_1518,N_28810,N_29191);
nor UO_1519 (O_1519,N_29861,N_29402);
nand UO_1520 (O_1520,N_28894,N_29454);
or UO_1521 (O_1521,N_29184,N_28919);
nor UO_1522 (O_1522,N_29776,N_29515);
or UO_1523 (O_1523,N_29296,N_28834);
nand UO_1524 (O_1524,N_29802,N_29441);
or UO_1525 (O_1525,N_29632,N_29283);
nor UO_1526 (O_1526,N_29445,N_28980);
nand UO_1527 (O_1527,N_28967,N_29428);
or UO_1528 (O_1528,N_28908,N_28875);
nor UO_1529 (O_1529,N_29313,N_29462);
nor UO_1530 (O_1530,N_28888,N_29751);
xor UO_1531 (O_1531,N_29367,N_29970);
nand UO_1532 (O_1532,N_29056,N_29014);
nor UO_1533 (O_1533,N_28809,N_29393);
xor UO_1534 (O_1534,N_29263,N_28944);
or UO_1535 (O_1535,N_29359,N_28956);
or UO_1536 (O_1536,N_29477,N_29055);
nor UO_1537 (O_1537,N_29428,N_29129);
nor UO_1538 (O_1538,N_29170,N_28882);
or UO_1539 (O_1539,N_28878,N_29713);
nor UO_1540 (O_1540,N_29080,N_29962);
xnor UO_1541 (O_1541,N_29913,N_29332);
or UO_1542 (O_1542,N_29505,N_29097);
nor UO_1543 (O_1543,N_29077,N_28997);
or UO_1544 (O_1544,N_29334,N_29289);
and UO_1545 (O_1545,N_29335,N_29637);
or UO_1546 (O_1546,N_28883,N_29799);
nor UO_1547 (O_1547,N_29387,N_29334);
xnor UO_1548 (O_1548,N_29510,N_29945);
nor UO_1549 (O_1549,N_29880,N_29314);
xor UO_1550 (O_1550,N_29304,N_29623);
xor UO_1551 (O_1551,N_29535,N_29855);
nand UO_1552 (O_1552,N_29786,N_28967);
nor UO_1553 (O_1553,N_29075,N_29106);
or UO_1554 (O_1554,N_29854,N_29180);
or UO_1555 (O_1555,N_29856,N_29054);
xnor UO_1556 (O_1556,N_29429,N_29592);
and UO_1557 (O_1557,N_29274,N_29476);
and UO_1558 (O_1558,N_29401,N_29616);
nor UO_1559 (O_1559,N_29849,N_29749);
xnor UO_1560 (O_1560,N_29525,N_29076);
or UO_1561 (O_1561,N_28926,N_28912);
or UO_1562 (O_1562,N_28819,N_29954);
nor UO_1563 (O_1563,N_29076,N_29509);
nor UO_1564 (O_1564,N_29521,N_29667);
and UO_1565 (O_1565,N_29115,N_29567);
and UO_1566 (O_1566,N_29828,N_29431);
or UO_1567 (O_1567,N_29652,N_29163);
and UO_1568 (O_1568,N_29155,N_28825);
nand UO_1569 (O_1569,N_29423,N_29871);
or UO_1570 (O_1570,N_29484,N_29231);
nand UO_1571 (O_1571,N_29953,N_29313);
and UO_1572 (O_1572,N_29547,N_29993);
or UO_1573 (O_1573,N_29973,N_29007);
and UO_1574 (O_1574,N_29674,N_29858);
nand UO_1575 (O_1575,N_28902,N_29261);
nor UO_1576 (O_1576,N_29668,N_29980);
nor UO_1577 (O_1577,N_28818,N_29277);
xnor UO_1578 (O_1578,N_29413,N_29344);
nor UO_1579 (O_1579,N_29883,N_29202);
or UO_1580 (O_1580,N_29938,N_29164);
nand UO_1581 (O_1581,N_29965,N_29931);
and UO_1582 (O_1582,N_29632,N_29177);
xor UO_1583 (O_1583,N_28869,N_29562);
or UO_1584 (O_1584,N_29338,N_29159);
xor UO_1585 (O_1585,N_28917,N_29956);
and UO_1586 (O_1586,N_29084,N_29130);
xnor UO_1587 (O_1587,N_29939,N_28952);
nor UO_1588 (O_1588,N_29931,N_29675);
nor UO_1589 (O_1589,N_29173,N_29760);
and UO_1590 (O_1590,N_29943,N_29248);
nand UO_1591 (O_1591,N_29325,N_28838);
nand UO_1592 (O_1592,N_29832,N_29221);
and UO_1593 (O_1593,N_29600,N_28921);
nand UO_1594 (O_1594,N_28860,N_29284);
nor UO_1595 (O_1595,N_29136,N_29481);
nor UO_1596 (O_1596,N_29340,N_29605);
nand UO_1597 (O_1597,N_29643,N_29351);
nand UO_1598 (O_1598,N_29985,N_29830);
xnor UO_1599 (O_1599,N_29598,N_28987);
xnor UO_1600 (O_1600,N_29908,N_29355);
or UO_1601 (O_1601,N_29111,N_29549);
xnor UO_1602 (O_1602,N_29970,N_29718);
xnor UO_1603 (O_1603,N_29110,N_28825);
nand UO_1604 (O_1604,N_29926,N_29113);
or UO_1605 (O_1605,N_29846,N_29349);
and UO_1606 (O_1606,N_29989,N_29593);
xnor UO_1607 (O_1607,N_29049,N_29583);
nand UO_1608 (O_1608,N_29968,N_29839);
and UO_1609 (O_1609,N_29027,N_29536);
xnor UO_1610 (O_1610,N_29651,N_29458);
xnor UO_1611 (O_1611,N_29924,N_29304);
and UO_1612 (O_1612,N_29253,N_29114);
nand UO_1613 (O_1613,N_29770,N_29708);
nand UO_1614 (O_1614,N_29447,N_29875);
xor UO_1615 (O_1615,N_29288,N_28935);
nor UO_1616 (O_1616,N_29541,N_29272);
xor UO_1617 (O_1617,N_29415,N_29136);
nand UO_1618 (O_1618,N_28870,N_29795);
and UO_1619 (O_1619,N_29299,N_28846);
nand UO_1620 (O_1620,N_29066,N_29948);
and UO_1621 (O_1621,N_29615,N_29981);
xnor UO_1622 (O_1622,N_29469,N_29349);
xnor UO_1623 (O_1623,N_29464,N_29396);
or UO_1624 (O_1624,N_29368,N_28940);
and UO_1625 (O_1625,N_29053,N_29927);
or UO_1626 (O_1626,N_29906,N_29214);
nor UO_1627 (O_1627,N_29254,N_29582);
and UO_1628 (O_1628,N_29557,N_29446);
or UO_1629 (O_1629,N_28887,N_29727);
and UO_1630 (O_1630,N_29289,N_29492);
nor UO_1631 (O_1631,N_29699,N_29772);
xnor UO_1632 (O_1632,N_29225,N_29584);
xor UO_1633 (O_1633,N_29498,N_29100);
xnor UO_1634 (O_1634,N_29290,N_29959);
and UO_1635 (O_1635,N_29188,N_29046);
and UO_1636 (O_1636,N_29499,N_29016);
and UO_1637 (O_1637,N_29004,N_29707);
and UO_1638 (O_1638,N_29814,N_29697);
nor UO_1639 (O_1639,N_29841,N_29065);
and UO_1640 (O_1640,N_28844,N_29912);
nand UO_1641 (O_1641,N_29871,N_28983);
nor UO_1642 (O_1642,N_28865,N_29244);
nor UO_1643 (O_1643,N_29167,N_29619);
or UO_1644 (O_1644,N_28955,N_28835);
or UO_1645 (O_1645,N_29380,N_29247);
nand UO_1646 (O_1646,N_29945,N_29782);
or UO_1647 (O_1647,N_29162,N_29557);
nand UO_1648 (O_1648,N_29888,N_29768);
or UO_1649 (O_1649,N_28839,N_29169);
xor UO_1650 (O_1650,N_29218,N_29872);
and UO_1651 (O_1651,N_29711,N_28843);
xnor UO_1652 (O_1652,N_29592,N_29009);
nand UO_1653 (O_1653,N_29744,N_29839);
nor UO_1654 (O_1654,N_29817,N_29171);
nand UO_1655 (O_1655,N_29464,N_29530);
nand UO_1656 (O_1656,N_28856,N_29152);
xor UO_1657 (O_1657,N_29310,N_29841);
or UO_1658 (O_1658,N_28952,N_29432);
and UO_1659 (O_1659,N_29251,N_29478);
nand UO_1660 (O_1660,N_29817,N_29295);
or UO_1661 (O_1661,N_28800,N_29622);
or UO_1662 (O_1662,N_28927,N_29651);
nor UO_1663 (O_1663,N_29621,N_29780);
nand UO_1664 (O_1664,N_29083,N_29035);
nand UO_1665 (O_1665,N_29957,N_29832);
nor UO_1666 (O_1666,N_29118,N_29131);
nor UO_1667 (O_1667,N_29085,N_29840);
and UO_1668 (O_1668,N_29283,N_28825);
xnor UO_1669 (O_1669,N_29199,N_29299);
nand UO_1670 (O_1670,N_29591,N_29907);
nand UO_1671 (O_1671,N_29468,N_29444);
nor UO_1672 (O_1672,N_29519,N_29340);
nand UO_1673 (O_1673,N_29172,N_29380);
and UO_1674 (O_1674,N_29926,N_29225);
and UO_1675 (O_1675,N_29351,N_29598);
nand UO_1676 (O_1676,N_29175,N_29864);
and UO_1677 (O_1677,N_29916,N_29683);
or UO_1678 (O_1678,N_29245,N_29047);
or UO_1679 (O_1679,N_28829,N_29031);
nand UO_1680 (O_1680,N_29592,N_29712);
and UO_1681 (O_1681,N_29504,N_28921);
and UO_1682 (O_1682,N_28952,N_29575);
nand UO_1683 (O_1683,N_29461,N_29964);
xnor UO_1684 (O_1684,N_29053,N_29928);
and UO_1685 (O_1685,N_29298,N_29539);
and UO_1686 (O_1686,N_28815,N_29510);
nand UO_1687 (O_1687,N_29507,N_29512);
or UO_1688 (O_1688,N_29597,N_28831);
and UO_1689 (O_1689,N_29781,N_28857);
xor UO_1690 (O_1690,N_29435,N_29827);
nand UO_1691 (O_1691,N_28820,N_29892);
or UO_1692 (O_1692,N_29625,N_29268);
nor UO_1693 (O_1693,N_29716,N_29470);
nand UO_1694 (O_1694,N_29334,N_29641);
and UO_1695 (O_1695,N_29854,N_29868);
xor UO_1696 (O_1696,N_29059,N_29801);
nor UO_1697 (O_1697,N_29389,N_29134);
and UO_1698 (O_1698,N_29309,N_29802);
or UO_1699 (O_1699,N_29670,N_29881);
nor UO_1700 (O_1700,N_28933,N_28844);
xor UO_1701 (O_1701,N_29269,N_29325);
nor UO_1702 (O_1702,N_29701,N_29403);
and UO_1703 (O_1703,N_29568,N_29881);
and UO_1704 (O_1704,N_29382,N_29868);
nor UO_1705 (O_1705,N_28983,N_29399);
xor UO_1706 (O_1706,N_28805,N_29477);
xor UO_1707 (O_1707,N_28988,N_29931);
nor UO_1708 (O_1708,N_29285,N_29790);
or UO_1709 (O_1709,N_29638,N_28868);
or UO_1710 (O_1710,N_29428,N_28997);
and UO_1711 (O_1711,N_29289,N_29659);
and UO_1712 (O_1712,N_29953,N_29368);
and UO_1713 (O_1713,N_29753,N_29267);
xor UO_1714 (O_1714,N_29698,N_29076);
or UO_1715 (O_1715,N_29334,N_29831);
nor UO_1716 (O_1716,N_28803,N_29131);
xor UO_1717 (O_1717,N_29259,N_28975);
nand UO_1718 (O_1718,N_29061,N_29746);
or UO_1719 (O_1719,N_29976,N_29871);
or UO_1720 (O_1720,N_29815,N_29606);
or UO_1721 (O_1721,N_29508,N_29494);
nand UO_1722 (O_1722,N_29380,N_29659);
nand UO_1723 (O_1723,N_29969,N_28920);
nor UO_1724 (O_1724,N_29888,N_29424);
and UO_1725 (O_1725,N_29947,N_29256);
and UO_1726 (O_1726,N_29210,N_29972);
xnor UO_1727 (O_1727,N_29378,N_28963);
nand UO_1728 (O_1728,N_28869,N_29323);
xnor UO_1729 (O_1729,N_29870,N_29491);
nor UO_1730 (O_1730,N_28901,N_29976);
nor UO_1731 (O_1731,N_29857,N_28942);
and UO_1732 (O_1732,N_29821,N_29315);
xnor UO_1733 (O_1733,N_29511,N_29793);
and UO_1734 (O_1734,N_29388,N_29058);
nor UO_1735 (O_1735,N_29658,N_29343);
xnor UO_1736 (O_1736,N_29022,N_29455);
or UO_1737 (O_1737,N_29265,N_28902);
nand UO_1738 (O_1738,N_29338,N_29555);
nand UO_1739 (O_1739,N_28952,N_29358);
nand UO_1740 (O_1740,N_29601,N_29417);
or UO_1741 (O_1741,N_29247,N_29786);
nor UO_1742 (O_1742,N_29648,N_29846);
nand UO_1743 (O_1743,N_29401,N_29393);
and UO_1744 (O_1744,N_29531,N_28845);
and UO_1745 (O_1745,N_29943,N_29429);
xnor UO_1746 (O_1746,N_29102,N_29371);
or UO_1747 (O_1747,N_29677,N_29104);
and UO_1748 (O_1748,N_29496,N_29433);
and UO_1749 (O_1749,N_29117,N_29808);
or UO_1750 (O_1750,N_29536,N_29265);
xnor UO_1751 (O_1751,N_29706,N_29440);
nand UO_1752 (O_1752,N_29305,N_29868);
nor UO_1753 (O_1753,N_29705,N_29339);
nor UO_1754 (O_1754,N_29249,N_29392);
nor UO_1755 (O_1755,N_29389,N_29905);
nor UO_1756 (O_1756,N_29457,N_29162);
nor UO_1757 (O_1757,N_29780,N_29928);
and UO_1758 (O_1758,N_29766,N_29839);
nand UO_1759 (O_1759,N_29069,N_28947);
nor UO_1760 (O_1760,N_29734,N_29159);
nor UO_1761 (O_1761,N_29301,N_29146);
nor UO_1762 (O_1762,N_28929,N_29070);
nor UO_1763 (O_1763,N_29791,N_29189);
nor UO_1764 (O_1764,N_29524,N_28958);
nand UO_1765 (O_1765,N_29319,N_29207);
and UO_1766 (O_1766,N_29413,N_29895);
xnor UO_1767 (O_1767,N_29357,N_29839);
or UO_1768 (O_1768,N_29095,N_29872);
xnor UO_1769 (O_1769,N_29090,N_29186);
nor UO_1770 (O_1770,N_29735,N_29858);
xor UO_1771 (O_1771,N_28822,N_28820);
or UO_1772 (O_1772,N_29196,N_29016);
and UO_1773 (O_1773,N_29136,N_29482);
nand UO_1774 (O_1774,N_29906,N_29007);
or UO_1775 (O_1775,N_29396,N_29536);
nor UO_1776 (O_1776,N_29927,N_28995);
and UO_1777 (O_1777,N_29993,N_29312);
nand UO_1778 (O_1778,N_29737,N_29580);
xor UO_1779 (O_1779,N_29576,N_29423);
nand UO_1780 (O_1780,N_29984,N_29356);
nand UO_1781 (O_1781,N_29488,N_29774);
nor UO_1782 (O_1782,N_29241,N_29883);
xor UO_1783 (O_1783,N_29292,N_29051);
nand UO_1784 (O_1784,N_29530,N_29586);
and UO_1785 (O_1785,N_29910,N_29994);
or UO_1786 (O_1786,N_29987,N_29520);
xor UO_1787 (O_1787,N_29419,N_28855);
nor UO_1788 (O_1788,N_29890,N_29711);
nor UO_1789 (O_1789,N_29626,N_29218);
xor UO_1790 (O_1790,N_29150,N_29712);
and UO_1791 (O_1791,N_28962,N_28878);
nor UO_1792 (O_1792,N_28915,N_29921);
xnor UO_1793 (O_1793,N_29064,N_29982);
nand UO_1794 (O_1794,N_29504,N_28903);
or UO_1795 (O_1795,N_28907,N_28849);
and UO_1796 (O_1796,N_28873,N_29967);
xor UO_1797 (O_1797,N_29883,N_29220);
or UO_1798 (O_1798,N_29828,N_29811);
nor UO_1799 (O_1799,N_29020,N_29565);
nand UO_1800 (O_1800,N_29843,N_29694);
and UO_1801 (O_1801,N_29345,N_29138);
and UO_1802 (O_1802,N_29591,N_29951);
and UO_1803 (O_1803,N_29462,N_29350);
or UO_1804 (O_1804,N_29507,N_28977);
or UO_1805 (O_1805,N_29180,N_29277);
nand UO_1806 (O_1806,N_28913,N_29597);
and UO_1807 (O_1807,N_29852,N_29003);
or UO_1808 (O_1808,N_28996,N_28825);
xnor UO_1809 (O_1809,N_29853,N_28931);
and UO_1810 (O_1810,N_29745,N_29860);
or UO_1811 (O_1811,N_28819,N_29305);
nor UO_1812 (O_1812,N_29446,N_29022);
nand UO_1813 (O_1813,N_29528,N_29425);
and UO_1814 (O_1814,N_29886,N_28955);
or UO_1815 (O_1815,N_29980,N_29421);
or UO_1816 (O_1816,N_29194,N_29846);
nand UO_1817 (O_1817,N_29597,N_28815);
or UO_1818 (O_1818,N_29185,N_28964);
or UO_1819 (O_1819,N_29356,N_29410);
nand UO_1820 (O_1820,N_29010,N_29539);
or UO_1821 (O_1821,N_29446,N_29396);
and UO_1822 (O_1822,N_29247,N_29712);
or UO_1823 (O_1823,N_28835,N_28976);
xor UO_1824 (O_1824,N_29143,N_29137);
or UO_1825 (O_1825,N_29723,N_29082);
nor UO_1826 (O_1826,N_29941,N_29246);
xnor UO_1827 (O_1827,N_29341,N_29837);
or UO_1828 (O_1828,N_29704,N_29062);
nand UO_1829 (O_1829,N_29854,N_29844);
and UO_1830 (O_1830,N_29471,N_29676);
xor UO_1831 (O_1831,N_29234,N_29677);
and UO_1832 (O_1832,N_29530,N_29201);
or UO_1833 (O_1833,N_29485,N_29543);
nor UO_1834 (O_1834,N_29494,N_29526);
nand UO_1835 (O_1835,N_29103,N_29236);
xor UO_1836 (O_1836,N_29331,N_28807);
nand UO_1837 (O_1837,N_29617,N_29108);
and UO_1838 (O_1838,N_29962,N_29299);
nand UO_1839 (O_1839,N_29778,N_29888);
and UO_1840 (O_1840,N_29805,N_29890);
nor UO_1841 (O_1841,N_29565,N_29705);
nor UO_1842 (O_1842,N_29579,N_29513);
or UO_1843 (O_1843,N_28932,N_29212);
and UO_1844 (O_1844,N_28884,N_29556);
and UO_1845 (O_1845,N_29117,N_29336);
or UO_1846 (O_1846,N_28972,N_29711);
or UO_1847 (O_1847,N_29295,N_29843);
nand UO_1848 (O_1848,N_29391,N_29288);
xor UO_1849 (O_1849,N_29330,N_28826);
or UO_1850 (O_1850,N_29559,N_29899);
xor UO_1851 (O_1851,N_29298,N_29920);
nor UO_1852 (O_1852,N_29933,N_29173);
xor UO_1853 (O_1853,N_29851,N_29563);
or UO_1854 (O_1854,N_29392,N_29696);
nand UO_1855 (O_1855,N_29253,N_29274);
nor UO_1856 (O_1856,N_29991,N_29901);
nor UO_1857 (O_1857,N_29855,N_28924);
nand UO_1858 (O_1858,N_29719,N_29312);
xor UO_1859 (O_1859,N_29250,N_29366);
nand UO_1860 (O_1860,N_29811,N_29078);
xor UO_1861 (O_1861,N_29933,N_29836);
nand UO_1862 (O_1862,N_29620,N_29607);
xnor UO_1863 (O_1863,N_29170,N_28856);
nand UO_1864 (O_1864,N_29450,N_29786);
xnor UO_1865 (O_1865,N_29565,N_29582);
or UO_1866 (O_1866,N_29093,N_29990);
nor UO_1867 (O_1867,N_29817,N_29403);
nor UO_1868 (O_1868,N_29420,N_29859);
or UO_1869 (O_1869,N_29950,N_29578);
or UO_1870 (O_1870,N_29791,N_29480);
nor UO_1871 (O_1871,N_29479,N_29422);
and UO_1872 (O_1872,N_29301,N_29795);
and UO_1873 (O_1873,N_29046,N_28997);
xnor UO_1874 (O_1874,N_29296,N_29984);
xor UO_1875 (O_1875,N_28948,N_29303);
nor UO_1876 (O_1876,N_29974,N_29568);
nor UO_1877 (O_1877,N_28829,N_29518);
nand UO_1878 (O_1878,N_29240,N_29187);
and UO_1879 (O_1879,N_29193,N_28988);
nand UO_1880 (O_1880,N_29824,N_29378);
or UO_1881 (O_1881,N_29075,N_29906);
xor UO_1882 (O_1882,N_29452,N_29768);
xor UO_1883 (O_1883,N_29998,N_29259);
or UO_1884 (O_1884,N_29572,N_28909);
xor UO_1885 (O_1885,N_28967,N_28991);
nand UO_1886 (O_1886,N_29952,N_29121);
nor UO_1887 (O_1887,N_28882,N_29273);
nor UO_1888 (O_1888,N_29616,N_29289);
and UO_1889 (O_1889,N_29413,N_29411);
xnor UO_1890 (O_1890,N_29607,N_29122);
nor UO_1891 (O_1891,N_29553,N_28996);
and UO_1892 (O_1892,N_29983,N_29707);
nor UO_1893 (O_1893,N_29518,N_29418);
nand UO_1894 (O_1894,N_28976,N_29463);
xor UO_1895 (O_1895,N_29921,N_28921);
or UO_1896 (O_1896,N_29242,N_29759);
nand UO_1897 (O_1897,N_28838,N_29608);
nor UO_1898 (O_1898,N_29404,N_29164);
nor UO_1899 (O_1899,N_29032,N_29066);
xor UO_1900 (O_1900,N_29089,N_29875);
xor UO_1901 (O_1901,N_29117,N_28845);
xor UO_1902 (O_1902,N_28905,N_28901);
and UO_1903 (O_1903,N_29816,N_29765);
xnor UO_1904 (O_1904,N_29681,N_29765);
nand UO_1905 (O_1905,N_29331,N_29210);
nand UO_1906 (O_1906,N_29099,N_29441);
and UO_1907 (O_1907,N_29883,N_29578);
or UO_1908 (O_1908,N_28908,N_29993);
or UO_1909 (O_1909,N_29480,N_28941);
nor UO_1910 (O_1910,N_29466,N_29736);
or UO_1911 (O_1911,N_29743,N_29506);
nor UO_1912 (O_1912,N_29225,N_28931);
xnor UO_1913 (O_1913,N_29502,N_29058);
xor UO_1914 (O_1914,N_29774,N_28990);
and UO_1915 (O_1915,N_29939,N_29554);
nand UO_1916 (O_1916,N_29700,N_29926);
nand UO_1917 (O_1917,N_29743,N_28882);
nor UO_1918 (O_1918,N_28932,N_29056);
nor UO_1919 (O_1919,N_29829,N_28852);
nand UO_1920 (O_1920,N_28965,N_28932);
or UO_1921 (O_1921,N_28825,N_29680);
nor UO_1922 (O_1922,N_29411,N_29242);
nand UO_1923 (O_1923,N_29894,N_29694);
nand UO_1924 (O_1924,N_29404,N_29730);
nand UO_1925 (O_1925,N_29165,N_28894);
or UO_1926 (O_1926,N_29202,N_29502);
nand UO_1927 (O_1927,N_29995,N_29210);
and UO_1928 (O_1928,N_29560,N_29529);
nor UO_1929 (O_1929,N_29197,N_29053);
and UO_1930 (O_1930,N_28861,N_29330);
nand UO_1931 (O_1931,N_29531,N_29593);
nand UO_1932 (O_1932,N_29209,N_29863);
xor UO_1933 (O_1933,N_28930,N_29968);
nor UO_1934 (O_1934,N_29031,N_29721);
and UO_1935 (O_1935,N_29810,N_29657);
or UO_1936 (O_1936,N_29105,N_29991);
and UO_1937 (O_1937,N_29064,N_29019);
or UO_1938 (O_1938,N_29240,N_29657);
xor UO_1939 (O_1939,N_29082,N_29687);
or UO_1940 (O_1940,N_29147,N_29258);
or UO_1941 (O_1941,N_29948,N_29634);
and UO_1942 (O_1942,N_29553,N_29796);
nor UO_1943 (O_1943,N_29510,N_28894);
xor UO_1944 (O_1944,N_29191,N_29423);
and UO_1945 (O_1945,N_29881,N_29503);
nor UO_1946 (O_1946,N_29069,N_29206);
xnor UO_1947 (O_1947,N_29209,N_29817);
xnor UO_1948 (O_1948,N_28869,N_29435);
and UO_1949 (O_1949,N_29624,N_29390);
xor UO_1950 (O_1950,N_28956,N_29941);
xnor UO_1951 (O_1951,N_29268,N_29463);
or UO_1952 (O_1952,N_29126,N_29700);
and UO_1953 (O_1953,N_29521,N_29130);
nand UO_1954 (O_1954,N_29960,N_29235);
nand UO_1955 (O_1955,N_28990,N_29167);
nor UO_1956 (O_1956,N_28843,N_29134);
or UO_1957 (O_1957,N_29887,N_29547);
nand UO_1958 (O_1958,N_28819,N_29957);
xnor UO_1959 (O_1959,N_29286,N_29428);
nand UO_1960 (O_1960,N_29163,N_29260);
xor UO_1961 (O_1961,N_29828,N_29966);
xor UO_1962 (O_1962,N_29971,N_29712);
nand UO_1963 (O_1963,N_29617,N_29542);
xnor UO_1964 (O_1964,N_29123,N_28865);
nor UO_1965 (O_1965,N_29315,N_28855);
or UO_1966 (O_1966,N_29693,N_28850);
or UO_1967 (O_1967,N_29548,N_29781);
xnor UO_1968 (O_1968,N_29140,N_29201);
nor UO_1969 (O_1969,N_28854,N_29360);
xnor UO_1970 (O_1970,N_28834,N_29407);
or UO_1971 (O_1971,N_29667,N_29216);
and UO_1972 (O_1972,N_29741,N_29408);
nor UO_1973 (O_1973,N_29173,N_29008);
or UO_1974 (O_1974,N_28911,N_29161);
xnor UO_1975 (O_1975,N_29333,N_29936);
nor UO_1976 (O_1976,N_29437,N_29646);
xor UO_1977 (O_1977,N_29630,N_29322);
xnor UO_1978 (O_1978,N_29553,N_29108);
and UO_1979 (O_1979,N_29364,N_29185);
xor UO_1980 (O_1980,N_29900,N_29574);
and UO_1981 (O_1981,N_29661,N_28922);
or UO_1982 (O_1982,N_29333,N_28902);
nand UO_1983 (O_1983,N_29290,N_29517);
xnor UO_1984 (O_1984,N_29857,N_29400);
xnor UO_1985 (O_1985,N_28832,N_29396);
nor UO_1986 (O_1986,N_29720,N_28944);
nor UO_1987 (O_1987,N_29201,N_29387);
and UO_1988 (O_1988,N_28943,N_29917);
xor UO_1989 (O_1989,N_29093,N_29022);
or UO_1990 (O_1990,N_29217,N_29816);
nand UO_1991 (O_1991,N_29613,N_29529);
nand UO_1992 (O_1992,N_29880,N_29721);
xor UO_1993 (O_1993,N_28858,N_28919);
nor UO_1994 (O_1994,N_28905,N_28856);
xor UO_1995 (O_1995,N_29262,N_29099);
and UO_1996 (O_1996,N_29783,N_28835);
xor UO_1997 (O_1997,N_29218,N_29561);
nand UO_1998 (O_1998,N_28909,N_28923);
and UO_1999 (O_1999,N_29185,N_29209);
nand UO_2000 (O_2000,N_29739,N_29771);
or UO_2001 (O_2001,N_28854,N_29602);
nand UO_2002 (O_2002,N_29348,N_29816);
nor UO_2003 (O_2003,N_29680,N_28877);
and UO_2004 (O_2004,N_29693,N_29578);
nor UO_2005 (O_2005,N_28800,N_29764);
nand UO_2006 (O_2006,N_29559,N_29924);
nor UO_2007 (O_2007,N_29872,N_29515);
and UO_2008 (O_2008,N_29185,N_29981);
or UO_2009 (O_2009,N_29420,N_29378);
xor UO_2010 (O_2010,N_29322,N_29929);
nor UO_2011 (O_2011,N_29272,N_29456);
or UO_2012 (O_2012,N_29176,N_29548);
nand UO_2013 (O_2013,N_29623,N_29680);
or UO_2014 (O_2014,N_29844,N_29147);
or UO_2015 (O_2015,N_29073,N_28849);
nor UO_2016 (O_2016,N_29405,N_29513);
xor UO_2017 (O_2017,N_28903,N_29758);
and UO_2018 (O_2018,N_29810,N_29881);
nand UO_2019 (O_2019,N_29083,N_28810);
and UO_2020 (O_2020,N_29398,N_28889);
and UO_2021 (O_2021,N_29361,N_29547);
nand UO_2022 (O_2022,N_29381,N_29712);
nand UO_2023 (O_2023,N_29158,N_29100);
xnor UO_2024 (O_2024,N_29689,N_29786);
and UO_2025 (O_2025,N_29894,N_29333);
nand UO_2026 (O_2026,N_29881,N_28904);
nor UO_2027 (O_2027,N_28861,N_29706);
nor UO_2028 (O_2028,N_29523,N_29010);
and UO_2029 (O_2029,N_29208,N_29978);
or UO_2030 (O_2030,N_29187,N_29891);
nand UO_2031 (O_2031,N_29951,N_29964);
nor UO_2032 (O_2032,N_29986,N_29807);
xnor UO_2033 (O_2033,N_28931,N_29655);
xnor UO_2034 (O_2034,N_28888,N_29178);
xor UO_2035 (O_2035,N_29120,N_29689);
nand UO_2036 (O_2036,N_29227,N_29681);
nor UO_2037 (O_2037,N_28882,N_29346);
nor UO_2038 (O_2038,N_29922,N_29250);
nand UO_2039 (O_2039,N_29164,N_29111);
nor UO_2040 (O_2040,N_29651,N_29137);
nor UO_2041 (O_2041,N_29965,N_28892);
xor UO_2042 (O_2042,N_29649,N_28851);
xnor UO_2043 (O_2043,N_28889,N_29124);
or UO_2044 (O_2044,N_29227,N_28829);
nor UO_2045 (O_2045,N_28881,N_29766);
nor UO_2046 (O_2046,N_29262,N_29286);
and UO_2047 (O_2047,N_29459,N_29331);
and UO_2048 (O_2048,N_29855,N_29024);
nand UO_2049 (O_2049,N_29521,N_29067);
nand UO_2050 (O_2050,N_29286,N_29847);
nand UO_2051 (O_2051,N_29040,N_29744);
and UO_2052 (O_2052,N_29584,N_29627);
nand UO_2053 (O_2053,N_29184,N_29031);
nand UO_2054 (O_2054,N_29314,N_29695);
and UO_2055 (O_2055,N_29944,N_29190);
xnor UO_2056 (O_2056,N_28834,N_29230);
nand UO_2057 (O_2057,N_29321,N_28971);
nor UO_2058 (O_2058,N_29952,N_29755);
or UO_2059 (O_2059,N_29767,N_28909);
nand UO_2060 (O_2060,N_28889,N_29627);
xnor UO_2061 (O_2061,N_29589,N_29510);
xor UO_2062 (O_2062,N_29062,N_28820);
nor UO_2063 (O_2063,N_29251,N_29575);
nand UO_2064 (O_2064,N_29366,N_29438);
nand UO_2065 (O_2065,N_29261,N_29467);
or UO_2066 (O_2066,N_29010,N_29107);
and UO_2067 (O_2067,N_29034,N_29569);
and UO_2068 (O_2068,N_29388,N_29750);
and UO_2069 (O_2069,N_28864,N_29617);
and UO_2070 (O_2070,N_29202,N_29277);
or UO_2071 (O_2071,N_29207,N_29221);
and UO_2072 (O_2072,N_29990,N_29293);
and UO_2073 (O_2073,N_29471,N_29531);
nand UO_2074 (O_2074,N_28836,N_29137);
xnor UO_2075 (O_2075,N_29429,N_29713);
nor UO_2076 (O_2076,N_29525,N_29178);
nor UO_2077 (O_2077,N_29525,N_29739);
nor UO_2078 (O_2078,N_28846,N_29879);
and UO_2079 (O_2079,N_29167,N_29612);
and UO_2080 (O_2080,N_29620,N_29032);
nand UO_2081 (O_2081,N_29339,N_28819);
or UO_2082 (O_2082,N_29541,N_28825);
and UO_2083 (O_2083,N_28963,N_29985);
or UO_2084 (O_2084,N_29965,N_29403);
nand UO_2085 (O_2085,N_29890,N_29893);
and UO_2086 (O_2086,N_29668,N_29756);
nor UO_2087 (O_2087,N_28884,N_29430);
and UO_2088 (O_2088,N_29697,N_29140);
nand UO_2089 (O_2089,N_29887,N_29290);
xor UO_2090 (O_2090,N_29372,N_29763);
and UO_2091 (O_2091,N_29575,N_28868);
or UO_2092 (O_2092,N_29386,N_29158);
nor UO_2093 (O_2093,N_29593,N_29244);
nor UO_2094 (O_2094,N_29232,N_29300);
nor UO_2095 (O_2095,N_28830,N_29557);
and UO_2096 (O_2096,N_29054,N_28849);
or UO_2097 (O_2097,N_29853,N_28817);
or UO_2098 (O_2098,N_29773,N_29246);
xnor UO_2099 (O_2099,N_29748,N_29215);
nand UO_2100 (O_2100,N_29105,N_29657);
and UO_2101 (O_2101,N_29672,N_29605);
and UO_2102 (O_2102,N_29595,N_29341);
nand UO_2103 (O_2103,N_29989,N_29207);
and UO_2104 (O_2104,N_29018,N_29921);
or UO_2105 (O_2105,N_29248,N_29855);
nand UO_2106 (O_2106,N_29386,N_29470);
and UO_2107 (O_2107,N_29565,N_29153);
xnor UO_2108 (O_2108,N_29950,N_29498);
and UO_2109 (O_2109,N_29749,N_28872);
nor UO_2110 (O_2110,N_29771,N_29392);
nand UO_2111 (O_2111,N_29773,N_29446);
xor UO_2112 (O_2112,N_29066,N_29533);
nand UO_2113 (O_2113,N_29086,N_28847);
or UO_2114 (O_2114,N_29595,N_29964);
nor UO_2115 (O_2115,N_28832,N_29130);
xor UO_2116 (O_2116,N_29503,N_29368);
or UO_2117 (O_2117,N_29861,N_29578);
or UO_2118 (O_2118,N_29439,N_29868);
and UO_2119 (O_2119,N_29340,N_29187);
and UO_2120 (O_2120,N_29993,N_29263);
nor UO_2121 (O_2121,N_29425,N_29377);
nand UO_2122 (O_2122,N_29713,N_28823);
nand UO_2123 (O_2123,N_29965,N_29374);
nor UO_2124 (O_2124,N_29214,N_29999);
nand UO_2125 (O_2125,N_29203,N_29194);
nand UO_2126 (O_2126,N_29513,N_29909);
xor UO_2127 (O_2127,N_29857,N_29583);
or UO_2128 (O_2128,N_29843,N_29299);
or UO_2129 (O_2129,N_29714,N_29497);
nand UO_2130 (O_2130,N_29783,N_29764);
and UO_2131 (O_2131,N_28975,N_29142);
xor UO_2132 (O_2132,N_29393,N_28853);
xor UO_2133 (O_2133,N_29380,N_29028);
and UO_2134 (O_2134,N_29150,N_28857);
and UO_2135 (O_2135,N_29711,N_29217);
nor UO_2136 (O_2136,N_29489,N_29055);
xor UO_2137 (O_2137,N_29576,N_29566);
nand UO_2138 (O_2138,N_29046,N_28916);
xor UO_2139 (O_2139,N_29542,N_29622);
xnor UO_2140 (O_2140,N_29729,N_29125);
and UO_2141 (O_2141,N_29124,N_29873);
or UO_2142 (O_2142,N_29631,N_29811);
nor UO_2143 (O_2143,N_29946,N_28865);
nor UO_2144 (O_2144,N_29048,N_28860);
and UO_2145 (O_2145,N_29896,N_28943);
nand UO_2146 (O_2146,N_29579,N_29611);
nor UO_2147 (O_2147,N_29136,N_29792);
nand UO_2148 (O_2148,N_29301,N_29425);
or UO_2149 (O_2149,N_29177,N_29983);
or UO_2150 (O_2150,N_28849,N_29966);
nor UO_2151 (O_2151,N_29183,N_28841);
xnor UO_2152 (O_2152,N_28963,N_28940);
nand UO_2153 (O_2153,N_29818,N_29562);
nor UO_2154 (O_2154,N_29242,N_29351);
nand UO_2155 (O_2155,N_28899,N_29658);
nand UO_2156 (O_2156,N_29287,N_29850);
or UO_2157 (O_2157,N_29981,N_28831);
or UO_2158 (O_2158,N_29673,N_28927);
and UO_2159 (O_2159,N_29666,N_29100);
nor UO_2160 (O_2160,N_29737,N_29430);
xnor UO_2161 (O_2161,N_28938,N_29504);
xor UO_2162 (O_2162,N_28988,N_29057);
and UO_2163 (O_2163,N_29814,N_29229);
or UO_2164 (O_2164,N_29035,N_29613);
and UO_2165 (O_2165,N_29620,N_29141);
nand UO_2166 (O_2166,N_29187,N_29745);
xor UO_2167 (O_2167,N_29982,N_29133);
xor UO_2168 (O_2168,N_29227,N_29974);
nand UO_2169 (O_2169,N_29119,N_28843);
xnor UO_2170 (O_2170,N_29773,N_29979);
or UO_2171 (O_2171,N_29105,N_29156);
nor UO_2172 (O_2172,N_29508,N_29484);
nand UO_2173 (O_2173,N_28902,N_29514);
or UO_2174 (O_2174,N_29515,N_29418);
nor UO_2175 (O_2175,N_29222,N_29697);
xnor UO_2176 (O_2176,N_29035,N_29617);
and UO_2177 (O_2177,N_29989,N_29164);
nor UO_2178 (O_2178,N_29307,N_29944);
nand UO_2179 (O_2179,N_29353,N_29911);
or UO_2180 (O_2180,N_29792,N_29347);
xor UO_2181 (O_2181,N_29884,N_28987);
xnor UO_2182 (O_2182,N_29533,N_29552);
nand UO_2183 (O_2183,N_29586,N_29271);
xnor UO_2184 (O_2184,N_29612,N_29051);
nor UO_2185 (O_2185,N_29623,N_29889);
xor UO_2186 (O_2186,N_29920,N_29241);
nand UO_2187 (O_2187,N_29186,N_28984);
nand UO_2188 (O_2188,N_29798,N_29733);
nor UO_2189 (O_2189,N_28825,N_29345);
nand UO_2190 (O_2190,N_29428,N_29266);
or UO_2191 (O_2191,N_29800,N_29405);
and UO_2192 (O_2192,N_29485,N_29726);
nand UO_2193 (O_2193,N_29763,N_29956);
or UO_2194 (O_2194,N_29872,N_29999);
and UO_2195 (O_2195,N_28868,N_29641);
or UO_2196 (O_2196,N_28881,N_29466);
and UO_2197 (O_2197,N_29541,N_29156);
xnor UO_2198 (O_2198,N_29761,N_28803);
and UO_2199 (O_2199,N_29414,N_29010);
and UO_2200 (O_2200,N_29851,N_29653);
nand UO_2201 (O_2201,N_29861,N_29080);
and UO_2202 (O_2202,N_29409,N_29856);
nand UO_2203 (O_2203,N_29697,N_29830);
xnor UO_2204 (O_2204,N_28951,N_29924);
nor UO_2205 (O_2205,N_29069,N_29954);
nand UO_2206 (O_2206,N_28908,N_29019);
nor UO_2207 (O_2207,N_29743,N_28975);
and UO_2208 (O_2208,N_29509,N_28821);
and UO_2209 (O_2209,N_28992,N_29249);
nor UO_2210 (O_2210,N_29853,N_29792);
nand UO_2211 (O_2211,N_28963,N_29903);
nand UO_2212 (O_2212,N_29419,N_29098);
xnor UO_2213 (O_2213,N_29452,N_29214);
or UO_2214 (O_2214,N_29651,N_29096);
nor UO_2215 (O_2215,N_29746,N_29464);
or UO_2216 (O_2216,N_29715,N_29169);
xor UO_2217 (O_2217,N_29609,N_29754);
or UO_2218 (O_2218,N_29911,N_29122);
nand UO_2219 (O_2219,N_28874,N_28841);
nor UO_2220 (O_2220,N_29878,N_29303);
or UO_2221 (O_2221,N_29056,N_29461);
and UO_2222 (O_2222,N_29837,N_29502);
nor UO_2223 (O_2223,N_29745,N_28938);
nand UO_2224 (O_2224,N_29855,N_29802);
xnor UO_2225 (O_2225,N_29445,N_29636);
nor UO_2226 (O_2226,N_28978,N_29992);
and UO_2227 (O_2227,N_29439,N_29169);
nor UO_2228 (O_2228,N_29783,N_29131);
or UO_2229 (O_2229,N_29080,N_28935);
xor UO_2230 (O_2230,N_28809,N_29480);
xnor UO_2231 (O_2231,N_29775,N_28935);
and UO_2232 (O_2232,N_29004,N_29951);
nor UO_2233 (O_2233,N_29835,N_29543);
and UO_2234 (O_2234,N_29957,N_29888);
nor UO_2235 (O_2235,N_29218,N_28968);
nor UO_2236 (O_2236,N_28900,N_29774);
nand UO_2237 (O_2237,N_29931,N_29527);
and UO_2238 (O_2238,N_29523,N_28902);
and UO_2239 (O_2239,N_28818,N_29144);
or UO_2240 (O_2240,N_29426,N_29305);
nor UO_2241 (O_2241,N_28922,N_29943);
nand UO_2242 (O_2242,N_29087,N_29759);
and UO_2243 (O_2243,N_29625,N_29316);
nor UO_2244 (O_2244,N_28838,N_29796);
xnor UO_2245 (O_2245,N_29841,N_29001);
xnor UO_2246 (O_2246,N_29986,N_29141);
nor UO_2247 (O_2247,N_28838,N_28813);
and UO_2248 (O_2248,N_29322,N_29401);
xnor UO_2249 (O_2249,N_29007,N_28963);
nor UO_2250 (O_2250,N_29350,N_29674);
nor UO_2251 (O_2251,N_29101,N_29063);
xnor UO_2252 (O_2252,N_29906,N_29494);
or UO_2253 (O_2253,N_29931,N_28841);
and UO_2254 (O_2254,N_29228,N_28916);
nor UO_2255 (O_2255,N_29921,N_29678);
xnor UO_2256 (O_2256,N_29598,N_29239);
nand UO_2257 (O_2257,N_29898,N_29308);
or UO_2258 (O_2258,N_29433,N_29207);
and UO_2259 (O_2259,N_28906,N_29423);
nor UO_2260 (O_2260,N_29963,N_29595);
nand UO_2261 (O_2261,N_29048,N_29076);
nand UO_2262 (O_2262,N_29091,N_29803);
nor UO_2263 (O_2263,N_28851,N_29802);
nor UO_2264 (O_2264,N_29624,N_29667);
xor UO_2265 (O_2265,N_28801,N_29499);
or UO_2266 (O_2266,N_28890,N_29137);
nand UO_2267 (O_2267,N_29180,N_28939);
nand UO_2268 (O_2268,N_29636,N_29813);
and UO_2269 (O_2269,N_29680,N_28914);
nor UO_2270 (O_2270,N_29326,N_29621);
and UO_2271 (O_2271,N_29588,N_29273);
nor UO_2272 (O_2272,N_29478,N_29630);
or UO_2273 (O_2273,N_29411,N_29443);
or UO_2274 (O_2274,N_29814,N_29165);
xnor UO_2275 (O_2275,N_29299,N_29961);
xnor UO_2276 (O_2276,N_29831,N_29988);
xor UO_2277 (O_2277,N_28944,N_29313);
xnor UO_2278 (O_2278,N_29775,N_29611);
xor UO_2279 (O_2279,N_29258,N_29381);
or UO_2280 (O_2280,N_29502,N_29248);
or UO_2281 (O_2281,N_29311,N_29098);
and UO_2282 (O_2282,N_29641,N_29007);
or UO_2283 (O_2283,N_29940,N_28902);
nor UO_2284 (O_2284,N_29757,N_28815);
and UO_2285 (O_2285,N_29267,N_29603);
or UO_2286 (O_2286,N_29989,N_28937);
or UO_2287 (O_2287,N_29345,N_29109);
or UO_2288 (O_2288,N_29328,N_29191);
nor UO_2289 (O_2289,N_29739,N_28896);
or UO_2290 (O_2290,N_29482,N_28948);
or UO_2291 (O_2291,N_29849,N_29140);
nor UO_2292 (O_2292,N_28902,N_29888);
xor UO_2293 (O_2293,N_29578,N_29375);
nor UO_2294 (O_2294,N_29808,N_29399);
xnor UO_2295 (O_2295,N_29047,N_28821);
xnor UO_2296 (O_2296,N_29055,N_29535);
nand UO_2297 (O_2297,N_29176,N_28903);
or UO_2298 (O_2298,N_29517,N_29118);
nand UO_2299 (O_2299,N_29284,N_29695);
nor UO_2300 (O_2300,N_28948,N_29706);
nor UO_2301 (O_2301,N_29885,N_29356);
nand UO_2302 (O_2302,N_29306,N_29717);
nand UO_2303 (O_2303,N_29792,N_28932);
xnor UO_2304 (O_2304,N_29700,N_29303);
xnor UO_2305 (O_2305,N_29485,N_28866);
or UO_2306 (O_2306,N_29817,N_29397);
nand UO_2307 (O_2307,N_29582,N_29680);
nand UO_2308 (O_2308,N_29996,N_29589);
and UO_2309 (O_2309,N_29567,N_29476);
xnor UO_2310 (O_2310,N_28956,N_28854);
nor UO_2311 (O_2311,N_29271,N_28800);
nand UO_2312 (O_2312,N_29452,N_29096);
nor UO_2313 (O_2313,N_29804,N_28861);
nor UO_2314 (O_2314,N_28876,N_29515);
nand UO_2315 (O_2315,N_29066,N_29064);
and UO_2316 (O_2316,N_29916,N_29002);
nand UO_2317 (O_2317,N_29228,N_29731);
nand UO_2318 (O_2318,N_29514,N_29648);
nor UO_2319 (O_2319,N_29826,N_29090);
or UO_2320 (O_2320,N_29328,N_29855);
or UO_2321 (O_2321,N_28869,N_29544);
nor UO_2322 (O_2322,N_28902,N_28822);
or UO_2323 (O_2323,N_29660,N_29362);
and UO_2324 (O_2324,N_28846,N_29907);
nand UO_2325 (O_2325,N_29373,N_28842);
or UO_2326 (O_2326,N_29327,N_29434);
nand UO_2327 (O_2327,N_29922,N_28848);
or UO_2328 (O_2328,N_29087,N_29433);
and UO_2329 (O_2329,N_29314,N_29972);
and UO_2330 (O_2330,N_29994,N_29135);
xor UO_2331 (O_2331,N_29168,N_29465);
nor UO_2332 (O_2332,N_29848,N_29391);
nor UO_2333 (O_2333,N_29495,N_29063);
or UO_2334 (O_2334,N_28827,N_28861);
xnor UO_2335 (O_2335,N_29429,N_29916);
xor UO_2336 (O_2336,N_29055,N_29526);
or UO_2337 (O_2337,N_29947,N_28836);
nor UO_2338 (O_2338,N_28887,N_29565);
nor UO_2339 (O_2339,N_29432,N_29324);
xor UO_2340 (O_2340,N_29293,N_29588);
or UO_2341 (O_2341,N_29146,N_29852);
or UO_2342 (O_2342,N_29812,N_29258);
and UO_2343 (O_2343,N_29632,N_29402);
nand UO_2344 (O_2344,N_29010,N_29210);
or UO_2345 (O_2345,N_29442,N_29605);
nor UO_2346 (O_2346,N_29958,N_29393);
xnor UO_2347 (O_2347,N_29716,N_29660);
nor UO_2348 (O_2348,N_29951,N_29944);
nand UO_2349 (O_2349,N_29094,N_29309);
xor UO_2350 (O_2350,N_29161,N_29133);
nand UO_2351 (O_2351,N_29549,N_28813);
and UO_2352 (O_2352,N_28956,N_29113);
or UO_2353 (O_2353,N_29245,N_29971);
nand UO_2354 (O_2354,N_29012,N_29383);
and UO_2355 (O_2355,N_29763,N_29378);
and UO_2356 (O_2356,N_29139,N_29759);
or UO_2357 (O_2357,N_28830,N_29712);
xnor UO_2358 (O_2358,N_29453,N_28927);
and UO_2359 (O_2359,N_29618,N_29114);
and UO_2360 (O_2360,N_29244,N_28889);
or UO_2361 (O_2361,N_29488,N_28800);
nand UO_2362 (O_2362,N_29525,N_29603);
xor UO_2363 (O_2363,N_29126,N_29571);
nor UO_2364 (O_2364,N_28975,N_29086);
and UO_2365 (O_2365,N_29775,N_29904);
or UO_2366 (O_2366,N_29073,N_29158);
and UO_2367 (O_2367,N_29176,N_29197);
and UO_2368 (O_2368,N_29281,N_29002);
nor UO_2369 (O_2369,N_29535,N_29778);
nand UO_2370 (O_2370,N_28935,N_29394);
nor UO_2371 (O_2371,N_29997,N_29504);
nand UO_2372 (O_2372,N_29650,N_29112);
xnor UO_2373 (O_2373,N_28928,N_29075);
or UO_2374 (O_2374,N_29051,N_28800);
or UO_2375 (O_2375,N_29179,N_29257);
xor UO_2376 (O_2376,N_28845,N_29105);
nor UO_2377 (O_2377,N_29658,N_29033);
or UO_2378 (O_2378,N_28867,N_29982);
and UO_2379 (O_2379,N_29658,N_29228);
and UO_2380 (O_2380,N_28997,N_29241);
nand UO_2381 (O_2381,N_29307,N_29850);
and UO_2382 (O_2382,N_29447,N_29701);
nor UO_2383 (O_2383,N_29417,N_29422);
and UO_2384 (O_2384,N_29099,N_29050);
nand UO_2385 (O_2385,N_29845,N_29701);
nand UO_2386 (O_2386,N_28849,N_29339);
xnor UO_2387 (O_2387,N_29932,N_29619);
xor UO_2388 (O_2388,N_29435,N_29792);
xnor UO_2389 (O_2389,N_28996,N_29005);
or UO_2390 (O_2390,N_29285,N_29996);
and UO_2391 (O_2391,N_29039,N_28868);
and UO_2392 (O_2392,N_29826,N_29108);
nor UO_2393 (O_2393,N_29085,N_29517);
nor UO_2394 (O_2394,N_28809,N_29259);
and UO_2395 (O_2395,N_29554,N_28965);
and UO_2396 (O_2396,N_29934,N_29334);
nand UO_2397 (O_2397,N_29255,N_29810);
nor UO_2398 (O_2398,N_29649,N_29921);
xor UO_2399 (O_2399,N_29831,N_29630);
nor UO_2400 (O_2400,N_29939,N_29882);
or UO_2401 (O_2401,N_29980,N_29177);
xnor UO_2402 (O_2402,N_29312,N_29770);
or UO_2403 (O_2403,N_29170,N_29399);
xor UO_2404 (O_2404,N_29747,N_28832);
nor UO_2405 (O_2405,N_29772,N_29845);
nand UO_2406 (O_2406,N_29629,N_28948);
and UO_2407 (O_2407,N_29960,N_29070);
and UO_2408 (O_2408,N_29932,N_29104);
and UO_2409 (O_2409,N_29758,N_28851);
and UO_2410 (O_2410,N_29759,N_29877);
nor UO_2411 (O_2411,N_28854,N_29362);
xnor UO_2412 (O_2412,N_29313,N_28968);
xnor UO_2413 (O_2413,N_28906,N_29703);
nand UO_2414 (O_2414,N_29620,N_29943);
and UO_2415 (O_2415,N_29476,N_29857);
nand UO_2416 (O_2416,N_29120,N_29174);
nand UO_2417 (O_2417,N_29051,N_29890);
or UO_2418 (O_2418,N_29869,N_29833);
and UO_2419 (O_2419,N_29591,N_29400);
or UO_2420 (O_2420,N_29674,N_29463);
or UO_2421 (O_2421,N_29642,N_29735);
or UO_2422 (O_2422,N_29280,N_29933);
nand UO_2423 (O_2423,N_29064,N_29661);
nor UO_2424 (O_2424,N_29767,N_29244);
or UO_2425 (O_2425,N_29795,N_28940);
nand UO_2426 (O_2426,N_29572,N_29712);
nand UO_2427 (O_2427,N_29709,N_29995);
and UO_2428 (O_2428,N_29532,N_29398);
nor UO_2429 (O_2429,N_29121,N_29532);
xor UO_2430 (O_2430,N_29511,N_29245);
xor UO_2431 (O_2431,N_29752,N_29311);
and UO_2432 (O_2432,N_29255,N_28923);
and UO_2433 (O_2433,N_28916,N_29554);
nand UO_2434 (O_2434,N_29545,N_29715);
nor UO_2435 (O_2435,N_29776,N_29004);
nand UO_2436 (O_2436,N_29913,N_29681);
nand UO_2437 (O_2437,N_29328,N_29689);
nand UO_2438 (O_2438,N_29039,N_29403);
or UO_2439 (O_2439,N_29991,N_29657);
xor UO_2440 (O_2440,N_29060,N_29842);
nand UO_2441 (O_2441,N_28979,N_29856);
nor UO_2442 (O_2442,N_28877,N_29436);
nor UO_2443 (O_2443,N_29014,N_29815);
or UO_2444 (O_2444,N_29139,N_29461);
or UO_2445 (O_2445,N_29457,N_29864);
and UO_2446 (O_2446,N_29342,N_29272);
and UO_2447 (O_2447,N_29849,N_29251);
xnor UO_2448 (O_2448,N_29148,N_29950);
nand UO_2449 (O_2449,N_29334,N_29510);
and UO_2450 (O_2450,N_29406,N_29354);
nor UO_2451 (O_2451,N_29740,N_29216);
xnor UO_2452 (O_2452,N_28924,N_29966);
xnor UO_2453 (O_2453,N_29730,N_29694);
nand UO_2454 (O_2454,N_29126,N_29572);
or UO_2455 (O_2455,N_28987,N_29999);
nand UO_2456 (O_2456,N_29051,N_29447);
xnor UO_2457 (O_2457,N_29901,N_29475);
nand UO_2458 (O_2458,N_29319,N_28833);
and UO_2459 (O_2459,N_29694,N_29851);
nand UO_2460 (O_2460,N_29471,N_29908);
nor UO_2461 (O_2461,N_29114,N_29613);
xnor UO_2462 (O_2462,N_29101,N_29797);
nor UO_2463 (O_2463,N_29583,N_29269);
or UO_2464 (O_2464,N_29161,N_29114);
xnor UO_2465 (O_2465,N_29344,N_29637);
and UO_2466 (O_2466,N_29729,N_29142);
nor UO_2467 (O_2467,N_29185,N_29943);
xor UO_2468 (O_2468,N_28881,N_28854);
nand UO_2469 (O_2469,N_29517,N_29167);
xnor UO_2470 (O_2470,N_29906,N_28887);
nand UO_2471 (O_2471,N_29118,N_28865);
nor UO_2472 (O_2472,N_29482,N_29804);
and UO_2473 (O_2473,N_29894,N_29049);
xor UO_2474 (O_2474,N_29990,N_29035);
nor UO_2475 (O_2475,N_29328,N_29834);
or UO_2476 (O_2476,N_29716,N_28916);
nand UO_2477 (O_2477,N_29296,N_29727);
and UO_2478 (O_2478,N_29205,N_29793);
and UO_2479 (O_2479,N_29916,N_29550);
nor UO_2480 (O_2480,N_29014,N_29952);
nor UO_2481 (O_2481,N_29283,N_28932);
xnor UO_2482 (O_2482,N_29205,N_29593);
and UO_2483 (O_2483,N_29717,N_29598);
and UO_2484 (O_2484,N_29285,N_29848);
xnor UO_2485 (O_2485,N_29025,N_29149);
or UO_2486 (O_2486,N_29652,N_29993);
and UO_2487 (O_2487,N_29612,N_29510);
nor UO_2488 (O_2488,N_29445,N_29000);
or UO_2489 (O_2489,N_29222,N_29112);
or UO_2490 (O_2490,N_28811,N_29791);
nand UO_2491 (O_2491,N_29673,N_29785);
nor UO_2492 (O_2492,N_29079,N_29873);
and UO_2493 (O_2493,N_28873,N_29371);
xnor UO_2494 (O_2494,N_29447,N_29276);
and UO_2495 (O_2495,N_28824,N_29076);
xor UO_2496 (O_2496,N_29826,N_28888);
nor UO_2497 (O_2497,N_29897,N_29926);
or UO_2498 (O_2498,N_29632,N_29798);
or UO_2499 (O_2499,N_29190,N_29200);
xor UO_2500 (O_2500,N_29078,N_29845);
or UO_2501 (O_2501,N_29039,N_29495);
nor UO_2502 (O_2502,N_29209,N_29280);
and UO_2503 (O_2503,N_29518,N_28861);
nor UO_2504 (O_2504,N_28925,N_29511);
or UO_2505 (O_2505,N_29514,N_29328);
xnor UO_2506 (O_2506,N_29557,N_29383);
nor UO_2507 (O_2507,N_29519,N_29945);
and UO_2508 (O_2508,N_29177,N_29368);
or UO_2509 (O_2509,N_29320,N_29009);
xnor UO_2510 (O_2510,N_29050,N_29677);
xnor UO_2511 (O_2511,N_29119,N_29754);
xor UO_2512 (O_2512,N_29154,N_29152);
and UO_2513 (O_2513,N_29169,N_29322);
or UO_2514 (O_2514,N_29267,N_29301);
and UO_2515 (O_2515,N_29939,N_29753);
or UO_2516 (O_2516,N_28917,N_29754);
xnor UO_2517 (O_2517,N_29312,N_29425);
and UO_2518 (O_2518,N_29830,N_29465);
or UO_2519 (O_2519,N_28880,N_29338);
nand UO_2520 (O_2520,N_28975,N_29312);
xnor UO_2521 (O_2521,N_28893,N_29839);
or UO_2522 (O_2522,N_29041,N_29159);
and UO_2523 (O_2523,N_29792,N_29032);
xor UO_2524 (O_2524,N_29403,N_28945);
nand UO_2525 (O_2525,N_29317,N_29018);
or UO_2526 (O_2526,N_29394,N_29064);
and UO_2527 (O_2527,N_29502,N_29114);
xnor UO_2528 (O_2528,N_28964,N_29448);
xor UO_2529 (O_2529,N_29440,N_29474);
or UO_2530 (O_2530,N_29428,N_28928);
xor UO_2531 (O_2531,N_28865,N_28930);
nand UO_2532 (O_2532,N_29496,N_29329);
nor UO_2533 (O_2533,N_29033,N_29070);
nor UO_2534 (O_2534,N_29053,N_29696);
or UO_2535 (O_2535,N_28857,N_28957);
and UO_2536 (O_2536,N_29643,N_29719);
and UO_2537 (O_2537,N_29003,N_28985);
xor UO_2538 (O_2538,N_29131,N_29670);
nand UO_2539 (O_2539,N_29070,N_29112);
xor UO_2540 (O_2540,N_29909,N_28878);
and UO_2541 (O_2541,N_28832,N_29648);
and UO_2542 (O_2542,N_29688,N_29092);
nand UO_2543 (O_2543,N_29878,N_29734);
or UO_2544 (O_2544,N_29857,N_29839);
or UO_2545 (O_2545,N_29719,N_29708);
and UO_2546 (O_2546,N_29663,N_29809);
nor UO_2547 (O_2547,N_29627,N_28865);
or UO_2548 (O_2548,N_29995,N_29758);
nor UO_2549 (O_2549,N_29260,N_29785);
and UO_2550 (O_2550,N_28920,N_29201);
or UO_2551 (O_2551,N_29753,N_28975);
and UO_2552 (O_2552,N_29625,N_29805);
nor UO_2553 (O_2553,N_29972,N_29704);
and UO_2554 (O_2554,N_28994,N_29841);
nor UO_2555 (O_2555,N_29435,N_29682);
or UO_2556 (O_2556,N_29662,N_29927);
and UO_2557 (O_2557,N_29840,N_29694);
and UO_2558 (O_2558,N_29383,N_29058);
and UO_2559 (O_2559,N_29794,N_29488);
nand UO_2560 (O_2560,N_29188,N_29415);
and UO_2561 (O_2561,N_29735,N_29058);
xor UO_2562 (O_2562,N_28940,N_29439);
nor UO_2563 (O_2563,N_29341,N_28887);
and UO_2564 (O_2564,N_29257,N_29315);
nor UO_2565 (O_2565,N_29691,N_29043);
or UO_2566 (O_2566,N_29943,N_29773);
or UO_2567 (O_2567,N_29795,N_29539);
nand UO_2568 (O_2568,N_29643,N_29390);
or UO_2569 (O_2569,N_28929,N_29152);
nand UO_2570 (O_2570,N_29326,N_29947);
or UO_2571 (O_2571,N_29786,N_29724);
xnor UO_2572 (O_2572,N_29393,N_28983);
xnor UO_2573 (O_2573,N_29672,N_28967);
or UO_2574 (O_2574,N_29178,N_28913);
xor UO_2575 (O_2575,N_29857,N_29669);
xor UO_2576 (O_2576,N_29939,N_29120);
or UO_2577 (O_2577,N_29126,N_28994);
nor UO_2578 (O_2578,N_29701,N_29404);
nor UO_2579 (O_2579,N_29955,N_29979);
nor UO_2580 (O_2580,N_29905,N_28821);
nor UO_2581 (O_2581,N_29967,N_29348);
xor UO_2582 (O_2582,N_29745,N_29547);
nor UO_2583 (O_2583,N_29757,N_28842);
and UO_2584 (O_2584,N_29211,N_29813);
nand UO_2585 (O_2585,N_29463,N_28975);
and UO_2586 (O_2586,N_29910,N_29235);
and UO_2587 (O_2587,N_29574,N_29602);
nand UO_2588 (O_2588,N_29703,N_28875);
and UO_2589 (O_2589,N_28987,N_29046);
nor UO_2590 (O_2590,N_29494,N_29238);
nand UO_2591 (O_2591,N_29177,N_29652);
or UO_2592 (O_2592,N_29022,N_29651);
and UO_2593 (O_2593,N_29940,N_29797);
xnor UO_2594 (O_2594,N_29685,N_29711);
or UO_2595 (O_2595,N_29111,N_29588);
nand UO_2596 (O_2596,N_28906,N_29739);
nand UO_2597 (O_2597,N_29340,N_29969);
nand UO_2598 (O_2598,N_29979,N_29592);
xor UO_2599 (O_2599,N_29640,N_29010);
nor UO_2600 (O_2600,N_29456,N_29149);
and UO_2601 (O_2601,N_29187,N_29246);
xnor UO_2602 (O_2602,N_29094,N_29666);
nand UO_2603 (O_2603,N_28940,N_29171);
or UO_2604 (O_2604,N_29930,N_29265);
or UO_2605 (O_2605,N_29832,N_29483);
nor UO_2606 (O_2606,N_29402,N_29588);
or UO_2607 (O_2607,N_29541,N_28848);
and UO_2608 (O_2608,N_29839,N_29203);
nand UO_2609 (O_2609,N_28974,N_29575);
xor UO_2610 (O_2610,N_28928,N_29979);
xor UO_2611 (O_2611,N_29101,N_29341);
or UO_2612 (O_2612,N_28846,N_29212);
and UO_2613 (O_2613,N_29324,N_29930);
nand UO_2614 (O_2614,N_29183,N_29138);
xnor UO_2615 (O_2615,N_28819,N_29225);
nand UO_2616 (O_2616,N_29172,N_29066);
nor UO_2617 (O_2617,N_29502,N_29665);
nor UO_2618 (O_2618,N_29679,N_29057);
xnor UO_2619 (O_2619,N_29972,N_28829);
or UO_2620 (O_2620,N_29836,N_28819);
and UO_2621 (O_2621,N_29930,N_28879);
or UO_2622 (O_2622,N_29307,N_28902);
xnor UO_2623 (O_2623,N_29073,N_29569);
and UO_2624 (O_2624,N_28883,N_29559);
nand UO_2625 (O_2625,N_28916,N_28913);
nand UO_2626 (O_2626,N_29409,N_29010);
xnor UO_2627 (O_2627,N_29349,N_29287);
or UO_2628 (O_2628,N_28823,N_29984);
and UO_2629 (O_2629,N_29883,N_29630);
nand UO_2630 (O_2630,N_29450,N_29728);
nor UO_2631 (O_2631,N_29751,N_29750);
and UO_2632 (O_2632,N_29329,N_29147);
xnor UO_2633 (O_2633,N_29135,N_29243);
xnor UO_2634 (O_2634,N_28929,N_29048);
nand UO_2635 (O_2635,N_29541,N_29949);
or UO_2636 (O_2636,N_29853,N_29964);
nor UO_2637 (O_2637,N_29140,N_29180);
xnor UO_2638 (O_2638,N_29558,N_29918);
xor UO_2639 (O_2639,N_29152,N_29533);
xnor UO_2640 (O_2640,N_29473,N_29090);
or UO_2641 (O_2641,N_29729,N_29144);
or UO_2642 (O_2642,N_29096,N_29717);
and UO_2643 (O_2643,N_29004,N_29095);
or UO_2644 (O_2644,N_29772,N_29474);
or UO_2645 (O_2645,N_29049,N_29129);
nor UO_2646 (O_2646,N_28904,N_29135);
nor UO_2647 (O_2647,N_29381,N_29118);
xnor UO_2648 (O_2648,N_29142,N_28902);
or UO_2649 (O_2649,N_29284,N_29202);
nor UO_2650 (O_2650,N_28999,N_29618);
xor UO_2651 (O_2651,N_28848,N_29857);
and UO_2652 (O_2652,N_29286,N_29089);
nor UO_2653 (O_2653,N_29984,N_29698);
nor UO_2654 (O_2654,N_29162,N_29003);
nand UO_2655 (O_2655,N_28802,N_29376);
nand UO_2656 (O_2656,N_28818,N_29236);
or UO_2657 (O_2657,N_29752,N_29157);
and UO_2658 (O_2658,N_29680,N_29487);
nor UO_2659 (O_2659,N_29627,N_29624);
nor UO_2660 (O_2660,N_28918,N_29266);
nand UO_2661 (O_2661,N_29496,N_29778);
nor UO_2662 (O_2662,N_29998,N_29385);
and UO_2663 (O_2663,N_28897,N_29492);
nor UO_2664 (O_2664,N_29984,N_29406);
or UO_2665 (O_2665,N_29174,N_29226);
and UO_2666 (O_2666,N_28983,N_29493);
or UO_2667 (O_2667,N_29039,N_29125);
and UO_2668 (O_2668,N_29228,N_29517);
nor UO_2669 (O_2669,N_29108,N_29358);
xor UO_2670 (O_2670,N_29958,N_29044);
xor UO_2671 (O_2671,N_29833,N_28813);
and UO_2672 (O_2672,N_29859,N_29787);
or UO_2673 (O_2673,N_29448,N_29170);
nor UO_2674 (O_2674,N_29292,N_29637);
and UO_2675 (O_2675,N_28876,N_29894);
or UO_2676 (O_2676,N_29525,N_29370);
nand UO_2677 (O_2677,N_29667,N_28982);
or UO_2678 (O_2678,N_29061,N_29919);
or UO_2679 (O_2679,N_29829,N_28844);
or UO_2680 (O_2680,N_29582,N_29083);
nand UO_2681 (O_2681,N_29129,N_29528);
xnor UO_2682 (O_2682,N_29755,N_29026);
nand UO_2683 (O_2683,N_28805,N_29730);
nor UO_2684 (O_2684,N_29177,N_29492);
or UO_2685 (O_2685,N_29021,N_28808);
xor UO_2686 (O_2686,N_29548,N_29067);
or UO_2687 (O_2687,N_29841,N_29296);
nand UO_2688 (O_2688,N_29173,N_29979);
or UO_2689 (O_2689,N_29111,N_29904);
or UO_2690 (O_2690,N_29870,N_28805);
nand UO_2691 (O_2691,N_29762,N_29066);
xnor UO_2692 (O_2692,N_29105,N_29647);
xnor UO_2693 (O_2693,N_28872,N_29027);
and UO_2694 (O_2694,N_29070,N_28804);
xor UO_2695 (O_2695,N_29389,N_29975);
xor UO_2696 (O_2696,N_29108,N_29419);
xnor UO_2697 (O_2697,N_28869,N_29098);
nand UO_2698 (O_2698,N_29906,N_29916);
and UO_2699 (O_2699,N_29051,N_29594);
and UO_2700 (O_2700,N_29001,N_29410);
xor UO_2701 (O_2701,N_29324,N_29736);
and UO_2702 (O_2702,N_28844,N_29603);
nand UO_2703 (O_2703,N_29100,N_29668);
nor UO_2704 (O_2704,N_29369,N_29744);
and UO_2705 (O_2705,N_29521,N_29642);
nand UO_2706 (O_2706,N_29638,N_28841);
xor UO_2707 (O_2707,N_29064,N_29517);
xor UO_2708 (O_2708,N_28940,N_29495);
nor UO_2709 (O_2709,N_29816,N_29480);
nand UO_2710 (O_2710,N_29506,N_29571);
nor UO_2711 (O_2711,N_29334,N_29746);
xor UO_2712 (O_2712,N_29669,N_29177);
xnor UO_2713 (O_2713,N_29543,N_29338);
nand UO_2714 (O_2714,N_29827,N_29070);
xor UO_2715 (O_2715,N_29625,N_29187);
and UO_2716 (O_2716,N_28924,N_28843);
nor UO_2717 (O_2717,N_29483,N_29510);
or UO_2718 (O_2718,N_29330,N_28925);
nor UO_2719 (O_2719,N_29536,N_29137);
or UO_2720 (O_2720,N_29841,N_29825);
and UO_2721 (O_2721,N_29781,N_29461);
nand UO_2722 (O_2722,N_29549,N_29093);
and UO_2723 (O_2723,N_29516,N_29410);
or UO_2724 (O_2724,N_29012,N_29930);
xnor UO_2725 (O_2725,N_29713,N_29500);
and UO_2726 (O_2726,N_29676,N_29632);
xnor UO_2727 (O_2727,N_29347,N_29429);
xor UO_2728 (O_2728,N_29733,N_29654);
xnor UO_2729 (O_2729,N_29770,N_29825);
and UO_2730 (O_2730,N_29080,N_29757);
nor UO_2731 (O_2731,N_29132,N_29233);
and UO_2732 (O_2732,N_29266,N_29121);
nand UO_2733 (O_2733,N_29166,N_28849);
xor UO_2734 (O_2734,N_29144,N_29997);
xor UO_2735 (O_2735,N_29682,N_29055);
and UO_2736 (O_2736,N_29259,N_29970);
or UO_2737 (O_2737,N_29631,N_29238);
xnor UO_2738 (O_2738,N_29071,N_29448);
nand UO_2739 (O_2739,N_29547,N_29267);
xor UO_2740 (O_2740,N_29525,N_29512);
or UO_2741 (O_2741,N_29714,N_29328);
or UO_2742 (O_2742,N_28950,N_29454);
xnor UO_2743 (O_2743,N_28917,N_29923);
nor UO_2744 (O_2744,N_28846,N_29286);
nor UO_2745 (O_2745,N_29021,N_29404);
xor UO_2746 (O_2746,N_29542,N_29794);
or UO_2747 (O_2747,N_29871,N_29007);
nor UO_2748 (O_2748,N_29164,N_29225);
nor UO_2749 (O_2749,N_28976,N_29721);
nor UO_2750 (O_2750,N_29755,N_29060);
xnor UO_2751 (O_2751,N_28851,N_28854);
or UO_2752 (O_2752,N_28815,N_29365);
nand UO_2753 (O_2753,N_29273,N_29809);
nand UO_2754 (O_2754,N_29434,N_29142);
nand UO_2755 (O_2755,N_29433,N_29239);
xnor UO_2756 (O_2756,N_29609,N_28866);
or UO_2757 (O_2757,N_29285,N_29871);
nand UO_2758 (O_2758,N_29628,N_29464);
and UO_2759 (O_2759,N_29973,N_29229);
nor UO_2760 (O_2760,N_29194,N_29722);
xnor UO_2761 (O_2761,N_29197,N_28958);
or UO_2762 (O_2762,N_29801,N_29297);
nor UO_2763 (O_2763,N_29908,N_29414);
nor UO_2764 (O_2764,N_29890,N_29869);
or UO_2765 (O_2765,N_29500,N_29600);
nor UO_2766 (O_2766,N_28920,N_29050);
or UO_2767 (O_2767,N_29035,N_29498);
and UO_2768 (O_2768,N_29560,N_29358);
or UO_2769 (O_2769,N_29223,N_29610);
and UO_2770 (O_2770,N_28986,N_29762);
nor UO_2771 (O_2771,N_29393,N_29912);
or UO_2772 (O_2772,N_28988,N_29002);
or UO_2773 (O_2773,N_29754,N_29168);
xor UO_2774 (O_2774,N_29973,N_29915);
nor UO_2775 (O_2775,N_29021,N_29263);
or UO_2776 (O_2776,N_29627,N_29024);
nor UO_2777 (O_2777,N_28854,N_29746);
or UO_2778 (O_2778,N_29521,N_29660);
xnor UO_2779 (O_2779,N_28918,N_29123);
or UO_2780 (O_2780,N_29669,N_29346);
xnor UO_2781 (O_2781,N_29847,N_29639);
and UO_2782 (O_2782,N_29648,N_29188);
and UO_2783 (O_2783,N_29599,N_29443);
nand UO_2784 (O_2784,N_29800,N_29021);
xnor UO_2785 (O_2785,N_29219,N_28938);
nand UO_2786 (O_2786,N_29284,N_29525);
nor UO_2787 (O_2787,N_28851,N_29039);
or UO_2788 (O_2788,N_29791,N_29330);
and UO_2789 (O_2789,N_29171,N_29188);
and UO_2790 (O_2790,N_29104,N_29847);
nand UO_2791 (O_2791,N_29142,N_29430);
or UO_2792 (O_2792,N_29861,N_29574);
and UO_2793 (O_2793,N_29552,N_29794);
or UO_2794 (O_2794,N_29054,N_29463);
nand UO_2795 (O_2795,N_29908,N_29809);
xor UO_2796 (O_2796,N_29940,N_29175);
nor UO_2797 (O_2797,N_29120,N_29374);
nor UO_2798 (O_2798,N_28924,N_29655);
nand UO_2799 (O_2799,N_29110,N_29879);
nor UO_2800 (O_2800,N_29454,N_29125);
xor UO_2801 (O_2801,N_28857,N_29491);
nor UO_2802 (O_2802,N_29728,N_29855);
nand UO_2803 (O_2803,N_28999,N_29151);
nand UO_2804 (O_2804,N_28838,N_29780);
and UO_2805 (O_2805,N_29822,N_28872);
and UO_2806 (O_2806,N_29777,N_29134);
or UO_2807 (O_2807,N_29697,N_29612);
and UO_2808 (O_2808,N_29064,N_29009);
or UO_2809 (O_2809,N_29553,N_29515);
nand UO_2810 (O_2810,N_29604,N_29877);
xnor UO_2811 (O_2811,N_28939,N_29425);
nor UO_2812 (O_2812,N_29079,N_29880);
nor UO_2813 (O_2813,N_29520,N_29482);
xnor UO_2814 (O_2814,N_28820,N_29722);
xnor UO_2815 (O_2815,N_28967,N_29451);
nand UO_2816 (O_2816,N_29783,N_29078);
xor UO_2817 (O_2817,N_29060,N_29651);
and UO_2818 (O_2818,N_29227,N_29192);
xnor UO_2819 (O_2819,N_29664,N_28902);
nand UO_2820 (O_2820,N_29959,N_29644);
xnor UO_2821 (O_2821,N_28852,N_29324);
nand UO_2822 (O_2822,N_29625,N_29559);
nand UO_2823 (O_2823,N_29692,N_29355);
nand UO_2824 (O_2824,N_29463,N_29959);
xor UO_2825 (O_2825,N_29965,N_29148);
nand UO_2826 (O_2826,N_29919,N_28883);
xnor UO_2827 (O_2827,N_29487,N_29237);
nand UO_2828 (O_2828,N_29160,N_29729);
xnor UO_2829 (O_2829,N_29515,N_29570);
and UO_2830 (O_2830,N_29847,N_29411);
or UO_2831 (O_2831,N_29758,N_29767);
and UO_2832 (O_2832,N_29499,N_28982);
xnor UO_2833 (O_2833,N_29210,N_29480);
nand UO_2834 (O_2834,N_29254,N_28846);
or UO_2835 (O_2835,N_29957,N_29439);
nor UO_2836 (O_2836,N_29737,N_28939);
nor UO_2837 (O_2837,N_28837,N_28957);
nand UO_2838 (O_2838,N_29869,N_28829);
nand UO_2839 (O_2839,N_29838,N_29918);
nor UO_2840 (O_2840,N_29996,N_29502);
nor UO_2841 (O_2841,N_29257,N_29533);
nand UO_2842 (O_2842,N_29644,N_28849);
xor UO_2843 (O_2843,N_28839,N_29353);
and UO_2844 (O_2844,N_29276,N_29683);
or UO_2845 (O_2845,N_29094,N_29059);
or UO_2846 (O_2846,N_29239,N_29491);
and UO_2847 (O_2847,N_29106,N_29738);
and UO_2848 (O_2848,N_29589,N_29193);
and UO_2849 (O_2849,N_29480,N_29700);
and UO_2850 (O_2850,N_29291,N_29226);
xnor UO_2851 (O_2851,N_28932,N_29073);
nor UO_2852 (O_2852,N_29370,N_29256);
or UO_2853 (O_2853,N_29735,N_28956);
nor UO_2854 (O_2854,N_29525,N_28832);
or UO_2855 (O_2855,N_29780,N_28971);
nand UO_2856 (O_2856,N_29597,N_29524);
or UO_2857 (O_2857,N_29620,N_29203);
xnor UO_2858 (O_2858,N_29360,N_29436);
nor UO_2859 (O_2859,N_29166,N_28930);
nor UO_2860 (O_2860,N_29295,N_29795);
or UO_2861 (O_2861,N_29743,N_29343);
or UO_2862 (O_2862,N_29369,N_29472);
nand UO_2863 (O_2863,N_29279,N_29712);
and UO_2864 (O_2864,N_28949,N_29260);
xnor UO_2865 (O_2865,N_28825,N_29458);
or UO_2866 (O_2866,N_29508,N_29231);
xnor UO_2867 (O_2867,N_28910,N_29406);
nor UO_2868 (O_2868,N_29767,N_29920);
nand UO_2869 (O_2869,N_29913,N_29300);
nor UO_2870 (O_2870,N_29147,N_29387);
nand UO_2871 (O_2871,N_28846,N_29831);
and UO_2872 (O_2872,N_28858,N_28953);
nor UO_2873 (O_2873,N_29664,N_29059);
nand UO_2874 (O_2874,N_28840,N_29120);
or UO_2875 (O_2875,N_29592,N_29376);
xnor UO_2876 (O_2876,N_29571,N_29056);
or UO_2877 (O_2877,N_29795,N_29840);
and UO_2878 (O_2878,N_29162,N_29731);
or UO_2879 (O_2879,N_29854,N_29494);
or UO_2880 (O_2880,N_29904,N_29038);
and UO_2881 (O_2881,N_28917,N_29879);
nor UO_2882 (O_2882,N_29859,N_29019);
nand UO_2883 (O_2883,N_29743,N_29994);
or UO_2884 (O_2884,N_28807,N_28830);
or UO_2885 (O_2885,N_29653,N_28894);
xor UO_2886 (O_2886,N_29773,N_29217);
nand UO_2887 (O_2887,N_29608,N_29451);
or UO_2888 (O_2888,N_29721,N_28908);
nand UO_2889 (O_2889,N_29649,N_29006);
or UO_2890 (O_2890,N_29223,N_29636);
and UO_2891 (O_2891,N_29083,N_29439);
xnor UO_2892 (O_2892,N_29577,N_29275);
xnor UO_2893 (O_2893,N_29792,N_28978);
and UO_2894 (O_2894,N_29298,N_29406);
xor UO_2895 (O_2895,N_29174,N_28917);
and UO_2896 (O_2896,N_29697,N_29365);
and UO_2897 (O_2897,N_28815,N_29499);
xnor UO_2898 (O_2898,N_29425,N_29499);
xor UO_2899 (O_2899,N_29840,N_29350);
and UO_2900 (O_2900,N_29386,N_29714);
nor UO_2901 (O_2901,N_28964,N_29749);
or UO_2902 (O_2902,N_29102,N_29280);
nor UO_2903 (O_2903,N_29749,N_29794);
xor UO_2904 (O_2904,N_29256,N_29379);
nor UO_2905 (O_2905,N_29896,N_29939);
and UO_2906 (O_2906,N_29558,N_28829);
and UO_2907 (O_2907,N_28995,N_29115);
and UO_2908 (O_2908,N_28801,N_29968);
or UO_2909 (O_2909,N_28957,N_28800);
xnor UO_2910 (O_2910,N_29454,N_29991);
nor UO_2911 (O_2911,N_29618,N_29875);
and UO_2912 (O_2912,N_29792,N_29305);
xor UO_2913 (O_2913,N_29398,N_29613);
xnor UO_2914 (O_2914,N_29016,N_28946);
nor UO_2915 (O_2915,N_29118,N_29743);
or UO_2916 (O_2916,N_29955,N_28805);
or UO_2917 (O_2917,N_29907,N_29088);
nand UO_2918 (O_2918,N_29161,N_29751);
xnor UO_2919 (O_2919,N_29259,N_28858);
and UO_2920 (O_2920,N_29531,N_28803);
xor UO_2921 (O_2921,N_29882,N_29520);
xor UO_2922 (O_2922,N_29951,N_29895);
and UO_2923 (O_2923,N_29180,N_29328);
nor UO_2924 (O_2924,N_29416,N_29812);
nand UO_2925 (O_2925,N_29402,N_29273);
or UO_2926 (O_2926,N_29699,N_29507);
xor UO_2927 (O_2927,N_29115,N_29914);
or UO_2928 (O_2928,N_28813,N_29864);
xnor UO_2929 (O_2929,N_29714,N_29663);
nor UO_2930 (O_2930,N_29955,N_29069);
xor UO_2931 (O_2931,N_29956,N_29903);
nor UO_2932 (O_2932,N_28940,N_29754);
nor UO_2933 (O_2933,N_28817,N_29760);
xor UO_2934 (O_2934,N_29066,N_29038);
and UO_2935 (O_2935,N_29569,N_29667);
xnor UO_2936 (O_2936,N_29580,N_29727);
nand UO_2937 (O_2937,N_28880,N_29775);
xnor UO_2938 (O_2938,N_29178,N_29855);
nor UO_2939 (O_2939,N_28904,N_29194);
nand UO_2940 (O_2940,N_29137,N_29273);
nor UO_2941 (O_2941,N_29910,N_29155);
or UO_2942 (O_2942,N_29922,N_29212);
xnor UO_2943 (O_2943,N_29383,N_29097);
nor UO_2944 (O_2944,N_29192,N_29675);
or UO_2945 (O_2945,N_29033,N_29068);
or UO_2946 (O_2946,N_29508,N_29913);
nor UO_2947 (O_2947,N_28962,N_29218);
nand UO_2948 (O_2948,N_29371,N_29053);
xor UO_2949 (O_2949,N_29339,N_28845);
xnor UO_2950 (O_2950,N_29034,N_28925);
and UO_2951 (O_2951,N_29683,N_28907);
and UO_2952 (O_2952,N_29757,N_29130);
nor UO_2953 (O_2953,N_29832,N_29699);
or UO_2954 (O_2954,N_29563,N_29402);
nor UO_2955 (O_2955,N_28927,N_29218);
or UO_2956 (O_2956,N_29110,N_29725);
or UO_2957 (O_2957,N_29058,N_29033);
and UO_2958 (O_2958,N_28888,N_29660);
and UO_2959 (O_2959,N_29030,N_29672);
or UO_2960 (O_2960,N_29453,N_29107);
nor UO_2961 (O_2961,N_29385,N_29920);
xor UO_2962 (O_2962,N_29100,N_29210);
nor UO_2963 (O_2963,N_29549,N_28846);
nor UO_2964 (O_2964,N_29456,N_29442);
or UO_2965 (O_2965,N_29314,N_28900);
nand UO_2966 (O_2966,N_28871,N_29004);
xnor UO_2967 (O_2967,N_28941,N_29840);
nand UO_2968 (O_2968,N_29958,N_29527);
and UO_2969 (O_2969,N_29373,N_29356);
nor UO_2970 (O_2970,N_28965,N_29648);
and UO_2971 (O_2971,N_29579,N_28892);
and UO_2972 (O_2972,N_29273,N_28965);
nand UO_2973 (O_2973,N_29241,N_29550);
or UO_2974 (O_2974,N_29956,N_29426);
nor UO_2975 (O_2975,N_29679,N_29486);
xor UO_2976 (O_2976,N_29346,N_29211);
xnor UO_2977 (O_2977,N_29457,N_28998);
and UO_2978 (O_2978,N_29381,N_29329);
nor UO_2979 (O_2979,N_29825,N_29711);
xor UO_2980 (O_2980,N_29559,N_29129);
nand UO_2981 (O_2981,N_29960,N_29065);
and UO_2982 (O_2982,N_29046,N_29649);
and UO_2983 (O_2983,N_29722,N_29992);
nor UO_2984 (O_2984,N_29225,N_29421);
xor UO_2985 (O_2985,N_29460,N_29778);
xnor UO_2986 (O_2986,N_29240,N_29558);
nor UO_2987 (O_2987,N_29878,N_29551);
nor UO_2988 (O_2988,N_29742,N_29458);
nor UO_2989 (O_2989,N_29590,N_29417);
or UO_2990 (O_2990,N_28878,N_29111);
xor UO_2991 (O_2991,N_29828,N_29571);
nand UO_2992 (O_2992,N_29668,N_29448);
nor UO_2993 (O_2993,N_29800,N_29854);
and UO_2994 (O_2994,N_29607,N_29732);
or UO_2995 (O_2995,N_29448,N_29053);
and UO_2996 (O_2996,N_29039,N_28938);
nand UO_2997 (O_2997,N_29680,N_29848);
and UO_2998 (O_2998,N_29690,N_29715);
or UO_2999 (O_2999,N_29958,N_29015);
nor UO_3000 (O_3000,N_29197,N_29706);
xnor UO_3001 (O_3001,N_29564,N_29773);
and UO_3002 (O_3002,N_28915,N_28918);
nor UO_3003 (O_3003,N_29714,N_29005);
nor UO_3004 (O_3004,N_29768,N_28871);
or UO_3005 (O_3005,N_29148,N_29344);
or UO_3006 (O_3006,N_29119,N_29948);
or UO_3007 (O_3007,N_29902,N_29420);
and UO_3008 (O_3008,N_28822,N_29821);
or UO_3009 (O_3009,N_29113,N_28931);
nor UO_3010 (O_3010,N_29141,N_29274);
xor UO_3011 (O_3011,N_29599,N_29919);
nor UO_3012 (O_3012,N_29956,N_29793);
xor UO_3013 (O_3013,N_29937,N_29328);
nor UO_3014 (O_3014,N_29267,N_29338);
nand UO_3015 (O_3015,N_29399,N_29151);
and UO_3016 (O_3016,N_29373,N_29530);
nor UO_3017 (O_3017,N_28903,N_29457);
nor UO_3018 (O_3018,N_29985,N_29095);
nand UO_3019 (O_3019,N_28821,N_28890);
nand UO_3020 (O_3020,N_29367,N_28880);
and UO_3021 (O_3021,N_29270,N_29745);
and UO_3022 (O_3022,N_29839,N_29245);
nand UO_3023 (O_3023,N_28870,N_28853);
or UO_3024 (O_3024,N_29967,N_28986);
and UO_3025 (O_3025,N_29122,N_29137);
nand UO_3026 (O_3026,N_29239,N_29042);
nand UO_3027 (O_3027,N_28971,N_29832);
or UO_3028 (O_3028,N_29158,N_29241);
nor UO_3029 (O_3029,N_29734,N_28810);
xnor UO_3030 (O_3030,N_29952,N_29792);
or UO_3031 (O_3031,N_29999,N_29376);
or UO_3032 (O_3032,N_29616,N_29266);
and UO_3033 (O_3033,N_29084,N_29908);
and UO_3034 (O_3034,N_29832,N_28854);
nor UO_3035 (O_3035,N_28821,N_29593);
nand UO_3036 (O_3036,N_29138,N_28993);
nand UO_3037 (O_3037,N_29964,N_29648);
xnor UO_3038 (O_3038,N_29194,N_29155);
nor UO_3039 (O_3039,N_29499,N_29572);
nor UO_3040 (O_3040,N_29369,N_29745);
xor UO_3041 (O_3041,N_29064,N_28855);
xor UO_3042 (O_3042,N_28932,N_29575);
nand UO_3043 (O_3043,N_29631,N_29845);
nor UO_3044 (O_3044,N_28885,N_29939);
xor UO_3045 (O_3045,N_29396,N_29953);
nor UO_3046 (O_3046,N_28846,N_29029);
or UO_3047 (O_3047,N_29684,N_29419);
nor UO_3048 (O_3048,N_29177,N_29300);
xnor UO_3049 (O_3049,N_28889,N_29544);
or UO_3050 (O_3050,N_29894,N_28867);
xor UO_3051 (O_3051,N_29520,N_29574);
or UO_3052 (O_3052,N_28943,N_29178);
xor UO_3053 (O_3053,N_28830,N_29298);
and UO_3054 (O_3054,N_29777,N_29027);
or UO_3055 (O_3055,N_29029,N_29943);
xnor UO_3056 (O_3056,N_29616,N_29565);
or UO_3057 (O_3057,N_29458,N_29990);
nor UO_3058 (O_3058,N_29931,N_29366);
xnor UO_3059 (O_3059,N_29326,N_29597);
and UO_3060 (O_3060,N_28823,N_29291);
xor UO_3061 (O_3061,N_29282,N_28912);
nand UO_3062 (O_3062,N_29444,N_29722);
or UO_3063 (O_3063,N_29276,N_29444);
and UO_3064 (O_3064,N_29568,N_28987);
xnor UO_3065 (O_3065,N_29617,N_28951);
xnor UO_3066 (O_3066,N_28891,N_29377);
nor UO_3067 (O_3067,N_29351,N_29400);
xnor UO_3068 (O_3068,N_29256,N_29351);
xnor UO_3069 (O_3069,N_29660,N_29545);
xnor UO_3070 (O_3070,N_29253,N_29596);
nand UO_3071 (O_3071,N_29603,N_29851);
or UO_3072 (O_3072,N_29335,N_29319);
and UO_3073 (O_3073,N_29191,N_29787);
xnor UO_3074 (O_3074,N_29431,N_29174);
xnor UO_3075 (O_3075,N_29735,N_29912);
and UO_3076 (O_3076,N_29651,N_29717);
nor UO_3077 (O_3077,N_29429,N_29383);
and UO_3078 (O_3078,N_29053,N_29738);
nand UO_3079 (O_3079,N_29026,N_28860);
and UO_3080 (O_3080,N_29170,N_29390);
or UO_3081 (O_3081,N_29300,N_29696);
nand UO_3082 (O_3082,N_29201,N_29300);
xor UO_3083 (O_3083,N_29147,N_29554);
or UO_3084 (O_3084,N_29537,N_29250);
and UO_3085 (O_3085,N_29572,N_29621);
nor UO_3086 (O_3086,N_29851,N_29562);
xnor UO_3087 (O_3087,N_29756,N_29640);
nand UO_3088 (O_3088,N_29400,N_29715);
nand UO_3089 (O_3089,N_29736,N_29264);
nor UO_3090 (O_3090,N_29045,N_29077);
xor UO_3091 (O_3091,N_29241,N_29461);
and UO_3092 (O_3092,N_29724,N_29704);
xor UO_3093 (O_3093,N_29840,N_29844);
xnor UO_3094 (O_3094,N_29355,N_29581);
nand UO_3095 (O_3095,N_29027,N_29737);
nand UO_3096 (O_3096,N_29401,N_29975);
xor UO_3097 (O_3097,N_29823,N_29155);
xor UO_3098 (O_3098,N_28856,N_29988);
nor UO_3099 (O_3099,N_29399,N_29599);
or UO_3100 (O_3100,N_29140,N_28946);
nand UO_3101 (O_3101,N_29287,N_29771);
and UO_3102 (O_3102,N_29440,N_28920);
nor UO_3103 (O_3103,N_29682,N_29649);
or UO_3104 (O_3104,N_28815,N_29948);
and UO_3105 (O_3105,N_29763,N_29418);
and UO_3106 (O_3106,N_29795,N_29334);
nand UO_3107 (O_3107,N_29163,N_29150);
or UO_3108 (O_3108,N_29013,N_29185);
xor UO_3109 (O_3109,N_29318,N_29248);
and UO_3110 (O_3110,N_28838,N_29596);
nor UO_3111 (O_3111,N_29081,N_28873);
xor UO_3112 (O_3112,N_29419,N_29380);
nand UO_3113 (O_3113,N_29925,N_29230);
or UO_3114 (O_3114,N_29785,N_28845);
or UO_3115 (O_3115,N_29455,N_29469);
nor UO_3116 (O_3116,N_29535,N_29146);
nor UO_3117 (O_3117,N_29483,N_29057);
and UO_3118 (O_3118,N_29047,N_29297);
xor UO_3119 (O_3119,N_28834,N_29998);
xnor UO_3120 (O_3120,N_29153,N_29997);
or UO_3121 (O_3121,N_29955,N_29697);
or UO_3122 (O_3122,N_29590,N_29613);
nor UO_3123 (O_3123,N_29610,N_28888);
nor UO_3124 (O_3124,N_29113,N_28990);
and UO_3125 (O_3125,N_29978,N_29937);
xnor UO_3126 (O_3126,N_28948,N_29357);
and UO_3127 (O_3127,N_29944,N_29860);
xor UO_3128 (O_3128,N_29477,N_29257);
xor UO_3129 (O_3129,N_29438,N_29459);
or UO_3130 (O_3130,N_29078,N_29820);
and UO_3131 (O_3131,N_29418,N_29372);
xor UO_3132 (O_3132,N_29461,N_29062);
nand UO_3133 (O_3133,N_29597,N_28938);
and UO_3134 (O_3134,N_29576,N_28923);
nand UO_3135 (O_3135,N_29660,N_29171);
and UO_3136 (O_3136,N_29104,N_29669);
nor UO_3137 (O_3137,N_28962,N_29830);
xor UO_3138 (O_3138,N_29349,N_28904);
xnor UO_3139 (O_3139,N_29689,N_29683);
xor UO_3140 (O_3140,N_28809,N_29674);
or UO_3141 (O_3141,N_29225,N_29067);
and UO_3142 (O_3142,N_29327,N_29779);
or UO_3143 (O_3143,N_29879,N_29612);
or UO_3144 (O_3144,N_29130,N_29209);
and UO_3145 (O_3145,N_28901,N_29531);
or UO_3146 (O_3146,N_29013,N_28994);
and UO_3147 (O_3147,N_29150,N_29566);
nor UO_3148 (O_3148,N_29287,N_29280);
and UO_3149 (O_3149,N_29249,N_29207);
and UO_3150 (O_3150,N_29898,N_29105);
and UO_3151 (O_3151,N_29699,N_28855);
xnor UO_3152 (O_3152,N_29120,N_29348);
nor UO_3153 (O_3153,N_29878,N_29701);
nand UO_3154 (O_3154,N_29216,N_29729);
and UO_3155 (O_3155,N_28989,N_29559);
and UO_3156 (O_3156,N_29516,N_29807);
or UO_3157 (O_3157,N_28986,N_29873);
nand UO_3158 (O_3158,N_28880,N_29990);
xnor UO_3159 (O_3159,N_29482,N_29785);
and UO_3160 (O_3160,N_29200,N_29969);
nand UO_3161 (O_3161,N_29080,N_29256);
and UO_3162 (O_3162,N_29435,N_29139);
or UO_3163 (O_3163,N_29536,N_29841);
and UO_3164 (O_3164,N_29488,N_29629);
and UO_3165 (O_3165,N_29571,N_29030);
and UO_3166 (O_3166,N_29887,N_28998);
nand UO_3167 (O_3167,N_29157,N_28806);
nor UO_3168 (O_3168,N_28837,N_28976);
xnor UO_3169 (O_3169,N_29192,N_29136);
nor UO_3170 (O_3170,N_29703,N_29470);
xnor UO_3171 (O_3171,N_29663,N_29608);
and UO_3172 (O_3172,N_29504,N_28912);
or UO_3173 (O_3173,N_28866,N_29378);
nand UO_3174 (O_3174,N_29997,N_29973);
and UO_3175 (O_3175,N_28877,N_28805);
xnor UO_3176 (O_3176,N_29056,N_29832);
and UO_3177 (O_3177,N_29693,N_29544);
nand UO_3178 (O_3178,N_29079,N_29282);
or UO_3179 (O_3179,N_29212,N_29444);
nand UO_3180 (O_3180,N_29049,N_29501);
and UO_3181 (O_3181,N_29686,N_29335);
nand UO_3182 (O_3182,N_29839,N_28840);
xnor UO_3183 (O_3183,N_29675,N_28958);
nand UO_3184 (O_3184,N_29267,N_29935);
xor UO_3185 (O_3185,N_29634,N_28857);
and UO_3186 (O_3186,N_29611,N_29484);
nor UO_3187 (O_3187,N_29391,N_29625);
and UO_3188 (O_3188,N_29819,N_29697);
xnor UO_3189 (O_3189,N_29884,N_28806);
and UO_3190 (O_3190,N_29497,N_29586);
xnor UO_3191 (O_3191,N_29018,N_29081);
nor UO_3192 (O_3192,N_29708,N_29919);
and UO_3193 (O_3193,N_29147,N_29636);
and UO_3194 (O_3194,N_29153,N_29580);
nand UO_3195 (O_3195,N_29690,N_28961);
and UO_3196 (O_3196,N_29819,N_29144);
nand UO_3197 (O_3197,N_28925,N_29984);
nand UO_3198 (O_3198,N_29491,N_29217);
xor UO_3199 (O_3199,N_29557,N_29956);
xnor UO_3200 (O_3200,N_29189,N_29905);
nand UO_3201 (O_3201,N_29110,N_29928);
nand UO_3202 (O_3202,N_28821,N_29981);
nor UO_3203 (O_3203,N_29064,N_29185);
nand UO_3204 (O_3204,N_29062,N_29588);
nor UO_3205 (O_3205,N_29357,N_29412);
and UO_3206 (O_3206,N_29100,N_29540);
nand UO_3207 (O_3207,N_29118,N_29166);
and UO_3208 (O_3208,N_29710,N_28915);
nand UO_3209 (O_3209,N_29633,N_29161);
and UO_3210 (O_3210,N_29189,N_29095);
and UO_3211 (O_3211,N_29297,N_29071);
xnor UO_3212 (O_3212,N_29790,N_28840);
nor UO_3213 (O_3213,N_28999,N_28849);
and UO_3214 (O_3214,N_29797,N_29422);
nand UO_3215 (O_3215,N_29939,N_29761);
nor UO_3216 (O_3216,N_29202,N_29686);
or UO_3217 (O_3217,N_29619,N_29701);
nand UO_3218 (O_3218,N_29917,N_29468);
xnor UO_3219 (O_3219,N_29605,N_29511);
xnor UO_3220 (O_3220,N_28911,N_29884);
and UO_3221 (O_3221,N_29094,N_29791);
nand UO_3222 (O_3222,N_29861,N_28982);
nand UO_3223 (O_3223,N_28977,N_29499);
nand UO_3224 (O_3224,N_29175,N_29004);
xnor UO_3225 (O_3225,N_29168,N_29738);
nand UO_3226 (O_3226,N_29654,N_29828);
or UO_3227 (O_3227,N_29758,N_29323);
xor UO_3228 (O_3228,N_29661,N_29007);
or UO_3229 (O_3229,N_28873,N_29786);
or UO_3230 (O_3230,N_29325,N_29920);
or UO_3231 (O_3231,N_29566,N_29028);
nand UO_3232 (O_3232,N_28900,N_28816);
xor UO_3233 (O_3233,N_29676,N_29107);
nand UO_3234 (O_3234,N_29328,N_29598);
nor UO_3235 (O_3235,N_29647,N_29599);
or UO_3236 (O_3236,N_29173,N_29473);
nand UO_3237 (O_3237,N_28989,N_28894);
nor UO_3238 (O_3238,N_29032,N_28958);
xnor UO_3239 (O_3239,N_29359,N_29598);
nor UO_3240 (O_3240,N_29711,N_29953);
and UO_3241 (O_3241,N_29603,N_28819);
nand UO_3242 (O_3242,N_29256,N_29897);
nand UO_3243 (O_3243,N_28980,N_29627);
nand UO_3244 (O_3244,N_29196,N_28919);
or UO_3245 (O_3245,N_29496,N_29374);
or UO_3246 (O_3246,N_29320,N_28829);
or UO_3247 (O_3247,N_28891,N_29482);
and UO_3248 (O_3248,N_29672,N_29075);
or UO_3249 (O_3249,N_29377,N_29320);
and UO_3250 (O_3250,N_29961,N_29898);
or UO_3251 (O_3251,N_29143,N_29326);
nor UO_3252 (O_3252,N_29969,N_29737);
nand UO_3253 (O_3253,N_29065,N_29920);
nor UO_3254 (O_3254,N_29046,N_29616);
or UO_3255 (O_3255,N_29566,N_28928);
and UO_3256 (O_3256,N_29919,N_29161);
and UO_3257 (O_3257,N_28810,N_29261);
nor UO_3258 (O_3258,N_29978,N_29429);
xor UO_3259 (O_3259,N_29302,N_28921);
and UO_3260 (O_3260,N_29748,N_29440);
or UO_3261 (O_3261,N_29178,N_28970);
and UO_3262 (O_3262,N_29640,N_29584);
nor UO_3263 (O_3263,N_29639,N_29659);
and UO_3264 (O_3264,N_29312,N_29920);
nor UO_3265 (O_3265,N_29724,N_29715);
nand UO_3266 (O_3266,N_29741,N_28868);
xnor UO_3267 (O_3267,N_29399,N_29884);
nand UO_3268 (O_3268,N_29440,N_29062);
xor UO_3269 (O_3269,N_28868,N_29325);
and UO_3270 (O_3270,N_29285,N_29756);
and UO_3271 (O_3271,N_29951,N_29194);
and UO_3272 (O_3272,N_29345,N_29936);
nand UO_3273 (O_3273,N_28926,N_28849);
or UO_3274 (O_3274,N_29338,N_29014);
nor UO_3275 (O_3275,N_29934,N_29944);
or UO_3276 (O_3276,N_29989,N_29862);
and UO_3277 (O_3277,N_29034,N_29874);
nor UO_3278 (O_3278,N_29211,N_29311);
or UO_3279 (O_3279,N_28947,N_29607);
xnor UO_3280 (O_3280,N_29401,N_28968);
xnor UO_3281 (O_3281,N_28869,N_28978);
nor UO_3282 (O_3282,N_29903,N_28950);
xnor UO_3283 (O_3283,N_29516,N_29607);
nand UO_3284 (O_3284,N_29714,N_29122);
nand UO_3285 (O_3285,N_29893,N_29702);
or UO_3286 (O_3286,N_29068,N_29746);
or UO_3287 (O_3287,N_29824,N_29114);
nor UO_3288 (O_3288,N_29013,N_29578);
xnor UO_3289 (O_3289,N_29595,N_29988);
or UO_3290 (O_3290,N_29357,N_29032);
or UO_3291 (O_3291,N_29379,N_29719);
or UO_3292 (O_3292,N_29791,N_28989);
and UO_3293 (O_3293,N_29108,N_28928);
xor UO_3294 (O_3294,N_29636,N_29597);
xor UO_3295 (O_3295,N_29656,N_29353);
or UO_3296 (O_3296,N_29786,N_29148);
nor UO_3297 (O_3297,N_29051,N_29083);
or UO_3298 (O_3298,N_29327,N_29273);
or UO_3299 (O_3299,N_28825,N_29167);
nor UO_3300 (O_3300,N_29761,N_29203);
nand UO_3301 (O_3301,N_29851,N_29581);
or UO_3302 (O_3302,N_29080,N_29180);
and UO_3303 (O_3303,N_29424,N_29136);
or UO_3304 (O_3304,N_29885,N_29766);
and UO_3305 (O_3305,N_28958,N_29589);
nor UO_3306 (O_3306,N_29367,N_29068);
or UO_3307 (O_3307,N_29298,N_29694);
nor UO_3308 (O_3308,N_29383,N_28853);
xnor UO_3309 (O_3309,N_29944,N_29229);
and UO_3310 (O_3310,N_29614,N_29949);
nor UO_3311 (O_3311,N_29972,N_29437);
or UO_3312 (O_3312,N_29106,N_29998);
and UO_3313 (O_3313,N_29276,N_29126);
and UO_3314 (O_3314,N_29507,N_29073);
nor UO_3315 (O_3315,N_29075,N_29845);
and UO_3316 (O_3316,N_28932,N_28971);
or UO_3317 (O_3317,N_29108,N_29418);
nand UO_3318 (O_3318,N_29963,N_29666);
or UO_3319 (O_3319,N_29585,N_29559);
nor UO_3320 (O_3320,N_28998,N_29056);
nand UO_3321 (O_3321,N_29766,N_29486);
or UO_3322 (O_3322,N_29867,N_29226);
or UO_3323 (O_3323,N_28885,N_29216);
and UO_3324 (O_3324,N_29123,N_29964);
nor UO_3325 (O_3325,N_29948,N_29359);
and UO_3326 (O_3326,N_29355,N_29516);
or UO_3327 (O_3327,N_29989,N_29088);
nand UO_3328 (O_3328,N_29367,N_29898);
nor UO_3329 (O_3329,N_29651,N_29927);
and UO_3330 (O_3330,N_29977,N_29493);
nand UO_3331 (O_3331,N_29877,N_28924);
nand UO_3332 (O_3332,N_29105,N_28945);
and UO_3333 (O_3333,N_29041,N_29468);
xor UO_3334 (O_3334,N_29812,N_29545);
or UO_3335 (O_3335,N_29913,N_29590);
nand UO_3336 (O_3336,N_29819,N_29591);
and UO_3337 (O_3337,N_29763,N_29411);
xor UO_3338 (O_3338,N_29341,N_29704);
nor UO_3339 (O_3339,N_29679,N_29831);
xnor UO_3340 (O_3340,N_29589,N_29822);
nor UO_3341 (O_3341,N_29244,N_29455);
and UO_3342 (O_3342,N_29790,N_29914);
nand UO_3343 (O_3343,N_29980,N_29477);
nor UO_3344 (O_3344,N_29747,N_29739);
xor UO_3345 (O_3345,N_28830,N_29573);
nand UO_3346 (O_3346,N_29914,N_29276);
nand UO_3347 (O_3347,N_28952,N_29307);
or UO_3348 (O_3348,N_28965,N_29744);
xnor UO_3349 (O_3349,N_28962,N_29941);
nand UO_3350 (O_3350,N_29349,N_29096);
and UO_3351 (O_3351,N_29547,N_29191);
or UO_3352 (O_3352,N_29213,N_29252);
nand UO_3353 (O_3353,N_29970,N_28888);
xnor UO_3354 (O_3354,N_29661,N_29473);
nand UO_3355 (O_3355,N_29777,N_29961);
xnor UO_3356 (O_3356,N_29629,N_29303);
and UO_3357 (O_3357,N_28922,N_29197);
nor UO_3358 (O_3358,N_29220,N_29119);
and UO_3359 (O_3359,N_28890,N_28865);
nand UO_3360 (O_3360,N_29454,N_29437);
nor UO_3361 (O_3361,N_29361,N_28823);
nand UO_3362 (O_3362,N_29592,N_29221);
xor UO_3363 (O_3363,N_29636,N_28808);
or UO_3364 (O_3364,N_29092,N_29976);
nand UO_3365 (O_3365,N_28803,N_29870);
and UO_3366 (O_3366,N_29776,N_29643);
nor UO_3367 (O_3367,N_29757,N_29602);
nand UO_3368 (O_3368,N_29229,N_29680);
nor UO_3369 (O_3369,N_29584,N_29680);
xor UO_3370 (O_3370,N_29322,N_29754);
or UO_3371 (O_3371,N_29308,N_29214);
nand UO_3372 (O_3372,N_28900,N_29665);
and UO_3373 (O_3373,N_28848,N_28829);
nand UO_3374 (O_3374,N_29543,N_29589);
xnor UO_3375 (O_3375,N_29951,N_28819);
or UO_3376 (O_3376,N_29597,N_29425);
and UO_3377 (O_3377,N_29189,N_29896);
nand UO_3378 (O_3378,N_28914,N_29458);
nand UO_3379 (O_3379,N_29306,N_29323);
or UO_3380 (O_3380,N_29815,N_29038);
nand UO_3381 (O_3381,N_29344,N_28981);
or UO_3382 (O_3382,N_29366,N_28829);
xor UO_3383 (O_3383,N_29647,N_28977);
nand UO_3384 (O_3384,N_29678,N_28899);
nand UO_3385 (O_3385,N_29515,N_29246);
xnor UO_3386 (O_3386,N_28830,N_28861);
or UO_3387 (O_3387,N_29530,N_29929);
xnor UO_3388 (O_3388,N_29083,N_28930);
or UO_3389 (O_3389,N_29769,N_29038);
or UO_3390 (O_3390,N_29559,N_29680);
nand UO_3391 (O_3391,N_29344,N_28885);
nor UO_3392 (O_3392,N_29844,N_29404);
xor UO_3393 (O_3393,N_29874,N_28807);
xor UO_3394 (O_3394,N_29382,N_29000);
and UO_3395 (O_3395,N_29165,N_29053);
nand UO_3396 (O_3396,N_29299,N_29266);
nor UO_3397 (O_3397,N_29099,N_29568);
xnor UO_3398 (O_3398,N_28965,N_29845);
xnor UO_3399 (O_3399,N_29477,N_29929);
and UO_3400 (O_3400,N_29175,N_29847);
nor UO_3401 (O_3401,N_28912,N_29211);
and UO_3402 (O_3402,N_28852,N_29499);
and UO_3403 (O_3403,N_29244,N_29334);
or UO_3404 (O_3404,N_29410,N_29266);
and UO_3405 (O_3405,N_29957,N_29241);
nand UO_3406 (O_3406,N_28968,N_29343);
xnor UO_3407 (O_3407,N_29349,N_29726);
nand UO_3408 (O_3408,N_29724,N_29049);
or UO_3409 (O_3409,N_29635,N_29149);
nand UO_3410 (O_3410,N_29316,N_29871);
or UO_3411 (O_3411,N_28952,N_28891);
nor UO_3412 (O_3412,N_29916,N_29118);
and UO_3413 (O_3413,N_28853,N_29874);
and UO_3414 (O_3414,N_29548,N_28994);
nor UO_3415 (O_3415,N_29469,N_29648);
and UO_3416 (O_3416,N_28903,N_29077);
and UO_3417 (O_3417,N_29356,N_29295);
nand UO_3418 (O_3418,N_29086,N_28851);
nand UO_3419 (O_3419,N_29329,N_29518);
nor UO_3420 (O_3420,N_29891,N_29279);
or UO_3421 (O_3421,N_29483,N_29121);
and UO_3422 (O_3422,N_29651,N_29083);
or UO_3423 (O_3423,N_29705,N_29532);
xor UO_3424 (O_3424,N_29271,N_29004);
or UO_3425 (O_3425,N_28916,N_29959);
nor UO_3426 (O_3426,N_29513,N_29192);
nor UO_3427 (O_3427,N_29198,N_29192);
xnor UO_3428 (O_3428,N_29781,N_29449);
and UO_3429 (O_3429,N_28881,N_29069);
nand UO_3430 (O_3430,N_29587,N_29399);
nand UO_3431 (O_3431,N_29964,N_29793);
or UO_3432 (O_3432,N_29878,N_28890);
nor UO_3433 (O_3433,N_29292,N_29084);
and UO_3434 (O_3434,N_29095,N_29741);
xor UO_3435 (O_3435,N_29570,N_29105);
or UO_3436 (O_3436,N_29608,N_29837);
xnor UO_3437 (O_3437,N_29771,N_28841);
and UO_3438 (O_3438,N_29144,N_28890);
nor UO_3439 (O_3439,N_29895,N_29632);
xor UO_3440 (O_3440,N_28860,N_29686);
xnor UO_3441 (O_3441,N_29782,N_29249);
nor UO_3442 (O_3442,N_29127,N_29166);
xor UO_3443 (O_3443,N_29182,N_28940);
and UO_3444 (O_3444,N_29409,N_29557);
or UO_3445 (O_3445,N_28902,N_29692);
nor UO_3446 (O_3446,N_29874,N_29614);
or UO_3447 (O_3447,N_28848,N_28813);
and UO_3448 (O_3448,N_29273,N_28953);
or UO_3449 (O_3449,N_29808,N_29629);
and UO_3450 (O_3450,N_29102,N_29612);
xnor UO_3451 (O_3451,N_29894,N_29891);
nand UO_3452 (O_3452,N_29469,N_29878);
and UO_3453 (O_3453,N_29027,N_29271);
and UO_3454 (O_3454,N_29400,N_29223);
and UO_3455 (O_3455,N_29483,N_29878);
or UO_3456 (O_3456,N_29923,N_29318);
xnor UO_3457 (O_3457,N_29648,N_29356);
and UO_3458 (O_3458,N_28846,N_29938);
nor UO_3459 (O_3459,N_28858,N_29990);
nand UO_3460 (O_3460,N_29373,N_29860);
or UO_3461 (O_3461,N_29765,N_29280);
and UO_3462 (O_3462,N_29306,N_29599);
and UO_3463 (O_3463,N_29003,N_29824);
and UO_3464 (O_3464,N_29081,N_28838);
nand UO_3465 (O_3465,N_29052,N_29992);
xor UO_3466 (O_3466,N_28885,N_29360);
and UO_3467 (O_3467,N_29683,N_29522);
nand UO_3468 (O_3468,N_28923,N_29122);
nand UO_3469 (O_3469,N_29908,N_29260);
nand UO_3470 (O_3470,N_29320,N_29729);
and UO_3471 (O_3471,N_29509,N_29700);
nand UO_3472 (O_3472,N_29433,N_29336);
and UO_3473 (O_3473,N_29452,N_29339);
nand UO_3474 (O_3474,N_28877,N_28990);
nand UO_3475 (O_3475,N_29849,N_29745);
nand UO_3476 (O_3476,N_28951,N_28969);
nand UO_3477 (O_3477,N_29837,N_29971);
nor UO_3478 (O_3478,N_29626,N_29270);
and UO_3479 (O_3479,N_29519,N_29054);
xnor UO_3480 (O_3480,N_29709,N_29461);
xnor UO_3481 (O_3481,N_28951,N_29953);
and UO_3482 (O_3482,N_28944,N_29721);
nand UO_3483 (O_3483,N_29461,N_29261);
xor UO_3484 (O_3484,N_29895,N_29097);
and UO_3485 (O_3485,N_29160,N_29385);
and UO_3486 (O_3486,N_28996,N_29564);
nand UO_3487 (O_3487,N_29351,N_29855);
nand UO_3488 (O_3488,N_29530,N_29199);
or UO_3489 (O_3489,N_29259,N_29248);
or UO_3490 (O_3490,N_29990,N_29583);
nor UO_3491 (O_3491,N_29676,N_29190);
xnor UO_3492 (O_3492,N_29958,N_29029);
and UO_3493 (O_3493,N_29565,N_29325);
nor UO_3494 (O_3494,N_29230,N_29301);
nor UO_3495 (O_3495,N_29058,N_28837);
and UO_3496 (O_3496,N_29994,N_29104);
and UO_3497 (O_3497,N_28968,N_29973);
nand UO_3498 (O_3498,N_29995,N_29808);
and UO_3499 (O_3499,N_29734,N_29165);
endmodule