module basic_750_5000_1000_10_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_422,In_240);
xnor U1 (N_1,In_248,In_291);
nor U2 (N_2,In_563,In_288);
nor U3 (N_3,In_207,In_138);
or U4 (N_4,In_366,In_329);
nand U5 (N_5,In_727,In_224);
xor U6 (N_6,In_13,In_551);
nand U7 (N_7,In_544,In_312);
or U8 (N_8,In_638,In_424);
xnor U9 (N_9,In_25,In_453);
nor U10 (N_10,In_584,In_686);
or U11 (N_11,In_94,In_506);
or U12 (N_12,In_680,In_528);
nand U13 (N_13,In_324,In_83);
and U14 (N_14,In_123,In_667);
and U15 (N_15,In_494,In_262);
or U16 (N_16,In_327,In_533);
xor U17 (N_17,In_599,In_606);
or U18 (N_18,In_491,In_33);
nand U19 (N_19,In_610,In_696);
and U20 (N_20,In_173,In_79);
and U21 (N_21,In_443,In_616);
or U22 (N_22,In_97,In_404);
nand U23 (N_23,In_10,In_647);
nor U24 (N_24,In_605,In_187);
nor U25 (N_25,In_710,In_12);
and U26 (N_26,In_54,In_80);
nand U27 (N_27,In_595,In_532);
or U28 (N_28,In_249,In_624);
xor U29 (N_29,In_182,In_596);
nor U30 (N_30,In_447,In_472);
and U31 (N_31,In_482,In_631);
and U32 (N_32,In_322,In_474);
nor U33 (N_33,In_66,In_525);
nand U34 (N_34,In_590,In_625);
nor U35 (N_35,In_190,In_558);
nor U36 (N_36,In_174,In_62);
and U37 (N_37,In_516,In_611);
or U38 (N_38,In_729,In_635);
or U39 (N_39,In_734,In_451);
and U40 (N_40,In_163,In_577);
nor U41 (N_41,In_305,In_358);
nor U42 (N_42,In_340,In_156);
or U43 (N_43,In_53,In_698);
and U44 (N_44,In_261,In_529);
xor U45 (N_45,In_736,In_59);
or U46 (N_46,In_157,In_670);
nand U47 (N_47,In_378,In_444);
nor U48 (N_48,In_657,In_553);
nand U49 (N_49,In_20,In_67);
nand U50 (N_50,In_633,In_639);
nand U51 (N_51,In_649,In_268);
nor U52 (N_52,In_275,In_737);
or U53 (N_53,In_153,In_205);
nor U54 (N_54,In_620,In_653);
nand U55 (N_55,In_543,In_379);
xor U56 (N_56,In_211,In_317);
and U57 (N_57,In_400,In_258);
nor U58 (N_58,In_73,In_549);
nor U59 (N_59,In_345,In_50);
and U60 (N_60,In_298,In_93);
and U61 (N_61,In_343,In_226);
nor U62 (N_62,In_726,In_521);
or U63 (N_63,In_125,In_467);
or U64 (N_64,In_61,In_743);
or U65 (N_65,In_339,In_454);
nand U66 (N_66,In_722,In_14);
and U67 (N_67,In_320,In_176);
or U68 (N_68,In_143,In_391);
nand U69 (N_69,In_254,In_131);
or U70 (N_70,In_270,In_133);
nor U71 (N_71,In_6,In_403);
and U72 (N_72,In_277,In_744);
and U73 (N_73,In_180,In_387);
or U74 (N_74,In_711,In_384);
and U75 (N_75,In_65,In_32);
nand U76 (N_76,In_231,In_389);
nand U77 (N_77,In_542,In_665);
nor U78 (N_78,In_699,In_161);
and U79 (N_79,In_376,In_216);
and U80 (N_80,In_614,In_212);
nand U81 (N_81,In_420,In_655);
nor U82 (N_82,In_461,In_352);
nor U83 (N_83,In_367,In_185);
nor U84 (N_84,In_284,In_301);
and U85 (N_85,In_475,In_69);
nor U86 (N_86,In_200,In_552);
or U87 (N_87,In_477,In_483);
nand U88 (N_88,In_431,In_527);
nand U89 (N_89,In_508,In_242);
nor U90 (N_90,In_449,In_4);
nor U91 (N_91,In_707,In_489);
or U92 (N_92,In_332,In_661);
or U93 (N_93,In_417,In_114);
or U94 (N_94,In_437,In_372);
and U95 (N_95,In_683,In_406);
nor U96 (N_96,In_524,In_319);
or U97 (N_97,In_42,In_738);
and U98 (N_98,In_117,In_58);
nor U99 (N_99,In_547,In_354);
nor U100 (N_100,In_396,In_380);
nand U101 (N_101,In_382,In_583);
or U102 (N_102,In_194,In_336);
nand U103 (N_103,In_351,In_746);
xnor U104 (N_104,In_139,In_46);
nand U105 (N_105,In_589,In_31);
and U106 (N_106,In_225,In_158);
and U107 (N_107,In_468,In_423);
xor U108 (N_108,In_90,In_159);
nand U109 (N_109,In_559,In_105);
nand U110 (N_110,In_456,In_450);
or U111 (N_111,In_501,In_421);
or U112 (N_112,In_749,In_689);
or U113 (N_113,In_490,In_648);
nor U114 (N_114,In_199,In_723);
or U115 (N_115,In_507,In_446);
nand U116 (N_116,In_168,In_692);
nand U117 (N_117,In_656,In_162);
and U118 (N_118,In_705,In_392);
and U119 (N_119,In_412,In_292);
nand U120 (N_120,In_365,In_650);
nand U121 (N_121,In_742,In_18);
nand U122 (N_122,In_196,In_505);
and U123 (N_123,In_92,In_191);
or U124 (N_124,In_178,In_210);
or U125 (N_125,In_666,In_95);
and U126 (N_126,In_104,In_630);
and U127 (N_127,In_538,In_626);
or U128 (N_128,In_228,In_748);
nor U129 (N_129,In_269,In_747);
nand U130 (N_130,In_129,In_247);
nor U131 (N_131,In_230,In_333);
or U132 (N_132,In_175,In_578);
nand U133 (N_133,In_740,In_674);
and U134 (N_134,In_397,In_217);
xnor U135 (N_135,In_530,In_119);
nor U136 (N_136,In_604,In_356);
nor U137 (N_137,In_613,In_480);
and U138 (N_138,In_309,In_34);
and U139 (N_139,In_88,In_19);
or U140 (N_140,In_346,In_2);
or U141 (N_141,In_243,In_484);
nand U142 (N_142,In_427,In_654);
or U143 (N_143,In_659,In_75);
nor U144 (N_144,In_503,In_548);
or U145 (N_145,In_463,In_714);
nand U146 (N_146,In_98,In_272);
nor U147 (N_147,In_492,In_441);
or U148 (N_148,In_334,In_203);
or U149 (N_149,In_615,In_362);
and U150 (N_150,In_68,In_435);
nor U151 (N_151,In_436,In_569);
or U152 (N_152,In_509,In_581);
and U153 (N_153,In_592,In_260);
nand U154 (N_154,In_706,In_681);
nor U155 (N_155,In_290,In_252);
or U156 (N_156,In_349,In_363);
and U157 (N_157,In_238,In_428);
nand U158 (N_158,In_166,In_409);
xnor U159 (N_159,In_110,In_308);
nand U160 (N_160,In_360,In_321);
or U161 (N_161,In_264,In_323);
and U162 (N_162,In_385,In_671);
nand U163 (N_163,In_486,In_281);
and U164 (N_164,In_24,In_582);
or U165 (N_165,In_197,In_518);
nand U166 (N_166,In_641,In_251);
and U167 (N_167,In_643,In_520);
nor U168 (N_168,In_383,In_371);
nor U169 (N_169,In_687,In_130);
and U170 (N_170,In_357,In_562);
or U171 (N_171,In_410,In_287);
nor U172 (N_172,In_49,In_218);
and U173 (N_173,In_515,In_720);
nand U174 (N_174,In_580,In_607);
and U175 (N_175,In_390,In_44);
nand U176 (N_176,In_497,In_536);
and U177 (N_177,In_675,In_229);
nor U178 (N_178,In_370,In_154);
xnor U179 (N_179,In_405,In_87);
and U180 (N_180,In_43,In_337);
or U181 (N_181,In_219,In_364);
xnor U182 (N_182,In_120,In_38);
nand U183 (N_183,In_236,In_204);
and U184 (N_184,In_283,In_72);
and U185 (N_185,In_697,In_568);
and U186 (N_186,In_602,In_579);
nand U187 (N_187,In_498,In_608);
or U188 (N_188,In_668,In_145);
nand U189 (N_189,In_132,In_438);
or U190 (N_190,In_227,In_469);
or U191 (N_191,In_289,In_513);
and U192 (N_192,In_165,In_241);
or U193 (N_193,In_122,In_682);
nor U194 (N_194,In_77,In_537);
nor U195 (N_195,In_214,In_716);
nor U196 (N_196,In_500,In_11);
or U197 (N_197,In_150,In_74);
and U198 (N_198,In_171,In_223);
or U199 (N_199,In_106,In_297);
nand U200 (N_200,In_40,In_695);
and U201 (N_201,In_464,In_233);
nor U202 (N_202,In_684,In_566);
nor U203 (N_203,In_193,In_556);
nor U204 (N_204,In_267,In_222);
or U205 (N_205,In_672,In_246);
nor U206 (N_206,In_81,In_597);
and U207 (N_207,In_172,In_419);
nand U208 (N_208,In_432,In_70);
and U209 (N_209,In_1,In_198);
and U210 (N_210,In_17,In_135);
nor U211 (N_211,In_510,In_496);
xnor U212 (N_212,In_457,In_189);
or U213 (N_213,In_48,In_545);
or U214 (N_214,In_448,In_5);
nand U215 (N_215,In_411,In_539);
nor U216 (N_216,In_26,In_265);
or U217 (N_217,In_213,In_601);
nand U218 (N_218,In_293,In_282);
nor U219 (N_219,In_201,In_316);
or U220 (N_220,In_663,In_462);
xor U221 (N_221,In_560,In_646);
and U222 (N_222,In_148,In_554);
and U223 (N_223,In_700,In_587);
nand U224 (N_224,In_21,In_315);
or U225 (N_225,In_208,In_679);
and U226 (N_226,In_658,In_619);
nand U227 (N_227,In_644,In_426);
nand U228 (N_228,In_78,In_652);
and U229 (N_229,In_144,In_452);
or U230 (N_230,In_146,In_3);
nand U231 (N_231,In_164,In_84);
nor U232 (N_232,In_286,In_263);
and U233 (N_233,In_445,In_221);
nand U234 (N_234,In_41,In_306);
and U235 (N_235,In_22,In_202);
nand U236 (N_236,In_295,In_407);
nand U237 (N_237,In_0,In_459);
nand U238 (N_238,In_487,In_576);
and U239 (N_239,In_408,In_713);
nand U240 (N_240,In_519,In_550);
xnor U241 (N_241,In_593,In_621);
nor U242 (N_242,In_101,In_85);
or U243 (N_243,In_473,In_531);
nor U244 (N_244,In_121,In_458);
nor U245 (N_245,In_673,In_733);
or U246 (N_246,In_341,In_141);
or U247 (N_247,In_76,In_571);
nand U248 (N_248,In_499,In_134);
nor U249 (N_249,In_512,In_393);
and U250 (N_250,In_708,In_102);
nand U251 (N_251,In_302,In_476);
and U252 (N_252,In_118,In_628);
and U253 (N_253,In_721,In_618);
and U254 (N_254,In_485,In_694);
or U255 (N_255,In_86,In_276);
and U256 (N_256,In_188,In_669);
and U257 (N_257,In_600,In_245);
nor U258 (N_258,In_99,In_523);
and U259 (N_259,In_401,In_561);
and U260 (N_260,In_7,In_574);
nor U261 (N_261,In_313,In_167);
xnor U262 (N_262,In_28,In_398);
or U263 (N_263,In_206,In_96);
nand U264 (N_264,In_89,In_731);
or U265 (N_265,In_702,In_640);
or U266 (N_266,In_634,In_56);
and U267 (N_267,In_712,In_399);
nor U268 (N_268,In_266,In_30);
nand U269 (N_269,In_374,In_186);
nor U270 (N_270,In_386,In_585);
and U271 (N_271,In_326,In_693);
and U272 (N_272,In_124,In_465);
and U273 (N_273,In_381,In_442);
and U274 (N_274,In_573,In_414);
nor U275 (N_275,In_416,In_466);
and U276 (N_276,In_555,In_183);
nand U277 (N_277,In_540,In_739);
and U278 (N_278,In_636,In_715);
nor U279 (N_279,In_402,In_181);
or U280 (N_280,In_377,In_103);
nand U281 (N_281,In_271,In_331);
or U282 (N_282,In_570,In_373);
nand U283 (N_283,In_353,In_741);
and U284 (N_284,In_9,In_239);
or U285 (N_285,In_495,In_57);
or U286 (N_286,In_594,In_128);
nand U287 (N_287,In_688,In_603);
nand U288 (N_288,In_23,In_151);
nor U289 (N_289,In_622,In_318);
and U290 (N_290,In_250,In_355);
and U291 (N_291,In_60,In_63);
and U292 (N_292,In_126,In_678);
or U293 (N_293,In_645,In_195);
nor U294 (N_294,In_45,In_425);
nor U295 (N_295,In_310,In_415);
nand U296 (N_296,In_113,In_745);
or U297 (N_297,In_328,In_15);
or U298 (N_298,In_517,In_273);
or U299 (N_299,In_107,In_296);
or U300 (N_300,In_184,In_127);
nor U301 (N_301,In_481,In_709);
nor U302 (N_302,In_147,In_136);
nor U303 (N_303,In_91,In_137);
nor U304 (N_304,In_192,In_256);
and U305 (N_305,In_274,In_534);
nor U306 (N_306,In_369,In_27);
or U307 (N_307,In_623,In_116);
nor U308 (N_308,In_418,In_591);
and U309 (N_309,In_278,In_701);
nor U310 (N_310,In_279,In_237);
nor U311 (N_311,In_330,In_347);
and U312 (N_312,In_478,In_108);
nor U313 (N_313,In_342,In_511);
nor U314 (N_314,In_677,In_735);
nor U315 (N_315,In_470,In_155);
and U316 (N_316,In_685,In_586);
nor U317 (N_317,In_440,In_348);
or U318 (N_318,In_504,In_725);
xor U319 (N_319,In_177,In_567);
nor U320 (N_320,In_152,In_338);
and U321 (N_321,In_64,In_314);
nor U322 (N_322,In_588,In_637);
nor U323 (N_323,In_368,In_35);
nor U324 (N_324,In_609,In_335);
or U325 (N_325,In_557,In_111);
nand U326 (N_326,In_471,In_455);
nand U327 (N_327,In_169,In_325);
or U328 (N_328,In_29,In_220);
and U329 (N_329,In_47,In_535);
and U330 (N_330,In_257,In_304);
nand U331 (N_331,In_732,In_541);
nand U332 (N_332,In_234,In_253);
nand U333 (N_333,In_575,In_52);
nand U334 (N_334,In_526,In_140);
or U335 (N_335,In_502,In_717);
xor U336 (N_336,In_71,In_170);
nor U337 (N_337,In_703,In_394);
nand U338 (N_338,In_307,In_690);
and U339 (N_339,In_664,In_259);
or U340 (N_340,In_395,In_215);
nand U341 (N_341,In_598,In_37);
and U342 (N_342,In_299,In_294);
nor U343 (N_343,In_311,In_55);
and U344 (N_344,In_51,In_522);
xor U345 (N_345,In_660,In_361);
nor U346 (N_346,In_546,In_429);
nor U347 (N_347,In_285,In_662);
or U348 (N_348,In_642,In_719);
or U349 (N_349,In_244,In_375);
nor U350 (N_350,In_434,In_730);
or U351 (N_351,In_39,In_8);
and U352 (N_352,In_350,In_632);
nor U353 (N_353,In_344,In_439);
nor U354 (N_354,In_565,In_514);
nor U355 (N_355,In_115,In_255);
or U356 (N_356,In_160,In_413);
and U357 (N_357,In_430,In_617);
or U358 (N_358,In_235,In_300);
and U359 (N_359,In_479,In_232);
nand U360 (N_360,In_149,In_728);
nand U361 (N_361,In_718,In_36);
or U362 (N_362,In_100,In_493);
or U363 (N_363,In_691,In_142);
and U364 (N_364,In_627,In_651);
and U365 (N_365,In_572,In_612);
nand U366 (N_366,In_303,In_280);
nand U367 (N_367,In_359,In_388);
nor U368 (N_368,In_629,In_16);
nand U369 (N_369,In_179,In_488);
and U370 (N_370,In_676,In_724);
or U371 (N_371,In_112,In_82);
and U372 (N_372,In_433,In_704);
nor U373 (N_373,In_209,In_564);
and U374 (N_374,In_109,In_460);
nor U375 (N_375,In_263,In_498);
nor U376 (N_376,In_188,In_545);
or U377 (N_377,In_201,In_363);
nand U378 (N_378,In_63,In_424);
or U379 (N_379,In_500,In_397);
nand U380 (N_380,In_88,In_460);
and U381 (N_381,In_166,In_353);
nand U382 (N_382,In_353,In_403);
nand U383 (N_383,In_668,In_200);
or U384 (N_384,In_309,In_628);
nor U385 (N_385,In_561,In_45);
and U386 (N_386,In_614,In_724);
nand U387 (N_387,In_176,In_274);
or U388 (N_388,In_594,In_633);
nand U389 (N_389,In_68,In_122);
and U390 (N_390,In_480,In_383);
nand U391 (N_391,In_52,In_113);
or U392 (N_392,In_15,In_390);
or U393 (N_393,In_548,In_464);
and U394 (N_394,In_93,In_337);
and U395 (N_395,In_354,In_190);
nor U396 (N_396,In_297,In_435);
nand U397 (N_397,In_714,In_536);
and U398 (N_398,In_24,In_704);
xnor U399 (N_399,In_442,In_573);
nand U400 (N_400,In_167,In_170);
or U401 (N_401,In_300,In_24);
nor U402 (N_402,In_288,In_177);
or U403 (N_403,In_271,In_438);
or U404 (N_404,In_355,In_331);
nand U405 (N_405,In_620,In_147);
nand U406 (N_406,In_57,In_643);
and U407 (N_407,In_123,In_124);
and U408 (N_408,In_517,In_698);
and U409 (N_409,In_220,In_168);
or U410 (N_410,In_104,In_528);
or U411 (N_411,In_680,In_748);
nand U412 (N_412,In_638,In_162);
nor U413 (N_413,In_249,In_389);
or U414 (N_414,In_399,In_422);
nor U415 (N_415,In_99,In_141);
or U416 (N_416,In_200,In_563);
or U417 (N_417,In_98,In_58);
or U418 (N_418,In_415,In_302);
or U419 (N_419,In_110,In_652);
or U420 (N_420,In_498,In_117);
or U421 (N_421,In_184,In_393);
nand U422 (N_422,In_299,In_406);
nand U423 (N_423,In_465,In_277);
nand U424 (N_424,In_91,In_34);
or U425 (N_425,In_478,In_306);
nor U426 (N_426,In_620,In_290);
nand U427 (N_427,In_483,In_14);
nand U428 (N_428,In_109,In_544);
nand U429 (N_429,In_195,In_320);
and U430 (N_430,In_246,In_383);
or U431 (N_431,In_68,In_742);
and U432 (N_432,In_512,In_546);
nor U433 (N_433,In_510,In_605);
nand U434 (N_434,In_670,In_181);
or U435 (N_435,In_500,In_275);
and U436 (N_436,In_21,In_511);
or U437 (N_437,In_35,In_47);
nor U438 (N_438,In_199,In_467);
nand U439 (N_439,In_492,In_338);
nand U440 (N_440,In_224,In_108);
and U441 (N_441,In_294,In_246);
nor U442 (N_442,In_582,In_694);
nor U443 (N_443,In_155,In_601);
and U444 (N_444,In_591,In_708);
nand U445 (N_445,In_722,In_604);
nand U446 (N_446,In_614,In_482);
xor U447 (N_447,In_362,In_322);
xor U448 (N_448,In_463,In_391);
nand U449 (N_449,In_278,In_466);
nand U450 (N_450,In_597,In_117);
nand U451 (N_451,In_250,In_104);
or U452 (N_452,In_274,In_743);
and U453 (N_453,In_576,In_171);
and U454 (N_454,In_102,In_504);
xor U455 (N_455,In_331,In_127);
and U456 (N_456,In_295,In_79);
and U457 (N_457,In_691,In_463);
nand U458 (N_458,In_361,In_264);
and U459 (N_459,In_153,In_648);
nand U460 (N_460,In_569,In_421);
and U461 (N_461,In_568,In_514);
or U462 (N_462,In_316,In_100);
or U463 (N_463,In_746,In_113);
and U464 (N_464,In_184,In_724);
or U465 (N_465,In_514,In_431);
nand U466 (N_466,In_743,In_262);
and U467 (N_467,In_372,In_92);
and U468 (N_468,In_154,In_503);
or U469 (N_469,In_626,In_71);
and U470 (N_470,In_510,In_222);
nor U471 (N_471,In_347,In_309);
nor U472 (N_472,In_266,In_136);
and U473 (N_473,In_284,In_677);
nor U474 (N_474,In_425,In_181);
nor U475 (N_475,In_468,In_149);
and U476 (N_476,In_161,In_397);
or U477 (N_477,In_179,In_537);
or U478 (N_478,In_64,In_227);
or U479 (N_479,In_473,In_657);
and U480 (N_480,In_65,In_724);
nand U481 (N_481,In_427,In_264);
xor U482 (N_482,In_698,In_98);
nand U483 (N_483,In_698,In_48);
nor U484 (N_484,In_233,In_484);
nor U485 (N_485,In_741,In_266);
and U486 (N_486,In_44,In_145);
or U487 (N_487,In_644,In_32);
nand U488 (N_488,In_562,In_748);
nand U489 (N_489,In_642,In_339);
nor U490 (N_490,In_329,In_520);
or U491 (N_491,In_105,In_313);
nor U492 (N_492,In_23,In_101);
or U493 (N_493,In_378,In_566);
or U494 (N_494,In_509,In_336);
nand U495 (N_495,In_160,In_209);
or U496 (N_496,In_426,In_160);
or U497 (N_497,In_58,In_663);
and U498 (N_498,In_137,In_619);
and U499 (N_499,In_196,In_565);
and U500 (N_500,N_348,N_105);
or U501 (N_501,N_32,N_294);
nand U502 (N_502,N_435,N_109);
and U503 (N_503,N_383,N_25);
nor U504 (N_504,N_399,N_47);
nor U505 (N_505,N_329,N_289);
xor U506 (N_506,N_246,N_271);
or U507 (N_507,N_416,N_213);
nor U508 (N_508,N_48,N_287);
nand U509 (N_509,N_41,N_485);
nand U510 (N_510,N_172,N_312);
or U511 (N_511,N_317,N_366);
nor U512 (N_512,N_180,N_187);
nor U513 (N_513,N_355,N_147);
nand U514 (N_514,N_198,N_107);
or U515 (N_515,N_33,N_17);
nand U516 (N_516,N_481,N_438);
xnor U517 (N_517,N_133,N_402);
and U518 (N_518,N_376,N_184);
and U519 (N_519,N_459,N_77);
or U520 (N_520,N_212,N_309);
nor U521 (N_521,N_468,N_127);
and U522 (N_522,N_258,N_16);
nand U523 (N_523,N_363,N_283);
nor U524 (N_524,N_306,N_232);
nor U525 (N_525,N_297,N_342);
nor U526 (N_526,N_448,N_320);
nor U527 (N_527,N_465,N_131);
nor U528 (N_528,N_268,N_168);
nor U529 (N_529,N_205,N_266);
nand U530 (N_530,N_279,N_391);
nand U531 (N_531,N_66,N_207);
and U532 (N_532,N_265,N_301);
nor U533 (N_533,N_296,N_97);
and U534 (N_534,N_136,N_139);
nor U535 (N_535,N_362,N_423);
and U536 (N_536,N_252,N_71);
nor U537 (N_537,N_2,N_42);
nor U538 (N_538,N_194,N_494);
or U539 (N_539,N_454,N_189);
xor U540 (N_540,N_85,N_470);
or U541 (N_541,N_19,N_20);
nand U542 (N_542,N_324,N_98);
nand U543 (N_543,N_11,N_247);
and U544 (N_544,N_352,N_110);
and U545 (N_545,N_386,N_316);
and U546 (N_546,N_488,N_335);
nand U547 (N_547,N_349,N_123);
and U548 (N_548,N_118,N_344);
nor U549 (N_549,N_122,N_436);
nand U550 (N_550,N_197,N_364);
or U551 (N_551,N_144,N_460);
and U552 (N_552,N_290,N_298);
nand U553 (N_553,N_55,N_395);
or U554 (N_554,N_236,N_166);
nand U555 (N_555,N_149,N_281);
nand U556 (N_556,N_219,N_155);
or U557 (N_557,N_200,N_156);
nor U558 (N_558,N_379,N_418);
nor U559 (N_559,N_36,N_134);
nand U560 (N_560,N_313,N_472);
nand U561 (N_561,N_221,N_196);
or U562 (N_562,N_430,N_69);
nor U563 (N_563,N_241,N_95);
nand U564 (N_564,N_492,N_469);
and U565 (N_565,N_433,N_409);
nor U566 (N_566,N_330,N_201);
or U567 (N_567,N_463,N_115);
nand U568 (N_568,N_372,N_257);
nand U569 (N_569,N_327,N_457);
or U570 (N_570,N_169,N_401);
or U571 (N_571,N_173,N_35);
or U572 (N_572,N_151,N_114);
or U573 (N_573,N_199,N_275);
or U574 (N_574,N_230,N_239);
and U575 (N_575,N_319,N_22);
or U576 (N_576,N_286,N_461);
or U577 (N_577,N_14,N_458);
and U578 (N_578,N_140,N_410);
nand U579 (N_579,N_272,N_228);
nand U580 (N_580,N_373,N_256);
or U581 (N_581,N_34,N_152);
nand U582 (N_582,N_204,N_338);
or U583 (N_583,N_181,N_83);
and U584 (N_584,N_174,N_243);
nand U585 (N_585,N_428,N_489);
nor U586 (N_586,N_210,N_393);
xor U587 (N_587,N_394,N_190);
or U588 (N_588,N_245,N_453);
nand U589 (N_589,N_466,N_478);
or U590 (N_590,N_214,N_18);
and U591 (N_591,N_30,N_64);
nand U592 (N_592,N_462,N_80);
or U593 (N_593,N_273,N_274);
and U594 (N_594,N_99,N_79);
and U595 (N_595,N_100,N_81);
nand U596 (N_596,N_90,N_185);
and U597 (N_597,N_182,N_321);
nor U598 (N_598,N_371,N_455);
or U599 (N_599,N_129,N_427);
nand U600 (N_600,N_499,N_112);
or U601 (N_601,N_400,N_343);
or U602 (N_602,N_424,N_405);
nand U603 (N_603,N_103,N_354);
nand U604 (N_604,N_227,N_217);
and U605 (N_605,N_65,N_331);
nor U606 (N_606,N_135,N_153);
or U607 (N_607,N_218,N_484);
and U608 (N_608,N_482,N_381);
nor U609 (N_609,N_419,N_254);
and U610 (N_610,N_425,N_295);
or U611 (N_611,N_164,N_8);
and U612 (N_612,N_456,N_78);
or U613 (N_613,N_493,N_440);
nand U614 (N_614,N_452,N_387);
or U615 (N_615,N_367,N_292);
and U616 (N_616,N_62,N_323);
and U617 (N_617,N_191,N_59);
nor U618 (N_618,N_377,N_75);
and U619 (N_619,N_480,N_27);
or U620 (N_620,N_390,N_206);
and U621 (N_621,N_276,N_72);
nor U622 (N_622,N_229,N_420);
or U623 (N_623,N_175,N_439);
or U624 (N_624,N_491,N_111);
nand U625 (N_625,N_162,N_495);
nand U626 (N_626,N_163,N_238);
nor U627 (N_627,N_128,N_61);
and U628 (N_628,N_192,N_6);
or U629 (N_629,N_94,N_57);
and U630 (N_630,N_269,N_497);
or U631 (N_631,N_260,N_421);
or U632 (N_632,N_345,N_249);
nor U633 (N_633,N_93,N_177);
nand U634 (N_634,N_250,N_89);
nand U635 (N_635,N_186,N_96);
nand U636 (N_636,N_141,N_270);
nor U637 (N_637,N_308,N_356);
or U638 (N_638,N_259,N_261);
or U639 (N_639,N_403,N_53);
and U640 (N_640,N_76,N_336);
or U641 (N_641,N_159,N_483);
and U642 (N_642,N_347,N_178);
nand U643 (N_643,N_225,N_242);
or U644 (N_644,N_293,N_496);
or U645 (N_645,N_479,N_5);
nand U646 (N_646,N_86,N_248);
nand U647 (N_647,N_255,N_434);
and U648 (N_648,N_444,N_56);
and U649 (N_649,N_464,N_498);
or U650 (N_650,N_26,N_233);
and U651 (N_651,N_380,N_411);
and U652 (N_652,N_358,N_124);
and U653 (N_653,N_116,N_29);
and U654 (N_654,N_475,N_0);
and U655 (N_655,N_88,N_44);
nor U656 (N_656,N_339,N_130);
nand U657 (N_657,N_368,N_346);
or U658 (N_658,N_9,N_304);
and U659 (N_659,N_326,N_220);
nand U660 (N_660,N_31,N_52);
and U661 (N_661,N_333,N_132);
nand U662 (N_662,N_285,N_431);
nor U663 (N_663,N_137,N_150);
nor U664 (N_664,N_193,N_441);
and U665 (N_665,N_40,N_325);
or U666 (N_666,N_106,N_63);
or U667 (N_667,N_442,N_280);
nand U668 (N_668,N_121,N_361);
or U669 (N_669,N_4,N_91);
nand U670 (N_670,N_102,N_369);
or U671 (N_671,N_167,N_334);
xnor U672 (N_672,N_240,N_449);
and U673 (N_673,N_303,N_226);
and U674 (N_674,N_417,N_45);
nand U675 (N_675,N_117,N_211);
and U676 (N_676,N_3,N_486);
nor U677 (N_677,N_278,N_23);
nand U678 (N_678,N_7,N_51);
nor U679 (N_679,N_341,N_21);
and U680 (N_680,N_68,N_474);
and U681 (N_681,N_397,N_158);
or U682 (N_682,N_378,N_74);
xnor U683 (N_683,N_1,N_203);
and U684 (N_684,N_209,N_222);
nor U685 (N_685,N_38,N_165);
nor U686 (N_686,N_148,N_92);
nor U687 (N_687,N_54,N_385);
or U688 (N_688,N_412,N_125);
and U689 (N_689,N_476,N_328);
nand U690 (N_690,N_215,N_406);
nand U691 (N_691,N_350,N_473);
and U692 (N_692,N_277,N_82);
nor U693 (N_693,N_73,N_50);
xnor U694 (N_694,N_311,N_113);
or U695 (N_695,N_15,N_157);
nand U696 (N_696,N_108,N_101);
nand U697 (N_697,N_37,N_202);
or U698 (N_698,N_288,N_145);
nand U699 (N_699,N_398,N_87);
xnor U700 (N_700,N_307,N_471);
and U701 (N_701,N_332,N_337);
nand U702 (N_702,N_414,N_39);
or U703 (N_703,N_104,N_451);
nor U704 (N_704,N_300,N_357);
and U705 (N_705,N_404,N_67);
and U706 (N_706,N_291,N_119);
nand U707 (N_707,N_208,N_176);
nand U708 (N_708,N_370,N_360);
xor U709 (N_709,N_353,N_388);
nand U710 (N_710,N_138,N_359);
nand U711 (N_711,N_384,N_12);
and U712 (N_712,N_422,N_263);
nor U713 (N_713,N_264,N_322);
or U714 (N_714,N_450,N_195);
nor U715 (N_715,N_413,N_446);
or U716 (N_716,N_84,N_443);
nand U717 (N_717,N_244,N_60);
nor U718 (N_718,N_447,N_10);
nand U719 (N_719,N_188,N_235);
or U720 (N_720,N_445,N_154);
nor U721 (N_721,N_267,N_415);
nor U722 (N_722,N_432,N_43);
and U723 (N_723,N_224,N_171);
and U724 (N_724,N_143,N_142);
or U725 (N_725,N_310,N_467);
and U726 (N_726,N_314,N_179);
and U727 (N_727,N_216,N_223);
and U728 (N_728,N_389,N_396);
or U729 (N_729,N_253,N_13);
or U730 (N_730,N_351,N_284);
nor U731 (N_731,N_46,N_262);
nand U732 (N_732,N_299,N_477);
nor U733 (N_733,N_365,N_183);
nand U734 (N_734,N_170,N_231);
and U735 (N_735,N_407,N_318);
or U736 (N_736,N_487,N_408);
nand U737 (N_737,N_490,N_49);
nand U738 (N_738,N_234,N_120);
and U739 (N_739,N_437,N_161);
nor U740 (N_740,N_146,N_426);
nand U741 (N_741,N_237,N_374);
nor U742 (N_742,N_382,N_126);
nand U743 (N_743,N_340,N_251);
or U744 (N_744,N_70,N_282);
and U745 (N_745,N_392,N_315);
and U746 (N_746,N_302,N_429);
nand U747 (N_747,N_160,N_305);
nand U748 (N_748,N_375,N_58);
or U749 (N_749,N_24,N_28);
xor U750 (N_750,N_229,N_444);
or U751 (N_751,N_489,N_280);
nor U752 (N_752,N_8,N_250);
or U753 (N_753,N_439,N_275);
nand U754 (N_754,N_154,N_489);
and U755 (N_755,N_382,N_16);
nor U756 (N_756,N_351,N_290);
nor U757 (N_757,N_391,N_459);
nand U758 (N_758,N_181,N_199);
and U759 (N_759,N_104,N_454);
nand U760 (N_760,N_190,N_312);
xnor U761 (N_761,N_150,N_262);
or U762 (N_762,N_314,N_24);
or U763 (N_763,N_22,N_435);
and U764 (N_764,N_88,N_323);
or U765 (N_765,N_432,N_296);
and U766 (N_766,N_136,N_130);
and U767 (N_767,N_269,N_50);
or U768 (N_768,N_238,N_198);
nor U769 (N_769,N_158,N_460);
nand U770 (N_770,N_266,N_281);
or U771 (N_771,N_303,N_229);
and U772 (N_772,N_249,N_225);
or U773 (N_773,N_305,N_331);
or U774 (N_774,N_231,N_405);
and U775 (N_775,N_97,N_227);
and U776 (N_776,N_382,N_181);
and U777 (N_777,N_394,N_222);
and U778 (N_778,N_109,N_295);
or U779 (N_779,N_182,N_346);
nand U780 (N_780,N_52,N_234);
or U781 (N_781,N_403,N_314);
and U782 (N_782,N_341,N_356);
nor U783 (N_783,N_184,N_484);
and U784 (N_784,N_492,N_465);
nand U785 (N_785,N_132,N_263);
and U786 (N_786,N_43,N_7);
nand U787 (N_787,N_365,N_209);
nand U788 (N_788,N_274,N_224);
or U789 (N_789,N_344,N_71);
and U790 (N_790,N_60,N_368);
and U791 (N_791,N_0,N_334);
nand U792 (N_792,N_279,N_227);
and U793 (N_793,N_318,N_8);
and U794 (N_794,N_277,N_4);
or U795 (N_795,N_354,N_199);
nor U796 (N_796,N_290,N_244);
and U797 (N_797,N_279,N_78);
nand U798 (N_798,N_456,N_28);
and U799 (N_799,N_114,N_275);
nand U800 (N_800,N_122,N_247);
and U801 (N_801,N_115,N_310);
nor U802 (N_802,N_447,N_208);
nor U803 (N_803,N_389,N_345);
nand U804 (N_804,N_473,N_41);
or U805 (N_805,N_376,N_38);
or U806 (N_806,N_150,N_281);
nor U807 (N_807,N_347,N_325);
nand U808 (N_808,N_441,N_283);
and U809 (N_809,N_349,N_231);
nor U810 (N_810,N_82,N_149);
and U811 (N_811,N_267,N_307);
nand U812 (N_812,N_356,N_214);
nand U813 (N_813,N_33,N_310);
and U814 (N_814,N_465,N_295);
nor U815 (N_815,N_433,N_230);
and U816 (N_816,N_60,N_258);
nand U817 (N_817,N_34,N_325);
or U818 (N_818,N_148,N_244);
nand U819 (N_819,N_1,N_194);
and U820 (N_820,N_365,N_212);
nand U821 (N_821,N_480,N_271);
nor U822 (N_822,N_196,N_227);
nand U823 (N_823,N_104,N_457);
xnor U824 (N_824,N_361,N_228);
nand U825 (N_825,N_70,N_297);
and U826 (N_826,N_188,N_431);
or U827 (N_827,N_309,N_196);
nand U828 (N_828,N_309,N_380);
or U829 (N_829,N_195,N_53);
nor U830 (N_830,N_486,N_489);
nand U831 (N_831,N_295,N_73);
nor U832 (N_832,N_169,N_499);
or U833 (N_833,N_175,N_342);
or U834 (N_834,N_288,N_377);
nor U835 (N_835,N_406,N_325);
nand U836 (N_836,N_184,N_82);
or U837 (N_837,N_167,N_394);
or U838 (N_838,N_227,N_226);
nand U839 (N_839,N_204,N_446);
xnor U840 (N_840,N_335,N_412);
nand U841 (N_841,N_167,N_254);
nor U842 (N_842,N_355,N_344);
and U843 (N_843,N_194,N_8);
nor U844 (N_844,N_214,N_312);
and U845 (N_845,N_398,N_149);
nor U846 (N_846,N_223,N_240);
nor U847 (N_847,N_210,N_243);
nor U848 (N_848,N_104,N_172);
nand U849 (N_849,N_57,N_242);
and U850 (N_850,N_370,N_257);
nand U851 (N_851,N_440,N_437);
or U852 (N_852,N_54,N_473);
nor U853 (N_853,N_444,N_366);
or U854 (N_854,N_132,N_393);
and U855 (N_855,N_181,N_247);
nand U856 (N_856,N_366,N_2);
or U857 (N_857,N_397,N_283);
and U858 (N_858,N_5,N_311);
nand U859 (N_859,N_221,N_179);
nor U860 (N_860,N_155,N_73);
and U861 (N_861,N_244,N_266);
xor U862 (N_862,N_111,N_6);
or U863 (N_863,N_487,N_315);
nand U864 (N_864,N_30,N_140);
nor U865 (N_865,N_0,N_65);
and U866 (N_866,N_111,N_179);
or U867 (N_867,N_236,N_436);
nand U868 (N_868,N_127,N_382);
or U869 (N_869,N_119,N_45);
and U870 (N_870,N_0,N_171);
nor U871 (N_871,N_125,N_270);
nor U872 (N_872,N_26,N_232);
and U873 (N_873,N_272,N_159);
nor U874 (N_874,N_248,N_288);
nor U875 (N_875,N_340,N_217);
and U876 (N_876,N_184,N_398);
and U877 (N_877,N_389,N_216);
nand U878 (N_878,N_214,N_421);
xnor U879 (N_879,N_65,N_127);
or U880 (N_880,N_47,N_367);
and U881 (N_881,N_354,N_389);
nand U882 (N_882,N_244,N_165);
and U883 (N_883,N_45,N_418);
and U884 (N_884,N_480,N_454);
and U885 (N_885,N_121,N_78);
or U886 (N_886,N_368,N_2);
and U887 (N_887,N_20,N_415);
nor U888 (N_888,N_170,N_432);
and U889 (N_889,N_266,N_232);
or U890 (N_890,N_386,N_146);
or U891 (N_891,N_76,N_340);
nand U892 (N_892,N_496,N_137);
or U893 (N_893,N_79,N_340);
nand U894 (N_894,N_204,N_263);
or U895 (N_895,N_55,N_327);
nor U896 (N_896,N_246,N_230);
or U897 (N_897,N_141,N_22);
nor U898 (N_898,N_17,N_344);
nor U899 (N_899,N_255,N_61);
nor U900 (N_900,N_470,N_120);
nor U901 (N_901,N_290,N_131);
nand U902 (N_902,N_98,N_424);
nand U903 (N_903,N_70,N_380);
nand U904 (N_904,N_54,N_311);
or U905 (N_905,N_380,N_440);
nor U906 (N_906,N_36,N_252);
and U907 (N_907,N_399,N_132);
nand U908 (N_908,N_478,N_69);
xnor U909 (N_909,N_198,N_422);
xor U910 (N_910,N_233,N_423);
and U911 (N_911,N_107,N_238);
nand U912 (N_912,N_381,N_494);
or U913 (N_913,N_402,N_427);
or U914 (N_914,N_392,N_58);
nand U915 (N_915,N_249,N_381);
nand U916 (N_916,N_276,N_82);
nor U917 (N_917,N_403,N_163);
nand U918 (N_918,N_461,N_267);
nand U919 (N_919,N_146,N_365);
nand U920 (N_920,N_63,N_233);
nor U921 (N_921,N_58,N_216);
nor U922 (N_922,N_61,N_270);
and U923 (N_923,N_225,N_287);
and U924 (N_924,N_237,N_132);
xnor U925 (N_925,N_101,N_379);
nand U926 (N_926,N_495,N_94);
nor U927 (N_927,N_201,N_109);
nand U928 (N_928,N_242,N_161);
or U929 (N_929,N_488,N_426);
or U930 (N_930,N_457,N_160);
or U931 (N_931,N_389,N_1);
nand U932 (N_932,N_352,N_305);
nor U933 (N_933,N_273,N_350);
or U934 (N_934,N_153,N_487);
and U935 (N_935,N_21,N_193);
nor U936 (N_936,N_154,N_14);
nand U937 (N_937,N_294,N_124);
and U938 (N_938,N_286,N_231);
or U939 (N_939,N_387,N_257);
and U940 (N_940,N_264,N_387);
nand U941 (N_941,N_138,N_242);
xor U942 (N_942,N_303,N_25);
and U943 (N_943,N_447,N_18);
and U944 (N_944,N_473,N_104);
or U945 (N_945,N_44,N_63);
nand U946 (N_946,N_409,N_194);
and U947 (N_947,N_286,N_137);
or U948 (N_948,N_125,N_252);
nand U949 (N_949,N_213,N_349);
nor U950 (N_950,N_405,N_212);
or U951 (N_951,N_18,N_225);
or U952 (N_952,N_332,N_303);
or U953 (N_953,N_134,N_414);
and U954 (N_954,N_394,N_265);
nand U955 (N_955,N_467,N_221);
nor U956 (N_956,N_166,N_291);
nor U957 (N_957,N_320,N_41);
nand U958 (N_958,N_194,N_58);
nand U959 (N_959,N_127,N_450);
nor U960 (N_960,N_420,N_379);
and U961 (N_961,N_283,N_117);
nor U962 (N_962,N_11,N_189);
and U963 (N_963,N_98,N_100);
or U964 (N_964,N_0,N_392);
or U965 (N_965,N_41,N_215);
nand U966 (N_966,N_174,N_178);
nand U967 (N_967,N_21,N_126);
and U968 (N_968,N_339,N_399);
and U969 (N_969,N_93,N_489);
or U970 (N_970,N_45,N_29);
and U971 (N_971,N_244,N_393);
nor U972 (N_972,N_466,N_157);
nor U973 (N_973,N_34,N_48);
xor U974 (N_974,N_170,N_499);
nor U975 (N_975,N_52,N_163);
or U976 (N_976,N_128,N_109);
nor U977 (N_977,N_122,N_139);
nor U978 (N_978,N_143,N_316);
nor U979 (N_979,N_398,N_400);
nor U980 (N_980,N_463,N_379);
nand U981 (N_981,N_361,N_392);
nand U982 (N_982,N_118,N_206);
or U983 (N_983,N_334,N_393);
or U984 (N_984,N_390,N_170);
or U985 (N_985,N_98,N_9);
nor U986 (N_986,N_343,N_316);
nor U987 (N_987,N_424,N_441);
nand U988 (N_988,N_27,N_17);
nor U989 (N_989,N_176,N_294);
nand U990 (N_990,N_50,N_382);
nand U991 (N_991,N_101,N_401);
nor U992 (N_992,N_279,N_270);
xnor U993 (N_993,N_337,N_426);
and U994 (N_994,N_296,N_40);
or U995 (N_995,N_93,N_122);
nor U996 (N_996,N_234,N_394);
and U997 (N_997,N_142,N_155);
nand U998 (N_998,N_464,N_49);
or U999 (N_999,N_113,N_225);
nand U1000 (N_1000,N_625,N_581);
nand U1001 (N_1001,N_689,N_601);
nand U1002 (N_1002,N_740,N_569);
or U1003 (N_1003,N_656,N_950);
nand U1004 (N_1004,N_989,N_574);
nor U1005 (N_1005,N_712,N_788);
and U1006 (N_1006,N_960,N_813);
nand U1007 (N_1007,N_739,N_845);
and U1008 (N_1008,N_795,N_903);
and U1009 (N_1009,N_636,N_759);
or U1010 (N_1010,N_791,N_974);
nand U1011 (N_1011,N_825,N_541);
nor U1012 (N_1012,N_592,N_990);
nand U1013 (N_1013,N_724,N_725);
or U1014 (N_1014,N_688,N_786);
nor U1015 (N_1015,N_797,N_615);
nand U1016 (N_1016,N_567,N_627);
xor U1017 (N_1017,N_503,N_628);
or U1018 (N_1018,N_604,N_719);
xor U1019 (N_1019,N_629,N_777);
nand U1020 (N_1020,N_707,N_940);
nand U1021 (N_1021,N_622,N_742);
or U1022 (N_1022,N_736,N_545);
nor U1023 (N_1023,N_593,N_681);
nor U1024 (N_1024,N_561,N_898);
and U1025 (N_1025,N_958,N_512);
or U1026 (N_1026,N_506,N_927);
and U1027 (N_1027,N_917,N_954);
or U1028 (N_1028,N_649,N_873);
xor U1029 (N_1029,N_714,N_527);
or U1030 (N_1030,N_860,N_683);
nor U1031 (N_1031,N_697,N_618);
nor U1032 (N_1032,N_578,N_669);
and U1033 (N_1033,N_651,N_865);
xnor U1034 (N_1034,N_955,N_730);
nor U1035 (N_1035,N_921,N_508);
and U1036 (N_1036,N_660,N_691);
and U1037 (N_1037,N_533,N_716);
or U1038 (N_1038,N_539,N_584);
nor U1039 (N_1039,N_899,N_679);
and U1040 (N_1040,N_782,N_543);
nand U1041 (N_1041,N_762,N_765);
nand U1042 (N_1042,N_901,N_695);
or U1043 (N_1043,N_696,N_648);
and U1044 (N_1044,N_972,N_540);
nand U1045 (N_1045,N_672,N_744);
nor U1046 (N_1046,N_985,N_548);
nor U1047 (N_1047,N_872,N_753);
and U1048 (N_1048,N_801,N_729);
and U1049 (N_1049,N_877,N_980);
or U1050 (N_1050,N_986,N_757);
nand U1051 (N_1051,N_959,N_857);
or U1052 (N_1052,N_772,N_969);
and U1053 (N_1053,N_590,N_607);
nor U1054 (N_1054,N_774,N_993);
and U1055 (N_1055,N_947,N_694);
nand U1056 (N_1056,N_895,N_848);
xor U1057 (N_1057,N_882,N_823);
nor U1058 (N_1058,N_554,N_553);
nand U1059 (N_1059,N_853,N_665);
nor U1060 (N_1060,N_962,N_536);
or U1061 (N_1061,N_624,N_515);
nand U1062 (N_1062,N_907,N_807);
and U1063 (N_1063,N_994,N_926);
or U1064 (N_1064,N_605,N_677);
nor U1065 (N_1065,N_748,N_793);
or U1066 (N_1066,N_510,N_517);
or U1067 (N_1067,N_529,N_878);
and U1068 (N_1068,N_588,N_706);
and U1069 (N_1069,N_705,N_524);
or U1070 (N_1070,N_767,N_546);
nor U1071 (N_1071,N_996,N_968);
nand U1072 (N_1072,N_973,N_502);
or U1073 (N_1073,N_518,N_743);
nor U1074 (N_1074,N_531,N_826);
nand U1075 (N_1075,N_924,N_904);
or U1076 (N_1076,N_704,N_830);
or U1077 (N_1077,N_806,N_632);
and U1078 (N_1078,N_534,N_934);
or U1079 (N_1079,N_661,N_726);
and U1080 (N_1080,N_728,N_606);
nand U1081 (N_1081,N_698,N_770);
nor U1082 (N_1082,N_881,N_600);
or U1083 (N_1083,N_897,N_858);
nor U1084 (N_1084,N_840,N_559);
nor U1085 (N_1085,N_732,N_657);
and U1086 (N_1086,N_500,N_916);
and U1087 (N_1087,N_752,N_700);
nor U1088 (N_1088,N_789,N_951);
or U1089 (N_1089,N_535,N_981);
nor U1090 (N_1090,N_626,N_943);
or U1091 (N_1091,N_914,N_945);
nand U1092 (N_1092,N_771,N_875);
nand U1093 (N_1093,N_507,N_975);
and U1094 (N_1094,N_710,N_634);
nand U1095 (N_1095,N_889,N_982);
nand U1096 (N_1096,N_886,N_699);
nand U1097 (N_1097,N_796,N_711);
nor U1098 (N_1098,N_520,N_867);
nor U1099 (N_1099,N_760,N_738);
nand U1100 (N_1100,N_749,N_787);
nand U1101 (N_1101,N_756,N_741);
and U1102 (N_1102,N_864,N_894);
and U1103 (N_1103,N_769,N_971);
or U1104 (N_1104,N_572,N_784);
and U1105 (N_1105,N_861,N_623);
nand U1106 (N_1106,N_731,N_918);
nand U1107 (N_1107,N_976,N_866);
and U1108 (N_1108,N_599,N_977);
nand U1109 (N_1109,N_570,N_690);
and U1110 (N_1110,N_585,N_639);
and U1111 (N_1111,N_645,N_915);
and U1112 (N_1112,N_964,N_798);
or U1113 (N_1113,N_702,N_686);
and U1114 (N_1114,N_780,N_727);
nor U1115 (N_1115,N_558,N_619);
nor U1116 (N_1116,N_750,N_803);
and U1117 (N_1117,N_650,N_953);
and U1118 (N_1118,N_556,N_664);
or U1119 (N_1119,N_514,N_988);
xnor U1120 (N_1120,N_965,N_620);
and U1121 (N_1121,N_883,N_952);
and U1122 (N_1122,N_747,N_550);
xor U1123 (N_1123,N_602,N_850);
nor U1124 (N_1124,N_678,N_776);
or U1125 (N_1125,N_792,N_836);
nand U1126 (N_1126,N_885,N_995);
and U1127 (N_1127,N_876,N_908);
nand U1128 (N_1128,N_847,N_671);
nand U1129 (N_1129,N_598,N_715);
or U1130 (N_1130,N_862,N_999);
nand U1131 (N_1131,N_911,N_745);
or U1132 (N_1132,N_794,N_893);
or U1133 (N_1133,N_956,N_513);
or U1134 (N_1134,N_963,N_831);
nand U1135 (N_1135,N_828,N_763);
nor U1136 (N_1136,N_931,N_654);
nand U1137 (N_1137,N_997,N_936);
and U1138 (N_1138,N_984,N_551);
nor U1139 (N_1139,N_819,N_746);
and U1140 (N_1140,N_532,N_979);
and U1141 (N_1141,N_834,N_930);
or U1142 (N_1142,N_929,N_859);
or U1143 (N_1143,N_920,N_804);
or U1144 (N_1144,N_817,N_855);
or U1145 (N_1145,N_842,N_652);
or U1146 (N_1146,N_939,N_576);
nor U1147 (N_1147,N_687,N_575);
or U1148 (N_1148,N_912,N_863);
or U1149 (N_1149,N_583,N_670);
nor U1150 (N_1150,N_906,N_682);
and U1151 (N_1151,N_591,N_608);
or U1152 (N_1152,N_880,N_941);
nand U1153 (N_1153,N_755,N_966);
and U1154 (N_1154,N_560,N_887);
nand U1155 (N_1155,N_846,N_616);
nand U1156 (N_1156,N_809,N_563);
nand U1157 (N_1157,N_816,N_611);
or U1158 (N_1158,N_970,N_603);
and U1159 (N_1159,N_884,N_837);
and U1160 (N_1160,N_709,N_721);
nand U1161 (N_1161,N_668,N_516);
nor U1162 (N_1162,N_718,N_617);
and U1163 (N_1163,N_526,N_693);
and U1164 (N_1164,N_647,N_851);
nand U1165 (N_1165,N_856,N_948);
and U1166 (N_1166,N_754,N_557);
nor U1167 (N_1167,N_734,N_525);
nor U1168 (N_1168,N_662,N_905);
nor U1169 (N_1169,N_523,N_587);
xor U1170 (N_1170,N_902,N_562);
nand U1171 (N_1171,N_586,N_946);
nor U1172 (N_1172,N_854,N_839);
nor U1173 (N_1173,N_703,N_764);
xnor U1174 (N_1174,N_922,N_538);
and U1175 (N_1175,N_785,N_935);
nand U1176 (N_1176,N_589,N_824);
nand U1177 (N_1177,N_579,N_800);
nand U1178 (N_1178,N_635,N_612);
and U1179 (N_1179,N_549,N_987);
and U1180 (N_1180,N_613,N_835);
or U1181 (N_1181,N_720,N_811);
nand U1182 (N_1182,N_827,N_737);
or U1183 (N_1183,N_820,N_998);
and U1184 (N_1184,N_544,N_597);
nand U1185 (N_1185,N_675,N_501);
and U1186 (N_1186,N_910,N_949);
nand U1187 (N_1187,N_568,N_821);
nand U1188 (N_1188,N_768,N_815);
nor U1189 (N_1189,N_708,N_802);
nand U1190 (N_1190,N_937,N_829);
nand U1191 (N_1191,N_640,N_638);
nand U1192 (N_1192,N_667,N_595);
nand U1193 (N_1193,N_913,N_832);
nor U1194 (N_1194,N_621,N_565);
nand U1195 (N_1195,N_537,N_666);
or U1196 (N_1196,N_957,N_938);
and U1197 (N_1197,N_773,N_923);
or U1198 (N_1198,N_505,N_582);
and U1199 (N_1199,N_511,N_717);
or U1200 (N_1200,N_735,N_684);
nand U1201 (N_1201,N_814,N_992);
nand U1202 (N_1202,N_944,N_577);
nand U1203 (N_1203,N_519,N_564);
nor U1204 (N_1204,N_779,N_713);
and U1205 (N_1205,N_542,N_808);
and U1206 (N_1206,N_896,N_818);
and U1207 (N_1207,N_733,N_504);
nor U1208 (N_1208,N_723,N_566);
or U1209 (N_1209,N_644,N_596);
nand U1210 (N_1210,N_509,N_869);
nand U1211 (N_1211,N_701,N_673);
nand U1212 (N_1212,N_852,N_547);
and U1213 (N_1213,N_631,N_609);
nor U1214 (N_1214,N_751,N_642);
nand U1215 (N_1215,N_653,N_778);
or U1216 (N_1216,N_812,N_630);
nand U1217 (N_1217,N_530,N_932);
nand U1218 (N_1218,N_849,N_928);
or U1219 (N_1219,N_614,N_783);
and U1220 (N_1220,N_843,N_841);
or U1221 (N_1221,N_663,N_978);
and U1222 (N_1222,N_888,N_646);
and U1223 (N_1223,N_685,N_890);
nand U1224 (N_1224,N_552,N_528);
and U1225 (N_1225,N_571,N_805);
and U1226 (N_1226,N_874,N_942);
nor U1227 (N_1227,N_844,N_925);
nand U1228 (N_1228,N_799,N_637);
and U1229 (N_1229,N_892,N_909);
nand U1230 (N_1230,N_810,N_643);
xor U1231 (N_1231,N_775,N_633);
nand U1232 (N_1232,N_676,N_781);
and U1233 (N_1233,N_522,N_833);
nand U1234 (N_1234,N_879,N_658);
nor U1235 (N_1235,N_967,N_790);
or U1236 (N_1236,N_933,N_674);
or U1237 (N_1237,N_991,N_655);
xnor U1238 (N_1238,N_868,N_610);
nor U1239 (N_1239,N_680,N_659);
nor U1240 (N_1240,N_758,N_870);
nand U1241 (N_1241,N_983,N_919);
nand U1242 (N_1242,N_555,N_761);
or U1243 (N_1243,N_594,N_891);
and U1244 (N_1244,N_838,N_766);
and U1245 (N_1245,N_692,N_871);
nor U1246 (N_1246,N_521,N_900);
and U1247 (N_1247,N_580,N_722);
or U1248 (N_1248,N_641,N_822);
nand U1249 (N_1249,N_961,N_573);
nor U1250 (N_1250,N_768,N_797);
nor U1251 (N_1251,N_547,N_836);
or U1252 (N_1252,N_696,N_632);
nand U1253 (N_1253,N_698,N_969);
and U1254 (N_1254,N_975,N_755);
and U1255 (N_1255,N_564,N_610);
and U1256 (N_1256,N_608,N_858);
and U1257 (N_1257,N_687,N_993);
or U1258 (N_1258,N_533,N_766);
nor U1259 (N_1259,N_660,N_768);
or U1260 (N_1260,N_697,N_918);
nand U1261 (N_1261,N_506,N_853);
nor U1262 (N_1262,N_674,N_887);
nand U1263 (N_1263,N_814,N_996);
and U1264 (N_1264,N_623,N_602);
nand U1265 (N_1265,N_757,N_635);
and U1266 (N_1266,N_861,N_915);
and U1267 (N_1267,N_736,N_817);
or U1268 (N_1268,N_524,N_666);
and U1269 (N_1269,N_887,N_817);
and U1270 (N_1270,N_830,N_847);
and U1271 (N_1271,N_604,N_744);
nand U1272 (N_1272,N_917,N_589);
nor U1273 (N_1273,N_927,N_920);
nor U1274 (N_1274,N_867,N_805);
nor U1275 (N_1275,N_865,N_621);
nor U1276 (N_1276,N_941,N_573);
or U1277 (N_1277,N_856,N_936);
nor U1278 (N_1278,N_744,N_581);
nand U1279 (N_1279,N_521,N_675);
and U1280 (N_1280,N_827,N_577);
or U1281 (N_1281,N_935,N_522);
and U1282 (N_1282,N_705,N_889);
nor U1283 (N_1283,N_583,N_772);
nor U1284 (N_1284,N_620,N_736);
nand U1285 (N_1285,N_907,N_977);
or U1286 (N_1286,N_755,N_709);
nand U1287 (N_1287,N_535,N_614);
or U1288 (N_1288,N_603,N_802);
or U1289 (N_1289,N_593,N_747);
nand U1290 (N_1290,N_917,N_582);
nand U1291 (N_1291,N_682,N_809);
nand U1292 (N_1292,N_618,N_610);
and U1293 (N_1293,N_810,N_675);
and U1294 (N_1294,N_699,N_879);
and U1295 (N_1295,N_767,N_760);
or U1296 (N_1296,N_963,N_680);
nor U1297 (N_1297,N_895,N_759);
nor U1298 (N_1298,N_923,N_928);
xnor U1299 (N_1299,N_759,N_773);
nor U1300 (N_1300,N_980,N_981);
nand U1301 (N_1301,N_896,N_511);
nor U1302 (N_1302,N_918,N_609);
nor U1303 (N_1303,N_508,N_780);
nand U1304 (N_1304,N_588,N_865);
nor U1305 (N_1305,N_948,N_518);
or U1306 (N_1306,N_746,N_579);
nand U1307 (N_1307,N_968,N_742);
nand U1308 (N_1308,N_921,N_945);
nand U1309 (N_1309,N_937,N_822);
nor U1310 (N_1310,N_998,N_774);
or U1311 (N_1311,N_695,N_564);
nand U1312 (N_1312,N_900,N_728);
nor U1313 (N_1313,N_863,N_621);
or U1314 (N_1314,N_766,N_820);
and U1315 (N_1315,N_582,N_716);
nor U1316 (N_1316,N_911,N_915);
nand U1317 (N_1317,N_914,N_796);
and U1318 (N_1318,N_954,N_611);
or U1319 (N_1319,N_667,N_752);
nand U1320 (N_1320,N_512,N_615);
nand U1321 (N_1321,N_793,N_875);
and U1322 (N_1322,N_682,N_881);
xnor U1323 (N_1323,N_546,N_791);
and U1324 (N_1324,N_814,N_774);
nor U1325 (N_1325,N_509,N_786);
and U1326 (N_1326,N_640,N_700);
or U1327 (N_1327,N_554,N_773);
nand U1328 (N_1328,N_697,N_523);
nand U1329 (N_1329,N_703,N_581);
or U1330 (N_1330,N_603,N_817);
nand U1331 (N_1331,N_961,N_662);
nor U1332 (N_1332,N_511,N_687);
nor U1333 (N_1333,N_540,N_657);
and U1334 (N_1334,N_685,N_939);
nand U1335 (N_1335,N_594,N_614);
nor U1336 (N_1336,N_733,N_806);
and U1337 (N_1337,N_962,N_952);
nor U1338 (N_1338,N_950,N_696);
nor U1339 (N_1339,N_643,N_972);
and U1340 (N_1340,N_750,N_952);
xnor U1341 (N_1341,N_884,N_729);
nand U1342 (N_1342,N_509,N_802);
or U1343 (N_1343,N_805,N_860);
nor U1344 (N_1344,N_550,N_664);
nand U1345 (N_1345,N_793,N_595);
or U1346 (N_1346,N_503,N_805);
nor U1347 (N_1347,N_728,N_834);
or U1348 (N_1348,N_580,N_984);
xor U1349 (N_1349,N_914,N_691);
nor U1350 (N_1350,N_597,N_879);
or U1351 (N_1351,N_936,N_829);
nand U1352 (N_1352,N_590,N_976);
nand U1353 (N_1353,N_715,N_809);
nor U1354 (N_1354,N_876,N_670);
nand U1355 (N_1355,N_797,N_774);
or U1356 (N_1356,N_559,N_562);
or U1357 (N_1357,N_994,N_633);
or U1358 (N_1358,N_900,N_571);
nor U1359 (N_1359,N_863,N_696);
nor U1360 (N_1360,N_633,N_980);
or U1361 (N_1361,N_968,N_888);
nor U1362 (N_1362,N_634,N_872);
nand U1363 (N_1363,N_813,N_530);
and U1364 (N_1364,N_781,N_927);
nor U1365 (N_1365,N_667,N_855);
nor U1366 (N_1366,N_902,N_654);
nand U1367 (N_1367,N_837,N_771);
nor U1368 (N_1368,N_686,N_561);
or U1369 (N_1369,N_766,N_731);
and U1370 (N_1370,N_837,N_647);
nand U1371 (N_1371,N_531,N_607);
nand U1372 (N_1372,N_831,N_726);
nand U1373 (N_1373,N_666,N_808);
nor U1374 (N_1374,N_536,N_531);
or U1375 (N_1375,N_757,N_681);
or U1376 (N_1376,N_639,N_536);
nand U1377 (N_1377,N_919,N_541);
nor U1378 (N_1378,N_991,N_973);
xnor U1379 (N_1379,N_662,N_980);
nor U1380 (N_1380,N_763,N_500);
and U1381 (N_1381,N_790,N_798);
nand U1382 (N_1382,N_954,N_622);
nand U1383 (N_1383,N_611,N_616);
nand U1384 (N_1384,N_985,N_627);
and U1385 (N_1385,N_805,N_554);
or U1386 (N_1386,N_529,N_609);
nand U1387 (N_1387,N_543,N_528);
and U1388 (N_1388,N_773,N_669);
and U1389 (N_1389,N_789,N_697);
xor U1390 (N_1390,N_664,N_716);
nor U1391 (N_1391,N_752,N_717);
or U1392 (N_1392,N_897,N_626);
and U1393 (N_1393,N_765,N_840);
and U1394 (N_1394,N_790,N_587);
xnor U1395 (N_1395,N_622,N_741);
nand U1396 (N_1396,N_798,N_826);
or U1397 (N_1397,N_624,N_987);
nand U1398 (N_1398,N_986,N_651);
nor U1399 (N_1399,N_901,N_609);
or U1400 (N_1400,N_917,N_871);
nand U1401 (N_1401,N_811,N_901);
or U1402 (N_1402,N_958,N_509);
xor U1403 (N_1403,N_591,N_752);
nor U1404 (N_1404,N_894,N_511);
nand U1405 (N_1405,N_768,N_697);
or U1406 (N_1406,N_714,N_652);
xnor U1407 (N_1407,N_992,N_623);
nor U1408 (N_1408,N_991,N_949);
nand U1409 (N_1409,N_662,N_659);
and U1410 (N_1410,N_684,N_962);
nor U1411 (N_1411,N_652,N_807);
and U1412 (N_1412,N_634,N_519);
or U1413 (N_1413,N_826,N_536);
or U1414 (N_1414,N_528,N_787);
nand U1415 (N_1415,N_930,N_596);
nand U1416 (N_1416,N_965,N_865);
or U1417 (N_1417,N_509,N_754);
or U1418 (N_1418,N_932,N_807);
or U1419 (N_1419,N_605,N_822);
nand U1420 (N_1420,N_795,N_693);
nand U1421 (N_1421,N_957,N_784);
nand U1422 (N_1422,N_984,N_949);
and U1423 (N_1423,N_771,N_904);
nor U1424 (N_1424,N_612,N_673);
and U1425 (N_1425,N_896,N_960);
nor U1426 (N_1426,N_821,N_997);
or U1427 (N_1427,N_700,N_645);
or U1428 (N_1428,N_806,N_603);
or U1429 (N_1429,N_935,N_615);
nor U1430 (N_1430,N_655,N_796);
nor U1431 (N_1431,N_533,N_501);
nand U1432 (N_1432,N_589,N_758);
and U1433 (N_1433,N_825,N_814);
nand U1434 (N_1434,N_716,N_897);
nand U1435 (N_1435,N_867,N_996);
and U1436 (N_1436,N_724,N_845);
or U1437 (N_1437,N_718,N_603);
or U1438 (N_1438,N_884,N_947);
and U1439 (N_1439,N_956,N_967);
nor U1440 (N_1440,N_553,N_671);
or U1441 (N_1441,N_613,N_532);
or U1442 (N_1442,N_765,N_755);
nor U1443 (N_1443,N_942,N_599);
nand U1444 (N_1444,N_650,N_955);
nor U1445 (N_1445,N_647,N_649);
and U1446 (N_1446,N_561,N_948);
nor U1447 (N_1447,N_572,N_766);
nand U1448 (N_1448,N_544,N_556);
or U1449 (N_1449,N_917,N_720);
or U1450 (N_1450,N_791,N_633);
or U1451 (N_1451,N_987,N_938);
nand U1452 (N_1452,N_923,N_545);
or U1453 (N_1453,N_678,N_564);
or U1454 (N_1454,N_856,N_503);
nand U1455 (N_1455,N_604,N_749);
and U1456 (N_1456,N_674,N_926);
nand U1457 (N_1457,N_706,N_745);
and U1458 (N_1458,N_853,N_873);
or U1459 (N_1459,N_892,N_710);
xnor U1460 (N_1460,N_713,N_690);
xnor U1461 (N_1461,N_526,N_811);
nor U1462 (N_1462,N_937,N_979);
xor U1463 (N_1463,N_918,N_940);
nand U1464 (N_1464,N_647,N_571);
and U1465 (N_1465,N_806,N_582);
nor U1466 (N_1466,N_884,N_935);
nor U1467 (N_1467,N_517,N_827);
nand U1468 (N_1468,N_835,N_802);
nor U1469 (N_1469,N_903,N_832);
and U1470 (N_1470,N_517,N_768);
nor U1471 (N_1471,N_961,N_680);
nor U1472 (N_1472,N_984,N_532);
nand U1473 (N_1473,N_680,N_900);
and U1474 (N_1474,N_772,N_634);
xnor U1475 (N_1475,N_535,N_592);
or U1476 (N_1476,N_824,N_627);
nor U1477 (N_1477,N_619,N_852);
nand U1478 (N_1478,N_896,N_979);
nand U1479 (N_1479,N_751,N_833);
and U1480 (N_1480,N_703,N_905);
and U1481 (N_1481,N_925,N_516);
nand U1482 (N_1482,N_967,N_935);
nand U1483 (N_1483,N_722,N_800);
and U1484 (N_1484,N_895,N_878);
nand U1485 (N_1485,N_742,N_559);
or U1486 (N_1486,N_985,N_644);
and U1487 (N_1487,N_558,N_777);
nand U1488 (N_1488,N_510,N_923);
and U1489 (N_1489,N_714,N_974);
nand U1490 (N_1490,N_837,N_969);
or U1491 (N_1491,N_698,N_619);
nor U1492 (N_1492,N_618,N_784);
nor U1493 (N_1493,N_943,N_923);
and U1494 (N_1494,N_699,N_882);
or U1495 (N_1495,N_840,N_881);
and U1496 (N_1496,N_671,N_820);
nand U1497 (N_1497,N_537,N_565);
nand U1498 (N_1498,N_597,N_724);
nor U1499 (N_1499,N_831,N_766);
nand U1500 (N_1500,N_1427,N_1458);
nand U1501 (N_1501,N_1123,N_1037);
nor U1502 (N_1502,N_1159,N_1395);
or U1503 (N_1503,N_1069,N_1369);
nand U1504 (N_1504,N_1046,N_1317);
and U1505 (N_1505,N_1268,N_1213);
or U1506 (N_1506,N_1043,N_1156);
nor U1507 (N_1507,N_1264,N_1393);
and U1508 (N_1508,N_1426,N_1023);
or U1509 (N_1509,N_1236,N_1385);
nor U1510 (N_1510,N_1322,N_1184);
nor U1511 (N_1511,N_1402,N_1490);
and U1512 (N_1512,N_1176,N_1388);
nor U1513 (N_1513,N_1276,N_1495);
and U1514 (N_1514,N_1241,N_1047);
and U1515 (N_1515,N_1446,N_1051);
nand U1516 (N_1516,N_1094,N_1216);
nand U1517 (N_1517,N_1251,N_1075);
nor U1518 (N_1518,N_1468,N_1132);
nor U1519 (N_1519,N_1021,N_1074);
nand U1520 (N_1520,N_1137,N_1090);
and U1521 (N_1521,N_1163,N_1431);
or U1522 (N_1522,N_1259,N_1192);
and U1523 (N_1523,N_1497,N_1462);
and U1524 (N_1524,N_1136,N_1351);
nor U1525 (N_1525,N_1350,N_1048);
and U1526 (N_1526,N_1474,N_1027);
nor U1527 (N_1527,N_1188,N_1326);
and U1528 (N_1528,N_1076,N_1379);
nand U1529 (N_1529,N_1017,N_1275);
or U1530 (N_1530,N_1222,N_1151);
and U1531 (N_1531,N_1143,N_1339);
or U1532 (N_1532,N_1201,N_1135);
and U1533 (N_1533,N_1315,N_1300);
and U1534 (N_1534,N_1430,N_1429);
or U1535 (N_1535,N_1111,N_1425);
and U1536 (N_1536,N_1019,N_1318);
and U1537 (N_1537,N_1070,N_1496);
nand U1538 (N_1538,N_1091,N_1347);
and U1539 (N_1539,N_1072,N_1272);
nor U1540 (N_1540,N_1266,N_1104);
and U1541 (N_1541,N_1434,N_1432);
or U1542 (N_1542,N_1117,N_1316);
and U1543 (N_1543,N_1361,N_1340);
nor U1544 (N_1544,N_1063,N_1147);
and U1545 (N_1545,N_1185,N_1253);
nor U1546 (N_1546,N_1460,N_1146);
nor U1547 (N_1547,N_1308,N_1186);
nand U1548 (N_1548,N_1380,N_1145);
and U1549 (N_1549,N_1397,N_1482);
nor U1550 (N_1550,N_1270,N_1022);
or U1551 (N_1551,N_1126,N_1479);
and U1552 (N_1552,N_1193,N_1373);
nor U1553 (N_1553,N_1087,N_1071);
nand U1554 (N_1554,N_1119,N_1278);
nor U1555 (N_1555,N_1304,N_1148);
nor U1556 (N_1556,N_1089,N_1441);
or U1557 (N_1557,N_1486,N_1211);
and U1558 (N_1558,N_1194,N_1084);
nor U1559 (N_1559,N_1064,N_1436);
nor U1560 (N_1560,N_1455,N_1060);
or U1561 (N_1561,N_1416,N_1341);
xor U1562 (N_1562,N_1439,N_1245);
nand U1563 (N_1563,N_1144,N_1142);
nand U1564 (N_1564,N_1279,N_1025);
nand U1565 (N_1565,N_1453,N_1134);
nor U1566 (N_1566,N_1414,N_1115);
nand U1567 (N_1567,N_1269,N_1150);
nand U1568 (N_1568,N_1349,N_1165);
nor U1569 (N_1569,N_1169,N_1362);
nor U1570 (N_1570,N_1198,N_1483);
and U1571 (N_1571,N_1489,N_1418);
or U1572 (N_1572,N_1226,N_1312);
or U1573 (N_1573,N_1467,N_1381);
and U1574 (N_1574,N_1412,N_1372);
nor U1575 (N_1575,N_1271,N_1298);
or U1576 (N_1576,N_1499,N_1209);
and U1577 (N_1577,N_1422,N_1447);
and U1578 (N_1578,N_1195,N_1252);
nand U1579 (N_1579,N_1055,N_1190);
nor U1580 (N_1580,N_1086,N_1172);
nand U1581 (N_1581,N_1406,N_1153);
or U1582 (N_1582,N_1331,N_1191);
nor U1583 (N_1583,N_1386,N_1054);
or U1584 (N_1584,N_1413,N_1463);
nor U1585 (N_1585,N_1005,N_1428);
nand U1586 (N_1586,N_1327,N_1238);
nor U1587 (N_1587,N_1319,N_1199);
nor U1588 (N_1588,N_1139,N_1301);
and U1589 (N_1589,N_1020,N_1283);
nand U1590 (N_1590,N_1116,N_1102);
and U1591 (N_1591,N_1127,N_1344);
and U1592 (N_1592,N_1235,N_1109);
nor U1593 (N_1593,N_1012,N_1267);
and U1594 (N_1594,N_1470,N_1082);
or U1595 (N_1595,N_1358,N_1108);
and U1596 (N_1596,N_1256,N_1473);
or U1597 (N_1597,N_1212,N_1305);
nor U1598 (N_1598,N_1183,N_1067);
or U1599 (N_1599,N_1129,N_1049);
nand U1600 (N_1600,N_1174,N_1354);
or U1601 (N_1601,N_1178,N_1457);
or U1602 (N_1602,N_1099,N_1287);
or U1603 (N_1603,N_1461,N_1000);
nor U1604 (N_1604,N_1100,N_1481);
or U1605 (N_1605,N_1006,N_1103);
nor U1606 (N_1606,N_1477,N_1154);
nor U1607 (N_1607,N_1032,N_1417);
or U1608 (N_1608,N_1309,N_1208);
nor U1609 (N_1609,N_1478,N_1187);
nor U1610 (N_1610,N_1028,N_1130);
and U1611 (N_1611,N_1288,N_1166);
and U1612 (N_1612,N_1472,N_1387);
nor U1613 (N_1613,N_1491,N_1456);
nand U1614 (N_1614,N_1034,N_1400);
and U1615 (N_1615,N_1389,N_1263);
nor U1616 (N_1616,N_1175,N_1355);
nand U1617 (N_1617,N_1258,N_1015);
nor U1618 (N_1618,N_1262,N_1438);
or U1619 (N_1619,N_1036,N_1014);
and U1620 (N_1620,N_1371,N_1138);
nand U1621 (N_1621,N_1365,N_1376);
or U1622 (N_1622,N_1107,N_1407);
xor U1623 (N_1623,N_1110,N_1164);
nand U1624 (N_1624,N_1366,N_1242);
or U1625 (N_1625,N_1059,N_1040);
nor U1626 (N_1626,N_1367,N_1255);
xor U1627 (N_1627,N_1325,N_1133);
and U1628 (N_1628,N_1290,N_1336);
nor U1629 (N_1629,N_1405,N_1085);
or U1630 (N_1630,N_1415,N_1098);
or U1631 (N_1631,N_1273,N_1452);
or U1632 (N_1632,N_1122,N_1003);
or U1633 (N_1633,N_1112,N_1359);
or U1634 (N_1634,N_1357,N_1080);
nor U1635 (N_1635,N_1353,N_1485);
xor U1636 (N_1636,N_1443,N_1239);
or U1637 (N_1637,N_1128,N_1280);
nor U1638 (N_1638,N_1484,N_1228);
or U1639 (N_1639,N_1171,N_1469);
or U1640 (N_1640,N_1011,N_1092);
nor U1641 (N_1641,N_1050,N_1210);
or U1642 (N_1642,N_1487,N_1476);
xor U1643 (N_1643,N_1039,N_1338);
xor U1644 (N_1644,N_1437,N_1449);
nand U1645 (N_1645,N_1310,N_1056);
nand U1646 (N_1646,N_1261,N_1289);
or U1647 (N_1647,N_1205,N_1200);
nand U1648 (N_1648,N_1442,N_1281);
or U1649 (N_1649,N_1149,N_1311);
or U1650 (N_1650,N_1013,N_1364);
nor U1651 (N_1651,N_1291,N_1162);
or U1652 (N_1652,N_1155,N_1488);
nor U1653 (N_1653,N_1250,N_1282);
nand U1654 (N_1654,N_1314,N_1356);
and U1655 (N_1655,N_1424,N_1423);
and U1656 (N_1656,N_1120,N_1332);
nand U1657 (N_1657,N_1274,N_1403);
and U1658 (N_1658,N_1079,N_1494);
or U1659 (N_1659,N_1218,N_1324);
or U1660 (N_1660,N_1237,N_1173);
and U1661 (N_1661,N_1257,N_1161);
nor U1662 (N_1662,N_1044,N_1445);
and U1663 (N_1663,N_1152,N_1018);
and U1664 (N_1664,N_1420,N_1058);
nor U1665 (N_1665,N_1313,N_1010);
and U1666 (N_1666,N_1337,N_1454);
xnor U1667 (N_1667,N_1008,N_1330);
xnor U1668 (N_1668,N_1081,N_1065);
nor U1669 (N_1669,N_1292,N_1206);
nand U1670 (N_1670,N_1062,N_1328);
or U1671 (N_1671,N_1105,N_1181);
nand U1672 (N_1672,N_1382,N_1125);
and U1673 (N_1673,N_1234,N_1002);
and U1674 (N_1674,N_1342,N_1247);
nor U1675 (N_1675,N_1464,N_1296);
nor U1676 (N_1676,N_1384,N_1493);
nor U1677 (N_1677,N_1124,N_1217);
and U1678 (N_1678,N_1392,N_1243);
and U1679 (N_1679,N_1167,N_1480);
and U1680 (N_1680,N_1360,N_1118);
nand U1681 (N_1681,N_1374,N_1249);
and U1682 (N_1682,N_1009,N_1160);
or U1683 (N_1683,N_1223,N_1035);
nor U1684 (N_1684,N_1204,N_1303);
and U1685 (N_1685,N_1345,N_1399);
nand U1686 (N_1686,N_1302,N_1240);
and U1687 (N_1687,N_1227,N_1346);
nand U1688 (N_1688,N_1421,N_1073);
nor U1689 (N_1689,N_1260,N_1435);
and U1690 (N_1690,N_1401,N_1244);
nor U1691 (N_1691,N_1299,N_1293);
and U1692 (N_1692,N_1471,N_1229);
nor U1693 (N_1693,N_1207,N_1096);
nor U1694 (N_1694,N_1246,N_1335);
or U1695 (N_1695,N_1179,N_1277);
and U1696 (N_1696,N_1170,N_1265);
or U1697 (N_1697,N_1077,N_1320);
nand U1698 (N_1698,N_1294,N_1450);
nand U1699 (N_1699,N_1113,N_1114);
or U1700 (N_1700,N_1329,N_1042);
and U1701 (N_1701,N_1041,N_1232);
xnor U1702 (N_1702,N_1097,N_1492);
and U1703 (N_1703,N_1038,N_1307);
xnor U1704 (N_1704,N_1131,N_1408);
xor U1705 (N_1705,N_1377,N_1498);
and U1706 (N_1706,N_1088,N_1383);
nor U1707 (N_1707,N_1202,N_1220);
and U1708 (N_1708,N_1189,N_1370);
and U1709 (N_1709,N_1323,N_1121);
nand U1710 (N_1710,N_1158,N_1396);
or U1711 (N_1711,N_1285,N_1451);
nand U1712 (N_1712,N_1398,N_1045);
nand U1713 (N_1713,N_1219,N_1033);
nand U1714 (N_1714,N_1286,N_1016);
and U1715 (N_1715,N_1404,N_1391);
or U1716 (N_1716,N_1101,N_1203);
and U1717 (N_1717,N_1001,N_1093);
and U1718 (N_1718,N_1057,N_1053);
or U1719 (N_1719,N_1007,N_1410);
nand U1720 (N_1720,N_1168,N_1106);
or U1721 (N_1721,N_1475,N_1052);
nor U1722 (N_1722,N_1180,N_1409);
nor U1723 (N_1723,N_1177,N_1182);
or U1724 (N_1724,N_1368,N_1433);
or U1725 (N_1725,N_1214,N_1068);
nor U1726 (N_1726,N_1031,N_1459);
nor U1727 (N_1727,N_1378,N_1141);
nand U1728 (N_1728,N_1343,N_1061);
nand U1729 (N_1729,N_1224,N_1363);
nand U1730 (N_1730,N_1348,N_1248);
nor U1731 (N_1731,N_1221,N_1352);
and U1732 (N_1732,N_1419,N_1334);
and U1733 (N_1733,N_1024,N_1026);
and U1734 (N_1734,N_1230,N_1225);
or U1735 (N_1735,N_1197,N_1004);
nand U1736 (N_1736,N_1394,N_1306);
or U1737 (N_1737,N_1066,N_1321);
nand U1738 (N_1738,N_1231,N_1254);
nor U1739 (N_1739,N_1095,N_1297);
or U1740 (N_1740,N_1444,N_1157);
or U1741 (N_1741,N_1030,N_1233);
and U1742 (N_1742,N_1295,N_1284);
or U1743 (N_1743,N_1215,N_1440);
xnor U1744 (N_1744,N_1448,N_1390);
and U1745 (N_1745,N_1140,N_1078);
and U1746 (N_1746,N_1029,N_1083);
or U1747 (N_1747,N_1196,N_1466);
nor U1748 (N_1748,N_1333,N_1375);
and U1749 (N_1749,N_1465,N_1411);
and U1750 (N_1750,N_1353,N_1250);
or U1751 (N_1751,N_1344,N_1078);
nand U1752 (N_1752,N_1017,N_1449);
nor U1753 (N_1753,N_1463,N_1013);
nor U1754 (N_1754,N_1413,N_1088);
or U1755 (N_1755,N_1342,N_1337);
nand U1756 (N_1756,N_1430,N_1143);
nand U1757 (N_1757,N_1489,N_1120);
nand U1758 (N_1758,N_1302,N_1361);
nand U1759 (N_1759,N_1256,N_1109);
nor U1760 (N_1760,N_1464,N_1383);
or U1761 (N_1761,N_1071,N_1132);
nor U1762 (N_1762,N_1209,N_1160);
nor U1763 (N_1763,N_1028,N_1099);
nand U1764 (N_1764,N_1329,N_1450);
and U1765 (N_1765,N_1306,N_1122);
and U1766 (N_1766,N_1147,N_1217);
or U1767 (N_1767,N_1413,N_1029);
nand U1768 (N_1768,N_1471,N_1402);
and U1769 (N_1769,N_1187,N_1405);
and U1770 (N_1770,N_1426,N_1009);
and U1771 (N_1771,N_1342,N_1111);
nand U1772 (N_1772,N_1451,N_1169);
and U1773 (N_1773,N_1478,N_1487);
and U1774 (N_1774,N_1232,N_1218);
or U1775 (N_1775,N_1477,N_1326);
or U1776 (N_1776,N_1116,N_1010);
or U1777 (N_1777,N_1210,N_1039);
or U1778 (N_1778,N_1002,N_1431);
nor U1779 (N_1779,N_1022,N_1257);
or U1780 (N_1780,N_1121,N_1395);
and U1781 (N_1781,N_1298,N_1401);
or U1782 (N_1782,N_1140,N_1168);
nor U1783 (N_1783,N_1068,N_1141);
nand U1784 (N_1784,N_1071,N_1495);
or U1785 (N_1785,N_1490,N_1168);
and U1786 (N_1786,N_1299,N_1121);
nor U1787 (N_1787,N_1344,N_1389);
or U1788 (N_1788,N_1475,N_1351);
nor U1789 (N_1789,N_1202,N_1209);
or U1790 (N_1790,N_1387,N_1456);
nor U1791 (N_1791,N_1183,N_1271);
or U1792 (N_1792,N_1307,N_1253);
or U1793 (N_1793,N_1144,N_1252);
nand U1794 (N_1794,N_1017,N_1137);
and U1795 (N_1795,N_1404,N_1411);
and U1796 (N_1796,N_1406,N_1178);
nand U1797 (N_1797,N_1038,N_1257);
or U1798 (N_1798,N_1183,N_1105);
nand U1799 (N_1799,N_1424,N_1044);
or U1800 (N_1800,N_1096,N_1457);
or U1801 (N_1801,N_1044,N_1385);
nand U1802 (N_1802,N_1142,N_1247);
and U1803 (N_1803,N_1123,N_1270);
or U1804 (N_1804,N_1394,N_1150);
nor U1805 (N_1805,N_1067,N_1201);
nor U1806 (N_1806,N_1258,N_1444);
nand U1807 (N_1807,N_1477,N_1142);
nand U1808 (N_1808,N_1165,N_1009);
nor U1809 (N_1809,N_1468,N_1396);
and U1810 (N_1810,N_1029,N_1117);
or U1811 (N_1811,N_1038,N_1001);
and U1812 (N_1812,N_1384,N_1420);
nor U1813 (N_1813,N_1284,N_1406);
nor U1814 (N_1814,N_1090,N_1038);
nor U1815 (N_1815,N_1239,N_1412);
or U1816 (N_1816,N_1245,N_1040);
or U1817 (N_1817,N_1472,N_1058);
nor U1818 (N_1818,N_1187,N_1155);
nand U1819 (N_1819,N_1212,N_1036);
and U1820 (N_1820,N_1316,N_1199);
or U1821 (N_1821,N_1004,N_1315);
and U1822 (N_1822,N_1420,N_1328);
or U1823 (N_1823,N_1088,N_1346);
and U1824 (N_1824,N_1124,N_1197);
and U1825 (N_1825,N_1417,N_1345);
and U1826 (N_1826,N_1340,N_1256);
nand U1827 (N_1827,N_1358,N_1205);
nor U1828 (N_1828,N_1381,N_1295);
nor U1829 (N_1829,N_1226,N_1470);
or U1830 (N_1830,N_1404,N_1152);
nand U1831 (N_1831,N_1450,N_1245);
nand U1832 (N_1832,N_1389,N_1230);
and U1833 (N_1833,N_1466,N_1148);
nand U1834 (N_1834,N_1094,N_1071);
or U1835 (N_1835,N_1172,N_1291);
and U1836 (N_1836,N_1304,N_1057);
and U1837 (N_1837,N_1065,N_1061);
xor U1838 (N_1838,N_1274,N_1148);
or U1839 (N_1839,N_1016,N_1201);
nand U1840 (N_1840,N_1110,N_1438);
or U1841 (N_1841,N_1399,N_1298);
and U1842 (N_1842,N_1277,N_1138);
and U1843 (N_1843,N_1261,N_1299);
nand U1844 (N_1844,N_1149,N_1274);
and U1845 (N_1845,N_1451,N_1369);
nor U1846 (N_1846,N_1084,N_1315);
and U1847 (N_1847,N_1367,N_1323);
or U1848 (N_1848,N_1271,N_1065);
or U1849 (N_1849,N_1129,N_1446);
or U1850 (N_1850,N_1226,N_1025);
nand U1851 (N_1851,N_1099,N_1489);
or U1852 (N_1852,N_1444,N_1353);
and U1853 (N_1853,N_1080,N_1391);
or U1854 (N_1854,N_1189,N_1031);
nor U1855 (N_1855,N_1116,N_1179);
nand U1856 (N_1856,N_1119,N_1466);
nor U1857 (N_1857,N_1228,N_1311);
or U1858 (N_1858,N_1466,N_1445);
or U1859 (N_1859,N_1260,N_1478);
and U1860 (N_1860,N_1262,N_1498);
nor U1861 (N_1861,N_1482,N_1039);
or U1862 (N_1862,N_1421,N_1360);
or U1863 (N_1863,N_1262,N_1396);
nand U1864 (N_1864,N_1151,N_1369);
and U1865 (N_1865,N_1292,N_1386);
nand U1866 (N_1866,N_1220,N_1498);
or U1867 (N_1867,N_1410,N_1260);
and U1868 (N_1868,N_1218,N_1270);
nor U1869 (N_1869,N_1095,N_1404);
nor U1870 (N_1870,N_1028,N_1475);
and U1871 (N_1871,N_1397,N_1284);
nor U1872 (N_1872,N_1273,N_1483);
nand U1873 (N_1873,N_1304,N_1086);
nor U1874 (N_1874,N_1281,N_1449);
and U1875 (N_1875,N_1075,N_1240);
and U1876 (N_1876,N_1039,N_1424);
and U1877 (N_1877,N_1302,N_1067);
or U1878 (N_1878,N_1416,N_1110);
nand U1879 (N_1879,N_1258,N_1147);
and U1880 (N_1880,N_1093,N_1254);
nor U1881 (N_1881,N_1041,N_1358);
or U1882 (N_1882,N_1025,N_1394);
xnor U1883 (N_1883,N_1356,N_1124);
or U1884 (N_1884,N_1289,N_1052);
or U1885 (N_1885,N_1371,N_1192);
nor U1886 (N_1886,N_1415,N_1133);
or U1887 (N_1887,N_1275,N_1038);
xnor U1888 (N_1888,N_1214,N_1275);
nand U1889 (N_1889,N_1214,N_1322);
or U1890 (N_1890,N_1114,N_1052);
nor U1891 (N_1891,N_1022,N_1135);
nand U1892 (N_1892,N_1479,N_1442);
nand U1893 (N_1893,N_1312,N_1478);
and U1894 (N_1894,N_1459,N_1391);
and U1895 (N_1895,N_1338,N_1189);
nor U1896 (N_1896,N_1420,N_1070);
nand U1897 (N_1897,N_1013,N_1495);
or U1898 (N_1898,N_1247,N_1056);
or U1899 (N_1899,N_1321,N_1456);
or U1900 (N_1900,N_1440,N_1277);
nand U1901 (N_1901,N_1394,N_1489);
nand U1902 (N_1902,N_1194,N_1154);
nand U1903 (N_1903,N_1278,N_1218);
xnor U1904 (N_1904,N_1182,N_1152);
nand U1905 (N_1905,N_1252,N_1344);
and U1906 (N_1906,N_1047,N_1111);
nand U1907 (N_1907,N_1047,N_1082);
or U1908 (N_1908,N_1058,N_1005);
nor U1909 (N_1909,N_1208,N_1037);
or U1910 (N_1910,N_1348,N_1325);
nand U1911 (N_1911,N_1288,N_1033);
nand U1912 (N_1912,N_1110,N_1133);
and U1913 (N_1913,N_1244,N_1393);
nor U1914 (N_1914,N_1039,N_1303);
nand U1915 (N_1915,N_1108,N_1087);
xor U1916 (N_1916,N_1341,N_1182);
nand U1917 (N_1917,N_1267,N_1472);
or U1918 (N_1918,N_1412,N_1191);
or U1919 (N_1919,N_1095,N_1158);
nor U1920 (N_1920,N_1130,N_1499);
or U1921 (N_1921,N_1256,N_1284);
nand U1922 (N_1922,N_1300,N_1330);
or U1923 (N_1923,N_1031,N_1066);
or U1924 (N_1924,N_1396,N_1071);
nand U1925 (N_1925,N_1040,N_1459);
xor U1926 (N_1926,N_1372,N_1391);
xnor U1927 (N_1927,N_1370,N_1089);
nor U1928 (N_1928,N_1275,N_1134);
nor U1929 (N_1929,N_1055,N_1121);
and U1930 (N_1930,N_1197,N_1273);
and U1931 (N_1931,N_1337,N_1136);
nand U1932 (N_1932,N_1313,N_1295);
and U1933 (N_1933,N_1037,N_1034);
nand U1934 (N_1934,N_1338,N_1485);
nor U1935 (N_1935,N_1263,N_1401);
and U1936 (N_1936,N_1118,N_1388);
and U1937 (N_1937,N_1347,N_1358);
nor U1938 (N_1938,N_1085,N_1307);
and U1939 (N_1939,N_1238,N_1080);
or U1940 (N_1940,N_1393,N_1141);
or U1941 (N_1941,N_1025,N_1115);
and U1942 (N_1942,N_1055,N_1194);
nor U1943 (N_1943,N_1234,N_1328);
and U1944 (N_1944,N_1287,N_1144);
nor U1945 (N_1945,N_1292,N_1040);
nor U1946 (N_1946,N_1236,N_1240);
nand U1947 (N_1947,N_1281,N_1419);
nand U1948 (N_1948,N_1295,N_1232);
nand U1949 (N_1949,N_1425,N_1089);
nand U1950 (N_1950,N_1219,N_1348);
and U1951 (N_1951,N_1109,N_1075);
and U1952 (N_1952,N_1373,N_1114);
nand U1953 (N_1953,N_1407,N_1289);
or U1954 (N_1954,N_1027,N_1174);
or U1955 (N_1955,N_1312,N_1050);
nor U1956 (N_1956,N_1222,N_1297);
and U1957 (N_1957,N_1435,N_1410);
or U1958 (N_1958,N_1255,N_1257);
and U1959 (N_1959,N_1470,N_1419);
or U1960 (N_1960,N_1159,N_1434);
or U1961 (N_1961,N_1057,N_1218);
nor U1962 (N_1962,N_1266,N_1019);
nand U1963 (N_1963,N_1282,N_1026);
nor U1964 (N_1964,N_1343,N_1196);
and U1965 (N_1965,N_1475,N_1455);
nand U1966 (N_1966,N_1316,N_1479);
nor U1967 (N_1967,N_1345,N_1456);
and U1968 (N_1968,N_1309,N_1067);
or U1969 (N_1969,N_1474,N_1276);
nand U1970 (N_1970,N_1466,N_1000);
nand U1971 (N_1971,N_1303,N_1310);
nand U1972 (N_1972,N_1315,N_1055);
xor U1973 (N_1973,N_1359,N_1185);
and U1974 (N_1974,N_1455,N_1442);
nand U1975 (N_1975,N_1213,N_1440);
and U1976 (N_1976,N_1187,N_1368);
or U1977 (N_1977,N_1106,N_1298);
nor U1978 (N_1978,N_1201,N_1467);
or U1979 (N_1979,N_1363,N_1084);
nand U1980 (N_1980,N_1400,N_1110);
nand U1981 (N_1981,N_1306,N_1168);
or U1982 (N_1982,N_1493,N_1373);
and U1983 (N_1983,N_1068,N_1160);
or U1984 (N_1984,N_1044,N_1191);
and U1985 (N_1985,N_1148,N_1423);
nand U1986 (N_1986,N_1010,N_1169);
nand U1987 (N_1987,N_1184,N_1402);
and U1988 (N_1988,N_1033,N_1174);
nor U1989 (N_1989,N_1111,N_1136);
nor U1990 (N_1990,N_1297,N_1313);
nand U1991 (N_1991,N_1166,N_1289);
nor U1992 (N_1992,N_1174,N_1243);
nand U1993 (N_1993,N_1027,N_1078);
nand U1994 (N_1994,N_1284,N_1031);
or U1995 (N_1995,N_1221,N_1425);
or U1996 (N_1996,N_1301,N_1358);
nand U1997 (N_1997,N_1353,N_1235);
nand U1998 (N_1998,N_1483,N_1353);
nor U1999 (N_1999,N_1314,N_1453);
and U2000 (N_2000,N_1718,N_1655);
nand U2001 (N_2001,N_1566,N_1797);
nor U2002 (N_2002,N_1991,N_1968);
and U2003 (N_2003,N_1769,N_1876);
or U2004 (N_2004,N_1736,N_1780);
nor U2005 (N_2005,N_1530,N_1904);
and U2006 (N_2006,N_1843,N_1809);
nor U2007 (N_2007,N_1546,N_1726);
nor U2008 (N_2008,N_1686,N_1603);
xnor U2009 (N_2009,N_1649,N_1856);
and U2010 (N_2010,N_1709,N_1668);
or U2011 (N_2011,N_1994,N_1810);
and U2012 (N_2012,N_1969,N_1771);
or U2013 (N_2013,N_1798,N_1805);
nand U2014 (N_2014,N_1785,N_1784);
nor U2015 (N_2015,N_1695,N_1815);
xnor U2016 (N_2016,N_1567,N_1703);
or U2017 (N_2017,N_1953,N_1727);
and U2018 (N_2018,N_1976,N_1787);
xnor U2019 (N_2019,N_1658,N_1517);
or U2020 (N_2020,N_1552,N_1910);
nand U2021 (N_2021,N_1975,N_1939);
or U2022 (N_2022,N_1987,N_1540);
or U2023 (N_2023,N_1715,N_1515);
nand U2024 (N_2024,N_1898,N_1775);
or U2025 (N_2025,N_1622,N_1527);
nand U2026 (N_2026,N_1753,N_1738);
nor U2027 (N_2027,N_1503,N_1937);
nor U2028 (N_2028,N_1674,N_1841);
nor U2029 (N_2029,N_1593,N_1525);
or U2030 (N_2030,N_1516,N_1831);
nand U2031 (N_2031,N_1601,N_1906);
or U2032 (N_2032,N_1756,N_1547);
nand U2033 (N_2033,N_1807,N_1538);
nand U2034 (N_2034,N_1650,N_1730);
and U2035 (N_2035,N_1701,N_1721);
nor U2036 (N_2036,N_1893,N_1950);
and U2037 (N_2037,N_1694,N_1744);
and U2038 (N_2038,N_1544,N_1732);
nand U2039 (N_2039,N_1734,N_1852);
and U2040 (N_2040,N_1737,N_1513);
and U2041 (N_2041,N_1778,N_1571);
nor U2042 (N_2042,N_1642,N_1645);
nor U2043 (N_2043,N_1746,N_1681);
and U2044 (N_2044,N_1687,N_1750);
nor U2045 (N_2045,N_1887,N_1951);
nor U2046 (N_2046,N_1862,N_1811);
nor U2047 (N_2047,N_1510,N_1661);
or U2048 (N_2048,N_1886,N_1758);
and U2049 (N_2049,N_1980,N_1685);
and U2050 (N_2050,N_1929,N_1783);
and U2051 (N_2051,N_1691,N_1760);
nor U2052 (N_2052,N_1713,N_1712);
nand U2053 (N_2053,N_1764,N_1553);
or U2054 (N_2054,N_1639,N_1558);
and U2055 (N_2055,N_1648,N_1837);
nand U2056 (N_2056,N_1696,N_1500);
and U2057 (N_2057,N_1605,N_1936);
nor U2058 (N_2058,N_1542,N_1640);
nand U2059 (N_2059,N_1839,N_1946);
or U2060 (N_2060,N_1877,N_1609);
and U2061 (N_2061,N_1844,N_1617);
nor U2062 (N_2062,N_1702,N_1773);
nand U2063 (N_2063,N_1519,N_1960);
and U2064 (N_2064,N_1786,N_1801);
or U2065 (N_2065,N_1792,N_1847);
or U2066 (N_2066,N_1993,N_1526);
nor U2067 (N_2067,N_1990,N_1903);
or U2068 (N_2068,N_1874,N_1952);
and U2069 (N_2069,N_1618,N_1920);
nor U2070 (N_2070,N_1570,N_1644);
nand U2071 (N_2071,N_1997,N_1978);
nor U2072 (N_2072,N_1679,N_1620);
and U2073 (N_2073,N_1717,N_1914);
and U2074 (N_2074,N_1878,N_1708);
nand U2075 (N_2075,N_1625,N_1610);
nand U2076 (N_2076,N_1961,N_1537);
nor U2077 (N_2077,N_1791,N_1671);
nand U2078 (N_2078,N_1849,N_1666);
nand U2079 (N_2079,N_1999,N_1629);
nor U2080 (N_2080,N_1819,N_1949);
nor U2081 (N_2081,N_1740,N_1632);
nand U2082 (N_2082,N_1654,N_1659);
nor U2083 (N_2083,N_1556,N_1896);
and U2084 (N_2084,N_1590,N_1673);
nand U2085 (N_2085,N_1697,N_1591);
nand U2086 (N_2086,N_1521,N_1966);
or U2087 (N_2087,N_1782,N_1984);
nor U2088 (N_2088,N_1858,N_1665);
xor U2089 (N_2089,N_1885,N_1833);
and U2090 (N_2090,N_1834,N_1677);
and U2091 (N_2091,N_1619,N_1643);
nand U2092 (N_2092,N_1962,N_1594);
nand U2093 (N_2093,N_1635,N_1765);
nor U2094 (N_2094,N_1582,N_1514);
and U2095 (N_2095,N_1845,N_1508);
and U2096 (N_2096,N_1706,N_1930);
nand U2097 (N_2097,N_1502,N_1892);
nor U2098 (N_2098,N_1770,N_1985);
nand U2099 (N_2099,N_1762,N_1989);
nand U2100 (N_2100,N_1548,N_1549);
and U2101 (N_2101,N_1623,N_1828);
or U2102 (N_2102,N_1584,N_1955);
and U2103 (N_2103,N_1634,N_1690);
and U2104 (N_2104,N_1529,N_1647);
and U2105 (N_2105,N_1789,N_1859);
or U2106 (N_2106,N_1585,N_1743);
nor U2107 (N_2107,N_1631,N_1539);
nor U2108 (N_2108,N_1501,N_1842);
nand U2109 (N_2109,N_1922,N_1924);
nor U2110 (N_2110,N_1759,N_1931);
or U2111 (N_2111,N_1865,N_1722);
nand U2112 (N_2112,N_1875,N_1574);
and U2113 (N_2113,N_1522,N_1751);
xor U2114 (N_2114,N_1820,N_1698);
and U2115 (N_2115,N_1853,N_1505);
nor U2116 (N_2116,N_1871,N_1693);
nor U2117 (N_2117,N_1626,N_1755);
or U2118 (N_2118,N_1680,N_1818);
nor U2119 (N_2119,N_1506,N_1921);
nand U2120 (N_2120,N_1586,N_1915);
nor U2121 (N_2121,N_1672,N_1814);
nand U2122 (N_2122,N_1891,N_1919);
nor U2123 (N_2123,N_1664,N_1656);
nor U2124 (N_2124,N_1925,N_1534);
nand U2125 (N_2125,N_1869,N_1944);
xor U2126 (N_2126,N_1653,N_1804);
or U2127 (N_2127,N_1683,N_1675);
or U2128 (N_2128,N_1676,N_1559);
nor U2129 (N_2129,N_1550,N_1796);
nand U2130 (N_2130,N_1943,N_1900);
nor U2131 (N_2131,N_1739,N_1568);
nand U2132 (N_2132,N_1688,N_1776);
and U2133 (N_2133,N_1940,N_1562);
nor U2134 (N_2134,N_1909,N_1541);
or U2135 (N_2135,N_1684,N_1882);
or U2136 (N_2136,N_1870,N_1587);
nand U2137 (N_2137,N_1724,N_1954);
nand U2138 (N_2138,N_1748,N_1965);
and U2139 (N_2139,N_1829,N_1816);
and U2140 (N_2140,N_1614,N_1580);
nor U2141 (N_2141,N_1560,N_1627);
xor U2142 (N_2142,N_1646,N_1890);
or U2143 (N_2143,N_1860,N_1967);
or U2144 (N_2144,N_1995,N_1793);
nand U2145 (N_2145,N_1723,N_1512);
and U2146 (N_2146,N_1504,N_1868);
nor U2147 (N_2147,N_1699,N_1597);
nor U2148 (N_2148,N_1667,N_1509);
nand U2149 (N_2149,N_1602,N_1857);
or U2150 (N_2150,N_1689,N_1971);
or U2151 (N_2151,N_1604,N_1660);
nand U2152 (N_2152,N_1777,N_1557);
xnor U2153 (N_2153,N_1880,N_1678);
nand U2154 (N_2154,N_1799,N_1823);
or U2155 (N_2155,N_1523,N_1575);
nor U2156 (N_2156,N_1902,N_1728);
or U2157 (N_2157,N_1872,N_1941);
nor U2158 (N_2158,N_1908,N_1576);
nor U2159 (N_2159,N_1945,N_1827);
nand U2160 (N_2160,N_1926,N_1711);
and U2161 (N_2161,N_1774,N_1986);
nand U2162 (N_2162,N_1611,N_1670);
or U2163 (N_2163,N_1733,N_1754);
or U2164 (N_2164,N_1752,N_1535);
and U2165 (N_2165,N_1735,N_1628);
nand U2166 (N_2166,N_1923,N_1982);
or U2167 (N_2167,N_1867,N_1633);
nand U2168 (N_2168,N_1565,N_1918);
nor U2169 (N_2169,N_1824,N_1613);
or U2170 (N_2170,N_1573,N_1636);
and U2171 (N_2171,N_1608,N_1979);
and U2172 (N_2172,N_1731,N_1825);
nor U2173 (N_2173,N_1977,N_1577);
nand U2174 (N_2174,N_1884,N_1719);
and U2175 (N_2175,N_1600,N_1947);
nor U2176 (N_2176,N_1894,N_1864);
nand U2177 (N_2177,N_1772,N_1981);
nor U2178 (N_2178,N_1830,N_1964);
and U2179 (N_2179,N_1928,N_1911);
nor U2180 (N_2180,N_1912,N_1551);
or U2181 (N_2181,N_1963,N_1705);
or U2182 (N_2182,N_1897,N_1532);
xnor U2183 (N_2183,N_1790,N_1511);
nor U2184 (N_2184,N_1707,N_1996);
nor U2185 (N_2185,N_1564,N_1881);
nand U2186 (N_2186,N_1662,N_1934);
and U2187 (N_2187,N_1518,N_1927);
and U2188 (N_2188,N_1742,N_1795);
nand U2189 (N_2189,N_1832,N_1866);
or U2190 (N_2190,N_1888,N_1861);
or U2191 (N_2191,N_1913,N_1835);
nand U2192 (N_2192,N_1901,N_1958);
nand U2193 (N_2193,N_1873,N_1607);
xor U2194 (N_2194,N_1716,N_1763);
or U2195 (N_2195,N_1612,N_1592);
or U2196 (N_2196,N_1616,N_1779);
and U2197 (N_2197,N_1651,N_1581);
and U2198 (N_2198,N_1578,N_1531);
nor U2199 (N_2199,N_1794,N_1561);
or U2200 (N_2200,N_1745,N_1766);
nor U2201 (N_2201,N_1767,N_1595);
nor U2202 (N_2202,N_1879,N_1883);
nor U2203 (N_2203,N_1781,N_1528);
and U2204 (N_2204,N_1983,N_1932);
nor U2205 (N_2205,N_1589,N_1998);
nand U2206 (N_2206,N_1822,N_1579);
or U2207 (N_2207,N_1768,N_1641);
or U2208 (N_2208,N_1638,N_1714);
or U2209 (N_2209,N_1813,N_1851);
nand U2210 (N_2210,N_1899,N_1555);
nand U2211 (N_2211,N_1855,N_1916);
and U2212 (N_2212,N_1637,N_1554);
nand U2213 (N_2213,N_1729,N_1536);
or U2214 (N_2214,N_1583,N_1907);
nand U2215 (N_2215,N_1917,N_1757);
nor U2216 (N_2216,N_1572,N_1817);
nor U2217 (N_2217,N_1682,N_1970);
nor U2218 (N_2218,N_1854,N_1808);
nor U2219 (N_2219,N_1704,N_1692);
nor U2220 (N_2220,N_1948,N_1957);
nor U2221 (N_2221,N_1935,N_1889);
nor U2222 (N_2222,N_1850,N_1725);
nand U2223 (N_2223,N_1630,N_1588);
and U2224 (N_2224,N_1507,N_1710);
or U2225 (N_2225,N_1959,N_1598);
or U2226 (N_2226,N_1563,N_1826);
nor U2227 (N_2227,N_1974,N_1599);
nor U2228 (N_2228,N_1652,N_1520);
nor U2229 (N_2229,N_1596,N_1988);
or U2230 (N_2230,N_1615,N_1992);
xor U2231 (N_2231,N_1543,N_1621);
nor U2232 (N_2232,N_1720,N_1741);
or U2233 (N_2233,N_1942,N_1848);
and U2234 (N_2234,N_1806,N_1524);
or U2235 (N_2235,N_1812,N_1545);
and U2236 (N_2236,N_1800,N_1933);
nor U2237 (N_2237,N_1938,N_1972);
or U2238 (N_2238,N_1533,N_1840);
nand U2239 (N_2239,N_1749,N_1700);
nand U2240 (N_2240,N_1863,N_1803);
or U2241 (N_2241,N_1802,N_1761);
nand U2242 (N_2242,N_1838,N_1788);
nor U2243 (N_2243,N_1956,N_1836);
nor U2244 (N_2244,N_1606,N_1846);
nand U2245 (N_2245,N_1669,N_1895);
nor U2246 (N_2246,N_1747,N_1569);
or U2247 (N_2247,N_1821,N_1973);
nand U2248 (N_2248,N_1663,N_1624);
and U2249 (N_2249,N_1657,N_1905);
nand U2250 (N_2250,N_1841,N_1901);
or U2251 (N_2251,N_1756,N_1737);
nor U2252 (N_2252,N_1673,N_1507);
and U2253 (N_2253,N_1922,N_1834);
nand U2254 (N_2254,N_1662,N_1650);
and U2255 (N_2255,N_1991,N_1555);
nand U2256 (N_2256,N_1715,N_1756);
and U2257 (N_2257,N_1543,N_1964);
nor U2258 (N_2258,N_1709,N_1542);
and U2259 (N_2259,N_1537,N_1828);
and U2260 (N_2260,N_1889,N_1786);
or U2261 (N_2261,N_1513,N_1989);
or U2262 (N_2262,N_1924,N_1848);
or U2263 (N_2263,N_1713,N_1963);
and U2264 (N_2264,N_1960,N_1639);
and U2265 (N_2265,N_1509,N_1876);
nand U2266 (N_2266,N_1921,N_1856);
nand U2267 (N_2267,N_1617,N_1724);
nand U2268 (N_2268,N_1891,N_1500);
or U2269 (N_2269,N_1739,N_1513);
nand U2270 (N_2270,N_1958,N_1968);
or U2271 (N_2271,N_1537,N_1974);
nand U2272 (N_2272,N_1907,N_1838);
and U2273 (N_2273,N_1503,N_1915);
and U2274 (N_2274,N_1961,N_1546);
or U2275 (N_2275,N_1900,N_1957);
and U2276 (N_2276,N_1963,N_1544);
xor U2277 (N_2277,N_1961,N_1812);
nor U2278 (N_2278,N_1923,N_1651);
and U2279 (N_2279,N_1873,N_1623);
or U2280 (N_2280,N_1519,N_1591);
nand U2281 (N_2281,N_1798,N_1985);
and U2282 (N_2282,N_1971,N_1918);
or U2283 (N_2283,N_1846,N_1883);
or U2284 (N_2284,N_1917,N_1959);
and U2285 (N_2285,N_1503,N_1510);
nor U2286 (N_2286,N_1624,N_1823);
and U2287 (N_2287,N_1599,N_1568);
nand U2288 (N_2288,N_1834,N_1782);
nand U2289 (N_2289,N_1941,N_1620);
nand U2290 (N_2290,N_1945,N_1808);
nand U2291 (N_2291,N_1799,N_1524);
nor U2292 (N_2292,N_1592,N_1722);
or U2293 (N_2293,N_1635,N_1656);
or U2294 (N_2294,N_1528,N_1555);
and U2295 (N_2295,N_1717,N_1548);
nand U2296 (N_2296,N_1921,N_1977);
and U2297 (N_2297,N_1806,N_1942);
or U2298 (N_2298,N_1934,N_1730);
nand U2299 (N_2299,N_1737,N_1890);
nor U2300 (N_2300,N_1771,N_1501);
and U2301 (N_2301,N_1538,N_1533);
nor U2302 (N_2302,N_1903,N_1716);
or U2303 (N_2303,N_1890,N_1981);
or U2304 (N_2304,N_1507,N_1634);
nand U2305 (N_2305,N_1974,N_1802);
nor U2306 (N_2306,N_1667,N_1986);
nand U2307 (N_2307,N_1577,N_1947);
nor U2308 (N_2308,N_1755,N_1587);
nand U2309 (N_2309,N_1767,N_1656);
nand U2310 (N_2310,N_1991,N_1679);
nand U2311 (N_2311,N_1882,N_1594);
or U2312 (N_2312,N_1525,N_1984);
and U2313 (N_2313,N_1654,N_1835);
nor U2314 (N_2314,N_1937,N_1948);
and U2315 (N_2315,N_1877,N_1702);
or U2316 (N_2316,N_1994,N_1756);
nor U2317 (N_2317,N_1849,N_1766);
nor U2318 (N_2318,N_1757,N_1559);
or U2319 (N_2319,N_1679,N_1837);
or U2320 (N_2320,N_1508,N_1812);
nor U2321 (N_2321,N_1539,N_1521);
nor U2322 (N_2322,N_1830,N_1889);
nor U2323 (N_2323,N_1834,N_1509);
nor U2324 (N_2324,N_1901,N_1902);
xnor U2325 (N_2325,N_1558,N_1929);
nand U2326 (N_2326,N_1861,N_1807);
and U2327 (N_2327,N_1583,N_1596);
or U2328 (N_2328,N_1814,N_1819);
nand U2329 (N_2329,N_1858,N_1684);
nand U2330 (N_2330,N_1780,N_1719);
nor U2331 (N_2331,N_1684,N_1876);
nor U2332 (N_2332,N_1819,N_1665);
nand U2333 (N_2333,N_1840,N_1992);
nand U2334 (N_2334,N_1938,N_1645);
or U2335 (N_2335,N_1526,N_1653);
or U2336 (N_2336,N_1608,N_1551);
and U2337 (N_2337,N_1533,N_1521);
or U2338 (N_2338,N_1849,N_1546);
nor U2339 (N_2339,N_1844,N_1864);
nor U2340 (N_2340,N_1958,N_1891);
nand U2341 (N_2341,N_1692,N_1539);
or U2342 (N_2342,N_1722,N_1550);
and U2343 (N_2343,N_1732,N_1964);
nor U2344 (N_2344,N_1975,N_1698);
nand U2345 (N_2345,N_1583,N_1502);
and U2346 (N_2346,N_1558,N_1620);
nor U2347 (N_2347,N_1596,N_1570);
or U2348 (N_2348,N_1866,N_1769);
and U2349 (N_2349,N_1825,N_1586);
nand U2350 (N_2350,N_1659,N_1741);
nand U2351 (N_2351,N_1691,N_1585);
nand U2352 (N_2352,N_1546,N_1734);
nand U2353 (N_2353,N_1745,N_1950);
xor U2354 (N_2354,N_1705,N_1993);
or U2355 (N_2355,N_1884,N_1852);
nand U2356 (N_2356,N_1728,N_1972);
or U2357 (N_2357,N_1657,N_1743);
nand U2358 (N_2358,N_1740,N_1790);
nor U2359 (N_2359,N_1877,N_1663);
or U2360 (N_2360,N_1647,N_1962);
and U2361 (N_2361,N_1755,N_1736);
and U2362 (N_2362,N_1533,N_1562);
nand U2363 (N_2363,N_1731,N_1998);
nand U2364 (N_2364,N_1849,N_1929);
nand U2365 (N_2365,N_1955,N_1987);
and U2366 (N_2366,N_1798,N_1711);
and U2367 (N_2367,N_1793,N_1871);
and U2368 (N_2368,N_1963,N_1856);
nor U2369 (N_2369,N_1813,N_1696);
and U2370 (N_2370,N_1664,N_1803);
and U2371 (N_2371,N_1847,N_1934);
nand U2372 (N_2372,N_1879,N_1796);
nand U2373 (N_2373,N_1656,N_1519);
and U2374 (N_2374,N_1798,N_1539);
and U2375 (N_2375,N_1794,N_1935);
nand U2376 (N_2376,N_1589,N_1783);
nand U2377 (N_2377,N_1828,N_1827);
and U2378 (N_2378,N_1836,N_1640);
or U2379 (N_2379,N_1900,N_1787);
and U2380 (N_2380,N_1844,N_1578);
nand U2381 (N_2381,N_1924,N_1681);
nand U2382 (N_2382,N_1655,N_1542);
and U2383 (N_2383,N_1567,N_1755);
and U2384 (N_2384,N_1531,N_1829);
or U2385 (N_2385,N_1580,N_1990);
nor U2386 (N_2386,N_1846,N_1894);
or U2387 (N_2387,N_1905,N_1540);
and U2388 (N_2388,N_1835,N_1677);
nand U2389 (N_2389,N_1670,N_1560);
and U2390 (N_2390,N_1954,N_1910);
nor U2391 (N_2391,N_1992,N_1753);
nor U2392 (N_2392,N_1868,N_1723);
and U2393 (N_2393,N_1690,N_1842);
xor U2394 (N_2394,N_1548,N_1742);
nand U2395 (N_2395,N_1885,N_1635);
and U2396 (N_2396,N_1585,N_1870);
and U2397 (N_2397,N_1555,N_1972);
nor U2398 (N_2398,N_1686,N_1584);
or U2399 (N_2399,N_1558,N_1550);
and U2400 (N_2400,N_1634,N_1567);
and U2401 (N_2401,N_1949,N_1911);
nand U2402 (N_2402,N_1651,N_1994);
or U2403 (N_2403,N_1876,N_1505);
nor U2404 (N_2404,N_1776,N_1733);
nand U2405 (N_2405,N_1526,N_1650);
and U2406 (N_2406,N_1907,N_1774);
or U2407 (N_2407,N_1880,N_1999);
and U2408 (N_2408,N_1589,N_1850);
and U2409 (N_2409,N_1732,N_1999);
or U2410 (N_2410,N_1581,N_1897);
xor U2411 (N_2411,N_1945,N_1761);
xor U2412 (N_2412,N_1872,N_1825);
xor U2413 (N_2413,N_1774,N_1517);
or U2414 (N_2414,N_1884,N_1792);
nor U2415 (N_2415,N_1910,N_1782);
or U2416 (N_2416,N_1563,N_1912);
nand U2417 (N_2417,N_1695,N_1540);
nor U2418 (N_2418,N_1877,N_1562);
and U2419 (N_2419,N_1607,N_1509);
and U2420 (N_2420,N_1977,N_1643);
nand U2421 (N_2421,N_1844,N_1551);
or U2422 (N_2422,N_1986,N_1920);
or U2423 (N_2423,N_1653,N_1874);
and U2424 (N_2424,N_1741,N_1665);
or U2425 (N_2425,N_1764,N_1737);
nand U2426 (N_2426,N_1657,N_1855);
and U2427 (N_2427,N_1554,N_1922);
nand U2428 (N_2428,N_1829,N_1623);
nor U2429 (N_2429,N_1863,N_1873);
nand U2430 (N_2430,N_1849,N_1815);
nand U2431 (N_2431,N_1996,N_1711);
nand U2432 (N_2432,N_1822,N_1563);
nand U2433 (N_2433,N_1988,N_1524);
or U2434 (N_2434,N_1642,N_1823);
nor U2435 (N_2435,N_1962,N_1974);
nand U2436 (N_2436,N_1846,N_1805);
nand U2437 (N_2437,N_1854,N_1884);
and U2438 (N_2438,N_1722,N_1855);
nand U2439 (N_2439,N_1994,N_1809);
and U2440 (N_2440,N_1918,N_1579);
and U2441 (N_2441,N_1800,N_1520);
nor U2442 (N_2442,N_1647,N_1949);
and U2443 (N_2443,N_1544,N_1967);
or U2444 (N_2444,N_1940,N_1976);
and U2445 (N_2445,N_1766,N_1951);
and U2446 (N_2446,N_1911,N_1969);
or U2447 (N_2447,N_1874,N_1585);
nand U2448 (N_2448,N_1654,N_1852);
or U2449 (N_2449,N_1563,N_1559);
or U2450 (N_2450,N_1543,N_1775);
nor U2451 (N_2451,N_1513,N_1998);
nor U2452 (N_2452,N_1540,N_1518);
and U2453 (N_2453,N_1531,N_1538);
and U2454 (N_2454,N_1558,N_1529);
nand U2455 (N_2455,N_1835,N_1687);
nand U2456 (N_2456,N_1518,N_1516);
or U2457 (N_2457,N_1621,N_1679);
nor U2458 (N_2458,N_1807,N_1942);
nor U2459 (N_2459,N_1667,N_1734);
nand U2460 (N_2460,N_1835,N_1971);
and U2461 (N_2461,N_1727,N_1945);
and U2462 (N_2462,N_1670,N_1833);
nand U2463 (N_2463,N_1537,N_1939);
nor U2464 (N_2464,N_1940,N_1581);
or U2465 (N_2465,N_1881,N_1972);
and U2466 (N_2466,N_1858,N_1725);
nand U2467 (N_2467,N_1716,N_1938);
nor U2468 (N_2468,N_1990,N_1983);
nand U2469 (N_2469,N_1829,N_1530);
nor U2470 (N_2470,N_1555,N_1921);
nor U2471 (N_2471,N_1830,N_1713);
and U2472 (N_2472,N_1755,N_1680);
or U2473 (N_2473,N_1786,N_1564);
and U2474 (N_2474,N_1569,N_1802);
or U2475 (N_2475,N_1588,N_1763);
nor U2476 (N_2476,N_1546,N_1960);
nor U2477 (N_2477,N_1580,N_1979);
or U2478 (N_2478,N_1550,N_1922);
xnor U2479 (N_2479,N_1827,N_1798);
nand U2480 (N_2480,N_1728,N_1631);
or U2481 (N_2481,N_1505,N_1746);
nand U2482 (N_2482,N_1608,N_1783);
or U2483 (N_2483,N_1873,N_1554);
nor U2484 (N_2484,N_1530,N_1988);
xnor U2485 (N_2485,N_1858,N_1831);
nor U2486 (N_2486,N_1583,N_1660);
and U2487 (N_2487,N_1558,N_1955);
nor U2488 (N_2488,N_1716,N_1776);
nor U2489 (N_2489,N_1980,N_1940);
nand U2490 (N_2490,N_1777,N_1719);
and U2491 (N_2491,N_1938,N_1710);
nor U2492 (N_2492,N_1522,N_1688);
nor U2493 (N_2493,N_1515,N_1749);
nand U2494 (N_2494,N_1985,N_1570);
nor U2495 (N_2495,N_1790,N_1755);
nor U2496 (N_2496,N_1675,N_1909);
nand U2497 (N_2497,N_1551,N_1742);
nor U2498 (N_2498,N_1973,N_1833);
nand U2499 (N_2499,N_1905,N_1530);
nor U2500 (N_2500,N_2372,N_2075);
nor U2501 (N_2501,N_2485,N_2328);
nand U2502 (N_2502,N_2272,N_2217);
or U2503 (N_2503,N_2431,N_2071);
nand U2504 (N_2504,N_2214,N_2055);
nand U2505 (N_2505,N_2013,N_2203);
and U2506 (N_2506,N_2268,N_2245);
and U2507 (N_2507,N_2218,N_2024);
and U2508 (N_2508,N_2181,N_2137);
or U2509 (N_2509,N_2407,N_2248);
or U2510 (N_2510,N_2316,N_2096);
or U2511 (N_2511,N_2278,N_2048);
and U2512 (N_2512,N_2389,N_2116);
nor U2513 (N_2513,N_2348,N_2251);
or U2514 (N_2514,N_2145,N_2223);
nor U2515 (N_2515,N_2486,N_2000);
nor U2516 (N_2516,N_2001,N_2043);
and U2517 (N_2517,N_2022,N_2311);
nand U2518 (N_2518,N_2166,N_2383);
and U2519 (N_2519,N_2444,N_2056);
and U2520 (N_2520,N_2063,N_2113);
or U2521 (N_2521,N_2170,N_2498);
or U2522 (N_2522,N_2104,N_2072);
and U2523 (N_2523,N_2288,N_2090);
or U2524 (N_2524,N_2443,N_2495);
nor U2525 (N_2525,N_2310,N_2420);
or U2526 (N_2526,N_2171,N_2014);
nor U2527 (N_2527,N_2342,N_2338);
or U2528 (N_2528,N_2489,N_2294);
nor U2529 (N_2529,N_2415,N_2067);
nand U2530 (N_2530,N_2313,N_2239);
nand U2531 (N_2531,N_2180,N_2402);
nor U2532 (N_2532,N_2030,N_2280);
nand U2533 (N_2533,N_2483,N_2006);
xnor U2534 (N_2534,N_2073,N_2395);
and U2535 (N_2535,N_2032,N_2490);
nor U2536 (N_2536,N_2125,N_2035);
nor U2537 (N_2537,N_2345,N_2334);
or U2538 (N_2538,N_2253,N_2423);
or U2539 (N_2539,N_2270,N_2147);
nand U2540 (N_2540,N_2445,N_2153);
and U2541 (N_2541,N_2088,N_2461);
or U2542 (N_2542,N_2391,N_2428);
xnor U2543 (N_2543,N_2271,N_2205);
nor U2544 (N_2544,N_2267,N_2343);
and U2545 (N_2545,N_2244,N_2258);
and U2546 (N_2546,N_2156,N_2277);
nor U2547 (N_2547,N_2028,N_2482);
nor U2548 (N_2548,N_2186,N_2151);
or U2549 (N_2549,N_2276,N_2499);
nor U2550 (N_2550,N_2341,N_2478);
and U2551 (N_2551,N_2379,N_2121);
or U2552 (N_2552,N_2227,N_2152);
and U2553 (N_2553,N_2016,N_2064);
nand U2554 (N_2554,N_2111,N_2260);
nor U2555 (N_2555,N_2359,N_2307);
or U2556 (N_2556,N_2371,N_2015);
nand U2557 (N_2557,N_2034,N_2287);
nor U2558 (N_2558,N_2354,N_2209);
nand U2559 (N_2559,N_2254,N_2336);
nor U2560 (N_2560,N_2304,N_2143);
or U2561 (N_2561,N_2216,N_2179);
and U2562 (N_2562,N_2496,N_2408);
or U2563 (N_2563,N_2135,N_2264);
nand U2564 (N_2564,N_2285,N_2281);
or U2565 (N_2565,N_2448,N_2435);
nor U2566 (N_2566,N_2114,N_2213);
or U2567 (N_2567,N_2070,N_2293);
nor U2568 (N_2568,N_2099,N_2057);
nor U2569 (N_2569,N_2246,N_2106);
nor U2570 (N_2570,N_2173,N_2178);
nor U2571 (N_2571,N_2128,N_2273);
and U2572 (N_2572,N_2182,N_2002);
nor U2573 (N_2573,N_2394,N_2026);
nor U2574 (N_2574,N_2255,N_2038);
or U2575 (N_2575,N_2424,N_2319);
nor U2576 (N_2576,N_2092,N_2140);
or U2577 (N_2577,N_2101,N_2332);
nor U2578 (N_2578,N_2323,N_2052);
nand U2579 (N_2579,N_2089,N_2003);
nand U2580 (N_2580,N_2470,N_2301);
or U2581 (N_2581,N_2078,N_2119);
nor U2582 (N_2582,N_2466,N_2426);
or U2583 (N_2583,N_2331,N_2465);
nand U2584 (N_2584,N_2427,N_2105);
nor U2585 (N_2585,N_2210,N_2029);
nand U2586 (N_2586,N_2405,N_2400);
nor U2587 (N_2587,N_2358,N_2370);
nand U2588 (N_2588,N_2131,N_2403);
or U2589 (N_2589,N_2229,N_2017);
and U2590 (N_2590,N_2148,N_2100);
nor U2591 (N_2591,N_2086,N_2475);
and U2592 (N_2592,N_2350,N_2091);
nor U2593 (N_2593,N_2306,N_2107);
nand U2594 (N_2594,N_2161,N_2149);
xnor U2595 (N_2595,N_2237,N_2335);
nor U2596 (N_2596,N_2419,N_2068);
nand U2597 (N_2597,N_2291,N_2221);
nor U2598 (N_2598,N_2436,N_2007);
nand U2599 (N_2599,N_2375,N_2312);
nand U2600 (N_2600,N_2492,N_2409);
and U2601 (N_2601,N_2115,N_2451);
or U2602 (N_2602,N_2366,N_2487);
nor U2603 (N_2603,N_2228,N_2497);
or U2604 (N_2604,N_2290,N_2447);
nor U2605 (N_2605,N_2361,N_2346);
nor U2606 (N_2606,N_2042,N_2226);
and U2607 (N_2607,N_2187,N_2416);
nor U2608 (N_2608,N_2390,N_2110);
xnor U2609 (N_2609,N_2146,N_2077);
nand U2610 (N_2610,N_2165,N_2184);
or U2611 (N_2611,N_2356,N_2378);
nor U2612 (N_2612,N_2437,N_2202);
or U2613 (N_2613,N_2404,N_2455);
or U2614 (N_2614,N_2076,N_2102);
and U2615 (N_2615,N_2252,N_2103);
nand U2616 (N_2616,N_2176,N_2368);
and U2617 (N_2617,N_2011,N_2297);
nand U2618 (N_2618,N_2132,N_2094);
or U2619 (N_2619,N_2215,N_2357);
nor U2620 (N_2620,N_2450,N_2230);
and U2621 (N_2621,N_2292,N_2275);
and U2622 (N_2622,N_2120,N_2109);
and U2623 (N_2623,N_2446,N_2473);
and U2624 (N_2624,N_2397,N_2393);
nand U2625 (N_2625,N_2159,N_2386);
or U2626 (N_2626,N_2136,N_2241);
and U2627 (N_2627,N_2308,N_2185);
nand U2628 (N_2628,N_2355,N_2095);
or U2629 (N_2629,N_2429,N_2263);
nor U2630 (N_2630,N_2256,N_2249);
or U2631 (N_2631,N_2235,N_2004);
or U2632 (N_2632,N_2413,N_2054);
nand U2633 (N_2633,N_2265,N_2144);
nand U2634 (N_2634,N_2066,N_2162);
nor U2635 (N_2635,N_2192,N_2289);
and U2636 (N_2636,N_2044,N_2039);
xor U2637 (N_2637,N_2351,N_2330);
nand U2638 (N_2638,N_2023,N_2240);
nor U2639 (N_2639,N_2299,N_2009);
nand U2640 (N_2640,N_2484,N_2417);
and U2641 (N_2641,N_2238,N_2286);
and U2642 (N_2642,N_2480,N_2344);
or U2643 (N_2643,N_2033,N_2399);
nor U2644 (N_2644,N_2220,N_2041);
nor U2645 (N_2645,N_2141,N_2296);
and U2646 (N_2646,N_2191,N_2481);
nand U2647 (N_2647,N_2352,N_2138);
or U2648 (N_2648,N_2195,N_2479);
or U2649 (N_2649,N_2333,N_2112);
or U2650 (N_2650,N_2060,N_2385);
xnor U2651 (N_2651,N_2406,N_2468);
and U2652 (N_2652,N_2440,N_2488);
and U2653 (N_2653,N_2211,N_2469);
nand U2654 (N_2654,N_2084,N_2326);
nor U2655 (N_2655,N_2284,N_2021);
or U2656 (N_2656,N_2062,N_2061);
xnor U2657 (N_2657,N_2040,N_2083);
and U2658 (N_2658,N_2367,N_2183);
nor U2659 (N_2659,N_2027,N_2329);
nor U2660 (N_2660,N_2476,N_2369);
or U2661 (N_2661,N_2283,N_2020);
nor U2662 (N_2662,N_2374,N_2175);
and U2663 (N_2663,N_2158,N_2142);
or U2664 (N_2664,N_2108,N_2491);
and U2665 (N_2665,N_2373,N_2163);
or U2666 (N_2666,N_2080,N_2309);
nand U2667 (N_2667,N_2133,N_2477);
and U2668 (N_2668,N_2414,N_2462);
nor U2669 (N_2669,N_2177,N_2471);
or U2670 (N_2670,N_2189,N_2317);
or U2671 (N_2671,N_2155,N_2257);
nor U2672 (N_2672,N_2172,N_2045);
nand U2673 (N_2673,N_2222,N_2458);
and U2674 (N_2674,N_2339,N_2388);
or U2675 (N_2675,N_2314,N_2449);
or U2676 (N_2676,N_2347,N_2079);
nor U2677 (N_2677,N_2097,N_2303);
or U2678 (N_2678,N_2442,N_2438);
nor U2679 (N_2679,N_2204,N_2049);
or U2680 (N_2680,N_2164,N_2224);
or U2681 (N_2681,N_2434,N_2259);
nand U2682 (N_2682,N_2194,N_2047);
and U2683 (N_2683,N_2212,N_2200);
or U2684 (N_2684,N_2093,N_2122);
and U2685 (N_2685,N_2327,N_2453);
nor U2686 (N_2686,N_2082,N_2460);
nand U2687 (N_2687,N_2134,N_2322);
and U2688 (N_2688,N_2325,N_2117);
nor U2689 (N_2689,N_2190,N_2493);
nor U2690 (N_2690,N_2425,N_2364);
or U2691 (N_2691,N_2167,N_2382);
nor U2692 (N_2692,N_2236,N_2349);
nand U2693 (N_2693,N_2242,N_2454);
and U2694 (N_2694,N_2452,N_2433);
nor U2695 (N_2695,N_2412,N_2457);
or U2696 (N_2696,N_2376,N_2472);
nor U2697 (N_2697,N_2365,N_2225);
or U2698 (N_2698,N_2233,N_2127);
nor U2699 (N_2699,N_2360,N_2059);
or U2700 (N_2700,N_2363,N_2421);
nand U2701 (N_2701,N_2168,N_2069);
nand U2702 (N_2702,N_2459,N_2302);
nand U2703 (N_2703,N_2154,N_2282);
and U2704 (N_2704,N_2199,N_2439);
nand U2705 (N_2705,N_2208,N_2305);
and U2706 (N_2706,N_2123,N_2234);
nor U2707 (N_2707,N_2193,N_2337);
nand U2708 (N_2708,N_2196,N_2410);
nand U2709 (N_2709,N_2474,N_2019);
nor U2710 (N_2710,N_2315,N_2387);
and U2711 (N_2711,N_2025,N_2261);
or U2712 (N_2712,N_2380,N_2169);
nor U2713 (N_2713,N_2081,N_2422);
and U2714 (N_2714,N_2464,N_2430);
nand U2715 (N_2715,N_2298,N_2467);
and U2716 (N_2716,N_2219,N_2139);
or U2717 (N_2717,N_2494,N_2362);
and U2718 (N_2718,N_2037,N_2441);
or U2719 (N_2719,N_2074,N_2005);
nor U2720 (N_2720,N_2058,N_2274);
nor U2721 (N_2721,N_2247,N_2124);
nand U2722 (N_2722,N_2384,N_2432);
nor U2723 (N_2723,N_2065,N_2324);
and U2724 (N_2724,N_2377,N_2150);
nand U2725 (N_2725,N_2262,N_2085);
or U2726 (N_2726,N_2411,N_2051);
nor U2727 (N_2727,N_2295,N_2197);
and U2728 (N_2728,N_2207,N_2050);
nand U2729 (N_2729,N_2053,N_2418);
nand U2730 (N_2730,N_2243,N_2036);
nand U2731 (N_2731,N_2126,N_2456);
nor U2732 (N_2732,N_2318,N_2269);
or U2733 (N_2733,N_2174,N_2279);
or U2734 (N_2734,N_2398,N_2130);
nand U2735 (N_2735,N_2012,N_2353);
xnor U2736 (N_2736,N_2010,N_2046);
and U2737 (N_2737,N_2381,N_2392);
nand U2738 (N_2738,N_2300,N_2463);
and U2739 (N_2739,N_2098,N_2401);
or U2740 (N_2740,N_2198,N_2206);
nor U2741 (N_2741,N_2018,N_2087);
or U2742 (N_2742,N_2320,N_2008);
or U2743 (N_2743,N_2160,N_2231);
or U2744 (N_2744,N_2201,N_2266);
or U2745 (N_2745,N_2340,N_2188);
and U2746 (N_2746,N_2118,N_2031);
nand U2747 (N_2747,N_2396,N_2157);
nor U2748 (N_2748,N_2250,N_2129);
or U2749 (N_2749,N_2232,N_2321);
or U2750 (N_2750,N_2075,N_2325);
nor U2751 (N_2751,N_2486,N_2027);
and U2752 (N_2752,N_2420,N_2381);
nor U2753 (N_2753,N_2294,N_2472);
and U2754 (N_2754,N_2053,N_2323);
nand U2755 (N_2755,N_2122,N_2092);
or U2756 (N_2756,N_2332,N_2341);
or U2757 (N_2757,N_2270,N_2288);
and U2758 (N_2758,N_2204,N_2466);
and U2759 (N_2759,N_2422,N_2187);
or U2760 (N_2760,N_2454,N_2047);
and U2761 (N_2761,N_2025,N_2368);
or U2762 (N_2762,N_2093,N_2336);
nor U2763 (N_2763,N_2071,N_2112);
nor U2764 (N_2764,N_2463,N_2183);
or U2765 (N_2765,N_2251,N_2376);
or U2766 (N_2766,N_2167,N_2384);
and U2767 (N_2767,N_2299,N_2355);
xor U2768 (N_2768,N_2198,N_2015);
nor U2769 (N_2769,N_2040,N_2124);
nor U2770 (N_2770,N_2303,N_2050);
and U2771 (N_2771,N_2150,N_2127);
nand U2772 (N_2772,N_2223,N_2072);
and U2773 (N_2773,N_2457,N_2091);
nand U2774 (N_2774,N_2085,N_2252);
and U2775 (N_2775,N_2121,N_2206);
and U2776 (N_2776,N_2425,N_2376);
and U2777 (N_2777,N_2174,N_2101);
and U2778 (N_2778,N_2133,N_2104);
nor U2779 (N_2779,N_2022,N_2064);
and U2780 (N_2780,N_2408,N_2019);
or U2781 (N_2781,N_2437,N_2482);
nor U2782 (N_2782,N_2192,N_2355);
nand U2783 (N_2783,N_2368,N_2306);
nand U2784 (N_2784,N_2146,N_2024);
nor U2785 (N_2785,N_2489,N_2055);
and U2786 (N_2786,N_2274,N_2389);
or U2787 (N_2787,N_2428,N_2085);
nor U2788 (N_2788,N_2224,N_2209);
and U2789 (N_2789,N_2308,N_2186);
and U2790 (N_2790,N_2232,N_2420);
nand U2791 (N_2791,N_2379,N_2155);
and U2792 (N_2792,N_2176,N_2393);
xor U2793 (N_2793,N_2204,N_2157);
or U2794 (N_2794,N_2410,N_2018);
nand U2795 (N_2795,N_2474,N_2000);
nand U2796 (N_2796,N_2072,N_2364);
or U2797 (N_2797,N_2151,N_2181);
nor U2798 (N_2798,N_2278,N_2300);
nor U2799 (N_2799,N_2394,N_2073);
nor U2800 (N_2800,N_2205,N_2457);
xor U2801 (N_2801,N_2059,N_2331);
nor U2802 (N_2802,N_2013,N_2223);
nand U2803 (N_2803,N_2191,N_2210);
xnor U2804 (N_2804,N_2167,N_2163);
or U2805 (N_2805,N_2078,N_2215);
and U2806 (N_2806,N_2278,N_2074);
or U2807 (N_2807,N_2058,N_2353);
or U2808 (N_2808,N_2445,N_2227);
nor U2809 (N_2809,N_2475,N_2203);
nand U2810 (N_2810,N_2089,N_2051);
nor U2811 (N_2811,N_2234,N_2314);
xnor U2812 (N_2812,N_2442,N_2223);
and U2813 (N_2813,N_2317,N_2214);
and U2814 (N_2814,N_2438,N_2497);
nor U2815 (N_2815,N_2230,N_2177);
nand U2816 (N_2816,N_2289,N_2336);
xor U2817 (N_2817,N_2381,N_2449);
nand U2818 (N_2818,N_2129,N_2290);
or U2819 (N_2819,N_2323,N_2120);
or U2820 (N_2820,N_2084,N_2201);
nand U2821 (N_2821,N_2297,N_2226);
nor U2822 (N_2822,N_2080,N_2041);
nand U2823 (N_2823,N_2444,N_2113);
nor U2824 (N_2824,N_2418,N_2471);
and U2825 (N_2825,N_2319,N_2041);
or U2826 (N_2826,N_2444,N_2244);
nand U2827 (N_2827,N_2123,N_2131);
xor U2828 (N_2828,N_2322,N_2443);
nand U2829 (N_2829,N_2353,N_2146);
nor U2830 (N_2830,N_2187,N_2239);
nor U2831 (N_2831,N_2046,N_2409);
nand U2832 (N_2832,N_2343,N_2245);
or U2833 (N_2833,N_2439,N_2015);
nand U2834 (N_2834,N_2342,N_2208);
nor U2835 (N_2835,N_2465,N_2429);
nor U2836 (N_2836,N_2475,N_2054);
nand U2837 (N_2837,N_2219,N_2400);
nand U2838 (N_2838,N_2170,N_2475);
xor U2839 (N_2839,N_2404,N_2320);
and U2840 (N_2840,N_2332,N_2465);
nor U2841 (N_2841,N_2463,N_2430);
and U2842 (N_2842,N_2452,N_2090);
or U2843 (N_2843,N_2257,N_2110);
nand U2844 (N_2844,N_2260,N_2296);
nand U2845 (N_2845,N_2175,N_2065);
nand U2846 (N_2846,N_2196,N_2147);
and U2847 (N_2847,N_2311,N_2240);
or U2848 (N_2848,N_2088,N_2499);
nand U2849 (N_2849,N_2369,N_2089);
nor U2850 (N_2850,N_2018,N_2270);
or U2851 (N_2851,N_2139,N_2328);
nor U2852 (N_2852,N_2025,N_2373);
nor U2853 (N_2853,N_2152,N_2284);
nand U2854 (N_2854,N_2428,N_2002);
nor U2855 (N_2855,N_2439,N_2413);
or U2856 (N_2856,N_2136,N_2015);
nand U2857 (N_2857,N_2268,N_2140);
nand U2858 (N_2858,N_2369,N_2073);
or U2859 (N_2859,N_2423,N_2421);
nand U2860 (N_2860,N_2456,N_2420);
nor U2861 (N_2861,N_2358,N_2101);
and U2862 (N_2862,N_2244,N_2314);
nand U2863 (N_2863,N_2028,N_2147);
nand U2864 (N_2864,N_2081,N_2233);
nor U2865 (N_2865,N_2240,N_2356);
and U2866 (N_2866,N_2459,N_2140);
or U2867 (N_2867,N_2159,N_2147);
and U2868 (N_2868,N_2103,N_2053);
nand U2869 (N_2869,N_2103,N_2401);
nor U2870 (N_2870,N_2245,N_2215);
nor U2871 (N_2871,N_2200,N_2290);
nor U2872 (N_2872,N_2220,N_2065);
nand U2873 (N_2873,N_2100,N_2326);
nand U2874 (N_2874,N_2406,N_2307);
nand U2875 (N_2875,N_2032,N_2402);
xor U2876 (N_2876,N_2307,N_2194);
nor U2877 (N_2877,N_2404,N_2247);
and U2878 (N_2878,N_2338,N_2335);
nand U2879 (N_2879,N_2109,N_2176);
nor U2880 (N_2880,N_2123,N_2414);
or U2881 (N_2881,N_2049,N_2284);
or U2882 (N_2882,N_2440,N_2104);
and U2883 (N_2883,N_2264,N_2145);
and U2884 (N_2884,N_2058,N_2037);
and U2885 (N_2885,N_2458,N_2109);
nor U2886 (N_2886,N_2314,N_2387);
nand U2887 (N_2887,N_2291,N_2420);
nand U2888 (N_2888,N_2113,N_2319);
or U2889 (N_2889,N_2029,N_2253);
nand U2890 (N_2890,N_2104,N_2139);
or U2891 (N_2891,N_2142,N_2260);
nor U2892 (N_2892,N_2090,N_2274);
or U2893 (N_2893,N_2260,N_2353);
and U2894 (N_2894,N_2065,N_2083);
and U2895 (N_2895,N_2234,N_2316);
nand U2896 (N_2896,N_2079,N_2055);
and U2897 (N_2897,N_2271,N_2265);
nand U2898 (N_2898,N_2222,N_2133);
nand U2899 (N_2899,N_2465,N_2079);
nand U2900 (N_2900,N_2258,N_2059);
nand U2901 (N_2901,N_2380,N_2339);
nand U2902 (N_2902,N_2424,N_2348);
nand U2903 (N_2903,N_2116,N_2101);
and U2904 (N_2904,N_2045,N_2454);
nand U2905 (N_2905,N_2034,N_2385);
nor U2906 (N_2906,N_2015,N_2479);
and U2907 (N_2907,N_2462,N_2237);
nor U2908 (N_2908,N_2280,N_2020);
nor U2909 (N_2909,N_2085,N_2187);
or U2910 (N_2910,N_2248,N_2191);
and U2911 (N_2911,N_2203,N_2041);
nand U2912 (N_2912,N_2157,N_2158);
or U2913 (N_2913,N_2116,N_2028);
nor U2914 (N_2914,N_2001,N_2373);
and U2915 (N_2915,N_2010,N_2181);
nor U2916 (N_2916,N_2412,N_2031);
and U2917 (N_2917,N_2298,N_2023);
or U2918 (N_2918,N_2088,N_2212);
nor U2919 (N_2919,N_2395,N_2043);
and U2920 (N_2920,N_2095,N_2279);
nand U2921 (N_2921,N_2430,N_2482);
nor U2922 (N_2922,N_2364,N_2478);
nor U2923 (N_2923,N_2175,N_2023);
nor U2924 (N_2924,N_2325,N_2010);
nor U2925 (N_2925,N_2121,N_2185);
or U2926 (N_2926,N_2403,N_2448);
nor U2927 (N_2927,N_2308,N_2024);
nor U2928 (N_2928,N_2146,N_2478);
xor U2929 (N_2929,N_2089,N_2230);
or U2930 (N_2930,N_2369,N_2222);
or U2931 (N_2931,N_2179,N_2493);
nor U2932 (N_2932,N_2465,N_2483);
nor U2933 (N_2933,N_2457,N_2446);
nand U2934 (N_2934,N_2425,N_2164);
nand U2935 (N_2935,N_2138,N_2198);
nand U2936 (N_2936,N_2358,N_2490);
and U2937 (N_2937,N_2051,N_2277);
and U2938 (N_2938,N_2357,N_2420);
or U2939 (N_2939,N_2315,N_2392);
and U2940 (N_2940,N_2432,N_2393);
or U2941 (N_2941,N_2142,N_2406);
and U2942 (N_2942,N_2483,N_2215);
nand U2943 (N_2943,N_2310,N_2374);
nand U2944 (N_2944,N_2307,N_2371);
xnor U2945 (N_2945,N_2401,N_2231);
and U2946 (N_2946,N_2483,N_2222);
nor U2947 (N_2947,N_2003,N_2461);
nor U2948 (N_2948,N_2342,N_2212);
nand U2949 (N_2949,N_2358,N_2218);
nand U2950 (N_2950,N_2293,N_2104);
nor U2951 (N_2951,N_2278,N_2149);
nor U2952 (N_2952,N_2336,N_2012);
nor U2953 (N_2953,N_2174,N_2063);
and U2954 (N_2954,N_2147,N_2237);
or U2955 (N_2955,N_2159,N_2266);
nand U2956 (N_2956,N_2238,N_2133);
or U2957 (N_2957,N_2491,N_2326);
and U2958 (N_2958,N_2418,N_2092);
nand U2959 (N_2959,N_2125,N_2462);
nor U2960 (N_2960,N_2338,N_2350);
and U2961 (N_2961,N_2260,N_2420);
and U2962 (N_2962,N_2221,N_2210);
or U2963 (N_2963,N_2111,N_2272);
nand U2964 (N_2964,N_2314,N_2062);
and U2965 (N_2965,N_2480,N_2161);
nand U2966 (N_2966,N_2028,N_2361);
and U2967 (N_2967,N_2361,N_2282);
nor U2968 (N_2968,N_2243,N_2120);
nor U2969 (N_2969,N_2281,N_2380);
nor U2970 (N_2970,N_2129,N_2379);
nor U2971 (N_2971,N_2209,N_2446);
nand U2972 (N_2972,N_2424,N_2024);
and U2973 (N_2973,N_2010,N_2411);
nor U2974 (N_2974,N_2255,N_2284);
and U2975 (N_2975,N_2080,N_2066);
or U2976 (N_2976,N_2392,N_2325);
nor U2977 (N_2977,N_2026,N_2171);
nand U2978 (N_2978,N_2422,N_2086);
or U2979 (N_2979,N_2288,N_2075);
or U2980 (N_2980,N_2128,N_2144);
and U2981 (N_2981,N_2138,N_2251);
nand U2982 (N_2982,N_2098,N_2329);
or U2983 (N_2983,N_2353,N_2381);
nor U2984 (N_2984,N_2490,N_2408);
xnor U2985 (N_2985,N_2215,N_2042);
nand U2986 (N_2986,N_2493,N_2199);
nor U2987 (N_2987,N_2031,N_2467);
nand U2988 (N_2988,N_2138,N_2378);
or U2989 (N_2989,N_2149,N_2383);
nand U2990 (N_2990,N_2121,N_2442);
and U2991 (N_2991,N_2020,N_2354);
xor U2992 (N_2992,N_2096,N_2235);
nand U2993 (N_2993,N_2463,N_2399);
or U2994 (N_2994,N_2097,N_2437);
nor U2995 (N_2995,N_2105,N_2211);
nor U2996 (N_2996,N_2185,N_2123);
or U2997 (N_2997,N_2282,N_2374);
or U2998 (N_2998,N_2311,N_2342);
nor U2999 (N_2999,N_2239,N_2275);
nor U3000 (N_3000,N_2919,N_2626);
nand U3001 (N_3001,N_2955,N_2789);
nand U3002 (N_3002,N_2971,N_2945);
or U3003 (N_3003,N_2908,N_2530);
nand U3004 (N_3004,N_2763,N_2977);
or U3005 (N_3005,N_2627,N_2931);
nor U3006 (N_3006,N_2628,N_2927);
nand U3007 (N_3007,N_2906,N_2715);
and U3008 (N_3008,N_2539,N_2837);
nand U3009 (N_3009,N_2509,N_2683);
and U3010 (N_3010,N_2845,N_2810);
and U3011 (N_3011,N_2982,N_2925);
or U3012 (N_3012,N_2872,N_2847);
or U3013 (N_3013,N_2795,N_2663);
nor U3014 (N_3014,N_2973,N_2885);
nor U3015 (N_3015,N_2727,N_2644);
nor U3016 (N_3016,N_2732,N_2710);
or U3017 (N_3017,N_2929,N_2711);
and U3018 (N_3018,N_2829,N_2529);
or U3019 (N_3019,N_2999,N_2900);
nor U3020 (N_3020,N_2704,N_2609);
xnor U3021 (N_3021,N_2915,N_2522);
nand U3022 (N_3022,N_2934,N_2868);
nand U3023 (N_3023,N_2717,N_2714);
nand U3024 (N_3024,N_2857,N_2508);
and U3025 (N_3025,N_2511,N_2596);
and U3026 (N_3026,N_2698,N_2702);
nor U3027 (N_3027,N_2685,N_2691);
nor U3028 (N_3028,N_2897,N_2779);
nand U3029 (N_3029,N_2749,N_2618);
nor U3030 (N_3030,N_2712,N_2788);
or U3031 (N_3031,N_2593,N_2639);
nand U3032 (N_3032,N_2625,N_2733);
nor U3033 (N_3033,N_2883,N_2921);
nor U3034 (N_3034,N_2928,N_2963);
nor U3035 (N_3035,N_2791,N_2518);
or U3036 (N_3036,N_2540,N_2670);
nor U3037 (N_3037,N_2780,N_2607);
or U3038 (N_3038,N_2998,N_2585);
and U3039 (N_3039,N_2541,N_2592);
nor U3040 (N_3040,N_2806,N_2597);
nor U3041 (N_3041,N_2759,N_2603);
nand U3042 (N_3042,N_2838,N_2990);
nor U3043 (N_3043,N_2828,N_2787);
nand U3044 (N_3044,N_2694,N_2831);
nor U3045 (N_3045,N_2561,N_2695);
nand U3046 (N_3046,N_2622,N_2944);
nor U3047 (N_3047,N_2756,N_2681);
nand U3048 (N_3048,N_2563,N_2504);
nor U3049 (N_3049,N_2718,N_2745);
and U3050 (N_3050,N_2692,N_2634);
nand U3051 (N_3051,N_2550,N_2635);
nand U3052 (N_3052,N_2677,N_2825);
nor U3053 (N_3053,N_2768,N_2578);
nand U3054 (N_3054,N_2972,N_2551);
nand U3055 (N_3055,N_2909,N_2661);
and U3056 (N_3056,N_2818,N_2599);
and U3057 (N_3057,N_2700,N_2752);
and U3058 (N_3058,N_2743,N_2730);
nor U3059 (N_3059,N_2836,N_2564);
nand U3060 (N_3060,N_2967,N_2546);
nor U3061 (N_3061,N_2907,N_2974);
nand U3062 (N_3062,N_2520,N_2744);
nand U3063 (N_3063,N_2542,N_2797);
or U3064 (N_3064,N_2862,N_2796);
and U3065 (N_3065,N_2848,N_2753);
nor U3066 (N_3066,N_2764,N_2722);
nor U3067 (N_3067,N_2668,N_2519);
and U3068 (N_3068,N_2874,N_2591);
or U3069 (N_3069,N_2948,N_2980);
nor U3070 (N_3070,N_2782,N_2901);
or U3071 (N_3071,N_2547,N_2935);
nand U3072 (N_3072,N_2992,N_2920);
nand U3073 (N_3073,N_2893,N_2871);
and U3074 (N_3074,N_2926,N_2606);
or U3075 (N_3075,N_2849,N_2569);
and U3076 (N_3076,N_2673,N_2951);
or U3077 (N_3077,N_2770,N_2760);
nor U3078 (N_3078,N_2884,N_2505);
and U3079 (N_3079,N_2570,N_2751);
nand U3080 (N_3080,N_2738,N_2619);
or U3081 (N_3081,N_2549,N_2721);
nor U3082 (N_3082,N_2731,N_2521);
nor U3083 (N_3083,N_2720,N_2545);
nor U3084 (N_3084,N_2556,N_2911);
xnor U3085 (N_3085,N_2559,N_2608);
nor U3086 (N_3086,N_2664,N_2724);
nor U3087 (N_3087,N_2543,N_2807);
or U3088 (N_3088,N_2696,N_2723);
and U3089 (N_3089,N_2769,N_2572);
and U3090 (N_3090,N_2669,N_2794);
or U3091 (N_3091,N_2595,N_2555);
and U3092 (N_3092,N_2594,N_2962);
nor U3093 (N_3093,N_2693,N_2953);
nor U3094 (N_3094,N_2558,N_2514);
or U3095 (N_3095,N_2958,N_2898);
and U3096 (N_3096,N_2641,N_2947);
and U3097 (N_3097,N_2923,N_2758);
and U3098 (N_3098,N_2856,N_2537);
nand U3099 (N_3099,N_2707,N_2647);
nand U3100 (N_3100,N_2579,N_2701);
nand U3101 (N_3101,N_2950,N_2834);
and U3102 (N_3102,N_2590,N_2983);
and U3103 (N_3103,N_2879,N_2894);
nand U3104 (N_3104,N_2560,N_2824);
or U3105 (N_3105,N_2614,N_2799);
nor U3106 (N_3106,N_2772,N_2880);
and U3107 (N_3107,N_2716,N_2943);
nor U3108 (N_3108,N_2895,N_2860);
and U3109 (N_3109,N_2913,N_2899);
or U3110 (N_3110,N_2778,N_2742);
or U3111 (N_3111,N_2703,N_2665);
nor U3112 (N_3112,N_2598,N_2930);
xor U3113 (N_3113,N_2655,N_2575);
nand U3114 (N_3114,N_2811,N_2666);
or U3115 (N_3115,N_2725,N_2652);
nand U3116 (N_3116,N_2699,N_2851);
nand U3117 (N_3117,N_2686,N_2936);
nor U3118 (N_3118,N_2844,N_2993);
and U3119 (N_3119,N_2544,N_2822);
nor U3120 (N_3120,N_2823,N_2922);
nand U3121 (N_3121,N_2531,N_2896);
nor U3122 (N_3122,N_2910,N_2678);
or U3123 (N_3123,N_2617,N_2873);
nor U3124 (N_3124,N_2775,N_2932);
or U3125 (N_3125,N_2638,N_2587);
nor U3126 (N_3126,N_2538,N_2832);
nor U3127 (N_3127,N_2937,N_2916);
or U3128 (N_3128,N_2820,N_2602);
xor U3129 (N_3129,N_2869,N_2584);
nor U3130 (N_3130,N_2528,N_2513);
or U3131 (N_3131,N_2675,N_2502);
or U3132 (N_3132,N_2623,N_2552);
and U3133 (N_3133,N_2600,N_2781);
or U3134 (N_3134,N_2777,N_2876);
nand U3135 (N_3135,N_2839,N_2589);
nand U3136 (N_3136,N_2580,N_2881);
nand U3137 (N_3137,N_2631,N_2814);
and U3138 (N_3138,N_2819,N_2525);
nor U3139 (N_3139,N_2888,N_2846);
nor U3140 (N_3140,N_2988,N_2583);
or U3141 (N_3141,N_2952,N_2985);
and U3142 (N_3142,N_2870,N_2997);
and U3143 (N_3143,N_2757,N_2688);
xnor U3144 (N_3144,N_2940,N_2658);
nand U3145 (N_3145,N_2765,N_2882);
or U3146 (N_3146,N_2903,N_2979);
or U3147 (N_3147,N_2803,N_2802);
nor U3148 (N_3148,N_2970,N_2527);
nand U3149 (N_3149,N_2503,N_2941);
nand U3150 (N_3150,N_2956,N_2776);
and U3151 (N_3151,N_2960,N_2728);
nand U3152 (N_3152,N_2612,N_2833);
or U3153 (N_3153,N_2610,N_2630);
nand U3154 (N_3154,N_2633,N_2792);
nand U3155 (N_3155,N_2645,N_2976);
or U3156 (N_3156,N_2949,N_2548);
or U3157 (N_3157,N_2755,N_2805);
nor U3158 (N_3158,N_2994,N_2889);
and U3159 (N_3159,N_2984,N_2709);
xor U3160 (N_3160,N_2968,N_2905);
and U3161 (N_3161,N_2861,N_2969);
and U3162 (N_3162,N_2774,N_2642);
and U3163 (N_3163,N_2676,N_2636);
and U3164 (N_3164,N_2705,N_2646);
nor U3165 (N_3165,N_2987,N_2662);
and U3166 (N_3166,N_2942,N_2887);
nor U3167 (N_3167,N_2826,N_2761);
nor U3168 (N_3168,N_2643,N_2510);
and U3169 (N_3169,N_2729,N_2816);
nor U3170 (N_3170,N_2914,N_2996);
nand U3171 (N_3171,N_2800,N_2516);
and U3172 (N_3172,N_2843,N_2739);
nor U3173 (N_3173,N_2878,N_2620);
or U3174 (N_3174,N_2746,N_2517);
or U3175 (N_3175,N_2801,N_2954);
nand U3176 (N_3176,N_2524,N_2902);
or U3177 (N_3177,N_2534,N_2588);
nand U3178 (N_3178,N_2991,N_2850);
nor U3179 (N_3179,N_2790,N_2854);
or U3180 (N_3180,N_2708,N_2650);
nor U3181 (N_3181,N_2853,N_2866);
and U3182 (N_3182,N_2891,N_2917);
and U3183 (N_3183,N_2875,N_2656);
nor U3184 (N_3184,N_2637,N_2684);
or U3185 (N_3185,N_2865,N_2817);
nor U3186 (N_3186,N_2601,N_2535);
nand U3187 (N_3187,N_2975,N_2690);
nand U3188 (N_3188,N_2737,N_2536);
or U3189 (N_3189,N_2667,N_2680);
nand U3190 (N_3190,N_2697,N_2939);
or U3191 (N_3191,N_2892,N_2827);
and U3192 (N_3192,N_2815,N_2835);
and U3193 (N_3193,N_2640,N_2786);
or U3194 (N_3194,N_2809,N_2852);
and U3195 (N_3195,N_2605,N_2812);
xnor U3196 (N_3196,N_2784,N_2582);
xnor U3197 (N_3197,N_2798,N_2762);
nand U3198 (N_3198,N_2793,N_2735);
nor U3199 (N_3199,N_2651,N_2783);
nor U3200 (N_3200,N_2632,N_2553);
and U3201 (N_3201,N_2989,N_2659);
nand U3202 (N_3202,N_2500,N_2629);
and U3203 (N_3203,N_2741,N_2532);
and U3204 (N_3204,N_2736,N_2959);
and U3205 (N_3205,N_2964,N_2523);
nor U3206 (N_3206,N_2566,N_2842);
or U3207 (N_3207,N_2574,N_2719);
and U3208 (N_3208,N_2571,N_2841);
or U3209 (N_3209,N_2740,N_2557);
nand U3210 (N_3210,N_2624,N_2526);
and U3211 (N_3211,N_2565,N_2660);
nand U3212 (N_3212,N_2813,N_2877);
nor U3213 (N_3213,N_2918,N_2785);
nand U3214 (N_3214,N_2747,N_2771);
nand U3215 (N_3215,N_2734,N_2904);
and U3216 (N_3216,N_2515,N_2657);
or U3217 (N_3217,N_2890,N_2981);
nand U3218 (N_3218,N_2754,N_2611);
and U3219 (N_3219,N_2912,N_2682);
nand U3220 (N_3220,N_2773,N_2726);
and U3221 (N_3221,N_2830,N_2648);
and U3222 (N_3222,N_2512,N_2750);
nand U3223 (N_3223,N_2507,N_2859);
nor U3224 (N_3224,N_2978,N_2581);
nand U3225 (N_3225,N_2604,N_2674);
nor U3226 (N_3226,N_2562,N_2804);
xor U3227 (N_3227,N_2748,N_2966);
and U3228 (N_3228,N_2689,N_2621);
nor U3229 (N_3229,N_2946,N_2766);
nor U3230 (N_3230,N_2924,N_2938);
and U3231 (N_3231,N_2616,N_2864);
or U3232 (N_3232,N_2863,N_2533);
and U3233 (N_3233,N_2821,N_2706);
nor U3234 (N_3234,N_2577,N_2568);
and U3235 (N_3235,N_2986,N_2679);
nor U3236 (N_3236,N_2654,N_2713);
nor U3237 (N_3237,N_2767,N_2867);
or U3238 (N_3238,N_2573,N_2886);
and U3239 (N_3239,N_2961,N_2808);
nor U3240 (N_3240,N_2554,N_2586);
nor U3241 (N_3241,N_2501,N_2858);
and U3242 (N_3242,N_2957,N_2995);
or U3243 (N_3243,N_2687,N_2576);
nor U3244 (N_3244,N_2671,N_2672);
nor U3245 (N_3245,N_2506,N_2855);
and U3246 (N_3246,N_2965,N_2567);
nand U3247 (N_3247,N_2933,N_2653);
nor U3248 (N_3248,N_2649,N_2615);
or U3249 (N_3249,N_2840,N_2613);
xnor U3250 (N_3250,N_2695,N_2980);
nand U3251 (N_3251,N_2500,N_2786);
and U3252 (N_3252,N_2629,N_2848);
nand U3253 (N_3253,N_2696,N_2643);
or U3254 (N_3254,N_2903,N_2845);
or U3255 (N_3255,N_2755,N_2525);
nand U3256 (N_3256,N_2652,N_2981);
nand U3257 (N_3257,N_2666,N_2984);
or U3258 (N_3258,N_2644,N_2764);
and U3259 (N_3259,N_2625,N_2756);
and U3260 (N_3260,N_2816,N_2872);
and U3261 (N_3261,N_2724,N_2828);
nor U3262 (N_3262,N_2733,N_2683);
and U3263 (N_3263,N_2680,N_2584);
nor U3264 (N_3264,N_2761,N_2737);
nand U3265 (N_3265,N_2999,N_2661);
nor U3266 (N_3266,N_2616,N_2723);
xor U3267 (N_3267,N_2901,N_2807);
or U3268 (N_3268,N_2725,N_2870);
and U3269 (N_3269,N_2761,N_2937);
nand U3270 (N_3270,N_2631,N_2605);
nor U3271 (N_3271,N_2955,N_2903);
or U3272 (N_3272,N_2579,N_2953);
nor U3273 (N_3273,N_2878,N_2831);
nand U3274 (N_3274,N_2707,N_2679);
nor U3275 (N_3275,N_2956,N_2542);
nand U3276 (N_3276,N_2700,N_2909);
nor U3277 (N_3277,N_2839,N_2643);
or U3278 (N_3278,N_2752,N_2568);
and U3279 (N_3279,N_2951,N_2646);
and U3280 (N_3280,N_2604,N_2875);
nand U3281 (N_3281,N_2837,N_2686);
or U3282 (N_3282,N_2928,N_2859);
and U3283 (N_3283,N_2810,N_2803);
or U3284 (N_3284,N_2870,N_2685);
and U3285 (N_3285,N_2838,N_2783);
and U3286 (N_3286,N_2892,N_2746);
or U3287 (N_3287,N_2734,N_2769);
nor U3288 (N_3288,N_2775,N_2525);
nor U3289 (N_3289,N_2523,N_2930);
or U3290 (N_3290,N_2775,N_2658);
and U3291 (N_3291,N_2611,N_2757);
or U3292 (N_3292,N_2893,N_2863);
nor U3293 (N_3293,N_2513,N_2512);
nor U3294 (N_3294,N_2898,N_2697);
or U3295 (N_3295,N_2511,N_2679);
xor U3296 (N_3296,N_2914,N_2711);
or U3297 (N_3297,N_2520,N_2779);
or U3298 (N_3298,N_2968,N_2860);
nand U3299 (N_3299,N_2539,N_2518);
or U3300 (N_3300,N_2923,N_2580);
nor U3301 (N_3301,N_2791,N_2676);
nand U3302 (N_3302,N_2787,N_2994);
or U3303 (N_3303,N_2624,N_2865);
nor U3304 (N_3304,N_2691,N_2877);
nand U3305 (N_3305,N_2949,N_2911);
nand U3306 (N_3306,N_2536,N_2841);
nand U3307 (N_3307,N_2657,N_2749);
and U3308 (N_3308,N_2937,N_2910);
and U3309 (N_3309,N_2591,N_2863);
or U3310 (N_3310,N_2720,N_2995);
nor U3311 (N_3311,N_2743,N_2780);
nor U3312 (N_3312,N_2571,N_2826);
and U3313 (N_3313,N_2946,N_2855);
nand U3314 (N_3314,N_2937,N_2930);
nand U3315 (N_3315,N_2573,N_2829);
nor U3316 (N_3316,N_2908,N_2755);
or U3317 (N_3317,N_2772,N_2528);
or U3318 (N_3318,N_2896,N_2952);
nor U3319 (N_3319,N_2851,N_2593);
nor U3320 (N_3320,N_2940,N_2636);
nor U3321 (N_3321,N_2707,N_2746);
nor U3322 (N_3322,N_2649,N_2527);
nor U3323 (N_3323,N_2546,N_2782);
and U3324 (N_3324,N_2570,N_2821);
or U3325 (N_3325,N_2782,N_2528);
nand U3326 (N_3326,N_2974,N_2680);
nor U3327 (N_3327,N_2632,N_2945);
nand U3328 (N_3328,N_2591,N_2597);
or U3329 (N_3329,N_2586,N_2831);
and U3330 (N_3330,N_2905,N_2607);
nand U3331 (N_3331,N_2921,N_2676);
nand U3332 (N_3332,N_2835,N_2603);
or U3333 (N_3333,N_2520,N_2831);
nor U3334 (N_3334,N_2783,N_2674);
xor U3335 (N_3335,N_2804,N_2805);
nor U3336 (N_3336,N_2807,N_2994);
or U3337 (N_3337,N_2631,N_2598);
nand U3338 (N_3338,N_2831,N_2826);
and U3339 (N_3339,N_2700,N_2957);
nand U3340 (N_3340,N_2731,N_2612);
nor U3341 (N_3341,N_2865,N_2600);
or U3342 (N_3342,N_2603,N_2971);
xor U3343 (N_3343,N_2953,N_2545);
nor U3344 (N_3344,N_2946,N_2717);
or U3345 (N_3345,N_2959,N_2753);
and U3346 (N_3346,N_2915,N_2832);
nor U3347 (N_3347,N_2984,N_2668);
nor U3348 (N_3348,N_2570,N_2609);
nand U3349 (N_3349,N_2705,N_2637);
nand U3350 (N_3350,N_2604,N_2769);
nand U3351 (N_3351,N_2967,N_2722);
nor U3352 (N_3352,N_2560,N_2657);
nand U3353 (N_3353,N_2857,N_2748);
nand U3354 (N_3354,N_2863,N_2852);
or U3355 (N_3355,N_2658,N_2509);
nand U3356 (N_3356,N_2698,N_2696);
nor U3357 (N_3357,N_2730,N_2734);
nor U3358 (N_3358,N_2533,N_2559);
and U3359 (N_3359,N_2931,N_2890);
nand U3360 (N_3360,N_2856,N_2681);
or U3361 (N_3361,N_2917,N_2623);
or U3362 (N_3362,N_2817,N_2606);
nand U3363 (N_3363,N_2706,N_2625);
or U3364 (N_3364,N_2728,N_2704);
and U3365 (N_3365,N_2746,N_2938);
or U3366 (N_3366,N_2636,N_2727);
nor U3367 (N_3367,N_2532,N_2876);
nand U3368 (N_3368,N_2854,N_2763);
nand U3369 (N_3369,N_2684,N_2986);
xnor U3370 (N_3370,N_2665,N_2513);
nand U3371 (N_3371,N_2554,N_2543);
or U3372 (N_3372,N_2954,N_2728);
xnor U3373 (N_3373,N_2758,N_2575);
and U3374 (N_3374,N_2722,N_2610);
and U3375 (N_3375,N_2644,N_2610);
nor U3376 (N_3376,N_2632,N_2664);
nand U3377 (N_3377,N_2709,N_2752);
nor U3378 (N_3378,N_2734,N_2526);
nor U3379 (N_3379,N_2811,N_2689);
or U3380 (N_3380,N_2800,N_2756);
and U3381 (N_3381,N_2974,N_2531);
or U3382 (N_3382,N_2575,N_2532);
and U3383 (N_3383,N_2937,N_2885);
nand U3384 (N_3384,N_2525,N_2572);
nand U3385 (N_3385,N_2993,N_2894);
and U3386 (N_3386,N_2647,N_2543);
or U3387 (N_3387,N_2834,N_2893);
and U3388 (N_3388,N_2827,N_2642);
and U3389 (N_3389,N_2652,N_2674);
xnor U3390 (N_3390,N_2588,N_2615);
nor U3391 (N_3391,N_2893,N_2615);
nor U3392 (N_3392,N_2967,N_2503);
nor U3393 (N_3393,N_2837,N_2620);
nor U3394 (N_3394,N_2578,N_2680);
or U3395 (N_3395,N_2989,N_2511);
and U3396 (N_3396,N_2708,N_2507);
and U3397 (N_3397,N_2567,N_2754);
or U3398 (N_3398,N_2959,N_2579);
nor U3399 (N_3399,N_2613,N_2937);
or U3400 (N_3400,N_2974,N_2868);
or U3401 (N_3401,N_2656,N_2567);
nand U3402 (N_3402,N_2889,N_2614);
or U3403 (N_3403,N_2840,N_2532);
nand U3404 (N_3404,N_2755,N_2693);
and U3405 (N_3405,N_2623,N_2801);
and U3406 (N_3406,N_2976,N_2790);
nor U3407 (N_3407,N_2666,N_2665);
nor U3408 (N_3408,N_2712,N_2554);
nand U3409 (N_3409,N_2697,N_2855);
or U3410 (N_3410,N_2857,N_2955);
nand U3411 (N_3411,N_2808,N_2851);
nor U3412 (N_3412,N_2563,N_2911);
nand U3413 (N_3413,N_2530,N_2569);
nor U3414 (N_3414,N_2751,N_2588);
or U3415 (N_3415,N_2533,N_2987);
and U3416 (N_3416,N_2646,N_2543);
or U3417 (N_3417,N_2929,N_2997);
and U3418 (N_3418,N_2652,N_2663);
and U3419 (N_3419,N_2768,N_2539);
nor U3420 (N_3420,N_2674,N_2756);
and U3421 (N_3421,N_2660,N_2932);
nor U3422 (N_3422,N_2579,N_2509);
and U3423 (N_3423,N_2745,N_2691);
and U3424 (N_3424,N_2507,N_2852);
nor U3425 (N_3425,N_2546,N_2830);
or U3426 (N_3426,N_2623,N_2540);
nand U3427 (N_3427,N_2539,N_2849);
or U3428 (N_3428,N_2769,N_2812);
and U3429 (N_3429,N_2872,N_2640);
or U3430 (N_3430,N_2875,N_2649);
nor U3431 (N_3431,N_2934,N_2824);
or U3432 (N_3432,N_2872,N_2757);
xnor U3433 (N_3433,N_2701,N_2920);
nand U3434 (N_3434,N_2948,N_2706);
xnor U3435 (N_3435,N_2748,N_2809);
nand U3436 (N_3436,N_2624,N_2751);
or U3437 (N_3437,N_2928,N_2802);
nand U3438 (N_3438,N_2764,N_2626);
and U3439 (N_3439,N_2881,N_2733);
and U3440 (N_3440,N_2798,N_2577);
nor U3441 (N_3441,N_2556,N_2914);
or U3442 (N_3442,N_2550,N_2627);
and U3443 (N_3443,N_2581,N_2566);
and U3444 (N_3444,N_2900,N_2838);
nand U3445 (N_3445,N_2751,N_2981);
and U3446 (N_3446,N_2937,N_2625);
xnor U3447 (N_3447,N_2585,N_2986);
or U3448 (N_3448,N_2958,N_2922);
and U3449 (N_3449,N_2802,N_2829);
or U3450 (N_3450,N_2592,N_2746);
nor U3451 (N_3451,N_2744,N_2961);
nand U3452 (N_3452,N_2766,N_2521);
and U3453 (N_3453,N_2584,N_2679);
and U3454 (N_3454,N_2537,N_2501);
and U3455 (N_3455,N_2657,N_2768);
nand U3456 (N_3456,N_2904,N_2970);
or U3457 (N_3457,N_2876,N_2640);
nand U3458 (N_3458,N_2557,N_2632);
nand U3459 (N_3459,N_2967,N_2540);
nor U3460 (N_3460,N_2657,N_2800);
nand U3461 (N_3461,N_2553,N_2837);
nand U3462 (N_3462,N_2538,N_2762);
and U3463 (N_3463,N_2622,N_2634);
nor U3464 (N_3464,N_2963,N_2878);
and U3465 (N_3465,N_2613,N_2976);
and U3466 (N_3466,N_2689,N_2902);
or U3467 (N_3467,N_2767,N_2649);
or U3468 (N_3468,N_2727,N_2987);
and U3469 (N_3469,N_2955,N_2842);
or U3470 (N_3470,N_2788,N_2932);
nor U3471 (N_3471,N_2794,N_2596);
nand U3472 (N_3472,N_2962,N_2559);
or U3473 (N_3473,N_2708,N_2822);
nor U3474 (N_3474,N_2869,N_2791);
and U3475 (N_3475,N_2572,N_2842);
nor U3476 (N_3476,N_2570,N_2797);
nand U3477 (N_3477,N_2901,N_2961);
or U3478 (N_3478,N_2942,N_2929);
nor U3479 (N_3479,N_2901,N_2648);
and U3480 (N_3480,N_2759,N_2815);
nor U3481 (N_3481,N_2948,N_2772);
nand U3482 (N_3482,N_2623,N_2513);
or U3483 (N_3483,N_2981,N_2512);
nor U3484 (N_3484,N_2917,N_2781);
nand U3485 (N_3485,N_2987,N_2674);
or U3486 (N_3486,N_2805,N_2802);
and U3487 (N_3487,N_2571,N_2605);
or U3488 (N_3488,N_2873,N_2762);
nand U3489 (N_3489,N_2643,N_2599);
and U3490 (N_3490,N_2536,N_2680);
nand U3491 (N_3491,N_2647,N_2990);
or U3492 (N_3492,N_2605,N_2841);
or U3493 (N_3493,N_2612,N_2576);
nor U3494 (N_3494,N_2940,N_2538);
or U3495 (N_3495,N_2559,N_2801);
nor U3496 (N_3496,N_2820,N_2507);
or U3497 (N_3497,N_2574,N_2882);
nor U3498 (N_3498,N_2915,N_2704);
nor U3499 (N_3499,N_2954,N_2885);
nand U3500 (N_3500,N_3210,N_3289);
nand U3501 (N_3501,N_3466,N_3155);
or U3502 (N_3502,N_3420,N_3045);
and U3503 (N_3503,N_3318,N_3224);
nand U3504 (N_3504,N_3342,N_3140);
nor U3505 (N_3505,N_3195,N_3379);
nand U3506 (N_3506,N_3041,N_3256);
nand U3507 (N_3507,N_3075,N_3095);
nor U3508 (N_3508,N_3356,N_3015);
or U3509 (N_3509,N_3108,N_3294);
and U3510 (N_3510,N_3232,N_3286);
nand U3511 (N_3511,N_3479,N_3246);
nor U3512 (N_3512,N_3101,N_3206);
and U3513 (N_3513,N_3085,N_3281);
or U3514 (N_3514,N_3414,N_3300);
or U3515 (N_3515,N_3486,N_3469);
or U3516 (N_3516,N_3497,N_3396);
and U3517 (N_3517,N_3129,N_3311);
nor U3518 (N_3518,N_3495,N_3453);
or U3519 (N_3519,N_3442,N_3080);
and U3520 (N_3520,N_3407,N_3054);
or U3521 (N_3521,N_3038,N_3242);
nand U3522 (N_3522,N_3384,N_3128);
or U3523 (N_3523,N_3399,N_3274);
or U3524 (N_3524,N_3416,N_3471);
and U3525 (N_3525,N_3005,N_3426);
nand U3526 (N_3526,N_3099,N_3487);
and U3527 (N_3527,N_3457,N_3068);
and U3528 (N_3528,N_3081,N_3402);
nor U3529 (N_3529,N_3354,N_3348);
and U3530 (N_3530,N_3197,N_3389);
and U3531 (N_3531,N_3103,N_3371);
and U3532 (N_3532,N_3102,N_3124);
nand U3533 (N_3533,N_3222,N_3106);
and U3534 (N_3534,N_3316,N_3186);
nor U3535 (N_3535,N_3317,N_3199);
nand U3536 (N_3536,N_3233,N_3474);
nand U3537 (N_3537,N_3401,N_3137);
and U3538 (N_3538,N_3024,N_3205);
nor U3539 (N_3539,N_3069,N_3488);
nand U3540 (N_3540,N_3044,N_3309);
nor U3541 (N_3541,N_3033,N_3121);
nand U3542 (N_3542,N_3392,N_3091);
nor U3543 (N_3543,N_3208,N_3018);
or U3544 (N_3544,N_3404,N_3134);
nor U3545 (N_3545,N_3008,N_3415);
and U3546 (N_3546,N_3056,N_3386);
or U3547 (N_3547,N_3174,N_3329);
or U3548 (N_3548,N_3461,N_3340);
or U3549 (N_3549,N_3359,N_3200);
nor U3550 (N_3550,N_3492,N_3111);
or U3551 (N_3551,N_3136,N_3336);
nand U3552 (N_3552,N_3169,N_3219);
and U3553 (N_3553,N_3436,N_3296);
or U3554 (N_3554,N_3409,N_3283);
nor U3555 (N_3555,N_3123,N_3025);
nor U3556 (N_3556,N_3084,N_3373);
nand U3557 (N_3557,N_3393,N_3427);
nor U3558 (N_3558,N_3417,N_3422);
nand U3559 (N_3559,N_3353,N_3484);
nor U3560 (N_3560,N_3451,N_3395);
nor U3561 (N_3561,N_3273,N_3230);
and U3562 (N_3562,N_3258,N_3363);
and U3563 (N_3563,N_3429,N_3170);
xnor U3564 (N_3564,N_3268,N_3221);
nand U3565 (N_3565,N_3007,N_3262);
or U3566 (N_3566,N_3446,N_3034);
xor U3567 (N_3567,N_3064,N_3467);
or U3568 (N_3568,N_3398,N_3066);
or U3569 (N_3569,N_3345,N_3027);
nor U3570 (N_3570,N_3308,N_3010);
and U3571 (N_3571,N_3026,N_3439);
nor U3572 (N_3572,N_3368,N_3198);
and U3573 (N_3573,N_3096,N_3153);
and U3574 (N_3574,N_3328,N_3423);
and U3575 (N_3575,N_3382,N_3113);
or U3576 (N_3576,N_3473,N_3369);
or U3577 (N_3577,N_3241,N_3278);
nand U3578 (N_3578,N_3297,N_3410);
or U3579 (N_3579,N_3358,N_3254);
nand U3580 (N_3580,N_3158,N_3046);
nand U3581 (N_3581,N_3196,N_3364);
nor U3582 (N_3582,N_3039,N_3352);
nor U3583 (N_3583,N_3138,N_3092);
nand U3584 (N_3584,N_3441,N_3370);
nor U3585 (N_3585,N_3483,N_3139);
and U3586 (N_3586,N_3157,N_3154);
nand U3587 (N_3587,N_3413,N_3491);
nand U3588 (N_3588,N_3141,N_3421);
or U3589 (N_3589,N_3164,N_3459);
nor U3590 (N_3590,N_3490,N_3076);
and U3591 (N_3591,N_3152,N_3288);
and U3592 (N_3592,N_3260,N_3263);
and U3593 (N_3593,N_3387,N_3276);
nand U3594 (N_3594,N_3133,N_3463);
and U3595 (N_3595,N_3062,N_3207);
nor U3596 (N_3596,N_3408,N_3225);
nand U3597 (N_3597,N_3072,N_3179);
xnor U3598 (N_3598,N_3234,N_3482);
or U3599 (N_3599,N_3259,N_3468);
nand U3600 (N_3600,N_3144,N_3073);
nand U3601 (N_3601,N_3160,N_3029);
nor U3602 (N_3602,N_3333,N_3462);
or U3603 (N_3603,N_3265,N_3238);
or U3604 (N_3604,N_3023,N_3394);
nand U3605 (N_3605,N_3285,N_3397);
and U3606 (N_3606,N_3209,N_3452);
and U3607 (N_3607,N_3424,N_3330);
xor U3608 (N_3608,N_3435,N_3456);
nand U3609 (N_3609,N_3334,N_3177);
nand U3610 (N_3610,N_3390,N_3019);
nor U3611 (N_3611,N_3269,N_3063);
or U3612 (N_3612,N_3455,N_3312);
nand U3613 (N_3613,N_3212,N_3086);
or U3614 (N_3614,N_3496,N_3322);
nand U3615 (N_3615,N_3264,N_3118);
and U3616 (N_3616,N_3295,N_3251);
or U3617 (N_3617,N_3163,N_3002);
or U3618 (N_3618,N_3105,N_3070);
nand U3619 (N_3619,N_3245,N_3282);
nor U3620 (N_3620,N_3303,N_3248);
or U3621 (N_3621,N_3290,N_3252);
nand U3622 (N_3622,N_3165,N_3301);
nor U3623 (N_3623,N_3302,N_3009);
or U3624 (N_3624,N_3065,N_3151);
and U3625 (N_3625,N_3217,N_3112);
and U3626 (N_3626,N_3449,N_3050);
or U3627 (N_3627,N_3257,N_3189);
or U3628 (N_3628,N_3305,N_3057);
nor U3629 (N_3629,N_3173,N_3465);
nand U3630 (N_3630,N_3425,N_3437);
or U3631 (N_3631,N_3287,N_3337);
and U3632 (N_3632,N_3114,N_3040);
xor U3633 (N_3633,N_3403,N_3047);
nand U3634 (N_3634,N_3020,N_3343);
nand U3635 (N_3635,N_3377,N_3203);
nand U3636 (N_3636,N_3476,N_3097);
and U3637 (N_3637,N_3012,N_3381);
nand U3638 (N_3638,N_3194,N_3104);
and U3639 (N_3639,N_3226,N_3182);
or U3640 (N_3640,N_3279,N_3087);
and U3641 (N_3641,N_3411,N_3166);
nor U3642 (N_3642,N_3385,N_3349);
xor U3643 (N_3643,N_3093,N_3214);
nand U3644 (N_3644,N_3418,N_3115);
nor U3645 (N_3645,N_3376,N_3176);
nand U3646 (N_3646,N_3351,N_3237);
and U3647 (N_3647,N_3172,N_3130);
or U3648 (N_3648,N_3324,N_3499);
nand U3649 (N_3649,N_3431,N_3339);
xnor U3650 (N_3650,N_3161,N_3321);
nand U3651 (N_3651,N_3307,N_3053);
nand U3652 (N_3652,N_3255,N_3185);
nor U3653 (N_3653,N_3247,N_3098);
or U3654 (N_3654,N_3277,N_3250);
or U3655 (N_3655,N_3119,N_3167);
or U3656 (N_3656,N_3231,N_3135);
or U3657 (N_3657,N_3021,N_3036);
nor U3658 (N_3658,N_3261,N_3310);
or U3659 (N_3659,N_3481,N_3372);
nand U3660 (N_3660,N_3458,N_3017);
and U3661 (N_3661,N_3314,N_3156);
nor U3662 (N_3662,N_3227,N_3454);
and U3663 (N_3663,N_3275,N_3052);
nand U3664 (N_3664,N_3145,N_3272);
and U3665 (N_3665,N_3074,N_3299);
nand U3666 (N_3666,N_3146,N_3148);
or U3667 (N_3667,N_3088,N_3071);
nor U3668 (N_3668,N_3006,N_3228);
nand U3669 (N_3669,N_3323,N_3178);
or U3670 (N_3670,N_3215,N_3320);
and U3671 (N_3671,N_3043,N_3444);
or U3672 (N_3672,N_3443,N_3201);
nor U3673 (N_3673,N_3315,N_3122);
nand U3674 (N_3674,N_3346,N_3357);
and U3675 (N_3675,N_3235,N_3031);
nor U3676 (N_3676,N_3478,N_3168);
and U3677 (N_3677,N_3022,N_3460);
and U3678 (N_3678,N_3191,N_3132);
nor U3679 (N_3679,N_3110,N_3082);
and U3680 (N_3680,N_3109,N_3058);
xor U3681 (N_3681,N_3445,N_3366);
nand U3682 (N_3682,N_3059,N_3216);
nand U3683 (N_3683,N_3107,N_3100);
nand U3684 (N_3684,N_3035,N_3298);
nor U3685 (N_3685,N_3438,N_3266);
nand U3686 (N_3686,N_3051,N_3480);
nand U3687 (N_3687,N_3190,N_3338);
or U3688 (N_3688,N_3406,N_3188);
nand U3689 (N_3689,N_3477,N_3094);
nand U3690 (N_3690,N_3204,N_3131);
nor U3691 (N_3691,N_3313,N_3360);
nor U3692 (N_3692,N_3048,N_3470);
or U3693 (N_3693,N_3150,N_3223);
nor U3694 (N_3694,N_3028,N_3055);
or U3695 (N_3695,N_3464,N_3253);
and U3696 (N_3696,N_3220,N_3037);
and U3697 (N_3697,N_3236,N_3412);
and U3698 (N_3698,N_3331,N_3159);
nor U3699 (N_3699,N_3147,N_3347);
or U3700 (N_3700,N_3011,N_3249);
nor U3701 (N_3701,N_3089,N_3375);
nor U3702 (N_3702,N_3493,N_3293);
and U3703 (N_3703,N_3291,N_3117);
nor U3704 (N_3704,N_3187,N_3432);
and U3705 (N_3705,N_3494,N_3125);
nor U3706 (N_3706,N_3284,N_3400);
or U3707 (N_3707,N_3270,N_3430);
or U3708 (N_3708,N_3183,N_3327);
or U3709 (N_3709,N_3171,N_3365);
or U3710 (N_3710,N_3202,N_3042);
or U3711 (N_3711,N_3448,N_3447);
nand U3712 (N_3712,N_3292,N_3014);
xnor U3713 (N_3713,N_3001,N_3361);
or U3714 (N_3714,N_3243,N_3142);
and U3715 (N_3715,N_3060,N_3355);
and U3716 (N_3716,N_3061,N_3120);
or U3717 (N_3717,N_3485,N_3350);
nor U3718 (N_3718,N_3049,N_3374);
nor U3719 (N_3719,N_3489,N_3218);
or U3720 (N_3720,N_3180,N_3332);
or U3721 (N_3721,N_3083,N_3433);
or U3722 (N_3722,N_3362,N_3267);
nand U3723 (N_3723,N_3388,N_3271);
or U3724 (N_3724,N_3383,N_3149);
or U3725 (N_3725,N_3440,N_3143);
or U3726 (N_3726,N_3240,N_3326);
or U3727 (N_3727,N_3030,N_3078);
nor U3728 (N_3728,N_3498,N_3067);
nor U3729 (N_3729,N_3335,N_3181);
or U3730 (N_3730,N_3032,N_3367);
and U3731 (N_3731,N_3175,N_3116);
and U3732 (N_3732,N_3419,N_3378);
nand U3733 (N_3733,N_3380,N_3184);
nand U3734 (N_3734,N_3450,N_3306);
and U3735 (N_3735,N_3013,N_3341);
or U3736 (N_3736,N_3162,N_3229);
xor U3737 (N_3737,N_3405,N_3127);
nand U3738 (N_3738,N_3325,N_3090);
nor U3739 (N_3739,N_3077,N_3004);
or U3740 (N_3740,N_3244,N_3434);
nand U3741 (N_3741,N_3391,N_3213);
and U3742 (N_3742,N_3000,N_3319);
nor U3743 (N_3743,N_3016,N_3428);
nand U3744 (N_3744,N_3280,N_3211);
or U3745 (N_3745,N_3344,N_3475);
nand U3746 (N_3746,N_3192,N_3193);
nand U3747 (N_3747,N_3304,N_3079);
nand U3748 (N_3748,N_3126,N_3472);
nand U3749 (N_3749,N_3003,N_3239);
and U3750 (N_3750,N_3132,N_3411);
nand U3751 (N_3751,N_3326,N_3372);
and U3752 (N_3752,N_3134,N_3433);
or U3753 (N_3753,N_3290,N_3129);
nor U3754 (N_3754,N_3433,N_3487);
and U3755 (N_3755,N_3393,N_3435);
or U3756 (N_3756,N_3324,N_3174);
nand U3757 (N_3757,N_3075,N_3120);
nand U3758 (N_3758,N_3283,N_3253);
or U3759 (N_3759,N_3256,N_3418);
and U3760 (N_3760,N_3143,N_3313);
nand U3761 (N_3761,N_3122,N_3098);
and U3762 (N_3762,N_3287,N_3052);
nor U3763 (N_3763,N_3025,N_3092);
nand U3764 (N_3764,N_3270,N_3277);
nor U3765 (N_3765,N_3269,N_3133);
nor U3766 (N_3766,N_3337,N_3191);
nor U3767 (N_3767,N_3481,N_3457);
nand U3768 (N_3768,N_3245,N_3205);
nand U3769 (N_3769,N_3428,N_3346);
nand U3770 (N_3770,N_3499,N_3249);
and U3771 (N_3771,N_3183,N_3024);
or U3772 (N_3772,N_3174,N_3367);
nand U3773 (N_3773,N_3362,N_3442);
nor U3774 (N_3774,N_3058,N_3186);
nand U3775 (N_3775,N_3383,N_3479);
and U3776 (N_3776,N_3315,N_3251);
or U3777 (N_3777,N_3499,N_3043);
nand U3778 (N_3778,N_3084,N_3439);
nand U3779 (N_3779,N_3482,N_3396);
and U3780 (N_3780,N_3439,N_3210);
nor U3781 (N_3781,N_3122,N_3286);
nand U3782 (N_3782,N_3102,N_3473);
and U3783 (N_3783,N_3050,N_3459);
nand U3784 (N_3784,N_3298,N_3272);
and U3785 (N_3785,N_3286,N_3307);
nor U3786 (N_3786,N_3388,N_3328);
and U3787 (N_3787,N_3319,N_3244);
nand U3788 (N_3788,N_3160,N_3352);
nor U3789 (N_3789,N_3053,N_3234);
and U3790 (N_3790,N_3347,N_3482);
and U3791 (N_3791,N_3351,N_3112);
and U3792 (N_3792,N_3008,N_3139);
xor U3793 (N_3793,N_3256,N_3171);
nor U3794 (N_3794,N_3172,N_3113);
nand U3795 (N_3795,N_3402,N_3219);
and U3796 (N_3796,N_3326,N_3120);
or U3797 (N_3797,N_3044,N_3323);
xor U3798 (N_3798,N_3325,N_3427);
xor U3799 (N_3799,N_3146,N_3038);
or U3800 (N_3800,N_3166,N_3264);
nor U3801 (N_3801,N_3109,N_3318);
and U3802 (N_3802,N_3381,N_3453);
xor U3803 (N_3803,N_3418,N_3275);
nor U3804 (N_3804,N_3270,N_3151);
or U3805 (N_3805,N_3008,N_3215);
nand U3806 (N_3806,N_3023,N_3140);
nor U3807 (N_3807,N_3191,N_3201);
nand U3808 (N_3808,N_3071,N_3320);
xor U3809 (N_3809,N_3052,N_3263);
xor U3810 (N_3810,N_3462,N_3430);
and U3811 (N_3811,N_3482,N_3405);
nand U3812 (N_3812,N_3471,N_3402);
and U3813 (N_3813,N_3446,N_3090);
nor U3814 (N_3814,N_3157,N_3287);
and U3815 (N_3815,N_3180,N_3439);
or U3816 (N_3816,N_3308,N_3192);
nand U3817 (N_3817,N_3257,N_3480);
nand U3818 (N_3818,N_3405,N_3473);
nand U3819 (N_3819,N_3023,N_3273);
and U3820 (N_3820,N_3266,N_3021);
nand U3821 (N_3821,N_3234,N_3207);
nor U3822 (N_3822,N_3123,N_3419);
or U3823 (N_3823,N_3063,N_3191);
and U3824 (N_3824,N_3188,N_3403);
or U3825 (N_3825,N_3149,N_3066);
or U3826 (N_3826,N_3335,N_3090);
nor U3827 (N_3827,N_3355,N_3171);
nand U3828 (N_3828,N_3088,N_3335);
or U3829 (N_3829,N_3453,N_3066);
or U3830 (N_3830,N_3068,N_3093);
nor U3831 (N_3831,N_3361,N_3296);
nor U3832 (N_3832,N_3498,N_3231);
nor U3833 (N_3833,N_3115,N_3474);
nand U3834 (N_3834,N_3204,N_3109);
or U3835 (N_3835,N_3226,N_3151);
nor U3836 (N_3836,N_3418,N_3083);
or U3837 (N_3837,N_3021,N_3156);
and U3838 (N_3838,N_3487,N_3079);
and U3839 (N_3839,N_3016,N_3147);
nand U3840 (N_3840,N_3498,N_3417);
nand U3841 (N_3841,N_3158,N_3296);
and U3842 (N_3842,N_3065,N_3467);
nand U3843 (N_3843,N_3248,N_3013);
nand U3844 (N_3844,N_3248,N_3436);
and U3845 (N_3845,N_3072,N_3495);
or U3846 (N_3846,N_3348,N_3319);
nor U3847 (N_3847,N_3032,N_3003);
and U3848 (N_3848,N_3243,N_3414);
nand U3849 (N_3849,N_3017,N_3042);
nand U3850 (N_3850,N_3347,N_3405);
or U3851 (N_3851,N_3496,N_3284);
nand U3852 (N_3852,N_3388,N_3094);
or U3853 (N_3853,N_3024,N_3042);
nand U3854 (N_3854,N_3063,N_3366);
and U3855 (N_3855,N_3026,N_3430);
and U3856 (N_3856,N_3454,N_3494);
or U3857 (N_3857,N_3122,N_3403);
or U3858 (N_3858,N_3151,N_3374);
nor U3859 (N_3859,N_3129,N_3348);
nor U3860 (N_3860,N_3240,N_3320);
nand U3861 (N_3861,N_3350,N_3351);
nand U3862 (N_3862,N_3299,N_3321);
nand U3863 (N_3863,N_3270,N_3149);
or U3864 (N_3864,N_3230,N_3202);
and U3865 (N_3865,N_3361,N_3031);
nor U3866 (N_3866,N_3446,N_3342);
or U3867 (N_3867,N_3258,N_3329);
nand U3868 (N_3868,N_3088,N_3251);
or U3869 (N_3869,N_3496,N_3340);
nand U3870 (N_3870,N_3241,N_3083);
or U3871 (N_3871,N_3011,N_3417);
or U3872 (N_3872,N_3406,N_3017);
and U3873 (N_3873,N_3398,N_3018);
nand U3874 (N_3874,N_3442,N_3181);
nand U3875 (N_3875,N_3136,N_3135);
or U3876 (N_3876,N_3401,N_3399);
nand U3877 (N_3877,N_3162,N_3164);
and U3878 (N_3878,N_3239,N_3470);
nand U3879 (N_3879,N_3147,N_3465);
nor U3880 (N_3880,N_3147,N_3061);
nand U3881 (N_3881,N_3185,N_3328);
or U3882 (N_3882,N_3131,N_3497);
nand U3883 (N_3883,N_3478,N_3419);
nor U3884 (N_3884,N_3400,N_3285);
nand U3885 (N_3885,N_3288,N_3034);
and U3886 (N_3886,N_3446,N_3137);
or U3887 (N_3887,N_3028,N_3062);
nor U3888 (N_3888,N_3170,N_3342);
or U3889 (N_3889,N_3451,N_3438);
or U3890 (N_3890,N_3139,N_3329);
or U3891 (N_3891,N_3064,N_3293);
nor U3892 (N_3892,N_3388,N_3406);
nor U3893 (N_3893,N_3049,N_3011);
nand U3894 (N_3894,N_3361,N_3067);
or U3895 (N_3895,N_3451,N_3343);
nand U3896 (N_3896,N_3023,N_3162);
or U3897 (N_3897,N_3136,N_3045);
or U3898 (N_3898,N_3404,N_3298);
or U3899 (N_3899,N_3038,N_3425);
nand U3900 (N_3900,N_3152,N_3340);
and U3901 (N_3901,N_3440,N_3429);
or U3902 (N_3902,N_3393,N_3108);
nand U3903 (N_3903,N_3205,N_3101);
nand U3904 (N_3904,N_3305,N_3172);
nor U3905 (N_3905,N_3159,N_3425);
xor U3906 (N_3906,N_3324,N_3306);
and U3907 (N_3907,N_3033,N_3498);
xor U3908 (N_3908,N_3092,N_3142);
nand U3909 (N_3909,N_3020,N_3296);
nor U3910 (N_3910,N_3162,N_3252);
or U3911 (N_3911,N_3491,N_3401);
and U3912 (N_3912,N_3193,N_3085);
or U3913 (N_3913,N_3257,N_3332);
or U3914 (N_3914,N_3007,N_3296);
or U3915 (N_3915,N_3156,N_3057);
and U3916 (N_3916,N_3133,N_3448);
and U3917 (N_3917,N_3305,N_3457);
or U3918 (N_3918,N_3462,N_3181);
nand U3919 (N_3919,N_3187,N_3011);
or U3920 (N_3920,N_3153,N_3375);
or U3921 (N_3921,N_3065,N_3262);
nand U3922 (N_3922,N_3345,N_3411);
nand U3923 (N_3923,N_3314,N_3126);
xnor U3924 (N_3924,N_3219,N_3454);
or U3925 (N_3925,N_3449,N_3226);
or U3926 (N_3926,N_3252,N_3161);
or U3927 (N_3927,N_3397,N_3167);
nor U3928 (N_3928,N_3029,N_3468);
nand U3929 (N_3929,N_3322,N_3181);
nand U3930 (N_3930,N_3068,N_3371);
nor U3931 (N_3931,N_3215,N_3364);
and U3932 (N_3932,N_3425,N_3457);
nor U3933 (N_3933,N_3473,N_3297);
xor U3934 (N_3934,N_3305,N_3029);
nand U3935 (N_3935,N_3032,N_3102);
nor U3936 (N_3936,N_3040,N_3105);
nor U3937 (N_3937,N_3333,N_3038);
nor U3938 (N_3938,N_3369,N_3409);
nor U3939 (N_3939,N_3490,N_3051);
and U3940 (N_3940,N_3447,N_3205);
nor U3941 (N_3941,N_3319,N_3284);
and U3942 (N_3942,N_3443,N_3109);
nor U3943 (N_3943,N_3219,N_3145);
or U3944 (N_3944,N_3402,N_3495);
nand U3945 (N_3945,N_3493,N_3062);
nor U3946 (N_3946,N_3013,N_3116);
nand U3947 (N_3947,N_3171,N_3029);
xor U3948 (N_3948,N_3432,N_3256);
nand U3949 (N_3949,N_3025,N_3120);
and U3950 (N_3950,N_3079,N_3025);
or U3951 (N_3951,N_3151,N_3141);
nor U3952 (N_3952,N_3272,N_3299);
and U3953 (N_3953,N_3419,N_3218);
or U3954 (N_3954,N_3413,N_3392);
nand U3955 (N_3955,N_3281,N_3011);
or U3956 (N_3956,N_3355,N_3398);
or U3957 (N_3957,N_3458,N_3336);
nand U3958 (N_3958,N_3226,N_3249);
or U3959 (N_3959,N_3064,N_3097);
and U3960 (N_3960,N_3123,N_3358);
and U3961 (N_3961,N_3318,N_3091);
and U3962 (N_3962,N_3044,N_3145);
nand U3963 (N_3963,N_3006,N_3454);
and U3964 (N_3964,N_3050,N_3040);
xnor U3965 (N_3965,N_3442,N_3464);
nor U3966 (N_3966,N_3410,N_3227);
nor U3967 (N_3967,N_3222,N_3000);
and U3968 (N_3968,N_3322,N_3128);
and U3969 (N_3969,N_3377,N_3019);
and U3970 (N_3970,N_3298,N_3273);
nor U3971 (N_3971,N_3012,N_3277);
or U3972 (N_3972,N_3202,N_3255);
and U3973 (N_3973,N_3004,N_3278);
and U3974 (N_3974,N_3481,N_3355);
or U3975 (N_3975,N_3047,N_3048);
nand U3976 (N_3976,N_3068,N_3108);
nand U3977 (N_3977,N_3103,N_3322);
nor U3978 (N_3978,N_3008,N_3308);
and U3979 (N_3979,N_3100,N_3178);
or U3980 (N_3980,N_3475,N_3094);
or U3981 (N_3981,N_3153,N_3075);
nand U3982 (N_3982,N_3138,N_3427);
xnor U3983 (N_3983,N_3281,N_3353);
or U3984 (N_3984,N_3123,N_3041);
or U3985 (N_3985,N_3132,N_3162);
and U3986 (N_3986,N_3148,N_3483);
nand U3987 (N_3987,N_3173,N_3356);
nand U3988 (N_3988,N_3317,N_3201);
nor U3989 (N_3989,N_3392,N_3477);
nor U3990 (N_3990,N_3416,N_3417);
or U3991 (N_3991,N_3058,N_3134);
nor U3992 (N_3992,N_3098,N_3279);
or U3993 (N_3993,N_3379,N_3257);
and U3994 (N_3994,N_3341,N_3006);
nand U3995 (N_3995,N_3098,N_3467);
and U3996 (N_3996,N_3228,N_3351);
nor U3997 (N_3997,N_3484,N_3189);
nand U3998 (N_3998,N_3405,N_3142);
or U3999 (N_3999,N_3474,N_3008);
and U4000 (N_4000,N_3554,N_3574);
nand U4001 (N_4001,N_3994,N_3535);
and U4002 (N_4002,N_3753,N_3548);
or U4003 (N_4003,N_3807,N_3969);
and U4004 (N_4004,N_3926,N_3594);
nand U4005 (N_4005,N_3788,N_3938);
nor U4006 (N_4006,N_3913,N_3771);
nor U4007 (N_4007,N_3539,N_3579);
nor U4008 (N_4008,N_3756,N_3501);
nor U4009 (N_4009,N_3931,N_3744);
nor U4010 (N_4010,N_3989,N_3860);
nand U4011 (N_4011,N_3734,N_3655);
nor U4012 (N_4012,N_3722,N_3985);
nand U4013 (N_4013,N_3766,N_3506);
or U4014 (N_4014,N_3615,N_3859);
nor U4015 (N_4015,N_3853,N_3557);
nand U4016 (N_4016,N_3808,N_3778);
and U4017 (N_4017,N_3703,N_3769);
xnor U4018 (N_4018,N_3811,N_3891);
nor U4019 (N_4019,N_3805,N_3743);
and U4020 (N_4020,N_3897,N_3698);
and U4021 (N_4021,N_3683,N_3503);
and U4022 (N_4022,N_3510,N_3632);
nor U4023 (N_4023,N_3881,N_3694);
nor U4024 (N_4024,N_3532,N_3739);
nor U4025 (N_4025,N_3874,N_3563);
and U4026 (N_4026,N_3907,N_3841);
nor U4027 (N_4027,N_3820,N_3512);
and U4028 (N_4028,N_3710,N_3616);
or U4029 (N_4029,N_3542,N_3997);
nor U4030 (N_4030,N_3957,N_3815);
nand U4031 (N_4031,N_3697,N_3849);
and U4032 (N_4032,N_3592,N_3861);
nor U4033 (N_4033,N_3544,N_3568);
or U4034 (N_4034,N_3593,N_3573);
nand U4035 (N_4035,N_3831,N_3970);
nand U4036 (N_4036,N_3966,N_3791);
nor U4037 (N_4037,N_3757,N_3732);
or U4038 (N_4038,N_3814,N_3755);
or U4039 (N_4039,N_3726,N_3680);
and U4040 (N_4040,N_3719,N_3876);
and U4041 (N_4041,N_3928,N_3991);
nor U4042 (N_4042,N_3656,N_3644);
or U4043 (N_4043,N_3772,N_3924);
or U4044 (N_4044,N_3792,N_3585);
or U4045 (N_4045,N_3519,N_3937);
nor U4046 (N_4046,N_3652,N_3664);
nand U4047 (N_4047,N_3671,N_3536);
or U4048 (N_4048,N_3785,N_3882);
and U4049 (N_4049,N_3962,N_3500);
nand U4050 (N_4050,N_3647,N_3560);
or U4051 (N_4051,N_3699,N_3550);
nand U4052 (N_4052,N_3848,N_3668);
nand U4053 (N_4053,N_3687,N_3827);
nor U4054 (N_4054,N_3906,N_3638);
nor U4055 (N_4055,N_3953,N_3529);
and U4056 (N_4056,N_3528,N_3727);
or U4057 (N_4057,N_3566,N_3975);
nor U4058 (N_4058,N_3794,N_3718);
nor U4059 (N_4059,N_3916,N_3598);
nor U4060 (N_4060,N_3576,N_3803);
and U4061 (N_4061,N_3624,N_3783);
nand U4062 (N_4062,N_3714,N_3603);
nor U4063 (N_4063,N_3625,N_3992);
and U4064 (N_4064,N_3707,N_3915);
nand U4065 (N_4065,N_3717,N_3621);
or U4066 (N_4066,N_3902,N_3677);
xor U4067 (N_4067,N_3949,N_3705);
or U4068 (N_4068,N_3741,N_3750);
nand U4069 (N_4069,N_3526,N_3672);
nand U4070 (N_4070,N_3582,N_3998);
nor U4071 (N_4071,N_3667,N_3978);
or U4072 (N_4072,N_3940,N_3782);
and U4073 (N_4073,N_3885,N_3922);
and U4074 (N_4074,N_3731,N_3684);
or U4075 (N_4075,N_3516,N_3821);
nor U4076 (N_4076,N_3565,N_3927);
or U4077 (N_4077,N_3908,N_3980);
nor U4078 (N_4078,N_3875,N_3552);
nor U4079 (N_4079,N_3702,N_3765);
or U4080 (N_4080,N_3654,N_3724);
nand U4081 (N_4081,N_3903,N_3990);
and U4082 (N_4082,N_3581,N_3754);
nor U4083 (N_4083,N_3633,N_3596);
nor U4084 (N_4084,N_3781,N_3511);
nor U4085 (N_4085,N_3762,N_3575);
or U4086 (N_4086,N_3999,N_3641);
or U4087 (N_4087,N_3838,N_3745);
and U4088 (N_4088,N_3917,N_3900);
or U4089 (N_4089,N_3706,N_3823);
nand U4090 (N_4090,N_3643,N_3879);
and U4091 (N_4091,N_3619,N_3629);
nand U4092 (N_4092,N_3716,N_3610);
and U4093 (N_4093,N_3767,N_3899);
nor U4094 (N_4094,N_3651,N_3547);
nand U4095 (N_4095,N_3972,N_3843);
and U4096 (N_4096,N_3746,N_3884);
or U4097 (N_4097,N_3936,N_3558);
and U4098 (N_4098,N_3971,N_3932);
or U4099 (N_4099,N_3862,N_3824);
and U4100 (N_4100,N_3967,N_3840);
and U4101 (N_4101,N_3649,N_3946);
nand U4102 (N_4102,N_3645,N_3965);
or U4103 (N_4103,N_3636,N_3919);
nor U4104 (N_4104,N_3695,N_3742);
nor U4105 (N_4105,N_3779,N_3872);
or U4106 (N_4106,N_3894,N_3770);
nor U4107 (N_4107,N_3798,N_3836);
or U4108 (N_4108,N_3774,N_3842);
nor U4109 (N_4109,N_3736,N_3693);
and U4110 (N_4110,N_3630,N_3800);
and U4111 (N_4111,N_3961,N_3870);
xnor U4112 (N_4112,N_3889,N_3704);
and U4113 (N_4113,N_3696,N_3611);
nand U4114 (N_4114,N_3733,N_3835);
nand U4115 (N_4115,N_3887,N_3752);
nor U4116 (N_4116,N_3773,N_3674);
nand U4117 (N_4117,N_3597,N_3521);
and U4118 (N_4118,N_3634,N_3845);
or U4119 (N_4119,N_3572,N_3983);
and U4120 (N_4120,N_3730,N_3570);
or U4121 (N_4121,N_3631,N_3586);
nor U4122 (N_4122,N_3987,N_3604);
and U4123 (N_4123,N_3748,N_3896);
nor U4124 (N_4124,N_3858,N_3540);
and U4125 (N_4125,N_3768,N_3981);
and U4126 (N_4126,N_3578,N_3751);
or U4127 (N_4127,N_3819,N_3883);
or U4128 (N_4128,N_3945,N_3832);
nand U4129 (N_4129,N_3583,N_3601);
or U4130 (N_4130,N_3893,N_3691);
nand U4131 (N_4131,N_3974,N_3627);
or U4132 (N_4132,N_3725,N_3559);
nor U4133 (N_4133,N_3729,N_3888);
and U4134 (N_4134,N_3564,N_3640);
or U4135 (N_4135,N_3681,N_3986);
nand U4136 (N_4136,N_3923,N_3648);
nor U4137 (N_4137,N_3657,N_3609);
and U4138 (N_4138,N_3660,N_3850);
nand U4139 (N_4139,N_3786,N_3963);
and U4140 (N_4140,N_3780,N_3721);
and U4141 (N_4141,N_3712,N_3720);
or U4142 (N_4142,N_3761,N_3984);
nor U4143 (N_4143,N_3968,N_3549);
nand U4144 (N_4144,N_3837,N_3555);
nor U4145 (N_4145,N_3665,N_3878);
nor U4146 (N_4146,N_3912,N_3605);
nand U4147 (N_4147,N_3622,N_3877);
nand U4148 (N_4148,N_3826,N_3759);
and U4149 (N_4149,N_3670,N_3905);
and U4150 (N_4150,N_3934,N_3700);
nor U4151 (N_4151,N_3809,N_3587);
nor U4152 (N_4152,N_3607,N_3628);
nand U4153 (N_4153,N_3517,N_3747);
or U4154 (N_4154,N_3639,N_3688);
or U4155 (N_4155,N_3737,N_3749);
nand U4156 (N_4156,N_3663,N_3538);
nor U4157 (N_4157,N_3642,N_3941);
or U4158 (N_4158,N_3846,N_3816);
and U4159 (N_4159,N_3543,N_3646);
or U4160 (N_4160,N_3514,N_3910);
nor U4161 (N_4161,N_3728,N_3869);
or U4162 (N_4162,N_3973,N_3892);
nand U4163 (N_4163,N_3553,N_3804);
nand U4164 (N_4164,N_3777,N_3600);
nor U4165 (N_4165,N_3618,N_3738);
nand U4166 (N_4166,N_3964,N_3577);
and U4167 (N_4167,N_3676,N_3612);
nand U4168 (N_4168,N_3522,N_3833);
or U4169 (N_4169,N_3935,N_3589);
nand U4170 (N_4170,N_3520,N_3531);
or U4171 (N_4171,N_3551,N_3867);
and U4172 (N_4172,N_3508,N_3951);
nor U4173 (N_4173,N_3797,N_3669);
nand U4174 (N_4174,N_3909,N_3689);
nand U4175 (N_4175,N_3829,N_3679);
or U4176 (N_4176,N_3933,N_3709);
xnor U4177 (N_4177,N_3678,N_3686);
nand U4178 (N_4178,N_3673,N_3939);
xor U4179 (N_4179,N_3534,N_3977);
nor U4180 (N_4180,N_3614,N_3839);
nand U4181 (N_4181,N_3541,N_3806);
nand U4182 (N_4182,N_3828,N_3569);
nand U4183 (N_4183,N_3650,N_3515);
nor U4184 (N_4184,N_3617,N_3787);
nor U4185 (N_4185,N_3954,N_3776);
nor U4186 (N_4186,N_3960,N_3556);
nand U4187 (N_4187,N_3822,N_3758);
and U4188 (N_4188,N_3523,N_3890);
or U4189 (N_4189,N_3996,N_3851);
and U4190 (N_4190,N_3911,N_3871);
nor U4191 (N_4191,N_3740,N_3659);
and U4192 (N_4192,N_3979,N_3584);
xor U4193 (N_4193,N_3590,N_3944);
xor U4194 (N_4194,N_3847,N_3518);
and U4195 (N_4195,N_3713,N_3606);
and U4196 (N_4196,N_3799,N_3591);
nor U4197 (N_4197,N_3795,N_3571);
and U4198 (N_4198,N_3658,N_3561);
and U4199 (N_4199,N_3825,N_3546);
xor U4200 (N_4200,N_3502,N_3929);
nor U4201 (N_4201,N_3857,N_3958);
nor U4202 (N_4202,N_3533,N_3504);
and U4203 (N_4203,N_3947,N_3637);
and U4204 (N_4204,N_3545,N_3817);
nor U4205 (N_4205,N_3993,N_3901);
nor U4206 (N_4206,N_3580,N_3711);
nor U4207 (N_4207,N_3790,N_3868);
or U4208 (N_4208,N_3856,N_3952);
or U4209 (N_4209,N_3775,N_3764);
and U4210 (N_4210,N_3813,N_3959);
or U4211 (N_4211,N_3864,N_3834);
nand U4212 (N_4212,N_3763,N_3701);
xnor U4213 (N_4213,N_3920,N_3796);
nor U4214 (N_4214,N_3666,N_3801);
nand U4215 (N_4215,N_3810,N_3898);
and U4216 (N_4216,N_3623,N_3505);
and U4217 (N_4217,N_3865,N_3904);
nand U4218 (N_4218,N_3789,N_3956);
or U4219 (N_4219,N_3793,N_3818);
nand U4220 (N_4220,N_3895,N_3863);
and U4221 (N_4221,N_3886,N_3588);
or U4222 (N_4222,N_3524,N_3855);
and U4223 (N_4223,N_3682,N_3562);
xnor U4224 (N_4224,N_3955,N_3661);
and U4225 (N_4225,N_3525,N_3509);
or U4226 (N_4226,N_3988,N_3507);
nand U4227 (N_4227,N_3943,N_3918);
nand U4228 (N_4228,N_3844,N_3613);
or U4229 (N_4229,N_3995,N_3942);
nand U4230 (N_4230,N_3527,N_3982);
and U4231 (N_4231,N_3690,N_3784);
or U4232 (N_4232,N_3880,N_3537);
or U4233 (N_4233,N_3930,N_3925);
nand U4234 (N_4234,N_3708,N_3852);
and U4235 (N_4235,N_3812,N_3662);
nand U4236 (N_4236,N_3735,N_3866);
nor U4237 (N_4237,N_3723,N_3948);
xor U4238 (N_4238,N_3873,N_3608);
nor U4239 (N_4239,N_3635,N_3530);
or U4240 (N_4240,N_3626,N_3620);
nor U4241 (N_4241,N_3653,N_3602);
nor U4242 (N_4242,N_3567,N_3599);
nand U4243 (N_4243,N_3854,N_3675);
and U4244 (N_4244,N_3692,N_3950);
xor U4245 (N_4245,N_3595,N_3914);
or U4246 (N_4246,N_3685,N_3802);
and U4247 (N_4247,N_3830,N_3760);
and U4248 (N_4248,N_3976,N_3921);
and U4249 (N_4249,N_3513,N_3715);
or U4250 (N_4250,N_3572,N_3562);
nand U4251 (N_4251,N_3679,N_3794);
or U4252 (N_4252,N_3956,N_3770);
or U4253 (N_4253,N_3538,N_3642);
or U4254 (N_4254,N_3749,N_3585);
and U4255 (N_4255,N_3830,N_3536);
nand U4256 (N_4256,N_3752,N_3725);
and U4257 (N_4257,N_3562,N_3625);
and U4258 (N_4258,N_3816,N_3584);
and U4259 (N_4259,N_3909,N_3585);
nand U4260 (N_4260,N_3519,N_3547);
nand U4261 (N_4261,N_3529,N_3779);
nor U4262 (N_4262,N_3708,N_3570);
nand U4263 (N_4263,N_3615,N_3614);
and U4264 (N_4264,N_3692,N_3569);
nand U4265 (N_4265,N_3799,N_3901);
nor U4266 (N_4266,N_3690,N_3547);
nor U4267 (N_4267,N_3804,N_3890);
nand U4268 (N_4268,N_3743,N_3826);
nor U4269 (N_4269,N_3721,N_3871);
or U4270 (N_4270,N_3722,N_3745);
or U4271 (N_4271,N_3910,N_3620);
and U4272 (N_4272,N_3753,N_3925);
nand U4273 (N_4273,N_3574,N_3587);
and U4274 (N_4274,N_3989,N_3896);
or U4275 (N_4275,N_3783,N_3678);
and U4276 (N_4276,N_3781,N_3675);
and U4277 (N_4277,N_3712,N_3687);
and U4278 (N_4278,N_3834,N_3672);
nand U4279 (N_4279,N_3993,N_3561);
nor U4280 (N_4280,N_3607,N_3825);
and U4281 (N_4281,N_3985,N_3843);
and U4282 (N_4282,N_3664,N_3604);
and U4283 (N_4283,N_3572,N_3587);
and U4284 (N_4284,N_3741,N_3800);
and U4285 (N_4285,N_3828,N_3640);
nand U4286 (N_4286,N_3889,N_3955);
nor U4287 (N_4287,N_3911,N_3659);
nor U4288 (N_4288,N_3824,N_3871);
or U4289 (N_4289,N_3783,N_3775);
nor U4290 (N_4290,N_3564,N_3994);
nand U4291 (N_4291,N_3781,N_3661);
and U4292 (N_4292,N_3954,N_3643);
and U4293 (N_4293,N_3990,N_3595);
nor U4294 (N_4294,N_3724,N_3627);
and U4295 (N_4295,N_3760,N_3739);
and U4296 (N_4296,N_3580,N_3526);
nor U4297 (N_4297,N_3891,N_3804);
and U4298 (N_4298,N_3915,N_3984);
and U4299 (N_4299,N_3730,N_3866);
nor U4300 (N_4300,N_3883,N_3530);
xor U4301 (N_4301,N_3730,N_3783);
nor U4302 (N_4302,N_3938,N_3573);
nor U4303 (N_4303,N_3683,N_3981);
nand U4304 (N_4304,N_3524,N_3906);
or U4305 (N_4305,N_3914,N_3922);
or U4306 (N_4306,N_3810,N_3892);
or U4307 (N_4307,N_3683,N_3610);
nor U4308 (N_4308,N_3667,N_3955);
nor U4309 (N_4309,N_3932,N_3738);
and U4310 (N_4310,N_3658,N_3914);
nor U4311 (N_4311,N_3618,N_3810);
nor U4312 (N_4312,N_3905,N_3698);
nor U4313 (N_4313,N_3898,N_3712);
nand U4314 (N_4314,N_3611,N_3638);
and U4315 (N_4315,N_3834,N_3745);
nor U4316 (N_4316,N_3518,N_3870);
nor U4317 (N_4317,N_3871,N_3852);
or U4318 (N_4318,N_3833,N_3928);
nand U4319 (N_4319,N_3553,N_3592);
nor U4320 (N_4320,N_3869,N_3695);
and U4321 (N_4321,N_3539,N_3804);
or U4322 (N_4322,N_3777,N_3747);
or U4323 (N_4323,N_3618,N_3587);
and U4324 (N_4324,N_3580,N_3753);
nand U4325 (N_4325,N_3719,N_3655);
and U4326 (N_4326,N_3647,N_3649);
or U4327 (N_4327,N_3771,N_3755);
nand U4328 (N_4328,N_3672,N_3509);
or U4329 (N_4329,N_3907,N_3794);
nor U4330 (N_4330,N_3696,N_3644);
nand U4331 (N_4331,N_3768,N_3984);
nor U4332 (N_4332,N_3503,N_3530);
nor U4333 (N_4333,N_3833,N_3924);
nor U4334 (N_4334,N_3659,N_3748);
and U4335 (N_4335,N_3570,N_3797);
or U4336 (N_4336,N_3967,N_3620);
nor U4337 (N_4337,N_3973,N_3708);
and U4338 (N_4338,N_3781,N_3906);
nor U4339 (N_4339,N_3663,N_3807);
or U4340 (N_4340,N_3707,N_3899);
or U4341 (N_4341,N_3871,N_3710);
nor U4342 (N_4342,N_3834,N_3510);
or U4343 (N_4343,N_3603,N_3882);
nand U4344 (N_4344,N_3695,N_3553);
nand U4345 (N_4345,N_3500,N_3727);
nand U4346 (N_4346,N_3994,N_3578);
or U4347 (N_4347,N_3819,N_3764);
nor U4348 (N_4348,N_3503,N_3562);
nor U4349 (N_4349,N_3790,N_3886);
nand U4350 (N_4350,N_3546,N_3717);
nor U4351 (N_4351,N_3765,N_3543);
nand U4352 (N_4352,N_3504,N_3978);
nand U4353 (N_4353,N_3504,N_3636);
and U4354 (N_4354,N_3544,N_3891);
or U4355 (N_4355,N_3768,N_3947);
nor U4356 (N_4356,N_3617,N_3862);
or U4357 (N_4357,N_3587,N_3934);
and U4358 (N_4358,N_3971,N_3664);
xor U4359 (N_4359,N_3761,N_3982);
or U4360 (N_4360,N_3625,N_3723);
nand U4361 (N_4361,N_3978,N_3770);
and U4362 (N_4362,N_3978,N_3633);
or U4363 (N_4363,N_3891,N_3941);
and U4364 (N_4364,N_3626,N_3618);
nand U4365 (N_4365,N_3751,N_3985);
nor U4366 (N_4366,N_3826,N_3816);
nand U4367 (N_4367,N_3639,N_3809);
nor U4368 (N_4368,N_3555,N_3750);
nand U4369 (N_4369,N_3604,N_3808);
nand U4370 (N_4370,N_3549,N_3854);
nor U4371 (N_4371,N_3828,N_3938);
and U4372 (N_4372,N_3550,N_3697);
nand U4373 (N_4373,N_3664,N_3916);
or U4374 (N_4374,N_3946,N_3615);
and U4375 (N_4375,N_3918,N_3536);
and U4376 (N_4376,N_3761,N_3557);
and U4377 (N_4377,N_3832,N_3630);
and U4378 (N_4378,N_3557,N_3601);
or U4379 (N_4379,N_3840,N_3741);
and U4380 (N_4380,N_3939,N_3987);
or U4381 (N_4381,N_3594,N_3528);
nor U4382 (N_4382,N_3771,N_3994);
nand U4383 (N_4383,N_3888,N_3648);
nor U4384 (N_4384,N_3629,N_3833);
nor U4385 (N_4385,N_3683,N_3936);
or U4386 (N_4386,N_3523,N_3952);
or U4387 (N_4387,N_3632,N_3809);
nor U4388 (N_4388,N_3816,N_3680);
nand U4389 (N_4389,N_3541,N_3987);
and U4390 (N_4390,N_3650,N_3985);
and U4391 (N_4391,N_3931,N_3786);
or U4392 (N_4392,N_3910,N_3508);
nand U4393 (N_4393,N_3805,N_3593);
nand U4394 (N_4394,N_3643,N_3625);
nor U4395 (N_4395,N_3557,N_3519);
and U4396 (N_4396,N_3902,N_3851);
and U4397 (N_4397,N_3675,N_3795);
nand U4398 (N_4398,N_3754,N_3697);
and U4399 (N_4399,N_3906,N_3858);
or U4400 (N_4400,N_3635,N_3545);
and U4401 (N_4401,N_3741,N_3742);
or U4402 (N_4402,N_3659,N_3828);
and U4403 (N_4403,N_3868,N_3523);
nor U4404 (N_4404,N_3591,N_3618);
and U4405 (N_4405,N_3965,N_3818);
nor U4406 (N_4406,N_3555,N_3696);
nor U4407 (N_4407,N_3789,N_3541);
and U4408 (N_4408,N_3849,N_3780);
and U4409 (N_4409,N_3755,N_3902);
nor U4410 (N_4410,N_3518,N_3659);
and U4411 (N_4411,N_3724,N_3511);
and U4412 (N_4412,N_3865,N_3954);
nor U4413 (N_4413,N_3634,N_3685);
and U4414 (N_4414,N_3947,N_3562);
or U4415 (N_4415,N_3981,N_3810);
or U4416 (N_4416,N_3641,N_3915);
nor U4417 (N_4417,N_3906,N_3751);
nand U4418 (N_4418,N_3804,N_3823);
or U4419 (N_4419,N_3860,N_3805);
nor U4420 (N_4420,N_3734,N_3824);
nor U4421 (N_4421,N_3871,N_3534);
or U4422 (N_4422,N_3826,N_3527);
and U4423 (N_4423,N_3879,N_3701);
or U4424 (N_4424,N_3569,N_3703);
and U4425 (N_4425,N_3793,N_3567);
or U4426 (N_4426,N_3835,N_3550);
or U4427 (N_4427,N_3845,N_3713);
and U4428 (N_4428,N_3910,N_3682);
nand U4429 (N_4429,N_3516,N_3584);
nor U4430 (N_4430,N_3719,N_3720);
nand U4431 (N_4431,N_3822,N_3762);
or U4432 (N_4432,N_3555,N_3549);
nand U4433 (N_4433,N_3700,N_3532);
nor U4434 (N_4434,N_3822,N_3944);
nand U4435 (N_4435,N_3528,N_3600);
nand U4436 (N_4436,N_3615,N_3975);
nor U4437 (N_4437,N_3940,N_3623);
nand U4438 (N_4438,N_3798,N_3514);
and U4439 (N_4439,N_3895,N_3811);
or U4440 (N_4440,N_3974,N_3904);
nand U4441 (N_4441,N_3965,N_3880);
nand U4442 (N_4442,N_3772,N_3766);
and U4443 (N_4443,N_3629,N_3773);
xnor U4444 (N_4444,N_3694,N_3826);
or U4445 (N_4445,N_3683,N_3729);
and U4446 (N_4446,N_3583,N_3874);
nand U4447 (N_4447,N_3990,N_3810);
or U4448 (N_4448,N_3997,N_3889);
and U4449 (N_4449,N_3574,N_3923);
and U4450 (N_4450,N_3940,N_3538);
nor U4451 (N_4451,N_3547,N_3717);
nand U4452 (N_4452,N_3572,N_3776);
nor U4453 (N_4453,N_3723,N_3813);
nand U4454 (N_4454,N_3786,N_3929);
nand U4455 (N_4455,N_3768,N_3959);
and U4456 (N_4456,N_3945,N_3835);
or U4457 (N_4457,N_3554,N_3939);
or U4458 (N_4458,N_3592,N_3507);
or U4459 (N_4459,N_3552,N_3754);
nand U4460 (N_4460,N_3660,N_3941);
and U4461 (N_4461,N_3978,N_3914);
nand U4462 (N_4462,N_3679,N_3907);
or U4463 (N_4463,N_3566,N_3650);
and U4464 (N_4464,N_3699,N_3949);
nor U4465 (N_4465,N_3824,N_3919);
and U4466 (N_4466,N_3624,N_3564);
or U4467 (N_4467,N_3513,N_3994);
and U4468 (N_4468,N_3623,N_3905);
and U4469 (N_4469,N_3975,N_3692);
nor U4470 (N_4470,N_3635,N_3938);
nand U4471 (N_4471,N_3964,N_3943);
or U4472 (N_4472,N_3502,N_3715);
nor U4473 (N_4473,N_3925,N_3657);
nand U4474 (N_4474,N_3938,N_3887);
nand U4475 (N_4475,N_3534,N_3695);
or U4476 (N_4476,N_3531,N_3724);
nand U4477 (N_4477,N_3735,N_3548);
or U4478 (N_4478,N_3783,N_3514);
or U4479 (N_4479,N_3525,N_3548);
nand U4480 (N_4480,N_3704,N_3630);
and U4481 (N_4481,N_3747,N_3871);
or U4482 (N_4482,N_3940,N_3542);
nor U4483 (N_4483,N_3622,N_3892);
and U4484 (N_4484,N_3638,N_3912);
or U4485 (N_4485,N_3703,N_3927);
xor U4486 (N_4486,N_3818,N_3877);
xnor U4487 (N_4487,N_3518,N_3866);
nand U4488 (N_4488,N_3878,N_3716);
nand U4489 (N_4489,N_3608,N_3511);
and U4490 (N_4490,N_3940,N_3798);
nor U4491 (N_4491,N_3808,N_3617);
xor U4492 (N_4492,N_3581,N_3997);
nand U4493 (N_4493,N_3866,N_3939);
or U4494 (N_4494,N_3773,N_3929);
and U4495 (N_4495,N_3808,N_3880);
and U4496 (N_4496,N_3700,N_3621);
or U4497 (N_4497,N_3819,N_3533);
or U4498 (N_4498,N_3610,N_3746);
or U4499 (N_4499,N_3773,N_3987);
xnor U4500 (N_4500,N_4161,N_4188);
or U4501 (N_4501,N_4211,N_4220);
nand U4502 (N_4502,N_4190,N_4359);
and U4503 (N_4503,N_4287,N_4465);
and U4504 (N_4504,N_4295,N_4327);
and U4505 (N_4505,N_4145,N_4095);
or U4506 (N_4506,N_4444,N_4456);
or U4507 (N_4507,N_4490,N_4072);
nand U4508 (N_4508,N_4343,N_4322);
nor U4509 (N_4509,N_4329,N_4044);
nor U4510 (N_4510,N_4158,N_4280);
nand U4511 (N_4511,N_4411,N_4470);
or U4512 (N_4512,N_4149,N_4071);
nand U4513 (N_4513,N_4417,N_4455);
and U4514 (N_4514,N_4132,N_4251);
nor U4515 (N_4515,N_4139,N_4283);
nor U4516 (N_4516,N_4005,N_4457);
nor U4517 (N_4517,N_4438,N_4334);
nand U4518 (N_4518,N_4309,N_4213);
nand U4519 (N_4519,N_4227,N_4113);
or U4520 (N_4520,N_4405,N_4195);
nand U4521 (N_4521,N_4377,N_4066);
nor U4522 (N_4522,N_4437,N_4200);
nor U4523 (N_4523,N_4410,N_4221);
or U4524 (N_4524,N_4019,N_4086);
and U4525 (N_4525,N_4033,N_4125);
nand U4526 (N_4526,N_4319,N_4469);
nand U4527 (N_4527,N_4431,N_4089);
or U4528 (N_4528,N_4124,N_4349);
nand U4529 (N_4529,N_4351,N_4433);
or U4530 (N_4530,N_4244,N_4320);
nor U4531 (N_4531,N_4300,N_4021);
nand U4532 (N_4532,N_4385,N_4478);
or U4533 (N_4533,N_4013,N_4263);
or U4534 (N_4534,N_4228,N_4306);
nor U4535 (N_4535,N_4069,N_4084);
nor U4536 (N_4536,N_4142,N_4192);
nand U4537 (N_4537,N_4129,N_4153);
and U4538 (N_4538,N_4184,N_4157);
nor U4539 (N_4539,N_4097,N_4464);
nor U4540 (N_4540,N_4474,N_4141);
and U4541 (N_4541,N_4079,N_4046);
nor U4542 (N_4542,N_4240,N_4102);
nor U4543 (N_4543,N_4103,N_4290);
or U4544 (N_4544,N_4302,N_4399);
or U4545 (N_4545,N_4321,N_4460);
xor U4546 (N_4546,N_4494,N_4182);
or U4547 (N_4547,N_4432,N_4077);
nand U4548 (N_4548,N_4006,N_4270);
nand U4549 (N_4549,N_4488,N_4011);
nor U4550 (N_4550,N_4056,N_4483);
nor U4551 (N_4551,N_4029,N_4247);
nand U4552 (N_4552,N_4216,N_4369);
and U4553 (N_4553,N_4229,N_4219);
and U4554 (N_4554,N_4037,N_4232);
and U4555 (N_4555,N_4144,N_4259);
nor U4556 (N_4556,N_4186,N_4026);
nand U4557 (N_4557,N_4067,N_4471);
nand U4558 (N_4558,N_4344,N_4206);
and U4559 (N_4559,N_4212,N_4246);
or U4560 (N_4560,N_4180,N_4271);
nor U4561 (N_4561,N_4418,N_4168);
or U4562 (N_4562,N_4191,N_4355);
and U4563 (N_4563,N_4307,N_4045);
nand U4564 (N_4564,N_4374,N_4185);
nand U4565 (N_4565,N_4123,N_4285);
nand U4566 (N_4566,N_4496,N_4367);
or U4567 (N_4567,N_4250,N_4256);
nor U4568 (N_4568,N_4238,N_4394);
nand U4569 (N_4569,N_4426,N_4252);
nand U4570 (N_4570,N_4092,N_4378);
nand U4571 (N_4571,N_4382,N_4371);
or U4572 (N_4572,N_4203,N_4181);
or U4573 (N_4573,N_4023,N_4274);
or U4574 (N_4574,N_4040,N_4201);
nor U4575 (N_4575,N_4434,N_4160);
nor U4576 (N_4576,N_4311,N_4315);
xor U4577 (N_4577,N_4347,N_4118);
or U4578 (N_4578,N_4324,N_4204);
nor U4579 (N_4579,N_4172,N_4094);
and U4580 (N_4580,N_4392,N_4435);
nor U4581 (N_4581,N_4004,N_4083);
nand U4582 (N_4582,N_4202,N_4273);
and U4583 (N_4583,N_4038,N_4208);
nand U4584 (N_4584,N_4258,N_4062);
xor U4585 (N_4585,N_4098,N_4128);
nand U4586 (N_4586,N_4171,N_4379);
and U4587 (N_4587,N_4467,N_4049);
and U4588 (N_4588,N_4462,N_4177);
or U4589 (N_4589,N_4364,N_4108);
or U4590 (N_4590,N_4454,N_4105);
nor U4591 (N_4591,N_4458,N_4050);
nor U4592 (N_4592,N_4299,N_4368);
nand U4593 (N_4593,N_4116,N_4015);
and U4594 (N_4594,N_4391,N_4179);
nand U4595 (N_4595,N_4131,N_4441);
and U4596 (N_4596,N_4337,N_4073);
and U4597 (N_4597,N_4257,N_4032);
or U4598 (N_4598,N_4439,N_4042);
or U4599 (N_4599,N_4120,N_4249);
nor U4600 (N_4600,N_4130,N_4241);
nand U4601 (N_4601,N_4027,N_4115);
nand U4602 (N_4602,N_4277,N_4022);
or U4603 (N_4603,N_4284,N_4057);
nor U4604 (N_4604,N_4197,N_4370);
nand U4605 (N_4605,N_4112,N_4384);
nor U4606 (N_4606,N_4296,N_4024);
or U4607 (N_4607,N_4366,N_4225);
nand U4608 (N_4608,N_4492,N_4036);
xnor U4609 (N_4609,N_4375,N_4233);
nor U4610 (N_4610,N_4498,N_4140);
and U4611 (N_4611,N_4301,N_4253);
and U4612 (N_4612,N_4152,N_4354);
and U4613 (N_4613,N_4065,N_4396);
nand U4614 (N_4614,N_4305,N_4356);
nor U4615 (N_4615,N_4348,N_4169);
nor U4616 (N_4616,N_4331,N_4101);
and U4617 (N_4617,N_4261,N_4122);
nor U4618 (N_4618,N_4215,N_4167);
and U4619 (N_4619,N_4291,N_4034);
nand U4620 (N_4620,N_4265,N_4147);
nor U4621 (N_4621,N_4443,N_4173);
nand U4622 (N_4622,N_4262,N_4237);
or U4623 (N_4623,N_4310,N_4199);
or U4624 (N_4624,N_4318,N_4163);
nor U4625 (N_4625,N_4423,N_4289);
and U4626 (N_4626,N_4166,N_4001);
xor U4627 (N_4627,N_4081,N_4292);
or U4628 (N_4628,N_4205,N_4484);
and U4629 (N_4629,N_4093,N_4020);
or U4630 (N_4630,N_4217,N_4395);
nor U4631 (N_4631,N_4119,N_4352);
nand U4632 (N_4632,N_4126,N_4111);
nor U4633 (N_4633,N_4298,N_4209);
or U4634 (N_4634,N_4075,N_4014);
and U4635 (N_4635,N_4170,N_4178);
and U4636 (N_4636,N_4175,N_4468);
nand U4637 (N_4637,N_4150,N_4332);
nand U4638 (N_4638,N_4475,N_4107);
or U4639 (N_4639,N_4148,N_4387);
or U4640 (N_4640,N_4245,N_4063);
or U4641 (N_4641,N_4018,N_4031);
nand U4642 (N_4642,N_4419,N_4421);
nor U4643 (N_4643,N_4282,N_4198);
and U4644 (N_4644,N_4279,N_4012);
or U4645 (N_4645,N_4407,N_4362);
nor U4646 (N_4646,N_4002,N_4060);
and U4647 (N_4647,N_4146,N_4424);
nor U4648 (N_4648,N_4008,N_4183);
and U4649 (N_4649,N_4480,N_4372);
or U4650 (N_4650,N_4409,N_4380);
or U4651 (N_4651,N_4390,N_4239);
nor U4652 (N_4652,N_4493,N_4472);
nor U4653 (N_4653,N_4448,N_4236);
or U4654 (N_4654,N_4230,N_4269);
nand U4655 (N_4655,N_4064,N_4078);
or U4656 (N_4656,N_4223,N_4009);
xor U4657 (N_4657,N_4497,N_4422);
xnor U4658 (N_4658,N_4412,N_4449);
nor U4659 (N_4659,N_4193,N_4428);
nand U4660 (N_4660,N_4400,N_4248);
nor U4661 (N_4661,N_4117,N_4174);
xnor U4662 (N_4662,N_4286,N_4333);
or U4663 (N_4663,N_4313,N_4453);
xnor U4664 (N_4664,N_4138,N_4459);
or U4665 (N_4665,N_4135,N_4254);
nand U4666 (N_4666,N_4342,N_4415);
or U4667 (N_4667,N_4187,N_4485);
and U4668 (N_4668,N_4275,N_4447);
xor U4669 (N_4669,N_4137,N_4427);
and U4670 (N_4670,N_4341,N_4133);
or U4671 (N_4671,N_4430,N_4099);
xor U4672 (N_4672,N_4070,N_4406);
nand U4673 (N_4673,N_4226,N_4136);
or U4674 (N_4674,N_4486,N_4068);
nor U4675 (N_4675,N_4028,N_4127);
and U4676 (N_4676,N_4267,N_4058);
and U4677 (N_4677,N_4055,N_4312);
xor U4678 (N_4678,N_4473,N_4260);
nor U4679 (N_4679,N_4121,N_4477);
nor U4680 (N_4680,N_4463,N_4461);
nor U4681 (N_4681,N_4231,N_4340);
or U4682 (N_4682,N_4491,N_4451);
nor U4683 (N_4683,N_4440,N_4466);
and U4684 (N_4684,N_4100,N_4048);
nand U4685 (N_4685,N_4082,N_4338);
nor U4686 (N_4686,N_4039,N_4294);
nor U4687 (N_4687,N_4090,N_4242);
nand U4688 (N_4688,N_4363,N_4350);
or U4689 (N_4689,N_4425,N_4266);
xnor U4690 (N_4690,N_4030,N_4268);
or U4691 (N_4691,N_4047,N_4194);
nand U4692 (N_4692,N_4328,N_4281);
nand U4693 (N_4693,N_4104,N_4151);
or U4694 (N_4694,N_4293,N_4189);
and U4695 (N_4695,N_4288,N_4304);
and U4696 (N_4696,N_4376,N_4154);
nor U4697 (N_4697,N_4143,N_4303);
nor U4698 (N_4698,N_4074,N_4389);
nand U4699 (N_4699,N_4016,N_4445);
or U4700 (N_4700,N_4420,N_4017);
and U4701 (N_4701,N_4162,N_4397);
xnor U4702 (N_4702,N_4041,N_4487);
xor U4703 (N_4703,N_4235,N_4080);
nand U4704 (N_4704,N_4276,N_4076);
or U4705 (N_4705,N_4383,N_4159);
or U4706 (N_4706,N_4361,N_4059);
nor U4707 (N_4707,N_4388,N_4164);
and U4708 (N_4708,N_4446,N_4413);
nand U4709 (N_4709,N_4155,N_4043);
or U4710 (N_4710,N_4243,N_4007);
nor U4711 (N_4711,N_4401,N_4035);
nor U4712 (N_4712,N_4326,N_4404);
nor U4713 (N_4713,N_4398,N_4323);
nand U4714 (N_4714,N_4345,N_4381);
and U4715 (N_4715,N_4365,N_4450);
or U4716 (N_4716,N_4234,N_4357);
and U4717 (N_4717,N_4335,N_4317);
nand U4718 (N_4718,N_4414,N_4481);
nor U4719 (N_4719,N_4436,N_4106);
or U4720 (N_4720,N_4114,N_4051);
nor U4721 (N_4721,N_4207,N_4091);
nor U4722 (N_4722,N_4429,N_4386);
nor U4723 (N_4723,N_4053,N_4316);
nor U4724 (N_4724,N_4087,N_4134);
nor U4725 (N_4725,N_4339,N_4489);
or U4726 (N_4726,N_4416,N_4109);
and U4727 (N_4727,N_4442,N_4308);
nor U4728 (N_4728,N_4297,N_4222);
nor U4729 (N_4729,N_4408,N_4346);
nand U4730 (N_4730,N_4482,N_4360);
nor U4731 (N_4731,N_4499,N_4061);
and U4732 (N_4732,N_4176,N_4224);
nand U4733 (N_4733,N_4264,N_4452);
nand U4734 (N_4734,N_4476,N_4403);
xor U4735 (N_4735,N_4393,N_4054);
nor U4736 (N_4736,N_4353,N_4000);
or U4737 (N_4737,N_4085,N_4255);
nor U4738 (N_4738,N_4010,N_4025);
or U4739 (N_4739,N_4214,N_4003);
or U4740 (N_4740,N_4052,N_4272);
nand U4741 (N_4741,N_4165,N_4196);
and U4742 (N_4742,N_4358,N_4088);
nor U4743 (N_4743,N_4278,N_4314);
or U4744 (N_4744,N_4218,N_4495);
xnor U4745 (N_4745,N_4325,N_4096);
nor U4746 (N_4746,N_4479,N_4402);
nand U4747 (N_4747,N_4330,N_4336);
and U4748 (N_4748,N_4156,N_4210);
and U4749 (N_4749,N_4373,N_4110);
nand U4750 (N_4750,N_4020,N_4462);
or U4751 (N_4751,N_4385,N_4228);
nand U4752 (N_4752,N_4498,N_4342);
nor U4753 (N_4753,N_4451,N_4191);
nor U4754 (N_4754,N_4249,N_4264);
or U4755 (N_4755,N_4485,N_4307);
and U4756 (N_4756,N_4266,N_4312);
nand U4757 (N_4757,N_4171,N_4237);
or U4758 (N_4758,N_4127,N_4264);
nor U4759 (N_4759,N_4315,N_4237);
nor U4760 (N_4760,N_4415,N_4289);
nand U4761 (N_4761,N_4118,N_4093);
and U4762 (N_4762,N_4316,N_4471);
or U4763 (N_4763,N_4491,N_4409);
or U4764 (N_4764,N_4275,N_4092);
nand U4765 (N_4765,N_4043,N_4014);
nor U4766 (N_4766,N_4258,N_4227);
nor U4767 (N_4767,N_4056,N_4198);
and U4768 (N_4768,N_4282,N_4476);
or U4769 (N_4769,N_4272,N_4349);
xor U4770 (N_4770,N_4032,N_4273);
nand U4771 (N_4771,N_4040,N_4179);
nand U4772 (N_4772,N_4411,N_4021);
xnor U4773 (N_4773,N_4459,N_4126);
nor U4774 (N_4774,N_4243,N_4324);
nor U4775 (N_4775,N_4145,N_4329);
nor U4776 (N_4776,N_4301,N_4262);
nor U4777 (N_4777,N_4457,N_4248);
nand U4778 (N_4778,N_4453,N_4042);
and U4779 (N_4779,N_4379,N_4465);
nand U4780 (N_4780,N_4108,N_4425);
and U4781 (N_4781,N_4420,N_4412);
nor U4782 (N_4782,N_4121,N_4219);
or U4783 (N_4783,N_4028,N_4306);
nor U4784 (N_4784,N_4425,N_4194);
and U4785 (N_4785,N_4148,N_4131);
and U4786 (N_4786,N_4334,N_4281);
nand U4787 (N_4787,N_4397,N_4245);
or U4788 (N_4788,N_4070,N_4397);
or U4789 (N_4789,N_4047,N_4293);
xnor U4790 (N_4790,N_4433,N_4317);
nor U4791 (N_4791,N_4269,N_4363);
nor U4792 (N_4792,N_4480,N_4431);
nor U4793 (N_4793,N_4492,N_4008);
and U4794 (N_4794,N_4205,N_4159);
nand U4795 (N_4795,N_4377,N_4097);
or U4796 (N_4796,N_4108,N_4433);
xnor U4797 (N_4797,N_4390,N_4323);
nand U4798 (N_4798,N_4083,N_4111);
nand U4799 (N_4799,N_4318,N_4491);
nor U4800 (N_4800,N_4435,N_4183);
nor U4801 (N_4801,N_4105,N_4269);
or U4802 (N_4802,N_4003,N_4192);
and U4803 (N_4803,N_4063,N_4167);
and U4804 (N_4804,N_4327,N_4416);
and U4805 (N_4805,N_4425,N_4476);
nor U4806 (N_4806,N_4272,N_4190);
and U4807 (N_4807,N_4457,N_4355);
nand U4808 (N_4808,N_4049,N_4218);
nand U4809 (N_4809,N_4499,N_4161);
nand U4810 (N_4810,N_4336,N_4094);
and U4811 (N_4811,N_4004,N_4155);
and U4812 (N_4812,N_4289,N_4368);
nor U4813 (N_4813,N_4328,N_4357);
or U4814 (N_4814,N_4116,N_4278);
nor U4815 (N_4815,N_4468,N_4199);
nand U4816 (N_4816,N_4319,N_4375);
or U4817 (N_4817,N_4228,N_4324);
nand U4818 (N_4818,N_4202,N_4220);
nor U4819 (N_4819,N_4020,N_4173);
nand U4820 (N_4820,N_4023,N_4497);
or U4821 (N_4821,N_4314,N_4232);
or U4822 (N_4822,N_4362,N_4081);
nand U4823 (N_4823,N_4382,N_4315);
and U4824 (N_4824,N_4291,N_4053);
and U4825 (N_4825,N_4123,N_4463);
nand U4826 (N_4826,N_4278,N_4186);
and U4827 (N_4827,N_4286,N_4308);
nand U4828 (N_4828,N_4163,N_4150);
or U4829 (N_4829,N_4278,N_4177);
or U4830 (N_4830,N_4099,N_4086);
or U4831 (N_4831,N_4127,N_4013);
nor U4832 (N_4832,N_4181,N_4401);
nor U4833 (N_4833,N_4325,N_4393);
and U4834 (N_4834,N_4105,N_4064);
nand U4835 (N_4835,N_4339,N_4225);
nor U4836 (N_4836,N_4032,N_4216);
or U4837 (N_4837,N_4154,N_4187);
or U4838 (N_4838,N_4463,N_4230);
and U4839 (N_4839,N_4437,N_4142);
nor U4840 (N_4840,N_4142,N_4148);
and U4841 (N_4841,N_4254,N_4117);
nand U4842 (N_4842,N_4224,N_4423);
or U4843 (N_4843,N_4004,N_4469);
and U4844 (N_4844,N_4491,N_4478);
or U4845 (N_4845,N_4157,N_4244);
nor U4846 (N_4846,N_4170,N_4272);
and U4847 (N_4847,N_4204,N_4168);
or U4848 (N_4848,N_4117,N_4372);
nor U4849 (N_4849,N_4163,N_4436);
nor U4850 (N_4850,N_4285,N_4299);
nand U4851 (N_4851,N_4415,N_4388);
nor U4852 (N_4852,N_4379,N_4083);
nor U4853 (N_4853,N_4181,N_4327);
nand U4854 (N_4854,N_4272,N_4463);
nand U4855 (N_4855,N_4232,N_4254);
nand U4856 (N_4856,N_4036,N_4073);
nand U4857 (N_4857,N_4476,N_4351);
or U4858 (N_4858,N_4455,N_4097);
nand U4859 (N_4859,N_4010,N_4499);
and U4860 (N_4860,N_4308,N_4496);
and U4861 (N_4861,N_4370,N_4499);
nand U4862 (N_4862,N_4264,N_4332);
and U4863 (N_4863,N_4302,N_4467);
or U4864 (N_4864,N_4304,N_4494);
nor U4865 (N_4865,N_4483,N_4491);
or U4866 (N_4866,N_4147,N_4054);
and U4867 (N_4867,N_4118,N_4279);
nor U4868 (N_4868,N_4250,N_4193);
nand U4869 (N_4869,N_4144,N_4322);
or U4870 (N_4870,N_4438,N_4073);
nand U4871 (N_4871,N_4016,N_4177);
and U4872 (N_4872,N_4026,N_4426);
nor U4873 (N_4873,N_4349,N_4433);
or U4874 (N_4874,N_4201,N_4391);
nor U4875 (N_4875,N_4226,N_4200);
and U4876 (N_4876,N_4137,N_4338);
nand U4877 (N_4877,N_4287,N_4388);
and U4878 (N_4878,N_4327,N_4076);
nor U4879 (N_4879,N_4066,N_4075);
and U4880 (N_4880,N_4279,N_4410);
nor U4881 (N_4881,N_4386,N_4210);
or U4882 (N_4882,N_4239,N_4398);
or U4883 (N_4883,N_4092,N_4023);
nand U4884 (N_4884,N_4371,N_4112);
and U4885 (N_4885,N_4364,N_4334);
nand U4886 (N_4886,N_4220,N_4198);
nor U4887 (N_4887,N_4170,N_4129);
nor U4888 (N_4888,N_4294,N_4023);
or U4889 (N_4889,N_4369,N_4176);
or U4890 (N_4890,N_4060,N_4280);
and U4891 (N_4891,N_4103,N_4413);
xnor U4892 (N_4892,N_4415,N_4069);
nor U4893 (N_4893,N_4436,N_4321);
and U4894 (N_4894,N_4064,N_4461);
nor U4895 (N_4895,N_4026,N_4463);
nor U4896 (N_4896,N_4423,N_4170);
nand U4897 (N_4897,N_4008,N_4349);
nor U4898 (N_4898,N_4247,N_4300);
or U4899 (N_4899,N_4236,N_4110);
nor U4900 (N_4900,N_4123,N_4335);
nor U4901 (N_4901,N_4422,N_4306);
and U4902 (N_4902,N_4428,N_4094);
and U4903 (N_4903,N_4422,N_4322);
xor U4904 (N_4904,N_4385,N_4017);
nand U4905 (N_4905,N_4197,N_4424);
nand U4906 (N_4906,N_4195,N_4129);
or U4907 (N_4907,N_4080,N_4019);
nor U4908 (N_4908,N_4488,N_4368);
xor U4909 (N_4909,N_4226,N_4107);
or U4910 (N_4910,N_4468,N_4266);
nor U4911 (N_4911,N_4180,N_4493);
and U4912 (N_4912,N_4140,N_4480);
nor U4913 (N_4913,N_4054,N_4279);
and U4914 (N_4914,N_4368,N_4029);
xnor U4915 (N_4915,N_4076,N_4073);
or U4916 (N_4916,N_4086,N_4246);
nand U4917 (N_4917,N_4285,N_4272);
or U4918 (N_4918,N_4487,N_4085);
nor U4919 (N_4919,N_4291,N_4115);
and U4920 (N_4920,N_4038,N_4336);
or U4921 (N_4921,N_4211,N_4454);
nand U4922 (N_4922,N_4108,N_4267);
nand U4923 (N_4923,N_4033,N_4061);
nor U4924 (N_4924,N_4279,N_4222);
or U4925 (N_4925,N_4192,N_4162);
and U4926 (N_4926,N_4280,N_4001);
nor U4927 (N_4927,N_4145,N_4416);
and U4928 (N_4928,N_4053,N_4385);
nand U4929 (N_4929,N_4386,N_4026);
nand U4930 (N_4930,N_4409,N_4458);
xor U4931 (N_4931,N_4491,N_4022);
and U4932 (N_4932,N_4284,N_4409);
and U4933 (N_4933,N_4425,N_4492);
and U4934 (N_4934,N_4213,N_4409);
nor U4935 (N_4935,N_4226,N_4150);
nor U4936 (N_4936,N_4054,N_4390);
or U4937 (N_4937,N_4172,N_4370);
nor U4938 (N_4938,N_4035,N_4365);
nor U4939 (N_4939,N_4251,N_4487);
and U4940 (N_4940,N_4328,N_4331);
nand U4941 (N_4941,N_4315,N_4434);
nor U4942 (N_4942,N_4077,N_4448);
nand U4943 (N_4943,N_4448,N_4129);
xor U4944 (N_4944,N_4105,N_4179);
or U4945 (N_4945,N_4331,N_4168);
xor U4946 (N_4946,N_4138,N_4173);
nand U4947 (N_4947,N_4465,N_4112);
and U4948 (N_4948,N_4348,N_4016);
or U4949 (N_4949,N_4403,N_4295);
nor U4950 (N_4950,N_4197,N_4348);
or U4951 (N_4951,N_4425,N_4348);
and U4952 (N_4952,N_4082,N_4031);
nand U4953 (N_4953,N_4187,N_4020);
nor U4954 (N_4954,N_4291,N_4347);
nand U4955 (N_4955,N_4056,N_4464);
nand U4956 (N_4956,N_4033,N_4370);
nand U4957 (N_4957,N_4183,N_4089);
and U4958 (N_4958,N_4079,N_4145);
xor U4959 (N_4959,N_4183,N_4095);
nor U4960 (N_4960,N_4107,N_4232);
nor U4961 (N_4961,N_4057,N_4311);
nand U4962 (N_4962,N_4429,N_4348);
nand U4963 (N_4963,N_4121,N_4243);
nand U4964 (N_4964,N_4418,N_4449);
nand U4965 (N_4965,N_4481,N_4324);
and U4966 (N_4966,N_4270,N_4016);
nor U4967 (N_4967,N_4281,N_4174);
and U4968 (N_4968,N_4363,N_4088);
or U4969 (N_4969,N_4046,N_4367);
or U4970 (N_4970,N_4123,N_4035);
or U4971 (N_4971,N_4349,N_4464);
or U4972 (N_4972,N_4427,N_4240);
or U4973 (N_4973,N_4056,N_4279);
nor U4974 (N_4974,N_4311,N_4005);
and U4975 (N_4975,N_4237,N_4212);
or U4976 (N_4976,N_4230,N_4290);
or U4977 (N_4977,N_4039,N_4432);
nand U4978 (N_4978,N_4119,N_4156);
nor U4979 (N_4979,N_4049,N_4321);
nor U4980 (N_4980,N_4173,N_4456);
or U4981 (N_4981,N_4000,N_4250);
nand U4982 (N_4982,N_4090,N_4141);
or U4983 (N_4983,N_4388,N_4031);
nand U4984 (N_4984,N_4151,N_4285);
xor U4985 (N_4985,N_4178,N_4251);
or U4986 (N_4986,N_4136,N_4456);
nand U4987 (N_4987,N_4496,N_4414);
or U4988 (N_4988,N_4413,N_4484);
or U4989 (N_4989,N_4240,N_4266);
nand U4990 (N_4990,N_4340,N_4263);
nor U4991 (N_4991,N_4169,N_4444);
nor U4992 (N_4992,N_4289,N_4202);
nand U4993 (N_4993,N_4191,N_4077);
and U4994 (N_4994,N_4263,N_4249);
nand U4995 (N_4995,N_4003,N_4327);
nand U4996 (N_4996,N_4312,N_4434);
xor U4997 (N_4997,N_4326,N_4120);
and U4998 (N_4998,N_4366,N_4272);
and U4999 (N_4999,N_4394,N_4105);
or UO_0 (O_0,N_4957,N_4937);
nor UO_1 (O_1,N_4572,N_4557);
nor UO_2 (O_2,N_4641,N_4853);
nor UO_3 (O_3,N_4769,N_4516);
nand UO_4 (O_4,N_4560,N_4526);
or UO_5 (O_5,N_4571,N_4966);
nand UO_6 (O_6,N_4562,N_4776);
or UO_7 (O_7,N_4553,N_4955);
and UO_8 (O_8,N_4511,N_4952);
or UO_9 (O_9,N_4594,N_4991);
nand UO_10 (O_10,N_4900,N_4944);
or UO_11 (O_11,N_4634,N_4984);
nand UO_12 (O_12,N_4884,N_4743);
or UO_13 (O_13,N_4783,N_4994);
and UO_14 (O_14,N_4896,N_4842);
and UO_15 (O_15,N_4576,N_4950);
nor UO_16 (O_16,N_4518,N_4872);
and UO_17 (O_17,N_4792,N_4870);
and UO_18 (O_18,N_4917,N_4764);
and UO_19 (O_19,N_4649,N_4927);
nor UO_20 (O_20,N_4628,N_4617);
or UO_21 (O_21,N_4928,N_4715);
xor UO_22 (O_22,N_4780,N_4808);
and UO_23 (O_23,N_4901,N_4602);
or UO_24 (O_24,N_4903,N_4814);
or UO_25 (O_25,N_4573,N_4710);
or UO_26 (O_26,N_4721,N_4926);
xor UO_27 (O_27,N_4567,N_4822);
nor UO_28 (O_28,N_4754,N_4677);
or UO_29 (O_29,N_4569,N_4890);
nand UO_30 (O_30,N_4804,N_4757);
and UO_31 (O_31,N_4575,N_4534);
nand UO_32 (O_32,N_4606,N_4510);
nor UO_33 (O_33,N_4585,N_4861);
or UO_34 (O_34,N_4623,N_4902);
nor UO_35 (O_35,N_4529,N_4865);
and UO_36 (O_36,N_4707,N_4543);
and UO_37 (O_37,N_4748,N_4753);
nand UO_38 (O_38,N_4687,N_4979);
or UO_39 (O_39,N_4733,N_4940);
nor UO_40 (O_40,N_4741,N_4895);
nor UO_41 (O_41,N_4811,N_4997);
nand UO_42 (O_42,N_4660,N_4790);
or UO_43 (O_43,N_4506,N_4770);
nand UO_44 (O_44,N_4666,N_4988);
or UO_45 (O_45,N_4761,N_4507);
and UO_46 (O_46,N_4815,N_4859);
nor UO_47 (O_47,N_4751,N_4750);
nand UO_48 (O_48,N_4945,N_4542);
nor UO_49 (O_49,N_4604,N_4845);
nand UO_50 (O_50,N_4868,N_4973);
or UO_51 (O_51,N_4911,N_4637);
nor UO_52 (O_52,N_4893,N_4722);
nand UO_53 (O_53,N_4598,N_4786);
nor UO_54 (O_54,N_4942,N_4580);
or UO_55 (O_55,N_4836,N_4877);
or UO_56 (O_56,N_4558,N_4514);
or UO_57 (O_57,N_4925,N_4974);
nor UO_58 (O_58,N_4656,N_4930);
nand UO_59 (O_59,N_4712,N_4866);
and UO_60 (O_60,N_4760,N_4679);
or UO_61 (O_61,N_4638,N_4839);
nand UO_62 (O_62,N_4883,N_4589);
or UO_63 (O_63,N_4972,N_4517);
or UO_64 (O_64,N_4527,N_4934);
or UO_65 (O_65,N_4608,N_4881);
or UO_66 (O_66,N_4744,N_4501);
and UO_67 (O_67,N_4696,N_4626);
and UO_68 (O_68,N_4995,N_4746);
or UO_69 (O_69,N_4657,N_4912);
or UO_70 (O_70,N_4844,N_4662);
nor UO_71 (O_71,N_4971,N_4676);
nand UO_72 (O_72,N_4673,N_4904);
and UO_73 (O_73,N_4788,N_4913);
nor UO_74 (O_74,N_4989,N_4880);
or UO_75 (O_75,N_4919,N_4600);
or UO_76 (O_76,N_4803,N_4668);
nor UO_77 (O_77,N_4702,N_4898);
nand UO_78 (O_78,N_4782,N_4785);
nor UO_79 (O_79,N_4923,N_4706);
nand UO_80 (O_80,N_4867,N_4593);
nor UO_81 (O_81,N_4767,N_4716);
and UO_82 (O_82,N_4834,N_4664);
nor UO_83 (O_83,N_4752,N_4559);
and UO_84 (O_84,N_4652,N_4835);
and UO_85 (O_85,N_4536,N_4658);
or UO_86 (O_86,N_4990,N_4591);
or UO_87 (O_87,N_4946,N_4871);
and UO_88 (O_88,N_4789,N_4694);
nand UO_89 (O_89,N_4779,N_4690);
and UO_90 (O_90,N_4964,N_4539);
nor UO_91 (O_91,N_4695,N_4530);
and UO_92 (O_92,N_4661,N_4654);
or UO_93 (O_93,N_4680,N_4519);
and UO_94 (O_94,N_4978,N_4907);
or UO_95 (O_95,N_4833,N_4813);
or UO_96 (O_96,N_4967,N_4947);
nor UO_97 (O_97,N_4635,N_4705);
nor UO_98 (O_98,N_4728,N_4650);
and UO_99 (O_99,N_4711,N_4618);
nor UO_100 (O_100,N_4578,N_4920);
or UO_101 (O_101,N_4772,N_4686);
xor UO_102 (O_102,N_4693,N_4985);
nor UO_103 (O_103,N_4681,N_4851);
nor UO_104 (O_104,N_4932,N_4855);
or UO_105 (O_105,N_4675,N_4943);
nor UO_106 (O_106,N_4546,N_4682);
and UO_107 (O_107,N_4781,N_4731);
and UO_108 (O_108,N_4791,N_4667);
nor UO_109 (O_109,N_4563,N_4975);
or UO_110 (O_110,N_4931,N_4500);
or UO_111 (O_111,N_4503,N_4936);
or UO_112 (O_112,N_4819,N_4512);
nand UO_113 (O_113,N_4535,N_4799);
nand UO_114 (O_114,N_4784,N_4581);
and UO_115 (O_115,N_4631,N_4802);
or UO_116 (O_116,N_4605,N_4688);
xnor UO_117 (O_117,N_4611,N_4863);
or UO_118 (O_118,N_4929,N_4840);
nand UO_119 (O_119,N_4899,N_4875);
and UO_120 (O_120,N_4889,N_4999);
nor UO_121 (O_121,N_4810,N_4981);
nand UO_122 (O_122,N_4939,N_4771);
nor UO_123 (O_123,N_4807,N_4620);
nand UO_124 (O_124,N_4905,N_4524);
and UO_125 (O_125,N_4998,N_4763);
nor UO_126 (O_126,N_4601,N_4787);
nand UO_127 (O_127,N_4847,N_4607);
and UO_128 (O_128,N_4831,N_4798);
or UO_129 (O_129,N_4592,N_4579);
nor UO_130 (O_130,N_4885,N_4565);
nand UO_131 (O_131,N_4888,N_4574);
xnor UO_132 (O_132,N_4713,N_4672);
and UO_133 (O_133,N_4832,N_4795);
nand UO_134 (O_134,N_4909,N_4726);
and UO_135 (O_135,N_4980,N_4806);
nand UO_136 (O_136,N_4671,N_4830);
or UO_137 (O_137,N_4699,N_4849);
xor UO_138 (O_138,N_4857,N_4692);
nand UO_139 (O_139,N_4570,N_4590);
nor UO_140 (O_140,N_4996,N_4596);
or UO_141 (O_141,N_4963,N_4599);
xor UO_142 (O_142,N_4829,N_4525);
nor UO_143 (O_143,N_4674,N_4921);
or UO_144 (O_144,N_4992,N_4820);
nand UO_145 (O_145,N_4640,N_4643);
nand UO_146 (O_146,N_4949,N_4869);
nand UO_147 (O_147,N_4838,N_4887);
xor UO_148 (O_148,N_4561,N_4545);
and UO_149 (O_149,N_4850,N_4513);
nor UO_150 (O_150,N_4703,N_4556);
nand UO_151 (O_151,N_4765,N_4737);
and UO_152 (O_152,N_4520,N_4970);
nand UO_153 (O_153,N_4962,N_4745);
nand UO_154 (O_154,N_4841,N_4509);
nand UO_155 (O_155,N_4910,N_4597);
or UO_156 (O_156,N_4734,N_4689);
nand UO_157 (O_157,N_4515,N_4961);
and UO_158 (O_158,N_4976,N_4700);
or UO_159 (O_159,N_4582,N_4532);
or UO_160 (O_160,N_4528,N_4773);
or UO_161 (O_161,N_4645,N_4817);
nor UO_162 (O_162,N_4522,N_4718);
nand UO_163 (O_163,N_4828,N_4725);
nor UO_164 (O_164,N_4959,N_4801);
nor UO_165 (O_165,N_4742,N_4629);
nor UO_166 (O_166,N_4683,N_4505);
nor UO_167 (O_167,N_4723,N_4670);
or UO_168 (O_168,N_4701,N_4775);
nand UO_169 (O_169,N_4924,N_4547);
nand UO_170 (O_170,N_4698,N_4938);
or UO_171 (O_171,N_4595,N_4568);
and UO_172 (O_172,N_4876,N_4502);
nor UO_173 (O_173,N_4848,N_4537);
xor UO_174 (O_174,N_4727,N_4610);
nor UO_175 (O_175,N_4747,N_4755);
or UO_176 (O_176,N_4918,N_4685);
nor UO_177 (O_177,N_4642,N_4951);
or UO_178 (O_178,N_4759,N_4630);
nor UO_179 (O_179,N_4812,N_4821);
or UO_180 (O_180,N_4619,N_4691);
nand UO_181 (O_181,N_4724,N_4566);
nand UO_182 (O_182,N_4941,N_4541);
nor UO_183 (O_183,N_4653,N_4621);
nor UO_184 (O_184,N_4794,N_4983);
or UO_185 (O_185,N_4632,N_4555);
and UO_186 (O_186,N_4708,N_4588);
nand UO_187 (O_187,N_4874,N_4616);
and UO_188 (O_188,N_4843,N_4809);
and UO_189 (O_189,N_4862,N_4886);
nand UO_190 (O_190,N_4969,N_4531);
or UO_191 (O_191,N_4758,N_4800);
or UO_192 (O_192,N_4603,N_4627);
or UO_193 (O_193,N_4533,N_4892);
or UO_194 (O_194,N_4659,N_4982);
and UO_195 (O_195,N_4878,N_4953);
nand UO_196 (O_196,N_4625,N_4564);
or UO_197 (O_197,N_4777,N_4735);
and UO_198 (O_198,N_4554,N_4615);
nor UO_199 (O_199,N_4540,N_4824);
and UO_200 (O_200,N_4647,N_4504);
nand UO_201 (O_201,N_4648,N_4987);
nor UO_202 (O_202,N_4879,N_4894);
nand UO_203 (O_203,N_4583,N_4873);
or UO_204 (O_204,N_4774,N_4816);
or UO_205 (O_205,N_4613,N_4915);
nand UO_206 (O_206,N_4577,N_4818);
and UO_207 (O_207,N_4684,N_4732);
or UO_208 (O_208,N_4825,N_4663);
or UO_209 (O_209,N_4954,N_4854);
nand UO_210 (O_210,N_4709,N_4756);
and UO_211 (O_211,N_4935,N_4768);
xor UO_212 (O_212,N_4636,N_4827);
or UO_213 (O_213,N_4523,N_4882);
or UO_214 (O_214,N_4651,N_4678);
and UO_215 (O_215,N_4852,N_4908);
nand UO_216 (O_216,N_4793,N_4846);
nand UO_217 (O_217,N_4823,N_4697);
nand UO_218 (O_218,N_4916,N_4736);
nor UO_219 (O_219,N_4762,N_4644);
xnor UO_220 (O_220,N_4612,N_4552);
nand UO_221 (O_221,N_4993,N_4858);
and UO_222 (O_222,N_4958,N_4796);
or UO_223 (O_223,N_4549,N_4587);
and UO_224 (O_224,N_4729,N_4948);
or UO_225 (O_225,N_4646,N_4977);
and UO_226 (O_226,N_4805,N_4665);
nand UO_227 (O_227,N_4986,N_4922);
and UO_228 (O_228,N_4717,N_4655);
nor UO_229 (O_229,N_4622,N_4704);
and UO_230 (O_230,N_4624,N_4740);
and UO_231 (O_231,N_4778,N_4826);
nand UO_232 (O_232,N_4550,N_4720);
nor UO_233 (O_233,N_4960,N_4544);
and UO_234 (O_234,N_4614,N_4548);
nor UO_235 (O_235,N_4584,N_4508);
nor UO_236 (O_236,N_4965,N_4766);
nor UO_237 (O_237,N_4856,N_4730);
nand UO_238 (O_238,N_4521,N_4714);
nor UO_239 (O_239,N_4914,N_4897);
nor UO_240 (O_240,N_4968,N_4639);
nor UO_241 (O_241,N_4669,N_4956);
and UO_242 (O_242,N_4933,N_4860);
nand UO_243 (O_243,N_4538,N_4906);
and UO_244 (O_244,N_4749,N_4633);
nor UO_245 (O_245,N_4719,N_4797);
or UO_246 (O_246,N_4739,N_4586);
nor UO_247 (O_247,N_4609,N_4891);
and UO_248 (O_248,N_4864,N_4551);
nor UO_249 (O_249,N_4837,N_4738);
or UO_250 (O_250,N_4739,N_4867);
or UO_251 (O_251,N_4599,N_4671);
nand UO_252 (O_252,N_4880,N_4979);
and UO_253 (O_253,N_4600,N_4595);
nand UO_254 (O_254,N_4934,N_4755);
and UO_255 (O_255,N_4583,N_4645);
or UO_256 (O_256,N_4900,N_4808);
nand UO_257 (O_257,N_4872,N_4992);
nand UO_258 (O_258,N_4889,N_4624);
nand UO_259 (O_259,N_4888,N_4569);
nand UO_260 (O_260,N_4642,N_4554);
nand UO_261 (O_261,N_4574,N_4599);
or UO_262 (O_262,N_4995,N_4657);
and UO_263 (O_263,N_4997,N_4847);
and UO_264 (O_264,N_4569,N_4970);
nor UO_265 (O_265,N_4751,N_4918);
nor UO_266 (O_266,N_4624,N_4910);
or UO_267 (O_267,N_4704,N_4660);
or UO_268 (O_268,N_4871,N_4676);
or UO_269 (O_269,N_4896,N_4530);
nand UO_270 (O_270,N_4656,N_4995);
nand UO_271 (O_271,N_4652,N_4863);
nand UO_272 (O_272,N_4971,N_4755);
or UO_273 (O_273,N_4799,N_4946);
and UO_274 (O_274,N_4852,N_4771);
and UO_275 (O_275,N_4957,N_4984);
or UO_276 (O_276,N_4647,N_4882);
or UO_277 (O_277,N_4908,N_4975);
nor UO_278 (O_278,N_4985,N_4788);
nor UO_279 (O_279,N_4815,N_4672);
nor UO_280 (O_280,N_4705,N_4752);
and UO_281 (O_281,N_4509,N_4754);
nor UO_282 (O_282,N_4916,N_4515);
nand UO_283 (O_283,N_4840,N_4665);
or UO_284 (O_284,N_4644,N_4506);
nor UO_285 (O_285,N_4819,N_4949);
nand UO_286 (O_286,N_4875,N_4577);
or UO_287 (O_287,N_4695,N_4535);
or UO_288 (O_288,N_4819,N_4899);
nand UO_289 (O_289,N_4983,N_4674);
and UO_290 (O_290,N_4810,N_4876);
and UO_291 (O_291,N_4689,N_4654);
nand UO_292 (O_292,N_4762,N_4893);
or UO_293 (O_293,N_4997,N_4828);
and UO_294 (O_294,N_4592,N_4804);
nand UO_295 (O_295,N_4732,N_4935);
and UO_296 (O_296,N_4780,N_4728);
and UO_297 (O_297,N_4612,N_4862);
or UO_298 (O_298,N_4588,N_4911);
or UO_299 (O_299,N_4536,N_4849);
nor UO_300 (O_300,N_4781,N_4802);
nand UO_301 (O_301,N_4813,N_4659);
or UO_302 (O_302,N_4557,N_4989);
nor UO_303 (O_303,N_4805,N_4698);
nand UO_304 (O_304,N_4910,N_4732);
and UO_305 (O_305,N_4960,N_4894);
and UO_306 (O_306,N_4663,N_4639);
nand UO_307 (O_307,N_4871,N_4898);
nor UO_308 (O_308,N_4717,N_4788);
and UO_309 (O_309,N_4662,N_4977);
or UO_310 (O_310,N_4862,N_4707);
nor UO_311 (O_311,N_4925,N_4870);
nand UO_312 (O_312,N_4826,N_4593);
nand UO_313 (O_313,N_4975,N_4559);
nand UO_314 (O_314,N_4607,N_4633);
xnor UO_315 (O_315,N_4717,N_4925);
nand UO_316 (O_316,N_4967,N_4849);
and UO_317 (O_317,N_4512,N_4620);
or UO_318 (O_318,N_4659,N_4795);
nor UO_319 (O_319,N_4643,N_4667);
nand UO_320 (O_320,N_4519,N_4867);
or UO_321 (O_321,N_4664,N_4925);
and UO_322 (O_322,N_4567,N_4543);
or UO_323 (O_323,N_4512,N_4864);
or UO_324 (O_324,N_4603,N_4848);
nor UO_325 (O_325,N_4746,N_4775);
nor UO_326 (O_326,N_4975,N_4788);
and UO_327 (O_327,N_4535,N_4783);
and UO_328 (O_328,N_4846,N_4554);
nand UO_329 (O_329,N_4984,N_4972);
or UO_330 (O_330,N_4536,N_4843);
nor UO_331 (O_331,N_4590,N_4933);
nor UO_332 (O_332,N_4689,N_4683);
and UO_333 (O_333,N_4780,N_4740);
nor UO_334 (O_334,N_4654,N_4523);
nor UO_335 (O_335,N_4861,N_4779);
or UO_336 (O_336,N_4814,N_4682);
or UO_337 (O_337,N_4607,N_4566);
nand UO_338 (O_338,N_4922,N_4797);
nand UO_339 (O_339,N_4790,N_4976);
nor UO_340 (O_340,N_4520,N_4666);
nor UO_341 (O_341,N_4605,N_4600);
nand UO_342 (O_342,N_4907,N_4746);
nand UO_343 (O_343,N_4814,N_4840);
nand UO_344 (O_344,N_4974,N_4859);
nor UO_345 (O_345,N_4650,N_4686);
nor UO_346 (O_346,N_4906,N_4728);
xor UO_347 (O_347,N_4956,N_4916);
nor UO_348 (O_348,N_4718,N_4592);
or UO_349 (O_349,N_4723,N_4843);
nand UO_350 (O_350,N_4719,N_4532);
nand UO_351 (O_351,N_4801,N_4856);
nand UO_352 (O_352,N_4840,N_4603);
nand UO_353 (O_353,N_4988,N_4575);
nor UO_354 (O_354,N_4818,N_4883);
nand UO_355 (O_355,N_4695,N_4776);
and UO_356 (O_356,N_4726,N_4928);
nand UO_357 (O_357,N_4713,N_4540);
or UO_358 (O_358,N_4840,N_4768);
nor UO_359 (O_359,N_4982,N_4686);
or UO_360 (O_360,N_4813,N_4934);
nand UO_361 (O_361,N_4571,N_4777);
nand UO_362 (O_362,N_4899,N_4552);
and UO_363 (O_363,N_4553,N_4518);
and UO_364 (O_364,N_4502,N_4709);
and UO_365 (O_365,N_4942,N_4775);
nor UO_366 (O_366,N_4939,N_4505);
and UO_367 (O_367,N_4735,N_4983);
or UO_368 (O_368,N_4514,N_4513);
nand UO_369 (O_369,N_4716,N_4924);
nor UO_370 (O_370,N_4532,N_4561);
and UO_371 (O_371,N_4646,N_4704);
and UO_372 (O_372,N_4957,N_4553);
nor UO_373 (O_373,N_4672,N_4932);
and UO_374 (O_374,N_4802,N_4730);
nand UO_375 (O_375,N_4858,N_4840);
and UO_376 (O_376,N_4631,N_4890);
nand UO_377 (O_377,N_4665,N_4588);
nor UO_378 (O_378,N_4622,N_4947);
and UO_379 (O_379,N_4955,N_4584);
or UO_380 (O_380,N_4702,N_4682);
and UO_381 (O_381,N_4775,N_4972);
nor UO_382 (O_382,N_4699,N_4622);
nand UO_383 (O_383,N_4699,N_4619);
xor UO_384 (O_384,N_4924,N_4744);
or UO_385 (O_385,N_4929,N_4654);
and UO_386 (O_386,N_4954,N_4889);
and UO_387 (O_387,N_4867,N_4503);
nand UO_388 (O_388,N_4861,N_4565);
nand UO_389 (O_389,N_4663,N_4919);
or UO_390 (O_390,N_4806,N_4510);
and UO_391 (O_391,N_4853,N_4999);
nand UO_392 (O_392,N_4634,N_4501);
and UO_393 (O_393,N_4929,N_4648);
nand UO_394 (O_394,N_4903,N_4878);
or UO_395 (O_395,N_4709,N_4550);
nand UO_396 (O_396,N_4810,N_4827);
nand UO_397 (O_397,N_4734,N_4828);
xnor UO_398 (O_398,N_4828,N_4683);
and UO_399 (O_399,N_4995,N_4962);
nand UO_400 (O_400,N_4509,N_4558);
nor UO_401 (O_401,N_4921,N_4615);
nor UO_402 (O_402,N_4625,N_4546);
xnor UO_403 (O_403,N_4598,N_4888);
and UO_404 (O_404,N_4655,N_4757);
and UO_405 (O_405,N_4961,N_4791);
or UO_406 (O_406,N_4888,N_4913);
nand UO_407 (O_407,N_4847,N_4664);
or UO_408 (O_408,N_4521,N_4981);
nand UO_409 (O_409,N_4890,N_4996);
and UO_410 (O_410,N_4909,N_4731);
nor UO_411 (O_411,N_4759,N_4929);
nand UO_412 (O_412,N_4551,N_4680);
or UO_413 (O_413,N_4834,N_4537);
and UO_414 (O_414,N_4954,N_4714);
nor UO_415 (O_415,N_4808,N_4711);
or UO_416 (O_416,N_4630,N_4683);
and UO_417 (O_417,N_4803,N_4509);
and UO_418 (O_418,N_4973,N_4534);
nand UO_419 (O_419,N_4827,N_4803);
or UO_420 (O_420,N_4953,N_4664);
and UO_421 (O_421,N_4875,N_4558);
nand UO_422 (O_422,N_4620,N_4525);
and UO_423 (O_423,N_4502,N_4645);
or UO_424 (O_424,N_4583,N_4627);
and UO_425 (O_425,N_4784,N_4855);
or UO_426 (O_426,N_4877,N_4654);
and UO_427 (O_427,N_4514,N_4716);
nand UO_428 (O_428,N_4879,N_4583);
or UO_429 (O_429,N_4637,N_4705);
nor UO_430 (O_430,N_4955,N_4680);
xor UO_431 (O_431,N_4938,N_4703);
or UO_432 (O_432,N_4991,N_4932);
or UO_433 (O_433,N_4753,N_4828);
or UO_434 (O_434,N_4636,N_4966);
and UO_435 (O_435,N_4858,N_4861);
or UO_436 (O_436,N_4898,N_4864);
and UO_437 (O_437,N_4834,N_4672);
xnor UO_438 (O_438,N_4833,N_4500);
and UO_439 (O_439,N_4802,N_4880);
or UO_440 (O_440,N_4779,N_4512);
or UO_441 (O_441,N_4500,N_4532);
nand UO_442 (O_442,N_4884,N_4780);
or UO_443 (O_443,N_4968,N_4813);
or UO_444 (O_444,N_4945,N_4878);
nor UO_445 (O_445,N_4918,N_4729);
or UO_446 (O_446,N_4842,N_4817);
and UO_447 (O_447,N_4663,N_4914);
nor UO_448 (O_448,N_4773,N_4946);
and UO_449 (O_449,N_4702,N_4814);
or UO_450 (O_450,N_4752,N_4678);
nor UO_451 (O_451,N_4690,N_4981);
nand UO_452 (O_452,N_4717,N_4566);
nand UO_453 (O_453,N_4944,N_4575);
and UO_454 (O_454,N_4573,N_4924);
and UO_455 (O_455,N_4677,N_4923);
xnor UO_456 (O_456,N_4509,N_4572);
and UO_457 (O_457,N_4635,N_4836);
nand UO_458 (O_458,N_4846,N_4565);
nor UO_459 (O_459,N_4583,N_4938);
nand UO_460 (O_460,N_4531,N_4545);
nor UO_461 (O_461,N_4885,N_4783);
or UO_462 (O_462,N_4552,N_4949);
and UO_463 (O_463,N_4725,N_4805);
nand UO_464 (O_464,N_4938,N_4611);
nor UO_465 (O_465,N_4676,N_4522);
and UO_466 (O_466,N_4752,N_4902);
nor UO_467 (O_467,N_4518,N_4776);
nand UO_468 (O_468,N_4643,N_4890);
nand UO_469 (O_469,N_4776,N_4903);
xor UO_470 (O_470,N_4851,N_4746);
nor UO_471 (O_471,N_4917,N_4742);
nand UO_472 (O_472,N_4613,N_4636);
and UO_473 (O_473,N_4778,N_4825);
or UO_474 (O_474,N_4983,N_4878);
and UO_475 (O_475,N_4862,N_4879);
nor UO_476 (O_476,N_4965,N_4632);
nor UO_477 (O_477,N_4879,N_4786);
and UO_478 (O_478,N_4568,N_4635);
or UO_479 (O_479,N_4611,N_4919);
nor UO_480 (O_480,N_4729,N_4667);
and UO_481 (O_481,N_4765,N_4666);
nand UO_482 (O_482,N_4596,N_4794);
nand UO_483 (O_483,N_4828,N_4560);
nand UO_484 (O_484,N_4943,N_4924);
and UO_485 (O_485,N_4823,N_4779);
nor UO_486 (O_486,N_4808,N_4634);
or UO_487 (O_487,N_4764,N_4950);
nor UO_488 (O_488,N_4863,N_4984);
nor UO_489 (O_489,N_4590,N_4545);
or UO_490 (O_490,N_4897,N_4700);
nor UO_491 (O_491,N_4953,N_4543);
and UO_492 (O_492,N_4878,N_4908);
nor UO_493 (O_493,N_4817,N_4949);
and UO_494 (O_494,N_4792,N_4676);
nand UO_495 (O_495,N_4737,N_4601);
and UO_496 (O_496,N_4603,N_4642);
and UO_497 (O_497,N_4944,N_4888);
or UO_498 (O_498,N_4556,N_4646);
and UO_499 (O_499,N_4973,N_4914);
and UO_500 (O_500,N_4666,N_4897);
xor UO_501 (O_501,N_4523,N_4758);
and UO_502 (O_502,N_4795,N_4641);
nor UO_503 (O_503,N_4691,N_4669);
or UO_504 (O_504,N_4633,N_4817);
xor UO_505 (O_505,N_4822,N_4790);
or UO_506 (O_506,N_4857,N_4897);
nand UO_507 (O_507,N_4925,N_4804);
and UO_508 (O_508,N_4710,N_4625);
nor UO_509 (O_509,N_4641,N_4701);
and UO_510 (O_510,N_4749,N_4752);
nor UO_511 (O_511,N_4748,N_4881);
or UO_512 (O_512,N_4535,N_4984);
nor UO_513 (O_513,N_4950,N_4908);
nand UO_514 (O_514,N_4630,N_4520);
nand UO_515 (O_515,N_4836,N_4875);
and UO_516 (O_516,N_4634,N_4718);
or UO_517 (O_517,N_4564,N_4922);
or UO_518 (O_518,N_4562,N_4810);
nand UO_519 (O_519,N_4663,N_4769);
and UO_520 (O_520,N_4537,N_4950);
or UO_521 (O_521,N_4701,N_4809);
nand UO_522 (O_522,N_4748,N_4605);
nor UO_523 (O_523,N_4641,N_4691);
nor UO_524 (O_524,N_4588,N_4549);
and UO_525 (O_525,N_4881,N_4596);
or UO_526 (O_526,N_4649,N_4844);
and UO_527 (O_527,N_4512,N_4850);
nor UO_528 (O_528,N_4544,N_4659);
and UO_529 (O_529,N_4642,N_4637);
nor UO_530 (O_530,N_4610,N_4696);
nand UO_531 (O_531,N_4512,N_4800);
and UO_532 (O_532,N_4720,N_4884);
xnor UO_533 (O_533,N_4564,N_4983);
and UO_534 (O_534,N_4885,N_4825);
nand UO_535 (O_535,N_4586,N_4526);
nand UO_536 (O_536,N_4765,N_4995);
or UO_537 (O_537,N_4919,N_4753);
nand UO_538 (O_538,N_4720,N_4703);
nor UO_539 (O_539,N_4780,N_4616);
and UO_540 (O_540,N_4904,N_4953);
or UO_541 (O_541,N_4790,N_4904);
nand UO_542 (O_542,N_4531,N_4707);
nor UO_543 (O_543,N_4963,N_4565);
or UO_544 (O_544,N_4759,N_4812);
nor UO_545 (O_545,N_4675,N_4645);
or UO_546 (O_546,N_4737,N_4955);
and UO_547 (O_547,N_4896,N_4718);
nor UO_548 (O_548,N_4512,N_4517);
and UO_549 (O_549,N_4984,N_4995);
nor UO_550 (O_550,N_4549,N_4668);
and UO_551 (O_551,N_4765,N_4841);
or UO_552 (O_552,N_4676,N_4580);
and UO_553 (O_553,N_4906,N_4655);
or UO_554 (O_554,N_4713,N_4981);
xor UO_555 (O_555,N_4865,N_4602);
nand UO_556 (O_556,N_4607,N_4774);
and UO_557 (O_557,N_4603,N_4652);
nor UO_558 (O_558,N_4857,N_4674);
and UO_559 (O_559,N_4512,N_4810);
or UO_560 (O_560,N_4649,N_4794);
or UO_561 (O_561,N_4595,N_4980);
and UO_562 (O_562,N_4923,N_4966);
or UO_563 (O_563,N_4650,N_4558);
nor UO_564 (O_564,N_4576,N_4915);
nor UO_565 (O_565,N_4930,N_4820);
nand UO_566 (O_566,N_4927,N_4594);
nor UO_567 (O_567,N_4512,N_4983);
nand UO_568 (O_568,N_4992,N_4879);
or UO_569 (O_569,N_4676,N_4882);
and UO_570 (O_570,N_4674,N_4546);
nand UO_571 (O_571,N_4953,N_4972);
nor UO_572 (O_572,N_4689,N_4712);
or UO_573 (O_573,N_4783,N_4610);
nand UO_574 (O_574,N_4880,N_4686);
and UO_575 (O_575,N_4832,N_4921);
and UO_576 (O_576,N_4713,N_4580);
and UO_577 (O_577,N_4504,N_4502);
nand UO_578 (O_578,N_4615,N_4888);
nand UO_579 (O_579,N_4540,N_4573);
nand UO_580 (O_580,N_4624,N_4741);
nand UO_581 (O_581,N_4570,N_4731);
and UO_582 (O_582,N_4937,N_4536);
and UO_583 (O_583,N_4929,N_4928);
nor UO_584 (O_584,N_4659,N_4938);
and UO_585 (O_585,N_4739,N_4964);
and UO_586 (O_586,N_4935,N_4735);
nor UO_587 (O_587,N_4543,N_4546);
xor UO_588 (O_588,N_4567,N_4811);
or UO_589 (O_589,N_4889,N_4923);
nand UO_590 (O_590,N_4619,N_4809);
nor UO_591 (O_591,N_4643,N_4993);
nand UO_592 (O_592,N_4620,N_4996);
nand UO_593 (O_593,N_4840,N_4620);
nand UO_594 (O_594,N_4827,N_4984);
nand UO_595 (O_595,N_4729,N_4595);
or UO_596 (O_596,N_4573,N_4652);
xor UO_597 (O_597,N_4657,N_4620);
nand UO_598 (O_598,N_4758,N_4560);
and UO_599 (O_599,N_4864,N_4592);
or UO_600 (O_600,N_4561,N_4675);
or UO_601 (O_601,N_4952,N_4929);
or UO_602 (O_602,N_4887,N_4756);
and UO_603 (O_603,N_4838,N_4717);
nor UO_604 (O_604,N_4636,N_4609);
nand UO_605 (O_605,N_4637,N_4717);
nor UO_606 (O_606,N_4536,N_4586);
nand UO_607 (O_607,N_4719,N_4990);
or UO_608 (O_608,N_4972,N_4715);
and UO_609 (O_609,N_4889,N_4876);
nand UO_610 (O_610,N_4691,N_4775);
or UO_611 (O_611,N_4903,N_4572);
nor UO_612 (O_612,N_4923,N_4993);
nand UO_613 (O_613,N_4590,N_4758);
nor UO_614 (O_614,N_4554,N_4741);
nand UO_615 (O_615,N_4662,N_4830);
or UO_616 (O_616,N_4593,N_4993);
nand UO_617 (O_617,N_4967,N_4716);
and UO_618 (O_618,N_4608,N_4704);
and UO_619 (O_619,N_4592,N_4806);
nand UO_620 (O_620,N_4582,N_4684);
or UO_621 (O_621,N_4716,N_4614);
nand UO_622 (O_622,N_4633,N_4685);
nor UO_623 (O_623,N_4609,N_4884);
nand UO_624 (O_624,N_4529,N_4541);
xnor UO_625 (O_625,N_4829,N_4632);
nor UO_626 (O_626,N_4682,N_4716);
nand UO_627 (O_627,N_4662,N_4660);
and UO_628 (O_628,N_4665,N_4788);
nor UO_629 (O_629,N_4607,N_4833);
and UO_630 (O_630,N_4793,N_4715);
and UO_631 (O_631,N_4779,N_4791);
nand UO_632 (O_632,N_4939,N_4958);
nor UO_633 (O_633,N_4771,N_4987);
nor UO_634 (O_634,N_4901,N_4823);
and UO_635 (O_635,N_4532,N_4648);
nand UO_636 (O_636,N_4523,N_4864);
or UO_637 (O_637,N_4756,N_4882);
nand UO_638 (O_638,N_4645,N_4980);
or UO_639 (O_639,N_4916,N_4513);
nand UO_640 (O_640,N_4927,N_4893);
and UO_641 (O_641,N_4882,N_4705);
or UO_642 (O_642,N_4667,N_4665);
nor UO_643 (O_643,N_4967,N_4662);
or UO_644 (O_644,N_4559,N_4823);
nor UO_645 (O_645,N_4800,N_4716);
or UO_646 (O_646,N_4674,N_4860);
or UO_647 (O_647,N_4804,N_4661);
nor UO_648 (O_648,N_4678,N_4748);
and UO_649 (O_649,N_4577,N_4797);
and UO_650 (O_650,N_4935,N_4529);
nor UO_651 (O_651,N_4856,N_4842);
and UO_652 (O_652,N_4665,N_4640);
nand UO_653 (O_653,N_4803,N_4745);
and UO_654 (O_654,N_4630,N_4646);
or UO_655 (O_655,N_4792,N_4783);
or UO_656 (O_656,N_4721,N_4860);
nor UO_657 (O_657,N_4843,N_4624);
nor UO_658 (O_658,N_4541,N_4685);
and UO_659 (O_659,N_4686,N_4946);
nor UO_660 (O_660,N_4949,N_4602);
nand UO_661 (O_661,N_4511,N_4582);
and UO_662 (O_662,N_4754,N_4767);
xor UO_663 (O_663,N_4507,N_4605);
or UO_664 (O_664,N_4655,N_4674);
or UO_665 (O_665,N_4630,N_4657);
or UO_666 (O_666,N_4588,N_4775);
or UO_667 (O_667,N_4690,N_4990);
or UO_668 (O_668,N_4569,N_4996);
nand UO_669 (O_669,N_4673,N_4582);
nor UO_670 (O_670,N_4774,N_4713);
or UO_671 (O_671,N_4673,N_4891);
nand UO_672 (O_672,N_4923,N_4552);
and UO_673 (O_673,N_4721,N_4768);
and UO_674 (O_674,N_4699,N_4979);
nor UO_675 (O_675,N_4611,N_4921);
and UO_676 (O_676,N_4519,N_4829);
and UO_677 (O_677,N_4603,N_4753);
and UO_678 (O_678,N_4531,N_4554);
nor UO_679 (O_679,N_4812,N_4845);
and UO_680 (O_680,N_4799,N_4591);
nand UO_681 (O_681,N_4910,N_4924);
nand UO_682 (O_682,N_4818,N_4753);
nand UO_683 (O_683,N_4886,N_4626);
nor UO_684 (O_684,N_4944,N_4845);
nand UO_685 (O_685,N_4719,N_4638);
or UO_686 (O_686,N_4587,N_4917);
and UO_687 (O_687,N_4802,N_4596);
nand UO_688 (O_688,N_4874,N_4597);
and UO_689 (O_689,N_4776,N_4862);
nor UO_690 (O_690,N_4840,N_4958);
and UO_691 (O_691,N_4676,N_4675);
nor UO_692 (O_692,N_4503,N_4792);
nor UO_693 (O_693,N_4999,N_4701);
nand UO_694 (O_694,N_4829,N_4529);
and UO_695 (O_695,N_4663,N_4504);
and UO_696 (O_696,N_4538,N_4865);
and UO_697 (O_697,N_4805,N_4743);
nand UO_698 (O_698,N_4737,N_4670);
nor UO_699 (O_699,N_4575,N_4786);
nor UO_700 (O_700,N_4510,N_4826);
nor UO_701 (O_701,N_4629,N_4884);
or UO_702 (O_702,N_4875,N_4753);
and UO_703 (O_703,N_4902,N_4846);
and UO_704 (O_704,N_4718,N_4834);
nand UO_705 (O_705,N_4580,N_4726);
nor UO_706 (O_706,N_4672,N_4773);
nand UO_707 (O_707,N_4848,N_4689);
or UO_708 (O_708,N_4813,N_4923);
and UO_709 (O_709,N_4807,N_4826);
or UO_710 (O_710,N_4690,N_4606);
or UO_711 (O_711,N_4670,N_4531);
xnor UO_712 (O_712,N_4893,N_4752);
and UO_713 (O_713,N_4699,N_4967);
or UO_714 (O_714,N_4569,N_4840);
nand UO_715 (O_715,N_4926,N_4914);
nand UO_716 (O_716,N_4511,N_4768);
and UO_717 (O_717,N_4645,N_4787);
and UO_718 (O_718,N_4692,N_4540);
nand UO_719 (O_719,N_4945,N_4665);
and UO_720 (O_720,N_4782,N_4953);
nor UO_721 (O_721,N_4539,N_4830);
or UO_722 (O_722,N_4734,N_4632);
nand UO_723 (O_723,N_4814,N_4539);
nand UO_724 (O_724,N_4878,N_4666);
and UO_725 (O_725,N_4890,N_4902);
nand UO_726 (O_726,N_4718,N_4590);
nand UO_727 (O_727,N_4641,N_4988);
nand UO_728 (O_728,N_4511,N_4972);
and UO_729 (O_729,N_4640,N_4590);
or UO_730 (O_730,N_4702,N_4816);
nor UO_731 (O_731,N_4743,N_4834);
nand UO_732 (O_732,N_4578,N_4932);
nand UO_733 (O_733,N_4899,N_4915);
or UO_734 (O_734,N_4569,N_4726);
and UO_735 (O_735,N_4784,N_4687);
nor UO_736 (O_736,N_4910,N_4528);
and UO_737 (O_737,N_4655,N_4779);
or UO_738 (O_738,N_4555,N_4602);
and UO_739 (O_739,N_4519,N_4791);
or UO_740 (O_740,N_4859,N_4731);
or UO_741 (O_741,N_4799,N_4701);
nor UO_742 (O_742,N_4708,N_4568);
or UO_743 (O_743,N_4931,N_4618);
or UO_744 (O_744,N_4915,N_4860);
nand UO_745 (O_745,N_4695,N_4750);
nand UO_746 (O_746,N_4619,N_4676);
nor UO_747 (O_747,N_4629,N_4812);
and UO_748 (O_748,N_4996,N_4676);
nor UO_749 (O_749,N_4607,N_4818);
nor UO_750 (O_750,N_4784,N_4748);
and UO_751 (O_751,N_4578,N_4626);
or UO_752 (O_752,N_4505,N_4526);
and UO_753 (O_753,N_4997,N_4640);
nand UO_754 (O_754,N_4699,N_4826);
and UO_755 (O_755,N_4836,N_4794);
and UO_756 (O_756,N_4963,N_4583);
and UO_757 (O_757,N_4903,N_4606);
or UO_758 (O_758,N_4616,N_4758);
nand UO_759 (O_759,N_4609,N_4971);
nand UO_760 (O_760,N_4511,N_4887);
and UO_761 (O_761,N_4591,N_4894);
and UO_762 (O_762,N_4796,N_4713);
or UO_763 (O_763,N_4688,N_4974);
nand UO_764 (O_764,N_4939,N_4632);
nand UO_765 (O_765,N_4536,N_4853);
nand UO_766 (O_766,N_4777,N_4644);
nor UO_767 (O_767,N_4861,N_4697);
nor UO_768 (O_768,N_4716,N_4522);
or UO_769 (O_769,N_4641,N_4511);
or UO_770 (O_770,N_4777,N_4677);
nand UO_771 (O_771,N_4845,N_4585);
nand UO_772 (O_772,N_4925,N_4635);
or UO_773 (O_773,N_4629,N_4994);
or UO_774 (O_774,N_4968,N_4623);
or UO_775 (O_775,N_4550,N_4764);
nand UO_776 (O_776,N_4730,N_4967);
nor UO_777 (O_777,N_4879,N_4572);
or UO_778 (O_778,N_4930,N_4717);
or UO_779 (O_779,N_4785,N_4741);
or UO_780 (O_780,N_4808,N_4602);
nor UO_781 (O_781,N_4942,N_4800);
or UO_782 (O_782,N_4740,N_4744);
and UO_783 (O_783,N_4988,N_4548);
nand UO_784 (O_784,N_4693,N_4899);
or UO_785 (O_785,N_4777,N_4975);
and UO_786 (O_786,N_4504,N_4776);
or UO_787 (O_787,N_4832,N_4947);
or UO_788 (O_788,N_4628,N_4758);
xnor UO_789 (O_789,N_4914,N_4632);
xor UO_790 (O_790,N_4661,N_4793);
nor UO_791 (O_791,N_4501,N_4671);
and UO_792 (O_792,N_4721,N_4863);
nor UO_793 (O_793,N_4621,N_4560);
nor UO_794 (O_794,N_4597,N_4659);
nor UO_795 (O_795,N_4786,N_4556);
and UO_796 (O_796,N_4925,N_4797);
nand UO_797 (O_797,N_4956,N_4987);
and UO_798 (O_798,N_4939,N_4698);
or UO_799 (O_799,N_4754,N_4879);
nor UO_800 (O_800,N_4979,N_4607);
nand UO_801 (O_801,N_4983,N_4820);
or UO_802 (O_802,N_4514,N_4616);
nand UO_803 (O_803,N_4679,N_4557);
or UO_804 (O_804,N_4961,N_4674);
and UO_805 (O_805,N_4591,N_4941);
or UO_806 (O_806,N_4789,N_4525);
and UO_807 (O_807,N_4923,N_4681);
nor UO_808 (O_808,N_4863,N_4521);
nand UO_809 (O_809,N_4647,N_4834);
nand UO_810 (O_810,N_4844,N_4931);
nand UO_811 (O_811,N_4794,N_4997);
nor UO_812 (O_812,N_4904,N_4613);
or UO_813 (O_813,N_4561,N_4668);
nor UO_814 (O_814,N_4603,N_4878);
nand UO_815 (O_815,N_4999,N_4954);
and UO_816 (O_816,N_4676,N_4961);
or UO_817 (O_817,N_4966,N_4696);
nor UO_818 (O_818,N_4777,N_4792);
and UO_819 (O_819,N_4789,N_4917);
and UO_820 (O_820,N_4905,N_4999);
or UO_821 (O_821,N_4955,N_4596);
nand UO_822 (O_822,N_4854,N_4639);
or UO_823 (O_823,N_4702,N_4887);
nor UO_824 (O_824,N_4910,N_4810);
or UO_825 (O_825,N_4558,N_4569);
nand UO_826 (O_826,N_4764,N_4633);
and UO_827 (O_827,N_4561,N_4764);
nand UO_828 (O_828,N_4688,N_4908);
nor UO_829 (O_829,N_4748,N_4948);
nand UO_830 (O_830,N_4919,N_4851);
nand UO_831 (O_831,N_4699,N_4848);
nand UO_832 (O_832,N_4892,N_4768);
and UO_833 (O_833,N_4633,N_4683);
nor UO_834 (O_834,N_4916,N_4943);
nand UO_835 (O_835,N_4912,N_4581);
nor UO_836 (O_836,N_4962,N_4758);
and UO_837 (O_837,N_4737,N_4992);
nor UO_838 (O_838,N_4704,N_4839);
or UO_839 (O_839,N_4573,N_4762);
nor UO_840 (O_840,N_4564,N_4830);
nand UO_841 (O_841,N_4981,N_4938);
and UO_842 (O_842,N_4951,N_4899);
nand UO_843 (O_843,N_4961,N_4977);
or UO_844 (O_844,N_4591,N_4933);
nor UO_845 (O_845,N_4820,N_4640);
or UO_846 (O_846,N_4621,N_4799);
nor UO_847 (O_847,N_4527,N_4534);
or UO_848 (O_848,N_4791,N_4855);
nand UO_849 (O_849,N_4799,N_4723);
and UO_850 (O_850,N_4684,N_4907);
nor UO_851 (O_851,N_4973,N_4563);
and UO_852 (O_852,N_4899,N_4707);
xor UO_853 (O_853,N_4611,N_4637);
and UO_854 (O_854,N_4715,N_4805);
or UO_855 (O_855,N_4816,N_4759);
and UO_856 (O_856,N_4562,N_4646);
and UO_857 (O_857,N_4556,N_4873);
and UO_858 (O_858,N_4511,N_4703);
nor UO_859 (O_859,N_4649,N_4936);
or UO_860 (O_860,N_4773,N_4915);
nor UO_861 (O_861,N_4868,N_4948);
and UO_862 (O_862,N_4947,N_4744);
nand UO_863 (O_863,N_4646,N_4707);
or UO_864 (O_864,N_4553,N_4531);
and UO_865 (O_865,N_4981,N_4788);
nor UO_866 (O_866,N_4979,N_4889);
or UO_867 (O_867,N_4842,N_4823);
nor UO_868 (O_868,N_4746,N_4583);
xor UO_869 (O_869,N_4550,N_4867);
and UO_870 (O_870,N_4546,N_4827);
or UO_871 (O_871,N_4862,N_4868);
and UO_872 (O_872,N_4952,N_4764);
and UO_873 (O_873,N_4896,N_4726);
and UO_874 (O_874,N_4920,N_4694);
nor UO_875 (O_875,N_4681,N_4919);
nor UO_876 (O_876,N_4939,N_4795);
and UO_877 (O_877,N_4676,N_4976);
and UO_878 (O_878,N_4699,N_4661);
and UO_879 (O_879,N_4952,N_4780);
and UO_880 (O_880,N_4770,N_4750);
nor UO_881 (O_881,N_4898,N_4788);
and UO_882 (O_882,N_4988,N_4511);
and UO_883 (O_883,N_4540,N_4861);
nor UO_884 (O_884,N_4553,N_4570);
nor UO_885 (O_885,N_4914,N_4935);
nor UO_886 (O_886,N_4879,N_4939);
nand UO_887 (O_887,N_4866,N_4561);
and UO_888 (O_888,N_4512,N_4773);
nand UO_889 (O_889,N_4777,N_4807);
or UO_890 (O_890,N_4963,N_4973);
or UO_891 (O_891,N_4835,N_4841);
nor UO_892 (O_892,N_4561,N_4985);
nand UO_893 (O_893,N_4565,N_4732);
nor UO_894 (O_894,N_4851,N_4565);
or UO_895 (O_895,N_4540,N_4799);
and UO_896 (O_896,N_4745,N_4501);
nor UO_897 (O_897,N_4758,N_4600);
nand UO_898 (O_898,N_4836,N_4740);
nand UO_899 (O_899,N_4970,N_4972);
nand UO_900 (O_900,N_4696,N_4706);
nor UO_901 (O_901,N_4999,N_4641);
nor UO_902 (O_902,N_4945,N_4608);
nand UO_903 (O_903,N_4938,N_4809);
or UO_904 (O_904,N_4830,N_4711);
and UO_905 (O_905,N_4518,N_4988);
nor UO_906 (O_906,N_4645,N_4877);
or UO_907 (O_907,N_4659,N_4630);
or UO_908 (O_908,N_4998,N_4750);
and UO_909 (O_909,N_4544,N_4984);
nand UO_910 (O_910,N_4754,N_4810);
or UO_911 (O_911,N_4907,N_4974);
nor UO_912 (O_912,N_4526,N_4851);
and UO_913 (O_913,N_4836,N_4523);
or UO_914 (O_914,N_4731,N_4631);
or UO_915 (O_915,N_4709,N_4722);
nor UO_916 (O_916,N_4678,N_4914);
nand UO_917 (O_917,N_4895,N_4893);
or UO_918 (O_918,N_4684,N_4826);
nand UO_919 (O_919,N_4631,N_4847);
and UO_920 (O_920,N_4978,N_4521);
nor UO_921 (O_921,N_4880,N_4845);
and UO_922 (O_922,N_4924,N_4989);
nor UO_923 (O_923,N_4971,N_4546);
nor UO_924 (O_924,N_4944,N_4806);
or UO_925 (O_925,N_4934,N_4522);
nor UO_926 (O_926,N_4731,N_4708);
or UO_927 (O_927,N_4593,N_4530);
and UO_928 (O_928,N_4671,N_4701);
or UO_929 (O_929,N_4777,N_4952);
nor UO_930 (O_930,N_4685,N_4501);
xor UO_931 (O_931,N_4771,N_4630);
xnor UO_932 (O_932,N_4739,N_4601);
and UO_933 (O_933,N_4812,N_4583);
nor UO_934 (O_934,N_4562,N_4571);
nor UO_935 (O_935,N_4756,N_4799);
or UO_936 (O_936,N_4677,N_4580);
nor UO_937 (O_937,N_4869,N_4988);
or UO_938 (O_938,N_4610,N_4534);
and UO_939 (O_939,N_4664,N_4702);
and UO_940 (O_940,N_4948,N_4529);
nand UO_941 (O_941,N_4552,N_4993);
and UO_942 (O_942,N_4650,N_4646);
nand UO_943 (O_943,N_4693,N_4972);
and UO_944 (O_944,N_4503,N_4581);
and UO_945 (O_945,N_4564,N_4656);
nor UO_946 (O_946,N_4997,N_4991);
nor UO_947 (O_947,N_4990,N_4900);
or UO_948 (O_948,N_4563,N_4990);
nor UO_949 (O_949,N_4610,N_4644);
xnor UO_950 (O_950,N_4657,N_4504);
or UO_951 (O_951,N_4688,N_4579);
nand UO_952 (O_952,N_4646,N_4561);
and UO_953 (O_953,N_4514,N_4548);
nand UO_954 (O_954,N_4966,N_4502);
nor UO_955 (O_955,N_4671,N_4797);
and UO_956 (O_956,N_4766,N_4748);
nand UO_957 (O_957,N_4623,N_4670);
nand UO_958 (O_958,N_4542,N_4778);
or UO_959 (O_959,N_4549,N_4519);
and UO_960 (O_960,N_4979,N_4723);
nor UO_961 (O_961,N_4877,N_4918);
and UO_962 (O_962,N_4850,N_4500);
or UO_963 (O_963,N_4935,N_4928);
nor UO_964 (O_964,N_4955,N_4882);
nand UO_965 (O_965,N_4811,N_4564);
or UO_966 (O_966,N_4759,N_4591);
nor UO_967 (O_967,N_4922,N_4760);
nand UO_968 (O_968,N_4531,N_4535);
and UO_969 (O_969,N_4773,N_4763);
nor UO_970 (O_970,N_4987,N_4937);
nor UO_971 (O_971,N_4905,N_4824);
and UO_972 (O_972,N_4529,N_4623);
nor UO_973 (O_973,N_4882,N_4837);
or UO_974 (O_974,N_4872,N_4967);
nor UO_975 (O_975,N_4579,N_4509);
xor UO_976 (O_976,N_4582,N_4734);
nor UO_977 (O_977,N_4761,N_4886);
nand UO_978 (O_978,N_4757,N_4678);
nand UO_979 (O_979,N_4992,N_4814);
nor UO_980 (O_980,N_4615,N_4840);
nand UO_981 (O_981,N_4788,N_4726);
nand UO_982 (O_982,N_4744,N_4990);
and UO_983 (O_983,N_4857,N_4891);
or UO_984 (O_984,N_4749,N_4581);
nor UO_985 (O_985,N_4556,N_4690);
and UO_986 (O_986,N_4662,N_4953);
nand UO_987 (O_987,N_4957,N_4737);
nor UO_988 (O_988,N_4756,N_4870);
xor UO_989 (O_989,N_4748,N_4863);
nor UO_990 (O_990,N_4571,N_4631);
and UO_991 (O_991,N_4896,N_4948);
nand UO_992 (O_992,N_4779,N_4974);
nand UO_993 (O_993,N_4570,N_4921);
nor UO_994 (O_994,N_4980,N_4948);
or UO_995 (O_995,N_4592,N_4697);
nand UO_996 (O_996,N_4704,N_4526);
nor UO_997 (O_997,N_4864,N_4908);
nor UO_998 (O_998,N_4736,N_4606);
or UO_999 (O_999,N_4915,N_4517);
endmodule