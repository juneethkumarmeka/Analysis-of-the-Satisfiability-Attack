module basic_5000_50000_5000_10_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_1893,In_1178);
xnor U1 (N_1,In_4572,In_2636);
nor U2 (N_2,In_798,In_2158);
or U3 (N_3,In_2623,In_3781);
nand U4 (N_4,In_4633,In_4521);
xnor U5 (N_5,In_3402,In_2490);
or U6 (N_6,In_2909,In_3252);
and U7 (N_7,In_1203,In_2778);
or U8 (N_8,In_1008,In_2420);
or U9 (N_9,In_3344,In_1022);
xor U10 (N_10,In_2143,In_582);
xor U11 (N_11,In_2065,In_415);
nand U12 (N_12,In_4517,In_2779);
and U13 (N_13,In_3112,In_2245);
and U14 (N_14,In_3241,In_932);
nand U15 (N_15,In_4417,In_3040);
and U16 (N_16,In_631,In_4072);
nor U17 (N_17,In_4801,In_4411);
and U18 (N_18,In_3139,In_1176);
xnor U19 (N_19,In_2436,In_16);
xor U20 (N_20,In_803,In_2456);
nor U21 (N_21,In_1113,In_2237);
or U22 (N_22,In_1272,In_3833);
or U23 (N_23,In_2645,In_3789);
nor U24 (N_24,In_32,In_4172);
nor U25 (N_25,In_407,In_1586);
and U26 (N_26,In_209,In_2206);
nand U27 (N_27,In_164,In_672);
nand U28 (N_28,In_3347,In_4933);
and U29 (N_29,In_1296,In_4452);
xnor U30 (N_30,In_1096,In_756);
or U31 (N_31,In_3596,In_2032);
nor U32 (N_32,In_4445,In_4765);
nor U33 (N_33,In_2685,In_1835);
nor U34 (N_34,In_3435,In_2507);
xor U35 (N_35,In_3963,In_1352);
xor U36 (N_36,In_1124,In_2125);
nand U37 (N_37,In_1450,In_670);
nor U38 (N_38,In_1307,In_1392);
nor U39 (N_39,In_982,In_4114);
xor U40 (N_40,In_3934,In_3991);
nor U41 (N_41,In_1923,In_2928);
xnor U42 (N_42,In_1066,In_2982);
or U43 (N_43,In_1942,In_1711);
xnor U44 (N_44,In_3981,In_2362);
nor U45 (N_45,In_3788,In_4885);
nand U46 (N_46,In_1384,In_810);
nand U47 (N_47,In_3427,In_2568);
xor U48 (N_48,In_2062,In_4512);
xor U49 (N_49,In_3911,In_4320);
xnor U50 (N_50,In_4814,In_1471);
or U51 (N_51,In_2268,In_1299);
xor U52 (N_52,In_3356,In_3135);
nor U53 (N_53,In_2298,In_1836);
nand U54 (N_54,In_4919,In_4273);
or U55 (N_55,In_3971,In_4668);
or U56 (N_56,In_4753,In_2885);
or U57 (N_57,In_2642,In_524);
or U58 (N_58,In_4429,In_1201);
and U59 (N_59,In_2825,In_436);
nor U60 (N_60,In_2677,In_2051);
nor U61 (N_61,In_267,In_2147);
nand U62 (N_62,In_2458,In_910);
nand U63 (N_63,In_4901,In_1441);
nor U64 (N_64,In_508,In_663);
xnor U65 (N_65,In_4524,In_3632);
nand U66 (N_66,In_198,In_3742);
or U67 (N_67,In_4370,In_1199);
xnor U68 (N_68,In_4745,In_4364);
nand U69 (N_69,In_4711,In_3228);
and U70 (N_70,In_103,In_3671);
nand U71 (N_71,In_3281,In_2790);
or U72 (N_72,In_4091,In_4568);
and U73 (N_73,In_1379,In_2750);
xor U74 (N_74,In_378,In_423);
and U75 (N_75,In_3469,In_2983);
nor U76 (N_76,In_1579,In_4421);
xnor U77 (N_77,In_1398,In_657);
nand U78 (N_78,In_27,In_2566);
nor U79 (N_79,In_4913,In_3797);
xor U80 (N_80,In_2075,In_2653);
xnor U81 (N_81,In_3711,In_4880);
nor U82 (N_82,In_3350,In_943);
nor U83 (N_83,In_2647,In_2441);
nand U84 (N_84,In_3495,In_3216);
or U85 (N_85,In_909,In_1727);
or U86 (N_86,In_2678,In_1062);
nand U87 (N_87,In_2700,In_1157);
nand U88 (N_88,In_466,In_4463);
or U89 (N_89,In_2788,In_2227);
or U90 (N_90,In_97,In_4466);
xor U91 (N_91,In_5,In_2011);
and U92 (N_92,In_2730,In_763);
or U93 (N_93,In_3527,In_1475);
and U94 (N_94,In_3816,In_2046);
nand U95 (N_95,In_4790,In_695);
nor U96 (N_96,In_2500,In_2088);
nor U97 (N_97,In_79,In_4026);
nand U98 (N_98,In_3052,In_2893);
and U99 (N_99,In_2090,In_2590);
nor U100 (N_100,In_2680,In_3085);
nand U101 (N_101,In_2621,In_3403);
and U102 (N_102,In_1361,In_3461);
nor U103 (N_103,In_2320,In_971);
and U104 (N_104,In_4870,In_2749);
or U105 (N_105,In_1101,In_3813);
nand U106 (N_106,In_4247,In_4194);
xnor U107 (N_107,In_3902,In_3299);
or U108 (N_108,In_3201,In_3206);
xor U109 (N_109,In_937,In_2810);
nand U110 (N_110,In_1954,In_231);
and U111 (N_111,In_912,In_1969);
nand U112 (N_112,In_1269,In_1216);
nand U113 (N_113,In_404,In_1154);
nor U114 (N_114,In_282,In_4553);
or U115 (N_115,In_4966,In_3587);
nor U116 (N_116,In_2817,In_4991);
nor U117 (N_117,In_17,In_3222);
nand U118 (N_118,In_2084,In_2388);
nand U119 (N_119,In_690,In_4415);
and U120 (N_120,In_2694,In_1280);
or U121 (N_121,In_3412,In_1487);
xnor U122 (N_122,In_1140,In_3317);
xnor U123 (N_123,In_2965,In_3338);
xor U124 (N_124,In_2048,In_4268);
xnor U125 (N_125,In_3978,In_2403);
or U126 (N_126,In_111,In_2005);
or U127 (N_127,In_2676,In_2247);
and U128 (N_128,In_1063,In_2401);
nand U129 (N_129,In_1552,In_1184);
and U130 (N_130,In_2987,In_202);
xor U131 (N_131,In_235,In_2714);
nand U132 (N_132,In_3232,In_1055);
xor U133 (N_133,In_641,In_1052);
nor U134 (N_134,In_4506,In_1736);
nand U135 (N_135,In_3472,In_705);
xnor U136 (N_136,In_2275,In_789);
and U137 (N_137,In_1015,In_4890);
and U138 (N_138,In_1111,In_3582);
and U139 (N_139,In_1224,In_3101);
nor U140 (N_140,In_921,In_3354);
and U141 (N_141,In_2086,In_3834);
xnor U142 (N_142,In_1051,In_792);
nor U143 (N_143,In_4462,In_2657);
nor U144 (N_144,In_479,In_454);
and U145 (N_145,In_1625,In_1229);
and U146 (N_146,In_2408,In_4944);
nand U147 (N_147,In_4059,In_2555);
or U148 (N_148,In_176,In_3968);
nand U149 (N_149,In_1328,In_1356);
and U150 (N_150,In_2070,In_3415);
xnor U151 (N_151,In_4089,In_4135);
nor U152 (N_152,In_1911,In_1597);
nor U153 (N_153,In_4938,In_295);
xor U154 (N_154,In_3882,In_658);
nor U155 (N_155,In_3523,In_2469);
nand U156 (N_156,In_96,In_3308);
or U157 (N_157,In_2951,In_775);
nand U158 (N_158,In_1035,In_2731);
or U159 (N_159,In_4625,In_129);
xnor U160 (N_160,In_4844,In_1568);
and U161 (N_161,In_880,In_4086);
xnor U162 (N_162,In_4929,In_3726);
and U163 (N_163,In_2493,In_4393);
nand U164 (N_164,In_2703,In_2650);
xnor U165 (N_165,In_4839,In_2930);
nor U166 (N_166,In_2226,In_1455);
or U167 (N_167,In_1630,In_1653);
and U168 (N_168,In_579,In_4490);
nand U169 (N_169,In_2850,In_529);
nor U170 (N_170,In_2785,In_519);
xor U171 (N_171,In_4627,In_3183);
and U172 (N_172,In_1150,In_1145);
or U173 (N_173,In_2682,In_4994);
or U174 (N_174,In_289,In_2382);
nand U175 (N_175,In_1517,In_4332);
nand U176 (N_176,In_714,In_2061);
and U177 (N_177,In_911,In_3001);
and U178 (N_178,In_2486,In_4518);
xor U179 (N_179,In_1849,In_3930);
xor U180 (N_180,In_685,In_4094);
or U181 (N_181,In_3369,In_1223);
and U182 (N_182,In_4055,In_2066);
nor U183 (N_183,In_1857,In_1615);
and U184 (N_184,In_4593,In_4315);
nand U185 (N_185,In_2586,In_3310);
nor U186 (N_186,In_2472,In_4063);
and U187 (N_187,In_2905,In_3832);
nor U188 (N_188,In_9,In_4592);
xnor U189 (N_189,In_3449,In_443);
xnor U190 (N_190,In_884,In_1276);
nand U191 (N_191,In_4514,In_3236);
and U192 (N_192,In_1335,In_2457);
and U193 (N_193,In_3856,In_874);
nor U194 (N_194,In_1745,In_1360);
nor U195 (N_195,In_310,In_4990);
nand U196 (N_196,In_1030,In_1695);
nor U197 (N_197,In_2243,In_2018);
or U198 (N_198,In_1365,In_3055);
or U199 (N_199,In_4961,In_3429);
nand U200 (N_200,In_2414,In_424);
and U201 (N_201,In_1612,In_1827);
and U202 (N_202,In_2522,In_2721);
or U203 (N_203,In_486,In_3740);
or U204 (N_204,In_2350,In_563);
nand U205 (N_205,In_3257,In_1733);
nand U206 (N_206,In_456,In_2877);
nor U207 (N_207,In_681,In_550);
nor U208 (N_208,In_2324,In_1758);
nand U209 (N_209,In_1875,In_4000);
nand U210 (N_210,In_4178,In_3096);
nand U211 (N_211,In_1075,In_1872);
and U212 (N_212,In_1249,In_3368);
xnor U213 (N_213,In_2985,In_481);
or U214 (N_214,In_1231,In_3887);
nor U215 (N_215,In_2935,In_4726);
and U216 (N_216,In_1924,In_4478);
or U217 (N_217,In_1316,In_1795);
nand U218 (N_218,In_3130,In_3876);
nand U219 (N_219,In_457,In_2199);
nor U220 (N_220,In_1886,In_3842);
nand U221 (N_221,In_2034,In_1342);
nand U222 (N_222,In_718,In_4326);
or U223 (N_223,In_1033,In_4103);
or U224 (N_224,In_938,In_3168);
nand U225 (N_225,In_3825,In_3056);
nor U226 (N_226,In_2156,In_1207);
xor U227 (N_227,In_4508,In_1898);
xnor U228 (N_228,In_854,In_852);
nor U229 (N_229,In_553,In_419);
nor U230 (N_230,In_460,In_3197);
xor U231 (N_231,In_4049,In_3117);
and U232 (N_232,In_3548,In_3549);
and U233 (N_233,In_967,In_2686);
or U234 (N_234,In_108,In_3697);
and U235 (N_235,In_1003,In_2525);
or U236 (N_236,In_2105,In_2166);
nand U237 (N_237,In_4276,In_1071);
and U238 (N_238,In_3649,In_2962);
xor U239 (N_239,In_3709,In_141);
nor U240 (N_240,In_3374,In_3702);
nand U241 (N_241,In_1247,In_3627);
xor U242 (N_242,In_338,In_4316);
nand U243 (N_243,In_4825,In_761);
nand U244 (N_244,In_1681,In_3831);
or U245 (N_245,In_1825,In_1599);
and U246 (N_246,In_1206,In_2589);
nand U247 (N_247,In_1925,In_2196);
or U248 (N_248,In_1409,In_356);
and U249 (N_249,In_3535,In_4954);
or U250 (N_250,In_1170,In_4789);
xnor U251 (N_251,In_2054,In_4116);
nor U252 (N_252,In_418,In_4614);
and U253 (N_253,In_2567,In_3185);
nand U254 (N_254,In_998,In_4024);
xor U255 (N_255,In_3772,In_4029);
nor U256 (N_256,In_397,In_3717);
and U257 (N_257,In_1067,In_342);
xnor U258 (N_258,In_3720,In_3125);
nor U259 (N_259,In_279,In_588);
nor U260 (N_260,In_3962,In_3556);
and U261 (N_261,In_170,In_1992);
nor U262 (N_262,In_2036,In_2771);
nand U263 (N_263,In_3852,In_1864);
nor U264 (N_264,In_4720,In_3014);
nor U265 (N_265,In_2480,In_2704);
nor U266 (N_266,In_4341,In_1038);
nand U267 (N_267,In_1029,In_3030);
nor U268 (N_268,In_1481,In_1059);
nor U269 (N_269,In_2079,In_1283);
nor U270 (N_270,In_1452,In_788);
and U271 (N_271,In_134,In_3677);
nor U272 (N_272,In_3540,In_4905);
nand U273 (N_273,In_776,In_4098);
or U274 (N_274,In_520,In_1548);
and U275 (N_275,In_1533,In_935);
or U276 (N_276,In_2768,In_4848);
xor U277 (N_277,In_4181,In_1326);
nand U278 (N_278,In_3361,In_3353);
nand U279 (N_279,In_1019,In_376);
nor U280 (N_280,In_99,In_3817);
and U281 (N_281,In_3625,In_2820);
or U282 (N_282,In_3163,In_2805);
nor U283 (N_283,In_2151,In_2174);
nor U284 (N_284,In_765,In_250);
or U285 (N_285,In_2379,In_4239);
nand U286 (N_286,In_2937,In_4387);
xor U287 (N_287,In_74,In_4792);
and U288 (N_288,In_455,In_497);
or U289 (N_289,In_3046,In_4390);
nand U290 (N_290,In_1814,In_4125);
nand U291 (N_291,In_2518,In_573);
or U292 (N_292,In_2977,In_4382);
nor U293 (N_293,In_505,In_3157);
nor U294 (N_294,In_1563,In_4106);
or U295 (N_295,In_22,In_1948);
nand U296 (N_296,In_3073,In_3173);
nor U297 (N_297,In_4959,In_1740);
and U298 (N_298,In_671,In_121);
and U299 (N_299,In_4199,In_1763);
xor U300 (N_300,In_3610,In_1882);
or U301 (N_301,In_3716,In_1265);
nor U302 (N_302,In_512,In_1865);
and U303 (N_303,In_251,In_1028);
and U304 (N_304,In_173,In_3107);
xor U305 (N_305,In_3918,In_2656);
xor U306 (N_306,In_4799,In_4940);
or U307 (N_307,In_1430,In_1473);
or U308 (N_308,In_1844,In_3868);
or U309 (N_309,In_1832,In_3850);
or U310 (N_310,In_2624,In_417);
and U311 (N_311,In_2841,In_35);
nor U312 (N_312,In_61,In_4591);
nor U313 (N_313,In_4299,In_2437);
nor U314 (N_314,In_4538,In_1306);
nand U315 (N_315,In_4437,In_4511);
and U316 (N_316,In_511,In_1012);
and U317 (N_317,In_19,In_3590);
nor U318 (N_318,In_2921,In_2000);
and U319 (N_319,In_783,In_1090);
nand U320 (N_320,In_4278,In_4051);
nand U321 (N_321,In_3000,In_1057);
and U322 (N_322,In_4872,In_3384);
or U323 (N_323,In_219,In_2816);
or U324 (N_324,In_1232,In_228);
and U325 (N_325,In_1501,In_4489);
nand U326 (N_326,In_2146,In_204);
nor U327 (N_327,In_374,In_3995);
or U328 (N_328,In_1649,In_2322);
xor U329 (N_329,In_4808,In_2178);
nor U330 (N_330,In_2803,In_2244);
nand U331 (N_331,In_2912,In_1404);
nor U332 (N_332,In_2934,In_1345);
nand U333 (N_333,In_3494,In_822);
or U334 (N_334,In_1155,In_1482);
or U335 (N_335,In_3459,In_3922);
and U336 (N_336,In_1321,In_1444);
or U337 (N_337,In_908,In_3329);
or U338 (N_338,In_3316,In_4681);
nor U339 (N_339,In_3857,In_504);
nand U340 (N_340,In_3,In_1126);
nor U341 (N_341,In_1241,In_814);
or U342 (N_342,In_1086,In_687);
and U343 (N_343,In_1191,In_4997);
nor U344 (N_344,In_4409,In_2052);
xnor U345 (N_345,In_2614,In_1670);
xor U346 (N_346,In_4155,In_883);
nor U347 (N_347,In_738,In_3682);
and U348 (N_348,In_4854,In_1589);
or U349 (N_349,In_2310,In_2213);
and U350 (N_350,In_72,In_2136);
and U351 (N_351,In_4384,In_4920);
nand U352 (N_352,In_829,In_2871);
nor U353 (N_353,In_3049,In_3804);
and U354 (N_354,In_3961,In_1935);
xnor U355 (N_355,In_147,In_1451);
nand U356 (N_356,In_1098,In_402);
nor U357 (N_357,In_4241,In_985);
nand U358 (N_358,In_3624,In_2451);
nand U359 (N_359,In_1797,In_3484);
and U360 (N_360,In_2762,In_4093);
or U361 (N_361,In_3862,In_1855);
nand U362 (N_362,In_2239,In_3947);
xor U363 (N_363,In_1436,In_3997);
xnor U364 (N_364,In_26,In_4504);
nor U365 (N_365,In_127,In_3805);
nor U366 (N_366,In_1107,In_3480);
nand U367 (N_367,In_522,In_3642);
xnor U368 (N_368,In_4294,In_3009);
xnor U369 (N_369,In_4142,In_2431);
and U370 (N_370,In_3277,In_4877);
and U371 (N_371,In_1856,In_740);
nor U372 (N_372,In_2992,In_4112);
nand U373 (N_373,In_4245,In_2017);
nand U374 (N_374,In_2946,In_1957);
nor U375 (N_375,In_1660,In_4611);
or U376 (N_376,In_3877,In_3089);
xor U377 (N_377,In_3929,In_4846);
nor U378 (N_378,In_886,In_2570);
or U379 (N_379,In_1054,In_1689);
and U380 (N_380,In_3331,In_1685);
and U381 (N_381,In_2786,In_4263);
nor U382 (N_382,In_4557,In_2924);
and U383 (N_383,In_1424,In_2377);
xor U384 (N_384,In_2684,In_3803);
nand U385 (N_385,In_3767,In_467);
and U386 (N_386,In_1747,In_655);
or U387 (N_387,In_49,In_3217);
and U388 (N_388,In_1142,In_1734);
or U389 (N_389,In_1391,In_4833);
or U390 (N_390,In_905,In_161);
nor U391 (N_391,In_78,In_3529);
or U392 (N_392,In_4884,In_1791);
or U393 (N_393,In_3136,In_1694);
nor U394 (N_394,In_4201,In_3820);
nor U395 (N_395,In_1091,In_2932);
and U396 (N_396,In_4660,In_3345);
nor U397 (N_397,In_4220,In_757);
or U398 (N_398,In_1407,In_469);
nand U399 (N_399,In_2706,In_1655);
and U400 (N_400,In_955,In_4036);
xnor U401 (N_401,In_628,In_3386);
or U402 (N_402,In_2221,In_3010);
xnor U403 (N_403,In_3482,In_2240);
and U404 (N_404,In_4875,In_632);
and U405 (N_405,In_2192,In_363);
and U406 (N_406,In_4987,In_1792);
and U407 (N_407,In_733,In_1959);
nor U408 (N_408,In_4470,In_1897);
or U409 (N_409,In_1921,In_772);
nand U410 (N_410,In_4134,In_3796);
nand U411 (N_411,In_1399,In_4868);
or U412 (N_412,In_2033,In_1687);
and U413 (N_413,In_4453,In_1524);
and U414 (N_414,In_1162,In_2015);
or U415 (N_415,In_4897,In_1813);
and U416 (N_416,In_2529,In_4371);
nor U417 (N_417,In_3885,In_1354);
and U418 (N_418,In_4910,In_2792);
nor U419 (N_419,In_3524,In_2455);
xor U420 (N_420,In_95,In_192);
and U421 (N_421,In_293,In_1601);
and U422 (N_422,In_1785,In_4418);
nor U423 (N_423,In_1159,In_3793);
nand U424 (N_424,In_3132,In_1755);
and U425 (N_425,In_1584,In_1175);
nor U426 (N_426,In_4007,In_2246);
xor U427 (N_427,In_797,In_2847);
or U428 (N_428,In_3387,In_1072);
or U429 (N_429,In_120,In_1918);
nand U430 (N_430,In_3253,In_3668);
and U431 (N_431,In_100,In_4275);
or U432 (N_432,In_3770,In_835);
nand U433 (N_433,In_2565,In_970);
or U434 (N_434,In_1671,In_3972);
or U435 (N_435,In_4658,In_3628);
nor U436 (N_436,In_3244,In_562);
nand U437 (N_437,In_3640,In_2520);
and U438 (N_438,In_3218,In_2095);
or U439 (N_439,In_3120,In_264);
xor U440 (N_440,In_4812,In_2628);
and U441 (N_441,In_3898,In_3810);
and U442 (N_442,In_2961,In_2398);
and U443 (N_443,In_3110,In_4031);
and U444 (N_444,In_4529,In_1303);
and U445 (N_445,In_4841,In_2444);
xor U446 (N_446,In_3641,In_433);
nand U447 (N_447,In_3174,In_3571);
nand U448 (N_448,In_75,In_1919);
xor U449 (N_449,In_4669,In_4824);
nor U450 (N_450,In_370,In_2220);
xor U451 (N_451,In_960,In_4756);
nand U452 (N_452,In_2394,In_2479);
nand U453 (N_453,In_4561,In_2972);
nand U454 (N_454,In_2641,In_2559);
or U455 (N_455,In_3661,In_680);
nand U456 (N_456,In_850,In_3166);
and U457 (N_457,In_851,In_537);
and U458 (N_458,In_427,In_386);
nor U459 (N_459,In_1330,In_3637);
and U460 (N_460,In_1275,In_3982);
or U461 (N_461,In_979,In_3974);
and U462 (N_462,In_3956,In_2157);
and U463 (N_463,In_2974,In_4865);
xor U464 (N_464,In_3076,In_1828);
nor U465 (N_465,In_3178,In_3220);
nand U466 (N_466,In_1393,In_215);
nor U467 (N_467,In_3563,In_2023);
xnor U468 (N_468,In_1783,In_495);
nand U469 (N_469,In_3269,In_411);
and U470 (N_470,In_1417,In_1885);
or U471 (N_471,In_1423,In_4852);
and U472 (N_472,In_2963,In_4531);
nor U473 (N_473,In_4535,In_360);
and U474 (N_474,In_493,In_4314);
or U475 (N_475,In_2836,In_3029);
nor U476 (N_476,In_1106,In_2269);
nand U477 (N_477,In_4795,In_2920);
or U478 (N_478,In_2223,In_2736);
or U479 (N_479,In_296,In_294);
nor U480 (N_480,In_371,In_4878);
or U481 (N_481,In_918,In_4207);
nor U482 (N_482,In_2898,In_4640);
and U483 (N_483,In_4968,In_1214);
and U484 (N_484,In_1217,In_2609);
or U485 (N_485,In_1138,In_904);
or U486 (N_486,In_216,In_569);
or U487 (N_487,In_4436,In_1427);
nand U488 (N_488,In_3235,In_3195);
nand U489 (N_489,In_3342,In_2553);
xnor U490 (N_490,In_2533,In_976);
xor U491 (N_491,In_1525,In_4132);
nor U492 (N_492,In_2519,In_1408);
or U493 (N_493,In_1812,In_1731);
and U494 (N_494,In_1757,In_1429);
or U495 (N_495,In_2367,In_2276);
or U496 (N_496,In_1811,In_3156);
or U497 (N_497,In_891,In_4649);
xnor U498 (N_498,In_2238,In_575);
nand U499 (N_499,In_2640,In_1820);
nor U500 (N_500,In_4482,In_3408);
and U501 (N_501,In_4908,In_3613);
or U502 (N_502,In_4564,In_4879);
nand U503 (N_503,In_1325,In_3519);
xnor U504 (N_504,In_389,In_3490);
and U505 (N_505,In_2901,In_1353);
xnor U506 (N_506,In_3901,In_2384);
and U507 (N_507,In_3093,In_4683);
nand U508 (N_508,In_2257,In_3520);
and U509 (N_509,In_845,In_2425);
or U510 (N_510,In_2463,In_3028);
xnor U511 (N_511,In_3855,In_4972);
nand U512 (N_512,In_2008,In_2167);
nor U513 (N_513,In_1389,In_4617);
nand U514 (N_514,In_358,In_1195);
nor U515 (N_515,In_4632,In_3609);
or U516 (N_516,In_1566,In_4934);
xor U517 (N_517,In_2025,In_4659);
xor U518 (N_518,In_688,In_2184);
and U519 (N_519,In_1973,In_574);
nor U520 (N_520,In_3565,In_1002);
nand U521 (N_521,In_4027,In_254);
nand U522 (N_522,In_1026,In_2094);
xnor U523 (N_523,In_700,In_1901);
nand U524 (N_524,In_4266,In_3151);
nand U525 (N_525,In_2719,In_1684);
xnor U526 (N_526,In_1706,In_4474);
nand U527 (N_527,In_82,In_2042);
nand U528 (N_528,In_3088,In_2561);
or U529 (N_529,In_4694,In_150);
nor U530 (N_530,In_3394,In_3414);
nand U531 (N_531,In_782,In_853);
or U532 (N_532,In_2083,In_2688);
or U533 (N_533,In_1956,In_2193);
or U534 (N_534,In_1021,In_893);
nor U535 (N_535,In_2524,In_777);
or U536 (N_536,In_2552,In_3692);
or U537 (N_537,In_2272,In_2675);
or U538 (N_538,In_956,In_1889);
and U539 (N_539,In_102,In_3300);
nand U540 (N_540,In_4601,In_2317);
nand U541 (N_541,In_1245,In_306);
or U542 (N_542,In_3900,In_952);
xor U543 (N_543,In_2916,In_1023);
xnor U544 (N_544,In_3614,In_807);
nor U545 (N_545,In_1818,In_3271);
xor U546 (N_546,In_4766,In_4661);
nand U547 (N_547,In_4546,In_1768);
nand U548 (N_548,In_1967,In_1236);
nor U549 (N_549,In_1531,In_3504);
or U550 (N_550,In_1603,In_2572);
nand U551 (N_551,In_459,In_2484);
xor U552 (N_552,In_1558,In_4237);
nand U553 (N_553,In_2056,In_1318);
xnor U554 (N_554,In_2128,In_2702);
nand U555 (N_555,In_1215,In_1633);
xor U556 (N_556,In_1461,In_333);
nand U557 (N_557,In_1709,In_2540);
or U558 (N_558,In_2225,In_3708);
and U559 (N_559,In_3889,In_4308);
nor U560 (N_560,In_4495,In_90);
nand U561 (N_561,In_4702,In_1380);
nor U562 (N_562,In_794,In_1725);
and U563 (N_563,In_1103,In_3577);
nand U564 (N_564,In_3809,In_2513);
nand U565 (N_565,In_3154,In_3434);
and U566 (N_566,In_4405,In_1977);
nor U567 (N_567,In_4404,In_3936);
or U568 (N_568,In_530,In_3240);
and U569 (N_569,In_4343,In_3026);
nor U570 (N_570,In_4590,In_276);
xor U571 (N_571,In_686,In_4376);
nand U572 (N_572,In_4685,In_4952);
or U573 (N_573,In_667,In_4779);
nor U574 (N_574,In_3420,In_2564);
xor U575 (N_575,In_4942,In_2148);
and U576 (N_576,In_2996,In_3388);
and U577 (N_577,In_4012,In_4050);
or U578 (N_578,In_4565,In_4610);
nor U579 (N_579,In_1628,In_1036);
and U580 (N_580,In_531,In_226);
nand U581 (N_581,In_2228,In_3359);
xor U582 (N_582,In_848,In_3367);
and U583 (N_583,In_4784,In_1981);
nor U584 (N_584,In_1133,In_2517);
nand U585 (N_585,In_2417,In_4113);
and U586 (N_586,In_4457,In_4510);
or U587 (N_587,In_2305,In_2689);
nand U588 (N_588,In_3672,In_1165);
nor U589 (N_589,In_4216,In_2181);
xnor U590 (N_590,In_1798,In_2899);
nand U591 (N_591,In_2573,In_369);
xnor U592 (N_592,In_1402,In_615);
xnor U593 (N_593,In_4810,In_3312);
nor U594 (N_594,In_4486,In_2777);
or U595 (N_595,In_448,In_2154);
and U596 (N_596,In_1610,In_1432);
nand U597 (N_597,In_2735,In_4057);
nor U598 (N_598,In_325,In_2860);
nand U599 (N_599,In_1717,In_2511);
nor U600 (N_600,In_4149,In_3293);
nor U601 (N_601,In_726,In_4227);
or U602 (N_602,In_4301,In_4708);
nor U603 (N_603,In_3558,In_2569);
or U604 (N_604,In_273,In_662);
nor U605 (N_605,In_864,In_1535);
nand U606 (N_606,In_1200,In_4560);
or U607 (N_607,In_1105,In_4243);
or U608 (N_608,In_4709,In_4337);
nand U609 (N_609,In_3378,In_3605);
nand U610 (N_610,In_2818,In_652);
nor U611 (N_611,In_329,In_332);
or U612 (N_612,In_3274,In_4566);
and U613 (N_613,In_2405,In_4331);
xnor U614 (N_614,In_372,In_4876);
nor U615 (N_615,In_1377,In_2997);
nand U616 (N_616,In_4804,In_2986);
and U617 (N_617,In_13,In_3410);
nor U618 (N_618,In_1068,In_824);
and U619 (N_619,In_2875,In_4076);
xnor U620 (N_620,In_1004,In_2772);
nand U621 (N_621,In_3048,In_3575);
nor U622 (N_622,In_2163,In_4580);
or U623 (N_623,In_1189,In_3680);
nand U624 (N_624,In_1697,In_2829);
nand U625 (N_625,In_3542,In_4458);
and U626 (N_626,In_1772,In_838);
and U627 (N_627,In_200,In_2823);
and U628 (N_628,In_3828,In_3486);
nor U629 (N_629,In_1373,In_499);
or U630 (N_630,In_335,In_3392);
xnor U631 (N_631,In_4762,In_3920);
or U632 (N_632,In_2085,In_560);
xnor U633 (N_633,In_4224,In_2826);
and U634 (N_634,In_3572,In_142);
nor U635 (N_635,In_1723,In_4999);
nor U636 (N_636,In_3501,In_1372);
nand U637 (N_637,In_4161,In_2800);
nor U638 (N_638,In_2863,In_4375);
nand U639 (N_639,In_940,In_4500);
and U640 (N_640,In_3074,In_4180);
or U641 (N_641,In_3870,In_3618);
or U642 (N_642,In_4618,In_2231);
xnor U643 (N_643,In_890,In_203);
nand U644 (N_644,In_2030,In_2053);
and U645 (N_645,In_4070,In_1940);
nor U646 (N_646,In_3396,In_3811);
nor U647 (N_647,In_832,In_4269);
xnor U648 (N_648,In_3899,In_4209);
or U649 (N_649,In_2376,In_354);
and U650 (N_650,In_1622,In_4330);
xnor U651 (N_651,In_34,In_817);
and U652 (N_652,In_4912,In_242);
and U653 (N_653,In_2280,In_4200);
nor U654 (N_654,In_4911,In_4479);
nor U655 (N_655,In_1841,In_3999);
nor U656 (N_656,In_30,In_380);
or U657 (N_657,In_4575,In_4533);
or U658 (N_658,In_130,In_4700);
and U659 (N_659,In_808,In_4352);
xor U660 (N_660,In_3114,In_2006);
and U661 (N_661,In_1963,In_4396);
nand U662 (N_662,In_4988,In_184);
nor U663 (N_663,In_3700,In_2655);
nand U664 (N_664,In_2319,In_4802);
xnor U665 (N_665,In_2399,In_1210);
nand U666 (N_666,In_3123,In_2633);
nor U667 (N_667,In_145,In_3884);
xor U668 (N_668,In_3925,In_713);
nor U669 (N_669,In_1580,In_2576);
and U670 (N_670,In_3443,In_758);
xor U671 (N_671,In_4431,In_4675);
or U672 (N_672,In_4927,In_4206);
or U673 (N_673,In_4283,In_1128);
xor U674 (N_674,In_1860,In_4736);
nor U675 (N_675,In_1616,In_255);
nand U676 (N_676,In_157,In_3798);
xor U677 (N_677,In_185,In_666);
and U678 (N_678,In_2421,In_3493);
nand U679 (N_679,In_1808,In_2595);
nand U680 (N_680,In_3807,In_1721);
and U681 (N_681,In_4715,In_983);
xnor U682 (N_682,In_4813,In_1800);
nor U683 (N_683,In_4230,In_4515);
or U684 (N_684,In_2074,In_2440);
nor U685 (N_685,In_2432,In_1198);
and U686 (N_686,In_924,In_1095);
nor U687 (N_687,In_2619,In_4791);
nor U688 (N_688,In_207,In_1137);
nor U689 (N_689,In_1459,In_4122);
nor U690 (N_690,In_2169,In_4052);
and U691 (N_691,In_1569,In_4129);
or U692 (N_692,In_3799,In_2681);
nor U693 (N_693,In_3254,In_897);
nand U694 (N_694,In_3090,In_4300);
nor U695 (N_695,In_88,In_3215);
nor U696 (N_696,In_3497,In_18);
nand U697 (N_697,In_2794,In_1400);
or U698 (N_698,In_1930,In_3349);
nor U699 (N_699,In_4123,In_1212);
and U700 (N_700,In_968,In_939);
or U701 (N_701,In_2216,In_866);
or U702 (N_702,In_3083,In_381);
xnor U703 (N_703,In_3646,In_1996);
xor U704 (N_704,In_936,In_1109);
xnor U705 (N_705,In_2232,In_823);
nand U706 (N_706,In_262,In_2371);
xnor U707 (N_707,In_361,In_4008);
and U708 (N_708,In_4109,In_1833);
nor U709 (N_709,In_1146,In_2830);
nor U710 (N_710,In_1712,In_1337);
nor U711 (N_711,In_2330,In_4061);
and U712 (N_712,In_2236,In_4395);
xnor U713 (N_713,In_4842,In_4062);
nand U714 (N_714,In_679,In_458);
and U715 (N_715,In_4088,In_2212);
nand U716 (N_716,In_4537,In_3315);
and U717 (N_717,In_4748,In_2959);
xnor U718 (N_718,In_1457,In_1688);
or U719 (N_719,In_2683,In_2262);
nor U720 (N_720,In_473,In_900);
xor U721 (N_721,In_113,In_3533);
xor U722 (N_722,In_2542,In_3778);
nor U723 (N_723,In_1253,In_4329);
or U724 (N_724,In_2009,In_735);
or U725 (N_725,In_1139,In_731);
or U726 (N_726,In_2938,In_195);
xor U727 (N_727,In_996,In_1896);
xor U728 (N_728,In_4797,In_2004);
xor U729 (N_729,In_313,In_3986);
and U730 (N_730,In_165,In_4357);
or U731 (N_731,In_2855,In_532);
or U732 (N_732,In_4612,In_4423);
nand U733 (N_733,In_2654,In_4090);
nor U734 (N_734,In_4697,In_1031);
or U735 (N_735,In_1547,In_345);
and U736 (N_736,In_305,In_65);
and U737 (N_737,In_1559,In_4171);
or U738 (N_738,In_619,In_3715);
or U739 (N_739,In_3103,In_4484);
nand U740 (N_740,In_3644,In_357);
xor U741 (N_741,In_3404,In_2814);
xor U742 (N_742,In_3018,In_373);
nand U743 (N_743,In_4187,In_1225);
and U744 (N_744,In_1779,In_445);
xnor U745 (N_745,In_2325,In_2098);
or U746 (N_746,In_1268,In_3383);
and U747 (N_747,In_2112,In_3021);
and U748 (N_748,In_1264,In_2264);
nand U749 (N_749,In_3562,In_2604);
nor U750 (N_750,In_4407,In_1780);
nor U751 (N_751,In_4728,In_1390);
or U752 (N_752,In_4831,In_3522);
nor U753 (N_753,In_4576,In_1907);
xnor U754 (N_754,In_4277,In_576);
nor U755 (N_755,In_1490,In_3814);
nor U756 (N_756,In_3229,In_1928);
or U757 (N_757,In_3044,In_4713);
nor U758 (N_758,In_3588,In_1528);
xor U759 (N_759,In_2316,In_3741);
or U760 (N_760,In_4214,In_2072);
or U761 (N_761,In_4830,In_4656);
and U762 (N_762,In_4555,In_4290);
or U763 (N_763,In_2208,In_501);
and U764 (N_764,In_3916,In_2477);
nand U765 (N_765,In_4353,In_2669);
xnor U766 (N_766,In_2798,In_3366);
xnor U767 (N_767,In_2019,In_58);
or U768 (N_768,In_1770,In_3639);
or U769 (N_769,In_1317,In_3508);
or U770 (N_770,In_568,In_2092);
xor U771 (N_771,In_4252,In_2648);
or U772 (N_772,In_2195,In_2523);
or U773 (N_773,In_4723,In_2326);
xnor U774 (N_774,In_3438,In_1504);
or U775 (N_775,In_2883,In_3225);
or U776 (N_776,In_1131,In_3467);
or U777 (N_777,In_561,In_3979);
nand U778 (N_778,In_3905,In_3451);
xor U779 (N_779,In_4491,In_799);
nor U780 (N_780,In_4127,In_4054);
nand U781 (N_781,In_263,In_3591);
nor U782 (N_782,In_536,In_2423);
xnor U783 (N_783,In_2179,In_240);
nor U784 (N_784,In_1756,In_1190);
and U785 (N_785,In_1594,In_4446);
xnor U786 (N_786,In_36,In_366);
nand U787 (N_787,In_4962,In_1152);
and U788 (N_788,In_806,In_425);
or U789 (N_789,In_62,In_1016);
nand U790 (N_790,In_3039,In_421);
nor U791 (N_791,In_128,In_1344);
nor U792 (N_792,In_3525,In_2488);
and U793 (N_793,In_862,In_2925);
nor U794 (N_794,In_300,In_3883);
and U795 (N_795,In_409,In_4430);
nand U796 (N_796,In_4347,In_3045);
and U797 (N_797,In_4361,In_3745);
and U798 (N_798,In_1946,In_3612);
and U799 (N_799,In_875,In_3854);
and U800 (N_800,In_2415,In_2029);
and U801 (N_801,In_1479,In_3481);
and U802 (N_802,In_1110,In_4344);
and U803 (N_803,In_4749,In_1862);
nor U804 (N_804,In_2252,In_4229);
xor U805 (N_805,In_139,In_1485);
xor U806 (N_806,In_1279,In_1073);
nand U807 (N_807,In_4803,In_4643);
nand U808 (N_808,In_4888,In_4536);
nor U809 (N_809,In_2661,In_1017);
and U810 (N_810,In_234,In_438);
nand U811 (N_811,In_4434,In_1499);
nand U812 (N_812,In_2386,In_3304);
or U813 (N_813,In_2759,In_1185);
nand U814 (N_814,In_3409,In_3204);
xor U815 (N_815,In_2744,In_872);
or U816 (N_816,In_3800,In_3036);
nor U817 (N_817,In_1238,In_4179);
and U818 (N_818,In_4860,In_4271);
and U819 (N_819,In_3261,In_2082);
or U820 (N_820,In_1064,In_1842);
nand U821 (N_821,In_3777,In_2265);
nor U822 (N_822,In_826,In_3430);
or U823 (N_823,In_2311,In_4288);
and U824 (N_824,In_1312,In_2577);
xnor U825 (N_825,In_2370,In_1984);
or U826 (N_826,In_624,In_793);
or U827 (N_827,In_1604,In_1136);
nor U828 (N_828,In_416,In_2738);
and U829 (N_829,In_269,In_67);
nor U830 (N_830,In_594,In_4483);
xor U831 (N_831,In_1256,In_1553);
nor U832 (N_832,In_830,In_4585);
or U833 (N_833,In_3147,In_4293);
nor U834 (N_834,In_4130,In_950);
xnor U835 (N_835,In_3072,In_2349);
and U836 (N_836,In_2958,In_3580);
nor U837 (N_837,In_2866,In_4903);
nor U838 (N_838,In_3500,In_1962);
and U839 (N_839,In_1102,In_1007);
xnor U840 (N_840,In_1169,In_4609);
and U841 (N_841,In_2964,In_2427);
xor U842 (N_842,In_2383,In_513);
nand U843 (N_843,In_2452,In_2635);
and U844 (N_844,In_2496,In_2560);
nand U845 (N_845,In_2287,In_426);
and U846 (N_846,In_1421,In_1425);
nand U847 (N_847,In_590,In_1874);
nand U848 (N_848,In_2312,In_3849);
or U849 (N_849,In_791,In_564);
nor U850 (N_850,In_4806,In_1053);
nor U851 (N_851,In_1507,In_1536);
xor U852 (N_852,In_155,In_3611);
xor U853 (N_853,In_1658,In_4670);
nand U854 (N_854,In_675,In_2617);
xor U855 (N_855,In_1088,In_4798);
nand U856 (N_856,In_41,In_3431);
xnor U857 (N_857,In_3418,In_516);
nand U858 (N_858,In_3873,In_3714);
nand U859 (N_859,In_597,In_3209);
xnor U860 (N_860,In_3053,In_2502);
or U861 (N_861,In_1796,In_3768);
nor U862 (N_862,In_387,In_3437);
nor U863 (N_863,In_1704,In_3517);
xnor U864 (N_864,In_2580,In_1732);
nand U865 (N_865,In_3907,In_106);
or U866 (N_866,In_3227,In_3025);
nor U867 (N_867,In_1348,In_3284);
or U868 (N_868,In_2435,In_633);
and U869 (N_869,In_498,In_1445);
xnor U870 (N_870,In_4420,In_648);
xor U871 (N_871,In_4467,In_1497);
or U872 (N_872,In_2294,In_1726);
or U873 (N_873,In_3783,In_439);
or U874 (N_874,In_4828,In_1233);
nor U875 (N_875,In_664,In_3600);
or U876 (N_876,In_2668,In_2359);
or U877 (N_877,In_1983,In_3511);
nor U878 (N_878,In_855,In_3129);
nor U879 (N_879,In_611,In_4953);
xor U880 (N_880,In_1551,In_1693);
and U881 (N_881,In_1115,In_4823);
nor U882 (N_882,In_638,In_1388);
nand U883 (N_883,In_1192,In_4960);
xor U884 (N_884,In_3673,In_2155);
and U885 (N_885,In_1149,In_4742);
and U886 (N_886,In_1519,In_2073);
nand U887 (N_887,In_860,In_3439);
nand U888 (N_888,In_3670,In_3007);
nor U889 (N_889,In_488,In_2481);
and U890 (N_890,In_2894,In_1331);
nand U891 (N_891,In_3035,In_3528);
and U892 (N_892,In_3774,In_4001);
xor U893 (N_893,In_697,In_1381);
and U894 (N_894,In_3466,In_3941);
nand U895 (N_895,In_3606,In_190);
and U896 (N_896,In_1900,In_2301);
and U897 (N_897,In_4444,In_800);
and U898 (N_898,In_3179,In_2039);
nor U899 (N_899,In_2428,In_4677);
xor U900 (N_900,In_3057,In_4587);
and U901 (N_901,In_795,In_1834);
nand U902 (N_902,In_748,In_4793);
or U903 (N_903,In_2791,In_2672);
nor U904 (N_904,In_3063,In_232);
nor U905 (N_905,In_3896,In_1647);
nor U906 (N_906,In_691,In_4718);
or U907 (N_907,In_2699,In_4095);
or U908 (N_908,In_3743,In_3080);
or U909 (N_909,In_3688,In_148);
xor U910 (N_910,In_171,In_2587);
and U911 (N_911,In_1512,In_2717);
xnor U912 (N_912,In_515,In_1252);
xor U913 (N_913,In_167,In_2903);
and U914 (N_914,In_965,In_1539);
nor U915 (N_915,In_1188,In_1966);
xor U916 (N_916,In_4205,In_3303);
and U917 (N_917,In_4957,In_214);
and U918 (N_918,In_4577,In_3267);
nor U919 (N_919,In_337,In_3311);
or U920 (N_920,In_4099,In_4862);
and U921 (N_921,In_1866,In_4251);
nor U922 (N_922,In_3584,In_400);
or U923 (N_923,In_4397,In_3578);
or U924 (N_924,In_3196,In_3695);
xnor U925 (N_925,In_4391,In_1867);
xor U926 (N_926,In_3546,In_2393);
nand U927 (N_927,In_1952,In_3450);
nand U928 (N_928,In_1509,In_1466);
and U929 (N_929,In_4248,In_4916);
xnor U930 (N_930,In_2872,In_4559);
nand U931 (N_931,In_4764,In_4185);
xor U932 (N_932,In_3054,In_432);
nand U933 (N_933,In_3247,In_1908);
nor U934 (N_934,In_645,In_4768);
or U935 (N_935,In_3874,In_2957);
nand U936 (N_936,In_1701,In_623);
xnor U937 (N_937,In_3515,In_736);
and U938 (N_938,In_3696,In_3823);
or U939 (N_939,In_3955,In_3966);
and U940 (N_940,In_1789,In_3752);
and U941 (N_941,In_4366,In_4849);
or U942 (N_942,In_676,In_2474);
xor U943 (N_943,In_3718,In_3314);
xor U944 (N_944,In_1340,In_2162);
nand U945 (N_945,In_4989,In_4983);
and U946 (N_946,In_931,In_4388);
nor U947 (N_947,In_4426,In_819);
nor U948 (N_948,In_3432,In_2271);
or U949 (N_949,In_4014,In_1741);
and U950 (N_950,In_526,In_3645);
and U951 (N_951,In_1985,In_3336);
or U952 (N_952,In_1018,In_3880);
nand U953 (N_953,In_975,In_1877);
or U954 (N_954,In_3290,In_2802);
and U955 (N_955,In_1458,In_3794);
nand U956 (N_956,In_3721,In_4324);
or U957 (N_957,In_1912,In_2598);
nor U958 (N_958,In_3917,In_1244);
xnor U959 (N_959,In_2837,In_2068);
nand U960 (N_960,In_804,In_4259);
and U961 (N_961,In_4809,In_2209);
or U962 (N_962,In_3536,In_218);
nand U963 (N_963,In_3681,In_1498);
and U964 (N_964,In_4368,In_4589);
or U965 (N_965,In_2409,In_3298);
nand U966 (N_966,In_1135,In_2881);
nand U967 (N_967,In_3008,In_4218);
or U968 (N_968,In_54,In_1767);
nand U969 (N_969,In_172,In_3626);
nand U970 (N_970,In_730,In_1554);
nor U971 (N_971,In_4053,In_2309);
xnor U972 (N_972,In_327,In_462);
nor U973 (N_973,In_3457,In_1151);
and U974 (N_974,In_1699,In_556);
nand U975 (N_975,In_4507,In_4755);
nor U976 (N_976,In_4183,In_2724);
nand U977 (N_977,In_4165,In_3294);
xor U978 (N_978,In_4448,In_1651);
nand U979 (N_979,In_1242,In_328);
or U980 (N_980,In_1617,In_2947);
xor U981 (N_981,In_3015,In_973);
or U982 (N_982,In_2991,In_3994);
xnor U983 (N_983,In_750,In_3231);
nand U984 (N_984,In_856,In_942);
or U985 (N_985,In_1148,In_2979);
and U986 (N_986,In_422,In_2622);
or U987 (N_987,In_2734,In_4815);
or U988 (N_988,In_4373,In_324);
nor U989 (N_989,In_1583,In_827);
or U990 (N_990,In_3737,In_83);
xor U991 (N_991,In_122,In_440);
and U992 (N_992,In_698,In_787);
nor U993 (N_993,In_3214,In_4232);
and U994 (N_994,In_3938,In_3499);
nand U995 (N_995,In_710,In_1119);
nor U996 (N_996,In_1394,In_1537);
or U997 (N_997,In_4235,In_4398);
xnor U998 (N_998,In_1270,In_3330);
nor U999 (N_999,In_474,In_3859);
or U1000 (N_1000,In_4077,In_1961);
and U1001 (N_1001,In_4210,In_1953);
or U1002 (N_1002,In_2202,In_2887);
nor U1003 (N_1003,In_3818,In_3570);
or U1004 (N_1004,In_316,In_1654);
and U1005 (N_1005,In_3541,In_4440);
and U1006 (N_1006,In_1209,In_4152);
nand U1007 (N_1007,In_1183,In_3784);
nand U1008 (N_1008,In_4551,In_3756);
nor U1009 (N_1009,In_4003,In_3335);
xnor U1010 (N_1010,In_2133,In_3140);
nor U1011 (N_1011,In_1782,In_626);
xor U1012 (N_1012,In_2188,In_643);
nand U1013 (N_1013,In_3327,In_334);
and U1014 (N_1014,In_2878,In_4945);
nor U1015 (N_1015,In_1989,In_482);
nand U1016 (N_1016,In_349,In_2365);
and U1017 (N_1017,In_1526,In_3011);
or U1018 (N_1018,In_1164,In_721);
xor U1019 (N_1019,In_2501,In_2433);
nand U1020 (N_1020,In_140,In_1636);
or U1021 (N_1021,In_2099,In_256);
nand U1022 (N_1022,In_2950,In_4763);
xor U1023 (N_1023,In_2763,In_4717);
or U1024 (N_1024,In_4380,In_2368);
or U1025 (N_1025,In_4620,In_651);
nand U1026 (N_1026,In_4674,In_429);
or U1027 (N_1027,In_725,In_4783);
xnor U1028 (N_1028,In_1905,In_4692);
nor U1029 (N_1029,In_3211,In_4772);
nor U1030 (N_1030,In_2579,In_4586);
xnor U1031 (N_1031,In_558,In_4193);
and U1032 (N_1032,In_1116,In_3333);
xor U1033 (N_1033,In_2637,In_4383);
and U1034 (N_1034,In_1805,In_1255);
nand U1035 (N_1035,In_3219,In_1285);
nor U1036 (N_1036,In_181,In_1034);
or U1037 (N_1037,In_4751,In_1565);
and U1038 (N_1038,In_237,In_2933);
and U1039 (N_1039,In_2801,In_4410);
or U1040 (N_1040,In_4040,In_3324);
nand U1041 (N_1041,In_3621,In_4065);
or U1042 (N_1042,In_4969,In_625);
xnor U1043 (N_1043,In_4948,In_3391);
xnor U1044 (N_1044,In_4909,In_4653);
or U1045 (N_1045,In_4733,In_4228);
and U1046 (N_1046,In_1083,In_2251);
nor U1047 (N_1047,In_199,In_957);
nand U1048 (N_1048,In_868,In_4758);
nor U1049 (N_1049,In_3732,In_4734);
xor U1050 (N_1050,In_2250,In_3643);
or U1051 (N_1051,In_2808,In_4986);
and U1052 (N_1052,In_4874,In_4498);
nor U1053 (N_1053,In_1705,In_2534);
nand U1054 (N_1054,In_3521,In_2670);
or U1055 (N_1055,In_15,In_2969);
xor U1056 (N_1056,In_992,In_4732);
nor U1057 (N_1057,In_1125,In_1802);
or U1058 (N_1058,In_2013,In_3594);
or U1059 (N_1059,In_441,In_4516);
nand U1060 (N_1060,In_1510,In_2339);
xnor U1061 (N_1061,In_4083,In_3701);
nand U1062 (N_1062,In_2016,In_2387);
nand U1063 (N_1063,In_3750,In_3212);
xor U1064 (N_1064,In_2404,In_3150);
and U1065 (N_1065,In_1163,In_4157);
nor U1066 (N_1066,In_820,In_3020);
xor U1067 (N_1067,In_3864,In_1363);
xor U1068 (N_1068,In_3731,In_3530);
xnor U1069 (N_1069,In_1114,In_2971);
xor U1070 (N_1070,In_4477,In_629);
and U1071 (N_1071,In_1753,In_3067);
xor U1072 (N_1072,In_1761,In_4894);
nor U1073 (N_1073,In_2254,In_3738);
nor U1074 (N_1074,In_2782,In_2929);
or U1075 (N_1075,In_1562,In_4899);
and U1076 (N_1076,In_2334,In_3358);
nand U1077 (N_1077,In_1991,In_3260);
xnor U1078 (N_1078,In_4698,In_653);
or U1079 (N_1079,In_4105,In_3633);
nor U1080 (N_1080,In_4322,In_25);
nand U1081 (N_1081,In_1801,In_3808);
nor U1082 (N_1082,In_3207,In_3766);
or U1083 (N_1083,In_2955,In_3739);
nand U1084 (N_1084,In_4226,In_2845);
and U1085 (N_1085,In_1227,In_4128);
nor U1086 (N_1086,In_4056,In_93);
or U1087 (N_1087,In_3503,In_1508);
or U1088 (N_1088,In_683,In_4488);
nor U1089 (N_1089,In_347,In_2418);
and U1090 (N_1090,In_3473,In_3318);
nand U1091 (N_1091,In_678,In_2273);
xor U1092 (N_1092,In_919,In_689);
or U1093 (N_1093,In_768,In_589);
nand U1094 (N_1094,In_2288,In_1254);
xor U1095 (N_1095,In_1112,In_3485);
nor U1096 (N_1096,In_2773,In_4191);
nand U1097 (N_1097,In_4296,In_3657);
nor U1098 (N_1098,In_2692,In_3061);
and U1099 (N_1099,In_3141,In_4258);
nand U1100 (N_1100,In_4,In_2419);
nor U1101 (N_1101,In_288,In_68);
nand U1102 (N_1102,In_43,In_1871);
or U1103 (N_1103,In_751,In_51);
xnor U1104 (N_1104,In_3753,In_3094);
nand U1105 (N_1105,In_2468,In_3676);
nand U1106 (N_1106,In_2140,In_69);
xnor U1107 (N_1107,In_4246,In_1840);
or U1108 (N_1108,In_1968,In_1850);
nand U1109 (N_1109,In_2356,In_4148);
nor U1110 (N_1110,In_4321,In_1894);
or U1111 (N_1111,In_640,In_3617);
xnor U1112 (N_1112,In_2115,In_2900);
nor U1113 (N_1113,In_8,In_2040);
and U1114 (N_1114,In_3650,In_3638);
nor U1115 (N_1115,In_4111,In_3498);
nand U1116 (N_1116,In_4438,In_3763);
nor U1117 (N_1117,In_1683,In_351);
nor U1118 (N_1118,In_2478,In_2106);
and U1119 (N_1119,In_3245,In_892);
and U1120 (N_1120,In_4857,In_364);
or U1121 (N_1121,In_4389,In_3016);
or U1122 (N_1122,In_3990,In_2176);
nor U1123 (N_1123,In_2693,In_771);
nand U1124 (N_1124,In_3910,In_1650);
nor U1125 (N_1125,In_3690,In_3923);
nor U1126 (N_1126,In_4861,In_510);
or U1127 (N_1127,In_1117,In_435);
nand U1128 (N_1128,In_84,In_4552);
nor U1129 (N_1129,In_815,In_4471);
and U1130 (N_1130,In_4540,In_431);
and U1131 (N_1131,In_3713,In_1614);
nand U1132 (N_1132,In_3116,In_3559);
xnor U1133 (N_1133,In_1606,In_2296);
or U1134 (N_1134,In_2438,In_913);
xor U1135 (N_1135,In_2191,In_4520);
or U1136 (N_1136,In_1434,In_4967);
nand U1137 (N_1137,In_2797,In_2941);
nand U1138 (N_1138,In_3423,In_2361);
nand U1139 (N_1139,In_2512,In_4724);
nand U1140 (N_1140,In_1938,In_2543);
xnor U1141 (N_1141,In_4298,In_3636);
and U1142 (N_1142,In_2995,In_3980);
and U1143 (N_1143,In_1435,In_44);
or U1144 (N_1144,In_1488,In_1308);
xnor U1145 (N_1145,In_1274,In_1301);
xnor U1146 (N_1146,In_1576,In_4737);
nand U1147 (N_1147,In_540,In_2058);
nand U1148 (N_1148,In_2795,In_1513);
and U1149 (N_1149,In_2541,In_2263);
nor U1150 (N_1150,In_2858,In_3965);
xor U1151 (N_1151,In_870,In_737);
xor U1152 (N_1152,In_586,In_4950);
and U1153 (N_1153,In_4196,In_1561);
or U1154 (N_1154,In_138,In_1643);
and U1155 (N_1155,In_3263,In_3256);
xnor U1156 (N_1156,In_2722,In_1824);
or U1157 (N_1157,In_1746,In_217);
xnor U1158 (N_1158,In_3478,In_3276);
xor U1159 (N_1159,In_2880,In_1817);
or U1160 (N_1160,In_3927,In_3262);
and U1161 (N_1161,In_3848,In_4042);
nand U1162 (N_1162,In_4339,In_4451);
nor U1163 (N_1163,In_2625,In_3471);
and U1164 (N_1164,In_2984,In_1932);
nand U1165 (N_1165,In_1846,In_1538);
xor U1166 (N_1166,In_744,In_4926);
nand U1167 (N_1167,In_1483,In_898);
and U1168 (N_1168,In_1595,In_2021);
xor U1169 (N_1169,In_261,In_3555);
nand U1170 (N_1170,In_3760,In_2528);
or U1171 (N_1171,In_1474,In_3704);
and U1172 (N_1172,In_4680,In_2746);
or U1173 (N_1173,In_2966,In_567);
nor U1174 (N_1174,In_2575,In_1374);
xor U1175 (N_1175,In_4837,In_2214);
nand U1176 (N_1176,In_4729,In_882);
xnor U1177 (N_1177,In_1631,In_3912);
nand U1178 (N_1178,In_984,In_4786);
xnor U1179 (N_1179,In_821,In_2705);
nand U1180 (N_1180,In_249,In_796);
nor U1181 (N_1181,In_4705,In_3186);
or U1182 (N_1182,In_2911,In_3815);
xor U1183 (N_1183,In_2279,In_4190);
nand U1184 (N_1184,In_4637,In_3379);
or U1185 (N_1185,In_915,In_3821);
xnor U1186 (N_1186,In_3042,In_1196);
and U1187 (N_1187,In_3302,In_3032);
and U1188 (N_1188,In_3355,In_2848);
nand U1189 (N_1189,In_3153,In_969);
nor U1190 (N_1190,In_3651,In_1890);
and U1191 (N_1191,In_4608,In_4033);
and U1192 (N_1192,In_4725,In_4345);
or U1193 (N_1193,In_3258,In_98);
or U1194 (N_1194,In_2895,In_4727);
nand U1195 (N_1195,In_600,In_336);
xnor U1196 (N_1196,In_2010,In_4121);
nand U1197 (N_1197,In_4468,In_1419);
nor U1198 (N_1198,In_3705,In_4892);
and U1199 (N_1199,In_2031,In_1970);
nand U1200 (N_1200,In_491,In_3082);
and U1201 (N_1201,In_4527,In_2412);
xor U1202 (N_1202,In_1282,In_2891);
nand U1203 (N_1203,In_70,In_1944);
nand U1204 (N_1204,In_2906,In_715);
nand U1205 (N_1205,In_2770,In_523);
nor U1206 (N_1206,In_4234,In_2843);
and U1207 (N_1207,In_2884,In_3635);
or U1208 (N_1208,In_2710,In_1078);
nor U1209 (N_1209,In_3933,In_4443);
xor U1210 (N_1210,In_1522,In_1515);
nand U1211 (N_1211,In_4886,In_3761);
nor U1212 (N_1212,In_4236,In_1618);
xnor U1213 (N_1213,In_7,In_2495);
and U1214 (N_1214,In_3002,In_2804);
nand U1215 (N_1215,In_197,In_492);
xor U1216 (N_1216,In_4835,In_1250);
nor U1217 (N_1217,In_1449,In_802);
or U1218 (N_1218,In_603,In_259);
nand U1219 (N_1219,In_2289,In_2293);
nor U1220 (N_1220,In_2793,In_2297);
nor U1221 (N_1221,In_2664,In_2978);
and U1222 (N_1222,In_277,In_283);
nand U1223 (N_1223,In_383,In_1082);
nor U1224 (N_1224,In_4219,In_3419);
xnor U1225 (N_1225,In_833,In_1696);
nor U1226 (N_1226,In_3509,In_475);
and U1227 (N_1227,In_4346,In_2663);
nor U1228 (N_1228,In_4595,In_790);
xor U1229 (N_1229,In_3187,In_4374);
or U1230 (N_1230,In_1288,In_627);
or U1231 (N_1231,In_1367,In_1204);
or U1232 (N_1232,In_4788,In_3790);
or U1233 (N_1233,In_2784,In_3765);
or U1234 (N_1234,In_3390,In_4372);
nor U1235 (N_1235,In_1700,In_2100);
and U1236 (N_1236,In_3060,In_80);
nand U1237 (N_1237,In_1122,In_4596);
or U1238 (N_1238,In_125,In_3550);
nor U1239 (N_1239,In_2748,In_286);
xor U1240 (N_1240,In_205,In_1378);
or U1241 (N_1241,In_39,In_2832);
nor U1242 (N_1242,In_4182,In_2498);
or U1243 (N_1243,In_1079,In_2892);
nor U1244 (N_1244,In_1246,In_1972);
nor U1245 (N_1245,In_3879,In_4102);
and U1246 (N_1246,In_3619,In_2482);
nor U1247 (N_1247,In_2282,In_755);
xor U1248 (N_1248,In_1046,In_131);
or U1249 (N_1249,In_587,In_1852);
nand U1250 (N_1250,In_2381,In_1278);
or U1251 (N_1251,In_3812,In_1640);
nand U1252 (N_1252,In_1910,In_934);
xor U1253 (N_1253,In_650,In_3988);
xor U1254 (N_1254,In_2012,In_1329);
or U1255 (N_1255,In_414,In_136);
or U1256 (N_1256,In_2902,In_3736);
or U1257 (N_1257,In_4177,In_2588);
nor U1258 (N_1258,In_4492,In_2888);
nand U1259 (N_1259,In_842,In_137);
xnor U1260 (N_1260,In_1418,In_1120);
and U1261 (N_1261,In_4279,In_109);
and U1262 (N_1262,In_4304,In_1773);
nor U1263 (N_1263,In_2007,In_1926);
nor U1264 (N_1264,In_1523,In_1092);
xor U1265 (N_1265,In_4323,In_2603);
nand U1266 (N_1266,In_4923,In_2114);
and U1267 (N_1267,In_2631,In_1009);
nand U1268 (N_1268,In_3400,In_3837);
or U1269 (N_1269,In_4819,In_895);
nor U1270 (N_1270,In_4385,In_4460);
xor U1271 (N_1271,In_3460,In_4613);
or U1272 (N_1272,In_545,In_4965);
or U1273 (N_1273,In_4043,In_4097);
xnor U1274 (N_1274,In_2660,In_962);
nor U1275 (N_1275,In_2741,In_3926);
nand U1276 (N_1276,In_1366,In_3958);
xor U1277 (N_1277,In_2442,In_1351);
nand U1278 (N_1278,In_4679,In_2189);
nor U1279 (N_1279,In_571,In_711);
nand U1280 (N_1280,In_2390,In_902);
nand U1281 (N_1281,In_3574,In_3078);
nor U1282 (N_1282,In_534,In_2299);
nor U1283 (N_1283,In_388,In_4074);
nand U1284 (N_1284,In_2198,In_1624);
nor U1285 (N_1285,In_2754,In_3146);
and U1286 (N_1286,In_2819,In_3019);
and U1287 (N_1287,In_4215,In_1540);
nand U1288 (N_1288,In_3119,In_665);
nand U1289 (N_1289,In_4932,In_2363);
nor U1290 (N_1290,In_953,In_85);
or U1291 (N_1291,In_3249,In_395);
xor U1292 (N_1292,In_4414,In_221);
or U1293 (N_1293,In_2139,In_2024);
nand U1294 (N_1294,In_1794,In_1044);
and U1295 (N_1295,In_2346,In_2922);
or U1296 (N_1296,In_2554,In_144);
and U1297 (N_1297,In_2385,In_1048);
and U1298 (N_1298,In_3514,In_4941);
nor U1299 (N_1299,In_1549,In_59);
xnor U1300 (N_1300,In_1305,In_4202);
nor U1301 (N_1301,In_3159,In_2968);
and U1302 (N_1302,In_4306,In_4496);
nor U1303 (N_1303,In_4425,In_3200);
nor U1304 (N_1304,In_3351,In_4363);
xnor U1305 (N_1305,In_1971,In_3064);
nand U1306 (N_1306,In_607,In_180);
xnor U1307 (N_1307,In_1591,In_2130);
nand U1308 (N_1308,In_1208,In_1947);
nand U1309 (N_1309,In_1891,In_894);
xor U1310 (N_1310,In_2876,In_3365);
xor U1311 (N_1311,In_4597,In_2494);
or U1312 (N_1312,In_348,In_1995);
and U1313 (N_1313,In_3860,In_1739);
xor U1314 (N_1314,In_2077,In_2718);
or U1315 (N_1315,In_2739,In_4811);
nand U1316 (N_1316,In_4092,In_535);
or U1317 (N_1317,In_1965,In_412);
nand U1318 (N_1318,In_3631,In_4403);
nand U1319 (N_1319,In_1226,In_20);
and U1320 (N_1320,In_3748,In_2259);
xor U1321 (N_1321,In_4548,In_3729);
and U1322 (N_1322,In_2760,In_836);
nor U1323 (N_1323,In_1343,In_2113);
and U1324 (N_1324,In_4943,In_0);
nand U1325 (N_1325,In_1941,In_3722);
xor U1326 (N_1326,In_274,In_4034);
and U1327 (N_1327,In_362,In_4006);
or U1328 (N_1328,In_2510,In_656);
xor U1329 (N_1329,In_3865,In_734);
xor U1330 (N_1330,In_1602,In_3924);
and U1331 (N_1331,In_809,In_514);
or U1332 (N_1332,In_1080,In_2321);
xor U1333 (N_1333,In_2306,In_1933);
and U1334 (N_1334,In_3566,In_2396);
xnor U1335 (N_1335,In_3557,In_2044);
and U1336 (N_1336,In_4544,In_4641);
nand U1337 (N_1337,In_3348,In_3622);
and U1338 (N_1338,In_2424,In_444);
nor U1339 (N_1339,In_1663,In_3694);
nand U1340 (N_1340,In_729,In_91);
xor U1341 (N_1341,In_2620,In_4469);
nor U1342 (N_1342,In_73,In_287);
or U1343 (N_1343,In_3401,In_4759);
nor U1344 (N_1344,In_1300,In_3775);
nand U1345 (N_1345,In_2402,In_275);
and U1346 (N_1346,In_21,In_4295);
or U1347 (N_1347,In_2338,In_4816);
and U1348 (N_1348,In_4085,In_2069);
xnor U1349 (N_1349,In_4871,In_4317);
nand U1350 (N_1350,In_4450,In_3237);
xnor U1351 (N_1351,In_3586,In_1406);
and U1352 (N_1352,In_3977,In_1472);
nor U1353 (N_1353,In_206,In_2632);
xor U1354 (N_1354,In_1370,In_1976);
and U1355 (N_1355,In_834,In_1577);
xnor U1356 (N_1356,In_3931,In_3604);
xor U1357 (N_1357,In_2873,In_4333);
or U1358 (N_1358,In_916,In_4009);
or U1359 (N_1359,In_3954,In_315);
xnor U1360 (N_1360,In_248,In_1593);
or U1361 (N_1361,In_4174,In_1186);
or U1362 (N_1362,In_546,In_1267);
or U1363 (N_1363,In_2126,In_1494);
xor U1364 (N_1364,In_4319,In_2217);
and U1365 (N_1365,In_4163,In_2215);
or U1366 (N_1366,In_4984,In_2122);
and U1367 (N_1367,In_2165,In_1194);
and U1368 (N_1368,In_4348,In_1416);
nand U1369 (N_1369,In_2360,In_1943);
xor U1370 (N_1370,In_865,In_2078);
and U1371 (N_1371,In_2422,In_3441);
and U1372 (N_1372,In_2374,In_4604);
nor U1373 (N_1373,In_3357,In_1219);
nor U1374 (N_1374,In_4807,In_2824);
nor U1375 (N_1375,In_3370,In_4563);
xor U1376 (N_1376,In_3079,In_3287);
xor U1377 (N_1377,In_636,In_2944);
nand U1378 (N_1378,In_4528,In_4166);
or U1379 (N_1379,In_1100,In_3160);
xor U1380 (N_1380,In_2331,In_572);
xnor U1381 (N_1381,In_152,In_2283);
and U1382 (N_1382,In_3492,In_2742);
nor U1383 (N_1383,In_225,In_3908);
and U1384 (N_1384,In_2200,In_1851);
xor U1385 (N_1385,In_430,In_1043);
and U1386 (N_1386,In_2753,In_2546);
nor U1387 (N_1387,In_1784,In_2594);
nor U1388 (N_1388,In_3453,In_3998);
and U1389 (N_1389,In_4493,In_52);
and U1390 (N_1390,In_2827,In_4231);
xnor U1391 (N_1391,In_914,In_4866);
and U1392 (N_1392,In_2740,In_749);
and U1393 (N_1393,In_1478,In_4015);
xor U1394 (N_1394,In_4011,In_903);
nand U1395 (N_1395,In_3951,In_1613);
nor U1396 (N_1396,In_162,In_4686);
or U1397 (N_1397,In_2849,In_753);
and U1398 (N_1398,In_2235,In_4794);
and U1399 (N_1399,In_2862,In_622);
nor U1400 (N_1400,In_94,In_614);
or U1401 (N_1401,In_2842,In_3243);
or U1402 (N_1402,In_1166,In_3155);
nand U1403 (N_1403,In_1240,In_1673);
nand U1404 (N_1404,In_331,In_2646);
xnor U1405 (N_1405,In_2341,In_2835);
xnor U1406 (N_1406,In_1141,In_1674);
and U1407 (N_1407,In_4977,In_4302);
nand U1408 (N_1408,In_4767,In_1743);
nor U1409 (N_1409,In_1776,In_3377);
xor U1410 (N_1410,In_3436,In_1775);
and U1411 (N_1411,In_307,In_478);
xor U1412 (N_1412,In_1964,In_1692);
and U1413 (N_1413,In_4334,In_229);
and U1414 (N_1414,In_1492,In_3964);
xor U1415 (N_1415,In_1108,In_4873);
or U1416 (N_1416,In_4212,In_3599);
xor U1417 (N_1417,In_4060,In_2989);
or U1418 (N_1418,In_3115,In_3534);
nand U1419 (N_1419,In_954,In_398);
and U1420 (N_1420,In_4760,In_489);
and U1421 (N_1421,In_3169,In_961);
xor U1422 (N_1422,In_4186,In_496);
and U1423 (N_1423,In_717,In_4714);
or U1424 (N_1424,In_2358,In_2787);
and U1425 (N_1425,In_4082,In_2608);
nor U1426 (N_1426,In_542,In_3043);
xor U1427 (N_1427,In_3507,In_1585);
xor U1428 (N_1428,In_4642,In_1672);
and U1429 (N_1429,In_926,In_4655);
nand U1430 (N_1430,In_3208,In_403);
nor U1431 (N_1431,In_1863,In_1703);
or U1432 (N_1432,In_945,In_2182);
and U1433 (N_1433,In_1978,In_999);
and U1434 (N_1434,In_3841,In_246);
and U1435 (N_1435,In_350,In_2913);
nand U1436 (N_1436,In_344,In_1177);
nand U1437 (N_1437,In_2728,In_2532);
nand U1438 (N_1438,In_3091,In_1570);
nand U1439 (N_1439,In_4264,In_3238);
or U1440 (N_1440,In_4356,In_4169);
nand U1441 (N_1441,In_4571,In_2539);
or U1442 (N_1442,In_1587,In_4605);
xor U1443 (N_1443,In_577,In_4898);
and U1444 (N_1444,In_3422,In_1464);
and U1445 (N_1445,In_4066,In_1916);
nor U1446 (N_1446,In_4081,In_3152);
or U1447 (N_1447,In_472,In_3827);
nand U1448 (N_1448,In_3824,In_1387);
nand U1449 (N_1449,In_4699,In_2487);
or U1450 (N_1450,In_1675,In_2712);
or U1451 (N_1451,In_4262,In_4922);
or U1452 (N_1452,In_1368,In_3138);
and U1453 (N_1453,In_4018,In_14);
xnor U1454 (N_1454,In_2041,In_322);
or U1455 (N_1455,In_2796,In_2752);
nand U1456 (N_1456,In_593,In_1642);
and U1457 (N_1457,In_1990,In_901);
or U1458 (N_1458,In_2160,In_887);
xor U1459 (N_1459,In_3454,In_270);
nand U1460 (N_1460,In_1915,In_3576);
or U1461 (N_1461,In_2596,In_1156);
and U1462 (N_1462,In_1521,In_1309);
and U1463 (N_1463,In_2141,In_2857);
or U1464 (N_1464,In_2038,In_1949);
or U1465 (N_1465,In_57,In_2725);
or U1466 (N_1466,In_1511,In_3248);
nor U1467 (N_1467,In_3428,In_4110);
and U1468 (N_1468,In_4644,In_2224);
xor U1469 (N_1469,In_4280,In_4995);
nor U1470 (N_1470,In_2665,In_2327);
or U1471 (N_1471,In_2284,In_1854);
nor U1472 (N_1472,In_4126,In_3246);
xnor U1473 (N_1473,In_2611,In_3099);
or U1474 (N_1474,In_4203,In_1765);
nand U1475 (N_1475,In_2610,In_2109);
and U1476 (N_1476,In_4465,In_3667);
xnor U1477 (N_1477,In_3337,In_3455);
nor U1478 (N_1478,In_4328,In_3802);
or U1479 (N_1479,In_4645,In_442);
xor U1480 (N_1480,In_3757,In_340);
xnor U1481 (N_1481,In_3144,In_4120);
nor U1482 (N_1482,In_1477,In_3446);
nor U1483 (N_1483,In_187,In_1787);
or U1484 (N_1484,In_2864,In_2127);
xnor U1485 (N_1485,In_3203,In_1);
nand U1486 (N_1486,In_4354,In_1621);
or U1487 (N_1487,In_2447,In_1716);
and U1488 (N_1488,In_2854,In_1197);
and U1489 (N_1489,In_1006,In_3698);
nor U1490 (N_1490,In_4406,In_4213);
and U1491 (N_1491,In_2354,In_2853);
nor U1492 (N_1492,In_1927,In_3914);
nand U1493 (N_1493,In_3268,In_4687);
xor U1494 (N_1494,In_2999,In_3744);
xor U1495 (N_1495,In_1682,In_703);
xnor U1496 (N_1496,In_3307,In_4282);
nor U1497 (N_1497,In_539,In_4195);
nor U1498 (N_1498,In_3678,In_2291);
nor U1499 (N_1499,In_746,In_2);
xnor U1500 (N_1500,In_637,In_343);
and U1501 (N_1501,In_2107,In_980);
and U1502 (N_1502,In_1880,In_153);
or U1503 (N_1503,In_3075,In_3973);
nor U1504 (N_1504,In_175,In_1322);
nand U1505 (N_1505,In_4902,In_3424);
or U1506 (N_1506,In_538,In_4292);
nor U1507 (N_1507,In_4188,In_3806);
nor U1508 (N_1508,In_3679,In_859);
or U1509 (N_1509,In_669,In_4735);
and U1510 (N_1510,In_3170,In_291);
xor U1511 (N_1511,In_1168,In_3447);
or U1512 (N_1512,In_2364,In_4041);
nand U1513 (N_1513,In_4921,In_1041);
nor U1514 (N_1514,In_3375,In_1676);
xnor U1515 (N_1515,In_634,In_4621);
nor U1516 (N_1516,In_1666,In_3886);
or U1517 (N_1517,In_3051,In_1960);
nor U1518 (N_1518,In_4703,In_3858);
or U1519 (N_1519,In_2673,In_247);
or U1520 (N_1520,In_2767,In_3513);
xnor U1521 (N_1521,In_4973,In_1087);
xor U1522 (N_1522,In_828,In_1293);
or U1523 (N_1523,In_3779,In_4101);
nand U1524 (N_1524,In_4355,In_1793);
and U1525 (N_1525,In_222,In_3771);
xnor U1526 (N_1526,In_2347,In_47);
nor U1527 (N_1527,In_3189,In_1347);
nor U1528 (N_1528,In_2711,In_3191);
nand U1529 (N_1529,In_3906,In_186);
and U1530 (N_1530,In_4847,In_3957);
xnor U1531 (N_1531,In_3270,In_1931);
and U1532 (N_1532,In_3960,In_3551);
nor U1533 (N_1533,In_365,In_4930);
nor U1534 (N_1534,In_1410,In_525);
nor U1535 (N_1535,In_3223,In_861);
xor U1536 (N_1536,In_2434,In_770);
nand U1537 (N_1537,In_972,In_3666);
nand U1538 (N_1538,In_4667,In_639);
nand U1539 (N_1539,In_4359,In_1468);
nor U1540 (N_1540,In_1020,In_3289);
and U1541 (N_1541,In_3413,In_193);
nand U1542 (N_1542,In_3288,In_3630);
or U1543 (N_1543,In_189,In_3105);
nand U1544 (N_1544,In_2491,In_3164);
and U1545 (N_1545,In_4744,In_4970);
nand U1546 (N_1546,In_847,In_3301);
or U1547 (N_1547,In_4441,In_993);
xnor U1548 (N_1548,In_2241,In_3840);
and U1549 (N_1549,In_55,In_4039);
nor U1550 (N_1550,In_2765,In_4550);
or U1551 (N_1551,In_2335,In_3038);
nand U1552 (N_1552,In_1396,In_3762);
nor U1553 (N_1553,In_4432,In_2260);
and U1554 (N_1554,In_3871,In_701);
nand U1555 (N_1555,In_2375,In_4629);
or U1556 (N_1556,In_4170,In_314);
or U1557 (N_1557,In_3069,In_3452);
or U1558 (N_1558,In_3407,In_2183);
xor U1559 (N_1559,In_4037,In_2600);
nand U1560 (N_1560,In_110,In_1934);
or U1561 (N_1561,In_92,In_1414);
nor U1562 (N_1562,In_1810,In_2980);
nor U1563 (N_1563,In_2450,In_2952);
and U1564 (N_1564,In_1218,In_4925);
or U1565 (N_1565,In_303,In_4035);
or U1566 (N_1566,In_1010,In_706);
or U1567 (N_1567,In_2454,In_1001);
and U1568 (N_1568,In_2020,In_2726);
nand U1569 (N_1569,In_2446,In_4461);
nor U1570 (N_1570,In_4133,In_1534);
nor U1571 (N_1571,In_2476,In_3343);
xor U1572 (N_1572,In_1369,In_24);
nor U1573 (N_1573,In_2602,In_4648);
or U1574 (N_1574,In_3122,In_4146);
or U1575 (N_1575,In_2278,In_2397);
nor U1576 (N_1576,In_3297,In_309);
xnor U1577 (N_1577,In_4958,In_238);
xor U1578 (N_1578,In_4455,In_554);
or U1579 (N_1579,In_517,In_2708);
nand U1580 (N_1580,In_1686,In_2591);
or U1581 (N_1581,In_6,In_3893);
nor U1582 (N_1582,In_158,In_4046);
or U1583 (N_1583,In_1678,In_154);
or U1584 (N_1584,In_527,In_392);
nand U1585 (N_1585,In_2755,In_2055);
xnor U1586 (N_1586,In_618,In_906);
xnor U1587 (N_1587,In_1076,In_1341);
nand U1588 (N_1588,In_2897,In_946);
nor U1589 (N_1589,In_3904,In_3487);
or U1590 (N_1590,In_1582,In_1691);
nand U1591 (N_1591,In_2861,In_3967);
and U1592 (N_1592,In_986,In_3755);
xnor U1593 (N_1593,In_3875,In_2690);
nand U1594 (N_1594,In_951,In_3475);
nand U1595 (N_1595,In_1158,In_1529);
and U1596 (N_1596,In_1202,In_3567);
and U1597 (N_1597,In_2449,In_1221);
and U1598 (N_1598,In_1320,In_4505);
nor U1599 (N_1599,In_4859,In_4918);
or U1600 (N_1600,In_3265,In_4013);
and U1601 (N_1601,In_271,In_4004);
xnor U1602 (N_1602,In_2679,In_105);
or U1603 (N_1603,In_1545,In_2644);
and U1604 (N_1604,In_4502,In_3286);
xor U1605 (N_1605,In_2407,In_3128);
nand U1606 (N_1606,In_114,In_4240);
or U1607 (N_1607,In_4581,In_723);
or U1608 (N_1608,In_2940,In_4891);
nand U1609 (N_1609,In_3346,In_2190);
or U1610 (N_1610,In_4197,In_1104);
and U1611 (N_1611,In_805,In_299);
nor U1612 (N_1612,In_1357,In_4539);
or U1613 (N_1613,In_2366,In_1819);
xnor U1614 (N_1614,In_3199,In_4032);
nand U1615 (N_1615,In_1873,In_470);
nor U1616 (N_1616,In_873,In_602);
xnor U1617 (N_1617,In_1284,In_3282);
or U1618 (N_1618,In_2583,In_2671);
or U1619 (N_1619,In_2659,In_4513);
or U1620 (N_1620,In_541,In_716);
nor U1621 (N_1621,In_245,In_613);
nor U1622 (N_1622,In_3405,In_1936);
nand U1623 (N_1623,In_1336,In_4904);
xor U1624 (N_1624,In_1489,In_3652);
or U1625 (N_1625,In_464,In_2270);
and U1626 (N_1626,In_3339,In_2781);
nor U1627 (N_1627,In_2597,In_4291);
or U1628 (N_1628,In_1011,In_4893);
nand U1629 (N_1629,In_2551,In_4044);
or U1630 (N_1630,In_591,In_2352);
or U1631 (N_1631,In_1469,In_317);
xnor U1632 (N_1632,In_3371,In_4829);
nand U1633 (N_1633,In_1605,In_126);
nand U1634 (N_1634,In_4980,In_616);
nand U1635 (N_1635,In_1762,In_2218);
and U1636 (N_1636,In_2022,In_933);
or U1637 (N_1637,In_257,In_1505);
and U1638 (N_1638,In_1879,In_3376);
nor U1639 (N_1639,In_3483,In_3919);
or U1640 (N_1640,In_1607,In_1560);
and U1641 (N_1641,In_2674,In_2230);
nor U1642 (N_1642,In_4058,In_4017);
and U1643 (N_1643,In_1127,In_4038);
nor U1644 (N_1644,In_2161,In_2508);
and U1645 (N_1645,In_2696,In_609);
nor U1646 (N_1646,In_4459,In_2256);
nand U1647 (N_1647,In_1291,In_2775);
nand U1648 (N_1648,In_194,In_3071);
nand U1649 (N_1649,In_2332,In_3458);
nor U1650 (N_1650,In_583,In_4554);
nand U1651 (N_1651,In_2315,In_1495);
nand U1652 (N_1652,In_4851,In_484);
and U1653 (N_1653,In_2411,In_1161);
xnor U1654 (N_1654,In_3573,In_1412);
and U1655 (N_1655,In_4800,In_2266);
and U1656 (N_1656,In_3801,In_3878);
xor U1657 (N_1657,In_1667,In_339);
and U1658 (N_1658,In_1611,In_48);
or U1659 (N_1659,In_4267,In_2769);
xor U1660 (N_1660,In_2709,In_4774);
and U1661 (N_1661,In_2064,In_1777);
nor U1662 (N_1662,In_3322,In_4602);
xor U1663 (N_1663,In_230,In_1718);
xor U1664 (N_1664,In_745,In_1600);
and U1665 (N_1665,In_4272,In_3853);
or U1666 (N_1666,In_1868,In_4351);
or U1667 (N_1667,In_4071,In_3465);
or U1668 (N_1668,In_1281,In_3109);
nor U1669 (N_1669,In_3034,In_1358);
xor U1670 (N_1670,In_292,In_4773);
xnor U1671 (N_1671,In_1831,In_831);
xor U1672 (N_1672,In_4665,In_1799);
or U1673 (N_1673,In_762,In_3084);
xnor U1674 (N_1674,In_326,In_1752);
and U1675 (N_1675,In_101,In_2973);
and U1676 (N_1676,In_4722,In_1839);
and U1677 (N_1677,In_1500,In_1619);
nor U1678 (N_1678,In_3058,In_1929);
and U1679 (N_1679,In_3892,In_1463);
xor U1680 (N_1680,In_2459,In_3266);
nand U1681 (N_1681,In_2111,In_2342);
nand U1682 (N_1682,In_2918,In_2807);
nor U1683 (N_1683,In_4242,In_1598);
nor U1684 (N_1684,In_888,In_2124);
nand U1685 (N_1685,In_2571,In_3491);
nand U1686 (N_1686,In_4297,In_494);
nand U1687 (N_1687,In_4016,In_2838);
and U1688 (N_1688,In_4646,In_2954);
nand U1689 (N_1689,In_1302,In_3983);
xnor U1690 (N_1690,In_3747,In_4678);
nand U1691 (N_1691,In_4671,In_2091);
and U1692 (N_1692,In_4075,In_3505);
xnor U1693 (N_1693,In_2194,In_4158);
nor U1694 (N_1694,In_2145,In_4781);
or U1695 (N_1695,In_4757,In_3417);
nand U1696 (N_1696,In_1516,In_3685);
nor U1697 (N_1697,In_2605,In_1822);
xor U1698 (N_1698,In_4827,In_584);
nor U1699 (N_1699,In_4064,In_1334);
xor U1700 (N_1700,In_2904,In_4222);
xnor U1701 (N_1701,In_2406,In_1637);
or U1702 (N_1702,In_2537,In_1632);
and U1703 (N_1703,In_2258,In_2203);
nor U1704 (N_1704,In_4752,In_4447);
xnor U1705 (N_1705,In_928,In_3177);
or U1706 (N_1706,In_178,In_1892);
nor U1707 (N_1707,In_2413,In_1744);
nor U1708 (N_1708,In_2939,In_927);
nand U1709 (N_1709,In_4145,In_1179);
xnor U1710 (N_1710,In_3496,In_2168);
nand U1711 (N_1711,In_4136,In_355);
nand U1712 (N_1712,In_1555,In_3251);
xor U1713 (N_1713,In_3656,In_3050);
nand U1714 (N_1714,In_3869,In_468);
and U1715 (N_1715,In_81,In_1039);
nand U1716 (N_1716,In_1298,In_3023);
xnor U1717 (N_1717,In_3421,In_1578);
and U1718 (N_1718,In_408,In_1895);
nand U1719 (N_1719,In_278,In_2592);
and U1720 (N_1720,In_4594,In_3950);
nand U1721 (N_1721,In_4652,In_241);
nor U1722 (N_1722,In_2249,In_684);
nand U1723 (N_1723,In_1069,In_4845);
nor U1724 (N_1724,In_2426,In_341);
nand U1725 (N_1725,In_4208,In_4693);
or U1726 (N_1726,In_507,In_2135);
or U1727 (N_1727,In_2993,In_4928);
and U1728 (N_1728,In_1719,In_1903);
nand U1729 (N_1729,In_1438,In_1042);
nand U1730 (N_1730,In_359,In_3382);
or U1731 (N_1731,In_4260,In_1257);
xor U1732 (N_1732,In_3724,In_4433);
xnor U1733 (N_1733,In_2378,In_2821);
nor U1734 (N_1734,In_1975,In_1790);
nand U1735 (N_1735,In_1546,In_2175);
or U1736 (N_1736,In_40,In_297);
nand U1737 (N_1737,In_3838,In_2392);
nand U1738 (N_1738,In_4782,In_4108);
nor U1739 (N_1739,In_352,In_4881);
or U1740 (N_1740,In_4978,In_4160);
and U1741 (N_1741,In_3749,In_2813);
xor U1742 (N_1742,In_647,In_3309);
nor U1743 (N_1743,In_2101,In_896);
and U1744 (N_1744,In_4543,In_840);
and U1745 (N_1745,In_2097,In_1888);
and U1746 (N_1746,In_1774,In_2601);
nor U1747 (N_1747,In_1413,In_2613);
nor U1748 (N_1748,In_958,In_4706);
nor U1749 (N_1749,In_3669,In_4379);
and U1750 (N_1750,In_4992,In_227);
xnor U1751 (N_1751,In_4600,In_1807);
xnor U1752 (N_1752,In_2780,In_31);
nor U1753 (N_1753,In_3360,In_825);
xnor U1754 (N_1754,In_4558,In_4567);
nand U1755 (N_1755,In_4951,In_1386);
nor U1756 (N_1756,In_461,In_2581);
or U1757 (N_1757,In_3975,In_997);
or U1758 (N_1758,In_1032,In_3295);
or U1759 (N_1759,In_4285,In_1094);
xor U1760 (N_1760,In_3897,In_4422);
and U1761 (N_1761,In_3658,In_2180);
or U1762 (N_1762,In_4078,In_1853);
or U1763 (N_1763,In_3791,In_476);
and U1764 (N_1764,In_2344,In_151);
xnor U1765 (N_1765,In_188,In_3867);
nor U1766 (N_1766,In_3092,In_2879);
or U1767 (N_1767,In_948,In_3890);
or U1768 (N_1768,In_4689,In_4481);
or U1769 (N_1769,In_2142,In_963);
or U1770 (N_1770,In_3564,In_754);
nor U1771 (N_1771,In_4979,In_3133);
nor U1772 (N_1772,In_1060,In_2255);
and U1773 (N_1773,In_2865,In_4746);
nor U1774 (N_1774,In_2713,In_1074);
nand U1775 (N_1775,In_1627,In_1205);
or U1776 (N_1776,In_33,In_4119);
nand U1777 (N_1777,In_899,In_2443);
or U1778 (N_1778,In_4651,In_3372);
xor U1779 (N_1779,In_728,In_2666);
xor U1780 (N_1780,In_644,In_4002);
nand U1781 (N_1781,In_4663,In_4549);
and U1782 (N_1782,In_2274,In_1870);
or U1783 (N_1783,In_2948,In_2521);
nand U1784 (N_1784,In_2667,In_1634);
nand U1785 (N_1785,In_786,In_784);
and U1786 (N_1786,In_1058,In_163);
and U1787 (N_1787,In_4340,In_995);
xnor U1788 (N_1788,In_1760,In_2187);
nand U1789 (N_1789,In_2131,In_2931);
nand U1790 (N_1790,In_280,In_4401);
nand U1791 (N_1791,In_881,In_1645);
and U1792 (N_1792,In_413,In_1081);
and U1793 (N_1793,In_2395,In_521);
or U1794 (N_1794,In_4156,In_346);
xor U1795 (N_1795,In_1350,In_3686);
and U1796 (N_1796,In_2132,In_2867);
xor U1797 (N_1797,In_2138,In_1690);
xnor U1798 (N_1798,In_2733,In_857);
nor U1799 (N_1799,In_2616,In_547);
or U1800 (N_1800,In_4615,In_1415);
nor U1801 (N_1801,In_1899,In_2701);
nor U1802 (N_1802,In_1447,In_4238);
xor U1803 (N_1803,In_1049,In_1239);
or U1804 (N_1804,In_1750,In_4662);
nor U1805 (N_1805,In_2923,In_3723);
nand U1806 (N_1806,In_3707,In_1749);
nor U1807 (N_1807,In_450,In_2336);
and U1808 (N_1808,In_3319,In_3615);
xor U1809 (N_1809,In_1635,In_320);
or U1810 (N_1810,In_177,In_1000);
or U1811 (N_1811,In_135,In_2729);
or U1812 (N_1812,In_4606,In_4914);
or U1813 (N_1813,In_3537,In_3664);
and U1814 (N_1814,In_3326,In_1248);
and U1815 (N_1815,In_3710,In_3233);
and U1816 (N_1816,In_2087,In_3362);
or U1817 (N_1817,In_502,In_2026);
and U1818 (N_1818,In_4287,In_213);
xor U1819 (N_1819,In_994,In_566);
nand U1820 (N_1820,In_38,In_871);
nor U1821 (N_1821,In_4947,In_4696);
and U1822 (N_1822,In_1677,In_4257);
and U1823 (N_1823,In_1465,In_4211);
xor U1824 (N_1824,In_1958,In_863);
xnor U1825 (N_1825,In_1710,In_233);
nor U1826 (N_1826,In_4335,In_1883);
xor U1827 (N_1827,In_2153,In_117);
nand U1828 (N_1828,In_3411,In_2047);
and U1829 (N_1829,In_4541,In_428);
and U1830 (N_1830,In_2173,In_1193);
nor U1831 (N_1831,In_2751,In_2822);
and U1832 (N_1832,In_4526,In_3041);
and U1833 (N_1833,In_773,In_3126);
or U1834 (N_1834,In_66,In_3193);
or U1835 (N_1835,In_4863,In_3003);
xnor U1836 (N_1836,In_1994,In_4654);
or U1837 (N_1837,In_266,In_2697);
nand U1838 (N_1838,In_2889,In_3442);
nor U1839 (N_1839,In_2698,In_2303);
and U1840 (N_1840,In_1289,In_2531);
nor U1841 (N_1841,In_236,In_2851);
nand U1842 (N_1842,In_3693,In_4853);
or U1843 (N_1843,In_123,In_774);
or U1844 (N_1844,In_3655,In_143);
nor U1845 (N_1845,In_4628,In_1097);
or U1846 (N_1846,In_191,In_304);
nand U1847 (N_1847,In_318,In_2060);
nor U1848 (N_1848,In_1382,In_2391);
nor U1849 (N_1849,In_2466,In_3545);
nor U1850 (N_1850,In_1258,In_4069);
nor U1851 (N_1851,In_1065,In_1638);
and U1852 (N_1852,In_42,In_3031);
nor U1853 (N_1853,In_1821,In_869);
and U1854 (N_1854,In_3888,In_2874);
or U1855 (N_1855,In_3137,In_3787);
or U1856 (N_1856,In_4530,In_3462);
nor U1857 (N_1857,In_2001,In_1431);
and U1858 (N_1858,In_3364,In_1047);
nor U1859 (N_1859,In_272,In_4982);
and U1860 (N_1860,In_483,In_2027);
or U1861 (N_1861,In_3935,In_2828);
or U1862 (N_1862,In_4710,In_4427);
nand U1863 (N_1863,In_1025,In_382);
and U1864 (N_1864,In_1574,In_533);
xor U1865 (N_1865,In_3100,In_3113);
nor U1866 (N_1866,In_1680,In_2809);
nand U1867 (N_1867,In_4365,In_308);
nand U1868 (N_1868,In_3943,In_4519);
and U1869 (N_1869,In_3479,In_1781);
and U1870 (N_1870,In_752,In_385);
or U1871 (N_1871,In_4005,In_3949);
xor U1872 (N_1872,In_551,In_4435);
xor U1873 (N_1873,In_3987,In_1467);
or U1874 (N_1874,In_4523,In_3730);
nand U1875 (N_1875,In_4616,In_1294);
nand U1876 (N_1876,In_769,In_3510);
nand U1877 (N_1877,In_747,In_451);
nor U1878 (N_1878,In_4647,In_107);
xor U1879 (N_1879,In_2956,In_3846);
nand U1880 (N_1880,In_2471,In_4775);
and U1881 (N_1881,In_3313,In_2248);
or U1882 (N_1882,In_3560,In_2975);
xnor U1883 (N_1883,In_4476,In_4305);
nand U1884 (N_1884,In_4578,In_1024);
and U1885 (N_1885,In_1945,In_3175);
and U1886 (N_1886,In_3070,In_3296);
nor U1887 (N_1887,In_3725,In_2059);
and U1888 (N_1888,In_104,In_1045);
and U1889 (N_1889,In_3161,In_877);
nand U1890 (N_1890,In_4349,In_169);
nor U1891 (N_1891,In_2557,In_2890);
nand U1892 (N_1892,In_1738,In_3589);
xor U1893 (N_1893,In_1339,In_837);
nor U1894 (N_1894,In_384,In_885);
or U1895 (N_1895,In_878,In_4164);
xor U1896 (N_1896,In_1443,In_1271);
nand U1897 (N_1897,In_1428,In_1243);
nand U1898 (N_1898,In_2290,In_1496);
nor U1899 (N_1899,In_544,In_3647);
xor U1900 (N_1900,In_2926,In_4198);
or U1901 (N_1901,In_1720,In_818);
and U1902 (N_1902,In_2295,In_4318);
and U1903 (N_1903,In_635,In_3285);
nand U1904 (N_1904,In_4981,In_3145);
nand U1905 (N_1905,In_843,In_1661);
or U1906 (N_1906,In_2080,In_4672);
nand U1907 (N_1907,In_2844,In_2117);
nor U1908 (N_1908,In_3984,In_3305);
and U1909 (N_1909,In_3373,In_1730);
or U1910 (N_1910,In_949,In_1134);
xor U1911 (N_1911,In_1609,In_2745);
nand U1912 (N_1912,In_2910,In_2475);
nor U1913 (N_1913,In_2430,In_3516);
and U1914 (N_1914,In_552,In_4312);
nor U1915 (N_1915,In_930,In_1359);
nand U1916 (N_1916,In_4047,In_1544);
xnor U1917 (N_1917,In_3399,In_1664);
and U1918 (N_1918,In_719,In_3180);
nor U1919 (N_1919,In_2516,In_3033);
and U1920 (N_1920,In_1324,In_284);
and U1921 (N_1921,In_2783,In_3782);
or U1922 (N_1922,In_3448,In_1420);
nand U1923 (N_1923,In_447,In_1848);
or U1924 (N_1924,In_4635,In_2990);
nand U1925 (N_1925,In_3598,In_4140);
nor U1926 (N_1926,In_132,In_1460);
nor U1927 (N_1927,In_3005,In_1295);
and U1928 (N_1928,In_4778,In_4769);
xnor U1929 (N_1929,In_844,In_1147);
nand U1930 (N_1930,In_396,In_224);
or U1931 (N_1931,In_12,In_379);
or U1932 (N_1932,In_2261,In_4509);
or U1933 (N_1933,In_1130,In_4048);
and U1934 (N_1934,In_330,In_920);
or U1935 (N_1935,In_4381,In_1735);
nor U1936 (N_1936,In_4895,In_3283);
and U1937 (N_1937,In_2313,In_4935);
and U1938 (N_1938,In_4777,In_2840);
xor U1939 (N_1939,In_2348,In_2002);
or U1940 (N_1940,In_4821,In_1766);
xor U1941 (N_1941,In_694,In_1542);
nand U1942 (N_1942,In_4603,In_3321);
nor U1943 (N_1943,In_2373,In_3097);
and U1944 (N_1944,In_4562,In_2547);
nand U1945 (N_1945,In_3142,In_3086);
xnor U1946 (N_1946,In_1173,In_4690);
and U1947 (N_1947,In_612,In_3751);
nand U1948 (N_1948,In_1493,In_1315);
or U1949 (N_1949,In_1327,In_4695);
nor U1950 (N_1950,In_2774,In_3273);
nor U1951 (N_1951,In_2103,In_578);
nand U1952 (N_1952,In_1453,In_2081);
or U1953 (N_1953,In_1829,In_4309);
nand U1954 (N_1954,In_3024,In_4416);
nor U1955 (N_1955,In_1914,In_319);
or U1956 (N_1956,In_991,In_2896);
and U1957 (N_1957,In_1532,In_2448);
or U1958 (N_1958,In_4730,In_2789);
nor U1959 (N_1959,In_977,In_2159);
xor U1960 (N_1960,In_4350,In_3531);
nor U1961 (N_1961,In_2389,In_1816);
xor U1962 (N_1962,In_1803,In_4473);
nor U1963 (N_1963,In_528,In_2556);
or U1964 (N_1964,In_4311,In_1974);
xnor U1965 (N_1965,In_3561,In_3065);
and U1966 (N_1966,In_2936,In_2764);
xnor U1967 (N_1967,In_4392,In_1085);
or U1968 (N_1968,In_4137,In_3894);
xor U1969 (N_1969,In_2758,In_3819);
xor U1970 (N_1970,In_4996,In_1027);
and U1971 (N_1971,In_1470,In_1333);
nand U1972 (N_1972,In_2467,In_1259);
nand U1973 (N_1973,In_1222,In_3616);
nand U1974 (N_1974,In_4976,In_2281);
nor U1975 (N_1975,In_3158,In_3210);
xnor U1976 (N_1976,In_4525,In_4153);
and U1977 (N_1977,In_4623,In_3124);
and U1978 (N_1978,In_2318,In_3940);
and U1979 (N_1979,In_290,In_3989);
nand U1980 (N_1980,In_4021,In_4485);
nand U1981 (N_1981,In_592,In_3939);
and U1982 (N_1982,In_4223,In_702);
or U1983 (N_1983,In_3620,In_2063);
or U1984 (N_1984,In_2732,In_2831);
nand U1985 (N_1985,In_4638,In_555);
or U1986 (N_1986,In_201,In_4631);
nor U1987 (N_1987,In_3278,In_1629);
and U1988 (N_1988,In_1040,In_4168);
or U1989 (N_1989,In_1262,In_390);
nand U1990 (N_1990,In_60,In_4998);
nand U1991 (N_1991,In_727,In_2812);
nand U1992 (N_1992,In_3684,In_4141);
and U1993 (N_1993,In_4442,In_3634);
nor U1994 (N_1994,In_944,In_4598);
nor U1995 (N_1995,In_4955,In_1005);
and U1996 (N_1996,In_2514,In_4838);
or U1997 (N_1997,In_3194,In_2102);
and U1998 (N_1998,In_1679,In_3506);
or U1999 (N_1999,In_989,In_659);
nor U2000 (N_2000,In_2846,In_3464);
and U2001 (N_2001,In_4284,In_2172);
xor U2002 (N_2002,In_4253,In_661);
nor U2003 (N_2003,In_4358,In_548);
xor U2004 (N_2004,In_4721,In_1171);
nor U2005 (N_2005,In_4150,In_4834);
nand U2006 (N_2006,In_2369,In_1061);
nand U2007 (N_2007,In_1869,In_4522);
xnor U2008 (N_2008,In_4843,In_3332);
xor U2009 (N_2009,In_1804,In_2638);
xor U2010 (N_2010,In_981,In_2960);
nand U2011 (N_2011,In_3675,In_1338);
or U2012 (N_2012,In_3733,In_4796);
and U2013 (N_2013,In_437,In_4634);
or U2014 (N_2014,In_3660,In_3111);
or U2015 (N_2015,In_1143,In_3162);
nor U2016 (N_2016,In_4619,In_4583);
nand U2017 (N_2017,In_2582,In_3474);
nor U2018 (N_2018,In_781,In_3785);
nand U2019 (N_2019,In_406,In_2465);
and U2020 (N_2020,In_3706,In_1180);
nor U2021 (N_2021,In_4682,In_4394);
xnor U2022 (N_2022,In_654,In_1405);
nand U2023 (N_2023,In_3872,In_3205);
and U2024 (N_2024,In_1403,In_1887);
xor U2025 (N_2025,In_4937,In_2615);
nand U2026 (N_2026,In_3188,In_37);
and U2027 (N_2027,In_3847,In_4204);
nand U2028 (N_2028,In_4704,In_4449);
nand U2029 (N_2029,In_2207,In_4336);
and U2030 (N_2030,In_2652,In_1937);
nand U2031 (N_2031,In_3992,In_1311);
and U2032 (N_2032,In_4045,In_3746);
and U2033 (N_2033,In_223,In_595);
nand U2034 (N_2034,In_53,In_3945);
or U2035 (N_2035,In_1287,In_3845);
nand U2036 (N_2036,In_115,In_3568);
nand U2037 (N_2037,In_1514,In_2201);
nor U2038 (N_2038,In_3603,In_3280);
and U2039 (N_2039,In_3148,In_166);
xor U2040 (N_2040,In_1462,In_4428);
or U2041 (N_2041,In_4664,In_2197);
xor U2042 (N_2042,In_2277,In_660);
or U2043 (N_2043,In_4542,In_471);
nor U2044 (N_2044,In_2045,In_2505);
xnor U2045 (N_2045,In_2915,In_1571);
nand U2046 (N_2046,In_673,In_2607);
and U2047 (N_2047,In_3279,In_3836);
or U2048 (N_2048,In_1722,In_174);
xnor U2049 (N_2049,In_2743,In_2869);
nor U2050 (N_2050,In_2116,In_3167);
nor U2051 (N_2051,In_4424,In_4131);
and U2052 (N_2052,In_4864,In_4817);
nor U2053 (N_2053,In_2222,In_3699);
and U2054 (N_2054,In_3171,In_3340);
or U2055 (N_2055,In_4367,In_490);
or U2056 (N_2056,In_2545,In_2908);
xnor U2057 (N_2057,In_3866,In_1228);
or U2058 (N_2058,In_4147,In_1859);
nor U2059 (N_2059,In_1917,In_4244);
and U2060 (N_2060,In_4588,In_302);
nor U2061 (N_2061,In_4412,In_4023);
nand U2062 (N_2062,In_1480,In_4956);
nand U2063 (N_2063,In_4107,In_858);
xnor U2064 (N_2064,In_2536,In_1656);
or U2065 (N_2065,In_2612,In_2834);
nor U2066 (N_2066,In_3835,In_1737);
or U2067 (N_2067,In_2550,In_3389);
or U2068 (N_2068,In_1121,In_1037);
xnor U2069 (N_2069,In_3477,In_3953);
and U2070 (N_2070,In_693,In_1476);
and U2071 (N_2071,In_4084,In_4310);
or U2072 (N_2072,In_3363,In_1433);
and U2073 (N_2073,In_1714,In_3687);
nand U2074 (N_2074,In_4906,In_4971);
or U2075 (N_2075,In_3583,In_811);
and U2076 (N_2076,In_3226,In_377);
nand U2077 (N_2077,In_1375,In_2538);
nor U2078 (N_2078,In_3663,In_506);
xor U2079 (N_2079,In_2852,In_707);
nand U2080 (N_2080,In_4650,In_118);
nor U2081 (N_2081,In_3607,In_4691);
xnor U2082 (N_2082,In_2584,In_1884);
or U2083 (N_2083,In_2970,In_3181);
nor U2084 (N_2084,In_907,In_1993);
or U2085 (N_2085,In_2089,In_1837);
and U2086 (N_2086,In_1596,In_446);
nor U2087 (N_2087,In_1652,In_11);
and U2088 (N_2088,In_2267,In_3792);
or U2089 (N_2089,In_45,In_4286);
or U2090 (N_2090,In_4740,In_4776);
and U2091 (N_2091,In_1260,In_1503);
nor U2092 (N_2092,In_3104,In_3839);
xor U2093 (N_2093,In_780,In_3913);
nor U2094 (N_2094,In_3406,In_739);
nand U2095 (N_2095,In_1764,In_1456);
or U2096 (N_2096,In_1788,In_3172);
nor U2097 (N_2097,In_4254,In_4836);
and U2098 (N_2098,In_3727,In_368);
nand U2099 (N_2099,In_4867,In_208);
nand U2100 (N_2100,In_1543,In_1332);
nand U2101 (N_2101,In_3928,In_1346);
or U2102 (N_2102,In_3425,In_4754);
xor U2103 (N_2103,In_4936,In_922);
nor U2104 (N_2104,In_212,In_3393);
or U2105 (N_2105,In_399,In_3795);
nand U2106 (N_2106,In_580,In_3047);
and U2107 (N_2107,In_1099,In_2337);
and U2108 (N_2108,In_2629,In_2549);
nand U2109 (N_2109,In_463,In_841);
nand U2110 (N_2110,In_2380,In_649);
nor U2111 (N_2111,In_2329,In_3595);
xnor U2112 (N_2112,In_2527,In_2057);
xnor U2113 (N_2113,In_2483,In_3381);
or U2114 (N_2114,In_3306,In_3728);
nand U2115 (N_2115,In_2691,In_3608);
xor U2116 (N_2116,In_3275,In_4124);
xnor U2117 (N_2117,In_2687,In_3440);
or U2118 (N_2118,In_2649,In_759);
or U2119 (N_2119,In_1648,In_1442);
and U2120 (N_2120,In_311,In_258);
nand U2121 (N_2121,In_3754,In_3601);
xor U2122 (N_2122,In_923,In_1713);
and U2123 (N_2123,In_3068,In_925);
nand U2124 (N_2124,In_549,In_2014);
xnor U2125 (N_2125,In_4400,In_2506);
and U2126 (N_2126,In_2445,In_1550);
nand U2127 (N_2127,In_1847,In_3993);
xnor U2128 (N_2128,In_2585,In_4342);
nand U2129 (N_2129,In_974,In_4115);
nor U2130 (N_2130,In_767,In_1440);
nand U2131 (N_2131,In_1174,In_2292);
or U2132 (N_2132,In_4840,In_452);
nand U2133 (N_2133,In_3579,In_1439);
nor U2134 (N_2134,In_1564,In_2355);
nand U2135 (N_2135,In_1950,In_3255);
xor U2136 (N_2136,In_849,In_604);
xor U2137 (N_2137,In_2071,In_846);
xor U2138 (N_2138,In_4599,In_1639);
nor U2139 (N_2139,In_1641,In_3844);
xnor U2140 (N_2140,In_3597,In_4747);
or U2141 (N_2141,In_1153,In_405);
nand U2142 (N_2142,In_3397,In_420);
or U2143 (N_2143,In_4712,In_4303);
nor U2144 (N_2144,In_4738,In_1132);
or U2145 (N_2145,In_1999,In_3176);
nor U2146 (N_2146,In_4464,In_1401);
nand U2147 (N_2147,In_3445,In_4402);
nor U2148 (N_2148,In_4454,In_2461);
or U2149 (N_2149,In_2504,In_3735);
and U2150 (N_2150,In_3121,In_2119);
or U2151 (N_2151,In_2123,In_608);
xnor U2152 (N_2152,In_1698,In_3915);
and U2153 (N_2153,In_2509,In_4785);
or U2154 (N_2154,In_990,In_1383);
xnor U2155 (N_2155,In_1646,In_2129);
nand U2156 (N_2156,In_3665,In_4787);
or U2157 (N_2157,In_2037,In_2626);
and U2158 (N_2158,In_77,In_2859);
xnor U2159 (N_2159,In_2907,In_2314);
nor U2160 (N_2160,In_1556,In_1988);
and U2161 (N_2161,In_2662,In_4274);
or U2162 (N_2162,In_2634,In_585);
and U2163 (N_2163,In_801,In_4716);
xor U2164 (N_2164,In_2630,In_2489);
or U2165 (N_2165,In_3143,In_2976);
xor U2166 (N_2166,In_2400,In_4630);
nor U2167 (N_2167,In_1876,In_1093);
nor U2168 (N_2168,In_2186,In_3544);
nand U2169 (N_2169,In_3734,In_3895);
nor U2170 (N_2170,In_4025,In_2473);
nor U2171 (N_2171,In_509,In_1702);
nor U2172 (N_2172,In_4096,In_4399);
nor U2173 (N_2173,In_704,In_2429);
xor U2174 (N_2174,In_812,In_485);
xnor U2175 (N_2175,In_3118,In_1904);
xnor U2176 (N_2176,In_785,In_3456);
and U2177 (N_2177,In_1297,In_4159);
and U2178 (N_2178,In_1823,In_3526);
nand U2179 (N_2179,In_3059,In_3539);
or U2180 (N_2180,In_3843,In_1707);
nor U2181 (N_2181,In_1592,In_2205);
nor U2182 (N_2182,In_3476,In_4820);
or U2183 (N_2183,In_1172,In_3518);
and U2184 (N_2184,In_3683,In_4307);
nor U2185 (N_2185,In_50,In_2776);
or U2186 (N_2186,In_4138,In_449);
or U2187 (N_2187,In_4964,In_674);
nand U2188 (N_2188,In_3334,In_1913);
or U2189 (N_2189,In_3786,In_4896);
or U2190 (N_2190,In_3027,In_1314);
xnor U2191 (N_2191,In_1486,In_1144);
and U2192 (N_2192,In_3602,In_182);
xor U2193 (N_2193,In_2868,In_4818);
xnor U2194 (N_2194,In_2593,In_1397);
and U2195 (N_2195,In_2806,In_3851);
or U2196 (N_2196,In_3758,In_211);
nor U2197 (N_2197,In_557,In_2219);
xor U2198 (N_2198,In_4176,In_3131);
or U2199 (N_2199,In_146,In_434);
nor U2200 (N_2200,In_696,In_1313);
and U2201 (N_2201,In_3013,In_2870);
or U2202 (N_2202,In_1230,In_1013);
and U2203 (N_2203,In_3629,In_947);
xor U2204 (N_2204,In_4327,In_1362);
nand U2205 (N_2205,In_4826,In_4167);
or U2206 (N_2206,In_2170,In_3489);
nor U2207 (N_2207,In_3903,In_1729);
nand U2208 (N_2208,In_3165,In_2720);
nor U2209 (N_2209,In_367,In_876);
xnor U2210 (N_2210,In_1668,In_1881);
and U2211 (N_2211,In_3764,In_4369);
nand U2212 (N_2212,In_4143,In_581);
or U2213 (N_2213,In_565,In_64);
nand U2214 (N_2214,In_3192,In_3292);
or U2215 (N_2215,In_244,In_4487);
or U2216 (N_2216,In_2343,In_1657);
nand U2217 (N_2217,In_1355,In_3230);
nand U2218 (N_2218,In_642,In_3184);
xor U2219 (N_2219,In_3106,In_1557);
and U2220 (N_2220,In_3341,In_2108);
and U2221 (N_2221,In_4497,In_1266);
and U2222 (N_2222,In_2606,In_2134);
and U2223 (N_2223,In_596,In_3554);
nand U2224 (N_2224,In_4501,In_4154);
nor U2225 (N_2225,In_2563,In_1858);
xnor U2226 (N_2226,In_2942,In_4255);
and U2227 (N_2227,In_889,In_1920);
and U2228 (N_2228,In_2766,In_1234);
nand U2229 (N_2229,In_353,In_3829);
nor U2230 (N_2230,In_1902,In_4858);
and U2231 (N_2231,In_2548,In_4480);
nand U2232 (N_2232,In_732,In_3066);
nor U2233 (N_2233,In_2242,In_1759);
or U2234 (N_2234,In_2707,In_1530);
nand U2235 (N_2235,In_917,In_4080);
nand U2236 (N_2236,In_1724,In_4684);
xor U2237 (N_2237,In_281,In_3921);
xnor U2238 (N_2238,In_2093,In_4408);
or U2239 (N_2239,In_4822,In_3654);
nor U2240 (N_2240,In_4249,In_1662);
xor U2241 (N_2241,In_2515,In_4856);
xnor U2242 (N_2242,In_1454,In_28);
nand U2243 (N_2243,In_1160,In_1771);
and U2244 (N_2244,In_3552,In_4386);
nand U2245 (N_2245,In_2716,In_1484);
nor U2246 (N_2246,In_1182,In_2757);
nor U2247 (N_2247,In_2211,In_2164);
nand U2248 (N_2248,In_4607,In_3543);
xnor U2249 (N_2249,In_2618,In_4192);
or U2250 (N_2250,In_119,In_4975);
nor U2251 (N_2251,In_1922,In_2953);
xnor U2252 (N_2252,In_2416,In_1261);
nand U2253 (N_2253,In_620,In_2562);
or U2254 (N_2254,In_2470,In_2815);
nand U2255 (N_2255,In_3830,In_1263);
nand U2256 (N_2256,In_2121,In_3773);
nand U2257 (N_2257,In_1437,In_1084);
or U2258 (N_2258,In_2308,In_3416);
and U2259 (N_2259,In_4547,In_1506);
and U2260 (N_2260,In_4676,In_4743);
or U2261 (N_2261,In_3585,In_2177);
and U2262 (N_2262,In_4030,In_2967);
nor U2263 (N_2263,In_4622,In_722);
nand U2264 (N_2264,In_1982,In_1422);
nor U2265 (N_2265,In_4584,In_1778);
nand U2266 (N_2266,In_4256,In_4771);
or U2267 (N_2267,In_3623,In_1826);
xnor U2268 (N_2268,In_1815,In_168);
nand U2269 (N_2269,In_4582,In_252);
xnor U2270 (N_2270,In_220,In_1290);
nand U2271 (N_2271,In_2372,In_1527);
and U2272 (N_2272,In_720,In_4770);
and U2273 (N_2273,In_4151,In_1319);
or U2274 (N_2274,In_1014,In_621);
nand U2275 (N_2275,In_2643,In_477);
nor U2276 (N_2276,In_559,In_3976);
xnor U2277 (N_2277,In_813,In_2185);
nand U2278 (N_2278,In_2118,In_4985);
nor U2279 (N_2279,In_149,In_159);
xor U2280 (N_2280,In_3948,In_4666);
nand U2281 (N_2281,In_2856,In_3291);
and U2282 (N_2282,In_3970,In_1567);
and U2283 (N_2283,In_2695,In_1588);
xor U2284 (N_2284,In_3239,In_1878);
and U2285 (N_2285,In_941,In_312);
or U2286 (N_2286,In_2927,In_3703);
and U2287 (N_2287,In_3081,In_1277);
nor U2288 (N_2288,In_2120,In_4377);
or U2289 (N_2289,In_3077,In_3719);
nor U2290 (N_2290,In_2353,In_4805);
nor U2291 (N_2291,In_682,In_1251);
nand U2292 (N_2292,In_2464,In_2152);
nor U2293 (N_2293,In_4882,In_1056);
and U2294 (N_2294,In_1754,In_4118);
or U2295 (N_2295,In_2627,In_86);
xor U2296 (N_2296,In_3776,In_4993);
nand U2297 (N_2297,In_4265,In_160);
nor U2298 (N_2298,In_1906,In_3242);
nand U2299 (N_2299,In_4688,In_2761);
and U2300 (N_2300,In_3468,In_1590);
and U2301 (N_2301,In_2096,In_4313);
and U2302 (N_2302,In_3909,In_1843);
and U2303 (N_2303,In_3095,In_978);
or U2304 (N_2304,In_1123,In_3004);
and U2305 (N_2305,In_2811,In_2050);
or U2306 (N_2306,In_4900,In_1349);
nand U2307 (N_2307,In_2076,In_3037);
and U2308 (N_2308,In_2304,In_4636);
nand U2309 (N_2309,In_3012,In_712);
nor U2310 (N_2310,In_1620,In_1708);
nand U2311 (N_2311,In_4889,In_3098);
nand U2312 (N_2312,In_2229,In_3659);
or U2313 (N_2313,In_2210,In_879);
nand U2314 (N_2314,In_3426,In_1644);
and U2315 (N_2315,In_3323,In_453);
or U2316 (N_2316,In_260,In_239);
and U2317 (N_2317,In_4362,In_2171);
nand U2318 (N_2318,In_3022,In_1187);
nor U2319 (N_2319,In_1573,In_699);
or U2320 (N_2320,In_480,In_764);
nor U2321 (N_2321,In_63,In_4022);
nor U2322 (N_2322,In_778,In_487);
and U2323 (N_2323,In_4073,In_3234);
or U2324 (N_2324,In_4019,In_1830);
nor U2325 (N_2325,In_112,In_2882);
nor U2326 (N_2326,In_3691,In_401);
nor U2327 (N_2327,In_959,In_606);
and U2328 (N_2328,In_2715,In_243);
and U2329 (N_2329,In_4360,In_10);
nor U2330 (N_2330,In_210,In_3134);
xnor U2331 (N_2331,In_2945,In_2302);
and U2332 (N_2332,In_3946,In_1376);
xnor U2333 (N_2333,In_4173,In_4579);
xor U2334 (N_2334,In_2357,In_3593);
and U2335 (N_2335,In_964,In_3325);
xnor U2336 (N_2336,In_1118,In_1861);
nand U2337 (N_2337,In_724,In_394);
or U2338 (N_2338,In_3648,In_987);
nor U2339 (N_2339,In_2485,In_4020);
nand U2340 (N_2340,In_1997,In_4739);
and U2341 (N_2341,In_668,In_4750);
or U2342 (N_2342,In_4144,In_183);
nor U2343 (N_2343,In_1748,In_4931);
xor U2344 (N_2344,In_2204,In_3328);
or U2345 (N_2345,In_285,In_4570);
xnor U2346 (N_2346,In_2043,In_2439);
xnor U2347 (N_2347,In_1939,In_1809);
xnor U2348 (N_2348,In_1909,In_3190);
and U2349 (N_2349,In_2886,In_2917);
nand U2350 (N_2350,In_391,In_4456);
or U2351 (N_2351,In_4719,In_2943);
or U2352 (N_2352,In_4494,In_3062);
nor U2353 (N_2353,In_3712,In_4067);
nand U2354 (N_2354,In_56,In_4946);
or U2355 (N_2355,In_4104,In_3127);
xor U2356 (N_2356,In_2981,In_3202);
and U2357 (N_2357,In_1659,In_3259);
and U2358 (N_2358,In_4574,In_4472);
xor U2359 (N_2359,In_2727,In_133);
nor U2360 (N_2360,In_2253,In_1665);
and U2361 (N_2361,In_1220,In_2003);
nor U2362 (N_2362,In_1237,In_4499);
and U2363 (N_2363,In_1769,In_2150);
or U2364 (N_2364,In_23,In_4162);
xor U2365 (N_2365,In_4639,In_605);
or U2366 (N_2366,In_4184,In_1955);
nand U2367 (N_2367,In_3932,In_2137);
xor U2368 (N_2368,In_4939,In_3108);
xnor U2369 (N_2369,In_4325,In_4573);
or U2370 (N_2370,In_2453,In_3264);
nand U2371 (N_2371,In_4217,In_3653);
xor U2372 (N_2372,In_2460,In_4378);
nand U2373 (N_2373,In_610,In_3380);
or U2374 (N_2374,In_1518,In_301);
nand U2375 (N_2375,In_3861,In_3674);
nand U2376 (N_2376,In_3221,In_2340);
xor U2377 (N_2377,In_3759,In_4289);
and U2378 (N_2378,In_2499,In_1385);
nand U2379 (N_2379,In_1987,In_2333);
nor U2380 (N_2380,In_4832,In_2307);
or U2381 (N_2381,In_3942,In_1623);
nor U2382 (N_2382,In_3512,In_1838);
nor U2383 (N_2383,In_1050,In_2149);
and U2384 (N_2384,In_760,In_4673);
and U2385 (N_2385,In_4701,In_1304);
or U2386 (N_2386,In_2747,In_3433);
nor U2387 (N_2387,In_3769,In_4503);
nor U2388 (N_2388,In_4924,In_4707);
xnor U2389 (N_2389,In_323,In_599);
nor U2390 (N_2390,In_3881,In_4907);
and U2391 (N_2391,In_2144,In_4949);
nand U2392 (N_2392,In_1715,In_1089);
and U2393 (N_2393,In_2998,In_3488);
nor U2394 (N_2394,In_156,In_1520);
xor U2395 (N_2395,In_779,In_4281);
xnor U2396 (N_2396,In_2497,In_4225);
nor U2397 (N_2397,In_2988,In_929);
xnor U2398 (N_2398,In_4010,In_708);
xnor U2399 (N_2399,In_543,In_2351);
or U2400 (N_2400,In_3581,In_2285);
and U2401 (N_2401,In_2028,In_988);
xor U2402 (N_2402,In_743,In_321);
nor U2403 (N_2403,In_966,In_1786);
nor U2404 (N_2404,In_2503,In_2833);
xor U2405 (N_2405,In_71,In_46);
xor U2406 (N_2406,In_839,In_4532);
and U2407 (N_2407,In_3553,In_2599);
and U2408 (N_2408,In_2233,In_465);
xor U2409 (N_2409,In_265,In_89);
nor U2410 (N_2410,In_3996,In_4270);
xnor U2411 (N_2411,In_4419,In_1181);
and U2412 (N_2412,In_2799,In_2300);
nor U2413 (N_2413,In_3320,In_1070);
and U2414 (N_2414,In_1581,In_3272);
nor U2415 (N_2415,In_4569,In_4087);
nand U2416 (N_2416,In_2723,In_179);
nor U2417 (N_2417,In_298,In_3592);
nand U2418 (N_2418,In_4731,In_253);
xnor U2419 (N_2419,In_2345,In_3985);
nand U2420 (N_2420,In_4657,In_692);
and U2421 (N_2421,In_1998,In_4250);
xnor U2422 (N_2422,In_2756,In_3213);
and U2423 (N_2423,In_2544,In_4761);
nor U2424 (N_2424,In_4139,In_3891);
nor U2425 (N_2425,In_3822,In_4475);
and U2426 (N_2426,In_2526,In_601);
xor U2427 (N_2427,In_2994,In_4175);
xor U2428 (N_2428,In_2323,In_3538);
xnor U2429 (N_2429,In_816,In_2839);
nor U2430 (N_2430,In_1213,In_742);
and U2431 (N_2431,In_4963,In_2328);
nor U2432 (N_2432,In_4855,In_1986);
xnor U2433 (N_2433,In_2067,In_1323);
nor U2434 (N_2434,In_3006,In_598);
or U2435 (N_2435,In_1669,In_2737);
nand U2436 (N_2436,In_4221,In_3224);
nor U2437 (N_2437,In_3937,In_4626);
nand U2438 (N_2438,In_3959,In_3662);
or U2439 (N_2439,In_3470,In_1572);
or U2440 (N_2440,In_2919,In_4233);
and U2441 (N_2441,In_2492,In_4741);
xnor U2442 (N_2442,In_4028,In_1980);
and U2443 (N_2443,In_1845,In_4068);
or U2444 (N_2444,In_3547,In_4261);
or U2445 (N_2445,In_4624,In_1626);
xnor U2446 (N_2446,In_3182,In_4917);
nand U2447 (N_2447,In_2530,In_570);
xor U2448 (N_2448,In_503,In_3102);
nor U2449 (N_2449,In_116,In_4780);
xnor U2450 (N_2450,In_2286,In_4413);
nor U2451 (N_2451,In_1806,In_3352);
xor U2452 (N_2452,In_1235,In_709);
nand U2453 (N_2453,In_1951,In_3969);
nand U2454 (N_2454,In_766,In_1575);
or U2455 (N_2455,In_1742,In_1286);
xnor U2456 (N_2456,In_1167,In_1491);
xor U2457 (N_2457,In_4117,In_268);
nand U2458 (N_2458,In_76,In_3569);
nor U2459 (N_2459,In_518,In_3149);
xor U2460 (N_2460,In_1728,In_3385);
nor U2461 (N_2461,In_1979,In_3250);
xnor U2462 (N_2462,In_196,In_4338);
xnor U2463 (N_2463,In_1541,In_3532);
and U2464 (N_2464,In_2110,In_1395);
nand U2465 (N_2465,In_87,In_3198);
xnor U2466 (N_2466,In_1292,In_2104);
nand U2467 (N_2467,In_4850,In_741);
nor U2468 (N_2468,In_3826,In_2558);
and U2469 (N_2469,In_2574,In_1211);
nor U2470 (N_2470,In_3395,In_1364);
and U2471 (N_2471,In_3689,In_1751);
nand U2472 (N_2472,In_1310,In_1446);
and U2473 (N_2473,In_4189,In_867);
or U2474 (N_2474,In_2639,In_124);
nor U2475 (N_2475,In_3952,In_677);
or U2476 (N_2476,In_3017,In_393);
or U2477 (N_2477,In_4915,In_4883);
nor U2478 (N_2478,In_1608,In_630);
xnor U2479 (N_2479,In_3863,In_4079);
nand U2480 (N_2480,In_4869,In_3444);
nand U2481 (N_2481,In_4439,In_2651);
nand U2482 (N_2482,In_2462,In_1129);
xor U2483 (N_2483,In_3780,In_2035);
nor U2484 (N_2484,In_2914,In_410);
or U2485 (N_2485,In_1448,In_3944);
nand U2486 (N_2486,In_2049,In_2949);
or U2487 (N_2487,In_29,In_4534);
nand U2488 (N_2488,In_2535,In_1426);
or U2489 (N_2489,In_3398,In_2234);
xor U2490 (N_2490,In_3463,In_617);
xnor U2491 (N_2491,In_1371,In_3502);
xor U2492 (N_2492,In_2658,In_2410);
nand U2493 (N_2493,In_4100,In_500);
and U2494 (N_2494,In_3087,In_375);
and U2495 (N_2495,In_1411,In_2578);
and U2496 (N_2496,In_4974,In_4556);
nor U2497 (N_2497,In_646,In_1502);
and U2498 (N_2498,In_4545,In_4887);
and U2499 (N_2499,In_1077,In_1273);
nand U2500 (N_2500,In_254,In_4342);
or U2501 (N_2501,In_1151,In_3946);
nand U2502 (N_2502,In_1372,In_3084);
nor U2503 (N_2503,In_1940,In_981);
and U2504 (N_2504,In_518,In_990);
and U2505 (N_2505,In_4903,In_221);
and U2506 (N_2506,In_3128,In_18);
nand U2507 (N_2507,In_2728,In_4487);
or U2508 (N_2508,In_3428,In_4564);
and U2509 (N_2509,In_1370,In_163);
or U2510 (N_2510,In_3655,In_4917);
nand U2511 (N_2511,In_4326,In_728);
or U2512 (N_2512,In_3188,In_1869);
and U2513 (N_2513,In_43,In_3349);
nand U2514 (N_2514,In_4405,In_2265);
nand U2515 (N_2515,In_833,In_1539);
or U2516 (N_2516,In_4948,In_143);
or U2517 (N_2517,In_4643,In_1819);
and U2518 (N_2518,In_593,In_4180);
or U2519 (N_2519,In_4476,In_4264);
xnor U2520 (N_2520,In_1898,In_3628);
xor U2521 (N_2521,In_3696,In_4831);
nand U2522 (N_2522,In_1844,In_3996);
nor U2523 (N_2523,In_1152,In_3633);
nand U2524 (N_2524,In_1116,In_2172);
or U2525 (N_2525,In_1005,In_3918);
or U2526 (N_2526,In_4324,In_1059);
or U2527 (N_2527,In_2563,In_2004);
or U2528 (N_2528,In_2449,In_4044);
or U2529 (N_2529,In_475,In_4960);
nor U2530 (N_2530,In_2474,In_2928);
xnor U2531 (N_2531,In_2654,In_3466);
nor U2532 (N_2532,In_2876,In_229);
nor U2533 (N_2533,In_1902,In_4435);
nor U2534 (N_2534,In_2386,In_1612);
nand U2535 (N_2535,In_2405,In_2110);
and U2536 (N_2536,In_3934,In_899);
and U2537 (N_2537,In_2128,In_3088);
and U2538 (N_2538,In_2470,In_4274);
and U2539 (N_2539,In_3412,In_4158);
and U2540 (N_2540,In_4031,In_1780);
or U2541 (N_2541,In_4468,In_2982);
or U2542 (N_2542,In_944,In_4445);
or U2543 (N_2543,In_3879,In_3992);
nand U2544 (N_2544,In_2518,In_4500);
xor U2545 (N_2545,In_4411,In_4784);
and U2546 (N_2546,In_3333,In_267);
xor U2547 (N_2547,In_695,In_4866);
xnor U2548 (N_2548,In_1877,In_2990);
xnor U2549 (N_2549,In_2436,In_2132);
nand U2550 (N_2550,In_4620,In_2985);
or U2551 (N_2551,In_4409,In_4640);
or U2552 (N_2552,In_2415,In_930);
xor U2553 (N_2553,In_204,In_4229);
nand U2554 (N_2554,In_3214,In_4669);
nand U2555 (N_2555,In_4840,In_1930);
and U2556 (N_2556,In_2401,In_2456);
nor U2557 (N_2557,In_780,In_864);
nor U2558 (N_2558,In_4679,In_3802);
nand U2559 (N_2559,In_821,In_970);
xor U2560 (N_2560,In_3966,In_2067);
nand U2561 (N_2561,In_4883,In_4567);
nor U2562 (N_2562,In_4539,In_1324);
and U2563 (N_2563,In_2882,In_3070);
nor U2564 (N_2564,In_2956,In_469);
nor U2565 (N_2565,In_805,In_2855);
and U2566 (N_2566,In_63,In_4713);
xnor U2567 (N_2567,In_3769,In_3060);
nand U2568 (N_2568,In_4899,In_3062);
xnor U2569 (N_2569,In_3750,In_1983);
and U2570 (N_2570,In_2512,In_118);
xnor U2571 (N_2571,In_2315,In_746);
nor U2572 (N_2572,In_355,In_2495);
nand U2573 (N_2573,In_1467,In_4036);
and U2574 (N_2574,In_3493,In_1522);
nor U2575 (N_2575,In_125,In_4154);
nand U2576 (N_2576,In_4279,In_2455);
and U2577 (N_2577,In_496,In_1557);
or U2578 (N_2578,In_3300,In_1871);
and U2579 (N_2579,In_2557,In_370);
nand U2580 (N_2580,In_2802,In_3865);
or U2581 (N_2581,In_3614,In_4303);
nand U2582 (N_2582,In_1724,In_1317);
nor U2583 (N_2583,In_3692,In_1646);
nor U2584 (N_2584,In_238,In_4149);
nand U2585 (N_2585,In_4501,In_2166);
nand U2586 (N_2586,In_4301,In_2244);
or U2587 (N_2587,In_2094,In_4382);
xnor U2588 (N_2588,In_928,In_1486);
nand U2589 (N_2589,In_4987,In_2393);
nor U2590 (N_2590,In_2556,In_4338);
nand U2591 (N_2591,In_4598,In_268);
nand U2592 (N_2592,In_2502,In_4059);
nand U2593 (N_2593,In_3863,In_4681);
nor U2594 (N_2594,In_213,In_724);
nor U2595 (N_2595,In_2754,In_3724);
and U2596 (N_2596,In_743,In_178);
and U2597 (N_2597,In_2370,In_3403);
and U2598 (N_2598,In_4741,In_4215);
or U2599 (N_2599,In_4349,In_2662);
nand U2600 (N_2600,In_2542,In_971);
xor U2601 (N_2601,In_3032,In_2321);
and U2602 (N_2602,In_1897,In_2499);
or U2603 (N_2603,In_3503,In_3871);
or U2604 (N_2604,In_3109,In_509);
nand U2605 (N_2605,In_3355,In_3139);
nor U2606 (N_2606,In_1952,In_2043);
and U2607 (N_2607,In_3402,In_2645);
or U2608 (N_2608,In_899,In_2405);
xor U2609 (N_2609,In_96,In_409);
and U2610 (N_2610,In_555,In_485);
and U2611 (N_2611,In_992,In_4984);
xor U2612 (N_2612,In_3267,In_4898);
and U2613 (N_2613,In_2232,In_4938);
nor U2614 (N_2614,In_3633,In_3327);
or U2615 (N_2615,In_1943,In_4312);
nand U2616 (N_2616,In_1581,In_4380);
or U2617 (N_2617,In_2444,In_3726);
and U2618 (N_2618,In_1470,In_923);
or U2619 (N_2619,In_910,In_3119);
nor U2620 (N_2620,In_4345,In_3305);
nor U2621 (N_2621,In_3366,In_724);
xnor U2622 (N_2622,In_3282,In_4110);
nor U2623 (N_2623,In_4240,In_4648);
or U2624 (N_2624,In_4215,In_4013);
nor U2625 (N_2625,In_80,In_1615);
xnor U2626 (N_2626,In_1510,In_2049);
nand U2627 (N_2627,In_2132,In_4132);
xnor U2628 (N_2628,In_475,In_1059);
nand U2629 (N_2629,In_1233,In_1371);
nor U2630 (N_2630,In_3196,In_2795);
or U2631 (N_2631,In_1490,In_1564);
nor U2632 (N_2632,In_4659,In_1109);
xnor U2633 (N_2633,In_3902,In_545);
and U2634 (N_2634,In_1646,In_2391);
nor U2635 (N_2635,In_302,In_4455);
or U2636 (N_2636,In_1057,In_4760);
nand U2637 (N_2637,In_4432,In_1336);
nand U2638 (N_2638,In_217,In_1524);
or U2639 (N_2639,In_825,In_2900);
xnor U2640 (N_2640,In_3591,In_3954);
or U2641 (N_2641,In_4992,In_1860);
or U2642 (N_2642,In_3080,In_4738);
nor U2643 (N_2643,In_2321,In_4778);
and U2644 (N_2644,In_370,In_1660);
or U2645 (N_2645,In_664,In_4249);
nor U2646 (N_2646,In_3423,In_1100);
xnor U2647 (N_2647,In_1573,In_4608);
nor U2648 (N_2648,In_3521,In_333);
xor U2649 (N_2649,In_2126,In_747);
xnor U2650 (N_2650,In_1241,In_4767);
and U2651 (N_2651,In_1521,In_3877);
nor U2652 (N_2652,In_1182,In_4201);
xnor U2653 (N_2653,In_1805,In_1856);
and U2654 (N_2654,In_4277,In_2174);
or U2655 (N_2655,In_3434,In_3849);
xor U2656 (N_2656,In_609,In_1094);
or U2657 (N_2657,In_3075,In_4000);
nor U2658 (N_2658,In_1749,In_3573);
or U2659 (N_2659,In_830,In_4389);
nand U2660 (N_2660,In_2568,In_2362);
and U2661 (N_2661,In_1624,In_3314);
nor U2662 (N_2662,In_3476,In_1183);
or U2663 (N_2663,In_2217,In_2582);
and U2664 (N_2664,In_4234,In_222);
xor U2665 (N_2665,In_1879,In_4682);
or U2666 (N_2666,In_4227,In_4033);
or U2667 (N_2667,In_976,In_3091);
or U2668 (N_2668,In_1470,In_2464);
and U2669 (N_2669,In_2774,In_614);
xnor U2670 (N_2670,In_94,In_3776);
nand U2671 (N_2671,In_4657,In_1634);
xnor U2672 (N_2672,In_3752,In_467);
nand U2673 (N_2673,In_890,In_108);
or U2674 (N_2674,In_1167,In_4066);
nor U2675 (N_2675,In_728,In_4505);
and U2676 (N_2676,In_4066,In_1025);
nor U2677 (N_2677,In_2197,In_3879);
and U2678 (N_2678,In_777,In_3815);
and U2679 (N_2679,In_3599,In_3901);
nand U2680 (N_2680,In_3134,In_4260);
nor U2681 (N_2681,In_1889,In_2872);
and U2682 (N_2682,In_1238,In_1962);
nand U2683 (N_2683,In_2274,In_1700);
or U2684 (N_2684,In_1633,In_3536);
nor U2685 (N_2685,In_4794,In_3704);
and U2686 (N_2686,In_2128,In_3757);
nor U2687 (N_2687,In_1613,In_40);
and U2688 (N_2688,In_2440,In_3971);
and U2689 (N_2689,In_2861,In_3989);
and U2690 (N_2690,In_1920,In_4694);
xor U2691 (N_2691,In_2063,In_984);
or U2692 (N_2692,In_2231,In_4266);
and U2693 (N_2693,In_2561,In_3849);
and U2694 (N_2694,In_1118,In_1424);
nand U2695 (N_2695,In_3262,In_107);
xnor U2696 (N_2696,In_514,In_2304);
nand U2697 (N_2697,In_402,In_3679);
and U2698 (N_2698,In_3028,In_4423);
xnor U2699 (N_2699,In_1623,In_4227);
and U2700 (N_2700,In_1506,In_1364);
or U2701 (N_2701,In_2560,In_2793);
nand U2702 (N_2702,In_4606,In_2888);
nand U2703 (N_2703,In_2842,In_291);
nor U2704 (N_2704,In_3622,In_3982);
nor U2705 (N_2705,In_2980,In_2841);
or U2706 (N_2706,In_266,In_3065);
nand U2707 (N_2707,In_1288,In_4247);
nor U2708 (N_2708,In_1391,In_91);
nor U2709 (N_2709,In_1324,In_2085);
nor U2710 (N_2710,In_3636,In_3873);
nand U2711 (N_2711,In_4828,In_4283);
xor U2712 (N_2712,In_701,In_3513);
nand U2713 (N_2713,In_3281,In_3988);
nor U2714 (N_2714,In_4257,In_2105);
nor U2715 (N_2715,In_3144,In_4612);
or U2716 (N_2716,In_3844,In_1695);
or U2717 (N_2717,In_848,In_898);
xnor U2718 (N_2718,In_4221,In_4141);
nor U2719 (N_2719,In_3291,In_4102);
xor U2720 (N_2720,In_4385,In_4682);
nor U2721 (N_2721,In_4366,In_1290);
or U2722 (N_2722,In_1074,In_1082);
or U2723 (N_2723,In_4794,In_4191);
nor U2724 (N_2724,In_366,In_729);
xnor U2725 (N_2725,In_2055,In_2407);
or U2726 (N_2726,In_2591,In_2989);
or U2727 (N_2727,In_4637,In_3303);
nor U2728 (N_2728,In_3733,In_3947);
nand U2729 (N_2729,In_3037,In_4569);
nor U2730 (N_2730,In_1718,In_1792);
and U2731 (N_2731,In_3499,In_1720);
and U2732 (N_2732,In_2573,In_2897);
nor U2733 (N_2733,In_699,In_4238);
nor U2734 (N_2734,In_980,In_4166);
xor U2735 (N_2735,In_2030,In_2361);
nor U2736 (N_2736,In_3820,In_451);
nand U2737 (N_2737,In_484,In_269);
or U2738 (N_2738,In_1607,In_3186);
and U2739 (N_2739,In_1324,In_4608);
or U2740 (N_2740,In_1245,In_2048);
or U2741 (N_2741,In_3739,In_3865);
nand U2742 (N_2742,In_4776,In_480);
or U2743 (N_2743,In_4319,In_466);
nand U2744 (N_2744,In_3218,In_1845);
and U2745 (N_2745,In_1663,In_4516);
and U2746 (N_2746,In_4221,In_1109);
or U2747 (N_2747,In_4732,In_4554);
xor U2748 (N_2748,In_2869,In_3701);
or U2749 (N_2749,In_4633,In_2856);
nand U2750 (N_2750,In_1132,In_658);
or U2751 (N_2751,In_1672,In_3720);
nor U2752 (N_2752,In_1827,In_1326);
xor U2753 (N_2753,In_2850,In_1738);
and U2754 (N_2754,In_1775,In_3553);
nand U2755 (N_2755,In_4552,In_3915);
nor U2756 (N_2756,In_2475,In_3394);
xor U2757 (N_2757,In_692,In_3346);
nand U2758 (N_2758,In_2411,In_3218);
nor U2759 (N_2759,In_2982,In_4662);
and U2760 (N_2760,In_594,In_191);
and U2761 (N_2761,In_2414,In_1045);
or U2762 (N_2762,In_4662,In_1856);
or U2763 (N_2763,In_956,In_48);
or U2764 (N_2764,In_638,In_1632);
nand U2765 (N_2765,In_2633,In_2966);
nor U2766 (N_2766,In_1392,In_1478);
nand U2767 (N_2767,In_1028,In_2036);
and U2768 (N_2768,In_244,In_2980);
nor U2769 (N_2769,In_518,In_1439);
xor U2770 (N_2770,In_4162,In_1360);
nor U2771 (N_2771,In_567,In_389);
nor U2772 (N_2772,In_711,In_4131);
or U2773 (N_2773,In_3942,In_599);
nor U2774 (N_2774,In_3271,In_1566);
xnor U2775 (N_2775,In_3534,In_4418);
and U2776 (N_2776,In_1521,In_2128);
or U2777 (N_2777,In_1169,In_3069);
or U2778 (N_2778,In_4156,In_889);
nor U2779 (N_2779,In_2021,In_4861);
and U2780 (N_2780,In_1093,In_438);
or U2781 (N_2781,In_4096,In_4495);
nor U2782 (N_2782,In_1185,In_2138);
nor U2783 (N_2783,In_399,In_4519);
and U2784 (N_2784,In_4731,In_3398);
or U2785 (N_2785,In_343,In_1324);
nor U2786 (N_2786,In_3898,In_4171);
and U2787 (N_2787,In_1526,In_4258);
xnor U2788 (N_2788,In_2121,In_3757);
or U2789 (N_2789,In_3162,In_818);
or U2790 (N_2790,In_2806,In_547);
or U2791 (N_2791,In_4218,In_2332);
or U2792 (N_2792,In_2594,In_4124);
and U2793 (N_2793,In_3365,In_3467);
and U2794 (N_2794,In_3649,In_2515);
and U2795 (N_2795,In_3923,In_679);
xnor U2796 (N_2796,In_4438,In_756);
nand U2797 (N_2797,In_4477,In_4149);
or U2798 (N_2798,In_1726,In_3711);
nand U2799 (N_2799,In_4768,In_438);
xor U2800 (N_2800,In_3677,In_3626);
and U2801 (N_2801,In_1785,In_3191);
nand U2802 (N_2802,In_1846,In_3359);
and U2803 (N_2803,In_598,In_4127);
and U2804 (N_2804,In_1844,In_2975);
and U2805 (N_2805,In_74,In_1712);
or U2806 (N_2806,In_1278,In_4979);
nor U2807 (N_2807,In_1920,In_4370);
nor U2808 (N_2808,In_1293,In_2999);
and U2809 (N_2809,In_3656,In_1447);
nor U2810 (N_2810,In_1337,In_1484);
nand U2811 (N_2811,In_1354,In_2433);
or U2812 (N_2812,In_3964,In_2061);
or U2813 (N_2813,In_2633,In_3244);
or U2814 (N_2814,In_1197,In_1701);
nor U2815 (N_2815,In_145,In_611);
nor U2816 (N_2816,In_3218,In_4336);
and U2817 (N_2817,In_1389,In_4068);
nand U2818 (N_2818,In_2399,In_2899);
xnor U2819 (N_2819,In_1052,In_4069);
nor U2820 (N_2820,In_718,In_715);
nand U2821 (N_2821,In_3986,In_1154);
or U2822 (N_2822,In_3335,In_3569);
or U2823 (N_2823,In_3066,In_3144);
nor U2824 (N_2824,In_2108,In_2617);
or U2825 (N_2825,In_4675,In_1485);
nor U2826 (N_2826,In_2746,In_1623);
xor U2827 (N_2827,In_185,In_1468);
nand U2828 (N_2828,In_2943,In_1698);
nor U2829 (N_2829,In_103,In_4345);
nand U2830 (N_2830,In_4422,In_3017);
and U2831 (N_2831,In_1945,In_2091);
xor U2832 (N_2832,In_1093,In_62);
or U2833 (N_2833,In_2076,In_1148);
nand U2834 (N_2834,In_1498,In_1894);
and U2835 (N_2835,In_896,In_1232);
and U2836 (N_2836,In_3564,In_2220);
nand U2837 (N_2837,In_4433,In_236);
xnor U2838 (N_2838,In_809,In_1839);
nand U2839 (N_2839,In_4742,In_4146);
and U2840 (N_2840,In_1294,In_61);
or U2841 (N_2841,In_2899,In_1905);
xnor U2842 (N_2842,In_2383,In_648);
and U2843 (N_2843,In_575,In_3917);
nand U2844 (N_2844,In_2925,In_2124);
nand U2845 (N_2845,In_593,In_2508);
and U2846 (N_2846,In_2389,In_4078);
nand U2847 (N_2847,In_387,In_1839);
xnor U2848 (N_2848,In_2766,In_1995);
or U2849 (N_2849,In_213,In_3246);
xnor U2850 (N_2850,In_4472,In_4427);
xnor U2851 (N_2851,In_1341,In_3244);
xnor U2852 (N_2852,In_2814,In_311);
and U2853 (N_2853,In_3205,In_918);
and U2854 (N_2854,In_4105,In_566);
and U2855 (N_2855,In_1368,In_4988);
and U2856 (N_2856,In_882,In_4550);
and U2857 (N_2857,In_4886,In_4437);
or U2858 (N_2858,In_2463,In_4110);
or U2859 (N_2859,In_2,In_642);
or U2860 (N_2860,In_2865,In_2475);
or U2861 (N_2861,In_4929,In_4973);
and U2862 (N_2862,In_3856,In_675);
and U2863 (N_2863,In_420,In_4835);
or U2864 (N_2864,In_3492,In_2892);
nor U2865 (N_2865,In_4541,In_1390);
nand U2866 (N_2866,In_528,In_695);
nand U2867 (N_2867,In_3263,In_301);
or U2868 (N_2868,In_1139,In_1312);
nand U2869 (N_2869,In_1573,In_1494);
nand U2870 (N_2870,In_2775,In_3333);
nand U2871 (N_2871,In_234,In_1799);
and U2872 (N_2872,In_3442,In_513);
xor U2873 (N_2873,In_1142,In_713);
nor U2874 (N_2874,In_4785,In_2644);
nor U2875 (N_2875,In_2997,In_1899);
xor U2876 (N_2876,In_4680,In_3862);
nor U2877 (N_2877,In_891,In_3685);
nand U2878 (N_2878,In_4528,In_1124);
xnor U2879 (N_2879,In_2074,In_3795);
nor U2880 (N_2880,In_2478,In_804);
nand U2881 (N_2881,In_4666,In_1928);
nand U2882 (N_2882,In_3309,In_2364);
and U2883 (N_2883,In_2697,In_2848);
nand U2884 (N_2884,In_949,In_4006);
or U2885 (N_2885,In_4796,In_339);
xnor U2886 (N_2886,In_1052,In_1519);
nand U2887 (N_2887,In_4119,In_2081);
and U2888 (N_2888,In_1354,In_4815);
xnor U2889 (N_2889,In_4516,In_4985);
nor U2890 (N_2890,In_495,In_853);
xnor U2891 (N_2891,In_3008,In_3783);
xnor U2892 (N_2892,In_360,In_3335);
nor U2893 (N_2893,In_2826,In_592);
or U2894 (N_2894,In_1909,In_1071);
or U2895 (N_2895,In_3474,In_2287);
xor U2896 (N_2896,In_401,In_1695);
xor U2897 (N_2897,In_1860,In_1491);
xor U2898 (N_2898,In_3637,In_1871);
or U2899 (N_2899,In_4698,In_1110);
and U2900 (N_2900,In_199,In_4382);
nor U2901 (N_2901,In_2344,In_541);
and U2902 (N_2902,In_3088,In_6);
and U2903 (N_2903,In_3818,In_2059);
nand U2904 (N_2904,In_2423,In_1789);
and U2905 (N_2905,In_2601,In_2613);
nand U2906 (N_2906,In_4787,In_2438);
nor U2907 (N_2907,In_2979,In_3729);
nor U2908 (N_2908,In_1623,In_679);
nor U2909 (N_2909,In_4103,In_3069);
or U2910 (N_2910,In_3972,In_515);
xnor U2911 (N_2911,In_1231,In_3141);
or U2912 (N_2912,In_2319,In_3122);
nor U2913 (N_2913,In_3353,In_4395);
or U2914 (N_2914,In_3989,In_1733);
or U2915 (N_2915,In_2598,In_3032);
or U2916 (N_2916,In_1022,In_597);
nand U2917 (N_2917,In_3666,In_4162);
nor U2918 (N_2918,In_4597,In_415);
nand U2919 (N_2919,In_2650,In_4550);
and U2920 (N_2920,In_2901,In_1012);
and U2921 (N_2921,In_4913,In_3662);
and U2922 (N_2922,In_959,In_1332);
or U2923 (N_2923,In_285,In_1781);
and U2924 (N_2924,In_2145,In_0);
or U2925 (N_2925,In_4137,In_1864);
and U2926 (N_2926,In_231,In_828);
and U2927 (N_2927,In_4433,In_3927);
nor U2928 (N_2928,In_2176,In_67);
nor U2929 (N_2929,In_1847,In_2305);
xor U2930 (N_2930,In_3259,In_1612);
or U2931 (N_2931,In_2187,In_2423);
nand U2932 (N_2932,In_3847,In_3391);
nand U2933 (N_2933,In_3661,In_2466);
nor U2934 (N_2934,In_2174,In_2759);
nor U2935 (N_2935,In_3389,In_3751);
nand U2936 (N_2936,In_4380,In_4941);
and U2937 (N_2937,In_854,In_15);
nor U2938 (N_2938,In_1556,In_3334);
nor U2939 (N_2939,In_4727,In_1587);
nand U2940 (N_2940,In_1181,In_3115);
or U2941 (N_2941,In_3379,In_1435);
and U2942 (N_2942,In_1482,In_3308);
nor U2943 (N_2943,In_3068,In_4127);
nand U2944 (N_2944,In_4027,In_2454);
xnor U2945 (N_2945,In_3213,In_4869);
nor U2946 (N_2946,In_2883,In_582);
xor U2947 (N_2947,In_3205,In_1202);
nor U2948 (N_2948,In_782,In_2610);
xor U2949 (N_2949,In_2467,In_2925);
nor U2950 (N_2950,In_2926,In_3079);
nor U2951 (N_2951,In_302,In_4016);
or U2952 (N_2952,In_1656,In_2501);
and U2953 (N_2953,In_2652,In_1694);
nor U2954 (N_2954,In_2892,In_1562);
xor U2955 (N_2955,In_100,In_3301);
xor U2956 (N_2956,In_58,In_2928);
or U2957 (N_2957,In_4872,In_2976);
nand U2958 (N_2958,In_174,In_2180);
or U2959 (N_2959,In_4753,In_1718);
and U2960 (N_2960,In_4660,In_597);
nand U2961 (N_2961,In_2166,In_3587);
or U2962 (N_2962,In_3286,In_763);
xor U2963 (N_2963,In_2043,In_3802);
or U2964 (N_2964,In_4142,In_4225);
or U2965 (N_2965,In_582,In_846);
and U2966 (N_2966,In_2299,In_1175);
nor U2967 (N_2967,In_695,In_2389);
or U2968 (N_2968,In_1398,In_4986);
xor U2969 (N_2969,In_658,In_700);
or U2970 (N_2970,In_532,In_2572);
nand U2971 (N_2971,In_994,In_3654);
nor U2972 (N_2972,In_1404,In_2462);
xnor U2973 (N_2973,In_126,In_4310);
nand U2974 (N_2974,In_912,In_3876);
or U2975 (N_2975,In_3758,In_2202);
nor U2976 (N_2976,In_166,In_1450);
nor U2977 (N_2977,In_2276,In_3268);
or U2978 (N_2978,In_2810,In_3026);
and U2979 (N_2979,In_4710,In_2314);
nand U2980 (N_2980,In_783,In_467);
and U2981 (N_2981,In_3100,In_4845);
and U2982 (N_2982,In_9,In_4575);
xor U2983 (N_2983,In_2299,In_2398);
or U2984 (N_2984,In_3869,In_290);
nor U2985 (N_2985,In_880,In_3712);
and U2986 (N_2986,In_4951,In_392);
or U2987 (N_2987,In_2855,In_2219);
xor U2988 (N_2988,In_2824,In_394);
nand U2989 (N_2989,In_1364,In_2905);
nor U2990 (N_2990,In_4961,In_3656);
nor U2991 (N_2991,In_1692,In_3635);
xnor U2992 (N_2992,In_640,In_4258);
nand U2993 (N_2993,In_2699,In_482);
xnor U2994 (N_2994,In_2205,In_4933);
xor U2995 (N_2995,In_2078,In_2934);
nand U2996 (N_2996,In_2862,In_3914);
or U2997 (N_2997,In_103,In_3136);
nor U2998 (N_2998,In_1825,In_232);
nor U2999 (N_2999,In_1438,In_1029);
or U3000 (N_3000,In_4722,In_2565);
and U3001 (N_3001,In_3000,In_3160);
and U3002 (N_3002,In_1046,In_1232);
nand U3003 (N_3003,In_4950,In_4803);
xnor U3004 (N_3004,In_2576,In_3050);
and U3005 (N_3005,In_4920,In_2789);
xor U3006 (N_3006,In_4682,In_2331);
or U3007 (N_3007,In_1638,In_4545);
or U3008 (N_3008,In_721,In_456);
and U3009 (N_3009,In_981,In_511);
or U3010 (N_3010,In_4773,In_2083);
or U3011 (N_3011,In_2349,In_2907);
xnor U3012 (N_3012,In_4493,In_3701);
or U3013 (N_3013,In_340,In_1531);
nand U3014 (N_3014,In_3054,In_1780);
nand U3015 (N_3015,In_4771,In_4608);
nand U3016 (N_3016,In_2420,In_1739);
and U3017 (N_3017,In_2923,In_294);
or U3018 (N_3018,In_526,In_3608);
nor U3019 (N_3019,In_3814,In_3505);
nand U3020 (N_3020,In_2610,In_4079);
and U3021 (N_3021,In_2630,In_4271);
and U3022 (N_3022,In_1428,In_1934);
and U3023 (N_3023,In_1083,In_327);
xnor U3024 (N_3024,In_4260,In_4295);
or U3025 (N_3025,In_3606,In_1783);
and U3026 (N_3026,In_3871,In_2968);
nor U3027 (N_3027,In_1256,In_1952);
and U3028 (N_3028,In_4635,In_300);
or U3029 (N_3029,In_4267,In_3018);
xnor U3030 (N_3030,In_4674,In_4417);
or U3031 (N_3031,In_2498,In_4725);
or U3032 (N_3032,In_2686,In_2439);
or U3033 (N_3033,In_748,In_1202);
nand U3034 (N_3034,In_536,In_2226);
xor U3035 (N_3035,In_70,In_4993);
nand U3036 (N_3036,In_2229,In_754);
or U3037 (N_3037,In_3129,In_2806);
and U3038 (N_3038,In_1890,In_3668);
and U3039 (N_3039,In_780,In_210);
nor U3040 (N_3040,In_4973,In_4510);
or U3041 (N_3041,In_2508,In_1286);
or U3042 (N_3042,In_3559,In_1455);
nand U3043 (N_3043,In_2334,In_936);
or U3044 (N_3044,In_3130,In_4570);
nor U3045 (N_3045,In_2620,In_456);
and U3046 (N_3046,In_1717,In_3040);
or U3047 (N_3047,In_907,In_501);
nor U3048 (N_3048,In_4641,In_3869);
or U3049 (N_3049,In_4489,In_432);
and U3050 (N_3050,In_4670,In_3549);
and U3051 (N_3051,In_695,In_4264);
nor U3052 (N_3052,In_367,In_2942);
or U3053 (N_3053,In_1643,In_2896);
and U3054 (N_3054,In_498,In_453);
nand U3055 (N_3055,In_4512,In_4350);
nor U3056 (N_3056,In_1278,In_3649);
or U3057 (N_3057,In_1520,In_1157);
or U3058 (N_3058,In_2474,In_4784);
and U3059 (N_3059,In_584,In_464);
and U3060 (N_3060,In_128,In_644);
xnor U3061 (N_3061,In_1657,In_520);
and U3062 (N_3062,In_1797,In_4940);
nand U3063 (N_3063,In_4873,In_557);
nor U3064 (N_3064,In_2624,In_411);
nand U3065 (N_3065,In_74,In_1501);
xor U3066 (N_3066,In_1805,In_498);
nand U3067 (N_3067,In_1138,In_1998);
nor U3068 (N_3068,In_1061,In_4612);
or U3069 (N_3069,In_2121,In_902);
nor U3070 (N_3070,In_4153,In_1300);
and U3071 (N_3071,In_566,In_25);
and U3072 (N_3072,In_4049,In_4563);
or U3073 (N_3073,In_630,In_601);
or U3074 (N_3074,In_660,In_412);
or U3075 (N_3075,In_607,In_2251);
xnor U3076 (N_3076,In_704,In_119);
nand U3077 (N_3077,In_3189,In_4698);
nor U3078 (N_3078,In_4044,In_4891);
nand U3079 (N_3079,In_4683,In_4599);
or U3080 (N_3080,In_144,In_791);
nand U3081 (N_3081,In_4259,In_2320);
and U3082 (N_3082,In_4843,In_3409);
and U3083 (N_3083,In_550,In_948);
nor U3084 (N_3084,In_4651,In_2846);
and U3085 (N_3085,In_4576,In_2657);
or U3086 (N_3086,In_4618,In_2355);
and U3087 (N_3087,In_4917,In_2549);
or U3088 (N_3088,In_4027,In_1614);
or U3089 (N_3089,In_3769,In_89);
or U3090 (N_3090,In_2674,In_4531);
nor U3091 (N_3091,In_1578,In_1355);
and U3092 (N_3092,In_1707,In_712);
nand U3093 (N_3093,In_1260,In_644);
or U3094 (N_3094,In_4185,In_400);
nand U3095 (N_3095,In_4575,In_4940);
xor U3096 (N_3096,In_1788,In_4511);
nand U3097 (N_3097,In_3492,In_707);
and U3098 (N_3098,In_2477,In_1238);
nand U3099 (N_3099,In_4960,In_2517);
nor U3100 (N_3100,In_4656,In_2140);
nand U3101 (N_3101,In_2727,In_2717);
xor U3102 (N_3102,In_4123,In_4874);
nor U3103 (N_3103,In_1242,In_4981);
or U3104 (N_3104,In_828,In_891);
and U3105 (N_3105,In_4566,In_2314);
xor U3106 (N_3106,In_835,In_531);
or U3107 (N_3107,In_3313,In_4628);
or U3108 (N_3108,In_4806,In_1558);
nor U3109 (N_3109,In_1819,In_222);
xnor U3110 (N_3110,In_3902,In_2083);
xnor U3111 (N_3111,In_1426,In_3761);
nand U3112 (N_3112,In_151,In_2909);
nor U3113 (N_3113,In_1263,In_3320);
or U3114 (N_3114,In_792,In_2315);
and U3115 (N_3115,In_4136,In_2323);
nand U3116 (N_3116,In_97,In_1025);
or U3117 (N_3117,In_1053,In_2571);
and U3118 (N_3118,In_2837,In_2467);
or U3119 (N_3119,In_3600,In_3236);
and U3120 (N_3120,In_1795,In_978);
and U3121 (N_3121,In_2015,In_4756);
nand U3122 (N_3122,In_3577,In_3622);
and U3123 (N_3123,In_3791,In_2140);
nand U3124 (N_3124,In_3471,In_1786);
nand U3125 (N_3125,In_1568,In_3502);
or U3126 (N_3126,In_3883,In_822);
or U3127 (N_3127,In_2149,In_2923);
and U3128 (N_3128,In_791,In_265);
xnor U3129 (N_3129,In_3,In_723);
nand U3130 (N_3130,In_4074,In_396);
nor U3131 (N_3131,In_2125,In_1764);
nor U3132 (N_3132,In_3658,In_3720);
or U3133 (N_3133,In_4080,In_2562);
and U3134 (N_3134,In_2656,In_3978);
nand U3135 (N_3135,In_4957,In_2911);
xnor U3136 (N_3136,In_3075,In_3762);
nand U3137 (N_3137,In_2295,In_2016);
xor U3138 (N_3138,In_915,In_1022);
and U3139 (N_3139,In_3024,In_4009);
nand U3140 (N_3140,In_525,In_1015);
and U3141 (N_3141,In_3214,In_1832);
xor U3142 (N_3142,In_1455,In_2370);
and U3143 (N_3143,In_4385,In_1937);
and U3144 (N_3144,In_1928,In_1878);
xnor U3145 (N_3145,In_1736,In_1254);
nor U3146 (N_3146,In_2433,In_4515);
nand U3147 (N_3147,In_2063,In_2917);
or U3148 (N_3148,In_4609,In_3287);
or U3149 (N_3149,In_3969,In_3145);
or U3150 (N_3150,In_3688,In_940);
nand U3151 (N_3151,In_3988,In_2076);
or U3152 (N_3152,In_3666,In_3047);
nor U3153 (N_3153,In_725,In_3277);
and U3154 (N_3154,In_4326,In_4769);
nand U3155 (N_3155,In_37,In_1199);
and U3156 (N_3156,In_2927,In_3462);
xor U3157 (N_3157,In_2635,In_3578);
nor U3158 (N_3158,In_41,In_140);
nand U3159 (N_3159,In_2301,In_2183);
and U3160 (N_3160,In_2014,In_4923);
and U3161 (N_3161,In_3548,In_4240);
nor U3162 (N_3162,In_4725,In_1768);
nand U3163 (N_3163,In_1369,In_1791);
or U3164 (N_3164,In_4176,In_2138);
nand U3165 (N_3165,In_1160,In_3379);
xor U3166 (N_3166,In_1806,In_4349);
nor U3167 (N_3167,In_4147,In_2639);
and U3168 (N_3168,In_4361,In_3657);
and U3169 (N_3169,In_3788,In_129);
and U3170 (N_3170,In_3009,In_3450);
xor U3171 (N_3171,In_1976,In_3290);
or U3172 (N_3172,In_2332,In_4012);
and U3173 (N_3173,In_3596,In_4398);
xnor U3174 (N_3174,In_1284,In_3662);
nor U3175 (N_3175,In_2217,In_88);
nor U3176 (N_3176,In_88,In_3426);
nor U3177 (N_3177,In_1858,In_3289);
nor U3178 (N_3178,In_3662,In_2302);
nand U3179 (N_3179,In_1080,In_240);
or U3180 (N_3180,In_1930,In_3682);
nand U3181 (N_3181,In_4116,In_2255);
and U3182 (N_3182,In_1961,In_3863);
nor U3183 (N_3183,In_1060,In_4559);
xor U3184 (N_3184,In_2436,In_3453);
and U3185 (N_3185,In_1423,In_4398);
or U3186 (N_3186,In_869,In_4562);
xnor U3187 (N_3187,In_3429,In_3628);
nand U3188 (N_3188,In_269,In_1514);
nand U3189 (N_3189,In_1138,In_4603);
xor U3190 (N_3190,In_2881,In_2068);
nor U3191 (N_3191,In_1620,In_4857);
and U3192 (N_3192,In_4137,In_1518);
and U3193 (N_3193,In_3134,In_4762);
xnor U3194 (N_3194,In_466,In_1506);
nand U3195 (N_3195,In_3807,In_1095);
nand U3196 (N_3196,In_4103,In_2303);
and U3197 (N_3197,In_4434,In_1154);
or U3198 (N_3198,In_1296,In_963);
xnor U3199 (N_3199,In_4200,In_2927);
xor U3200 (N_3200,In_4373,In_140);
or U3201 (N_3201,In_4243,In_3507);
nor U3202 (N_3202,In_4851,In_4535);
nor U3203 (N_3203,In_1802,In_875);
and U3204 (N_3204,In_1428,In_3115);
or U3205 (N_3205,In_1880,In_4658);
nand U3206 (N_3206,In_2520,In_2474);
nor U3207 (N_3207,In_1355,In_2726);
nor U3208 (N_3208,In_236,In_2232);
or U3209 (N_3209,In_1412,In_916);
or U3210 (N_3210,In_1347,In_3938);
and U3211 (N_3211,In_3051,In_459);
xor U3212 (N_3212,In_149,In_3965);
and U3213 (N_3213,In_3826,In_2427);
xnor U3214 (N_3214,In_1720,In_3795);
nor U3215 (N_3215,In_2927,In_4249);
nand U3216 (N_3216,In_4356,In_402);
xnor U3217 (N_3217,In_717,In_4830);
xor U3218 (N_3218,In_4618,In_3908);
xor U3219 (N_3219,In_4862,In_3687);
and U3220 (N_3220,In_559,In_3398);
and U3221 (N_3221,In_4046,In_3399);
or U3222 (N_3222,In_3913,In_3459);
nand U3223 (N_3223,In_2100,In_4115);
and U3224 (N_3224,In_4132,In_2544);
xnor U3225 (N_3225,In_4502,In_4378);
xnor U3226 (N_3226,In_1921,In_1881);
nor U3227 (N_3227,In_2638,In_2766);
and U3228 (N_3228,In_1042,In_2816);
or U3229 (N_3229,In_4767,In_84);
nand U3230 (N_3230,In_1570,In_1245);
nand U3231 (N_3231,In_2296,In_3087);
and U3232 (N_3232,In_3994,In_2139);
or U3233 (N_3233,In_4610,In_3652);
xor U3234 (N_3234,In_3133,In_3680);
nor U3235 (N_3235,In_3780,In_3470);
nand U3236 (N_3236,In_54,In_2121);
nor U3237 (N_3237,In_418,In_4773);
and U3238 (N_3238,In_4702,In_2496);
nand U3239 (N_3239,In_3832,In_4515);
and U3240 (N_3240,In_1779,In_2103);
nor U3241 (N_3241,In_2713,In_924);
or U3242 (N_3242,In_2658,In_4890);
nand U3243 (N_3243,In_4844,In_2805);
nand U3244 (N_3244,In_4123,In_1243);
xnor U3245 (N_3245,In_1169,In_2051);
and U3246 (N_3246,In_3990,In_4767);
or U3247 (N_3247,In_4544,In_633);
nand U3248 (N_3248,In_2177,In_570);
nand U3249 (N_3249,In_3977,In_3165);
and U3250 (N_3250,In_784,In_573);
and U3251 (N_3251,In_3348,In_2747);
nor U3252 (N_3252,In_4338,In_2761);
nand U3253 (N_3253,In_1834,In_417);
xnor U3254 (N_3254,In_2525,In_520);
nor U3255 (N_3255,In_4217,In_2926);
nor U3256 (N_3256,In_3777,In_2351);
and U3257 (N_3257,In_3429,In_3298);
nand U3258 (N_3258,In_1889,In_4674);
nor U3259 (N_3259,In_3955,In_2203);
or U3260 (N_3260,In_70,In_154);
or U3261 (N_3261,In_4634,In_2626);
nor U3262 (N_3262,In_289,In_2863);
nand U3263 (N_3263,In_2730,In_2094);
nand U3264 (N_3264,In_4150,In_1546);
nor U3265 (N_3265,In_1080,In_962);
nor U3266 (N_3266,In_3189,In_69);
or U3267 (N_3267,In_2791,In_3996);
nand U3268 (N_3268,In_1545,In_4384);
nand U3269 (N_3269,In_281,In_3824);
and U3270 (N_3270,In_4898,In_3237);
nor U3271 (N_3271,In_2310,In_4504);
nand U3272 (N_3272,In_4577,In_4778);
nand U3273 (N_3273,In_1075,In_4542);
nor U3274 (N_3274,In_4610,In_1721);
nor U3275 (N_3275,In_4338,In_1257);
or U3276 (N_3276,In_242,In_1327);
and U3277 (N_3277,In_2803,In_3993);
nand U3278 (N_3278,In_3454,In_4719);
and U3279 (N_3279,In_194,In_3850);
and U3280 (N_3280,In_1698,In_213);
nor U3281 (N_3281,In_2473,In_519);
and U3282 (N_3282,In_4828,In_4316);
nor U3283 (N_3283,In_1797,In_3799);
or U3284 (N_3284,In_1361,In_637);
or U3285 (N_3285,In_3779,In_1536);
nor U3286 (N_3286,In_1790,In_4459);
nor U3287 (N_3287,In_4013,In_1573);
and U3288 (N_3288,In_109,In_719);
or U3289 (N_3289,In_222,In_827);
xor U3290 (N_3290,In_4670,In_3072);
xor U3291 (N_3291,In_1437,In_490);
nor U3292 (N_3292,In_861,In_3245);
xnor U3293 (N_3293,In_2930,In_4290);
and U3294 (N_3294,In_1184,In_3108);
and U3295 (N_3295,In_4790,In_4374);
nor U3296 (N_3296,In_4771,In_1259);
and U3297 (N_3297,In_2822,In_4825);
nor U3298 (N_3298,In_1726,In_1497);
nor U3299 (N_3299,In_1410,In_343);
nor U3300 (N_3300,In_590,In_0);
and U3301 (N_3301,In_3420,In_3907);
nand U3302 (N_3302,In_2222,In_2364);
nand U3303 (N_3303,In_4629,In_1932);
or U3304 (N_3304,In_2115,In_2199);
nand U3305 (N_3305,In_1586,In_1384);
or U3306 (N_3306,In_4389,In_4466);
nor U3307 (N_3307,In_4809,In_827);
xnor U3308 (N_3308,In_3443,In_1102);
xor U3309 (N_3309,In_373,In_1175);
xnor U3310 (N_3310,In_3879,In_1173);
and U3311 (N_3311,In_298,In_4418);
nor U3312 (N_3312,In_3229,In_2169);
and U3313 (N_3313,In_2732,In_1095);
and U3314 (N_3314,In_479,In_1151);
and U3315 (N_3315,In_1229,In_3105);
xnor U3316 (N_3316,In_1633,In_235);
or U3317 (N_3317,In_3846,In_474);
xnor U3318 (N_3318,In_1049,In_118);
or U3319 (N_3319,In_3471,In_3544);
nand U3320 (N_3320,In_235,In_1666);
nand U3321 (N_3321,In_2007,In_871);
and U3322 (N_3322,In_1390,In_3273);
xnor U3323 (N_3323,In_104,In_2448);
and U3324 (N_3324,In_3097,In_4897);
nand U3325 (N_3325,In_602,In_2208);
nor U3326 (N_3326,In_4624,In_4634);
xnor U3327 (N_3327,In_1972,In_4452);
nor U3328 (N_3328,In_242,In_2796);
nand U3329 (N_3329,In_3661,In_3185);
and U3330 (N_3330,In_3554,In_2033);
and U3331 (N_3331,In_177,In_940);
and U3332 (N_3332,In_380,In_4672);
or U3333 (N_3333,In_340,In_4324);
xnor U3334 (N_3334,In_4533,In_1039);
or U3335 (N_3335,In_4818,In_3768);
xor U3336 (N_3336,In_2222,In_1203);
or U3337 (N_3337,In_2650,In_4206);
nor U3338 (N_3338,In_3107,In_1976);
or U3339 (N_3339,In_3512,In_3567);
xor U3340 (N_3340,In_3133,In_4293);
and U3341 (N_3341,In_3258,In_2678);
nand U3342 (N_3342,In_462,In_1717);
nor U3343 (N_3343,In_2566,In_4825);
xnor U3344 (N_3344,In_1968,In_4190);
or U3345 (N_3345,In_373,In_1543);
or U3346 (N_3346,In_3808,In_3836);
or U3347 (N_3347,In_4814,In_1264);
and U3348 (N_3348,In_678,In_3991);
and U3349 (N_3349,In_741,In_2954);
nand U3350 (N_3350,In_1520,In_2420);
nand U3351 (N_3351,In_4499,In_4257);
or U3352 (N_3352,In_3052,In_3706);
and U3353 (N_3353,In_679,In_230);
nand U3354 (N_3354,In_4410,In_4362);
and U3355 (N_3355,In_264,In_4297);
nand U3356 (N_3356,In_3259,In_1526);
and U3357 (N_3357,In_3469,In_3184);
and U3358 (N_3358,In_3713,In_4975);
and U3359 (N_3359,In_3005,In_140);
xnor U3360 (N_3360,In_4113,In_621);
nand U3361 (N_3361,In_4647,In_4557);
nor U3362 (N_3362,In_2048,In_1954);
nor U3363 (N_3363,In_3314,In_2878);
and U3364 (N_3364,In_348,In_1584);
nor U3365 (N_3365,In_2882,In_2001);
nor U3366 (N_3366,In_1058,In_4145);
and U3367 (N_3367,In_1966,In_1368);
and U3368 (N_3368,In_3137,In_786);
nand U3369 (N_3369,In_3867,In_4835);
nand U3370 (N_3370,In_3747,In_405);
nand U3371 (N_3371,In_1271,In_4359);
or U3372 (N_3372,In_1923,In_909);
or U3373 (N_3373,In_3350,In_3842);
or U3374 (N_3374,In_343,In_1054);
and U3375 (N_3375,In_1362,In_1716);
nor U3376 (N_3376,In_310,In_1715);
and U3377 (N_3377,In_3541,In_1682);
and U3378 (N_3378,In_4527,In_395);
xnor U3379 (N_3379,In_3472,In_2733);
or U3380 (N_3380,In_1529,In_3014);
nand U3381 (N_3381,In_3266,In_4103);
nor U3382 (N_3382,In_3354,In_2078);
nor U3383 (N_3383,In_4920,In_4159);
nand U3384 (N_3384,In_1769,In_1830);
nand U3385 (N_3385,In_669,In_1913);
nor U3386 (N_3386,In_1352,In_3567);
and U3387 (N_3387,In_1852,In_4876);
nor U3388 (N_3388,In_1800,In_3633);
xnor U3389 (N_3389,In_4762,In_2378);
nor U3390 (N_3390,In_2726,In_1791);
nand U3391 (N_3391,In_1949,In_1571);
xor U3392 (N_3392,In_618,In_280);
nor U3393 (N_3393,In_3474,In_4156);
and U3394 (N_3394,In_4315,In_877);
xnor U3395 (N_3395,In_14,In_3526);
and U3396 (N_3396,In_1898,In_1757);
nor U3397 (N_3397,In_612,In_2212);
and U3398 (N_3398,In_1092,In_343);
xor U3399 (N_3399,In_1027,In_3534);
nand U3400 (N_3400,In_3944,In_86);
and U3401 (N_3401,In_2028,In_2390);
xnor U3402 (N_3402,In_1097,In_4362);
nor U3403 (N_3403,In_2404,In_4239);
or U3404 (N_3404,In_1104,In_1186);
and U3405 (N_3405,In_4604,In_1260);
xnor U3406 (N_3406,In_2178,In_3033);
and U3407 (N_3407,In_3004,In_2712);
xnor U3408 (N_3408,In_2077,In_1371);
nor U3409 (N_3409,In_2173,In_3779);
nand U3410 (N_3410,In_130,In_3708);
nand U3411 (N_3411,In_4830,In_3829);
or U3412 (N_3412,In_996,In_3366);
or U3413 (N_3413,In_181,In_4761);
and U3414 (N_3414,In_3574,In_384);
or U3415 (N_3415,In_3109,In_3062);
or U3416 (N_3416,In_1981,In_4655);
or U3417 (N_3417,In_2283,In_570);
xor U3418 (N_3418,In_38,In_814);
nor U3419 (N_3419,In_4857,In_3796);
nand U3420 (N_3420,In_3059,In_2164);
or U3421 (N_3421,In_3188,In_3720);
and U3422 (N_3422,In_4918,In_1777);
and U3423 (N_3423,In_593,In_1313);
and U3424 (N_3424,In_3407,In_4644);
nand U3425 (N_3425,In_686,In_650);
nand U3426 (N_3426,In_1647,In_2058);
nor U3427 (N_3427,In_535,In_2055);
nand U3428 (N_3428,In_3260,In_42);
or U3429 (N_3429,In_279,In_1451);
xnor U3430 (N_3430,In_3699,In_2027);
and U3431 (N_3431,In_3894,In_311);
nand U3432 (N_3432,In_291,In_4861);
nand U3433 (N_3433,In_2627,In_2915);
xnor U3434 (N_3434,In_981,In_4933);
xnor U3435 (N_3435,In_3919,In_1111);
and U3436 (N_3436,In_4830,In_3268);
or U3437 (N_3437,In_4583,In_4664);
xnor U3438 (N_3438,In_2824,In_4297);
nand U3439 (N_3439,In_4751,In_457);
or U3440 (N_3440,In_4654,In_3407);
xor U3441 (N_3441,In_2782,In_4270);
xor U3442 (N_3442,In_2763,In_3793);
xor U3443 (N_3443,In_72,In_3514);
nand U3444 (N_3444,In_1430,In_1496);
and U3445 (N_3445,In_4785,In_2878);
and U3446 (N_3446,In_676,In_4112);
nand U3447 (N_3447,In_16,In_3851);
nand U3448 (N_3448,In_590,In_760);
nor U3449 (N_3449,In_4357,In_4849);
xnor U3450 (N_3450,In_2636,In_2139);
nand U3451 (N_3451,In_4115,In_1914);
xor U3452 (N_3452,In_4571,In_1959);
nor U3453 (N_3453,In_2038,In_595);
and U3454 (N_3454,In_3554,In_620);
nand U3455 (N_3455,In_500,In_2051);
or U3456 (N_3456,In_1133,In_3777);
nor U3457 (N_3457,In_3643,In_4654);
and U3458 (N_3458,In_2617,In_1014);
nor U3459 (N_3459,In_4849,In_901);
nand U3460 (N_3460,In_4587,In_4271);
nor U3461 (N_3461,In_336,In_3523);
or U3462 (N_3462,In_3145,In_1448);
nand U3463 (N_3463,In_2111,In_1237);
nor U3464 (N_3464,In_2543,In_2495);
xnor U3465 (N_3465,In_1736,In_3923);
xnor U3466 (N_3466,In_3816,In_2101);
xnor U3467 (N_3467,In_1798,In_1848);
xnor U3468 (N_3468,In_1996,In_4745);
and U3469 (N_3469,In_4524,In_4969);
and U3470 (N_3470,In_70,In_3979);
xnor U3471 (N_3471,In_3763,In_1791);
or U3472 (N_3472,In_876,In_3824);
and U3473 (N_3473,In_4330,In_2961);
xor U3474 (N_3474,In_2576,In_2997);
xor U3475 (N_3475,In_3315,In_1487);
or U3476 (N_3476,In_3296,In_527);
or U3477 (N_3477,In_3687,In_1130);
or U3478 (N_3478,In_1776,In_3618);
or U3479 (N_3479,In_2509,In_284);
or U3480 (N_3480,In_978,In_2048);
and U3481 (N_3481,In_1631,In_4805);
or U3482 (N_3482,In_2768,In_4053);
or U3483 (N_3483,In_4156,In_1674);
nand U3484 (N_3484,In_3988,In_4116);
nand U3485 (N_3485,In_706,In_3068);
nand U3486 (N_3486,In_4316,In_1764);
xnor U3487 (N_3487,In_2971,In_3236);
xnor U3488 (N_3488,In_2850,In_1661);
nor U3489 (N_3489,In_1608,In_4044);
or U3490 (N_3490,In_632,In_504);
or U3491 (N_3491,In_3479,In_4384);
nor U3492 (N_3492,In_187,In_3490);
or U3493 (N_3493,In_212,In_3242);
nor U3494 (N_3494,In_1328,In_1228);
xnor U3495 (N_3495,In_4667,In_4960);
and U3496 (N_3496,In_471,In_206);
nor U3497 (N_3497,In_4339,In_1582);
nor U3498 (N_3498,In_2110,In_4361);
or U3499 (N_3499,In_4178,In_2539);
and U3500 (N_3500,In_3750,In_400);
or U3501 (N_3501,In_1209,In_456);
and U3502 (N_3502,In_2901,In_4762);
or U3503 (N_3503,In_1667,In_3572);
nor U3504 (N_3504,In_1678,In_1878);
nand U3505 (N_3505,In_2489,In_3394);
nor U3506 (N_3506,In_4220,In_626);
and U3507 (N_3507,In_1599,In_423);
xor U3508 (N_3508,In_2624,In_3094);
xnor U3509 (N_3509,In_4275,In_4705);
xor U3510 (N_3510,In_2868,In_708);
nor U3511 (N_3511,In_1369,In_1670);
or U3512 (N_3512,In_3338,In_4432);
xor U3513 (N_3513,In_1934,In_3250);
or U3514 (N_3514,In_3335,In_4552);
or U3515 (N_3515,In_1968,In_3155);
xor U3516 (N_3516,In_1937,In_58);
xnor U3517 (N_3517,In_4112,In_1346);
and U3518 (N_3518,In_3061,In_2727);
or U3519 (N_3519,In_4655,In_1553);
nor U3520 (N_3520,In_4087,In_2837);
nor U3521 (N_3521,In_4146,In_1430);
or U3522 (N_3522,In_1738,In_4315);
xnor U3523 (N_3523,In_2696,In_2627);
nor U3524 (N_3524,In_4885,In_2543);
nor U3525 (N_3525,In_1920,In_2140);
and U3526 (N_3526,In_3768,In_4263);
nor U3527 (N_3527,In_767,In_3439);
or U3528 (N_3528,In_2568,In_1937);
and U3529 (N_3529,In_147,In_3657);
nand U3530 (N_3530,In_3088,In_1841);
nand U3531 (N_3531,In_4886,In_382);
nand U3532 (N_3532,In_3471,In_3330);
xnor U3533 (N_3533,In_1801,In_3660);
and U3534 (N_3534,In_4131,In_3001);
and U3535 (N_3535,In_3836,In_3455);
or U3536 (N_3536,In_4544,In_4129);
or U3537 (N_3537,In_4226,In_3581);
or U3538 (N_3538,In_3600,In_422);
nor U3539 (N_3539,In_379,In_2508);
or U3540 (N_3540,In_1982,In_389);
and U3541 (N_3541,In_1974,In_2291);
nand U3542 (N_3542,In_3064,In_4262);
xor U3543 (N_3543,In_3312,In_3401);
nand U3544 (N_3544,In_1011,In_4678);
xor U3545 (N_3545,In_4896,In_4628);
and U3546 (N_3546,In_4618,In_2487);
or U3547 (N_3547,In_1521,In_2313);
xor U3548 (N_3548,In_2391,In_2883);
xnor U3549 (N_3549,In_4803,In_4555);
and U3550 (N_3550,In_4267,In_2304);
and U3551 (N_3551,In_3150,In_4725);
nor U3552 (N_3552,In_4330,In_3234);
xor U3553 (N_3553,In_3985,In_4801);
nor U3554 (N_3554,In_338,In_441);
xor U3555 (N_3555,In_784,In_3708);
xor U3556 (N_3556,In_2608,In_1132);
and U3557 (N_3557,In_4422,In_226);
nor U3558 (N_3558,In_552,In_2471);
nor U3559 (N_3559,In_167,In_3590);
nor U3560 (N_3560,In_1001,In_966);
or U3561 (N_3561,In_4348,In_671);
nand U3562 (N_3562,In_633,In_2783);
nor U3563 (N_3563,In_2383,In_2505);
or U3564 (N_3564,In_4831,In_697);
nand U3565 (N_3565,In_2118,In_2051);
xnor U3566 (N_3566,In_103,In_2607);
xnor U3567 (N_3567,In_1321,In_1372);
nor U3568 (N_3568,In_3781,In_3631);
xor U3569 (N_3569,In_478,In_640);
or U3570 (N_3570,In_1403,In_1769);
and U3571 (N_3571,In_3159,In_3733);
and U3572 (N_3572,In_3295,In_871);
nor U3573 (N_3573,In_1477,In_4924);
nand U3574 (N_3574,In_105,In_2088);
nand U3575 (N_3575,In_1624,In_1125);
xnor U3576 (N_3576,In_79,In_431);
xnor U3577 (N_3577,In_3337,In_3710);
xor U3578 (N_3578,In_1640,In_3972);
nor U3579 (N_3579,In_1378,In_669);
xnor U3580 (N_3580,In_4823,In_4405);
and U3581 (N_3581,In_281,In_1257);
xnor U3582 (N_3582,In_3262,In_588);
nor U3583 (N_3583,In_3939,In_3918);
nor U3584 (N_3584,In_2604,In_681);
and U3585 (N_3585,In_688,In_0);
and U3586 (N_3586,In_3617,In_2790);
nand U3587 (N_3587,In_858,In_3290);
xor U3588 (N_3588,In_1564,In_1163);
nand U3589 (N_3589,In_375,In_3027);
or U3590 (N_3590,In_2756,In_4928);
and U3591 (N_3591,In_3427,In_959);
nand U3592 (N_3592,In_3810,In_2307);
nor U3593 (N_3593,In_4692,In_2957);
and U3594 (N_3594,In_4024,In_779);
xnor U3595 (N_3595,In_2428,In_1107);
nand U3596 (N_3596,In_3056,In_2779);
nand U3597 (N_3597,In_2562,In_1742);
nand U3598 (N_3598,In_2248,In_2741);
nor U3599 (N_3599,In_1285,In_1143);
nand U3600 (N_3600,In_1076,In_2907);
nor U3601 (N_3601,In_4094,In_4018);
xor U3602 (N_3602,In_3141,In_2466);
nand U3603 (N_3603,In_1624,In_4191);
and U3604 (N_3604,In_3449,In_1036);
xor U3605 (N_3605,In_3076,In_203);
and U3606 (N_3606,In_3454,In_2078);
nor U3607 (N_3607,In_1860,In_4747);
or U3608 (N_3608,In_3301,In_46);
and U3609 (N_3609,In_254,In_3724);
xor U3610 (N_3610,In_2007,In_3274);
nor U3611 (N_3611,In_3088,In_4536);
or U3612 (N_3612,In_1855,In_2122);
or U3613 (N_3613,In_2336,In_2083);
xnor U3614 (N_3614,In_3304,In_2241);
nand U3615 (N_3615,In_331,In_4066);
nand U3616 (N_3616,In_703,In_2825);
and U3617 (N_3617,In_1169,In_530);
nor U3618 (N_3618,In_285,In_2425);
nand U3619 (N_3619,In_3402,In_3481);
and U3620 (N_3620,In_1532,In_1744);
nand U3621 (N_3621,In_819,In_4945);
or U3622 (N_3622,In_699,In_816);
nor U3623 (N_3623,In_898,In_1165);
or U3624 (N_3624,In_314,In_3322);
nor U3625 (N_3625,In_4440,In_4813);
or U3626 (N_3626,In_788,In_4366);
and U3627 (N_3627,In_4918,In_892);
and U3628 (N_3628,In_2692,In_3447);
nand U3629 (N_3629,In_611,In_454);
or U3630 (N_3630,In_643,In_2450);
and U3631 (N_3631,In_1848,In_4212);
nand U3632 (N_3632,In_1403,In_1564);
xnor U3633 (N_3633,In_1628,In_3879);
xnor U3634 (N_3634,In_808,In_2596);
nor U3635 (N_3635,In_3418,In_4423);
nor U3636 (N_3636,In_4798,In_4331);
and U3637 (N_3637,In_3517,In_452);
nand U3638 (N_3638,In_548,In_2975);
nand U3639 (N_3639,In_2070,In_103);
nor U3640 (N_3640,In_4678,In_1848);
nand U3641 (N_3641,In_1900,In_763);
xnor U3642 (N_3642,In_1987,In_1221);
and U3643 (N_3643,In_3138,In_3155);
or U3644 (N_3644,In_1966,In_4880);
or U3645 (N_3645,In_4428,In_20);
or U3646 (N_3646,In_3834,In_4463);
nand U3647 (N_3647,In_1456,In_183);
xnor U3648 (N_3648,In_852,In_2932);
xor U3649 (N_3649,In_3525,In_453);
nand U3650 (N_3650,In_2541,In_1055);
nor U3651 (N_3651,In_4795,In_4866);
or U3652 (N_3652,In_2818,In_232);
and U3653 (N_3653,In_2312,In_615);
nor U3654 (N_3654,In_632,In_3835);
or U3655 (N_3655,In_4160,In_3904);
and U3656 (N_3656,In_3891,In_2005);
xnor U3657 (N_3657,In_2723,In_1500);
xnor U3658 (N_3658,In_1113,In_2119);
or U3659 (N_3659,In_1108,In_1608);
or U3660 (N_3660,In_1248,In_3947);
xor U3661 (N_3661,In_3634,In_4607);
nand U3662 (N_3662,In_1252,In_3321);
xnor U3663 (N_3663,In_3941,In_4260);
and U3664 (N_3664,In_1076,In_2951);
nand U3665 (N_3665,In_2974,In_3490);
xnor U3666 (N_3666,In_1313,In_3640);
xnor U3667 (N_3667,In_86,In_3242);
nand U3668 (N_3668,In_2648,In_1299);
nand U3669 (N_3669,In_4675,In_4625);
and U3670 (N_3670,In_3294,In_4499);
nor U3671 (N_3671,In_2985,In_2407);
or U3672 (N_3672,In_859,In_74);
nand U3673 (N_3673,In_950,In_775);
and U3674 (N_3674,In_611,In_3462);
and U3675 (N_3675,In_3682,In_4504);
nor U3676 (N_3676,In_2422,In_1662);
nand U3677 (N_3677,In_1458,In_4155);
or U3678 (N_3678,In_4106,In_387);
nor U3679 (N_3679,In_2454,In_2619);
and U3680 (N_3680,In_3652,In_4417);
xor U3681 (N_3681,In_80,In_2209);
xor U3682 (N_3682,In_4765,In_855);
nand U3683 (N_3683,In_242,In_211);
nor U3684 (N_3684,In_148,In_946);
xnor U3685 (N_3685,In_3689,In_2513);
xor U3686 (N_3686,In_2546,In_4963);
nand U3687 (N_3687,In_2,In_1146);
or U3688 (N_3688,In_4280,In_4564);
nand U3689 (N_3689,In_1304,In_602);
or U3690 (N_3690,In_1831,In_3817);
nor U3691 (N_3691,In_4632,In_1428);
nor U3692 (N_3692,In_2102,In_15);
nand U3693 (N_3693,In_2324,In_1241);
and U3694 (N_3694,In_697,In_1995);
or U3695 (N_3695,In_2106,In_638);
or U3696 (N_3696,In_2313,In_619);
or U3697 (N_3697,In_3720,In_4248);
nor U3698 (N_3698,In_3756,In_947);
and U3699 (N_3699,In_3293,In_3053);
xnor U3700 (N_3700,In_1681,In_2297);
or U3701 (N_3701,In_3891,In_267);
xor U3702 (N_3702,In_4148,In_2303);
xnor U3703 (N_3703,In_2225,In_463);
and U3704 (N_3704,In_3806,In_2547);
xor U3705 (N_3705,In_1297,In_4978);
or U3706 (N_3706,In_1129,In_3890);
nand U3707 (N_3707,In_4530,In_1272);
xor U3708 (N_3708,In_1867,In_393);
nand U3709 (N_3709,In_883,In_3303);
nand U3710 (N_3710,In_3509,In_2188);
or U3711 (N_3711,In_4358,In_1770);
nor U3712 (N_3712,In_1151,In_4875);
and U3713 (N_3713,In_2617,In_4340);
xnor U3714 (N_3714,In_1617,In_3791);
xnor U3715 (N_3715,In_1011,In_4987);
nor U3716 (N_3716,In_580,In_3326);
or U3717 (N_3717,In_4297,In_4585);
xor U3718 (N_3718,In_1330,In_4782);
nor U3719 (N_3719,In_3326,In_25);
nor U3720 (N_3720,In_2935,In_4725);
and U3721 (N_3721,In_4420,In_1327);
xnor U3722 (N_3722,In_4030,In_2750);
or U3723 (N_3723,In_3957,In_290);
nand U3724 (N_3724,In_4043,In_3315);
nor U3725 (N_3725,In_4332,In_4533);
nor U3726 (N_3726,In_1627,In_2556);
nand U3727 (N_3727,In_1347,In_2073);
and U3728 (N_3728,In_331,In_3329);
xor U3729 (N_3729,In_4980,In_2197);
and U3730 (N_3730,In_3296,In_4520);
and U3731 (N_3731,In_4444,In_1998);
or U3732 (N_3732,In_2054,In_3512);
nand U3733 (N_3733,In_1467,In_3433);
xor U3734 (N_3734,In_2405,In_1250);
nand U3735 (N_3735,In_151,In_1842);
and U3736 (N_3736,In_2314,In_2954);
xor U3737 (N_3737,In_1708,In_1252);
nor U3738 (N_3738,In_2407,In_3358);
nor U3739 (N_3739,In_4928,In_834);
or U3740 (N_3740,In_444,In_1432);
or U3741 (N_3741,In_838,In_3408);
nand U3742 (N_3742,In_1802,In_4980);
nand U3743 (N_3743,In_3671,In_2221);
or U3744 (N_3744,In_1550,In_4904);
and U3745 (N_3745,In_2309,In_2561);
and U3746 (N_3746,In_3380,In_18);
xor U3747 (N_3747,In_2001,In_4761);
xor U3748 (N_3748,In_2722,In_3925);
and U3749 (N_3749,In_4725,In_1272);
or U3750 (N_3750,In_653,In_1100);
nor U3751 (N_3751,In_2757,In_1180);
or U3752 (N_3752,In_3509,In_2504);
or U3753 (N_3753,In_3250,In_1836);
xnor U3754 (N_3754,In_3761,In_516);
xor U3755 (N_3755,In_1299,In_1114);
xor U3756 (N_3756,In_3678,In_1136);
and U3757 (N_3757,In_3631,In_2320);
nor U3758 (N_3758,In_615,In_1073);
nand U3759 (N_3759,In_2431,In_3807);
and U3760 (N_3760,In_683,In_1578);
and U3761 (N_3761,In_4271,In_2019);
xnor U3762 (N_3762,In_1106,In_3786);
nor U3763 (N_3763,In_4608,In_3149);
nor U3764 (N_3764,In_3711,In_3481);
and U3765 (N_3765,In_1443,In_2681);
and U3766 (N_3766,In_2400,In_4547);
xor U3767 (N_3767,In_3739,In_3233);
nor U3768 (N_3768,In_358,In_3076);
xor U3769 (N_3769,In_3908,In_3334);
xnor U3770 (N_3770,In_852,In_3165);
or U3771 (N_3771,In_2117,In_4566);
and U3772 (N_3772,In_3098,In_2747);
nor U3773 (N_3773,In_4753,In_4871);
nor U3774 (N_3774,In_1646,In_4031);
nor U3775 (N_3775,In_49,In_3013);
xor U3776 (N_3776,In_3133,In_4660);
or U3777 (N_3777,In_4759,In_3532);
or U3778 (N_3778,In_2889,In_4149);
xor U3779 (N_3779,In_2539,In_4135);
and U3780 (N_3780,In_1104,In_701);
or U3781 (N_3781,In_3343,In_1858);
xnor U3782 (N_3782,In_536,In_3938);
xor U3783 (N_3783,In_1345,In_2658);
and U3784 (N_3784,In_993,In_1384);
nand U3785 (N_3785,In_1207,In_3423);
or U3786 (N_3786,In_4258,In_626);
and U3787 (N_3787,In_3539,In_1691);
nand U3788 (N_3788,In_3818,In_331);
and U3789 (N_3789,In_341,In_2031);
nor U3790 (N_3790,In_3143,In_1843);
nor U3791 (N_3791,In_977,In_3114);
and U3792 (N_3792,In_3702,In_2066);
or U3793 (N_3793,In_2411,In_2060);
and U3794 (N_3794,In_4037,In_3982);
nor U3795 (N_3795,In_1619,In_1726);
nand U3796 (N_3796,In_1740,In_2354);
xor U3797 (N_3797,In_3542,In_4215);
nand U3798 (N_3798,In_1911,In_3980);
or U3799 (N_3799,In_4408,In_4622);
xnor U3800 (N_3800,In_1999,In_3248);
and U3801 (N_3801,In_2802,In_2758);
and U3802 (N_3802,In_4325,In_4745);
or U3803 (N_3803,In_2496,In_756);
nor U3804 (N_3804,In_1594,In_3213);
nor U3805 (N_3805,In_1591,In_2805);
or U3806 (N_3806,In_4575,In_2882);
xor U3807 (N_3807,In_2342,In_1910);
nor U3808 (N_3808,In_3132,In_1885);
nand U3809 (N_3809,In_1277,In_3808);
or U3810 (N_3810,In_3974,In_1162);
nand U3811 (N_3811,In_458,In_1832);
xnor U3812 (N_3812,In_4929,In_4648);
xor U3813 (N_3813,In_4238,In_4134);
nor U3814 (N_3814,In_3831,In_4942);
xor U3815 (N_3815,In_4752,In_3703);
xor U3816 (N_3816,In_2769,In_1850);
nor U3817 (N_3817,In_444,In_4630);
xnor U3818 (N_3818,In_409,In_567);
nand U3819 (N_3819,In_4569,In_2594);
nor U3820 (N_3820,In_3845,In_3183);
nand U3821 (N_3821,In_2836,In_1173);
xnor U3822 (N_3822,In_1489,In_500);
xor U3823 (N_3823,In_697,In_1334);
and U3824 (N_3824,In_1428,In_117);
and U3825 (N_3825,In_3119,In_1543);
or U3826 (N_3826,In_588,In_2366);
xnor U3827 (N_3827,In_2041,In_977);
nand U3828 (N_3828,In_4508,In_1544);
or U3829 (N_3829,In_730,In_709);
xnor U3830 (N_3830,In_2498,In_3775);
nor U3831 (N_3831,In_1465,In_1587);
xor U3832 (N_3832,In_3468,In_2720);
or U3833 (N_3833,In_1874,In_2130);
and U3834 (N_3834,In_4547,In_1396);
or U3835 (N_3835,In_1007,In_48);
nor U3836 (N_3836,In_3321,In_706);
or U3837 (N_3837,In_2554,In_4696);
or U3838 (N_3838,In_278,In_2979);
xor U3839 (N_3839,In_1922,In_3571);
nand U3840 (N_3840,In_973,In_1618);
and U3841 (N_3841,In_1127,In_1414);
and U3842 (N_3842,In_3808,In_3814);
and U3843 (N_3843,In_4495,In_4921);
nor U3844 (N_3844,In_1680,In_4988);
or U3845 (N_3845,In_4758,In_1759);
nor U3846 (N_3846,In_4338,In_654);
or U3847 (N_3847,In_3867,In_2772);
nand U3848 (N_3848,In_2571,In_3666);
nor U3849 (N_3849,In_4129,In_2941);
xor U3850 (N_3850,In_1112,In_1817);
xor U3851 (N_3851,In_2969,In_3159);
and U3852 (N_3852,In_505,In_770);
nor U3853 (N_3853,In_2147,In_3771);
xor U3854 (N_3854,In_4301,In_2893);
and U3855 (N_3855,In_1990,In_2797);
nor U3856 (N_3856,In_2712,In_1179);
nand U3857 (N_3857,In_3449,In_1515);
or U3858 (N_3858,In_4120,In_3819);
xor U3859 (N_3859,In_2776,In_3802);
or U3860 (N_3860,In_1132,In_3255);
xor U3861 (N_3861,In_4844,In_4597);
nand U3862 (N_3862,In_2829,In_4280);
and U3863 (N_3863,In_2144,In_45);
nand U3864 (N_3864,In_1504,In_2164);
and U3865 (N_3865,In_1249,In_1496);
nor U3866 (N_3866,In_2736,In_749);
nor U3867 (N_3867,In_4867,In_2829);
or U3868 (N_3868,In_3999,In_3606);
nor U3869 (N_3869,In_4105,In_1563);
xor U3870 (N_3870,In_2684,In_2236);
nand U3871 (N_3871,In_1646,In_4029);
nand U3872 (N_3872,In_4785,In_2212);
or U3873 (N_3873,In_2201,In_2607);
or U3874 (N_3874,In_1455,In_928);
or U3875 (N_3875,In_4664,In_4732);
and U3876 (N_3876,In_4961,In_1409);
or U3877 (N_3877,In_3197,In_1223);
or U3878 (N_3878,In_348,In_3418);
nand U3879 (N_3879,In_3743,In_3375);
xnor U3880 (N_3880,In_2144,In_4754);
or U3881 (N_3881,In_253,In_3408);
or U3882 (N_3882,In_1715,In_3269);
nor U3883 (N_3883,In_4604,In_260);
xnor U3884 (N_3884,In_2216,In_2830);
or U3885 (N_3885,In_2945,In_4787);
nor U3886 (N_3886,In_2065,In_3174);
nand U3887 (N_3887,In_885,In_3053);
xnor U3888 (N_3888,In_2976,In_2038);
xnor U3889 (N_3889,In_3978,In_1481);
and U3890 (N_3890,In_2520,In_2937);
nand U3891 (N_3891,In_2386,In_1645);
xnor U3892 (N_3892,In_2854,In_4417);
xor U3893 (N_3893,In_2223,In_3054);
or U3894 (N_3894,In_3055,In_3537);
nor U3895 (N_3895,In_3608,In_2869);
xor U3896 (N_3896,In_4710,In_4371);
or U3897 (N_3897,In_3210,In_414);
nor U3898 (N_3898,In_3434,In_4790);
xnor U3899 (N_3899,In_117,In_605);
nand U3900 (N_3900,In_2251,In_119);
and U3901 (N_3901,In_867,In_2170);
nor U3902 (N_3902,In_808,In_4606);
or U3903 (N_3903,In_4059,In_1163);
nand U3904 (N_3904,In_4015,In_1564);
and U3905 (N_3905,In_617,In_1532);
or U3906 (N_3906,In_4532,In_3512);
nand U3907 (N_3907,In_78,In_189);
and U3908 (N_3908,In_1490,In_684);
nand U3909 (N_3909,In_2124,In_4546);
nand U3910 (N_3910,In_3379,In_3139);
xor U3911 (N_3911,In_2861,In_187);
and U3912 (N_3912,In_4483,In_2478);
nor U3913 (N_3913,In_77,In_856);
and U3914 (N_3914,In_2183,In_3193);
xnor U3915 (N_3915,In_4277,In_2247);
xor U3916 (N_3916,In_3463,In_1322);
or U3917 (N_3917,In_1374,In_4393);
and U3918 (N_3918,In_2102,In_2861);
nand U3919 (N_3919,In_3673,In_674);
nand U3920 (N_3920,In_128,In_2613);
and U3921 (N_3921,In_3216,In_2515);
xnor U3922 (N_3922,In_4962,In_2098);
nor U3923 (N_3923,In_2313,In_587);
xnor U3924 (N_3924,In_883,In_2709);
xor U3925 (N_3925,In_89,In_1527);
or U3926 (N_3926,In_1548,In_3574);
nand U3927 (N_3927,In_620,In_1603);
xnor U3928 (N_3928,In_2262,In_4392);
nor U3929 (N_3929,In_2677,In_1143);
nor U3930 (N_3930,In_196,In_1572);
nor U3931 (N_3931,In_1630,In_2245);
nor U3932 (N_3932,In_3877,In_2038);
nor U3933 (N_3933,In_2787,In_2465);
or U3934 (N_3934,In_4610,In_4509);
or U3935 (N_3935,In_4067,In_3822);
xor U3936 (N_3936,In_553,In_4929);
and U3937 (N_3937,In_2918,In_4802);
and U3938 (N_3938,In_887,In_670);
nor U3939 (N_3939,In_622,In_3047);
nand U3940 (N_3940,In_720,In_3211);
nand U3941 (N_3941,In_117,In_1255);
or U3942 (N_3942,In_2671,In_1927);
nor U3943 (N_3943,In_1159,In_1344);
and U3944 (N_3944,In_645,In_3580);
nand U3945 (N_3945,In_3631,In_4819);
and U3946 (N_3946,In_3439,In_2005);
or U3947 (N_3947,In_4418,In_630);
xor U3948 (N_3948,In_2426,In_3117);
xnor U3949 (N_3949,In_2699,In_3287);
nor U3950 (N_3950,In_3030,In_1080);
and U3951 (N_3951,In_898,In_640);
and U3952 (N_3952,In_4600,In_914);
nor U3953 (N_3953,In_1572,In_288);
nor U3954 (N_3954,In_4422,In_3158);
or U3955 (N_3955,In_4286,In_1135);
nor U3956 (N_3956,In_2993,In_4673);
nor U3957 (N_3957,In_1897,In_2288);
nor U3958 (N_3958,In_3963,In_2195);
or U3959 (N_3959,In_1212,In_4126);
nor U3960 (N_3960,In_1072,In_3480);
and U3961 (N_3961,In_997,In_4216);
nor U3962 (N_3962,In_2065,In_4557);
nor U3963 (N_3963,In_2517,In_1011);
or U3964 (N_3964,In_3593,In_1897);
and U3965 (N_3965,In_3378,In_2807);
nor U3966 (N_3966,In_4748,In_2145);
nand U3967 (N_3967,In_3505,In_779);
nand U3968 (N_3968,In_3564,In_647);
and U3969 (N_3969,In_2089,In_1911);
and U3970 (N_3970,In_2005,In_3803);
xor U3971 (N_3971,In_3806,In_2322);
and U3972 (N_3972,In_1310,In_3577);
or U3973 (N_3973,In_578,In_1732);
nand U3974 (N_3974,In_1873,In_1667);
nor U3975 (N_3975,In_1351,In_2172);
nor U3976 (N_3976,In_3800,In_2626);
nand U3977 (N_3977,In_2067,In_3261);
or U3978 (N_3978,In_3512,In_1614);
or U3979 (N_3979,In_2421,In_269);
or U3980 (N_3980,In_3632,In_2134);
and U3981 (N_3981,In_1060,In_4754);
and U3982 (N_3982,In_2039,In_2060);
and U3983 (N_3983,In_2543,In_1841);
xor U3984 (N_3984,In_4471,In_3120);
or U3985 (N_3985,In_1758,In_2947);
and U3986 (N_3986,In_3854,In_1241);
xnor U3987 (N_3987,In_1942,In_2788);
nor U3988 (N_3988,In_862,In_1284);
xor U3989 (N_3989,In_1980,In_4944);
and U3990 (N_3990,In_2376,In_890);
and U3991 (N_3991,In_3943,In_1762);
or U3992 (N_3992,In_959,In_3007);
xnor U3993 (N_3993,In_1769,In_4104);
nand U3994 (N_3994,In_3847,In_1781);
xnor U3995 (N_3995,In_2354,In_1591);
and U3996 (N_3996,In_4942,In_1539);
nor U3997 (N_3997,In_4670,In_1506);
nand U3998 (N_3998,In_992,In_2476);
nor U3999 (N_3999,In_2977,In_533);
nand U4000 (N_4000,In_74,In_3398);
nor U4001 (N_4001,In_1951,In_1453);
nand U4002 (N_4002,In_4856,In_2576);
nor U4003 (N_4003,In_2862,In_4639);
or U4004 (N_4004,In_1786,In_5);
nand U4005 (N_4005,In_1738,In_107);
and U4006 (N_4006,In_718,In_4808);
xnor U4007 (N_4007,In_1888,In_746);
or U4008 (N_4008,In_2895,In_2251);
nand U4009 (N_4009,In_4753,In_4410);
and U4010 (N_4010,In_4178,In_1405);
xor U4011 (N_4011,In_152,In_621);
xnor U4012 (N_4012,In_3936,In_1130);
or U4013 (N_4013,In_1300,In_1725);
nor U4014 (N_4014,In_2251,In_2348);
or U4015 (N_4015,In_4827,In_1122);
and U4016 (N_4016,In_1335,In_998);
or U4017 (N_4017,In_2223,In_2691);
or U4018 (N_4018,In_2315,In_2826);
or U4019 (N_4019,In_2680,In_2386);
or U4020 (N_4020,In_3071,In_379);
nand U4021 (N_4021,In_4731,In_3937);
nand U4022 (N_4022,In_3023,In_1477);
nor U4023 (N_4023,In_3268,In_48);
nand U4024 (N_4024,In_4083,In_1929);
nand U4025 (N_4025,In_1926,In_4345);
nor U4026 (N_4026,In_3720,In_3775);
or U4027 (N_4027,In_3825,In_657);
nor U4028 (N_4028,In_469,In_4717);
or U4029 (N_4029,In_3015,In_3951);
xnor U4030 (N_4030,In_2891,In_2876);
and U4031 (N_4031,In_2415,In_525);
and U4032 (N_4032,In_1274,In_2293);
or U4033 (N_4033,In_3528,In_3360);
and U4034 (N_4034,In_4341,In_3072);
nand U4035 (N_4035,In_4164,In_1452);
xor U4036 (N_4036,In_474,In_4043);
nand U4037 (N_4037,In_1662,In_1953);
nor U4038 (N_4038,In_1849,In_1042);
nand U4039 (N_4039,In_4391,In_2413);
and U4040 (N_4040,In_1416,In_2979);
and U4041 (N_4041,In_3989,In_4909);
and U4042 (N_4042,In_3730,In_1093);
nor U4043 (N_4043,In_2636,In_918);
or U4044 (N_4044,In_220,In_345);
and U4045 (N_4045,In_3164,In_3286);
nor U4046 (N_4046,In_2973,In_2480);
nor U4047 (N_4047,In_3727,In_3308);
or U4048 (N_4048,In_1798,In_4460);
xor U4049 (N_4049,In_486,In_2813);
or U4050 (N_4050,In_4112,In_4870);
nand U4051 (N_4051,In_899,In_3625);
nand U4052 (N_4052,In_2991,In_1715);
nand U4053 (N_4053,In_4958,In_4077);
xor U4054 (N_4054,In_1341,In_4373);
and U4055 (N_4055,In_1052,In_3131);
xnor U4056 (N_4056,In_2756,In_2286);
xor U4057 (N_4057,In_4701,In_3531);
xnor U4058 (N_4058,In_755,In_2453);
and U4059 (N_4059,In_3987,In_3815);
or U4060 (N_4060,In_3918,In_3685);
nand U4061 (N_4061,In_2523,In_767);
or U4062 (N_4062,In_3151,In_236);
nand U4063 (N_4063,In_3921,In_1993);
nand U4064 (N_4064,In_3059,In_4630);
xnor U4065 (N_4065,In_2794,In_4309);
and U4066 (N_4066,In_4996,In_950);
nand U4067 (N_4067,In_109,In_1214);
and U4068 (N_4068,In_3665,In_3672);
nand U4069 (N_4069,In_617,In_3101);
nand U4070 (N_4070,In_2450,In_1275);
or U4071 (N_4071,In_1447,In_3401);
nand U4072 (N_4072,In_2040,In_3964);
xor U4073 (N_4073,In_3616,In_4215);
nor U4074 (N_4074,In_3369,In_283);
xor U4075 (N_4075,In_2471,In_3124);
xnor U4076 (N_4076,In_97,In_243);
or U4077 (N_4077,In_602,In_4967);
xnor U4078 (N_4078,In_4971,In_1470);
nand U4079 (N_4079,In_2981,In_2368);
nor U4080 (N_4080,In_4210,In_1678);
and U4081 (N_4081,In_1548,In_4627);
nor U4082 (N_4082,In_3756,In_1511);
or U4083 (N_4083,In_4886,In_3599);
nand U4084 (N_4084,In_2921,In_1876);
xnor U4085 (N_4085,In_4782,In_2265);
nand U4086 (N_4086,In_501,In_1435);
or U4087 (N_4087,In_1257,In_1191);
nor U4088 (N_4088,In_4693,In_2935);
xnor U4089 (N_4089,In_2491,In_2383);
xnor U4090 (N_4090,In_1428,In_2181);
and U4091 (N_4091,In_1034,In_470);
and U4092 (N_4092,In_131,In_2696);
and U4093 (N_4093,In_3847,In_2638);
nand U4094 (N_4094,In_224,In_1348);
or U4095 (N_4095,In_2372,In_201);
nand U4096 (N_4096,In_1587,In_2158);
xnor U4097 (N_4097,In_4756,In_3884);
and U4098 (N_4098,In_1348,In_1776);
nor U4099 (N_4099,In_4528,In_1566);
nand U4100 (N_4100,In_1955,In_4162);
nor U4101 (N_4101,In_1748,In_4710);
or U4102 (N_4102,In_1896,In_3546);
or U4103 (N_4103,In_717,In_1704);
and U4104 (N_4104,In_739,In_4008);
nand U4105 (N_4105,In_35,In_624);
xnor U4106 (N_4106,In_4021,In_3417);
nor U4107 (N_4107,In_3073,In_2476);
xnor U4108 (N_4108,In_3340,In_3132);
or U4109 (N_4109,In_3534,In_3946);
nand U4110 (N_4110,In_1190,In_911);
nand U4111 (N_4111,In_172,In_1209);
nor U4112 (N_4112,In_560,In_1346);
nand U4113 (N_4113,In_102,In_3161);
or U4114 (N_4114,In_3293,In_4709);
nand U4115 (N_4115,In_3445,In_4280);
xor U4116 (N_4116,In_4967,In_1606);
or U4117 (N_4117,In_1313,In_4066);
xnor U4118 (N_4118,In_223,In_1213);
and U4119 (N_4119,In_3417,In_3251);
xnor U4120 (N_4120,In_2342,In_1892);
nor U4121 (N_4121,In_1300,In_1677);
xor U4122 (N_4122,In_4058,In_2381);
and U4123 (N_4123,In_2879,In_1011);
nand U4124 (N_4124,In_3196,In_852);
xor U4125 (N_4125,In_3806,In_830);
and U4126 (N_4126,In_1666,In_4387);
nor U4127 (N_4127,In_15,In_4564);
xor U4128 (N_4128,In_2558,In_472);
xor U4129 (N_4129,In_3413,In_4037);
xnor U4130 (N_4130,In_2782,In_2397);
and U4131 (N_4131,In_1448,In_2775);
and U4132 (N_4132,In_3823,In_2345);
nand U4133 (N_4133,In_1049,In_4477);
nand U4134 (N_4134,In_4302,In_3991);
nor U4135 (N_4135,In_1301,In_424);
nand U4136 (N_4136,In_3428,In_3866);
xnor U4137 (N_4137,In_2110,In_535);
xor U4138 (N_4138,In_3854,In_4907);
or U4139 (N_4139,In_52,In_2699);
xor U4140 (N_4140,In_1623,In_2940);
and U4141 (N_4141,In_1598,In_1258);
and U4142 (N_4142,In_2430,In_4333);
nand U4143 (N_4143,In_4040,In_4290);
and U4144 (N_4144,In_2179,In_782);
nand U4145 (N_4145,In_1077,In_4845);
nand U4146 (N_4146,In_1167,In_3734);
nand U4147 (N_4147,In_2531,In_1269);
xnor U4148 (N_4148,In_3372,In_3650);
xor U4149 (N_4149,In_3572,In_1430);
nor U4150 (N_4150,In_4549,In_1813);
or U4151 (N_4151,In_827,In_682);
nor U4152 (N_4152,In_2673,In_2893);
nand U4153 (N_4153,In_3686,In_4782);
and U4154 (N_4154,In_4417,In_2422);
and U4155 (N_4155,In_1506,In_4069);
nand U4156 (N_4156,In_1694,In_923);
nand U4157 (N_4157,In_1703,In_2466);
xor U4158 (N_4158,In_3634,In_2777);
or U4159 (N_4159,In_1951,In_4327);
and U4160 (N_4160,In_4824,In_3649);
nand U4161 (N_4161,In_3091,In_4238);
nor U4162 (N_4162,In_4439,In_1424);
nand U4163 (N_4163,In_1955,In_3280);
nor U4164 (N_4164,In_2961,In_1936);
nor U4165 (N_4165,In_4853,In_4458);
and U4166 (N_4166,In_973,In_3726);
nor U4167 (N_4167,In_3525,In_4456);
and U4168 (N_4168,In_4475,In_2222);
and U4169 (N_4169,In_1012,In_4607);
or U4170 (N_4170,In_3184,In_2885);
or U4171 (N_4171,In_1799,In_4653);
xnor U4172 (N_4172,In_3875,In_2699);
nand U4173 (N_4173,In_920,In_1551);
nor U4174 (N_4174,In_2436,In_2846);
and U4175 (N_4175,In_4347,In_2073);
or U4176 (N_4176,In_3738,In_1532);
and U4177 (N_4177,In_2583,In_3367);
nor U4178 (N_4178,In_2575,In_3924);
xor U4179 (N_4179,In_3037,In_2484);
xor U4180 (N_4180,In_1632,In_2176);
nand U4181 (N_4181,In_3800,In_3554);
or U4182 (N_4182,In_2101,In_1589);
xnor U4183 (N_4183,In_4314,In_1674);
or U4184 (N_4184,In_1936,In_4123);
nor U4185 (N_4185,In_2193,In_3870);
xor U4186 (N_4186,In_3926,In_2955);
nand U4187 (N_4187,In_1704,In_3792);
xor U4188 (N_4188,In_2683,In_2503);
or U4189 (N_4189,In_4673,In_2247);
xor U4190 (N_4190,In_166,In_2414);
nor U4191 (N_4191,In_4934,In_2292);
nand U4192 (N_4192,In_4516,In_128);
nor U4193 (N_4193,In_1532,In_4879);
and U4194 (N_4194,In_1530,In_4948);
or U4195 (N_4195,In_1680,In_204);
nor U4196 (N_4196,In_242,In_3674);
xnor U4197 (N_4197,In_225,In_3562);
nand U4198 (N_4198,In_214,In_3809);
and U4199 (N_4199,In_2136,In_4339);
nor U4200 (N_4200,In_3271,In_3630);
xor U4201 (N_4201,In_2170,In_2349);
and U4202 (N_4202,In_2505,In_3434);
nand U4203 (N_4203,In_3310,In_899);
nor U4204 (N_4204,In_1526,In_1636);
nand U4205 (N_4205,In_2649,In_694);
xnor U4206 (N_4206,In_4761,In_681);
nand U4207 (N_4207,In_4226,In_4598);
and U4208 (N_4208,In_927,In_4133);
and U4209 (N_4209,In_1981,In_3657);
or U4210 (N_4210,In_3546,In_2457);
and U4211 (N_4211,In_617,In_3936);
xnor U4212 (N_4212,In_4151,In_4288);
xnor U4213 (N_4213,In_3356,In_4572);
or U4214 (N_4214,In_4272,In_3450);
or U4215 (N_4215,In_1170,In_1422);
nor U4216 (N_4216,In_736,In_370);
nand U4217 (N_4217,In_3799,In_120);
or U4218 (N_4218,In_4373,In_463);
and U4219 (N_4219,In_1887,In_3303);
nand U4220 (N_4220,In_2038,In_2965);
or U4221 (N_4221,In_4747,In_2999);
nor U4222 (N_4222,In_1543,In_1308);
nand U4223 (N_4223,In_2827,In_4130);
xnor U4224 (N_4224,In_4237,In_3824);
nand U4225 (N_4225,In_2005,In_3113);
xnor U4226 (N_4226,In_4445,In_1354);
nor U4227 (N_4227,In_4893,In_4810);
and U4228 (N_4228,In_3471,In_1159);
and U4229 (N_4229,In_3526,In_3136);
and U4230 (N_4230,In_2406,In_4390);
nand U4231 (N_4231,In_4660,In_74);
or U4232 (N_4232,In_1743,In_3214);
or U4233 (N_4233,In_2703,In_81);
or U4234 (N_4234,In_2442,In_3472);
xor U4235 (N_4235,In_4408,In_1037);
nor U4236 (N_4236,In_1912,In_4695);
and U4237 (N_4237,In_1779,In_4042);
nor U4238 (N_4238,In_2324,In_1023);
nor U4239 (N_4239,In_3468,In_3274);
nand U4240 (N_4240,In_2810,In_2351);
nand U4241 (N_4241,In_453,In_1380);
xnor U4242 (N_4242,In_669,In_493);
and U4243 (N_4243,In_4857,In_2404);
xor U4244 (N_4244,In_4826,In_3830);
or U4245 (N_4245,In_2864,In_2890);
and U4246 (N_4246,In_4404,In_2070);
and U4247 (N_4247,In_4248,In_2153);
and U4248 (N_4248,In_1330,In_4244);
xor U4249 (N_4249,In_3509,In_858);
and U4250 (N_4250,In_1554,In_705);
nor U4251 (N_4251,In_2403,In_3450);
or U4252 (N_4252,In_4986,In_4577);
xor U4253 (N_4253,In_3895,In_2094);
xnor U4254 (N_4254,In_1598,In_167);
or U4255 (N_4255,In_462,In_2349);
nor U4256 (N_4256,In_3444,In_4563);
or U4257 (N_4257,In_4729,In_1346);
or U4258 (N_4258,In_0,In_3698);
or U4259 (N_4259,In_737,In_3624);
nor U4260 (N_4260,In_2582,In_3151);
nand U4261 (N_4261,In_2592,In_4890);
nor U4262 (N_4262,In_1004,In_4598);
nand U4263 (N_4263,In_1799,In_483);
nor U4264 (N_4264,In_670,In_1137);
nand U4265 (N_4265,In_1081,In_2071);
nand U4266 (N_4266,In_1398,In_914);
or U4267 (N_4267,In_3419,In_847);
nor U4268 (N_4268,In_3891,In_1851);
nor U4269 (N_4269,In_3128,In_1709);
nor U4270 (N_4270,In_3039,In_4741);
xor U4271 (N_4271,In_4317,In_1865);
or U4272 (N_4272,In_2289,In_681);
nand U4273 (N_4273,In_4283,In_1812);
xor U4274 (N_4274,In_3453,In_3906);
or U4275 (N_4275,In_4830,In_652);
nand U4276 (N_4276,In_3617,In_4561);
nand U4277 (N_4277,In_4079,In_949);
or U4278 (N_4278,In_2875,In_3655);
or U4279 (N_4279,In_2884,In_2462);
xnor U4280 (N_4280,In_2802,In_1773);
or U4281 (N_4281,In_4499,In_463);
xor U4282 (N_4282,In_669,In_4);
nor U4283 (N_4283,In_2520,In_956);
xnor U4284 (N_4284,In_1859,In_626);
and U4285 (N_4285,In_2033,In_2762);
nand U4286 (N_4286,In_3631,In_1493);
or U4287 (N_4287,In_2128,In_1830);
xor U4288 (N_4288,In_2094,In_146);
nor U4289 (N_4289,In_1466,In_363);
or U4290 (N_4290,In_3835,In_269);
or U4291 (N_4291,In_4341,In_563);
and U4292 (N_4292,In_4097,In_20);
and U4293 (N_4293,In_2892,In_1636);
nand U4294 (N_4294,In_507,In_4481);
and U4295 (N_4295,In_4040,In_3844);
nor U4296 (N_4296,In_2290,In_171);
nor U4297 (N_4297,In_2373,In_4404);
nand U4298 (N_4298,In_3459,In_1735);
xor U4299 (N_4299,In_725,In_1641);
nand U4300 (N_4300,In_1055,In_4828);
and U4301 (N_4301,In_2819,In_2879);
nor U4302 (N_4302,In_4709,In_232);
or U4303 (N_4303,In_82,In_3944);
nor U4304 (N_4304,In_3477,In_1600);
xor U4305 (N_4305,In_226,In_914);
nand U4306 (N_4306,In_3893,In_441);
xnor U4307 (N_4307,In_2100,In_256);
or U4308 (N_4308,In_4793,In_1241);
or U4309 (N_4309,In_3954,In_3729);
xor U4310 (N_4310,In_4747,In_859);
or U4311 (N_4311,In_1149,In_4534);
and U4312 (N_4312,In_2452,In_588);
xor U4313 (N_4313,In_1219,In_4283);
xnor U4314 (N_4314,In_2947,In_1259);
nand U4315 (N_4315,In_1231,In_573);
xor U4316 (N_4316,In_1250,In_2185);
nand U4317 (N_4317,In_3597,In_2229);
xor U4318 (N_4318,In_4073,In_646);
xor U4319 (N_4319,In_3445,In_1232);
xnor U4320 (N_4320,In_4215,In_817);
and U4321 (N_4321,In_4680,In_3814);
nand U4322 (N_4322,In_3327,In_4396);
or U4323 (N_4323,In_2857,In_4804);
nand U4324 (N_4324,In_4358,In_1687);
and U4325 (N_4325,In_4377,In_1263);
or U4326 (N_4326,In_1422,In_572);
and U4327 (N_4327,In_1486,In_3666);
nor U4328 (N_4328,In_929,In_1907);
or U4329 (N_4329,In_565,In_3782);
nor U4330 (N_4330,In_1373,In_2571);
or U4331 (N_4331,In_2306,In_1119);
xor U4332 (N_4332,In_97,In_4900);
or U4333 (N_4333,In_490,In_3067);
nand U4334 (N_4334,In_1203,In_2371);
xor U4335 (N_4335,In_2416,In_3652);
nand U4336 (N_4336,In_1364,In_4833);
nor U4337 (N_4337,In_729,In_717);
or U4338 (N_4338,In_1252,In_1249);
and U4339 (N_4339,In_2627,In_3553);
or U4340 (N_4340,In_4987,In_4955);
or U4341 (N_4341,In_2234,In_3073);
xor U4342 (N_4342,In_4940,In_99);
xor U4343 (N_4343,In_308,In_627);
xor U4344 (N_4344,In_1386,In_3689);
xnor U4345 (N_4345,In_3886,In_2357);
or U4346 (N_4346,In_3323,In_3435);
nand U4347 (N_4347,In_1006,In_2565);
nand U4348 (N_4348,In_2531,In_603);
nor U4349 (N_4349,In_3325,In_1345);
nand U4350 (N_4350,In_749,In_2223);
nand U4351 (N_4351,In_3827,In_4383);
xnor U4352 (N_4352,In_3744,In_4113);
and U4353 (N_4353,In_2153,In_1493);
or U4354 (N_4354,In_1936,In_1443);
nand U4355 (N_4355,In_3340,In_3535);
xor U4356 (N_4356,In_3822,In_2244);
and U4357 (N_4357,In_4498,In_1560);
and U4358 (N_4358,In_3095,In_1423);
nand U4359 (N_4359,In_2298,In_583);
nor U4360 (N_4360,In_4715,In_2516);
or U4361 (N_4361,In_2951,In_1494);
and U4362 (N_4362,In_3143,In_2776);
or U4363 (N_4363,In_4968,In_4675);
nor U4364 (N_4364,In_1587,In_1124);
nor U4365 (N_4365,In_139,In_462);
or U4366 (N_4366,In_1054,In_741);
nor U4367 (N_4367,In_4149,In_4936);
nand U4368 (N_4368,In_1814,In_641);
xor U4369 (N_4369,In_2884,In_1427);
nand U4370 (N_4370,In_2324,In_1962);
and U4371 (N_4371,In_3086,In_158);
or U4372 (N_4372,In_1058,In_2912);
and U4373 (N_4373,In_1475,In_262);
nor U4374 (N_4374,In_216,In_3151);
and U4375 (N_4375,In_4187,In_2379);
and U4376 (N_4376,In_2642,In_1871);
xor U4377 (N_4377,In_2812,In_4269);
xnor U4378 (N_4378,In_1454,In_1684);
and U4379 (N_4379,In_3508,In_536);
or U4380 (N_4380,In_4698,In_3351);
and U4381 (N_4381,In_4209,In_3520);
or U4382 (N_4382,In_1284,In_4963);
or U4383 (N_4383,In_2710,In_2023);
or U4384 (N_4384,In_1914,In_2145);
nand U4385 (N_4385,In_712,In_4101);
xor U4386 (N_4386,In_2067,In_1088);
or U4387 (N_4387,In_2748,In_3288);
xor U4388 (N_4388,In_1683,In_1654);
xnor U4389 (N_4389,In_2873,In_2099);
xnor U4390 (N_4390,In_3280,In_1487);
and U4391 (N_4391,In_4586,In_4428);
nand U4392 (N_4392,In_1964,In_1430);
nand U4393 (N_4393,In_11,In_4921);
xnor U4394 (N_4394,In_1993,In_299);
nand U4395 (N_4395,In_3300,In_4538);
nand U4396 (N_4396,In_543,In_3411);
or U4397 (N_4397,In_2374,In_936);
or U4398 (N_4398,In_4706,In_4175);
and U4399 (N_4399,In_3665,In_1371);
or U4400 (N_4400,In_379,In_1252);
nand U4401 (N_4401,In_722,In_3291);
nand U4402 (N_4402,In_373,In_1925);
nand U4403 (N_4403,In_4699,In_4034);
nand U4404 (N_4404,In_2480,In_4300);
xor U4405 (N_4405,In_532,In_1875);
and U4406 (N_4406,In_4322,In_2738);
or U4407 (N_4407,In_1173,In_4097);
xnor U4408 (N_4408,In_1495,In_1671);
nor U4409 (N_4409,In_4796,In_3779);
nor U4410 (N_4410,In_598,In_1887);
nand U4411 (N_4411,In_2711,In_3029);
and U4412 (N_4412,In_1808,In_4416);
nor U4413 (N_4413,In_3846,In_469);
nand U4414 (N_4414,In_3053,In_566);
xor U4415 (N_4415,In_167,In_900);
or U4416 (N_4416,In_2495,In_2720);
or U4417 (N_4417,In_1262,In_638);
or U4418 (N_4418,In_2167,In_4388);
or U4419 (N_4419,In_1247,In_4768);
and U4420 (N_4420,In_3442,In_4757);
and U4421 (N_4421,In_4575,In_4251);
and U4422 (N_4422,In_4957,In_2534);
xor U4423 (N_4423,In_1039,In_3312);
and U4424 (N_4424,In_1472,In_2682);
or U4425 (N_4425,In_2117,In_3380);
and U4426 (N_4426,In_4224,In_99);
nand U4427 (N_4427,In_4148,In_4559);
or U4428 (N_4428,In_4867,In_911);
xnor U4429 (N_4429,In_4527,In_1779);
and U4430 (N_4430,In_4254,In_3380);
or U4431 (N_4431,In_2528,In_4593);
and U4432 (N_4432,In_142,In_3976);
or U4433 (N_4433,In_2770,In_1326);
nor U4434 (N_4434,In_544,In_4797);
and U4435 (N_4435,In_3475,In_2077);
xor U4436 (N_4436,In_2787,In_2775);
and U4437 (N_4437,In_4581,In_1913);
and U4438 (N_4438,In_670,In_3212);
nor U4439 (N_4439,In_3312,In_3800);
xor U4440 (N_4440,In_2592,In_4547);
or U4441 (N_4441,In_415,In_881);
xnor U4442 (N_4442,In_6,In_3304);
nor U4443 (N_4443,In_3489,In_523);
xor U4444 (N_4444,In_982,In_1648);
and U4445 (N_4445,In_13,In_4358);
nor U4446 (N_4446,In_1582,In_1341);
xnor U4447 (N_4447,In_3588,In_3789);
nand U4448 (N_4448,In_4689,In_2151);
xor U4449 (N_4449,In_4249,In_4126);
and U4450 (N_4450,In_2779,In_1412);
nor U4451 (N_4451,In_2582,In_1584);
nor U4452 (N_4452,In_4295,In_4604);
and U4453 (N_4453,In_1243,In_1726);
and U4454 (N_4454,In_477,In_3090);
nand U4455 (N_4455,In_4668,In_1681);
and U4456 (N_4456,In_2600,In_3166);
or U4457 (N_4457,In_4548,In_4631);
nand U4458 (N_4458,In_2583,In_4513);
and U4459 (N_4459,In_3974,In_2165);
nand U4460 (N_4460,In_2144,In_1371);
and U4461 (N_4461,In_1669,In_4841);
nor U4462 (N_4462,In_58,In_1677);
or U4463 (N_4463,In_4450,In_1012);
or U4464 (N_4464,In_3010,In_590);
and U4465 (N_4465,In_4683,In_3116);
and U4466 (N_4466,In_3019,In_3421);
or U4467 (N_4467,In_2913,In_3250);
or U4468 (N_4468,In_4780,In_610);
xor U4469 (N_4469,In_4832,In_406);
nand U4470 (N_4470,In_3254,In_4849);
nor U4471 (N_4471,In_4454,In_2039);
xnor U4472 (N_4472,In_185,In_3582);
nand U4473 (N_4473,In_483,In_2838);
or U4474 (N_4474,In_3236,In_1419);
and U4475 (N_4475,In_1476,In_2995);
and U4476 (N_4476,In_757,In_368);
and U4477 (N_4477,In_3172,In_3825);
nor U4478 (N_4478,In_4730,In_62);
xnor U4479 (N_4479,In_409,In_1972);
or U4480 (N_4480,In_1915,In_2913);
and U4481 (N_4481,In_4384,In_767);
xor U4482 (N_4482,In_3979,In_3005);
or U4483 (N_4483,In_741,In_2603);
xor U4484 (N_4484,In_980,In_3302);
xnor U4485 (N_4485,In_2888,In_4896);
xor U4486 (N_4486,In_1681,In_4210);
or U4487 (N_4487,In_1799,In_425);
nand U4488 (N_4488,In_780,In_4677);
nor U4489 (N_4489,In_264,In_32);
or U4490 (N_4490,In_3309,In_2819);
xor U4491 (N_4491,In_3243,In_1370);
and U4492 (N_4492,In_1053,In_3746);
nor U4493 (N_4493,In_1406,In_4910);
and U4494 (N_4494,In_866,In_2093);
xor U4495 (N_4495,In_3721,In_4809);
nand U4496 (N_4496,In_2548,In_3567);
or U4497 (N_4497,In_2917,In_1801);
nand U4498 (N_4498,In_2336,In_3895);
nor U4499 (N_4499,In_4168,In_4579);
and U4500 (N_4500,In_2144,In_4467);
nor U4501 (N_4501,In_3744,In_3423);
nor U4502 (N_4502,In_629,In_3545);
nand U4503 (N_4503,In_1931,In_1072);
or U4504 (N_4504,In_314,In_1699);
and U4505 (N_4505,In_1933,In_2858);
and U4506 (N_4506,In_4208,In_673);
nand U4507 (N_4507,In_339,In_4937);
nor U4508 (N_4508,In_3876,In_2525);
or U4509 (N_4509,In_1765,In_3142);
nor U4510 (N_4510,In_961,In_3060);
or U4511 (N_4511,In_2174,In_2731);
or U4512 (N_4512,In_9,In_2164);
or U4513 (N_4513,In_3087,In_1163);
and U4514 (N_4514,In_548,In_2358);
nor U4515 (N_4515,In_1047,In_499);
nor U4516 (N_4516,In_1560,In_3365);
nor U4517 (N_4517,In_2696,In_4490);
or U4518 (N_4518,In_2152,In_4529);
and U4519 (N_4519,In_2071,In_3195);
xnor U4520 (N_4520,In_4322,In_4421);
xnor U4521 (N_4521,In_183,In_1354);
nor U4522 (N_4522,In_3981,In_3291);
and U4523 (N_4523,In_4974,In_2138);
nand U4524 (N_4524,In_3431,In_3778);
nor U4525 (N_4525,In_1149,In_4269);
or U4526 (N_4526,In_1237,In_1755);
xnor U4527 (N_4527,In_732,In_4602);
nand U4528 (N_4528,In_2866,In_1665);
and U4529 (N_4529,In_909,In_1903);
nand U4530 (N_4530,In_760,In_2109);
or U4531 (N_4531,In_4598,In_1560);
nand U4532 (N_4532,In_374,In_676);
nand U4533 (N_4533,In_1144,In_413);
xor U4534 (N_4534,In_1080,In_4329);
or U4535 (N_4535,In_2026,In_1612);
and U4536 (N_4536,In_4072,In_2081);
nand U4537 (N_4537,In_2277,In_79);
xor U4538 (N_4538,In_2475,In_3274);
nor U4539 (N_4539,In_4023,In_1517);
nor U4540 (N_4540,In_1914,In_4447);
or U4541 (N_4541,In_2913,In_4912);
nand U4542 (N_4542,In_2668,In_3108);
nand U4543 (N_4543,In_3715,In_382);
nor U4544 (N_4544,In_449,In_1710);
nor U4545 (N_4545,In_3548,In_2228);
or U4546 (N_4546,In_399,In_207);
or U4547 (N_4547,In_49,In_703);
nor U4548 (N_4548,In_2635,In_3768);
or U4549 (N_4549,In_3749,In_3906);
and U4550 (N_4550,In_2964,In_1509);
or U4551 (N_4551,In_199,In_4575);
nor U4552 (N_4552,In_4080,In_3457);
and U4553 (N_4553,In_4424,In_1833);
nor U4554 (N_4554,In_4006,In_4095);
or U4555 (N_4555,In_1005,In_654);
or U4556 (N_4556,In_1820,In_1755);
and U4557 (N_4557,In_951,In_1372);
nor U4558 (N_4558,In_1206,In_3429);
and U4559 (N_4559,In_2097,In_1051);
xnor U4560 (N_4560,In_1278,In_684);
xor U4561 (N_4561,In_4963,In_4612);
xor U4562 (N_4562,In_2696,In_4780);
xnor U4563 (N_4563,In_441,In_4513);
nor U4564 (N_4564,In_1136,In_4595);
xor U4565 (N_4565,In_2313,In_2576);
and U4566 (N_4566,In_3166,In_2853);
nor U4567 (N_4567,In_1193,In_666);
nand U4568 (N_4568,In_3762,In_454);
or U4569 (N_4569,In_4211,In_3570);
xor U4570 (N_4570,In_2363,In_4090);
nor U4571 (N_4571,In_3292,In_4451);
nor U4572 (N_4572,In_2947,In_2320);
nor U4573 (N_4573,In_4128,In_3955);
nand U4574 (N_4574,In_1437,In_101);
and U4575 (N_4575,In_2335,In_3090);
nor U4576 (N_4576,In_2919,In_3612);
xnor U4577 (N_4577,In_4220,In_2424);
and U4578 (N_4578,In_3633,In_2532);
or U4579 (N_4579,In_4344,In_3840);
and U4580 (N_4580,In_1541,In_3684);
nand U4581 (N_4581,In_863,In_4985);
and U4582 (N_4582,In_4712,In_1487);
xor U4583 (N_4583,In_2963,In_382);
nand U4584 (N_4584,In_1986,In_1482);
and U4585 (N_4585,In_2616,In_3790);
nand U4586 (N_4586,In_2603,In_4990);
nor U4587 (N_4587,In_3577,In_4734);
and U4588 (N_4588,In_4076,In_1585);
nor U4589 (N_4589,In_1192,In_3282);
xor U4590 (N_4590,In_1859,In_3421);
xor U4591 (N_4591,In_3582,In_4973);
nand U4592 (N_4592,In_2151,In_3732);
xnor U4593 (N_4593,In_1889,In_2061);
nand U4594 (N_4594,In_3267,In_182);
xnor U4595 (N_4595,In_1125,In_4927);
or U4596 (N_4596,In_4810,In_1324);
nand U4597 (N_4597,In_625,In_3569);
nor U4598 (N_4598,In_3328,In_4089);
or U4599 (N_4599,In_3127,In_4547);
nor U4600 (N_4600,In_2671,In_3940);
nor U4601 (N_4601,In_4315,In_2222);
nor U4602 (N_4602,In_2322,In_1851);
xnor U4603 (N_4603,In_2407,In_4392);
or U4604 (N_4604,In_4700,In_3635);
nor U4605 (N_4605,In_1001,In_1978);
nand U4606 (N_4606,In_4907,In_584);
and U4607 (N_4607,In_1578,In_942);
nor U4608 (N_4608,In_58,In_2719);
nand U4609 (N_4609,In_842,In_3133);
nand U4610 (N_4610,In_3696,In_4294);
or U4611 (N_4611,In_965,In_3687);
or U4612 (N_4612,In_2763,In_1688);
nor U4613 (N_4613,In_2849,In_540);
nand U4614 (N_4614,In_1216,In_942);
nor U4615 (N_4615,In_4105,In_2531);
nand U4616 (N_4616,In_1278,In_4819);
nor U4617 (N_4617,In_3165,In_1000);
nor U4618 (N_4618,In_1830,In_1701);
and U4619 (N_4619,In_3289,In_1033);
nor U4620 (N_4620,In_1646,In_1045);
nand U4621 (N_4621,In_4049,In_3677);
xnor U4622 (N_4622,In_3955,In_2137);
and U4623 (N_4623,In_185,In_3084);
nand U4624 (N_4624,In_2468,In_3335);
nor U4625 (N_4625,In_3358,In_3231);
nand U4626 (N_4626,In_1614,In_1438);
nand U4627 (N_4627,In_4664,In_435);
nor U4628 (N_4628,In_1863,In_2182);
nand U4629 (N_4629,In_3441,In_906);
and U4630 (N_4630,In_124,In_4664);
xnor U4631 (N_4631,In_4120,In_2190);
and U4632 (N_4632,In_3694,In_52);
nor U4633 (N_4633,In_4675,In_1243);
nand U4634 (N_4634,In_1369,In_1256);
and U4635 (N_4635,In_4010,In_2309);
nand U4636 (N_4636,In_3896,In_2998);
nor U4637 (N_4637,In_1708,In_2040);
or U4638 (N_4638,In_1516,In_817);
xor U4639 (N_4639,In_574,In_1178);
nor U4640 (N_4640,In_2905,In_2761);
xor U4641 (N_4641,In_2786,In_1937);
xnor U4642 (N_4642,In_656,In_1457);
xor U4643 (N_4643,In_4410,In_244);
nor U4644 (N_4644,In_3662,In_2027);
xor U4645 (N_4645,In_3193,In_4038);
xor U4646 (N_4646,In_1048,In_2880);
xnor U4647 (N_4647,In_2323,In_4689);
xnor U4648 (N_4648,In_4419,In_3816);
nand U4649 (N_4649,In_3336,In_342);
or U4650 (N_4650,In_4801,In_304);
nand U4651 (N_4651,In_1197,In_240);
and U4652 (N_4652,In_1629,In_3159);
and U4653 (N_4653,In_713,In_2793);
xor U4654 (N_4654,In_1838,In_10);
or U4655 (N_4655,In_4845,In_3734);
or U4656 (N_4656,In_1549,In_4054);
nand U4657 (N_4657,In_2613,In_4163);
and U4658 (N_4658,In_56,In_1340);
and U4659 (N_4659,In_4195,In_2342);
nor U4660 (N_4660,In_3968,In_4942);
nor U4661 (N_4661,In_2867,In_4900);
and U4662 (N_4662,In_2571,In_3801);
and U4663 (N_4663,In_304,In_658);
nand U4664 (N_4664,In_2043,In_3548);
nor U4665 (N_4665,In_3718,In_1986);
and U4666 (N_4666,In_3900,In_1751);
and U4667 (N_4667,In_164,In_3997);
nor U4668 (N_4668,In_4167,In_297);
nor U4669 (N_4669,In_4406,In_3336);
nor U4670 (N_4670,In_3350,In_1338);
nand U4671 (N_4671,In_499,In_4862);
nand U4672 (N_4672,In_2824,In_888);
nor U4673 (N_4673,In_4091,In_302);
xor U4674 (N_4674,In_669,In_2561);
xor U4675 (N_4675,In_1983,In_4872);
and U4676 (N_4676,In_987,In_3575);
nand U4677 (N_4677,In_353,In_1468);
and U4678 (N_4678,In_4497,In_2695);
nor U4679 (N_4679,In_1613,In_2632);
or U4680 (N_4680,In_3969,In_4526);
or U4681 (N_4681,In_164,In_3644);
and U4682 (N_4682,In_350,In_1529);
and U4683 (N_4683,In_942,In_2484);
or U4684 (N_4684,In_890,In_3160);
xnor U4685 (N_4685,In_349,In_2554);
xnor U4686 (N_4686,In_3681,In_4110);
xnor U4687 (N_4687,In_812,In_2266);
nor U4688 (N_4688,In_4280,In_893);
and U4689 (N_4689,In_782,In_4292);
nand U4690 (N_4690,In_2949,In_4534);
xnor U4691 (N_4691,In_3641,In_4439);
or U4692 (N_4692,In_4910,In_4984);
or U4693 (N_4693,In_390,In_3219);
and U4694 (N_4694,In_1983,In_3070);
xnor U4695 (N_4695,In_2213,In_119);
and U4696 (N_4696,In_880,In_2794);
nand U4697 (N_4697,In_333,In_4862);
and U4698 (N_4698,In_662,In_230);
and U4699 (N_4699,In_4080,In_1849);
nor U4700 (N_4700,In_1704,In_4870);
or U4701 (N_4701,In_4154,In_2372);
or U4702 (N_4702,In_4550,In_2108);
and U4703 (N_4703,In_1996,In_772);
xnor U4704 (N_4704,In_1106,In_2101);
nand U4705 (N_4705,In_1875,In_2603);
xnor U4706 (N_4706,In_1672,In_883);
xor U4707 (N_4707,In_1706,In_3891);
nor U4708 (N_4708,In_3703,In_2431);
xor U4709 (N_4709,In_3676,In_2116);
xor U4710 (N_4710,In_4914,In_1586);
xor U4711 (N_4711,In_4599,In_3889);
and U4712 (N_4712,In_4455,In_3142);
or U4713 (N_4713,In_1091,In_341);
nand U4714 (N_4714,In_4059,In_3931);
and U4715 (N_4715,In_4725,In_508);
and U4716 (N_4716,In_4009,In_1076);
nand U4717 (N_4717,In_1092,In_2806);
nor U4718 (N_4718,In_3926,In_4821);
and U4719 (N_4719,In_4653,In_2924);
nor U4720 (N_4720,In_479,In_4318);
xor U4721 (N_4721,In_478,In_1480);
xnor U4722 (N_4722,In_4188,In_4065);
and U4723 (N_4723,In_2459,In_4146);
or U4724 (N_4724,In_4012,In_3528);
nand U4725 (N_4725,In_4539,In_1428);
nor U4726 (N_4726,In_3206,In_945);
nor U4727 (N_4727,In_3740,In_2241);
nand U4728 (N_4728,In_2799,In_3704);
xnor U4729 (N_4729,In_1700,In_1102);
or U4730 (N_4730,In_3483,In_1011);
xor U4731 (N_4731,In_2612,In_4988);
nand U4732 (N_4732,In_805,In_3161);
nor U4733 (N_4733,In_1013,In_3834);
nand U4734 (N_4734,In_1729,In_4622);
or U4735 (N_4735,In_4828,In_3416);
and U4736 (N_4736,In_4901,In_977);
and U4737 (N_4737,In_2479,In_2498);
nand U4738 (N_4738,In_4777,In_2823);
or U4739 (N_4739,In_140,In_213);
nor U4740 (N_4740,In_3082,In_4764);
xor U4741 (N_4741,In_1481,In_2594);
and U4742 (N_4742,In_4144,In_2316);
nor U4743 (N_4743,In_2194,In_274);
or U4744 (N_4744,In_4170,In_510);
and U4745 (N_4745,In_1198,In_3697);
nor U4746 (N_4746,In_2551,In_4625);
and U4747 (N_4747,In_4378,In_3799);
xnor U4748 (N_4748,In_4843,In_2803);
nor U4749 (N_4749,In_4004,In_1883);
and U4750 (N_4750,In_2000,In_1091);
and U4751 (N_4751,In_2670,In_3239);
nor U4752 (N_4752,In_3815,In_4106);
or U4753 (N_4753,In_568,In_1352);
or U4754 (N_4754,In_480,In_4229);
xnor U4755 (N_4755,In_2459,In_1904);
xor U4756 (N_4756,In_161,In_3090);
nor U4757 (N_4757,In_3493,In_1269);
xor U4758 (N_4758,In_4817,In_3242);
or U4759 (N_4759,In_3497,In_2718);
xnor U4760 (N_4760,In_2542,In_4217);
nor U4761 (N_4761,In_3475,In_2309);
nor U4762 (N_4762,In_1084,In_2272);
or U4763 (N_4763,In_3708,In_2331);
or U4764 (N_4764,In_918,In_3004);
and U4765 (N_4765,In_3192,In_1068);
nor U4766 (N_4766,In_524,In_181);
and U4767 (N_4767,In_4021,In_1433);
xor U4768 (N_4768,In_1273,In_4597);
and U4769 (N_4769,In_3055,In_1425);
xnor U4770 (N_4770,In_1245,In_4593);
and U4771 (N_4771,In_746,In_1167);
and U4772 (N_4772,In_2974,In_3783);
nor U4773 (N_4773,In_4022,In_2724);
xor U4774 (N_4774,In_1508,In_4384);
nor U4775 (N_4775,In_718,In_1682);
and U4776 (N_4776,In_2499,In_990);
nand U4777 (N_4777,In_1226,In_574);
xnor U4778 (N_4778,In_1072,In_316);
xnor U4779 (N_4779,In_2556,In_257);
nand U4780 (N_4780,In_2664,In_1764);
nor U4781 (N_4781,In_4331,In_1908);
and U4782 (N_4782,In_741,In_4086);
or U4783 (N_4783,In_1765,In_302);
nor U4784 (N_4784,In_4511,In_1820);
or U4785 (N_4785,In_272,In_2198);
nand U4786 (N_4786,In_3865,In_2246);
nor U4787 (N_4787,In_2169,In_2516);
nand U4788 (N_4788,In_2743,In_2245);
nor U4789 (N_4789,In_1537,In_3027);
xor U4790 (N_4790,In_2810,In_2958);
nor U4791 (N_4791,In_1783,In_1660);
and U4792 (N_4792,In_4123,In_617);
xor U4793 (N_4793,In_835,In_931);
xnor U4794 (N_4794,In_1559,In_2920);
and U4795 (N_4795,In_4621,In_3429);
and U4796 (N_4796,In_1565,In_2246);
nor U4797 (N_4797,In_3798,In_2505);
nor U4798 (N_4798,In_2020,In_3267);
xnor U4799 (N_4799,In_3877,In_4845);
nand U4800 (N_4800,In_2947,In_4914);
or U4801 (N_4801,In_20,In_4991);
xnor U4802 (N_4802,In_4501,In_564);
or U4803 (N_4803,In_2843,In_1145);
nand U4804 (N_4804,In_4948,In_1718);
xnor U4805 (N_4805,In_4014,In_3257);
or U4806 (N_4806,In_4377,In_2374);
nand U4807 (N_4807,In_3048,In_735);
xnor U4808 (N_4808,In_4799,In_3480);
or U4809 (N_4809,In_46,In_3832);
and U4810 (N_4810,In_3480,In_3894);
and U4811 (N_4811,In_963,In_918);
nor U4812 (N_4812,In_4877,In_2713);
nor U4813 (N_4813,In_3021,In_1043);
or U4814 (N_4814,In_1967,In_3968);
and U4815 (N_4815,In_4937,In_1100);
or U4816 (N_4816,In_3857,In_1401);
nor U4817 (N_4817,In_1241,In_4302);
or U4818 (N_4818,In_3886,In_2883);
nor U4819 (N_4819,In_2839,In_2731);
nand U4820 (N_4820,In_3838,In_2096);
nand U4821 (N_4821,In_3788,In_4535);
nand U4822 (N_4822,In_4705,In_2681);
or U4823 (N_4823,In_3867,In_3011);
xnor U4824 (N_4824,In_2384,In_666);
xor U4825 (N_4825,In_4806,In_385);
xnor U4826 (N_4826,In_1766,In_32);
and U4827 (N_4827,In_4079,In_2689);
and U4828 (N_4828,In_2411,In_1090);
or U4829 (N_4829,In_2290,In_1766);
nor U4830 (N_4830,In_2655,In_1212);
xor U4831 (N_4831,In_4816,In_4251);
or U4832 (N_4832,In_3364,In_644);
nand U4833 (N_4833,In_1081,In_4954);
nor U4834 (N_4834,In_3651,In_2642);
and U4835 (N_4835,In_4169,In_2026);
or U4836 (N_4836,In_3530,In_1394);
xor U4837 (N_4837,In_2438,In_3153);
or U4838 (N_4838,In_1800,In_3228);
nand U4839 (N_4839,In_3159,In_3897);
nand U4840 (N_4840,In_1121,In_1747);
xnor U4841 (N_4841,In_2444,In_439);
and U4842 (N_4842,In_3945,In_96);
nand U4843 (N_4843,In_1841,In_4691);
nor U4844 (N_4844,In_1477,In_525);
xnor U4845 (N_4845,In_1450,In_147);
xnor U4846 (N_4846,In_3673,In_4910);
xnor U4847 (N_4847,In_4354,In_2746);
nand U4848 (N_4848,In_3414,In_1067);
and U4849 (N_4849,In_1322,In_2022);
and U4850 (N_4850,In_3570,In_1010);
and U4851 (N_4851,In_4912,In_54);
nand U4852 (N_4852,In_4199,In_2607);
nand U4853 (N_4853,In_3450,In_3093);
nor U4854 (N_4854,In_4283,In_56);
xnor U4855 (N_4855,In_649,In_4265);
nor U4856 (N_4856,In_3662,In_3672);
nor U4857 (N_4857,In_1968,In_1314);
nand U4858 (N_4858,In_3091,In_2140);
xor U4859 (N_4859,In_4842,In_4915);
and U4860 (N_4860,In_4189,In_1096);
nor U4861 (N_4861,In_4798,In_4382);
nor U4862 (N_4862,In_2945,In_2134);
xnor U4863 (N_4863,In_3825,In_630);
nor U4864 (N_4864,In_4261,In_4159);
nor U4865 (N_4865,In_4014,In_3280);
or U4866 (N_4866,In_336,In_2984);
and U4867 (N_4867,In_37,In_2881);
and U4868 (N_4868,In_0,In_1485);
xnor U4869 (N_4869,In_4195,In_4226);
nand U4870 (N_4870,In_3851,In_4330);
nor U4871 (N_4871,In_2626,In_204);
and U4872 (N_4872,In_1176,In_3220);
and U4873 (N_4873,In_4346,In_2677);
nor U4874 (N_4874,In_2967,In_2974);
and U4875 (N_4875,In_1635,In_4607);
xor U4876 (N_4876,In_3242,In_4633);
nand U4877 (N_4877,In_1662,In_1089);
xor U4878 (N_4878,In_1847,In_4731);
or U4879 (N_4879,In_2699,In_1096);
nand U4880 (N_4880,In_176,In_162);
or U4881 (N_4881,In_1060,In_1306);
nor U4882 (N_4882,In_436,In_4247);
nor U4883 (N_4883,In_1268,In_4472);
nand U4884 (N_4884,In_1612,In_4280);
and U4885 (N_4885,In_3743,In_1956);
nor U4886 (N_4886,In_2254,In_4587);
nand U4887 (N_4887,In_4164,In_3968);
xor U4888 (N_4888,In_2292,In_4894);
and U4889 (N_4889,In_1190,In_2223);
and U4890 (N_4890,In_3271,In_1022);
nor U4891 (N_4891,In_2924,In_1178);
nor U4892 (N_4892,In_2147,In_2440);
xnor U4893 (N_4893,In_2469,In_194);
nor U4894 (N_4894,In_2257,In_2956);
or U4895 (N_4895,In_2791,In_841);
and U4896 (N_4896,In_4975,In_3433);
or U4897 (N_4897,In_1227,In_792);
nand U4898 (N_4898,In_866,In_3215);
nand U4899 (N_4899,In_2330,In_4359);
or U4900 (N_4900,In_4910,In_2719);
xnor U4901 (N_4901,In_1299,In_2450);
and U4902 (N_4902,In_1117,In_4379);
nor U4903 (N_4903,In_4578,In_2714);
xor U4904 (N_4904,In_2052,In_4823);
nand U4905 (N_4905,In_2482,In_482);
nand U4906 (N_4906,In_3649,In_3028);
or U4907 (N_4907,In_801,In_2495);
or U4908 (N_4908,In_3034,In_1827);
and U4909 (N_4909,In_2557,In_2710);
xnor U4910 (N_4910,In_1817,In_2055);
nor U4911 (N_4911,In_4895,In_2681);
xnor U4912 (N_4912,In_1600,In_69);
nor U4913 (N_4913,In_4978,In_1224);
nand U4914 (N_4914,In_2966,In_1836);
xnor U4915 (N_4915,In_2808,In_4438);
nand U4916 (N_4916,In_4112,In_2988);
and U4917 (N_4917,In_3598,In_4516);
nor U4918 (N_4918,In_3364,In_2865);
and U4919 (N_4919,In_511,In_1911);
and U4920 (N_4920,In_1744,In_2185);
and U4921 (N_4921,In_3810,In_585);
and U4922 (N_4922,In_3687,In_386);
xnor U4923 (N_4923,In_2649,In_2550);
and U4924 (N_4924,In_377,In_3751);
nand U4925 (N_4925,In_2630,In_4261);
and U4926 (N_4926,In_1680,In_4539);
xnor U4927 (N_4927,In_2144,In_2941);
xor U4928 (N_4928,In_387,In_4109);
nor U4929 (N_4929,In_1494,In_4024);
nor U4930 (N_4930,In_4222,In_3231);
xor U4931 (N_4931,In_2773,In_1497);
nor U4932 (N_4932,In_1831,In_3446);
xnor U4933 (N_4933,In_894,In_1394);
nand U4934 (N_4934,In_535,In_2492);
or U4935 (N_4935,In_4986,In_3885);
nor U4936 (N_4936,In_3496,In_2598);
nor U4937 (N_4937,In_2404,In_4141);
nand U4938 (N_4938,In_2892,In_2602);
nand U4939 (N_4939,In_2993,In_163);
xor U4940 (N_4940,In_2686,In_616);
nor U4941 (N_4941,In_2146,In_3290);
xnor U4942 (N_4942,In_1014,In_1771);
and U4943 (N_4943,In_3566,In_255);
xor U4944 (N_4944,In_671,In_2188);
xor U4945 (N_4945,In_204,In_2600);
or U4946 (N_4946,In_3279,In_1310);
nor U4947 (N_4947,In_1643,In_1359);
and U4948 (N_4948,In_1648,In_4323);
xor U4949 (N_4949,In_675,In_3688);
and U4950 (N_4950,In_2781,In_4643);
and U4951 (N_4951,In_451,In_1384);
or U4952 (N_4952,In_4785,In_2516);
nor U4953 (N_4953,In_4656,In_443);
or U4954 (N_4954,In_4291,In_2622);
nand U4955 (N_4955,In_4723,In_3335);
nor U4956 (N_4956,In_2004,In_2280);
and U4957 (N_4957,In_4775,In_4015);
or U4958 (N_4958,In_837,In_4424);
nor U4959 (N_4959,In_1250,In_1342);
xor U4960 (N_4960,In_279,In_2125);
xnor U4961 (N_4961,In_609,In_3387);
nand U4962 (N_4962,In_1864,In_3433);
or U4963 (N_4963,In_2306,In_2495);
xnor U4964 (N_4964,In_350,In_3668);
or U4965 (N_4965,In_1847,In_4183);
and U4966 (N_4966,In_1229,In_3950);
and U4967 (N_4967,In_3686,In_4376);
xor U4968 (N_4968,In_2763,In_1058);
nor U4969 (N_4969,In_1889,In_3812);
nor U4970 (N_4970,In_2998,In_294);
nand U4971 (N_4971,In_3702,In_1352);
and U4972 (N_4972,In_1034,In_4374);
xnor U4973 (N_4973,In_2060,In_2453);
nand U4974 (N_4974,In_3952,In_4552);
nor U4975 (N_4975,In_4754,In_4470);
xor U4976 (N_4976,In_3007,In_3077);
or U4977 (N_4977,In_3466,In_4978);
nand U4978 (N_4978,In_4561,In_2235);
and U4979 (N_4979,In_1715,In_4323);
xnor U4980 (N_4980,In_4550,In_34);
xor U4981 (N_4981,In_1771,In_3406);
and U4982 (N_4982,In_1548,In_3458);
nand U4983 (N_4983,In_3619,In_3394);
nor U4984 (N_4984,In_3032,In_53);
nand U4985 (N_4985,In_2064,In_287);
nand U4986 (N_4986,In_376,In_2741);
xnor U4987 (N_4987,In_3825,In_1467);
or U4988 (N_4988,In_113,In_4816);
xnor U4989 (N_4989,In_4038,In_3342);
nand U4990 (N_4990,In_3571,In_4113);
nor U4991 (N_4991,In_2317,In_1665);
nand U4992 (N_4992,In_2715,In_2716);
and U4993 (N_4993,In_2373,In_606);
and U4994 (N_4994,In_623,In_1344);
and U4995 (N_4995,In_4531,In_391);
nor U4996 (N_4996,In_3720,In_1041);
nor U4997 (N_4997,In_4919,In_4660);
and U4998 (N_4998,In_462,In_2345);
nand U4999 (N_4999,In_1159,In_3006);
or U5000 (N_5000,N_1844,N_2401);
xor U5001 (N_5001,N_886,N_4097);
nor U5002 (N_5002,N_3189,N_4324);
nand U5003 (N_5003,N_4904,N_16);
nand U5004 (N_5004,N_1376,N_4575);
nor U5005 (N_5005,N_3168,N_4426);
or U5006 (N_5006,N_1249,N_1384);
nand U5007 (N_5007,N_4429,N_4353);
nand U5008 (N_5008,N_2890,N_4184);
nand U5009 (N_5009,N_3524,N_1532);
nand U5010 (N_5010,N_3288,N_619);
xor U5011 (N_5011,N_898,N_1917);
nor U5012 (N_5012,N_2484,N_125);
xor U5013 (N_5013,N_2104,N_1943);
nor U5014 (N_5014,N_2871,N_3674);
and U5015 (N_5015,N_1057,N_3160);
and U5016 (N_5016,N_2861,N_3270);
and U5017 (N_5017,N_4349,N_3985);
and U5018 (N_5018,N_881,N_2606);
nand U5019 (N_5019,N_2506,N_4294);
and U5020 (N_5020,N_2553,N_2777);
and U5021 (N_5021,N_1297,N_4967);
or U5022 (N_5022,N_3476,N_299);
nor U5023 (N_5023,N_2279,N_3412);
nand U5024 (N_5024,N_767,N_4508);
nor U5025 (N_5025,N_4139,N_1149);
nand U5026 (N_5026,N_4132,N_867);
nor U5027 (N_5027,N_2978,N_2296);
and U5028 (N_5028,N_3907,N_995);
and U5029 (N_5029,N_906,N_567);
nor U5030 (N_5030,N_4057,N_3503);
nor U5031 (N_5031,N_1066,N_817);
nand U5032 (N_5032,N_1264,N_4092);
nand U5033 (N_5033,N_3194,N_1617);
and U5034 (N_5034,N_3931,N_3977);
or U5035 (N_5035,N_2788,N_3402);
xnor U5036 (N_5036,N_1675,N_4811);
xor U5037 (N_5037,N_690,N_3131);
nor U5038 (N_5038,N_775,N_3560);
or U5039 (N_5039,N_2999,N_4679);
nand U5040 (N_5040,N_3898,N_2151);
nand U5041 (N_5041,N_1131,N_1133);
or U5042 (N_5042,N_1932,N_195);
or U5043 (N_5043,N_2997,N_4912);
nor U5044 (N_5044,N_3355,N_2627);
xnor U5045 (N_5045,N_2274,N_4832);
nand U5046 (N_5046,N_1261,N_4185);
nand U5047 (N_5047,N_1010,N_89);
or U5048 (N_5048,N_2519,N_4628);
nand U5049 (N_5049,N_2432,N_4638);
nand U5050 (N_5050,N_1766,N_3403);
nor U5051 (N_5051,N_965,N_412);
xor U5052 (N_5052,N_3036,N_3046);
nand U5053 (N_5053,N_4277,N_3462);
xor U5054 (N_5054,N_3593,N_1341);
and U5055 (N_5055,N_897,N_929);
xor U5056 (N_5056,N_1649,N_116);
xnor U5057 (N_5057,N_2510,N_2042);
xnor U5058 (N_5058,N_3387,N_1797);
nor U5059 (N_5059,N_1948,N_2775);
and U5060 (N_5060,N_4228,N_4712);
nor U5061 (N_5061,N_3429,N_3438);
xnor U5062 (N_5062,N_2517,N_1478);
or U5063 (N_5063,N_4568,N_1007);
nor U5064 (N_5064,N_2940,N_978);
nor U5065 (N_5065,N_1112,N_4913);
nor U5066 (N_5066,N_1070,N_1317);
or U5067 (N_5067,N_2284,N_3865);
xnor U5068 (N_5068,N_3991,N_3130);
nand U5069 (N_5069,N_1431,N_3464);
nand U5070 (N_5070,N_2560,N_207);
nor U5071 (N_5071,N_1798,N_2847);
nand U5072 (N_5072,N_3006,N_2710);
and U5073 (N_5073,N_560,N_4141);
and U5074 (N_5074,N_2811,N_4510);
or U5075 (N_5075,N_1470,N_2898);
and U5076 (N_5076,N_592,N_1678);
and U5077 (N_5077,N_4987,N_1385);
or U5078 (N_5078,N_4741,N_1395);
and U5079 (N_5079,N_803,N_2239);
or U5080 (N_5080,N_4088,N_551);
xor U5081 (N_5081,N_3920,N_2782);
or U5082 (N_5082,N_4234,N_1138);
or U5083 (N_5083,N_1433,N_3125);
or U5084 (N_5084,N_3468,N_1580);
and U5085 (N_5085,N_4778,N_3950);
xnor U5086 (N_5086,N_3732,N_1342);
xnor U5087 (N_5087,N_2518,N_3143);
nor U5088 (N_5088,N_4048,N_2543);
xor U5089 (N_5089,N_1450,N_4491);
nand U5090 (N_5090,N_1747,N_1656);
nand U5091 (N_5091,N_1604,N_4166);
or U5092 (N_5092,N_2479,N_110);
nand U5093 (N_5093,N_3149,N_4817);
xor U5094 (N_5094,N_387,N_1979);
or U5095 (N_5095,N_3943,N_2497);
or U5096 (N_5096,N_1897,N_733);
and U5097 (N_5097,N_1463,N_1964);
nor U5098 (N_5098,N_3650,N_2013);
nand U5099 (N_5099,N_877,N_1880);
nand U5100 (N_5100,N_4337,N_4686);
nor U5101 (N_5101,N_3071,N_3894);
nand U5102 (N_5102,N_4915,N_918);
nand U5103 (N_5103,N_4026,N_2282);
and U5104 (N_5104,N_1816,N_430);
nor U5105 (N_5105,N_4067,N_3242);
nand U5106 (N_5106,N_3782,N_3836);
nand U5107 (N_5107,N_4954,N_4417);
and U5108 (N_5108,N_837,N_1988);
nand U5109 (N_5109,N_3932,N_3981);
and U5110 (N_5110,N_3871,N_3909);
and U5111 (N_5111,N_4539,N_2546);
nor U5112 (N_5112,N_4898,N_2623);
or U5113 (N_5113,N_4320,N_3652);
and U5114 (N_5114,N_4398,N_252);
xor U5115 (N_5115,N_1866,N_2188);
nor U5116 (N_5116,N_4620,N_153);
and U5117 (N_5117,N_4259,N_2758);
nor U5118 (N_5118,N_4746,N_3622);
and U5119 (N_5119,N_4480,N_1005);
xor U5120 (N_5120,N_4461,N_1037);
and U5121 (N_5121,N_925,N_2616);
xor U5122 (N_5122,N_92,N_1120);
nor U5123 (N_5123,N_413,N_1971);
nand U5124 (N_5124,N_1743,N_4482);
nor U5125 (N_5125,N_3775,N_732);
nor U5126 (N_5126,N_756,N_1740);
and U5127 (N_5127,N_4548,N_3364);
nor U5128 (N_5128,N_3849,N_4938);
nand U5129 (N_5129,N_708,N_392);
nor U5130 (N_5130,N_246,N_2807);
xnor U5131 (N_5131,N_1288,N_2554);
nor U5132 (N_5132,N_4814,N_3328);
and U5133 (N_5133,N_2026,N_631);
nor U5134 (N_5134,N_1344,N_3214);
and U5135 (N_5135,N_4069,N_4609);
or U5136 (N_5136,N_2786,N_4086);
and U5137 (N_5137,N_399,N_4897);
nor U5138 (N_5138,N_3266,N_1464);
nand U5139 (N_5139,N_1614,N_3773);
xnor U5140 (N_5140,N_3696,N_4050);
and U5141 (N_5141,N_1224,N_3064);
nand U5142 (N_5142,N_2095,N_1712);
or U5143 (N_5143,N_3972,N_1094);
nand U5144 (N_5144,N_4546,N_3724);
nand U5145 (N_5145,N_3376,N_2304);
or U5146 (N_5146,N_2671,N_4029);
and U5147 (N_5147,N_638,N_2242);
xnor U5148 (N_5148,N_4870,N_2684);
xor U5149 (N_5149,N_4891,N_992);
or U5150 (N_5150,N_300,N_4589);
xor U5151 (N_5151,N_4151,N_4160);
nand U5152 (N_5152,N_753,N_4616);
nand U5153 (N_5153,N_4601,N_4567);
nor U5154 (N_5154,N_3655,N_1926);
nor U5155 (N_5155,N_586,N_4505);
nand U5156 (N_5156,N_3134,N_313);
nand U5157 (N_5157,N_2755,N_564);
or U5158 (N_5158,N_1025,N_3016);
and U5159 (N_5159,N_913,N_1311);
nor U5160 (N_5160,N_4696,N_2590);
or U5161 (N_5161,N_4543,N_4405);
nand U5162 (N_5162,N_3716,N_131);
or U5163 (N_5163,N_2603,N_2727);
and U5164 (N_5164,N_1974,N_839);
or U5165 (N_5165,N_1505,N_2969);
and U5166 (N_5166,N_2383,N_1683);
nand U5167 (N_5167,N_1846,N_4867);
and U5168 (N_5168,N_4326,N_3368);
nand U5169 (N_5169,N_378,N_3679);
nor U5170 (N_5170,N_1837,N_4407);
or U5171 (N_5171,N_679,N_3868);
nor U5172 (N_5172,N_893,N_1673);
and U5173 (N_5173,N_821,N_2155);
xor U5174 (N_5174,N_2916,N_4200);
nor U5175 (N_5175,N_2478,N_4641);
and U5176 (N_5176,N_80,N_294);
nand U5177 (N_5177,N_3828,N_2542);
or U5178 (N_5178,N_3798,N_1719);
xnor U5179 (N_5179,N_868,N_1919);
nand U5180 (N_5180,N_2675,N_3037);
or U5181 (N_5181,N_1391,N_962);
xnor U5182 (N_5182,N_2670,N_3997);
nand U5183 (N_5183,N_1186,N_3161);
xnor U5184 (N_5184,N_4507,N_539);
nor U5185 (N_5185,N_3183,N_4794);
xor U5186 (N_5186,N_1128,N_4582);
nor U5187 (N_5187,N_394,N_627);
xnor U5188 (N_5188,N_3459,N_3731);
and U5189 (N_5189,N_956,N_84);
nand U5190 (N_5190,N_1011,N_1817);
nor U5191 (N_5191,N_478,N_4885);
and U5192 (N_5192,N_1290,N_2696);
or U5193 (N_5193,N_4564,N_2245);
and U5194 (N_5194,N_2505,N_444);
nor U5195 (N_5195,N_2077,N_4454);
or U5196 (N_5196,N_3658,N_341);
xnor U5197 (N_5197,N_168,N_4772);
nor U5198 (N_5198,N_4734,N_1893);
and U5199 (N_5199,N_2408,N_2162);
nand U5200 (N_5200,N_4905,N_4573);
or U5201 (N_5201,N_4312,N_1830);
or U5202 (N_5202,N_3174,N_4512);
nand U5203 (N_5203,N_2996,N_2536);
xor U5204 (N_5204,N_2885,N_4835);
nand U5205 (N_5205,N_3386,N_454);
nor U5206 (N_5206,N_1954,N_3435);
nor U5207 (N_5207,N_1033,N_2264);
and U5208 (N_5208,N_3852,N_4792);
xnor U5209 (N_5209,N_1246,N_3743);
or U5210 (N_5210,N_2318,N_432);
or U5211 (N_5211,N_1884,N_723);
and U5212 (N_5212,N_56,N_1853);
or U5213 (N_5213,N_340,N_880);
and U5214 (N_5214,N_1422,N_537);
or U5215 (N_5215,N_44,N_2713);
xor U5216 (N_5216,N_4753,N_1430);
xor U5217 (N_5217,N_526,N_3757);
or U5218 (N_5218,N_1393,N_1600);
and U5219 (N_5219,N_4947,N_4183);
nand U5220 (N_5220,N_39,N_973);
or U5221 (N_5221,N_4053,N_3610);
and U5222 (N_5222,N_1471,N_828);
xor U5223 (N_5223,N_1027,N_348);
nor U5224 (N_5224,N_3225,N_4571);
nor U5225 (N_5225,N_2976,N_438);
or U5226 (N_5226,N_2718,N_4066);
and U5227 (N_5227,N_2760,N_1935);
or U5228 (N_5228,N_4771,N_144);
or U5229 (N_5229,N_1708,N_4919);
xnor U5230 (N_5230,N_4708,N_2915);
and U5231 (N_5231,N_2843,N_327);
nand U5232 (N_5232,N_1557,N_2138);
xnor U5233 (N_5233,N_3564,N_494);
and U5234 (N_5234,N_2654,N_4873);
or U5235 (N_5235,N_1881,N_4605);
xor U5236 (N_5236,N_416,N_1204);
nor U5237 (N_5237,N_146,N_648);
nand U5238 (N_5238,N_1689,N_3017);
and U5239 (N_5239,N_4075,N_3025);
nor U5240 (N_5240,N_3608,N_2102);
xor U5241 (N_5241,N_2991,N_570);
nor U5242 (N_5242,N_4118,N_4127);
nand U5243 (N_5243,N_3007,N_3015);
and U5244 (N_5244,N_1568,N_725);
and U5245 (N_5245,N_4966,N_226);
or U5246 (N_5246,N_3955,N_4348);
or U5247 (N_5247,N_2125,N_3841);
nand U5248 (N_5248,N_1793,N_1534);
and U5249 (N_5249,N_1828,N_3499);
nand U5250 (N_5250,N_3291,N_2080);
nor U5251 (N_5251,N_576,N_3123);
or U5252 (N_5252,N_2043,N_2116);
or U5253 (N_5253,N_4789,N_4193);
or U5254 (N_5254,N_4338,N_281);
nor U5255 (N_5255,N_3649,N_1259);
and U5256 (N_5256,N_3013,N_4111);
or U5257 (N_5257,N_1542,N_2678);
and U5258 (N_5258,N_4803,N_2164);
nand U5259 (N_5259,N_3888,N_2000);
xnor U5260 (N_5260,N_3646,N_4718);
or U5261 (N_5261,N_4928,N_1918);
nor U5262 (N_5262,N_2656,N_1783);
nand U5263 (N_5263,N_4117,N_3752);
or U5264 (N_5264,N_2967,N_3745);
nor U5265 (N_5265,N_3688,N_3913);
or U5266 (N_5266,N_2930,N_295);
xor U5267 (N_5267,N_3942,N_1840);
xnor U5268 (N_5268,N_243,N_3445);
xnor U5269 (N_5269,N_583,N_4540);
nor U5270 (N_5270,N_1192,N_626);
nor U5271 (N_5271,N_451,N_3479);
nor U5272 (N_5272,N_991,N_417);
nand U5273 (N_5273,N_4666,N_4239);
and U5274 (N_5274,N_4557,N_71);
or U5275 (N_5275,N_393,N_3185);
and U5276 (N_5276,N_590,N_4464);
and U5277 (N_5277,N_3035,N_3177);
xnor U5278 (N_5278,N_1941,N_1592);
nor U5279 (N_5279,N_4336,N_2598);
xor U5280 (N_5280,N_3653,N_1564);
and U5281 (N_5281,N_1364,N_2280);
or U5282 (N_5282,N_3172,N_2762);
xnor U5283 (N_5283,N_774,N_740);
and U5284 (N_5284,N_191,N_3301);
and U5285 (N_5285,N_1914,N_4376);
xnor U5286 (N_5286,N_4040,N_442);
nor U5287 (N_5287,N_3851,N_4115);
or U5288 (N_5288,N_1273,N_1713);
and U5289 (N_5289,N_4187,N_3124);
nor U5290 (N_5290,N_1374,N_2513);
nor U5291 (N_5291,N_266,N_37);
nor U5292 (N_5292,N_35,N_3892);
and U5293 (N_5293,N_2866,N_2321);
and U5294 (N_5294,N_1252,N_2150);
xnor U5295 (N_5295,N_1605,N_278);
nand U5296 (N_5296,N_382,N_2740);
xnor U5297 (N_5297,N_267,N_2596);
and U5298 (N_5298,N_4927,N_200);
or U5299 (N_5299,N_1484,N_2664);
xor U5300 (N_5300,N_2311,N_4094);
nand U5301 (N_5301,N_1577,N_3069);
nand U5302 (N_5302,N_315,N_2826);
or U5303 (N_5303,N_2494,N_2023);
nor U5304 (N_5304,N_2703,N_1693);
or U5305 (N_5305,N_4144,N_3847);
or U5306 (N_5306,N_1581,N_874);
and U5307 (N_5307,N_170,N_3933);
and U5308 (N_5308,N_2285,N_3604);
nand U5309 (N_5309,N_1113,N_4600);
or U5310 (N_5310,N_656,N_1657);
nand U5311 (N_5311,N_3500,N_3897);
nor U5312 (N_5312,N_2988,N_1835);
nand U5313 (N_5313,N_4062,N_2391);
xnor U5314 (N_5314,N_2899,N_1791);
nor U5315 (N_5315,N_2131,N_3886);
and U5316 (N_5316,N_4860,N_3215);
nor U5317 (N_5317,N_1292,N_4442);
nand U5318 (N_5318,N_3207,N_2501);
nor U5319 (N_5319,N_3466,N_3366);
xor U5320 (N_5320,N_4989,N_3181);
nor U5321 (N_5321,N_1362,N_3737);
xnor U5322 (N_5322,N_3916,N_3581);
nand U5323 (N_5323,N_259,N_2745);
xnor U5324 (N_5324,N_38,N_1363);
and U5325 (N_5325,N_4780,N_1606);
or U5326 (N_5326,N_3606,N_968);
xor U5327 (N_5327,N_2856,N_979);
nand U5328 (N_5328,N_2694,N_4145);
nor U5329 (N_5329,N_2483,N_1895);
nand U5330 (N_5330,N_4285,N_3987);
xnor U5331 (N_5331,N_1811,N_149);
nor U5332 (N_5332,N_2317,N_4621);
and U5333 (N_5333,N_3184,N_3774);
and U5334 (N_5334,N_1286,N_2814);
xnor U5335 (N_5335,N_326,N_3795);
and U5336 (N_5336,N_4569,N_860);
and U5337 (N_5337,N_4411,N_1388);
or U5338 (N_5338,N_1124,N_4224);
nand U5339 (N_5339,N_3928,N_1697);
or U5340 (N_5340,N_4455,N_1524);
xnor U5341 (N_5341,N_1348,N_1142);
and U5342 (N_5342,N_4527,N_3585);
nor U5343 (N_5343,N_279,N_4503);
xnor U5344 (N_5344,N_2450,N_2926);
nor U5345 (N_5345,N_4982,N_4959);
nand U5346 (N_5346,N_3050,N_1404);
nor U5347 (N_5347,N_4196,N_2532);
xnor U5348 (N_5348,N_4673,N_1206);
nor U5349 (N_5349,N_4021,N_362);
and U5350 (N_5350,N_2669,N_1922);
nor U5351 (N_5351,N_875,N_4033);
nand U5352 (N_5352,N_351,N_948);
or U5353 (N_5353,N_1258,N_82);
xnor U5354 (N_5354,N_319,N_3570);
and U5355 (N_5355,N_3922,N_145);
nor U5356 (N_5356,N_2749,N_4852);
nor U5357 (N_5357,N_960,N_306);
nor U5358 (N_5358,N_2661,N_4242);
xor U5359 (N_5359,N_3979,N_783);
xor U5360 (N_5360,N_1143,N_1955);
nor U5361 (N_5361,N_4995,N_544);
and U5362 (N_5362,N_4106,N_2770);
and U5363 (N_5363,N_1190,N_558);
nand U5364 (N_5364,N_3212,N_4559);
and U5365 (N_5365,N_1942,N_3200);
nand U5366 (N_5366,N_709,N_1281);
nand U5367 (N_5367,N_97,N_2266);
and U5368 (N_5368,N_2429,N_3914);
xnor U5369 (N_5369,N_517,N_4976);
nand U5370 (N_5370,N_4866,N_2458);
xor U5371 (N_5371,N_2011,N_2416);
nor U5372 (N_5372,N_2277,N_2407);
xnor U5373 (N_5373,N_4041,N_3423);
xnor U5374 (N_5374,N_3236,N_4702);
nand U5375 (N_5375,N_1159,N_2717);
nor U5376 (N_5376,N_1235,N_3980);
and U5377 (N_5377,N_1792,N_3694);
xor U5378 (N_5378,N_4592,N_467);
nor U5379 (N_5379,N_1155,N_91);
xor U5380 (N_5380,N_1371,N_4102);
xor U5381 (N_5381,N_3224,N_744);
xor U5382 (N_5382,N_4921,N_2561);
or U5383 (N_5383,N_3874,N_923);
or U5384 (N_5384,N_1398,N_2937);
or U5385 (N_5385,N_1610,N_4310);
and U5386 (N_5386,N_4251,N_14);
and U5387 (N_5387,N_952,N_1343);
or U5388 (N_5388,N_2460,N_1491);
and U5389 (N_5389,N_2482,N_2336);
or U5390 (N_5390,N_4713,N_4245);
or U5391 (N_5391,N_2748,N_2132);
and U5392 (N_5392,N_2028,N_2674);
nand U5393 (N_5393,N_1907,N_4210);
nor U5394 (N_5394,N_318,N_1285);
or U5395 (N_5395,N_2445,N_2078);
xor U5396 (N_5396,N_3401,N_3491);
or U5397 (N_5397,N_4421,N_4191);
or U5398 (N_5398,N_1486,N_4198);
or U5399 (N_5399,N_4299,N_2168);
and U5400 (N_5400,N_4871,N_3032);
nor U5401 (N_5401,N_4602,N_4834);
nand U5402 (N_5402,N_4221,N_3811);
and U5403 (N_5403,N_825,N_350);
or U5404 (N_5404,N_2139,N_4039);
or U5405 (N_5405,N_269,N_461);
and U5406 (N_5406,N_3726,N_3263);
nor U5407 (N_5407,N_701,N_4468);
or U5408 (N_5408,N_3576,N_2766);
nor U5409 (N_5409,N_1223,N_2504);
and U5410 (N_5410,N_3887,N_2466);
nand U5411 (N_5411,N_3095,N_474);
or U5412 (N_5412,N_2035,N_3787);
xnor U5413 (N_5413,N_2251,N_4497);
nand U5414 (N_5414,N_3147,N_2275);
or U5415 (N_5415,N_547,N_3915);
or U5416 (N_5416,N_4109,N_1921);
and U5417 (N_5417,N_1603,N_4547);
and U5418 (N_5418,N_4926,N_312);
nor U5419 (N_5419,N_791,N_3504);
or U5420 (N_5420,N_3120,N_4888);
or U5421 (N_5421,N_4416,N_633);
and U5422 (N_5422,N_3294,N_794);
xor U5423 (N_5423,N_3169,N_4370);
and U5424 (N_5424,N_449,N_1541);
nor U5425 (N_5425,N_2452,N_488);
xnor U5426 (N_5426,N_3415,N_878);
or U5427 (N_5427,N_3447,N_4156);
and U5428 (N_5428,N_141,N_51);
nor U5429 (N_5429,N_645,N_4509);
or U5430 (N_5430,N_3605,N_383);
xnor U5431 (N_5431,N_3307,N_1308);
nor U5432 (N_5432,N_1150,N_1925);
xor U5433 (N_5433,N_782,N_3258);
nand U5434 (N_5434,N_2662,N_4177);
nor U5435 (N_5435,N_199,N_1939);
nor U5436 (N_5436,N_4828,N_1629);
and U5437 (N_5437,N_3245,N_2489);
nor U5438 (N_5438,N_357,N_83);
xor U5439 (N_5439,N_3953,N_1400);
or U5440 (N_5440,N_2581,N_2716);
and U5441 (N_5441,N_21,N_3102);
or U5442 (N_5442,N_2086,N_296);
or U5443 (N_5443,N_2995,N_4167);
nor U5444 (N_5444,N_1294,N_2276);
and U5445 (N_5445,N_2064,N_2835);
or U5446 (N_5446,N_1684,N_4603);
or U5447 (N_5447,N_4804,N_102);
nor U5448 (N_5448,N_808,N_3703);
or U5449 (N_5449,N_1399,N_1641);
nor U5450 (N_5450,N_317,N_3691);
and U5451 (N_5451,N_1157,N_30);
xnor U5452 (N_5452,N_3678,N_4855);
xor U5453 (N_5453,N_3218,N_1613);
or U5454 (N_5454,N_4841,N_4202);
or U5455 (N_5455,N_3052,N_1528);
and U5456 (N_5456,N_15,N_2014);
nor U5457 (N_5457,N_3094,N_1867);
xor U5458 (N_5458,N_4643,N_3000);
and U5459 (N_5459,N_4744,N_1100);
xnor U5460 (N_5460,N_2007,N_1358);
nand U5461 (N_5461,N_1130,N_2617);
or U5462 (N_5462,N_3148,N_1063);
xor U5463 (N_5463,N_2824,N_4674);
nor U5464 (N_5464,N_2213,N_336);
xnor U5465 (N_5465,N_4058,N_624);
xnor U5466 (N_5466,N_4844,N_248);
xnor U5467 (N_5467,N_2208,N_4531);
xnor U5468 (N_5468,N_46,N_1287);
nor U5469 (N_5469,N_1499,N_1800);
nor U5470 (N_5470,N_1489,N_764);
xnor U5471 (N_5471,N_426,N_2122);
nor U5472 (N_5472,N_2370,N_3011);
nor U5473 (N_5473,N_3128,N_4119);
nand U5474 (N_5474,N_2037,N_642);
nand U5475 (N_5475,N_1803,N_2910);
xnor U5476 (N_5476,N_4382,N_3937);
nand U5477 (N_5477,N_3896,N_3063);
nor U5478 (N_5478,N_4637,N_365);
and U5479 (N_5479,N_359,N_4225);
nor U5480 (N_5480,N_612,N_2081);
nor U5481 (N_5481,N_25,N_1824);
and U5482 (N_5482,N_3590,N_793);
and U5483 (N_5483,N_2462,N_997);
xor U5484 (N_5484,N_3586,N_4881);
nor U5485 (N_5485,N_3310,N_687);
or U5486 (N_5486,N_3284,N_2524);
or U5487 (N_5487,N_3076,N_2141);
nand U5488 (N_5488,N_3167,N_3690);
xnor U5489 (N_5489,N_2454,N_562);
and U5490 (N_5490,N_1134,N_1616);
nand U5491 (N_5491,N_2060,N_710);
and U5492 (N_5492,N_2263,N_2772);
or U5493 (N_5493,N_4387,N_1796);
and U5494 (N_5494,N_4189,N_2880);
nor U5495 (N_5495,N_4303,N_3390);
or U5496 (N_5496,N_4818,N_64);
nand U5497 (N_5497,N_213,N_1643);
xor U5498 (N_5498,N_4965,N_3664);
nand U5499 (N_5499,N_1115,N_3536);
and U5500 (N_5500,N_4884,N_873);
or U5501 (N_5501,N_843,N_2158);
nor U5502 (N_5502,N_3525,N_2048);
or U5503 (N_5503,N_1567,N_657);
or U5504 (N_5504,N_1379,N_2374);
nor U5505 (N_5505,N_404,N_2025);
nand U5506 (N_5506,N_4561,N_1561);
nor U5507 (N_5507,N_4163,N_3345);
or U5508 (N_5508,N_4313,N_1901);
and U5509 (N_5509,N_2205,N_1576);
xor U5510 (N_5510,N_2022,N_4652);
or U5511 (N_5511,N_3022,N_1161);
and U5512 (N_5512,N_4283,N_4676);
nor U5513 (N_5513,N_2451,N_3657);
and U5514 (N_5514,N_2534,N_1819);
nor U5515 (N_5515,N_4013,N_1808);
or U5516 (N_5516,N_2704,N_3643);
or U5517 (N_5517,N_1201,N_2877);
or U5518 (N_5518,N_2124,N_4916);
nand U5519 (N_5519,N_795,N_189);
and U5520 (N_5520,N_4711,N_3573);
nand U5521 (N_5521,N_3601,N_3666);
and U5522 (N_5522,N_1275,N_2714);
and U5523 (N_5523,N_3551,N_3505);
nor U5524 (N_5524,N_142,N_3385);
xor U5525 (N_5525,N_4932,N_2255);
or U5526 (N_5526,N_2929,N_4714);
xor U5527 (N_5527,N_3322,N_1177);
nand U5528 (N_5528,N_4038,N_4082);
nor U5529 (N_5529,N_2512,N_748);
or U5530 (N_5530,N_1533,N_4629);
nor U5531 (N_5531,N_489,N_3323);
xnor U5532 (N_5532,N_4023,N_4566);
and U5533 (N_5533,N_3004,N_1141);
xnor U5534 (N_5534,N_3289,N_2620);
xnor U5535 (N_5535,N_3946,N_1497);
nor U5536 (N_5536,N_3830,N_50);
xnor U5537 (N_5537,N_1785,N_736);
or U5538 (N_5538,N_4,N_1753);
or U5539 (N_5539,N_158,N_2500);
nor U5540 (N_5540,N_611,N_853);
nand U5541 (N_5541,N_2960,N_2806);
nand U5542 (N_5542,N_3526,N_3140);
xnor U5543 (N_5543,N_3472,N_2977);
xor U5544 (N_5544,N_4513,N_651);
or U5545 (N_5545,N_4528,N_3826);
xnor U5546 (N_5546,N_3676,N_4707);
nor U5547 (N_5547,N_2101,N_3144);
xor U5548 (N_5548,N_193,N_4112);
nand U5549 (N_5549,N_4864,N_3460);
and U5550 (N_5550,N_2328,N_4799);
and U5551 (N_5551,N_2281,N_3718);
nand U5552 (N_5552,N_4580,N_618);
or U5553 (N_5553,N_2110,N_3813);
nand U5554 (N_5554,N_6,N_4615);
xnor U5555 (N_5555,N_4810,N_1587);
xor U5556 (N_5556,N_2216,N_2093);
and U5557 (N_5557,N_591,N_4742);
xnor U5558 (N_5558,N_504,N_3162);
xnor U5559 (N_5559,N_4176,N_4051);
and U5560 (N_5560,N_1414,N_1751);
xnor U5561 (N_5561,N_4677,N_3842);
or U5562 (N_5562,N_2538,N_4447);
xor U5563 (N_5563,N_4759,N_2409);
nor U5564 (N_5564,N_3705,N_2257);
and U5565 (N_5565,N_3539,N_674);
or U5566 (N_5566,N_3966,N_2400);
and U5567 (N_5567,N_3701,N_1966);
or U5568 (N_5568,N_4630,N_4653);
and U5569 (N_5569,N_2901,N_389);
nand U5570 (N_5570,N_2556,N_4220);
nand U5571 (N_5571,N_3599,N_1085);
nor U5572 (N_5572,N_2943,N_1887);
and U5573 (N_5573,N_3518,N_1648);
or U5574 (N_5574,N_750,N_4315);
nor U5575 (N_5575,N_1507,N_1666);
or U5576 (N_5576,N_2514,N_1560);
xor U5577 (N_5577,N_1845,N_1276);
or U5578 (N_5578,N_2411,N_1016);
or U5579 (N_5579,N_934,N_1076);
or U5580 (N_5580,N_2498,N_2771);
xnor U5581 (N_5581,N_4074,N_3336);
xor U5582 (N_5582,N_4459,N_499);
and U5583 (N_5583,N_3940,N_2984);
nand U5584 (N_5584,N_4779,N_2186);
nor U5585 (N_5585,N_1823,N_2886);
and U5586 (N_5586,N_1553,N_242);
or U5587 (N_5587,N_4341,N_1466);
and U5588 (N_5588,N_1972,N_2575);
and U5589 (N_5589,N_3220,N_4549);
nand U5590 (N_5590,N_970,N_165);
or U5591 (N_5591,N_1212,N_615);
and U5592 (N_5592,N_2792,N_4152);
nor U5593 (N_5593,N_1957,N_2423);
or U5594 (N_5594,N_1772,N_630);
nand U5595 (N_5595,N_3889,N_2226);
nor U5596 (N_5596,N_518,N_3299);
and U5597 (N_5597,N_3112,N_3867);
nor U5598 (N_5598,N_26,N_3202);
and U5599 (N_5599,N_1199,N_3552);
or U5600 (N_5600,N_1970,N_4334);
or U5601 (N_5601,N_487,N_3347);
nor U5602 (N_5602,N_3092,N_2849);
nand U5603 (N_5603,N_731,N_4797);
or U5604 (N_5604,N_4766,N_78);
nand U5605 (N_5605,N_3815,N_3837);
nor U5606 (N_5606,N_4008,N_506);
xnor U5607 (N_5607,N_3636,N_2376);
nor U5608 (N_5608,N_2380,N_2818);
and U5609 (N_5609,N_1602,N_2791);
or U5610 (N_5610,N_2414,N_2261);
nand U5611 (N_5611,N_1301,N_2428);
nor U5612 (N_5612,N_1815,N_3444);
nand U5613 (N_5613,N_1207,N_250);
nand U5614 (N_5614,N_3136,N_2742);
nor U5615 (N_5615,N_2719,N_4378);
nand U5616 (N_5616,N_2225,N_3231);
or U5617 (N_5617,N_147,N_2410);
or U5618 (N_5618,N_1989,N_3165);
xor U5619 (N_5619,N_156,N_870);
nor U5620 (N_5620,N_613,N_2905);
xnor U5621 (N_5621,N_1107,N_2541);
nor U5622 (N_5622,N_409,N_1632);
nand U5623 (N_5623,N_667,N_2293);
or U5624 (N_5624,N_101,N_4036);
nor U5625 (N_5625,N_2046,N_1319);
xnor U5626 (N_5626,N_3371,N_502);
nand U5627 (N_5627,N_123,N_4875);
nor U5628 (N_5628,N_2619,N_3033);
or U5629 (N_5629,N_3449,N_4043);
or U5630 (N_5630,N_3317,N_3244);
or U5631 (N_5631,N_3359,N_431);
and U5632 (N_5632,N_545,N_1563);
or U5633 (N_5633,N_4142,N_1488);
and U5634 (N_5634,N_1668,N_3091);
and U5635 (N_5635,N_2523,N_2823);
or U5636 (N_5636,N_3062,N_67);
and U5637 (N_5637,N_2892,N_1034);
xor U5638 (N_5638,N_4577,N_4925);
or U5639 (N_5639,N_3252,N_1451);
or U5640 (N_5640,N_1805,N_3469);
or U5641 (N_5641,N_1164,N_778);
nand U5642 (N_5642,N_3517,N_1209);
nand U5643 (N_5643,N_3982,N_73);
xor U5644 (N_5644,N_2089,N_458);
and U5645 (N_5645,N_445,N_1526);
nor U5646 (N_5646,N_2785,N_3414);
and U5647 (N_5647,N_3925,N_1282);
nor U5648 (N_5648,N_3365,N_490);
and U5649 (N_5649,N_2088,N_4227);
xnor U5650 (N_5650,N_3721,N_4261);
and U5651 (N_5651,N_695,N_3758);
and U5652 (N_5652,N_2819,N_1295);
and U5653 (N_5653,N_2911,N_3992);
xor U5654 (N_5654,N_2828,N_4223);
xor U5655 (N_5655,N_4758,N_1825);
nand U5656 (N_5656,N_1296,N_634);
xnor U5657 (N_5657,N_4774,N_4699);
or U5658 (N_5658,N_253,N_4782);
or U5659 (N_5659,N_4084,N_1920);
nand U5660 (N_5660,N_2472,N_1706);
and U5661 (N_5661,N_594,N_4769);
xor U5662 (N_5662,N_1879,N_4035);
nor U5663 (N_5663,N_3073,N_4839);
and U5664 (N_5664,N_1102,N_3684);
nand U5665 (N_5665,N_879,N_4317);
nand U5666 (N_5666,N_2238,N_3059);
nand U5667 (N_5667,N_1013,N_2180);
xor U5668 (N_5668,N_4762,N_2525);
nand U5669 (N_5669,N_1459,N_408);
and U5670 (N_5670,N_2699,N_1762);
nand U5671 (N_5671,N_99,N_208);
nor U5672 (N_5672,N_711,N_4848);
and U5673 (N_5673,N_2375,N_4037);
nor U5674 (N_5674,N_2034,N_309);
or U5675 (N_5675,N_1111,N_1969);
nand U5676 (N_5676,N_2170,N_3750);
or U5677 (N_5677,N_183,N_2455);
and U5678 (N_5678,N_3964,N_4743);
and U5679 (N_5679,N_2228,N_2659);
xnor U5680 (N_5680,N_2630,N_4019);
nand U5681 (N_5681,N_1623,N_1555);
xor U5682 (N_5682,N_3733,N_1051);
nand U5683 (N_5683,N_2320,N_2070);
nand U5684 (N_5684,N_4647,N_2340);
or U5685 (N_5685,N_2726,N_4890);
nand U5686 (N_5686,N_2734,N_2913);
xor U5687 (N_5687,N_2272,N_3617);
and U5688 (N_5688,N_707,N_4878);
and U5689 (N_5689,N_2848,N_4660);
xnor U5690 (N_5690,N_1608,N_4980);
nand U5691 (N_5691,N_1014,N_1234);
xor U5692 (N_5692,N_1326,N_1847);
xnor U5693 (N_5693,N_2269,N_3146);
xor U5694 (N_5694,N_1779,N_1667);
and U5695 (N_5695,N_1638,N_702);
xnor U5696 (N_5696,N_2570,N_1537);
xnor U5697 (N_5697,N_3273,N_3494);
nor U5698 (N_5698,N_1927,N_4483);
xnor U5699 (N_5699,N_2608,N_55);
xor U5700 (N_5700,N_98,N_1672);
or U5701 (N_5701,N_446,N_60);
nor U5702 (N_5702,N_1365,N_2434);
nand U5703 (N_5703,N_1501,N_1833);
nor U5704 (N_5704,N_1008,N_3878);
and U5705 (N_5705,N_4325,N_3535);
and U5706 (N_5706,N_1423,N_678);
or U5707 (N_5707,N_1594,N_3338);
or U5708 (N_5708,N_781,N_366);
nand U5709 (N_5709,N_4598,N_2869);
and U5710 (N_5710,N_3580,N_2667);
or U5711 (N_5711,N_1182,N_9);
and U5712 (N_5712,N_2867,N_2144);
nor U5713 (N_5713,N_4882,N_2395);
nor U5714 (N_5714,N_1698,N_1215);
nor U5715 (N_5715,N_2840,N_2419);
and U5716 (N_5716,N_652,N_4463);
xnor U5717 (N_5717,N_3089,N_2938);
xnor U5718 (N_5718,N_2453,N_4252);
xnor U5719 (N_5719,N_4135,N_1325);
and U5720 (N_5720,N_192,N_3781);
nand U5721 (N_5721,N_4607,N_4164);
nor U5722 (N_5722,N_420,N_2887);
nor U5723 (N_5723,N_1053,N_364);
nand U5724 (N_5724,N_2114,N_255);
and U5725 (N_5725,N_1392,N_1447);
nand U5726 (N_5726,N_1316,N_4856);
and U5727 (N_5727,N_3039,N_2790);
or U5728 (N_5728,N_4379,N_4319);
or U5729 (N_5729,N_3192,N_4014);
nand U5730 (N_5730,N_3341,N_2865);
nand U5731 (N_5731,N_2422,N_4692);
or U5732 (N_5732,N_2218,N_3480);
nor U5733 (N_5733,N_4388,N_2424);
nand U5734 (N_5734,N_249,N_4715);
and U5735 (N_5735,N_1882,N_2587);
nor U5736 (N_5736,N_2822,N_4872);
and U5737 (N_5737,N_4136,N_2551);
or U5738 (N_5738,N_3735,N_3665);
nand U5739 (N_5739,N_2634,N_2952);
nor U5740 (N_5740,N_909,N_2767);
nor U5741 (N_5741,N_2545,N_136);
and U5742 (N_5742,N_324,N_174);
nor U5743 (N_5743,N_4933,N_3446);
nor U5744 (N_5744,N_1443,N_4530);
nor U5745 (N_5745,N_3197,N_734);
nor U5746 (N_5746,N_2480,N_143);
nand U5747 (N_5747,N_3014,N_1601);
nor U5748 (N_5748,N_3318,N_4061);
xor U5749 (N_5749,N_3647,N_1302);
nor U5750 (N_5750,N_22,N_4908);
or U5751 (N_5751,N_407,N_525);
nor U5752 (N_5752,N_988,N_373);
or U5753 (N_5753,N_3099,N_4383);
and U5754 (N_5754,N_4662,N_1733);
and U5755 (N_5755,N_2302,N_718);
or U5756 (N_5756,N_4433,N_2665);
nor U5757 (N_5757,N_3720,N_4845);
and U5758 (N_5758,N_230,N_792);
nor U5759 (N_5759,N_2858,N_1291);
and U5760 (N_5760,N_3483,N_4090);
or U5761 (N_5761,N_4764,N_680);
xor U5762 (N_5762,N_4281,N_4955);
xnor U5763 (N_5763,N_2879,N_3303);
and U5764 (N_5764,N_818,N_2342);
xnor U5765 (N_5765,N_1731,N_976);
nor U5766 (N_5766,N_2127,N_1571);
nand U5767 (N_5767,N_4806,N_4292);
xnor U5768 (N_5768,N_2256,N_1401);
or U5769 (N_5769,N_3680,N_3264);
or U5770 (N_5770,N_4434,N_1193);
nor U5771 (N_5771,N_4272,N_2431);
or U5772 (N_5772,N_1906,N_666);
nand U5773 (N_5773,N_2989,N_649);
nand U5774 (N_5774,N_1284,N_1208);
nor U5775 (N_5775,N_70,N_4861);
and U5776 (N_5776,N_2262,N_1198);
or U5777 (N_5777,N_2555,N_990);
or U5778 (N_5778,N_3698,N_1412);
nand U5779 (N_5779,N_3614,N_1937);
xnor U5780 (N_5780,N_2005,N_2628);
or U5781 (N_5781,N_4093,N_4990);
and U5782 (N_5782,N_2672,N_2673);
nand U5783 (N_5783,N_1407,N_787);
nand U5784 (N_5784,N_4488,N_3625);
and U5785 (N_5785,N_1173,N_4776);
or U5786 (N_5786,N_4649,N_4877);
xnor U5787 (N_5787,N_2692,N_4393);
and U5788 (N_5788,N_966,N_3870);
nand U5789 (N_5789,N_961,N_2087);
nand U5790 (N_5790,N_3051,N_2301);
nand U5791 (N_5791,N_4801,N_3122);
and U5792 (N_5792,N_3532,N_1630);
nor U5793 (N_5793,N_2360,N_1912);
or U5794 (N_5794,N_3511,N_3311);
or U5795 (N_5795,N_646,N_4672);
nand U5796 (N_5796,N_2465,N_3267);
and U5797 (N_5797,N_4519,N_4941);
and U5798 (N_5798,N_185,N_2846);
and U5799 (N_5799,N_2092,N_2975);
and U5800 (N_5800,N_1056,N_597);
and U5801 (N_5801,N_4606,N_2339);
nor U5802 (N_5802,N_607,N_4827);
nor U5803 (N_5803,N_1178,N_4101);
xor U5804 (N_5804,N_1624,N_2578);
or U5805 (N_5805,N_310,N_1493);
or U5806 (N_5806,N_3530,N_2121);
nand U5807 (N_5807,N_2039,N_983);
or U5808 (N_5808,N_2685,N_2172);
nor U5809 (N_5809,N_4618,N_4970);
nand U5810 (N_5810,N_724,N_4168);
nand U5811 (N_5811,N_2983,N_2558);
nand U5812 (N_5812,N_1730,N_1116);
nor U5813 (N_5813,N_477,N_974);
nand U5814 (N_5814,N_836,N_47);
xnor U5815 (N_5815,N_1749,N_1554);
xor U5816 (N_5816,N_4131,N_4004);
xor U5817 (N_5817,N_384,N_4162);
nand U5818 (N_5818,N_3261,N_3766);
and U5819 (N_5819,N_4581,N_34);
or U5820 (N_5820,N_1170,N_2833);
or U5821 (N_5821,N_851,N_2776);
or U5822 (N_5822,N_1965,N_2530);
nor U5823 (N_5823,N_3951,N_4646);
or U5824 (N_5824,N_1510,N_61);
nor U5825 (N_5825,N_2547,N_3514);
xor U5826 (N_5826,N_1839,N_1857);
or U5827 (N_5827,N_1998,N_342);
and U5828 (N_5828,N_2154,N_859);
and U5829 (N_5829,N_4663,N_2357);
and U5830 (N_5830,N_1331,N_3926);
nor U5831 (N_5831,N_629,N_3107);
or U5832 (N_5832,N_3563,N_4719);
xnor U5833 (N_5833,N_3234,N_1242);
nor U5834 (N_5834,N_1354,N_3204);
nand U5835 (N_5835,N_553,N_289);
or U5836 (N_5836,N_3150,N_2059);
nand U5837 (N_5837,N_2471,N_4737);
and U5838 (N_5838,N_3989,N_1003);
xnor U5839 (N_5839,N_4917,N_4678);
nor U5840 (N_5840,N_3049,N_3574);
nor U5841 (N_5841,N_2593,N_4288);
or U5842 (N_5842,N_1088,N_205);
and U5843 (N_5843,N_980,N_1818);
xor U5844 (N_5844,N_2250,N_3848);
xor U5845 (N_5845,N_2220,N_1574);
xor U5846 (N_5846,N_1758,N_2143);
or U5847 (N_5847,N_819,N_3553);
or U5848 (N_5848,N_2712,N_745);
nand U5849 (N_5849,N_1761,N_1090);
and U5850 (N_5850,N_3040,N_2802);
or U5851 (N_5851,N_4020,N_1069);
nor U5852 (N_5852,N_1782,N_167);
or U5853 (N_5853,N_4956,N_3769);
xor U5854 (N_5854,N_462,N_1442);
xnor U5855 (N_5855,N_273,N_3777);
and U5856 (N_5856,N_2217,N_683);
nand U5857 (N_5857,N_1048,N_741);
nor U5858 (N_5858,N_4948,N_3641);
nor U5859 (N_5859,N_993,N_2808);
nand U5860 (N_5860,N_768,N_3357);
or U5861 (N_5861,N_2981,N_4560);
xor U5862 (N_5862,N_672,N_3298);
or U5863 (N_5863,N_1938,N_4332);
and U5864 (N_5864,N_1512,N_2167);
nand U5865 (N_5865,N_4161,N_3210);
xnor U5866 (N_5866,N_4523,N_3361);
xor U5867 (N_5867,N_585,N_1891);
nor U5868 (N_5868,N_184,N_1963);
nor U5869 (N_5869,N_2437,N_2747);
and U5870 (N_5870,N_885,N_2591);
or U5871 (N_5871,N_3426,N_1087);
or U5872 (N_5872,N_3241,N_523);
nand U5873 (N_5873,N_1405,N_3380);
or U5874 (N_5874,N_3621,N_1127);
nand U5875 (N_5875,N_1763,N_4282);
and U5876 (N_5876,N_75,N_3900);
nand U5877 (N_5877,N_2234,N_2820);
or U5878 (N_5878,N_2928,N_1058);
nand U5879 (N_5879,N_4121,N_2299);
nand U5880 (N_5880,N_4444,N_473);
and U5881 (N_5881,N_3615,N_1031);
nor U5882 (N_5882,N_770,N_4403);
and U5883 (N_5883,N_3890,N_1086);
nand U5884 (N_5884,N_2464,N_4301);
nand U5885 (N_5885,N_944,N_1977);
xor U5886 (N_5886,N_2793,N_133);
and U5887 (N_5887,N_3789,N_1479);
and U5888 (N_5888,N_3908,N_4558);
or U5889 (N_5889,N_2676,N_1213);
xnor U5890 (N_5890,N_930,N_1030);
nor U5891 (N_5891,N_1660,N_4178);
nor U5892 (N_5892,N_620,N_333);
or U5893 (N_5893,N_2386,N_2842);
or U5894 (N_5894,N_3759,N_1425);
and U5895 (N_5895,N_4408,N_1615);
nor U5896 (N_5896,N_4495,N_4031);
xnor U5897 (N_5897,N_2544,N_2537);
nor U5898 (N_5898,N_3521,N_3369);
nand U5899 (N_5899,N_3806,N_951);
and U5900 (N_5900,N_3493,N_2058);
nor U5901 (N_5901,N_4626,N_2559);
xor U5902 (N_5902,N_985,N_829);
nand U5903 (N_5903,N_959,N_1994);
and U5904 (N_5904,N_3860,N_1618);
nand U5905 (N_5905,N_2907,N_4732);
nand U5906 (N_5906,N_2417,N_3306);
and U5907 (N_5907,N_4147,N_2182);
nor U5908 (N_5908,N_2954,N_4633);
and U5909 (N_5909,N_2600,N_424);
and U5910 (N_5910,N_2588,N_419);
xor U5911 (N_5911,N_2349,N_2175);
xor U5912 (N_5912,N_4893,N_1741);
or U5913 (N_5913,N_2564,N_1842);
nand U5914 (N_5914,N_1790,N_1547);
xnor U5915 (N_5915,N_4099,N_1469);
xnor U5916 (N_5916,N_1002,N_4892);
nand U5917 (N_5917,N_3962,N_4472);
nor U5918 (N_5918,N_3840,N_2736);
nor U5919 (N_5919,N_1612,N_2845);
nand U5920 (N_5920,N_3963,N_390);
nor U5921 (N_5921,N_4883,N_4409);
and U5922 (N_5922,N_2098,N_3846);
xnor U5923 (N_5923,N_676,N_3008);
or U5924 (N_5924,N_95,N_1902);
and U5925 (N_5925,N_4693,N_3748);
or U5926 (N_5926,N_4486,N_1968);
and U5927 (N_5927,N_19,N_4271);
and U5928 (N_5928,N_1556,N_1336);
nor U5929 (N_5929,N_2111,N_3398);
nand U5930 (N_5930,N_4962,N_3044);
or U5931 (N_5931,N_3249,N_1997);
nand U5932 (N_5932,N_1351,N_239);
or U5933 (N_5933,N_928,N_2056);
nand U5934 (N_5934,N_568,N_4756);
xnor U5935 (N_5935,N_2962,N_3949);
xnor U5936 (N_5936,N_660,N_2485);
nor U5937 (N_5937,N_869,N_3760);
nor U5938 (N_5938,N_1473,N_845);
nand U5939 (N_5939,N_4305,N_522);
or U5940 (N_5940,N_2119,N_1934);
or U5941 (N_5941,N_4431,N_4553);
xnor U5942 (N_5942,N_4485,N_3961);
or U5943 (N_5943,N_4645,N_2288);
nor U5944 (N_5944,N_4584,N_2961);
or U5945 (N_5945,N_4650,N_1032);
nor U5946 (N_5946,N_3282,N_1679);
nand U5947 (N_5947,N_3818,N_3632);
or U5948 (N_5948,N_2194,N_3278);
xnor U5949 (N_5949,N_4316,N_3602);
nor U5950 (N_5950,N_284,N_3616);
xnor U5951 (N_5951,N_1896,N_1642);
nand U5952 (N_5952,N_809,N_922);
and U5953 (N_5953,N_941,N_4195);
or U5954 (N_5954,N_94,N_1018);
xor U5955 (N_5955,N_227,N_1191);
xnor U5956 (N_5956,N_1269,N_1474);
nor U5957 (N_5957,N_1723,N_2072);
or U5958 (N_5958,N_800,N_3296);
nand U5959 (N_5959,N_4267,N_3045);
or U5960 (N_5960,N_2594,N_476);
or U5961 (N_5961,N_4182,N_3);
xnor U5962 (N_5962,N_1184,N_115);
nand U5963 (N_5963,N_2053,N_3516);
xor U5964 (N_5964,N_2337,N_435);
or U5965 (N_5965,N_2870,N_1408);
or U5966 (N_5966,N_810,N_4389);
nand U5967 (N_5967,N_830,N_3911);
nand U5968 (N_5968,N_2009,N_1788);
nor U5969 (N_5969,N_4757,N_2724);
and U5970 (N_5970,N_4005,N_4364);
or U5971 (N_5971,N_1784,N_2580);
nor U5972 (N_5972,N_3749,N_958);
nand U5973 (N_5973,N_771,N_4201);
and U5974 (N_5974,N_4138,N_4909);
xor U5975 (N_5975,N_2902,N_2966);
nor U5976 (N_5976,N_2406,N_1810);
nor U5977 (N_5977,N_4266,N_3740);
or U5978 (N_5978,N_3326,N_3348);
or U5979 (N_5979,N_840,N_1065);
nor U5980 (N_5980,N_4237,N_4735);
and U5981 (N_5981,N_3861,N_3998);
or U5982 (N_5982,N_4924,N_1531);
xnor U5983 (N_5983,N_514,N_493);
nor U5984 (N_5984,N_797,N_4335);
or U5985 (N_5985,N_4675,N_4006);
or U5986 (N_5986,N_3973,N_3854);
nand U5987 (N_5987,N_2721,N_4682);
nor U5988 (N_5988,N_321,N_2589);
nand U5989 (N_5989,N_2979,N_4906);
or U5990 (N_5990,N_1446,N_3708);
and U5991 (N_5991,N_410,N_2972);
nand U5992 (N_5992,N_1777,N_443);
nor U5993 (N_5993,N_2957,N_972);
xor U5994 (N_5994,N_4028,N_4357);
or U5995 (N_5995,N_2754,N_1084);
nand U5996 (N_5996,N_772,N_1240);
xor U5997 (N_5997,N_1746,N_3677);
nand U5998 (N_5998,N_670,N_2741);
and U5999 (N_5999,N_1009,N_2584);
xor U6000 (N_6000,N_2109,N_4492);
or U6001 (N_6001,N_2197,N_4209);
or U6002 (N_6002,N_2355,N_3891);
nor U6003 (N_6003,N_3770,N_4072);
xor U6004 (N_6004,N_939,N_2604);
xor U6005 (N_6005,N_2998,N_345);
xor U6006 (N_6006,N_1764,N_4920);
nand U6007 (N_6007,N_2207,N_4658);
and U6008 (N_6008,N_1646,N_696);
or U6009 (N_6009,N_4972,N_2068);
or U6010 (N_6010,N_3741,N_2050);
or U6011 (N_6011,N_1136,N_2373);
nand U6012 (N_6012,N_849,N_1477);
or U6013 (N_6013,N_4329,N_2377);
nor U6014 (N_6014,N_4640,N_1372);
nand U6015 (N_6015,N_12,N_4610);
xnor U6016 (N_6016,N_3793,N_3418);
xnor U6017 (N_6017,N_527,N_4203);
nand U6018 (N_6018,N_1467,N_4230);
nor U6019 (N_6019,N_1435,N_647);
nor U6020 (N_6020,N_4723,N_4504);
nand U6021 (N_6021,N_2057,N_789);
nand U6022 (N_6022,N_316,N_260);
nor U6023 (N_6023,N_240,N_1573);
nor U6024 (N_6024,N_1411,N_3675);
nor U6025 (N_6025,N_4556,N_4496);
xor U6026 (N_6026,N_1174,N_1357);
nand U6027 (N_6027,N_4795,N_1428);
nor U6028 (N_6028,N_3246,N_4747);
or U6029 (N_6029,N_4458,N_3934);
and U6030 (N_6030,N_173,N_3723);
nand U6031 (N_6031,N_806,N_943);
xor U6032 (N_6032,N_4110,N_3631);
nand U6033 (N_6033,N_2683,N_1386);
xor U6034 (N_6034,N_90,N_921);
nand U6035 (N_6035,N_3948,N_4343);
nand U6036 (N_6036,N_1991,N_2922);
and U6037 (N_6037,N_3497,N_322);
or U6038 (N_6038,N_605,N_4449);
xor U6039 (N_6039,N_4840,N_1913);
nand U6040 (N_6040,N_1579,N_4265);
and U6041 (N_6041,N_3208,N_4358);
and U6042 (N_6042,N_1950,N_3187);
nand U6043 (N_6043,N_496,N_2563);
xor U6044 (N_6044,N_2873,N_1634);
and U6045 (N_6045,N_4318,N_4964);
or U6046 (N_6046,N_2211,N_610);
or U6047 (N_6047,N_1046,N_2387);
and U6048 (N_6048,N_3687,N_4831);
nand U6049 (N_6049,N_831,N_4934);
nor U6050 (N_6050,N_3885,N_1999);
nor U6051 (N_6051,N_3471,N_1075);
and U6052 (N_6052,N_1338,N_4365);
or U6053 (N_6053,N_1359,N_4499);
nand U6054 (N_6054,N_111,N_119);
nor U6055 (N_6055,N_3827,N_368);
and U6056 (N_6056,N_4809,N_106);
xnor U6057 (N_6057,N_2800,N_1117);
and U6058 (N_6058,N_4625,N_3005);
or U6059 (N_6059,N_2283,N_3363);
xor U6060 (N_6060,N_159,N_1487);
xor U6061 (N_6061,N_4404,N_2322);
or U6062 (N_6062,N_3381,N_3315);
and U6063 (N_6063,N_2738,N_196);
nor U6064 (N_6064,N_4452,N_4502);
and U6065 (N_6065,N_2174,N_3180);
nand U6066 (N_6066,N_4107,N_2511);
and U6067 (N_6067,N_1180,N_3139);
nor U6068 (N_6068,N_4619,N_4644);
nand U6069 (N_6069,N_1437,N_832);
and U6070 (N_6070,N_2568,N_4474);
xor U6071 (N_6071,N_1722,N_3382);
or U6072 (N_6072,N_3339,N_63);
nor U6073 (N_6073,N_2701,N_777);
xor U6074 (N_6074,N_2769,N_4134);
nor U6075 (N_6075,N_1236,N_2189);
or U6076 (N_6076,N_1658,N_335);
nor U6077 (N_6077,N_2698,N_1415);
or U6078 (N_6078,N_2329,N_3927);
xnor U6079 (N_6079,N_1760,N_2073);
and U6080 (N_6080,N_2919,N_2235);
nand U6081 (N_6081,N_1589,N_2016);
and U6082 (N_6082,N_4514,N_2868);
xnor U6083 (N_6083,N_3802,N_3334);
xor U6084 (N_6084,N_1061,N_4751);
and U6085 (N_6085,N_1509,N_4001);
or U6086 (N_6086,N_2017,N_4728);
nor U6087 (N_6087,N_3686,N_4172);
and U6088 (N_6088,N_3784,N_4154);
nand U6089 (N_6089,N_982,N_3084);
xor U6090 (N_6090,N_1426,N_543);
or U6091 (N_6091,N_903,N_1500);
nor U6092 (N_6092,N_4500,N_3090);
nor U6093 (N_6093,N_2237,N_2878);
and U6094 (N_6094,N_3670,N_3809);
and U6095 (N_6095,N_472,N_4415);
nand U6096 (N_6096,N_3268,N_4328);
xor U6097 (N_6097,N_4478,N_4669);
nor U6098 (N_6098,N_3312,N_2265);
nor U6099 (N_6099,N_4709,N_1619);
or U6100 (N_6100,N_1875,N_3257);
or U6101 (N_6101,N_3508,N_4974);
nand U6102 (N_6102,N_4562,N_895);
nand U6103 (N_6103,N_1597,N_2106);
nor U6104 (N_6104,N_4798,N_212);
xnor U6105 (N_6105,N_2006,N_36);
nor U6106 (N_6106,N_746,N_1552);
nand U6107 (N_6107,N_276,N_949);
nor U6108 (N_6108,N_2278,N_358);
or U6109 (N_6109,N_3577,N_2204);
xor U6110 (N_6110,N_507,N_2473);
and U6111 (N_6111,N_220,N_1883);
nand U6112 (N_6112,N_3372,N_4688);
or U6113 (N_6113,N_3228,N_1305);
or U6114 (N_6114,N_421,N_135);
and U6115 (N_6115,N_2436,N_2354);
or U6116 (N_6116,N_3141,N_4280);
xor U6117 (N_6117,N_429,N_2137);
nand U6118 (N_6118,N_4489,N_3043);
xor U6119 (N_6119,N_3776,N_4590);
nor U6120 (N_6120,N_1162,N_1244);
or U6121 (N_6121,N_3108,N_2812);
and U6122 (N_6122,N_1742,N_4238);
nor U6123 (N_6123,N_788,N_2496);
xor U6124 (N_6124,N_62,N_114);
nand U6125 (N_6125,N_4278,N_3117);
nor U6126 (N_6126,N_4796,N_483);
nand U6127 (N_6127,N_2779,N_2313);
xnor U6128 (N_6128,N_2520,N_4525);
and U6129 (N_6129,N_2190,N_2120);
nor U6130 (N_6130,N_2442,N_3575);
or U6131 (N_6131,N_1095,N_2491);
or U6132 (N_6132,N_4859,N_4205);
nand U6133 (N_6133,N_799,N_1503);
nand U6134 (N_6134,N_3193,N_3523);
or U6135 (N_6135,N_3436,N_1982);
and U6136 (N_6136,N_4858,N_2768);
or U6137 (N_6137,N_625,N_13);
and U6138 (N_6138,N_32,N_4300);
nand U6139 (N_6139,N_3633,N_2074);
nand U6140 (N_6140,N_160,N_3105);
and U6141 (N_6141,N_4354,N_187);
or U6142 (N_6142,N_3232,N_841);
and U6143 (N_6143,N_2695,N_4484);
nor U6144 (N_6144,N_450,N_3041);
or U6145 (N_6145,N_2147,N_915);
nor U6146 (N_6146,N_4208,N_582);
or U6147 (N_6147,N_1538,N_4122);
xor U6148 (N_6148,N_464,N_1717);
or U6149 (N_6149,N_4304,N_2094);
nand U6150 (N_6150,N_1832,N_3295);
and U6151 (N_6151,N_3330,N_1229);
or U6152 (N_6152,N_3154,N_3884);
and U6153 (N_6153,N_4680,N_916);
xor U6154 (N_6154,N_4724,N_1599);
or U6155 (N_6155,N_127,N_4439);
or U6156 (N_6156,N_3941,N_760);
nand U6157 (N_6157,N_1029,N_2854);
nand U6158 (N_6158,N_4951,N_692);
nand U6159 (N_6159,N_856,N_2474);
xnor U6160 (N_6160,N_4596,N_739);
or U6161 (N_6161,N_1704,N_2797);
nor U6162 (N_6162,N_3967,N_3428);
or U6163 (N_6163,N_2633,N_1959);
and U6164 (N_6164,N_4722,N_3490);
xnor U6165 (N_6165,N_3337,N_4587);
nand U6166 (N_6166,N_1060,N_3269);
nand U6167 (N_6167,N_2642,N_1093);
xnor U6168 (N_6168,N_2941,N_4865);
or U6169 (N_6169,N_4070,N_1936);
or U6170 (N_6170,N_4830,N_2415);
and U6171 (N_6171,N_3976,N_3085);
or U6172 (N_6172,N_49,N_2635);
xor U6173 (N_6173,N_344,N_3343);
nor U6174 (N_6174,N_946,N_2198);
or U6175 (N_6175,N_2743,N_595);
or U6176 (N_6176,N_2066,N_3624);
xnor U6177 (N_6177,N_556,N_2896);
nand U6178 (N_6178,N_910,N_2310);
and U6179 (N_6179,N_3903,N_1105);
xor U6180 (N_6180,N_4716,N_3824);
and U6181 (N_6181,N_398,N_4369);
nand U6182 (N_6182,N_1409,N_2187);
nand U6183 (N_6183,N_4306,N_3053);
nor U6184 (N_6184,N_1768,N_1205);
xor U6185 (N_6185,N_2389,N_1662);
xor U6186 (N_6186,N_2160,N_4077);
xor U6187 (N_6187,N_3663,N_1);
nor U6188 (N_6188,N_2874,N_349);
xnor U6189 (N_6189,N_4473,N_3313);
or U6190 (N_6190,N_3304,N_1339);
and U6191 (N_6191,N_1831,N_917);
nand U6192 (N_6192,N_616,N_1462);
nand U6193 (N_6193,N_1145,N_4822);
and U6194 (N_6194,N_57,N_4217);
or U6195 (N_6195,N_3960,N_4494);
and U6196 (N_6196,N_600,N_4235);
xor U6197 (N_6197,N_3275,N_2540);
xor U6198 (N_6198,N_1529,N_4894);
nand U6199 (N_6199,N_4501,N_4786);
nor U6200 (N_6200,N_3659,N_4374);
or U6201 (N_6201,N_4148,N_1525);
xor U6202 (N_6202,N_2838,N_4949);
xnor U6203 (N_6203,N_104,N_3597);
nor U6204 (N_6204,N_1748,N_3603);
nor U6205 (N_6205,N_4565,N_4874);
nand U6206 (N_6206,N_1540,N_1986);
and U6207 (N_6207,N_1856,N_1892);
nand U6208 (N_6208,N_1944,N_3383);
or U6209 (N_6209,N_1908,N_3455);
xnor U6210 (N_6210,N_1976,N_4579);
nand U6211 (N_6211,N_1453,N_1692);
xor U6212 (N_6212,N_4022,N_4614);
nor U6213 (N_6213,N_2441,N_2990);
or U6214 (N_6214,N_4192,N_3222);
or U6215 (N_6215,N_3702,N_4396);
and U6216 (N_6216,N_1227,N_4767);
or U6217 (N_6217,N_3764,N_2347);
or U6218 (N_6218,N_3801,N_2240);
xnor U6219 (N_6219,N_3510,N_331);
nand U6220 (N_6220,N_2572,N_367);
xor U6221 (N_6221,N_4785,N_1725);
nor U6222 (N_6222,N_3374,N_2739);
xor U6223 (N_6223,N_4541,N_241);
and U6224 (N_6224,N_1767,N_3456);
nor U6225 (N_6225,N_4375,N_4854);
or U6226 (N_6226,N_3213,N_699);
and U6227 (N_6227,N_3156,N_3788);
nor U6228 (N_6228,N_3588,N_2521);
xnor U6229 (N_6229,N_889,N_4754);
or U6230 (N_6230,N_4060,N_2363);
xor U6231 (N_6231,N_403,N_4791);
nand U6232 (N_6232,N_3340,N_2254);
nor U6233 (N_6233,N_2875,N_3019);
xnor U6234 (N_6234,N_1759,N_4123);
xor U6235 (N_6235,N_2973,N_3954);
and U6236 (N_6236,N_3042,N_3100);
nor U6237 (N_6237,N_1262,N_852);
xor U6238 (N_6238,N_1232,N_920);
nand U6239 (N_6239,N_3388,N_176);
or U6240 (N_6240,N_3198,N_2925);
and U6241 (N_6241,N_1265,N_280);
nor U6242 (N_6242,N_395,N_1535);
nand U6243 (N_6243,N_1001,N_2385);
and U6244 (N_6244,N_4685,N_161);
nand U6245 (N_6245,N_3611,N_2592);
nand U6246 (N_6246,N_4279,N_2421);
nor U6247 (N_6247,N_3057,N_2148);
or U6248 (N_6248,N_1283,N_675);
and U6249 (N_6249,N_437,N_291);
nor U6250 (N_6250,N_668,N_901);
xnor U6251 (N_6251,N_3778,N_773);
nor U6252 (N_6252,N_2827,N_4381);
nor U6253 (N_6253,N_4937,N_2244);
and U6254 (N_6254,N_2872,N_1946);
xor U6255 (N_6255,N_388,N_1508);
nand U6256 (N_6256,N_1550,N_3127);
or U6257 (N_6257,N_4018,N_3707);
nand U6258 (N_6258,N_2459,N_1323);
nor U6259 (N_6259,N_3104,N_1862);
nand U6260 (N_6260,N_816,N_1653);
nand U6261 (N_6261,N_1888,N_3756);
xnor U6262 (N_6262,N_1734,N_2949);
and U6263 (N_6263,N_17,N_3566);
nand U6264 (N_6264,N_811,N_2690);
xor U6265 (N_6265,N_2045,N_4143);
or U6266 (N_6266,N_1521,N_1651);
nor U6267 (N_6267,N_3717,N_754);
xnor U6268 (N_6268,N_460,N_377);
nor U6269 (N_6269,N_4264,N_4309);
or U6270 (N_6270,N_40,N_2565);
nor U6271 (N_6271,N_244,N_891);
or U6272 (N_6272,N_2426,N_2569);
or U6273 (N_6273,N_1903,N_4030);
and U6274 (N_6274,N_3327,N_2908);
and U6275 (N_6275,N_1728,N_3753);
xor U6276 (N_6276,N_3373,N_1099);
xor U6277 (N_6277,N_3331,N_418);
and U6278 (N_6278,N_1181,N_2804);
xnor U6279 (N_6279,N_2051,N_2611);
or U6280 (N_6280,N_1885,N_2067);
nor U6281 (N_6281,N_1520,N_4460);
and U6282 (N_6282,N_4506,N_2796);
nor U6283 (N_6283,N_2829,N_1945);
or U6284 (N_6284,N_3810,N_2044);
xnor U6285 (N_6285,N_1519,N_4289);
nor U6286 (N_6286,N_4823,N_3728);
nand U6287 (N_6287,N_4422,N_3024);
or U6288 (N_6288,N_2488,N_1266);
and U6289 (N_6289,N_1794,N_3484);
nand U6290 (N_6290,N_1135,N_2932);
xnor U6291 (N_6291,N_4424,N_2691);
and U6292 (N_6292,N_210,N_3875);
or U6293 (N_6293,N_2049,N_2821);
and U6294 (N_6294,N_3929,N_3431);
or U6295 (N_6295,N_2794,N_2438);
and U6296 (N_6296,N_3527,N_4308);
nor U6297 (N_6297,N_812,N_2468);
nand U6298 (N_6298,N_233,N_3452);
or U6299 (N_6299,N_994,N_4027);
xnor U6300 (N_6300,N_3639,N_3706);
or U6301 (N_6301,N_3983,N_4516);
xor U6302 (N_6302,N_3482,N_3651);
xnor U6303 (N_6303,N_2958,N_2010);
or U6304 (N_6304,N_3056,N_72);
nor U6305 (N_6305,N_4400,N_3399);
or U6306 (N_6306,N_2723,N_4583);
or U6307 (N_6307,N_1322,N_4243);
or U6308 (N_6308,N_3714,N_3729);
or U6309 (N_6309,N_2018,N_221);
nand U6310 (N_6310,N_1303,N_1961);
xnor U6311 (N_6311,N_3882,N_42);
xnor U6312 (N_6312,N_3685,N_1438);
nor U6313 (N_6313,N_1346,N_805);
nor U6314 (N_6314,N_855,N_3814);
or U6315 (N_6315,N_386,N_1416);
nor U6316 (N_6316,N_2448,N_28);
or U6317 (N_6317,N_4248,N_2331);
and U6318 (N_6318,N_3893,N_4550);
or U6319 (N_6319,N_950,N_1078);
or U6320 (N_6320,N_2307,N_2688);
nand U6321 (N_6321,N_4721,N_4333);
nor U6322 (N_6322,N_2965,N_2702);
nand U6323 (N_6323,N_466,N_320);
nand U6324 (N_6324,N_4233,N_1017);
or U6325 (N_6325,N_361,N_4889);
xnor U6326 (N_6326,N_1940,N_3607);
nand U6327 (N_6327,N_4373,N_606);
and U6328 (N_6328,N_888,N_2609);
or U6329 (N_6329,N_1864,N_3817);
and U6330 (N_6330,N_4390,N_3081);
nor U6331 (N_6331,N_2573,N_2815);
and U6332 (N_6332,N_566,N_1449);
and U6333 (N_6333,N_2171,N_1910);
and U6334 (N_6334,N_1035,N_3938);
nand U6335 (N_6335,N_2810,N_1703);
nand U6336 (N_6336,N_271,N_698);
nand U6337 (N_6337,N_3883,N_4671);
nor U6338 (N_6338,N_1307,N_3863);
or U6339 (N_6339,N_863,N_2192);
and U6340 (N_6340,N_422,N_43);
nand U6341 (N_6341,N_3474,N_1021);
and U6342 (N_6342,N_4973,N_2294);
nand U6343 (N_6343,N_1119,N_2193);
or U6344 (N_6344,N_3595,N_3211);
nor U6345 (N_6345,N_1582,N_4448);
nand U6346 (N_6346,N_2381,N_4544);
or U6347 (N_6347,N_1140,N_1980);
xor U6348 (N_6348,N_862,N_712);
nand U6349 (N_6349,N_3253,N_3427);
xnor U6350 (N_6350,N_2934,N_4342);
nand U6351 (N_6351,N_2071,N_4518);
or U6352 (N_6352,N_4960,N_4683);
or U6353 (N_6353,N_2399,N_3142);
or U6354 (N_6354,N_573,N_3329);
xnor U6355 (N_6355,N_3804,N_3791);
nand U6356 (N_6356,N_1894,N_3029);
xnor U6357 (N_6357,N_3467,N_4805);
or U6358 (N_6358,N_1163,N_3223);
or U6359 (N_6359,N_1067,N_834);
nand U6360 (N_6360,N_2904,N_3808);
xor U6361 (N_6361,N_4720,N_4174);
or U6362 (N_6362,N_4055,N_2803);
and U6363 (N_6363,N_3796,N_3170);
and U6364 (N_6364,N_1417,N_637);
and U6365 (N_6365,N_2566,N_180);
and U6366 (N_6366,N_2130,N_53);
and U6367 (N_6367,N_604,N_1439);
or U6368 (N_6368,N_2396,N_3873);
xor U6369 (N_6369,N_126,N_2798);
and U6370 (N_6370,N_2364,N_3578);
and U6371 (N_6371,N_469,N_3558);
and U6372 (N_6372,N_801,N_2176);
nor U6373 (N_6373,N_4214,N_2652);
nand U6374 (N_6374,N_3489,N_2731);
and U6375 (N_6375,N_4155,N_3975);
and U6376 (N_6376,N_665,N_2508);
or U6377 (N_6377,N_1390,N_1559);
xnor U6378 (N_6378,N_4521,N_3219);
nand U6379 (N_6379,N_463,N_500);
nand U6380 (N_6380,N_2601,N_3243);
nand U6381 (N_6381,N_308,N_334);
or U6382 (N_6382,N_256,N_4768);
and U6383 (N_6383,N_4465,N_4998);
or U6384 (N_6384,N_2403,N_1361);
nand U6385 (N_6385,N_3930,N_96);
xnor U6386 (N_6386,N_4515,N_563);
and U6387 (N_6387,N_2001,N_3722);
nor U6388 (N_6388,N_1650,N_1931);
and U6389 (N_6389,N_3276,N_103);
nor U6390 (N_6390,N_3751,N_204);
nor U6391 (N_6391,N_1838,N_2457);
and U6392 (N_6392,N_1539,N_1289);
or U6393 (N_6393,N_4825,N_2382);
or U6394 (N_6394,N_1123,N_858);
nand U6395 (N_6395,N_1611,N_2697);
nand U6396 (N_6396,N_1092,N_4730);
xnor U6397 (N_6397,N_987,N_2763);
xnor U6398 (N_6398,N_1572,N_4322);
nand U6399 (N_6399,N_4095,N_3730);
xor U6400 (N_6400,N_1355,N_957);
nand U6401 (N_6401,N_1247,N_376);
or U6402 (N_6402,N_2223,N_3902);
nor U6403 (N_6403,N_1039,N_3862);
nand U6404 (N_6404,N_1737,N_4986);
nand U6405 (N_6405,N_1661,N_3834);
and U6406 (N_6406,N_986,N_2677);
nand U6407 (N_6407,N_598,N_2778);
and U6408 (N_6408,N_3522,N_3661);
nor U6409 (N_6409,N_4731,N_569);
nor U6410 (N_6410,N_953,N_1795);
nand U6411 (N_6411,N_2987,N_2268);
or U6412 (N_6412,N_4481,N_4526);
nand U6413 (N_6413,N_4851,N_1321);
xor U6414 (N_6414,N_2862,N_3031);
and U6415 (N_6415,N_360,N_1444);
xnor U6416 (N_6416,N_4207,N_2117);
xor U6417 (N_6417,N_3394,N_129);
nor U6418 (N_6418,N_4537,N_2184);
nor U6419 (N_6419,N_3279,N_1000);
nand U6420 (N_6420,N_2924,N_3308);
or U6421 (N_6421,N_659,N_4096);
and U6422 (N_6422,N_4194,N_3544);
nand U6423 (N_6423,N_1176,N_1947);
xor U6424 (N_6424,N_1148,N_2348);
and U6425 (N_6425,N_4250,N_1257);
xnor U6426 (N_6426,N_2735,N_3293);
or U6427 (N_6427,N_2956,N_372);
nor U6428 (N_6428,N_4833,N_3999);
xnor U6429 (N_6429,N_2487,N_2783);
xnor U6430 (N_6430,N_3939,N_4169);
nor U6431 (N_6431,N_1146,N_1221);
xor U6432 (N_6432,N_3859,N_1517);
and U6433 (N_6433,N_3416,N_1546);
nor U6434 (N_6434,N_2341,N_565);
nor U6435 (N_6435,N_2980,N_3481);
nor U6436 (N_6436,N_3408,N_68);
xor U6437 (N_6437,N_4532,N_3958);
nand U6438 (N_6438,N_1147,N_479);
or U6439 (N_6439,N_1110,N_339);
nor U6440 (N_6440,N_3375,N_1834);
and U6441 (N_6441,N_3754,N_3725);
and U6442 (N_6442,N_3901,N_3367);
nand U6443 (N_6443,N_4380,N_2526);
nand U6444 (N_6444,N_4406,N_3857);
and U6445 (N_6445,N_3506,N_231);
and U6446 (N_6446,N_4297,N_3673);
xor U6447 (N_6447,N_1502,N_3314);
and U6448 (N_6448,N_4689,N_3640);
or U6449 (N_6449,N_1062,N_396);
nand U6450 (N_6450,N_706,N_902);
nand U6451 (N_6451,N_1729,N_2369);
and U6452 (N_6452,N_1952,N_3097);
or U6453 (N_6453,N_2651,N_989);
xnor U6454 (N_6454,N_2259,N_4622);
nand U6455 (N_6455,N_2963,N_2021);
xnor U6456 (N_6456,N_871,N_1253);
nor U6457 (N_6457,N_2851,N_513);
nor U6458 (N_6458,N_1434,N_1378);
nor U6459 (N_6459,N_3054,N_1626);
nor U6460 (N_6460,N_1738,N_1739);
nor U6461 (N_6461,N_3549,N_3377);
and U6462 (N_6462,N_1125,N_4114);
nand U6463 (N_6463,N_515,N_1780);
xor U6464 (N_6464,N_3747,N_4091);
xor U6465 (N_6465,N_2834,N_2730);
or U6466 (N_6466,N_1465,N_714);
and U6467 (N_6467,N_4423,N_3512);
xor U6468 (N_6468,N_4950,N_3668);
nand U6469 (N_6469,N_924,N_1367);
and U6470 (N_6470,N_2836,N_697);
and U6471 (N_6471,N_1019,N_4697);
xnor U6472 (N_6472,N_4635,N_201);
or U6473 (N_6473,N_1137,N_4441);
nand U6474 (N_6474,N_1098,N_4273);
nand U6475 (N_6475,N_3251,N_1312);
nor U6476 (N_6476,N_2047,N_4003);
nand U6477 (N_6477,N_2801,N_304);
nor U6478 (N_6478,N_528,N_4360);
nor U6479 (N_6479,N_1219,N_1049);
nand U6480 (N_6480,N_1226,N_3816);
nand U6481 (N_6481,N_1676,N_3609);
and U6482 (N_6482,N_4113,N_1992);
xor U6483 (N_6483,N_3103,N_682);
or U6484 (N_6484,N_3058,N_1869);
and U6485 (N_6485,N_402,N_251);
nand U6486 (N_6486,N_1699,N_298);
nand U6487 (N_6487,N_3320,N_1978);
nor U6488 (N_6488,N_554,N_4634);
or U6489 (N_6489,N_1397,N_1006);
or U6490 (N_6490,N_3248,N_4862);
nor U6491 (N_6491,N_2019,N_4538);
and U6492 (N_6492,N_1139,N_491);
or U6493 (N_6493,N_4729,N_3417);
and U6494 (N_6494,N_2831,N_3693);
xor U6495 (N_6495,N_3556,N_3028);
and U6496 (N_6496,N_109,N_4063);
nand U6497 (N_6497,N_1144,N_1179);
or U6498 (N_6498,N_536,N_3487);
nand U6499 (N_6499,N_2232,N_1973);
and U6500 (N_6500,N_1769,N_2839);
and U6501 (N_6501,N_3065,N_3171);
and U6502 (N_6502,N_2481,N_2405);
nor U6503 (N_6503,N_3935,N_557);
xor U6504 (N_6504,N_423,N_1736);
or U6505 (N_6505,N_3709,N_3587);
nor U6506 (N_6506,N_1498,N_4632);
or U6507 (N_6507,N_4836,N_2115);
nand U6508 (N_6508,N_2618,N_2456);
and U6509 (N_6509,N_4659,N_1628);
and U6510 (N_6510,N_1826,N_3559);
nor U6511 (N_6511,N_3660,N_332);
and U6512 (N_6512,N_4146,N_425);
nor U6513 (N_6513,N_428,N_3178);
xnor U6514 (N_6514,N_2394,N_4816);
xor U6515 (N_6515,N_3984,N_2964);
or U6516 (N_6516,N_3021,N_2312);
or U6517 (N_6517,N_2435,N_2708);
nand U6518 (N_6518,N_2165,N_1575);
xnor U6519 (N_6519,N_2069,N_4529);
or U6520 (N_6520,N_1329,N_2863);
or U6521 (N_6521,N_1911,N_2817);
nor U6522 (N_6522,N_1203,N_181);
xor U6523 (N_6523,N_297,N_1299);
or U6524 (N_6524,N_1217,N_4438);
xor U6525 (N_6525,N_1691,N_1480);
nand U6526 (N_6526,N_3785,N_1210);
nand U6527 (N_6527,N_4274,N_3704);
xor U6528 (N_6528,N_1310,N_270);
xor U6529 (N_6529,N_3807,N_79);
and U6530 (N_6530,N_4456,N_2210);
or U6531 (N_6531,N_3344,N_4080);
and U6532 (N_6532,N_3121,N_2477);
nand U6533 (N_6533,N_4597,N_971);
or U6534 (N_6534,N_887,N_198);
nor U6535 (N_6535,N_3565,N_1621);
and U6536 (N_6536,N_3744,N_3543);
and U6537 (N_6537,N_2273,N_1012);
and U6538 (N_6538,N_4755,N_3155);
and U6539 (N_6539,N_4761,N_1727);
xor U6540 (N_6540,N_815,N_4790);
or U6541 (N_6541,N_4219,N_762);
or U6542 (N_6542,N_3654,N_717);
and U6543 (N_6543,N_1189,N_411);
nor U6544 (N_6544,N_3409,N_3277);
nor U6545 (N_6545,N_1827,N_3993);
or U6546 (N_6546,N_2679,N_1590);
xor U6547 (N_6547,N_1454,N_1987);
or U6548 (N_6548,N_4876,N_3550);
nand U6549 (N_6549,N_3823,N_468);
xor U6550 (N_6550,N_1055,N_3133);
xor U6551 (N_6551,N_4869,N_3406);
xor U6552 (N_6552,N_3302,N_3569);
nand U6553 (N_6553,N_1878,N_3470);
xnor U6554 (N_6554,N_2,N_1268);
or U6555 (N_6555,N_3411,N_1413);
and U6556 (N_6556,N_3689,N_4654);
or U6557 (N_6557,N_4899,N_3356);
nor U6558 (N_6558,N_4984,N_2860);
nand U6559 (N_6559,N_3082,N_1732);
nor U6560 (N_6560,N_2249,N_436);
and U6561 (N_6561,N_884,N_3630);
and U6562 (N_6562,N_4552,N_2319);
nand U6563 (N_6563,N_3378,N_3335);
xnor U6564 (N_6564,N_1436,N_1334);
nor U6565 (N_6565,N_2201,N_2085);
and U6566 (N_6566,N_4436,N_814);
xor U6567 (N_6567,N_2968,N_4181);
and U6568 (N_6568,N_4257,N_1456);
or U6569 (N_6569,N_4432,N_3458);
and U6570 (N_6570,N_4000,N_52);
and U6571 (N_6571,N_3488,N_3434);
nor U6572 (N_6572,N_2038,N_4371);
nand U6573 (N_6573,N_4690,N_3203);
xor U6574 (N_6574,N_4996,N_684);
or U6575 (N_6575,N_3546,N_4781);
or U6576 (N_6576,N_4236,N_2936);
and U6577 (N_6577,N_415,N_4624);
nand U6578 (N_6578,N_2177,N_3763);
or U6579 (N_6579,N_1598,N_1631);
and U6580 (N_6580,N_2227,N_4298);
and U6581 (N_6581,N_2658,N_4838);
nor U6582 (N_6582,N_2123,N_2629);
and U6583 (N_6583,N_4367,N_69);
and U6584 (N_6584,N_4922,N_4763);
xor U6585 (N_6585,N_4846,N_4009);
nand U6586 (N_6586,N_3755,N_3209);
nor U6587 (N_6587,N_4533,N_2040);
nand U6588 (N_6588,N_3240,N_4820);
nor U6589 (N_6589,N_3419,N_4563);
nand U6590 (N_6590,N_1327,N_2358);
or U6591 (N_6591,N_2746,N_865);
xor U6592 (N_6592,N_2948,N_137);
xnor U6593 (N_6593,N_4216,N_937);
nand U6594 (N_6594,N_540,N_218);
and U6595 (N_6595,N_3425,N_3235);
nand U6596 (N_6596,N_1309,N_1492);
nor U6597 (N_6597,N_914,N_2705);
nor U6598 (N_6598,N_3612,N_4366);
or U6599 (N_6599,N_3352,N_807);
xor U6600 (N_6600,N_2243,N_3835);
or U6601 (N_6601,N_352,N_2248);
and U6602 (N_6602,N_4978,N_1482);
xnor U6603 (N_6603,N_826,N_1694);
or U6604 (N_6604,N_1716,N_596);
and U6605 (N_6605,N_4498,N_2921);
nand U6606 (N_6606,N_3422,N_2614);
nor U6607 (N_6607,N_1160,N_2923);
nor U6608 (N_6608,N_4627,N_1859);
xor U6609 (N_6609,N_3879,N_4453);
xor U6610 (N_6610,N_2388,N_3667);
and U6611 (N_6611,N_2607,N_3259);
or U6612 (N_6612,N_4551,N_1089);
and U6613 (N_6613,N_4350,N_2196);
xor U6614 (N_6614,N_776,N_1744);
or U6615 (N_6615,N_182,N_4687);
and U6616 (N_6616,N_4752,N_4961);
nor U6617 (N_6617,N_427,N_2214);
nand U6618 (N_6618,N_3531,N_677);
or U6619 (N_6619,N_1079,N_693);
or U6620 (N_6620,N_3038,N_1633);
xnor U6621 (N_6621,N_3618,N_1506);
and U6622 (N_6622,N_223,N_363);
or U6623 (N_6623,N_900,N_3843);
nand U6624 (N_6624,N_379,N_48);
nand U6625 (N_6625,N_780,N_4826);
nand U6626 (N_6626,N_4997,N_3384);
xnor U6627 (N_6627,N_3600,N_2305);
xor U6628 (N_6628,N_2345,N_2308);
and U6629 (N_6629,N_105,N_3283);
nor U6630 (N_6630,N_4412,N_3634);
or U6631 (N_6631,N_1081,N_1967);
xnor U6632 (N_6632,N_3018,N_4800);
xor U6633 (N_6633,N_580,N_632);
or U6634 (N_6634,N_4157,N_4631);
nor U6635 (N_6635,N_4056,N_237);
xor U6636 (N_6636,N_1654,N_4657);
or U6637 (N_6637,N_3529,N_1735);
or U6638 (N_6638,N_3644,N_2271);
nand U6639 (N_6639,N_2982,N_3623);
and U6640 (N_6640,N_1710,N_3855);
and U6641 (N_6641,N_650,N_3309);
or U6642 (N_6642,N_2825,N_508);
nor U6643 (N_6643,N_338,N_761);
xor U6644 (N_6644,N_124,N_3101);
nor U6645 (N_6645,N_945,N_257);
nand U6646 (N_6646,N_3010,N_1165);
nand U6647 (N_6647,N_3396,N_1874);
nor U6648 (N_6648,N_4670,N_3048);
or U6649 (N_6649,N_4936,N_2286);
or U6650 (N_6650,N_599,N_4611);
and U6651 (N_6651,N_1382,N_1073);
and U6652 (N_6652,N_283,N_1332);
and U6653 (N_6653,N_662,N_353);
or U6654 (N_6654,N_766,N_475);
or U6655 (N_6655,N_1231,N_4736);
or U6656 (N_6656,N_3175,N_3196);
nand U6657 (N_6657,N_3354,N_1004);
nor U6658 (N_6658,N_727,N_380);
nand U6659 (N_6659,N_931,N_3003);
or U6660 (N_6660,N_1340,N_4270);
or U6661 (N_6661,N_2129,N_1754);
nand U6662 (N_6662,N_2316,N_3845);
nand U6663 (N_6663,N_743,N_1778);
nor U6664 (N_6664,N_2112,N_704);
xnor U6665 (N_6665,N_2103,N_3262);
nand U6666 (N_6666,N_4130,N_134);
xnor U6667 (N_6667,N_2882,N_3910);
and U6668 (N_6668,N_2888,N_784);
xor U6669 (N_6669,N_33,N_1396);
and U6670 (N_6670,N_2883,N_1995);
nor U6671 (N_6671,N_1551,N_3719);
or U6672 (N_6672,N_700,N_4089);
nand U6673 (N_6673,N_1045,N_4992);
nand U6674 (N_6674,N_3571,N_3075);
and U6675 (N_6675,N_151,N_3271);
or U6676 (N_6676,N_3738,N_835);
and U6677 (N_6677,N_1238,N_190);
nand U6678 (N_6678,N_1664,N_3391);
nor U6679 (N_6679,N_3638,N_3346);
or U6680 (N_6680,N_4150,N_1250);
xnor U6681 (N_6681,N_833,N_4698);
nor U6682 (N_6682,N_628,N_3216);
nand U6683 (N_6683,N_290,N_1475);
nand U6684 (N_6684,N_2715,N_846);
or U6685 (N_6685,N_4667,N_3821);
nor U6686 (N_6686,N_3432,N_4180);
xnor U6687 (N_6687,N_3825,N_1200);
nor U6688 (N_6688,N_850,N_1106);
xnor U6689 (N_6689,N_857,N_4017);
nand U6690 (N_6690,N_3023,N_904);
xnor U6691 (N_6691,N_963,N_4125);
xnor U6692 (N_6692,N_4064,N_4081);
xor U6693 (N_6693,N_996,N_4085);
and U6694 (N_6694,N_2640,N_2054);
nor U6695 (N_6695,N_2784,N_171);
xnor U6696 (N_6696,N_1609,N_3439);
or U6697 (N_6697,N_2146,N_726);
nor U6698 (N_6698,N_1975,N_1172);
nor U6699 (N_6699,N_2169,N_4918);
or U6700 (N_6700,N_1670,N_3093);
xor U6701 (N_6701,N_2579,N_4819);
or U6702 (N_6702,N_2895,N_2805);
nand U6703 (N_6703,N_1274,N_4748);
and U6704 (N_6704,N_2152,N_2229);
nor U6705 (N_6705,N_2832,N_285);
and U6706 (N_6706,N_2970,N_4668);
or U6707 (N_6707,N_4555,N_1185);
nor U6708 (N_6708,N_1686,N_1514);
nor U6709 (N_6709,N_1770,N_3179);
nand U6710 (N_6710,N_661,N_263);
or U6711 (N_6711,N_1171,N_118);
nand U6712 (N_6712,N_4604,N_2728);
xnor U6713 (N_6713,N_511,N_24);
xnor U6714 (N_6714,N_3554,N_2528);
or U6715 (N_6715,N_3850,N_4783);
nand U6716 (N_6716,N_1197,N_2657);
xor U6717 (N_6717,N_307,N_2390);
nand U6718 (N_6718,N_140,N_2427);
or U6719 (N_6719,N_1330,N_4286);
nand U6720 (N_6720,N_2090,N_3448);
or U6721 (N_6721,N_3583,N_2646);
or U6722 (N_6722,N_2469,N_4330);
or U6723 (N_6723,N_1781,N_2246);
or U6724 (N_6724,N_896,N_2660);
xor U6725 (N_6725,N_3584,N_1607);
nand U6726 (N_6726,N_4476,N_4059);
and U6727 (N_6727,N_20,N_1900);
or U6728 (N_6728,N_4591,N_1858);
xor U6729 (N_6729,N_3555,N_735);
nand U6730 (N_6730,N_3589,N_4078);
and U6731 (N_6731,N_3395,N_3265);
or U6732 (N_6732,N_2323,N_3844);
or U6733 (N_6733,N_1047,N_2909);
or U6734 (N_6734,N_2813,N_3001);
nor U6735 (N_6735,N_2384,N_2099);
nand U6736 (N_6736,N_765,N_1750);
nor U6737 (N_6737,N_2470,N_4419);
xnor U6738 (N_6738,N_4083,N_3201);
or U6739 (N_6739,N_206,N_4188);
xnor U6740 (N_6740,N_4331,N_197);
nand U6741 (N_6741,N_4608,N_4394);
and U6742 (N_6742,N_148,N_1394);
or U6743 (N_6743,N_4988,N_2055);
nand U6744 (N_6744,N_3404,N_1104);
xor U6745 (N_6745,N_2927,N_1044);
xor U6746 (N_6746,N_2502,N_2939);
and U6747 (N_6747,N_4524,N_685);
and U6748 (N_6748,N_2946,N_3473);
nand U6749 (N_6749,N_274,N_2145);
xor U6750 (N_6750,N_919,N_2203);
nand U6751 (N_6751,N_470,N_2625);
nor U6752 (N_6752,N_4104,N_3113);
and U6753 (N_6753,N_3895,N_498);
nand U6754 (N_6754,N_265,N_29);
nor U6755 (N_6755,N_2199,N_3780);
nor U6756 (N_6756,N_3838,N_3557);
nor U6757 (N_6757,N_1455,N_2449);
xnor U6758 (N_6758,N_2476,N_2031);
xnor U6759 (N_6759,N_3533,N_758);
and U6760 (N_6760,N_175,N_1928);
nor U6761 (N_6761,N_1068,N_2859);
nand U6762 (N_6762,N_4725,N_4985);
xnor U6763 (N_6763,N_4963,N_2096);
or U6764 (N_6764,N_3138,N_1851);
xnor U6765 (N_6765,N_1028,N_686);
nand U6766 (N_6766,N_1263,N_3420);
nor U6767 (N_6767,N_3519,N_2737);
nor U6768 (N_6768,N_529,N_3812);
nand U6769 (N_6769,N_1636,N_3568);
nor U6770 (N_6770,N_4430,N_4469);
xnor U6771 (N_6771,N_1645,N_785);
and U6772 (N_6772,N_311,N_2097);
and U6773 (N_6773,N_1804,N_4749);
nand U6774 (N_6774,N_2951,N_2230);
and U6775 (N_6775,N_27,N_1280);
nor U6776 (N_6776,N_1132,N_1663);
and U6777 (N_6777,N_2222,N_4599);
nand U6778 (N_6778,N_2334,N_2585);
or U6779 (N_6779,N_872,N_2200);
nand U6780 (N_6780,N_4623,N_4133);
nand U6781 (N_6781,N_4321,N_3765);
xnor U6782 (N_6782,N_4340,N_4902);
nor U6783 (N_6783,N_1188,N_4895);
and U6784 (N_6784,N_128,N_4981);
nor U6785 (N_6785,N_1054,N_254);
xor U6786 (N_6786,N_3635,N_2649);
and U6787 (N_6787,N_1765,N_4815);
nand U6788 (N_6788,N_4462,N_4975);
nand U6789 (N_6789,N_4413,N_3869);
xnor U6790 (N_6790,N_3994,N_4701);
nor U6791 (N_6791,N_4793,N_926);
or U6792 (N_6792,N_2893,N_4229);
xor U6793 (N_6793,N_905,N_4445);
xor U6794 (N_6794,N_584,N_484);
xor U6795 (N_6795,N_120,N_3799);
xor U6796 (N_6796,N_3205,N_2844);
and U6797 (N_6797,N_4777,N_4386);
and U6798 (N_6798,N_2855,N_4457);
nor U6799 (N_6799,N_3286,N_2647);
nor U6800 (N_6800,N_546,N_3978);
nor U6801 (N_6801,N_3832,N_640);
nand U6802 (N_6802,N_3002,N_1256);
nand U6803 (N_6803,N_3407,N_66);
or U6804 (N_6804,N_3410,N_4886);
or U6805 (N_6805,N_4661,N_2693);
or U6806 (N_6806,N_150,N_1187);
xnor U6807 (N_6807,N_177,N_2352);
and U6808 (N_6808,N_3496,N_139);
nor U6809 (N_6809,N_1983,N_155);
nand U6810 (N_6810,N_282,N_1373);
nand U6811 (N_6811,N_3088,N_4475);
nor U6812 (N_6812,N_2365,N_4377);
nor U6813 (N_6813,N_4511,N_3400);
nor U6814 (N_6814,N_3370,N_4427);
and U6815 (N_6815,N_88,N_721);
and U6816 (N_6816,N_1771,N_715);
or U6817 (N_6817,N_229,N_2562);
and U6818 (N_6818,N_1239,N_4977);
nor U6819 (N_6819,N_2041,N_10);
nor U6820 (N_6820,N_3537,N_486);
nand U6821 (N_6821,N_305,N_2128);
xnor U6822 (N_6822,N_1776,N_1195);
nand U6823 (N_6823,N_1421,N_2371);
nor U6824 (N_6824,N_4574,N_964);
nand U6825 (N_6825,N_1202,N_4128);
nand U6826 (N_6826,N_1406,N_2191);
or U6827 (N_6827,N_3230,N_838);
nand U6828 (N_6828,N_813,N_1214);
xor U6829 (N_6829,N_1072,N_217);
xnor U6830 (N_6830,N_4490,N_2624);
and U6831 (N_6831,N_749,N_4065);
xnor U6832 (N_6832,N_1799,N_3173);
or U6833 (N_6833,N_4428,N_222);
xnor U6834 (N_6834,N_2971,N_2209);
and U6835 (N_6835,N_3020,N_2297);
nor U6836 (N_6836,N_3109,N_4536);
and U6837 (N_6837,N_2113,N_1293);
nor U6838 (N_6838,N_4076,N_3502);
or U6839 (N_6839,N_1527,N_1156);
xnor U6840 (N_6840,N_501,N_3628);
and U6841 (N_6841,N_2079,N_1043);
nand U6842 (N_6842,N_1536,N_3822);
xor U6843 (N_6843,N_1167,N_3060);
nand U6844 (N_6844,N_4414,N_4206);
and U6845 (N_6845,N_4244,N_4368);
or U6846 (N_6846,N_4231,N_588);
nor U6847 (N_6847,N_4648,N_1865);
nand U6848 (N_6848,N_480,N_3433);
nand U6849 (N_6849,N_1701,N_1169);
and U6850 (N_6850,N_1481,N_1153);
nor U6851 (N_6851,N_3572,N_1158);
or U6852 (N_6852,N_4170,N_4158);
nor U6853 (N_6853,N_4717,N_4813);
xor U6854 (N_6854,N_385,N_984);
nor U6855 (N_6855,N_3792,N_2173);
or U6856 (N_6856,N_2012,N_3783);
nor U6857 (N_6857,N_130,N_3671);
and U6858 (N_6858,N_643,N_1682);
nor U6859 (N_6859,N_1904,N_2507);
or U6860 (N_6860,N_2689,N_2857);
and U6861 (N_6861,N_2527,N_3899);
nand U6862 (N_6862,N_824,N_4999);
and U6863 (N_6863,N_2711,N_2463);
nand U6864 (N_6864,N_4284,N_4979);
or U6865 (N_6865,N_3319,N_2499);
nor U6866 (N_6866,N_2752,N_2140);
or U6867 (N_6867,N_4738,N_4991);
nand U6868 (N_6868,N_1687,N_2668);
nand U6869 (N_6869,N_2613,N_2361);
xor U6870 (N_6870,N_375,N_2891);
and U6871 (N_6871,N_899,N_369);
nand U6872 (N_6872,N_751,N_4339);
nor U6873 (N_6873,N_293,N_3055);
or U6874 (N_6874,N_4190,N_1898);
and U6875 (N_6875,N_4775,N_3579);
nor U6876 (N_6876,N_790,N_578);
and U6877 (N_6877,N_2136,N_1814);
xor U6878 (N_6878,N_3349,N_2644);
nor U6879 (N_6879,N_1121,N_4291);
nor U6880 (N_6880,N_1152,N_3068);
or U6881 (N_6881,N_820,N_337);
and U6882 (N_6882,N_4930,N_1588);
nand U6883 (N_6883,N_3163,N_3534);
nand U6884 (N_6884,N_209,N_1807);
xnor U6885 (N_6885,N_301,N_4857);
nand U6886 (N_6886,N_854,N_7);
and U6887 (N_6887,N_4535,N_2185);
and U6888 (N_6888,N_639,N_2315);
xnor U6889 (N_6889,N_4880,N_2118);
and U6890 (N_6890,N_3715,N_2030);
and U6891 (N_6891,N_4254,N_3700);
nand U6892 (N_6892,N_2236,N_516);
and U6893 (N_6893,N_4784,N_1345);
or U6894 (N_6894,N_138,N_3877);
nand U6895 (N_6895,N_303,N_4879);
or U6896 (N_6896,N_4586,N_609);
or U6897 (N_6897,N_3881,N_4694);
nand U6898 (N_6898,N_3074,N_154);
xnor U6899 (N_6899,N_3450,N_447);
nand U6900 (N_6900,N_2576,N_1175);
and U6901 (N_6901,N_1530,N_1366);
nand U6902 (N_6902,N_4124,N_3761);
or U6903 (N_6903,N_4821,N_4971);
xor U6904 (N_6904,N_623,N_1254);
nor U6905 (N_6905,N_1714,N_1424);
xnor U6906 (N_6906,N_1951,N_3620);
nor U6907 (N_6907,N_742,N_2753);
xnor U6908 (N_6908,N_2327,N_531);
or U6909 (N_6909,N_188,N_287);
xor U6910 (N_6910,N_4010,N_2195);
xor U6911 (N_6911,N_3683,N_541);
and U6912 (N_6912,N_272,N_520);
and U6913 (N_6913,N_2343,N_4290);
and U6914 (N_6914,N_1522,N_2291);
and U6915 (N_6915,N_1923,N_3547);
nor U6916 (N_6916,N_2258,N_535);
or U6917 (N_6917,N_178,N_4247);
xnor U6918 (N_6918,N_505,N_3629);
xor U6919 (N_6919,N_2577,N_1627);
or U6920 (N_6920,N_1260,N_4952);
and U6921 (N_6921,N_4843,N_669);
xor U6922 (N_6922,N_3250,N_663);
nor U6923 (N_6923,N_1775,N_3853);
nand U6924 (N_6924,N_3734,N_2061);
or U6925 (N_6925,N_107,N_2231);
and U6926 (N_6926,N_3819,N_286);
xor U6927 (N_6927,N_211,N_4140);
or U6928 (N_6928,N_552,N_575);
nor U6929 (N_6929,N_730,N_355);
nand U6930 (N_6930,N_3562,N_1377);
and U6931 (N_6931,N_2515,N_2004);
xor U6932 (N_6932,N_691,N_4837);
nand U6933 (N_6933,N_1709,N_4636);
xor U6934 (N_6934,N_1389,N_4171);
and U6935 (N_6935,N_4812,N_4327);
and U6936 (N_6936,N_4446,N_1915);
nand U6937 (N_6937,N_3321,N_542);
xnor U6938 (N_6938,N_441,N_2398);
and U6939 (N_6939,N_1659,N_4923);
nand U6940 (N_6940,N_4197,N_4129);
xor U6941 (N_6941,N_3767,N_4969);
and U6942 (N_6942,N_2638,N_2215);
nor U6943 (N_6943,N_3027,N_827);
and U6944 (N_6944,N_4684,N_694);
and U6945 (N_6945,N_2420,N_2325);
or U6946 (N_6946,N_288,N_4356);
nor U6947 (N_6947,N_1129,N_1328);
or U6948 (N_6948,N_3736,N_933);
or U6949 (N_6949,N_1984,N_2889);
xnor U6950 (N_6950,N_1122,N_1688);
xnor U6951 (N_6951,N_4103,N_179);
or U6952 (N_6952,N_3797,N_3280);
nor U6953 (N_6953,N_4268,N_1916);
and U6954 (N_6954,N_247,N_3805);
and U6955 (N_6955,N_4681,N_981);
xor U6956 (N_6956,N_911,N_4054);
or U6957 (N_6957,N_414,N_1548);
nor U6958 (N_6958,N_3475,N_2567);
nor U6959 (N_6959,N_4068,N_4847);
nor U6960 (N_6960,N_1806,N_2894);
and U6961 (N_6961,N_3971,N_3096);
nand U6962 (N_6962,N_4773,N_4808);
and U6963 (N_6963,N_2412,N_0);
xor U6964 (N_6964,N_1504,N_2219);
nor U6965 (N_6965,N_4344,N_622);
and U6966 (N_6966,N_74,N_2663);
and U6967 (N_6967,N_533,N_2799);
nand U6968 (N_6968,N_440,N_3118);
xor U6969 (N_6969,N_370,N_2393);
nand U6970 (N_6970,N_2906,N_3956);
nand U6971 (N_6971,N_844,N_3829);
nor U6972 (N_6972,N_3561,N_3443);
or U6973 (N_6973,N_3711,N_3945);
xnor U6974 (N_6974,N_1786,N_3292);
nor U6975 (N_6975,N_4940,N_503);
nand U6976 (N_6976,N_3324,N_1990);
and U6977 (N_6977,N_3904,N_3970);
nor U6978 (N_6978,N_2467,N_848);
xor U6979 (N_6979,N_2015,N_4361);
nand U6980 (N_6980,N_759,N_4418);
or U6981 (N_6981,N_4098,N_4126);
and U6982 (N_6982,N_4665,N_2986);
nand U6983 (N_6983,N_2953,N_391);
nand U6984 (N_6984,N_1429,N_4016);
nor U6985 (N_6985,N_688,N_292);
or U6986 (N_6986,N_2751,N_1448);
or U6987 (N_6987,N_2346,N_2645);
xor U6988 (N_6988,N_2622,N_1114);
nor U6989 (N_6989,N_3839,N_769);
or U6990 (N_6990,N_1460,N_1715);
nand U6991 (N_6991,N_4287,N_2379);
and U6992 (N_6992,N_1578,N_4479);
or U6993 (N_6993,N_457,N_636);
xnor U6994 (N_6994,N_381,N_152);
nand U6995 (N_6995,N_2289,N_3454);
or U6996 (N_6996,N_555,N_1495);
nand U6997 (N_6997,N_574,N_883);
and U6998 (N_6998,N_2781,N_635);
xnor U6999 (N_6999,N_4868,N_3393);
nor U7000 (N_7000,N_302,N_1168);
xor U7001 (N_7001,N_3858,N_1441);
or U7002 (N_7002,N_2615,N_3712);
nand U7003 (N_7003,N_1375,N_1228);
nand U7004 (N_7004,N_3453,N_459);
nand U7005 (N_7005,N_4534,N_3800);
or U7006 (N_7006,N_1277,N_1812);
and U7007 (N_7007,N_2583,N_1196);
xor U7008 (N_7008,N_172,N_4260);
nand U7009 (N_7009,N_4907,N_3135);
nand U7010 (N_7010,N_1652,N_3762);
or U7011 (N_7011,N_1452,N_2183);
nand U7012 (N_7012,N_548,N_2134);
and U7013 (N_7013,N_3116,N_1166);
nor U7014 (N_7014,N_4007,N_1929);
nand U7015 (N_7015,N_2253,N_2931);
and U7016 (N_7016,N_3070,N_1868);
and U7017 (N_7017,N_4993,N_86);
xnor U7018 (N_7018,N_4471,N_400);
nand U7019 (N_7019,N_3272,N_2083);
and U7020 (N_7020,N_842,N_1996);
xor U7021 (N_7021,N_3746,N_3699);
nor U7022 (N_7022,N_3067,N_641);
xor U7023 (N_7023,N_164,N_1843);
and U7024 (N_7024,N_3695,N_2368);
or U7025 (N_7025,N_1889,N_4466);
nand U7026 (N_7026,N_3545,N_2212);
xnor U7027 (N_7027,N_1752,N_4863);
and U7028 (N_7028,N_4253,N_2950);
nand U7029 (N_7029,N_23,N_325);
nor U7030 (N_7030,N_1850,N_3191);
or U7031 (N_7031,N_3437,N_3461);
nor U7032 (N_7032,N_969,N_4520);
nand U7033 (N_7033,N_3619,N_3351);
or U7034 (N_7034,N_2367,N_4391);
nand U7035 (N_7035,N_1583,N_1036);
and U7036 (N_7036,N_1809,N_2884);
xor U7037 (N_7037,N_1543,N_4347);
xor U7038 (N_7038,N_932,N_1083);
and U7039 (N_7039,N_4945,N_4740);
nand U7040 (N_7040,N_3077,N_947);
nand U7041 (N_7041,N_4642,N_1403);
and U7042 (N_7042,N_4345,N_4958);
nand U7043 (N_7043,N_3596,N_1886);
or U7044 (N_7044,N_908,N_4842);
or U7045 (N_7045,N_482,N_1052);
nor U7046 (N_7046,N_1108,N_4293);
nand U7047 (N_7047,N_2084,N_3501);
and U7048 (N_7048,N_2757,N_3969);
and U7049 (N_7049,N_4049,N_330);
nor U7050 (N_7050,N_2643,N_2765);
or U7051 (N_7051,N_4765,N_3106);
and U7052 (N_7052,N_1230,N_4931);
nand U7053 (N_7053,N_1458,N_1337);
xnor U7054 (N_7054,N_673,N_268);
and U7055 (N_7055,N_31,N_2149);
xnor U7056 (N_7056,N_3360,N_85);
xnor U7057 (N_7057,N_1801,N_2602);
nor U7058 (N_7058,N_4570,N_4410);
nand U7059 (N_7059,N_1591,N_1126);
nand U7060 (N_7060,N_752,N_2733);
or U7061 (N_7061,N_942,N_654);
or U7062 (N_7062,N_323,N_2142);
and U7063 (N_7063,N_4450,N_4807);
or U7064 (N_7064,N_1222,N_1298);
nor U7065 (N_7065,N_4588,N_1241);
xnor U7066 (N_7066,N_108,N_3697);
xor U7067 (N_7067,N_4739,N_1353);
xnor U7068 (N_7068,N_1432,N_2653);
or U7069 (N_7069,N_3710,N_1813);
nand U7070 (N_7070,N_1680,N_3080);
or U7071 (N_7071,N_2052,N_2430);
or U7072 (N_7072,N_112,N_439);
xor U7073 (N_7073,N_3157,N_3669);
xnor U7074 (N_7074,N_4363,N_4042);
and U7075 (N_7075,N_1074,N_3957);
and U7076 (N_7076,N_1023,N_4849);
and U7077 (N_7077,N_2495,N_4385);
nand U7078 (N_7078,N_3919,N_3066);
or U7079 (N_7079,N_653,N_1154);
and U7080 (N_7080,N_3119,N_4212);
nand U7081 (N_7081,N_4853,N_1255);
nand U7082 (N_7082,N_3206,N_601);
and U7083 (N_7083,N_2290,N_1360);
nand U7084 (N_7084,N_4726,N_3542);
nor U7085 (N_7085,N_512,N_3739);
nor U7086 (N_7086,N_2918,N_4770);
xor U7087 (N_7087,N_3254,N_4545);
nor U7088 (N_7088,N_999,N_3281);
nand U7089 (N_7089,N_495,N_892);
nand U7090 (N_7090,N_2425,N_2789);
xnor U7091 (N_7091,N_1595,N_4443);
and U7092 (N_7092,N_747,N_1584);
nand U7093 (N_7093,N_3918,N_4829);
xor U7094 (N_7094,N_3856,N_2332);
or U7095 (N_7095,N_1549,N_1352);
nor U7096 (N_7096,N_3637,N_2443);
and U7097 (N_7097,N_3627,N_235);
xnor U7098 (N_7098,N_705,N_1248);
xnor U7099 (N_7099,N_2700,N_261);
xnor U7100 (N_7100,N_1724,N_786);
nor U7101 (N_7101,N_3297,N_3507);
nand U7102 (N_7102,N_4012,N_4384);
xnor U7103 (N_7103,N_1022,N_1854);
nor U7104 (N_7104,N_2605,N_1565);
nand U7105 (N_7105,N_4487,N_4105);
nand U7106 (N_7106,N_117,N_1518);
and U7107 (N_7107,N_3485,N_587);
or U7108 (N_7108,N_4437,N_2686);
nor U7109 (N_7109,N_397,N_2492);
or U7110 (N_7110,N_3350,N_1194);
and U7111 (N_7111,N_2397,N_3876);
and U7112 (N_7112,N_371,N_1622);
xor U7113 (N_7113,N_1251,N_510);
nor U7114 (N_7114,N_3582,N_1494);
nand U7115 (N_7115,N_2706,N_2063);
or U7116 (N_7116,N_2306,N_1702);
nor U7117 (N_7117,N_2944,N_1243);
nand U7118 (N_7118,N_2233,N_1958);
or U7119 (N_7119,N_497,N_2773);
and U7120 (N_7120,N_559,N_755);
or U7121 (N_7121,N_1671,N_530);
nand U7122 (N_7122,N_716,N_729);
or U7123 (N_7123,N_2091,N_3260);
and U7124 (N_7124,N_2912,N_703);
or U7125 (N_7125,N_2666,N_4656);
xnor U7126 (N_7126,N_4750,N_2338);
nand U7127 (N_7127,N_3030,N_3300);
and U7128 (N_7128,N_534,N_4942);
xnor U7129 (N_7129,N_216,N_2876);
xnor U7130 (N_7130,N_2447,N_4477);
nand U7131 (N_7131,N_1829,N_4788);
or U7132 (N_7132,N_1711,N_3996);
xor U7133 (N_7133,N_4241,N_3917);
xor U7134 (N_7134,N_1476,N_1419);
and U7135 (N_7135,N_3486,N_621);
xor U7136 (N_7136,N_4651,N_453);
nand U7137 (N_7137,N_169,N_3026);
xnor U7138 (N_7138,N_2853,N_433);
nor U7139 (N_7139,N_54,N_3768);
and U7140 (N_7140,N_2795,N_4943);
xor U7141 (N_7141,N_264,N_3229);
nand U7142 (N_7142,N_448,N_58);
xor U7143 (N_7143,N_4994,N_2574);
and U7144 (N_7144,N_3477,N_3233);
xor U7145 (N_7145,N_779,N_2372);
xnor U7146 (N_7146,N_2881,N_4240);
nor U7147 (N_7147,N_3548,N_1271);
nand U7148 (N_7148,N_356,N_2366);
and U7149 (N_7149,N_4953,N_3905);
xor U7150 (N_7150,N_3528,N_1225);
xnor U7151 (N_7151,N_3803,N_3424);
or U7152 (N_7152,N_4071,N_3936);
and U7153 (N_7153,N_4420,N_1756);
nand U7154 (N_7154,N_4222,N_2335);
and U7155 (N_7155,N_4887,N_2356);
or U7156 (N_7156,N_2378,N_967);
nor U7157 (N_7157,N_2599,N_1387);
nand U7158 (N_7158,N_4401,N_2586);
nor U7159 (N_7159,N_894,N_3152);
nor U7160 (N_7160,N_2764,N_1962);
xor U7161 (N_7161,N_2550,N_1873);
xor U7162 (N_7162,N_1871,N_4617);
xnor U7163 (N_7163,N_2153,N_4944);
xor U7164 (N_7164,N_1848,N_2024);
or U7165 (N_7165,N_328,N_4402);
nand U7166 (N_7166,N_1700,N_4957);
xor U7167 (N_7167,N_2075,N_1279);
nor U7168 (N_7168,N_757,N_3413);
nor U7169 (N_7169,N_236,N_671);
or U7170 (N_7170,N_658,N_3594);
or U7171 (N_7171,N_1306,N_4554);
nand U7172 (N_7172,N_2326,N_2440);
and U7173 (N_7173,N_2082,N_4215);
xor U7174 (N_7174,N_3463,N_1091);
or U7175 (N_7175,N_132,N_1822);
nand U7176 (N_7176,N_2157,N_245);
nor U7177 (N_7177,N_2549,N_538);
nor U7178 (N_7178,N_2610,N_4087);
and U7179 (N_7179,N_1024,N_1640);
and U7180 (N_7180,N_4108,N_4032);
and U7181 (N_7181,N_2809,N_1370);
or U7182 (N_7182,N_2461,N_4572);
xor U7183 (N_7183,N_2062,N_907);
or U7184 (N_7184,N_1872,N_1233);
xnor U7185 (N_7185,N_713,N_2830);
xor U7186 (N_7186,N_4352,N_3176);
nand U7187 (N_7187,N_2065,N_2032);
nand U7188 (N_7188,N_1960,N_3316);
and U7189 (N_7189,N_3110,N_3392);
xor U7190 (N_7190,N_1566,N_2404);
nor U7191 (N_7191,N_1320,N_3613);
or U7192 (N_7192,N_3959,N_4395);
or U7193 (N_7193,N_4901,N_4467);
and U7194 (N_7194,N_3182,N_2166);
nand U7195 (N_7195,N_4399,N_912);
nor U7196 (N_7196,N_3509,N_2903);
nor U7197 (N_7197,N_3421,N_4911);
nor U7198 (N_7198,N_3831,N_2529);
and U7199 (N_7199,N_4186,N_3405);
or U7200 (N_7200,N_2732,N_3353);
xnor U7201 (N_7201,N_4213,N_1755);
nor U7202 (N_7202,N_4100,N_4595);
xor U7203 (N_7203,N_798,N_864);
xnor U7204 (N_7204,N_1485,N_4034);
nand U7205 (N_7205,N_1569,N_1855);
nand U7206 (N_7206,N_76,N_3012);
nor U7207 (N_7207,N_3520,N_3924);
nand U7208 (N_7208,N_1516,N_1585);
nor U7209 (N_7209,N_1836,N_1383);
nor U7210 (N_7210,N_4425,N_3342);
and U7211 (N_7211,N_2008,N_1696);
and U7212 (N_7212,N_2897,N_3430);
xor U7213 (N_7213,N_3921,N_1369);
nor U7214 (N_7214,N_2985,N_481);
nor U7215 (N_7215,N_1596,N_18);
xnor U7216 (N_7216,N_3199,N_59);
nand U7217 (N_7217,N_4073,N_2533);
or U7218 (N_7218,N_720,N_3912);
xnor U7219 (N_7219,N_2539,N_2720);
nor U7220 (N_7220,N_4470,N_3451);
and U7221 (N_7221,N_3086,N_2626);
xnor U7222 (N_7222,N_3626,N_1270);
xor U7223 (N_7223,N_1905,N_822);
nand U7224 (N_7224,N_1096,N_927);
nand U7225 (N_7225,N_186,N_1356);
nor U7226 (N_7226,N_2076,N_4935);
nor U7227 (N_7227,N_4760,N_4153);
or U7228 (N_7228,N_1313,N_2595);
and U7229 (N_7229,N_2850,N_194);
nand U7230 (N_7230,N_4025,N_1220);
nand U7231 (N_7231,N_3221,N_4824);
or U7232 (N_7232,N_4116,N_2682);
nand U7233 (N_7233,N_2759,N_1721);
nor U7234 (N_7234,N_3238,N_2493);
or U7235 (N_7235,N_936,N_561);
or U7236 (N_7236,N_3255,N_593);
nand U7237 (N_7237,N_3567,N_2955);
nor U7238 (N_7238,N_2020,N_1038);
and U7239 (N_7239,N_2267,N_3137);
xor U7240 (N_7240,N_940,N_4255);
or U7241 (N_7241,N_738,N_4493);
nor U7242 (N_7242,N_1849,N_1118);
or U7243 (N_7243,N_1026,N_1440);
xnor U7244 (N_7244,N_3153,N_347);
xnor U7245 (N_7245,N_1690,N_1949);
xnor U7246 (N_7246,N_3237,N_1020);
xor U7247 (N_7247,N_4362,N_3126);
and U7248 (N_7248,N_1647,N_4249);
nand U7249 (N_7249,N_405,N_4046);
nor U7250 (N_7250,N_3779,N_2178);
nor U7251 (N_7251,N_1490,N_1570);
and U7252 (N_7252,N_1644,N_1877);
nand U7253 (N_7253,N_3285,N_1956);
xor U7254 (N_7254,N_4165,N_2161);
nor U7255 (N_7255,N_3790,N_2816);
and U7256 (N_7256,N_1082,N_1483);
or U7257 (N_7257,N_3513,N_4269);
or U7258 (N_7258,N_2841,N_890);
xor U7259 (N_7259,N_1445,N_3441);
nor U7260 (N_7260,N_93,N_234);
xnor U7261 (N_7261,N_2135,N_4578);
nand U7262 (N_7262,N_4914,N_3305);
nand U7263 (N_7263,N_1071,N_2612);
nand U7264 (N_7264,N_1496,N_4044);
nand U7265 (N_7265,N_4204,N_166);
xnor U7266 (N_7266,N_1655,N_572);
or U7267 (N_7267,N_2402,N_3440);
or U7268 (N_7268,N_3492,N_1333);
xor U7269 (N_7269,N_3332,N_3115);
xnor U7270 (N_7270,N_1109,N_2433);
or U7271 (N_7271,N_3866,N_2247);
and U7272 (N_7272,N_2503,N_3129);
nor U7273 (N_7273,N_162,N_4733);
or U7274 (N_7274,N_163,N_1097);
or U7275 (N_7275,N_3662,N_3132);
and U7276 (N_7276,N_1586,N_3727);
or U7277 (N_7277,N_763,N_2582);
xnor U7278 (N_7278,N_1861,N_2722);
or U7279 (N_7279,N_4440,N_804);
nand U7280 (N_7280,N_2947,N_3034);
nand U7281 (N_7281,N_603,N_4024);
nor U7282 (N_7282,N_3672,N_45);
xor U7283 (N_7283,N_617,N_1930);
or U7284 (N_7284,N_2324,N_157);
xnor U7285 (N_7285,N_203,N_1267);
or U7286 (N_7286,N_2206,N_2756);
and U7287 (N_7287,N_4218,N_4946);
xnor U7288 (N_7288,N_3498,N_3833);
and U7289 (N_7289,N_1237,N_2636);
nor U7290 (N_7290,N_4359,N_4704);
nand U7291 (N_7291,N_2392,N_1245);
nor U7292 (N_7292,N_1410,N_3648);
nand U7293 (N_7293,N_2900,N_2202);
or U7294 (N_7294,N_796,N_3274);
and U7295 (N_7295,N_3880,N_4745);
or U7296 (N_7296,N_3079,N_3158);
and U7297 (N_7297,N_4585,N_1637);
xnor U7298 (N_7298,N_4703,N_1820);
nand U7299 (N_7299,N_3692,N_4159);
or U7300 (N_7300,N_3772,N_3592);
nand U7301 (N_7301,N_2221,N_1899);
xor U7302 (N_7302,N_3988,N_4705);
xor U7303 (N_7303,N_354,N_1981);
nand U7304 (N_7304,N_3145,N_1315);
nor U7305 (N_7305,N_4002,N_1064);
or U7306 (N_7306,N_1639,N_737);
nor U7307 (N_7307,N_1080,N_1513);
or U7308 (N_7308,N_4691,N_2993);
xor U7309 (N_7309,N_2552,N_1511);
or U7310 (N_7310,N_3965,N_3098);
and U7311 (N_7311,N_4522,N_571);
or U7312 (N_7312,N_1860,N_689);
and U7313 (N_7313,N_614,N_1685);
and U7314 (N_7314,N_3379,N_2750);
nor U7315 (N_7315,N_3923,N_3047);
or U7316 (N_7316,N_4435,N_4211);
and U7317 (N_7317,N_2945,N_1350);
and U7318 (N_7318,N_3111,N_2107);
or U7319 (N_7319,N_2303,N_2333);
or U7320 (N_7320,N_1545,N_3226);
or U7321 (N_7321,N_4295,N_1620);
or U7322 (N_7322,N_2522,N_1457);
nand U7323 (N_7323,N_3247,N_579);
or U7324 (N_7324,N_3515,N_4263);
or U7325 (N_7325,N_1059,N_3159);
xor U7326 (N_7326,N_2650,N_2631);
or U7327 (N_7327,N_1461,N_3541);
xnor U7328 (N_7328,N_121,N_2241);
nor U7329 (N_7329,N_401,N_1707);
and U7330 (N_7330,N_4346,N_2413);
nand U7331 (N_7331,N_521,N_3087);
nor U7332 (N_7332,N_1418,N_1468);
and U7333 (N_7333,N_3906,N_4276);
nor U7334 (N_7334,N_2761,N_3682);
xor U7335 (N_7335,N_1774,N_3952);
and U7336 (N_7336,N_4968,N_2359);
xor U7337 (N_7337,N_3986,N_1681);
nor U7338 (N_7338,N_3478,N_4323);
and U7339 (N_7339,N_3974,N_998);
nand U7340 (N_7340,N_1635,N_2787);
or U7341 (N_7341,N_1720,N_2548);
and U7342 (N_7342,N_681,N_2920);
or U7343 (N_7343,N_1985,N_2270);
nor U7344 (N_7344,N_2105,N_2353);
nand U7345 (N_7345,N_2033,N_1272);
and U7346 (N_7346,N_977,N_655);
and U7347 (N_7347,N_343,N_4372);
or U7348 (N_7348,N_4664,N_2298);
nand U7349 (N_7349,N_3598,N_2036);
nand U7350 (N_7350,N_1211,N_644);
or U7351 (N_7351,N_434,N_1472);
nor U7352 (N_7352,N_955,N_277);
or U7353 (N_7353,N_3397,N_4392);
nor U7354 (N_7354,N_1870,N_2933);
or U7355 (N_7355,N_4047,N_452);
nand U7356 (N_7356,N_1558,N_4929);
nand U7357 (N_7357,N_1993,N_3995);
xor U7358 (N_7358,N_2252,N_2707);
and U7359 (N_7359,N_3072,N_3239);
or U7360 (N_7360,N_3287,N_1335);
and U7361 (N_7361,N_549,N_602);
xor U7362 (N_7362,N_258,N_2003);
xor U7363 (N_7363,N_4700,N_3333);
nand U7364 (N_7364,N_3786,N_876);
or U7365 (N_7365,N_3290,N_1677);
xor U7366 (N_7366,N_1890,N_1924);
nand U7367 (N_7367,N_4903,N_4015);
xor U7368 (N_7368,N_532,N_219);
or U7369 (N_7369,N_4011,N_2744);
or U7370 (N_7370,N_550,N_100);
or U7371 (N_7371,N_65,N_4311);
xor U7372 (N_7372,N_1909,N_2942);
or U7373 (N_7373,N_314,N_4045);
xor U7374 (N_7374,N_4910,N_3164);
and U7375 (N_7375,N_3358,N_329);
nand U7376 (N_7376,N_1625,N_2780);
nand U7377 (N_7377,N_509,N_1515);
nand U7378 (N_7378,N_1718,N_2639);
or U7379 (N_7379,N_214,N_262);
xnor U7380 (N_7380,N_3495,N_2535);
nand U7381 (N_7381,N_2330,N_3656);
xor U7382 (N_7382,N_1050,N_2439);
or U7383 (N_7383,N_4900,N_2531);
xor U7384 (N_7384,N_2490,N_3325);
xor U7385 (N_7385,N_1523,N_577);
nor U7386 (N_7386,N_4710,N_1041);
nand U7387 (N_7387,N_2300,N_2027);
nand U7388 (N_7388,N_3188,N_2725);
xor U7389 (N_7389,N_4397,N_2774);
nand U7390 (N_7390,N_2509,N_3195);
or U7391 (N_7391,N_2974,N_1314);
and U7392 (N_7392,N_3457,N_1669);
nand U7393 (N_7393,N_2475,N_5);
xnor U7394 (N_7394,N_1787,N_456);
nor U7395 (N_7395,N_4612,N_8);
and U7396 (N_7396,N_2914,N_471);
and U7397 (N_7397,N_3389,N_4175);
and U7398 (N_7398,N_1368,N_465);
xor U7399 (N_7399,N_3820,N_2287);
nor U7400 (N_7400,N_4314,N_2351);
nor U7401 (N_7401,N_1300,N_3540);
xnor U7402 (N_7402,N_3061,N_938);
nand U7403 (N_7403,N_2224,N_224);
and U7404 (N_7404,N_2362,N_2709);
nand U7405 (N_7405,N_1863,N_4787);
or U7406 (N_7406,N_346,N_847);
nand U7407 (N_7407,N_2864,N_4275);
and U7408 (N_7408,N_2917,N_4302);
and U7409 (N_7409,N_2444,N_3151);
nand U7410 (N_7410,N_1852,N_1103);
and U7411 (N_7411,N_861,N_2029);
nand U7412 (N_7412,N_2108,N_2992);
nor U7413 (N_7413,N_3947,N_1745);
or U7414 (N_7414,N_3256,N_2680);
xnor U7415 (N_7415,N_1876,N_4199);
or U7416 (N_7416,N_3227,N_589);
or U7417 (N_7417,N_4179,N_1216);
nor U7418 (N_7418,N_3872,N_4542);
nand U7419 (N_7419,N_2994,N_3642);
xnor U7420 (N_7420,N_1593,N_2935);
or U7421 (N_7421,N_1420,N_3083);
nor U7422 (N_7422,N_4355,N_1278);
and U7423 (N_7423,N_2159,N_228);
nand U7424 (N_7424,N_1381,N_1821);
nand U7425 (N_7425,N_4517,N_2179);
and U7426 (N_7426,N_882,N_1544);
nand U7427 (N_7427,N_3742,N_492);
nand U7428 (N_7428,N_2156,N_1151);
and U7429 (N_7429,N_2350,N_4802);
nand U7430 (N_7430,N_485,N_2648);
and U7431 (N_7431,N_1953,N_1427);
and U7432 (N_7432,N_4850,N_2632);
nor U7433 (N_7433,N_3166,N_1773);
and U7434 (N_7434,N_406,N_3538);
and U7435 (N_7435,N_3794,N_4639);
nand U7436 (N_7436,N_2637,N_2597);
or U7437 (N_7437,N_2163,N_4226);
and U7438 (N_7438,N_1802,N_1695);
nor U7439 (N_7439,N_3114,N_2181);
or U7440 (N_7440,N_3362,N_41);
and U7441 (N_7441,N_2133,N_2260);
nor U7442 (N_7442,N_2571,N_3990);
nand U7443 (N_7443,N_1349,N_1218);
and U7444 (N_7444,N_4149,N_2655);
and U7445 (N_7445,N_823,N_1380);
nand U7446 (N_7446,N_608,N_3442);
or U7447 (N_7447,N_728,N_2837);
and U7448 (N_7448,N_2344,N_2292);
nor U7449 (N_7449,N_1304,N_4262);
nand U7450 (N_7450,N_1077,N_3944);
nor U7451 (N_7451,N_113,N_3190);
or U7452 (N_7452,N_2100,N_1705);
and U7453 (N_7453,N_4052,N_4613);
and U7454 (N_7454,N_3681,N_1841);
nand U7455 (N_7455,N_1789,N_455);
nand U7456 (N_7456,N_581,N_215);
and U7457 (N_7457,N_519,N_275);
or U7458 (N_7458,N_1665,N_122);
and U7459 (N_7459,N_2486,N_4727);
and U7460 (N_7460,N_4655,N_4896);
xnor U7461 (N_7461,N_4307,N_4594);
or U7462 (N_7462,N_3078,N_2681);
xor U7463 (N_7463,N_3713,N_2314);
xnor U7464 (N_7464,N_2309,N_1726);
nor U7465 (N_7465,N_4246,N_2729);
and U7466 (N_7466,N_954,N_3771);
xnor U7467 (N_7467,N_1040,N_3217);
nor U7468 (N_7468,N_1318,N_2852);
nand U7469 (N_7469,N_4296,N_1674);
xor U7470 (N_7470,N_1042,N_2126);
nor U7471 (N_7471,N_2621,N_866);
nor U7472 (N_7472,N_1183,N_1757);
nand U7473 (N_7473,N_4137,N_87);
and U7474 (N_7474,N_4079,N_4351);
xnor U7475 (N_7475,N_4695,N_2002);
nand U7476 (N_7476,N_1101,N_2687);
nand U7477 (N_7477,N_4451,N_2959);
nor U7478 (N_7478,N_4939,N_3009);
xor U7479 (N_7479,N_1562,N_664);
xor U7480 (N_7480,N_2641,N_524);
nand U7481 (N_7481,N_1933,N_4120);
nand U7482 (N_7482,N_2418,N_802);
nand U7483 (N_7483,N_4256,N_3186);
xor U7484 (N_7484,N_1402,N_238);
nor U7485 (N_7485,N_2557,N_4173);
nor U7486 (N_7486,N_4593,N_1015);
xnor U7487 (N_7487,N_4706,N_81);
and U7488 (N_7488,N_935,N_3864);
nand U7489 (N_7489,N_77,N_4258);
and U7490 (N_7490,N_1324,N_2446);
and U7491 (N_7491,N_225,N_232);
or U7492 (N_7492,N_2516,N_2295);
or U7493 (N_7493,N_4232,N_374);
nand U7494 (N_7494,N_3645,N_202);
nor U7495 (N_7495,N_719,N_3591);
nand U7496 (N_7496,N_3465,N_1347);
nor U7497 (N_7497,N_3968,N_975);
xor U7498 (N_7498,N_4576,N_4983);
nand U7499 (N_7499,N_11,N_722);
nand U7500 (N_7500,N_179,N_3193);
nand U7501 (N_7501,N_3927,N_4325);
nor U7502 (N_7502,N_2083,N_1586);
xnor U7503 (N_7503,N_964,N_1461);
or U7504 (N_7504,N_385,N_4320);
xnor U7505 (N_7505,N_1179,N_3749);
and U7506 (N_7506,N_1347,N_4408);
nor U7507 (N_7507,N_3326,N_3528);
nand U7508 (N_7508,N_2706,N_3548);
nor U7509 (N_7509,N_1344,N_2312);
nor U7510 (N_7510,N_979,N_3778);
nand U7511 (N_7511,N_3726,N_2594);
or U7512 (N_7512,N_1014,N_3629);
nand U7513 (N_7513,N_18,N_2542);
and U7514 (N_7514,N_479,N_3293);
and U7515 (N_7515,N_2916,N_2834);
nor U7516 (N_7516,N_4565,N_3899);
and U7517 (N_7517,N_1397,N_1057);
and U7518 (N_7518,N_1892,N_1779);
nand U7519 (N_7519,N_936,N_4871);
and U7520 (N_7520,N_1215,N_4230);
xor U7521 (N_7521,N_3489,N_4618);
nor U7522 (N_7522,N_4453,N_556);
nand U7523 (N_7523,N_1100,N_3045);
and U7524 (N_7524,N_3815,N_717);
or U7525 (N_7525,N_235,N_609);
and U7526 (N_7526,N_3938,N_1075);
xor U7527 (N_7527,N_3738,N_3775);
or U7528 (N_7528,N_2738,N_37);
or U7529 (N_7529,N_4280,N_3571);
and U7530 (N_7530,N_4889,N_4897);
or U7531 (N_7531,N_4398,N_1868);
nor U7532 (N_7532,N_3003,N_4742);
nor U7533 (N_7533,N_1244,N_542);
nor U7534 (N_7534,N_3622,N_4130);
or U7535 (N_7535,N_2169,N_293);
or U7536 (N_7536,N_178,N_3231);
and U7537 (N_7537,N_449,N_3021);
nand U7538 (N_7538,N_3644,N_3605);
xnor U7539 (N_7539,N_133,N_2352);
nor U7540 (N_7540,N_2252,N_1564);
nand U7541 (N_7541,N_1145,N_965);
xor U7542 (N_7542,N_1165,N_727);
or U7543 (N_7543,N_1194,N_1756);
xor U7544 (N_7544,N_4356,N_3415);
xor U7545 (N_7545,N_3086,N_4142);
or U7546 (N_7546,N_1849,N_481);
nor U7547 (N_7547,N_631,N_2058);
xnor U7548 (N_7548,N_3550,N_1501);
nor U7549 (N_7549,N_1117,N_1681);
nor U7550 (N_7550,N_3915,N_2808);
nor U7551 (N_7551,N_375,N_501);
nand U7552 (N_7552,N_324,N_365);
xor U7553 (N_7553,N_2869,N_3284);
and U7554 (N_7554,N_4776,N_4399);
and U7555 (N_7555,N_1852,N_4707);
or U7556 (N_7556,N_1769,N_225);
xor U7557 (N_7557,N_3224,N_4923);
and U7558 (N_7558,N_3549,N_298);
nor U7559 (N_7559,N_3030,N_3322);
and U7560 (N_7560,N_724,N_2101);
xnor U7561 (N_7561,N_1671,N_2760);
nand U7562 (N_7562,N_2785,N_3000);
or U7563 (N_7563,N_4159,N_345);
and U7564 (N_7564,N_1925,N_1596);
nand U7565 (N_7565,N_195,N_1754);
and U7566 (N_7566,N_4924,N_4832);
and U7567 (N_7567,N_3583,N_2750);
nor U7568 (N_7568,N_2190,N_622);
xor U7569 (N_7569,N_1710,N_2829);
or U7570 (N_7570,N_1991,N_1373);
or U7571 (N_7571,N_4656,N_4462);
and U7572 (N_7572,N_3892,N_3755);
or U7573 (N_7573,N_3226,N_2396);
or U7574 (N_7574,N_21,N_781);
xnor U7575 (N_7575,N_3935,N_852);
and U7576 (N_7576,N_4864,N_1828);
xor U7577 (N_7577,N_3932,N_4202);
nand U7578 (N_7578,N_3038,N_4899);
nand U7579 (N_7579,N_1074,N_3209);
or U7580 (N_7580,N_117,N_3538);
nand U7581 (N_7581,N_450,N_2013);
and U7582 (N_7582,N_3433,N_3664);
nor U7583 (N_7583,N_1104,N_1737);
nand U7584 (N_7584,N_1936,N_3744);
nand U7585 (N_7585,N_3245,N_2693);
nand U7586 (N_7586,N_2069,N_2485);
nor U7587 (N_7587,N_2341,N_1654);
and U7588 (N_7588,N_4147,N_3323);
or U7589 (N_7589,N_967,N_690);
and U7590 (N_7590,N_1997,N_3190);
xor U7591 (N_7591,N_4580,N_4177);
and U7592 (N_7592,N_3873,N_3833);
or U7593 (N_7593,N_2884,N_1777);
xor U7594 (N_7594,N_2344,N_2362);
nand U7595 (N_7595,N_4974,N_599);
nand U7596 (N_7596,N_3356,N_2095);
or U7597 (N_7597,N_4540,N_4828);
xnor U7598 (N_7598,N_4460,N_2646);
or U7599 (N_7599,N_3739,N_4641);
xnor U7600 (N_7600,N_2242,N_569);
or U7601 (N_7601,N_4924,N_3628);
and U7602 (N_7602,N_4709,N_4660);
and U7603 (N_7603,N_111,N_523);
and U7604 (N_7604,N_503,N_2261);
xnor U7605 (N_7605,N_3914,N_3666);
nand U7606 (N_7606,N_1949,N_893);
and U7607 (N_7607,N_2650,N_905);
and U7608 (N_7608,N_2651,N_2607);
nor U7609 (N_7609,N_3504,N_2341);
or U7610 (N_7610,N_3289,N_2399);
nand U7611 (N_7611,N_2883,N_4132);
and U7612 (N_7612,N_4880,N_783);
nand U7613 (N_7613,N_2340,N_916);
or U7614 (N_7614,N_3857,N_3566);
nor U7615 (N_7615,N_3892,N_2670);
nand U7616 (N_7616,N_34,N_2438);
xor U7617 (N_7617,N_278,N_4627);
or U7618 (N_7618,N_4240,N_3114);
nand U7619 (N_7619,N_64,N_2329);
nand U7620 (N_7620,N_4115,N_4299);
and U7621 (N_7621,N_1930,N_1426);
or U7622 (N_7622,N_216,N_2815);
nor U7623 (N_7623,N_420,N_3728);
nand U7624 (N_7624,N_1493,N_2208);
nand U7625 (N_7625,N_3144,N_107);
xor U7626 (N_7626,N_4315,N_1295);
and U7627 (N_7627,N_2231,N_3056);
and U7628 (N_7628,N_4431,N_2458);
and U7629 (N_7629,N_2821,N_3864);
and U7630 (N_7630,N_3087,N_147);
xnor U7631 (N_7631,N_711,N_870);
nor U7632 (N_7632,N_4347,N_4691);
nand U7633 (N_7633,N_3403,N_1729);
xnor U7634 (N_7634,N_2783,N_227);
nor U7635 (N_7635,N_2691,N_3958);
nand U7636 (N_7636,N_4201,N_243);
or U7637 (N_7637,N_3248,N_3208);
nand U7638 (N_7638,N_2628,N_256);
or U7639 (N_7639,N_2959,N_591);
xor U7640 (N_7640,N_1279,N_127);
and U7641 (N_7641,N_4139,N_1147);
or U7642 (N_7642,N_4427,N_1881);
nor U7643 (N_7643,N_3980,N_1268);
and U7644 (N_7644,N_4553,N_4778);
or U7645 (N_7645,N_3247,N_3327);
nand U7646 (N_7646,N_1822,N_1816);
xnor U7647 (N_7647,N_1977,N_574);
and U7648 (N_7648,N_3243,N_2327);
nor U7649 (N_7649,N_3133,N_951);
xor U7650 (N_7650,N_678,N_1529);
or U7651 (N_7651,N_2946,N_1637);
nand U7652 (N_7652,N_799,N_4719);
and U7653 (N_7653,N_4292,N_4149);
xnor U7654 (N_7654,N_1075,N_3292);
xnor U7655 (N_7655,N_38,N_3915);
and U7656 (N_7656,N_3019,N_2642);
nor U7657 (N_7657,N_4926,N_872);
and U7658 (N_7658,N_2168,N_1546);
or U7659 (N_7659,N_946,N_2727);
or U7660 (N_7660,N_110,N_2532);
xor U7661 (N_7661,N_4528,N_4695);
xnor U7662 (N_7662,N_2496,N_3103);
nand U7663 (N_7663,N_2032,N_497);
nor U7664 (N_7664,N_2249,N_4272);
and U7665 (N_7665,N_3078,N_2314);
nand U7666 (N_7666,N_2650,N_930);
xnor U7667 (N_7667,N_3298,N_4325);
nand U7668 (N_7668,N_2065,N_208);
or U7669 (N_7669,N_2443,N_1282);
xor U7670 (N_7670,N_3559,N_1419);
nor U7671 (N_7671,N_4617,N_3471);
nand U7672 (N_7672,N_386,N_1156);
nand U7673 (N_7673,N_1495,N_3014);
or U7674 (N_7674,N_230,N_1411);
nor U7675 (N_7675,N_878,N_1581);
and U7676 (N_7676,N_471,N_2405);
or U7677 (N_7677,N_2647,N_2065);
nor U7678 (N_7678,N_4088,N_840);
and U7679 (N_7679,N_42,N_2654);
xnor U7680 (N_7680,N_3696,N_526);
xnor U7681 (N_7681,N_1981,N_1070);
and U7682 (N_7682,N_208,N_2844);
xnor U7683 (N_7683,N_1648,N_100);
and U7684 (N_7684,N_1281,N_2699);
nand U7685 (N_7685,N_4794,N_2522);
or U7686 (N_7686,N_4187,N_1678);
xnor U7687 (N_7687,N_670,N_3775);
xnor U7688 (N_7688,N_2712,N_642);
xnor U7689 (N_7689,N_4706,N_4912);
xnor U7690 (N_7690,N_3981,N_3895);
nand U7691 (N_7691,N_4616,N_1128);
and U7692 (N_7692,N_1030,N_933);
and U7693 (N_7693,N_1879,N_1288);
nor U7694 (N_7694,N_4191,N_2645);
or U7695 (N_7695,N_606,N_90);
nand U7696 (N_7696,N_2842,N_1083);
nor U7697 (N_7697,N_1237,N_2024);
nand U7698 (N_7698,N_585,N_4460);
and U7699 (N_7699,N_637,N_4698);
and U7700 (N_7700,N_3477,N_2212);
nor U7701 (N_7701,N_2921,N_968);
nor U7702 (N_7702,N_4023,N_2062);
and U7703 (N_7703,N_686,N_1766);
and U7704 (N_7704,N_3284,N_3876);
or U7705 (N_7705,N_1919,N_1363);
and U7706 (N_7706,N_2670,N_459);
nor U7707 (N_7707,N_4337,N_308);
nor U7708 (N_7708,N_2953,N_4885);
xor U7709 (N_7709,N_3075,N_236);
and U7710 (N_7710,N_2276,N_2747);
or U7711 (N_7711,N_3343,N_580);
or U7712 (N_7712,N_4777,N_4977);
and U7713 (N_7713,N_3710,N_4750);
or U7714 (N_7714,N_4582,N_893);
xnor U7715 (N_7715,N_4608,N_2928);
and U7716 (N_7716,N_404,N_1097);
nor U7717 (N_7717,N_4237,N_672);
and U7718 (N_7718,N_438,N_1133);
nand U7719 (N_7719,N_2711,N_156);
xnor U7720 (N_7720,N_3308,N_443);
xor U7721 (N_7721,N_943,N_8);
or U7722 (N_7722,N_1979,N_2972);
nor U7723 (N_7723,N_3460,N_3350);
or U7724 (N_7724,N_4191,N_1431);
xnor U7725 (N_7725,N_445,N_3987);
and U7726 (N_7726,N_3507,N_1215);
or U7727 (N_7727,N_3771,N_4397);
xor U7728 (N_7728,N_3130,N_26);
xnor U7729 (N_7729,N_274,N_2612);
xnor U7730 (N_7730,N_206,N_35);
xor U7731 (N_7731,N_233,N_919);
or U7732 (N_7732,N_2591,N_1960);
nor U7733 (N_7733,N_4634,N_2620);
or U7734 (N_7734,N_3382,N_2984);
nand U7735 (N_7735,N_159,N_3123);
nand U7736 (N_7736,N_1325,N_2018);
or U7737 (N_7737,N_4270,N_3370);
or U7738 (N_7738,N_4387,N_3324);
xor U7739 (N_7739,N_1826,N_517);
nor U7740 (N_7740,N_2661,N_1870);
and U7741 (N_7741,N_1063,N_954);
xor U7742 (N_7742,N_2535,N_2618);
nor U7743 (N_7743,N_3433,N_4971);
xor U7744 (N_7744,N_1315,N_3788);
nand U7745 (N_7745,N_3990,N_2622);
nand U7746 (N_7746,N_3971,N_4683);
and U7747 (N_7747,N_155,N_2541);
nor U7748 (N_7748,N_248,N_3433);
nand U7749 (N_7749,N_4348,N_2975);
xor U7750 (N_7750,N_248,N_4095);
nand U7751 (N_7751,N_3299,N_3482);
or U7752 (N_7752,N_2432,N_2194);
and U7753 (N_7753,N_3092,N_4898);
xor U7754 (N_7754,N_1738,N_2597);
xnor U7755 (N_7755,N_744,N_10);
xnor U7756 (N_7756,N_1335,N_1422);
xnor U7757 (N_7757,N_3524,N_3827);
nor U7758 (N_7758,N_3481,N_2544);
or U7759 (N_7759,N_3186,N_1330);
xnor U7760 (N_7760,N_3935,N_1987);
nor U7761 (N_7761,N_4731,N_1554);
or U7762 (N_7762,N_2322,N_4107);
or U7763 (N_7763,N_3745,N_2567);
or U7764 (N_7764,N_128,N_1596);
xnor U7765 (N_7765,N_4557,N_1629);
xnor U7766 (N_7766,N_1463,N_2622);
and U7767 (N_7767,N_4849,N_3930);
xnor U7768 (N_7768,N_3432,N_371);
and U7769 (N_7769,N_1539,N_4595);
nand U7770 (N_7770,N_3866,N_1613);
xor U7771 (N_7771,N_2861,N_630);
and U7772 (N_7772,N_3650,N_1117);
and U7773 (N_7773,N_1150,N_4772);
or U7774 (N_7774,N_1000,N_3160);
nor U7775 (N_7775,N_1777,N_3355);
and U7776 (N_7776,N_4097,N_4868);
nor U7777 (N_7777,N_4286,N_2040);
xnor U7778 (N_7778,N_226,N_968);
xor U7779 (N_7779,N_1214,N_613);
nand U7780 (N_7780,N_4311,N_4703);
and U7781 (N_7781,N_1067,N_1805);
and U7782 (N_7782,N_3875,N_1748);
or U7783 (N_7783,N_3269,N_231);
or U7784 (N_7784,N_551,N_2016);
and U7785 (N_7785,N_4069,N_1213);
nor U7786 (N_7786,N_3448,N_3071);
nor U7787 (N_7787,N_634,N_537);
xor U7788 (N_7788,N_173,N_290);
nand U7789 (N_7789,N_1158,N_4230);
nand U7790 (N_7790,N_3652,N_2417);
and U7791 (N_7791,N_4807,N_3688);
nor U7792 (N_7792,N_2884,N_2894);
and U7793 (N_7793,N_750,N_3000);
nand U7794 (N_7794,N_4991,N_4480);
nor U7795 (N_7795,N_3644,N_228);
or U7796 (N_7796,N_2444,N_1469);
xnor U7797 (N_7797,N_3362,N_2261);
and U7798 (N_7798,N_3452,N_1534);
nor U7799 (N_7799,N_1901,N_995);
and U7800 (N_7800,N_4562,N_2985);
nor U7801 (N_7801,N_3689,N_3164);
nor U7802 (N_7802,N_866,N_2320);
and U7803 (N_7803,N_1346,N_4617);
nor U7804 (N_7804,N_1783,N_346);
and U7805 (N_7805,N_2099,N_4904);
nor U7806 (N_7806,N_2217,N_418);
nor U7807 (N_7807,N_4603,N_2674);
and U7808 (N_7808,N_4346,N_2268);
and U7809 (N_7809,N_575,N_882);
xor U7810 (N_7810,N_3038,N_2101);
or U7811 (N_7811,N_2974,N_70);
or U7812 (N_7812,N_3158,N_2105);
and U7813 (N_7813,N_3440,N_704);
nor U7814 (N_7814,N_4210,N_2586);
nand U7815 (N_7815,N_1303,N_4339);
xor U7816 (N_7816,N_3032,N_2879);
and U7817 (N_7817,N_2391,N_3211);
xor U7818 (N_7818,N_2709,N_3503);
nor U7819 (N_7819,N_2933,N_3537);
nand U7820 (N_7820,N_3546,N_4910);
nor U7821 (N_7821,N_4017,N_2726);
nand U7822 (N_7822,N_3376,N_2508);
or U7823 (N_7823,N_4801,N_2375);
nand U7824 (N_7824,N_901,N_4295);
nor U7825 (N_7825,N_864,N_338);
nor U7826 (N_7826,N_1669,N_4389);
or U7827 (N_7827,N_3745,N_1550);
nor U7828 (N_7828,N_199,N_2291);
and U7829 (N_7829,N_1974,N_4426);
nor U7830 (N_7830,N_3960,N_2656);
or U7831 (N_7831,N_591,N_3862);
or U7832 (N_7832,N_2939,N_3910);
nand U7833 (N_7833,N_2917,N_780);
xor U7834 (N_7834,N_2304,N_4215);
xor U7835 (N_7835,N_3152,N_2717);
nor U7836 (N_7836,N_3518,N_3525);
nand U7837 (N_7837,N_912,N_3568);
and U7838 (N_7838,N_1763,N_3247);
or U7839 (N_7839,N_2856,N_3286);
nand U7840 (N_7840,N_3209,N_2788);
and U7841 (N_7841,N_2907,N_4133);
xnor U7842 (N_7842,N_376,N_2778);
nand U7843 (N_7843,N_572,N_683);
nand U7844 (N_7844,N_4832,N_2744);
and U7845 (N_7845,N_1175,N_140);
and U7846 (N_7846,N_1324,N_545);
or U7847 (N_7847,N_4449,N_3275);
and U7848 (N_7848,N_2903,N_1151);
nor U7849 (N_7849,N_3937,N_1588);
nand U7850 (N_7850,N_147,N_4933);
nor U7851 (N_7851,N_1817,N_2063);
nand U7852 (N_7852,N_11,N_811);
nor U7853 (N_7853,N_749,N_206);
xor U7854 (N_7854,N_1637,N_3133);
or U7855 (N_7855,N_2049,N_4645);
nor U7856 (N_7856,N_3038,N_1284);
nand U7857 (N_7857,N_3495,N_4214);
or U7858 (N_7858,N_1508,N_2254);
xor U7859 (N_7859,N_889,N_3985);
and U7860 (N_7860,N_1399,N_145);
nand U7861 (N_7861,N_2968,N_1229);
or U7862 (N_7862,N_186,N_4844);
xnor U7863 (N_7863,N_4220,N_4293);
nand U7864 (N_7864,N_4901,N_1382);
nor U7865 (N_7865,N_1537,N_1081);
and U7866 (N_7866,N_4170,N_3547);
and U7867 (N_7867,N_3103,N_1723);
and U7868 (N_7868,N_2719,N_4529);
xnor U7869 (N_7869,N_4664,N_4660);
xor U7870 (N_7870,N_3168,N_4469);
nand U7871 (N_7871,N_3255,N_164);
nand U7872 (N_7872,N_4116,N_4674);
xnor U7873 (N_7873,N_4510,N_1861);
or U7874 (N_7874,N_4692,N_671);
nor U7875 (N_7875,N_1432,N_3371);
xnor U7876 (N_7876,N_1188,N_354);
and U7877 (N_7877,N_1335,N_4810);
and U7878 (N_7878,N_4784,N_3352);
and U7879 (N_7879,N_2488,N_3216);
nand U7880 (N_7880,N_1383,N_1239);
and U7881 (N_7881,N_1777,N_2913);
and U7882 (N_7882,N_3311,N_1706);
or U7883 (N_7883,N_966,N_2954);
nand U7884 (N_7884,N_776,N_2275);
and U7885 (N_7885,N_1908,N_3566);
nor U7886 (N_7886,N_4663,N_4913);
or U7887 (N_7887,N_926,N_535);
or U7888 (N_7888,N_1511,N_3376);
nor U7889 (N_7889,N_3590,N_454);
nor U7890 (N_7890,N_4880,N_4531);
or U7891 (N_7891,N_3583,N_1086);
or U7892 (N_7892,N_4862,N_4824);
or U7893 (N_7893,N_4180,N_2689);
nand U7894 (N_7894,N_2579,N_776);
nand U7895 (N_7895,N_3195,N_4841);
or U7896 (N_7896,N_4615,N_1834);
nor U7897 (N_7897,N_4189,N_680);
and U7898 (N_7898,N_615,N_4192);
nor U7899 (N_7899,N_3989,N_498);
nor U7900 (N_7900,N_604,N_4209);
nor U7901 (N_7901,N_3332,N_1407);
or U7902 (N_7902,N_4292,N_2336);
or U7903 (N_7903,N_482,N_836);
nor U7904 (N_7904,N_3321,N_2535);
xnor U7905 (N_7905,N_2414,N_66);
and U7906 (N_7906,N_2414,N_2899);
xor U7907 (N_7907,N_4885,N_321);
nor U7908 (N_7908,N_3134,N_3105);
and U7909 (N_7909,N_620,N_3688);
nand U7910 (N_7910,N_3606,N_407);
nor U7911 (N_7911,N_3620,N_1962);
xor U7912 (N_7912,N_4911,N_2625);
nor U7913 (N_7913,N_4298,N_4039);
nand U7914 (N_7914,N_4236,N_3248);
nand U7915 (N_7915,N_4230,N_3128);
nor U7916 (N_7916,N_3374,N_561);
nand U7917 (N_7917,N_1905,N_3905);
or U7918 (N_7918,N_4150,N_3280);
xor U7919 (N_7919,N_2786,N_3046);
or U7920 (N_7920,N_2998,N_1007);
nor U7921 (N_7921,N_3849,N_1897);
xor U7922 (N_7922,N_2378,N_1471);
nand U7923 (N_7923,N_2796,N_3319);
nor U7924 (N_7924,N_4916,N_27);
or U7925 (N_7925,N_3246,N_3611);
nor U7926 (N_7926,N_2202,N_2406);
nor U7927 (N_7927,N_4021,N_1764);
nor U7928 (N_7928,N_4209,N_2277);
nor U7929 (N_7929,N_3344,N_811);
or U7930 (N_7930,N_2758,N_2540);
nor U7931 (N_7931,N_882,N_3288);
nand U7932 (N_7932,N_2502,N_1360);
or U7933 (N_7933,N_1856,N_1595);
nor U7934 (N_7934,N_262,N_4305);
nor U7935 (N_7935,N_3907,N_1322);
and U7936 (N_7936,N_3836,N_4160);
nand U7937 (N_7937,N_3374,N_1785);
or U7938 (N_7938,N_2922,N_599);
xor U7939 (N_7939,N_1557,N_4221);
or U7940 (N_7940,N_2769,N_3303);
xor U7941 (N_7941,N_671,N_957);
and U7942 (N_7942,N_1010,N_4807);
nor U7943 (N_7943,N_3916,N_900);
nor U7944 (N_7944,N_2641,N_894);
nor U7945 (N_7945,N_2628,N_4886);
xnor U7946 (N_7946,N_1648,N_2233);
nand U7947 (N_7947,N_2993,N_3629);
xor U7948 (N_7948,N_1350,N_2971);
nand U7949 (N_7949,N_4695,N_4670);
xnor U7950 (N_7950,N_2130,N_3489);
nor U7951 (N_7951,N_1737,N_2747);
nor U7952 (N_7952,N_3114,N_498);
nor U7953 (N_7953,N_1459,N_3004);
or U7954 (N_7954,N_1007,N_1787);
nor U7955 (N_7955,N_4728,N_128);
or U7956 (N_7956,N_1449,N_4242);
nor U7957 (N_7957,N_4955,N_2029);
or U7958 (N_7958,N_1287,N_4240);
nand U7959 (N_7959,N_1934,N_3553);
and U7960 (N_7960,N_2566,N_4992);
xor U7961 (N_7961,N_2588,N_13);
or U7962 (N_7962,N_3887,N_4758);
or U7963 (N_7963,N_2144,N_145);
nand U7964 (N_7964,N_2934,N_3605);
nand U7965 (N_7965,N_43,N_3388);
nand U7966 (N_7966,N_2935,N_2285);
or U7967 (N_7967,N_662,N_673);
or U7968 (N_7968,N_2270,N_4401);
nand U7969 (N_7969,N_4236,N_2506);
nand U7970 (N_7970,N_3929,N_1614);
nand U7971 (N_7971,N_888,N_71);
nand U7972 (N_7972,N_200,N_3304);
nor U7973 (N_7973,N_4502,N_2161);
and U7974 (N_7974,N_722,N_2468);
or U7975 (N_7975,N_2379,N_2357);
nand U7976 (N_7976,N_3200,N_4807);
nor U7977 (N_7977,N_1484,N_1888);
and U7978 (N_7978,N_4198,N_3532);
and U7979 (N_7979,N_564,N_4479);
xor U7980 (N_7980,N_3406,N_2504);
and U7981 (N_7981,N_2730,N_4117);
xor U7982 (N_7982,N_3193,N_3596);
nor U7983 (N_7983,N_3468,N_2834);
nor U7984 (N_7984,N_920,N_2660);
or U7985 (N_7985,N_1275,N_614);
nand U7986 (N_7986,N_8,N_46);
or U7987 (N_7987,N_504,N_4552);
and U7988 (N_7988,N_2707,N_1643);
or U7989 (N_7989,N_72,N_19);
and U7990 (N_7990,N_4206,N_504);
or U7991 (N_7991,N_2694,N_715);
nor U7992 (N_7992,N_1863,N_3187);
xor U7993 (N_7993,N_4642,N_4261);
and U7994 (N_7994,N_3315,N_4110);
xnor U7995 (N_7995,N_2759,N_2621);
xor U7996 (N_7996,N_4497,N_3295);
or U7997 (N_7997,N_2266,N_2816);
xnor U7998 (N_7998,N_3698,N_2741);
nand U7999 (N_7999,N_3120,N_925);
nand U8000 (N_8000,N_1403,N_4377);
nor U8001 (N_8001,N_1365,N_3628);
and U8002 (N_8002,N_1612,N_4235);
or U8003 (N_8003,N_90,N_1673);
nand U8004 (N_8004,N_4126,N_2341);
nand U8005 (N_8005,N_2634,N_780);
nand U8006 (N_8006,N_3,N_2724);
and U8007 (N_8007,N_512,N_3968);
nand U8008 (N_8008,N_2278,N_3417);
or U8009 (N_8009,N_2081,N_3614);
and U8010 (N_8010,N_3486,N_1649);
and U8011 (N_8011,N_643,N_4985);
nand U8012 (N_8012,N_3435,N_3524);
nand U8013 (N_8013,N_3785,N_4710);
nand U8014 (N_8014,N_500,N_2132);
nor U8015 (N_8015,N_836,N_4899);
nand U8016 (N_8016,N_2269,N_1716);
and U8017 (N_8017,N_487,N_2056);
or U8018 (N_8018,N_4519,N_455);
nor U8019 (N_8019,N_1840,N_4445);
nand U8020 (N_8020,N_936,N_2831);
nor U8021 (N_8021,N_770,N_1769);
or U8022 (N_8022,N_2890,N_2113);
nand U8023 (N_8023,N_2696,N_58);
and U8024 (N_8024,N_2754,N_1995);
or U8025 (N_8025,N_1644,N_2989);
nand U8026 (N_8026,N_1894,N_1317);
nor U8027 (N_8027,N_2732,N_2604);
or U8028 (N_8028,N_622,N_1132);
nor U8029 (N_8029,N_1012,N_64);
xor U8030 (N_8030,N_1539,N_3324);
nand U8031 (N_8031,N_3583,N_4203);
or U8032 (N_8032,N_161,N_3024);
nand U8033 (N_8033,N_3015,N_4662);
or U8034 (N_8034,N_3410,N_4996);
or U8035 (N_8035,N_1000,N_847);
and U8036 (N_8036,N_2448,N_4203);
or U8037 (N_8037,N_1893,N_4220);
or U8038 (N_8038,N_3475,N_75);
nor U8039 (N_8039,N_1743,N_4248);
or U8040 (N_8040,N_1540,N_3613);
nand U8041 (N_8041,N_1680,N_1336);
and U8042 (N_8042,N_1775,N_2985);
xnor U8043 (N_8043,N_2509,N_937);
nor U8044 (N_8044,N_2416,N_1614);
and U8045 (N_8045,N_1195,N_380);
and U8046 (N_8046,N_230,N_450);
nand U8047 (N_8047,N_104,N_2446);
or U8048 (N_8048,N_816,N_1051);
xnor U8049 (N_8049,N_492,N_1474);
or U8050 (N_8050,N_2120,N_773);
and U8051 (N_8051,N_4763,N_4766);
nand U8052 (N_8052,N_1142,N_3062);
nor U8053 (N_8053,N_2812,N_2632);
xor U8054 (N_8054,N_3812,N_4089);
nand U8055 (N_8055,N_4251,N_4474);
nor U8056 (N_8056,N_1210,N_3156);
nor U8057 (N_8057,N_2471,N_1244);
or U8058 (N_8058,N_2560,N_4319);
and U8059 (N_8059,N_4061,N_3961);
nor U8060 (N_8060,N_772,N_4549);
or U8061 (N_8061,N_4734,N_4083);
or U8062 (N_8062,N_978,N_1579);
nor U8063 (N_8063,N_3643,N_2641);
nand U8064 (N_8064,N_2270,N_2923);
nand U8065 (N_8065,N_2817,N_3589);
and U8066 (N_8066,N_4195,N_1693);
nor U8067 (N_8067,N_1678,N_1726);
or U8068 (N_8068,N_2776,N_3638);
or U8069 (N_8069,N_3076,N_3698);
or U8070 (N_8070,N_1808,N_2506);
xnor U8071 (N_8071,N_2699,N_2196);
or U8072 (N_8072,N_1195,N_4050);
or U8073 (N_8073,N_4111,N_4689);
xor U8074 (N_8074,N_3980,N_869);
and U8075 (N_8075,N_4147,N_4311);
and U8076 (N_8076,N_1394,N_2000);
and U8077 (N_8077,N_3209,N_2391);
nor U8078 (N_8078,N_158,N_3702);
xor U8079 (N_8079,N_2818,N_612);
or U8080 (N_8080,N_1595,N_1397);
nor U8081 (N_8081,N_657,N_3083);
xor U8082 (N_8082,N_1791,N_2185);
nor U8083 (N_8083,N_4862,N_3010);
and U8084 (N_8084,N_538,N_3536);
or U8085 (N_8085,N_4531,N_2698);
or U8086 (N_8086,N_2316,N_4690);
nor U8087 (N_8087,N_2380,N_4163);
nand U8088 (N_8088,N_1460,N_3604);
nand U8089 (N_8089,N_567,N_4433);
and U8090 (N_8090,N_1008,N_4073);
and U8091 (N_8091,N_4444,N_4869);
xor U8092 (N_8092,N_1582,N_1132);
xor U8093 (N_8093,N_1113,N_88);
nand U8094 (N_8094,N_1119,N_345);
xor U8095 (N_8095,N_4049,N_3338);
nand U8096 (N_8096,N_3459,N_2462);
xor U8097 (N_8097,N_934,N_374);
or U8098 (N_8098,N_4968,N_4955);
and U8099 (N_8099,N_4869,N_2554);
nand U8100 (N_8100,N_749,N_2827);
and U8101 (N_8101,N_214,N_2866);
or U8102 (N_8102,N_697,N_2133);
or U8103 (N_8103,N_4610,N_3823);
and U8104 (N_8104,N_4933,N_4713);
or U8105 (N_8105,N_3049,N_2256);
or U8106 (N_8106,N_2142,N_3773);
and U8107 (N_8107,N_627,N_2446);
nand U8108 (N_8108,N_2695,N_1714);
xor U8109 (N_8109,N_3053,N_827);
nand U8110 (N_8110,N_2060,N_1578);
nor U8111 (N_8111,N_4107,N_1954);
or U8112 (N_8112,N_4199,N_3641);
and U8113 (N_8113,N_2415,N_2022);
xnor U8114 (N_8114,N_4137,N_2171);
nor U8115 (N_8115,N_2959,N_1431);
nor U8116 (N_8116,N_2913,N_2784);
nand U8117 (N_8117,N_1104,N_1879);
and U8118 (N_8118,N_3145,N_3418);
or U8119 (N_8119,N_3952,N_700);
and U8120 (N_8120,N_3609,N_315);
or U8121 (N_8121,N_2963,N_3769);
and U8122 (N_8122,N_3248,N_4041);
nand U8123 (N_8123,N_2035,N_3712);
nand U8124 (N_8124,N_2602,N_4221);
or U8125 (N_8125,N_3941,N_4250);
and U8126 (N_8126,N_1310,N_769);
xor U8127 (N_8127,N_4098,N_2734);
nor U8128 (N_8128,N_4787,N_1610);
or U8129 (N_8129,N_1698,N_1338);
or U8130 (N_8130,N_2575,N_595);
xor U8131 (N_8131,N_4013,N_2996);
and U8132 (N_8132,N_4444,N_4497);
nand U8133 (N_8133,N_2602,N_2168);
nand U8134 (N_8134,N_3512,N_4072);
nand U8135 (N_8135,N_968,N_2734);
and U8136 (N_8136,N_4192,N_1964);
or U8137 (N_8137,N_3993,N_4561);
xor U8138 (N_8138,N_3704,N_166);
and U8139 (N_8139,N_3766,N_1136);
nor U8140 (N_8140,N_1023,N_231);
nand U8141 (N_8141,N_2564,N_2632);
and U8142 (N_8142,N_1612,N_4376);
or U8143 (N_8143,N_4819,N_853);
and U8144 (N_8144,N_2747,N_1843);
nand U8145 (N_8145,N_4000,N_3983);
nand U8146 (N_8146,N_1561,N_4769);
nor U8147 (N_8147,N_4854,N_924);
nor U8148 (N_8148,N_2540,N_3683);
nor U8149 (N_8149,N_3731,N_2446);
and U8150 (N_8150,N_1035,N_4068);
nand U8151 (N_8151,N_2857,N_2995);
nand U8152 (N_8152,N_2845,N_1764);
or U8153 (N_8153,N_1736,N_76);
xor U8154 (N_8154,N_4838,N_2513);
or U8155 (N_8155,N_627,N_1757);
nor U8156 (N_8156,N_4994,N_845);
nor U8157 (N_8157,N_2315,N_3147);
xor U8158 (N_8158,N_3348,N_1167);
or U8159 (N_8159,N_278,N_1709);
and U8160 (N_8160,N_1625,N_2963);
or U8161 (N_8161,N_310,N_4945);
nand U8162 (N_8162,N_1458,N_304);
nor U8163 (N_8163,N_2881,N_2390);
or U8164 (N_8164,N_147,N_1367);
and U8165 (N_8165,N_3063,N_1370);
xor U8166 (N_8166,N_4978,N_327);
and U8167 (N_8167,N_436,N_1366);
or U8168 (N_8168,N_2411,N_4473);
nor U8169 (N_8169,N_3898,N_1275);
nor U8170 (N_8170,N_713,N_3727);
and U8171 (N_8171,N_1697,N_1514);
and U8172 (N_8172,N_390,N_2127);
nor U8173 (N_8173,N_2640,N_3334);
xnor U8174 (N_8174,N_2036,N_2525);
or U8175 (N_8175,N_1068,N_3749);
or U8176 (N_8176,N_4573,N_412);
or U8177 (N_8177,N_418,N_525);
or U8178 (N_8178,N_4829,N_152);
nand U8179 (N_8179,N_4289,N_4861);
or U8180 (N_8180,N_815,N_2834);
or U8181 (N_8181,N_4315,N_4623);
xnor U8182 (N_8182,N_1500,N_3000);
nor U8183 (N_8183,N_2611,N_2241);
and U8184 (N_8184,N_2226,N_2993);
and U8185 (N_8185,N_3959,N_3647);
nand U8186 (N_8186,N_4288,N_808);
and U8187 (N_8187,N_3238,N_1496);
and U8188 (N_8188,N_3546,N_3010);
nor U8189 (N_8189,N_1184,N_1858);
or U8190 (N_8190,N_3306,N_213);
and U8191 (N_8191,N_959,N_1011);
or U8192 (N_8192,N_3347,N_583);
or U8193 (N_8193,N_3888,N_1177);
nand U8194 (N_8194,N_1102,N_1910);
or U8195 (N_8195,N_572,N_2240);
nand U8196 (N_8196,N_1326,N_2822);
nand U8197 (N_8197,N_4320,N_1844);
and U8198 (N_8198,N_1491,N_832);
nor U8199 (N_8199,N_3735,N_4653);
xor U8200 (N_8200,N_1799,N_109);
or U8201 (N_8201,N_298,N_4357);
nand U8202 (N_8202,N_4508,N_3112);
nand U8203 (N_8203,N_4157,N_3732);
or U8204 (N_8204,N_4590,N_2876);
nor U8205 (N_8205,N_983,N_834);
and U8206 (N_8206,N_4438,N_3080);
or U8207 (N_8207,N_1482,N_4109);
and U8208 (N_8208,N_1093,N_180);
nor U8209 (N_8209,N_3591,N_3543);
and U8210 (N_8210,N_535,N_2878);
or U8211 (N_8211,N_1371,N_5);
and U8212 (N_8212,N_3680,N_1886);
nand U8213 (N_8213,N_2779,N_907);
nor U8214 (N_8214,N_1973,N_4030);
nor U8215 (N_8215,N_2325,N_1544);
and U8216 (N_8216,N_2147,N_1883);
or U8217 (N_8217,N_1251,N_3015);
nor U8218 (N_8218,N_2191,N_2409);
nand U8219 (N_8219,N_3237,N_740);
xor U8220 (N_8220,N_4523,N_3125);
nand U8221 (N_8221,N_2426,N_924);
nand U8222 (N_8222,N_2096,N_2180);
or U8223 (N_8223,N_1594,N_4675);
xnor U8224 (N_8224,N_3761,N_2093);
and U8225 (N_8225,N_4880,N_566);
and U8226 (N_8226,N_1273,N_4451);
and U8227 (N_8227,N_760,N_1508);
nand U8228 (N_8228,N_357,N_758);
or U8229 (N_8229,N_164,N_1207);
nand U8230 (N_8230,N_891,N_3298);
and U8231 (N_8231,N_2176,N_106);
nor U8232 (N_8232,N_4562,N_1178);
and U8233 (N_8233,N_1535,N_4997);
xnor U8234 (N_8234,N_3002,N_3113);
and U8235 (N_8235,N_1172,N_3956);
or U8236 (N_8236,N_3602,N_3861);
nor U8237 (N_8237,N_2220,N_610);
xor U8238 (N_8238,N_1609,N_1486);
nor U8239 (N_8239,N_1502,N_1640);
or U8240 (N_8240,N_2358,N_2089);
xor U8241 (N_8241,N_2964,N_1777);
and U8242 (N_8242,N_527,N_287);
and U8243 (N_8243,N_1756,N_3778);
nor U8244 (N_8244,N_2951,N_396);
xor U8245 (N_8245,N_244,N_2993);
nor U8246 (N_8246,N_2251,N_4015);
nor U8247 (N_8247,N_1891,N_4966);
nor U8248 (N_8248,N_282,N_3223);
nor U8249 (N_8249,N_374,N_2217);
xor U8250 (N_8250,N_4917,N_1109);
or U8251 (N_8251,N_1480,N_2446);
nand U8252 (N_8252,N_2896,N_3051);
nand U8253 (N_8253,N_3147,N_574);
nor U8254 (N_8254,N_4808,N_3615);
and U8255 (N_8255,N_101,N_640);
or U8256 (N_8256,N_1006,N_3141);
and U8257 (N_8257,N_1316,N_754);
nor U8258 (N_8258,N_3870,N_582);
and U8259 (N_8259,N_1640,N_3450);
and U8260 (N_8260,N_520,N_4858);
nor U8261 (N_8261,N_3888,N_3348);
or U8262 (N_8262,N_2501,N_214);
or U8263 (N_8263,N_900,N_3838);
or U8264 (N_8264,N_3482,N_3934);
or U8265 (N_8265,N_1427,N_3010);
nor U8266 (N_8266,N_4272,N_250);
xor U8267 (N_8267,N_2620,N_1029);
xnor U8268 (N_8268,N_2179,N_682);
nand U8269 (N_8269,N_2775,N_234);
or U8270 (N_8270,N_1783,N_3955);
nor U8271 (N_8271,N_3266,N_3196);
nand U8272 (N_8272,N_1134,N_132);
nand U8273 (N_8273,N_3584,N_183);
or U8274 (N_8274,N_354,N_3177);
and U8275 (N_8275,N_632,N_3073);
nand U8276 (N_8276,N_1009,N_1193);
xnor U8277 (N_8277,N_2661,N_2920);
or U8278 (N_8278,N_3110,N_176);
or U8279 (N_8279,N_1114,N_1227);
and U8280 (N_8280,N_427,N_1184);
nand U8281 (N_8281,N_3015,N_4783);
and U8282 (N_8282,N_1055,N_3412);
and U8283 (N_8283,N_2623,N_1750);
or U8284 (N_8284,N_227,N_1400);
nor U8285 (N_8285,N_3865,N_1578);
nor U8286 (N_8286,N_1076,N_1773);
nand U8287 (N_8287,N_2066,N_2766);
and U8288 (N_8288,N_1519,N_3436);
nand U8289 (N_8289,N_881,N_1881);
and U8290 (N_8290,N_3543,N_1280);
nor U8291 (N_8291,N_2622,N_1069);
nor U8292 (N_8292,N_2367,N_1685);
or U8293 (N_8293,N_4470,N_1785);
nor U8294 (N_8294,N_2227,N_360);
xor U8295 (N_8295,N_1518,N_762);
xnor U8296 (N_8296,N_2266,N_1536);
and U8297 (N_8297,N_4487,N_1919);
xnor U8298 (N_8298,N_4614,N_19);
or U8299 (N_8299,N_833,N_4107);
xnor U8300 (N_8300,N_2206,N_893);
xor U8301 (N_8301,N_3022,N_3684);
and U8302 (N_8302,N_365,N_3495);
and U8303 (N_8303,N_3459,N_1175);
or U8304 (N_8304,N_4386,N_4199);
nand U8305 (N_8305,N_3085,N_1960);
xor U8306 (N_8306,N_122,N_1750);
and U8307 (N_8307,N_778,N_94);
or U8308 (N_8308,N_3642,N_2375);
nand U8309 (N_8309,N_3207,N_2025);
xnor U8310 (N_8310,N_3948,N_2534);
or U8311 (N_8311,N_2533,N_1835);
nand U8312 (N_8312,N_2613,N_4715);
nand U8313 (N_8313,N_937,N_3977);
nand U8314 (N_8314,N_1121,N_508);
nor U8315 (N_8315,N_2889,N_905);
nor U8316 (N_8316,N_4986,N_144);
nor U8317 (N_8317,N_2260,N_4521);
or U8318 (N_8318,N_1011,N_152);
xnor U8319 (N_8319,N_15,N_292);
nor U8320 (N_8320,N_3891,N_2704);
or U8321 (N_8321,N_128,N_3502);
or U8322 (N_8322,N_2209,N_4637);
or U8323 (N_8323,N_171,N_1779);
and U8324 (N_8324,N_665,N_739);
nand U8325 (N_8325,N_3442,N_1324);
nand U8326 (N_8326,N_3309,N_4223);
xnor U8327 (N_8327,N_1264,N_4774);
and U8328 (N_8328,N_2273,N_2481);
nand U8329 (N_8329,N_811,N_1020);
xor U8330 (N_8330,N_2066,N_121);
or U8331 (N_8331,N_1663,N_1107);
and U8332 (N_8332,N_1630,N_4544);
or U8333 (N_8333,N_4620,N_4219);
nor U8334 (N_8334,N_1550,N_4062);
nand U8335 (N_8335,N_1942,N_2150);
nor U8336 (N_8336,N_186,N_3402);
and U8337 (N_8337,N_2818,N_3425);
nor U8338 (N_8338,N_4213,N_2710);
and U8339 (N_8339,N_1081,N_3911);
nor U8340 (N_8340,N_2762,N_952);
xnor U8341 (N_8341,N_2455,N_3879);
nand U8342 (N_8342,N_1401,N_1786);
or U8343 (N_8343,N_814,N_4464);
nand U8344 (N_8344,N_1960,N_3684);
nor U8345 (N_8345,N_2669,N_491);
xnor U8346 (N_8346,N_3345,N_3884);
nand U8347 (N_8347,N_4312,N_753);
nor U8348 (N_8348,N_1853,N_794);
xor U8349 (N_8349,N_1778,N_435);
and U8350 (N_8350,N_1346,N_1818);
nor U8351 (N_8351,N_2816,N_2836);
nand U8352 (N_8352,N_3273,N_4256);
xor U8353 (N_8353,N_1677,N_3734);
xor U8354 (N_8354,N_4251,N_1577);
nand U8355 (N_8355,N_880,N_2428);
and U8356 (N_8356,N_1417,N_4461);
xnor U8357 (N_8357,N_2727,N_814);
nor U8358 (N_8358,N_3649,N_4048);
xor U8359 (N_8359,N_4831,N_726);
nand U8360 (N_8360,N_2793,N_3270);
nand U8361 (N_8361,N_572,N_2196);
and U8362 (N_8362,N_3061,N_3938);
and U8363 (N_8363,N_1712,N_3516);
and U8364 (N_8364,N_3731,N_4011);
and U8365 (N_8365,N_3582,N_1486);
nor U8366 (N_8366,N_413,N_3533);
nor U8367 (N_8367,N_2692,N_4267);
and U8368 (N_8368,N_2343,N_1070);
xor U8369 (N_8369,N_593,N_2044);
nor U8370 (N_8370,N_2909,N_3656);
nor U8371 (N_8371,N_4850,N_2429);
nor U8372 (N_8372,N_2026,N_3334);
nand U8373 (N_8373,N_4039,N_2024);
or U8374 (N_8374,N_2208,N_769);
nor U8375 (N_8375,N_1497,N_2815);
nand U8376 (N_8376,N_1510,N_2324);
and U8377 (N_8377,N_3187,N_1104);
nor U8378 (N_8378,N_2767,N_4887);
or U8379 (N_8379,N_332,N_1549);
nor U8380 (N_8380,N_2835,N_2320);
xnor U8381 (N_8381,N_1197,N_485);
nor U8382 (N_8382,N_4834,N_1519);
xor U8383 (N_8383,N_1056,N_2264);
xor U8384 (N_8384,N_4256,N_4399);
xor U8385 (N_8385,N_3540,N_4845);
and U8386 (N_8386,N_4445,N_2474);
xor U8387 (N_8387,N_4482,N_4768);
nor U8388 (N_8388,N_2830,N_3836);
and U8389 (N_8389,N_1700,N_3001);
nor U8390 (N_8390,N_2490,N_1702);
nor U8391 (N_8391,N_4544,N_2383);
and U8392 (N_8392,N_1944,N_3316);
nand U8393 (N_8393,N_4584,N_3942);
nand U8394 (N_8394,N_408,N_1946);
xor U8395 (N_8395,N_2429,N_2539);
and U8396 (N_8396,N_1005,N_2860);
nor U8397 (N_8397,N_2559,N_3259);
nor U8398 (N_8398,N_2602,N_4368);
nand U8399 (N_8399,N_2830,N_2083);
and U8400 (N_8400,N_2946,N_1266);
xor U8401 (N_8401,N_4865,N_4676);
nand U8402 (N_8402,N_3141,N_2893);
xnor U8403 (N_8403,N_4894,N_664);
and U8404 (N_8404,N_11,N_1354);
nand U8405 (N_8405,N_3133,N_1000);
xnor U8406 (N_8406,N_4800,N_3120);
and U8407 (N_8407,N_2266,N_2441);
or U8408 (N_8408,N_2489,N_4779);
nand U8409 (N_8409,N_3166,N_1491);
and U8410 (N_8410,N_4269,N_3893);
xnor U8411 (N_8411,N_4827,N_2321);
or U8412 (N_8412,N_85,N_2549);
xor U8413 (N_8413,N_2255,N_1227);
xor U8414 (N_8414,N_2611,N_1183);
and U8415 (N_8415,N_3541,N_2571);
nand U8416 (N_8416,N_3294,N_4533);
nand U8417 (N_8417,N_4896,N_3813);
xor U8418 (N_8418,N_4669,N_4779);
or U8419 (N_8419,N_4582,N_4697);
nor U8420 (N_8420,N_2645,N_2011);
or U8421 (N_8421,N_4293,N_65);
nor U8422 (N_8422,N_1507,N_4266);
xnor U8423 (N_8423,N_1423,N_3726);
nand U8424 (N_8424,N_2814,N_4795);
or U8425 (N_8425,N_2641,N_4985);
and U8426 (N_8426,N_3820,N_1232);
nor U8427 (N_8427,N_2392,N_574);
nor U8428 (N_8428,N_1705,N_3266);
nand U8429 (N_8429,N_3787,N_528);
nand U8430 (N_8430,N_1283,N_1579);
and U8431 (N_8431,N_1059,N_2774);
nand U8432 (N_8432,N_1657,N_2557);
xor U8433 (N_8433,N_2048,N_4475);
and U8434 (N_8434,N_4187,N_660);
nand U8435 (N_8435,N_2178,N_3565);
xnor U8436 (N_8436,N_1013,N_2370);
and U8437 (N_8437,N_4884,N_966);
or U8438 (N_8438,N_3198,N_4934);
nor U8439 (N_8439,N_1825,N_4365);
nor U8440 (N_8440,N_4797,N_1138);
nor U8441 (N_8441,N_1713,N_3133);
or U8442 (N_8442,N_219,N_2328);
and U8443 (N_8443,N_4283,N_114);
nand U8444 (N_8444,N_4786,N_982);
xor U8445 (N_8445,N_4110,N_2682);
nor U8446 (N_8446,N_4200,N_3703);
or U8447 (N_8447,N_4976,N_303);
or U8448 (N_8448,N_2346,N_2812);
or U8449 (N_8449,N_4585,N_4366);
and U8450 (N_8450,N_356,N_697);
or U8451 (N_8451,N_4036,N_841);
nor U8452 (N_8452,N_3374,N_2472);
and U8453 (N_8453,N_156,N_3128);
and U8454 (N_8454,N_80,N_2608);
or U8455 (N_8455,N_3648,N_150);
nor U8456 (N_8456,N_3319,N_452);
or U8457 (N_8457,N_2030,N_4921);
or U8458 (N_8458,N_194,N_1077);
or U8459 (N_8459,N_805,N_4455);
xnor U8460 (N_8460,N_4704,N_4489);
nand U8461 (N_8461,N_1817,N_550);
nor U8462 (N_8462,N_866,N_1706);
and U8463 (N_8463,N_2936,N_1928);
or U8464 (N_8464,N_83,N_387);
and U8465 (N_8465,N_1207,N_4730);
or U8466 (N_8466,N_2139,N_3332);
and U8467 (N_8467,N_4730,N_1098);
nor U8468 (N_8468,N_1543,N_4370);
nand U8469 (N_8469,N_3682,N_2698);
nor U8470 (N_8470,N_2196,N_1254);
nor U8471 (N_8471,N_54,N_59);
nand U8472 (N_8472,N_2599,N_1038);
and U8473 (N_8473,N_1949,N_3315);
or U8474 (N_8474,N_3207,N_4095);
nand U8475 (N_8475,N_2273,N_4181);
xor U8476 (N_8476,N_2021,N_4023);
nand U8477 (N_8477,N_816,N_378);
or U8478 (N_8478,N_4914,N_3618);
and U8479 (N_8479,N_4497,N_3340);
and U8480 (N_8480,N_2495,N_18);
or U8481 (N_8481,N_1578,N_4422);
and U8482 (N_8482,N_823,N_1851);
xor U8483 (N_8483,N_3796,N_3536);
or U8484 (N_8484,N_2833,N_187);
nor U8485 (N_8485,N_3615,N_1898);
nand U8486 (N_8486,N_3518,N_3350);
xor U8487 (N_8487,N_2425,N_4446);
or U8488 (N_8488,N_4240,N_757);
nand U8489 (N_8489,N_2765,N_3061);
and U8490 (N_8490,N_4273,N_3502);
xor U8491 (N_8491,N_4951,N_3293);
or U8492 (N_8492,N_1026,N_4996);
xor U8493 (N_8493,N_3940,N_743);
and U8494 (N_8494,N_3502,N_3147);
nand U8495 (N_8495,N_2671,N_2259);
nor U8496 (N_8496,N_3970,N_1455);
or U8497 (N_8497,N_4863,N_1308);
and U8498 (N_8498,N_4150,N_2270);
nand U8499 (N_8499,N_1928,N_1525);
nor U8500 (N_8500,N_4719,N_1483);
nor U8501 (N_8501,N_1498,N_3006);
xor U8502 (N_8502,N_2771,N_1024);
and U8503 (N_8503,N_356,N_1852);
nor U8504 (N_8504,N_3651,N_4377);
or U8505 (N_8505,N_92,N_3337);
or U8506 (N_8506,N_1853,N_2113);
xor U8507 (N_8507,N_1468,N_969);
or U8508 (N_8508,N_2029,N_1653);
or U8509 (N_8509,N_2514,N_3788);
and U8510 (N_8510,N_2989,N_3529);
nand U8511 (N_8511,N_2010,N_3734);
and U8512 (N_8512,N_820,N_2878);
nor U8513 (N_8513,N_1111,N_2159);
xnor U8514 (N_8514,N_1099,N_4042);
or U8515 (N_8515,N_3229,N_2494);
or U8516 (N_8516,N_1591,N_3428);
nand U8517 (N_8517,N_3768,N_877);
nand U8518 (N_8518,N_835,N_942);
xor U8519 (N_8519,N_731,N_486);
nor U8520 (N_8520,N_1753,N_571);
xnor U8521 (N_8521,N_3474,N_169);
or U8522 (N_8522,N_4376,N_4286);
xor U8523 (N_8523,N_4033,N_2529);
nor U8524 (N_8524,N_12,N_292);
nand U8525 (N_8525,N_1804,N_4797);
nand U8526 (N_8526,N_4726,N_2284);
and U8527 (N_8527,N_1627,N_172);
or U8528 (N_8528,N_2333,N_1809);
xor U8529 (N_8529,N_3971,N_2146);
or U8530 (N_8530,N_1954,N_721);
or U8531 (N_8531,N_781,N_2385);
xnor U8532 (N_8532,N_2229,N_2312);
xor U8533 (N_8533,N_4243,N_3936);
nor U8534 (N_8534,N_3454,N_2325);
and U8535 (N_8535,N_4752,N_1709);
xnor U8536 (N_8536,N_3687,N_3839);
xnor U8537 (N_8537,N_1318,N_641);
or U8538 (N_8538,N_1649,N_2258);
and U8539 (N_8539,N_1753,N_3150);
nand U8540 (N_8540,N_2533,N_3069);
nand U8541 (N_8541,N_447,N_454);
nand U8542 (N_8542,N_2885,N_3488);
xnor U8543 (N_8543,N_2026,N_3824);
nor U8544 (N_8544,N_4281,N_3225);
or U8545 (N_8545,N_3307,N_2318);
or U8546 (N_8546,N_854,N_1853);
nand U8547 (N_8547,N_4795,N_1972);
nor U8548 (N_8548,N_750,N_2393);
or U8549 (N_8549,N_3068,N_1102);
nand U8550 (N_8550,N_886,N_687);
nor U8551 (N_8551,N_2754,N_1401);
nor U8552 (N_8552,N_4382,N_1488);
and U8553 (N_8553,N_4890,N_4265);
nand U8554 (N_8554,N_898,N_2868);
or U8555 (N_8555,N_1321,N_3);
or U8556 (N_8556,N_4083,N_530);
xor U8557 (N_8557,N_2631,N_3675);
or U8558 (N_8558,N_1506,N_314);
xnor U8559 (N_8559,N_2018,N_1868);
nor U8560 (N_8560,N_1772,N_1561);
and U8561 (N_8561,N_4516,N_3053);
nor U8562 (N_8562,N_2896,N_3797);
or U8563 (N_8563,N_3159,N_1747);
nand U8564 (N_8564,N_2673,N_320);
nor U8565 (N_8565,N_4804,N_2403);
or U8566 (N_8566,N_448,N_705);
nand U8567 (N_8567,N_579,N_749);
xnor U8568 (N_8568,N_4923,N_814);
or U8569 (N_8569,N_2183,N_2239);
or U8570 (N_8570,N_4463,N_3451);
nand U8571 (N_8571,N_1506,N_3373);
and U8572 (N_8572,N_761,N_2632);
or U8573 (N_8573,N_2067,N_4725);
and U8574 (N_8574,N_551,N_1392);
nand U8575 (N_8575,N_2825,N_906);
nor U8576 (N_8576,N_3022,N_2259);
nand U8577 (N_8577,N_4198,N_3073);
nor U8578 (N_8578,N_3278,N_4566);
nand U8579 (N_8579,N_1072,N_4588);
xor U8580 (N_8580,N_906,N_4229);
and U8581 (N_8581,N_453,N_348);
or U8582 (N_8582,N_4878,N_4223);
or U8583 (N_8583,N_366,N_1137);
nor U8584 (N_8584,N_1002,N_2402);
or U8585 (N_8585,N_1451,N_4985);
or U8586 (N_8586,N_2439,N_4036);
and U8587 (N_8587,N_2941,N_2505);
nor U8588 (N_8588,N_3360,N_4422);
nand U8589 (N_8589,N_1822,N_2725);
xor U8590 (N_8590,N_2373,N_4701);
nor U8591 (N_8591,N_3356,N_210);
xnor U8592 (N_8592,N_3532,N_4526);
or U8593 (N_8593,N_1951,N_3749);
or U8594 (N_8594,N_239,N_4766);
nor U8595 (N_8595,N_58,N_474);
xnor U8596 (N_8596,N_1967,N_1);
and U8597 (N_8597,N_2754,N_1035);
and U8598 (N_8598,N_4909,N_18);
or U8599 (N_8599,N_2382,N_4812);
or U8600 (N_8600,N_870,N_666);
or U8601 (N_8601,N_4302,N_1054);
and U8602 (N_8602,N_3356,N_1544);
nand U8603 (N_8603,N_1040,N_1715);
and U8604 (N_8604,N_4268,N_4963);
nor U8605 (N_8605,N_926,N_703);
or U8606 (N_8606,N_2251,N_414);
nand U8607 (N_8607,N_1554,N_1168);
xnor U8608 (N_8608,N_2229,N_2212);
xor U8609 (N_8609,N_3717,N_467);
xnor U8610 (N_8610,N_508,N_4487);
nand U8611 (N_8611,N_3839,N_4750);
nand U8612 (N_8612,N_1594,N_418);
nor U8613 (N_8613,N_1101,N_1774);
nor U8614 (N_8614,N_2717,N_2798);
nor U8615 (N_8615,N_1684,N_406);
nor U8616 (N_8616,N_4792,N_3380);
and U8617 (N_8617,N_4323,N_3453);
nand U8618 (N_8618,N_1717,N_321);
xor U8619 (N_8619,N_3188,N_1364);
nand U8620 (N_8620,N_4457,N_4239);
nand U8621 (N_8621,N_374,N_3448);
nand U8622 (N_8622,N_1665,N_1587);
xnor U8623 (N_8623,N_2427,N_1855);
nor U8624 (N_8624,N_2579,N_127);
or U8625 (N_8625,N_4335,N_1277);
nor U8626 (N_8626,N_4156,N_593);
or U8627 (N_8627,N_1927,N_3588);
or U8628 (N_8628,N_3142,N_841);
or U8629 (N_8629,N_4619,N_1147);
or U8630 (N_8630,N_3876,N_4457);
nor U8631 (N_8631,N_1306,N_3669);
and U8632 (N_8632,N_1900,N_4009);
nor U8633 (N_8633,N_2842,N_4923);
nand U8634 (N_8634,N_4835,N_2359);
nor U8635 (N_8635,N_2601,N_3031);
nor U8636 (N_8636,N_1879,N_696);
or U8637 (N_8637,N_3362,N_1416);
or U8638 (N_8638,N_2191,N_770);
xnor U8639 (N_8639,N_1719,N_2474);
or U8640 (N_8640,N_356,N_853);
and U8641 (N_8641,N_1688,N_1959);
or U8642 (N_8642,N_1908,N_2029);
nand U8643 (N_8643,N_3802,N_1002);
xor U8644 (N_8644,N_1704,N_2598);
and U8645 (N_8645,N_627,N_3639);
xor U8646 (N_8646,N_1493,N_1644);
nor U8647 (N_8647,N_4150,N_46);
nand U8648 (N_8648,N_1058,N_3762);
xnor U8649 (N_8649,N_2758,N_2167);
xor U8650 (N_8650,N_4887,N_4422);
xnor U8651 (N_8651,N_4416,N_4792);
and U8652 (N_8652,N_4745,N_4367);
nor U8653 (N_8653,N_3997,N_2015);
xor U8654 (N_8654,N_3347,N_1940);
and U8655 (N_8655,N_2998,N_3111);
and U8656 (N_8656,N_3598,N_4143);
nor U8657 (N_8657,N_2815,N_281);
xor U8658 (N_8658,N_1444,N_836);
and U8659 (N_8659,N_4822,N_150);
and U8660 (N_8660,N_1751,N_4450);
and U8661 (N_8661,N_4694,N_4544);
nand U8662 (N_8662,N_4885,N_3457);
and U8663 (N_8663,N_115,N_1805);
xnor U8664 (N_8664,N_2398,N_608);
nand U8665 (N_8665,N_3372,N_2283);
and U8666 (N_8666,N_4618,N_2900);
xor U8667 (N_8667,N_4763,N_2220);
and U8668 (N_8668,N_3360,N_4042);
nand U8669 (N_8669,N_2639,N_437);
nand U8670 (N_8670,N_1283,N_2111);
nand U8671 (N_8671,N_3949,N_4645);
or U8672 (N_8672,N_4551,N_1470);
or U8673 (N_8673,N_2217,N_3952);
and U8674 (N_8674,N_4828,N_4875);
xnor U8675 (N_8675,N_1526,N_1277);
and U8676 (N_8676,N_2897,N_576);
and U8677 (N_8677,N_846,N_2958);
nand U8678 (N_8678,N_2706,N_294);
nand U8679 (N_8679,N_4653,N_3595);
xor U8680 (N_8680,N_1594,N_4322);
nand U8681 (N_8681,N_4398,N_58);
xor U8682 (N_8682,N_624,N_3528);
and U8683 (N_8683,N_3226,N_3246);
and U8684 (N_8684,N_4829,N_1031);
xnor U8685 (N_8685,N_3923,N_1559);
or U8686 (N_8686,N_2175,N_3957);
nand U8687 (N_8687,N_2681,N_1540);
nand U8688 (N_8688,N_2010,N_2730);
xor U8689 (N_8689,N_4707,N_2567);
nand U8690 (N_8690,N_1953,N_3046);
nor U8691 (N_8691,N_784,N_3856);
nor U8692 (N_8692,N_3815,N_4083);
nand U8693 (N_8693,N_1772,N_2101);
and U8694 (N_8694,N_3900,N_745);
nor U8695 (N_8695,N_3380,N_1455);
nand U8696 (N_8696,N_4198,N_4428);
nor U8697 (N_8697,N_3975,N_3702);
nor U8698 (N_8698,N_1040,N_2442);
xnor U8699 (N_8699,N_1272,N_2191);
or U8700 (N_8700,N_4154,N_799);
nand U8701 (N_8701,N_4040,N_4961);
and U8702 (N_8702,N_1481,N_4195);
xor U8703 (N_8703,N_4610,N_422);
xnor U8704 (N_8704,N_59,N_4824);
nand U8705 (N_8705,N_501,N_2809);
xor U8706 (N_8706,N_646,N_1726);
xnor U8707 (N_8707,N_659,N_1563);
or U8708 (N_8708,N_2845,N_4006);
nand U8709 (N_8709,N_2479,N_3221);
and U8710 (N_8710,N_2491,N_3598);
xnor U8711 (N_8711,N_1943,N_3932);
and U8712 (N_8712,N_20,N_3852);
nor U8713 (N_8713,N_2560,N_2447);
xor U8714 (N_8714,N_4399,N_3157);
or U8715 (N_8715,N_1623,N_2345);
nor U8716 (N_8716,N_2775,N_463);
nand U8717 (N_8717,N_3452,N_182);
nand U8718 (N_8718,N_740,N_1256);
or U8719 (N_8719,N_785,N_1797);
nor U8720 (N_8720,N_1619,N_1007);
nand U8721 (N_8721,N_3950,N_4987);
or U8722 (N_8722,N_1667,N_43);
or U8723 (N_8723,N_1450,N_3392);
and U8724 (N_8724,N_1963,N_1195);
nor U8725 (N_8725,N_1176,N_3594);
or U8726 (N_8726,N_853,N_2186);
nand U8727 (N_8727,N_4072,N_1909);
xnor U8728 (N_8728,N_4451,N_1114);
nand U8729 (N_8729,N_1258,N_1450);
nor U8730 (N_8730,N_2301,N_2161);
nor U8731 (N_8731,N_622,N_2355);
nand U8732 (N_8732,N_2813,N_4301);
nor U8733 (N_8733,N_1784,N_1261);
or U8734 (N_8734,N_2514,N_3975);
nand U8735 (N_8735,N_4118,N_3823);
nand U8736 (N_8736,N_4685,N_1881);
xor U8737 (N_8737,N_4283,N_2819);
xor U8738 (N_8738,N_1160,N_424);
and U8739 (N_8739,N_398,N_3199);
xnor U8740 (N_8740,N_3627,N_2720);
nor U8741 (N_8741,N_1646,N_214);
or U8742 (N_8742,N_3125,N_1689);
nand U8743 (N_8743,N_3376,N_2858);
nor U8744 (N_8744,N_2981,N_1961);
nor U8745 (N_8745,N_37,N_2908);
xor U8746 (N_8746,N_197,N_4085);
nor U8747 (N_8747,N_2835,N_532);
xor U8748 (N_8748,N_3745,N_971);
nand U8749 (N_8749,N_564,N_2234);
xor U8750 (N_8750,N_3030,N_4429);
xor U8751 (N_8751,N_4624,N_4457);
xor U8752 (N_8752,N_4948,N_1073);
nor U8753 (N_8753,N_4211,N_1744);
and U8754 (N_8754,N_4901,N_1395);
and U8755 (N_8755,N_2145,N_3626);
and U8756 (N_8756,N_53,N_3147);
and U8757 (N_8757,N_4580,N_2290);
nor U8758 (N_8758,N_2092,N_251);
xnor U8759 (N_8759,N_2573,N_80);
or U8760 (N_8760,N_1202,N_794);
or U8761 (N_8761,N_3194,N_3699);
nand U8762 (N_8762,N_2712,N_2826);
nand U8763 (N_8763,N_3872,N_3314);
nand U8764 (N_8764,N_3254,N_2725);
xnor U8765 (N_8765,N_1995,N_4543);
nor U8766 (N_8766,N_2317,N_2301);
xor U8767 (N_8767,N_306,N_3056);
or U8768 (N_8768,N_11,N_1166);
nand U8769 (N_8769,N_3348,N_4507);
nor U8770 (N_8770,N_4106,N_355);
and U8771 (N_8771,N_1655,N_1212);
and U8772 (N_8772,N_576,N_4209);
nand U8773 (N_8773,N_4955,N_3304);
or U8774 (N_8774,N_349,N_210);
nand U8775 (N_8775,N_1015,N_1139);
xor U8776 (N_8776,N_2396,N_1351);
or U8777 (N_8777,N_2279,N_3800);
nor U8778 (N_8778,N_2209,N_3198);
xnor U8779 (N_8779,N_2395,N_4782);
and U8780 (N_8780,N_3232,N_102);
nor U8781 (N_8781,N_2085,N_559);
or U8782 (N_8782,N_4426,N_4288);
nor U8783 (N_8783,N_4717,N_4685);
or U8784 (N_8784,N_4641,N_2275);
and U8785 (N_8785,N_1984,N_3027);
nand U8786 (N_8786,N_2931,N_4646);
xnor U8787 (N_8787,N_4722,N_592);
xor U8788 (N_8788,N_2615,N_3272);
nor U8789 (N_8789,N_450,N_1435);
and U8790 (N_8790,N_2137,N_4226);
and U8791 (N_8791,N_4168,N_4240);
xor U8792 (N_8792,N_836,N_373);
xor U8793 (N_8793,N_2102,N_3111);
and U8794 (N_8794,N_1823,N_2659);
nor U8795 (N_8795,N_4290,N_1995);
nor U8796 (N_8796,N_1373,N_2672);
nand U8797 (N_8797,N_4802,N_2422);
or U8798 (N_8798,N_2279,N_2578);
nor U8799 (N_8799,N_770,N_871);
nor U8800 (N_8800,N_961,N_3447);
xnor U8801 (N_8801,N_1117,N_3984);
and U8802 (N_8802,N_3812,N_229);
xor U8803 (N_8803,N_3345,N_1279);
xor U8804 (N_8804,N_2898,N_914);
nand U8805 (N_8805,N_938,N_3021);
nand U8806 (N_8806,N_4340,N_3104);
or U8807 (N_8807,N_2958,N_198);
nor U8808 (N_8808,N_1328,N_2718);
xnor U8809 (N_8809,N_3144,N_828);
nor U8810 (N_8810,N_2959,N_2492);
nand U8811 (N_8811,N_4726,N_2223);
and U8812 (N_8812,N_1096,N_3541);
nand U8813 (N_8813,N_2171,N_3900);
nand U8814 (N_8814,N_1374,N_4540);
nand U8815 (N_8815,N_1710,N_2928);
xor U8816 (N_8816,N_1322,N_2945);
and U8817 (N_8817,N_242,N_4077);
or U8818 (N_8818,N_1222,N_1543);
and U8819 (N_8819,N_438,N_648);
nor U8820 (N_8820,N_803,N_2849);
nor U8821 (N_8821,N_3609,N_2375);
nand U8822 (N_8822,N_3665,N_1063);
nand U8823 (N_8823,N_329,N_94);
or U8824 (N_8824,N_3045,N_1958);
nor U8825 (N_8825,N_1536,N_1904);
nand U8826 (N_8826,N_188,N_4761);
or U8827 (N_8827,N_4699,N_2530);
nand U8828 (N_8828,N_1706,N_1685);
xnor U8829 (N_8829,N_4501,N_4254);
or U8830 (N_8830,N_4829,N_469);
and U8831 (N_8831,N_1740,N_2654);
nor U8832 (N_8832,N_3381,N_215);
nand U8833 (N_8833,N_2911,N_2775);
and U8834 (N_8834,N_3766,N_3907);
xnor U8835 (N_8835,N_1722,N_4982);
nand U8836 (N_8836,N_4665,N_3108);
nand U8837 (N_8837,N_360,N_2360);
nand U8838 (N_8838,N_4317,N_1257);
nor U8839 (N_8839,N_2153,N_2817);
nand U8840 (N_8840,N_3460,N_4526);
xor U8841 (N_8841,N_923,N_1853);
or U8842 (N_8842,N_4461,N_2813);
nor U8843 (N_8843,N_1496,N_2494);
nand U8844 (N_8844,N_4798,N_1096);
nor U8845 (N_8845,N_263,N_2589);
nand U8846 (N_8846,N_1751,N_1357);
or U8847 (N_8847,N_1187,N_4903);
nor U8848 (N_8848,N_153,N_2332);
nand U8849 (N_8849,N_2700,N_230);
xnor U8850 (N_8850,N_4994,N_976);
and U8851 (N_8851,N_3638,N_2868);
and U8852 (N_8852,N_1332,N_399);
xor U8853 (N_8853,N_2290,N_3990);
xnor U8854 (N_8854,N_2741,N_1388);
xor U8855 (N_8855,N_2825,N_516);
xnor U8856 (N_8856,N_2938,N_2852);
and U8857 (N_8857,N_686,N_2615);
nor U8858 (N_8858,N_1649,N_1560);
and U8859 (N_8859,N_1935,N_1369);
nand U8860 (N_8860,N_3891,N_1860);
xor U8861 (N_8861,N_122,N_4185);
nand U8862 (N_8862,N_2239,N_842);
xnor U8863 (N_8863,N_3119,N_2849);
nand U8864 (N_8864,N_1823,N_418);
xor U8865 (N_8865,N_414,N_348);
nand U8866 (N_8866,N_2981,N_4422);
xor U8867 (N_8867,N_2761,N_4057);
xor U8868 (N_8868,N_139,N_3777);
and U8869 (N_8869,N_1999,N_4735);
or U8870 (N_8870,N_2106,N_3929);
nand U8871 (N_8871,N_1970,N_146);
xnor U8872 (N_8872,N_2058,N_1738);
nand U8873 (N_8873,N_4886,N_1312);
nand U8874 (N_8874,N_2368,N_768);
and U8875 (N_8875,N_178,N_2581);
nor U8876 (N_8876,N_821,N_4428);
xor U8877 (N_8877,N_2304,N_57);
or U8878 (N_8878,N_1372,N_3148);
nand U8879 (N_8879,N_3051,N_1555);
and U8880 (N_8880,N_3596,N_134);
nand U8881 (N_8881,N_4312,N_2704);
nand U8882 (N_8882,N_3728,N_3139);
xor U8883 (N_8883,N_3655,N_4085);
xor U8884 (N_8884,N_1142,N_3083);
or U8885 (N_8885,N_2895,N_3851);
nor U8886 (N_8886,N_3157,N_2372);
nor U8887 (N_8887,N_3586,N_3481);
nand U8888 (N_8888,N_3683,N_21);
or U8889 (N_8889,N_2305,N_3731);
and U8890 (N_8890,N_2925,N_2812);
and U8891 (N_8891,N_149,N_3094);
xnor U8892 (N_8892,N_2063,N_847);
xor U8893 (N_8893,N_3958,N_1206);
or U8894 (N_8894,N_3468,N_4543);
or U8895 (N_8895,N_2905,N_596);
nand U8896 (N_8896,N_2368,N_1178);
or U8897 (N_8897,N_4889,N_2157);
xor U8898 (N_8898,N_1511,N_4292);
nand U8899 (N_8899,N_3929,N_2040);
nand U8900 (N_8900,N_4660,N_1365);
xor U8901 (N_8901,N_3200,N_3364);
xnor U8902 (N_8902,N_2693,N_3362);
nand U8903 (N_8903,N_2187,N_3486);
and U8904 (N_8904,N_1840,N_4775);
nor U8905 (N_8905,N_2408,N_1197);
and U8906 (N_8906,N_3667,N_4809);
nand U8907 (N_8907,N_4910,N_2546);
or U8908 (N_8908,N_2008,N_2017);
nor U8909 (N_8909,N_145,N_4897);
nor U8910 (N_8910,N_555,N_3444);
and U8911 (N_8911,N_3,N_2314);
and U8912 (N_8912,N_4188,N_4123);
nand U8913 (N_8913,N_2300,N_2551);
and U8914 (N_8914,N_2036,N_1103);
or U8915 (N_8915,N_4625,N_1941);
and U8916 (N_8916,N_2944,N_1048);
xnor U8917 (N_8917,N_3171,N_1017);
xor U8918 (N_8918,N_3252,N_2610);
nor U8919 (N_8919,N_545,N_1191);
nand U8920 (N_8920,N_2056,N_2312);
nor U8921 (N_8921,N_1332,N_541);
nand U8922 (N_8922,N_4074,N_311);
nor U8923 (N_8923,N_4276,N_1098);
nand U8924 (N_8924,N_258,N_3894);
xor U8925 (N_8925,N_2025,N_4785);
xnor U8926 (N_8926,N_4894,N_4976);
nor U8927 (N_8927,N_2233,N_4798);
nor U8928 (N_8928,N_3829,N_2468);
nand U8929 (N_8929,N_3991,N_4071);
or U8930 (N_8930,N_805,N_710);
and U8931 (N_8931,N_3654,N_1942);
and U8932 (N_8932,N_1310,N_3466);
and U8933 (N_8933,N_1172,N_4970);
nor U8934 (N_8934,N_2123,N_2953);
or U8935 (N_8935,N_1897,N_2427);
nand U8936 (N_8936,N_3719,N_1115);
nor U8937 (N_8937,N_136,N_2526);
xor U8938 (N_8938,N_873,N_4162);
nor U8939 (N_8939,N_3316,N_705);
xnor U8940 (N_8940,N_4704,N_4145);
nor U8941 (N_8941,N_2684,N_2754);
or U8942 (N_8942,N_1419,N_1209);
nor U8943 (N_8943,N_755,N_3732);
nor U8944 (N_8944,N_4386,N_3586);
xor U8945 (N_8945,N_4776,N_4845);
or U8946 (N_8946,N_2042,N_237);
nor U8947 (N_8947,N_254,N_4683);
xor U8948 (N_8948,N_4613,N_496);
xor U8949 (N_8949,N_4717,N_1808);
nor U8950 (N_8950,N_1663,N_4651);
nand U8951 (N_8951,N_1455,N_3797);
or U8952 (N_8952,N_4258,N_2003);
xnor U8953 (N_8953,N_4708,N_1240);
or U8954 (N_8954,N_4808,N_4322);
or U8955 (N_8955,N_3143,N_717);
nand U8956 (N_8956,N_1724,N_493);
nand U8957 (N_8957,N_4368,N_3567);
nand U8958 (N_8958,N_4775,N_3269);
nor U8959 (N_8959,N_2150,N_1952);
and U8960 (N_8960,N_3276,N_3383);
and U8961 (N_8961,N_203,N_2374);
nor U8962 (N_8962,N_1483,N_852);
nand U8963 (N_8963,N_1421,N_4706);
and U8964 (N_8964,N_4456,N_1924);
and U8965 (N_8965,N_3100,N_4227);
nor U8966 (N_8966,N_3941,N_3448);
and U8967 (N_8967,N_2466,N_3949);
nor U8968 (N_8968,N_1200,N_1436);
or U8969 (N_8969,N_4273,N_3507);
and U8970 (N_8970,N_1697,N_1848);
nand U8971 (N_8971,N_120,N_3434);
and U8972 (N_8972,N_1595,N_2412);
nor U8973 (N_8973,N_472,N_1103);
nand U8974 (N_8974,N_1203,N_997);
or U8975 (N_8975,N_1539,N_528);
and U8976 (N_8976,N_3066,N_3017);
nor U8977 (N_8977,N_3875,N_2137);
nand U8978 (N_8978,N_4431,N_2241);
and U8979 (N_8979,N_1700,N_3142);
nor U8980 (N_8980,N_1720,N_712);
nand U8981 (N_8981,N_4034,N_1005);
xor U8982 (N_8982,N_2699,N_1615);
nor U8983 (N_8983,N_4911,N_3837);
nor U8984 (N_8984,N_2008,N_4078);
xor U8985 (N_8985,N_3142,N_2689);
and U8986 (N_8986,N_4795,N_1419);
nand U8987 (N_8987,N_2781,N_4768);
nand U8988 (N_8988,N_1876,N_727);
and U8989 (N_8989,N_3484,N_2155);
and U8990 (N_8990,N_3543,N_1102);
nand U8991 (N_8991,N_1308,N_3689);
nand U8992 (N_8992,N_4837,N_1850);
or U8993 (N_8993,N_1120,N_2544);
xnor U8994 (N_8994,N_4713,N_4392);
nand U8995 (N_8995,N_759,N_3006);
and U8996 (N_8996,N_3622,N_59);
nor U8997 (N_8997,N_1969,N_940);
xnor U8998 (N_8998,N_1998,N_1729);
xor U8999 (N_8999,N_1250,N_1961);
or U9000 (N_9000,N_4305,N_45);
nand U9001 (N_9001,N_2183,N_4033);
or U9002 (N_9002,N_4171,N_3466);
or U9003 (N_9003,N_3309,N_3065);
and U9004 (N_9004,N_598,N_1638);
or U9005 (N_9005,N_4453,N_1228);
xnor U9006 (N_9006,N_4516,N_726);
nor U9007 (N_9007,N_1098,N_1072);
or U9008 (N_9008,N_4216,N_4232);
or U9009 (N_9009,N_1463,N_2038);
or U9010 (N_9010,N_1423,N_1513);
nand U9011 (N_9011,N_4572,N_635);
nand U9012 (N_9012,N_4140,N_1232);
nor U9013 (N_9013,N_1968,N_685);
xor U9014 (N_9014,N_4854,N_469);
xnor U9015 (N_9015,N_3971,N_3656);
xnor U9016 (N_9016,N_4447,N_1748);
or U9017 (N_9017,N_2638,N_1867);
nor U9018 (N_9018,N_381,N_4270);
xor U9019 (N_9019,N_830,N_1267);
nand U9020 (N_9020,N_125,N_1290);
nor U9021 (N_9021,N_4937,N_2379);
nor U9022 (N_9022,N_3241,N_47);
and U9023 (N_9023,N_3984,N_3351);
nand U9024 (N_9024,N_1044,N_600);
and U9025 (N_9025,N_398,N_3897);
and U9026 (N_9026,N_1233,N_1572);
xor U9027 (N_9027,N_3005,N_1668);
or U9028 (N_9028,N_145,N_246);
and U9029 (N_9029,N_580,N_1986);
and U9030 (N_9030,N_1031,N_3944);
nor U9031 (N_9031,N_4954,N_1736);
or U9032 (N_9032,N_1080,N_4508);
or U9033 (N_9033,N_3462,N_639);
or U9034 (N_9034,N_3601,N_4440);
xor U9035 (N_9035,N_4178,N_4241);
nand U9036 (N_9036,N_108,N_4319);
nand U9037 (N_9037,N_701,N_4416);
xor U9038 (N_9038,N_3024,N_881);
nand U9039 (N_9039,N_3407,N_651);
and U9040 (N_9040,N_500,N_246);
or U9041 (N_9041,N_1316,N_1562);
and U9042 (N_9042,N_2315,N_4184);
nand U9043 (N_9043,N_279,N_3572);
nor U9044 (N_9044,N_1026,N_4135);
nor U9045 (N_9045,N_18,N_19);
nand U9046 (N_9046,N_1888,N_384);
xnor U9047 (N_9047,N_91,N_871);
xor U9048 (N_9048,N_4799,N_4416);
or U9049 (N_9049,N_1732,N_626);
or U9050 (N_9050,N_732,N_2257);
nor U9051 (N_9051,N_2574,N_11);
nor U9052 (N_9052,N_829,N_367);
nand U9053 (N_9053,N_1228,N_2544);
nand U9054 (N_9054,N_1778,N_4132);
nand U9055 (N_9055,N_2881,N_2827);
nand U9056 (N_9056,N_1181,N_4448);
xnor U9057 (N_9057,N_4919,N_3248);
nand U9058 (N_9058,N_3155,N_3822);
nor U9059 (N_9059,N_1692,N_4160);
nand U9060 (N_9060,N_4319,N_1558);
xnor U9061 (N_9061,N_228,N_4486);
and U9062 (N_9062,N_1022,N_1642);
xnor U9063 (N_9063,N_4124,N_4177);
or U9064 (N_9064,N_1501,N_3222);
xnor U9065 (N_9065,N_3980,N_4313);
nand U9066 (N_9066,N_3045,N_2060);
xnor U9067 (N_9067,N_560,N_3689);
and U9068 (N_9068,N_4214,N_124);
xnor U9069 (N_9069,N_4302,N_778);
or U9070 (N_9070,N_2912,N_151);
xnor U9071 (N_9071,N_4769,N_732);
or U9072 (N_9072,N_3723,N_1943);
nand U9073 (N_9073,N_510,N_3402);
nor U9074 (N_9074,N_1851,N_1586);
nor U9075 (N_9075,N_3055,N_1189);
nand U9076 (N_9076,N_3942,N_1759);
xor U9077 (N_9077,N_1507,N_4437);
and U9078 (N_9078,N_1173,N_2801);
nand U9079 (N_9079,N_3893,N_176);
and U9080 (N_9080,N_408,N_1240);
or U9081 (N_9081,N_3930,N_4842);
nand U9082 (N_9082,N_2225,N_2676);
or U9083 (N_9083,N_4046,N_2457);
and U9084 (N_9084,N_1825,N_3080);
and U9085 (N_9085,N_445,N_2487);
nor U9086 (N_9086,N_3324,N_302);
or U9087 (N_9087,N_3769,N_2235);
nand U9088 (N_9088,N_3790,N_2200);
or U9089 (N_9089,N_1146,N_1532);
nor U9090 (N_9090,N_3444,N_980);
or U9091 (N_9091,N_4180,N_3832);
nor U9092 (N_9092,N_2222,N_269);
xnor U9093 (N_9093,N_2561,N_3797);
or U9094 (N_9094,N_2236,N_2113);
nor U9095 (N_9095,N_4928,N_510);
or U9096 (N_9096,N_959,N_3589);
xor U9097 (N_9097,N_1158,N_2773);
or U9098 (N_9098,N_206,N_4426);
nor U9099 (N_9099,N_1362,N_701);
xor U9100 (N_9100,N_3549,N_3995);
or U9101 (N_9101,N_4459,N_717);
and U9102 (N_9102,N_1693,N_1923);
xnor U9103 (N_9103,N_1756,N_2968);
or U9104 (N_9104,N_1631,N_839);
and U9105 (N_9105,N_2768,N_1516);
and U9106 (N_9106,N_4479,N_1051);
xnor U9107 (N_9107,N_42,N_1412);
or U9108 (N_9108,N_126,N_4453);
nand U9109 (N_9109,N_1984,N_4476);
xor U9110 (N_9110,N_345,N_2419);
or U9111 (N_9111,N_4957,N_4049);
xnor U9112 (N_9112,N_4711,N_340);
and U9113 (N_9113,N_3815,N_4137);
nor U9114 (N_9114,N_983,N_2817);
or U9115 (N_9115,N_3250,N_2548);
or U9116 (N_9116,N_330,N_437);
nor U9117 (N_9117,N_3630,N_3343);
xnor U9118 (N_9118,N_4689,N_4581);
nand U9119 (N_9119,N_455,N_2428);
or U9120 (N_9120,N_1362,N_3757);
or U9121 (N_9121,N_818,N_326);
or U9122 (N_9122,N_116,N_4692);
nand U9123 (N_9123,N_579,N_2006);
or U9124 (N_9124,N_4415,N_2457);
nor U9125 (N_9125,N_1386,N_1723);
or U9126 (N_9126,N_540,N_1112);
or U9127 (N_9127,N_4835,N_1162);
nand U9128 (N_9128,N_1027,N_4580);
nand U9129 (N_9129,N_2722,N_2250);
nand U9130 (N_9130,N_1565,N_3673);
and U9131 (N_9131,N_3099,N_3566);
and U9132 (N_9132,N_1815,N_2217);
nand U9133 (N_9133,N_2260,N_4432);
or U9134 (N_9134,N_3480,N_858);
nor U9135 (N_9135,N_402,N_2941);
nand U9136 (N_9136,N_2351,N_1851);
xnor U9137 (N_9137,N_3296,N_1309);
nor U9138 (N_9138,N_2237,N_836);
and U9139 (N_9139,N_3484,N_412);
or U9140 (N_9140,N_4789,N_1493);
or U9141 (N_9141,N_257,N_3838);
nand U9142 (N_9142,N_2762,N_2139);
nor U9143 (N_9143,N_4748,N_3308);
xnor U9144 (N_9144,N_3981,N_2543);
or U9145 (N_9145,N_2838,N_965);
nor U9146 (N_9146,N_4550,N_3001);
or U9147 (N_9147,N_3751,N_608);
nand U9148 (N_9148,N_1183,N_3582);
xor U9149 (N_9149,N_3409,N_499);
and U9150 (N_9150,N_998,N_4696);
nor U9151 (N_9151,N_1723,N_1207);
and U9152 (N_9152,N_2550,N_421);
nand U9153 (N_9153,N_4639,N_3876);
nor U9154 (N_9154,N_1750,N_4046);
nand U9155 (N_9155,N_4745,N_4746);
and U9156 (N_9156,N_1418,N_3669);
nor U9157 (N_9157,N_4234,N_1614);
or U9158 (N_9158,N_3622,N_1143);
nor U9159 (N_9159,N_2187,N_133);
and U9160 (N_9160,N_3797,N_505);
nor U9161 (N_9161,N_2504,N_3063);
nor U9162 (N_9162,N_502,N_3065);
and U9163 (N_9163,N_811,N_3185);
or U9164 (N_9164,N_2885,N_661);
xor U9165 (N_9165,N_1057,N_4502);
nand U9166 (N_9166,N_4155,N_716);
nor U9167 (N_9167,N_4940,N_175);
and U9168 (N_9168,N_1274,N_3747);
or U9169 (N_9169,N_3017,N_352);
nand U9170 (N_9170,N_215,N_1810);
nand U9171 (N_9171,N_4193,N_1102);
xnor U9172 (N_9172,N_4103,N_3674);
nor U9173 (N_9173,N_4233,N_808);
nor U9174 (N_9174,N_563,N_2022);
nor U9175 (N_9175,N_2026,N_4086);
nand U9176 (N_9176,N_2463,N_1429);
or U9177 (N_9177,N_4504,N_2843);
nor U9178 (N_9178,N_73,N_1551);
xor U9179 (N_9179,N_122,N_4792);
xnor U9180 (N_9180,N_2718,N_2481);
nor U9181 (N_9181,N_574,N_462);
nand U9182 (N_9182,N_2281,N_834);
or U9183 (N_9183,N_174,N_3321);
or U9184 (N_9184,N_1263,N_3560);
nand U9185 (N_9185,N_4145,N_1666);
xnor U9186 (N_9186,N_391,N_2123);
xor U9187 (N_9187,N_1571,N_1956);
xor U9188 (N_9188,N_4460,N_1326);
or U9189 (N_9189,N_502,N_4877);
nor U9190 (N_9190,N_1808,N_3456);
xor U9191 (N_9191,N_4596,N_2927);
and U9192 (N_9192,N_1634,N_1018);
or U9193 (N_9193,N_543,N_3530);
xnor U9194 (N_9194,N_3565,N_2688);
or U9195 (N_9195,N_1880,N_572);
and U9196 (N_9196,N_3677,N_2832);
nand U9197 (N_9197,N_984,N_3288);
xnor U9198 (N_9198,N_2121,N_4498);
nor U9199 (N_9199,N_4226,N_195);
or U9200 (N_9200,N_1883,N_2840);
xnor U9201 (N_9201,N_2078,N_4341);
and U9202 (N_9202,N_4099,N_833);
and U9203 (N_9203,N_3726,N_557);
and U9204 (N_9204,N_4777,N_227);
nor U9205 (N_9205,N_4820,N_723);
and U9206 (N_9206,N_1895,N_1114);
or U9207 (N_9207,N_1643,N_208);
and U9208 (N_9208,N_3854,N_1685);
and U9209 (N_9209,N_324,N_3468);
and U9210 (N_9210,N_4095,N_2698);
xor U9211 (N_9211,N_2546,N_2826);
xor U9212 (N_9212,N_4523,N_1557);
nor U9213 (N_9213,N_1780,N_3104);
xor U9214 (N_9214,N_384,N_2179);
xor U9215 (N_9215,N_3821,N_3622);
or U9216 (N_9216,N_924,N_2702);
nand U9217 (N_9217,N_4857,N_4866);
nor U9218 (N_9218,N_1257,N_4030);
xor U9219 (N_9219,N_3663,N_2926);
or U9220 (N_9220,N_3191,N_1842);
nand U9221 (N_9221,N_302,N_205);
nor U9222 (N_9222,N_2645,N_3989);
xnor U9223 (N_9223,N_1986,N_2283);
xnor U9224 (N_9224,N_4557,N_3169);
and U9225 (N_9225,N_1457,N_2448);
or U9226 (N_9226,N_1241,N_857);
nand U9227 (N_9227,N_504,N_4950);
or U9228 (N_9228,N_2123,N_3061);
or U9229 (N_9229,N_841,N_52);
and U9230 (N_9230,N_3659,N_4105);
nor U9231 (N_9231,N_739,N_4140);
or U9232 (N_9232,N_2600,N_2836);
or U9233 (N_9233,N_2462,N_1850);
or U9234 (N_9234,N_896,N_4251);
xor U9235 (N_9235,N_1673,N_1697);
nor U9236 (N_9236,N_200,N_2421);
and U9237 (N_9237,N_3684,N_1806);
xnor U9238 (N_9238,N_4133,N_702);
xor U9239 (N_9239,N_3024,N_2029);
nor U9240 (N_9240,N_2628,N_665);
nand U9241 (N_9241,N_2667,N_2307);
nor U9242 (N_9242,N_2290,N_1139);
nand U9243 (N_9243,N_2216,N_1686);
nor U9244 (N_9244,N_2592,N_3818);
nor U9245 (N_9245,N_3144,N_4925);
xor U9246 (N_9246,N_3006,N_4471);
nand U9247 (N_9247,N_1982,N_3354);
and U9248 (N_9248,N_2357,N_309);
xnor U9249 (N_9249,N_1048,N_512);
nand U9250 (N_9250,N_3034,N_1159);
nor U9251 (N_9251,N_4979,N_1474);
and U9252 (N_9252,N_64,N_4657);
nor U9253 (N_9253,N_581,N_3208);
or U9254 (N_9254,N_2717,N_2487);
nand U9255 (N_9255,N_1814,N_1877);
and U9256 (N_9256,N_3112,N_1871);
nor U9257 (N_9257,N_876,N_1936);
nor U9258 (N_9258,N_2276,N_2694);
xor U9259 (N_9259,N_2069,N_3696);
xor U9260 (N_9260,N_701,N_2019);
xnor U9261 (N_9261,N_1419,N_2113);
xnor U9262 (N_9262,N_2387,N_3480);
xnor U9263 (N_9263,N_2484,N_3641);
and U9264 (N_9264,N_4383,N_2948);
nand U9265 (N_9265,N_2125,N_103);
and U9266 (N_9266,N_4181,N_743);
nand U9267 (N_9267,N_110,N_3827);
and U9268 (N_9268,N_2611,N_2119);
nor U9269 (N_9269,N_227,N_1571);
nor U9270 (N_9270,N_283,N_1596);
nand U9271 (N_9271,N_1755,N_1871);
xnor U9272 (N_9272,N_3142,N_3262);
xnor U9273 (N_9273,N_1835,N_1041);
and U9274 (N_9274,N_4780,N_3069);
or U9275 (N_9275,N_739,N_4553);
and U9276 (N_9276,N_1306,N_982);
and U9277 (N_9277,N_2291,N_2559);
nor U9278 (N_9278,N_1116,N_4749);
nor U9279 (N_9279,N_622,N_4998);
xnor U9280 (N_9280,N_3815,N_4438);
nor U9281 (N_9281,N_1256,N_939);
nand U9282 (N_9282,N_4487,N_713);
nor U9283 (N_9283,N_286,N_380);
or U9284 (N_9284,N_1327,N_3769);
nand U9285 (N_9285,N_4506,N_3777);
and U9286 (N_9286,N_97,N_3957);
nor U9287 (N_9287,N_2643,N_4921);
nor U9288 (N_9288,N_1888,N_3028);
and U9289 (N_9289,N_4175,N_2113);
xnor U9290 (N_9290,N_2436,N_1775);
nand U9291 (N_9291,N_4414,N_2672);
xor U9292 (N_9292,N_1385,N_1634);
nor U9293 (N_9293,N_3873,N_4591);
and U9294 (N_9294,N_1482,N_4087);
or U9295 (N_9295,N_2294,N_4238);
nor U9296 (N_9296,N_2908,N_145);
nor U9297 (N_9297,N_3527,N_2244);
xnor U9298 (N_9298,N_362,N_528);
nor U9299 (N_9299,N_381,N_1353);
nand U9300 (N_9300,N_1700,N_3371);
nand U9301 (N_9301,N_2732,N_4216);
or U9302 (N_9302,N_4459,N_287);
nor U9303 (N_9303,N_2326,N_198);
nand U9304 (N_9304,N_45,N_1053);
nand U9305 (N_9305,N_304,N_4524);
nor U9306 (N_9306,N_3018,N_3675);
nand U9307 (N_9307,N_3628,N_1370);
or U9308 (N_9308,N_4076,N_552);
xor U9309 (N_9309,N_2114,N_3130);
and U9310 (N_9310,N_3029,N_2617);
nand U9311 (N_9311,N_912,N_4081);
nor U9312 (N_9312,N_3113,N_3775);
nand U9313 (N_9313,N_4762,N_1971);
nand U9314 (N_9314,N_163,N_3331);
nor U9315 (N_9315,N_4129,N_4223);
nand U9316 (N_9316,N_719,N_226);
nand U9317 (N_9317,N_3629,N_3684);
or U9318 (N_9318,N_732,N_3465);
and U9319 (N_9319,N_2284,N_348);
or U9320 (N_9320,N_2410,N_2819);
xnor U9321 (N_9321,N_1711,N_850);
nor U9322 (N_9322,N_1788,N_1658);
and U9323 (N_9323,N_1241,N_3246);
and U9324 (N_9324,N_1619,N_4041);
and U9325 (N_9325,N_427,N_3749);
and U9326 (N_9326,N_2238,N_387);
and U9327 (N_9327,N_2467,N_4688);
nor U9328 (N_9328,N_440,N_972);
or U9329 (N_9329,N_4436,N_3717);
nand U9330 (N_9330,N_4420,N_205);
and U9331 (N_9331,N_813,N_1570);
nor U9332 (N_9332,N_1379,N_4826);
xor U9333 (N_9333,N_4587,N_3916);
and U9334 (N_9334,N_4899,N_99);
or U9335 (N_9335,N_2307,N_2640);
or U9336 (N_9336,N_4038,N_2299);
nor U9337 (N_9337,N_3617,N_3321);
or U9338 (N_9338,N_3719,N_4846);
nor U9339 (N_9339,N_2376,N_324);
nand U9340 (N_9340,N_928,N_251);
nand U9341 (N_9341,N_148,N_3178);
or U9342 (N_9342,N_469,N_232);
or U9343 (N_9343,N_4139,N_4921);
or U9344 (N_9344,N_3462,N_1491);
nand U9345 (N_9345,N_1874,N_1616);
or U9346 (N_9346,N_4260,N_4199);
nand U9347 (N_9347,N_953,N_2976);
nand U9348 (N_9348,N_14,N_1481);
xor U9349 (N_9349,N_1263,N_716);
and U9350 (N_9350,N_1818,N_1052);
nor U9351 (N_9351,N_1758,N_622);
xor U9352 (N_9352,N_4678,N_4012);
xor U9353 (N_9353,N_4515,N_837);
or U9354 (N_9354,N_2583,N_1679);
or U9355 (N_9355,N_3626,N_3035);
nand U9356 (N_9356,N_4230,N_4853);
nand U9357 (N_9357,N_2557,N_2492);
and U9358 (N_9358,N_1385,N_4520);
nor U9359 (N_9359,N_563,N_780);
nor U9360 (N_9360,N_2311,N_3834);
and U9361 (N_9361,N_2840,N_2294);
or U9362 (N_9362,N_2601,N_89);
nand U9363 (N_9363,N_4359,N_4493);
nor U9364 (N_9364,N_1362,N_1728);
nand U9365 (N_9365,N_4970,N_992);
and U9366 (N_9366,N_1036,N_3977);
or U9367 (N_9367,N_2566,N_4913);
xor U9368 (N_9368,N_2171,N_1697);
and U9369 (N_9369,N_1214,N_474);
nand U9370 (N_9370,N_1778,N_4660);
xor U9371 (N_9371,N_3487,N_3116);
nor U9372 (N_9372,N_3915,N_4982);
or U9373 (N_9373,N_3090,N_3588);
nand U9374 (N_9374,N_1404,N_176);
nor U9375 (N_9375,N_2315,N_2846);
xor U9376 (N_9376,N_1941,N_3343);
nand U9377 (N_9377,N_702,N_2966);
or U9378 (N_9378,N_2554,N_4586);
nand U9379 (N_9379,N_1916,N_429);
xor U9380 (N_9380,N_4359,N_2619);
or U9381 (N_9381,N_3355,N_2137);
or U9382 (N_9382,N_4162,N_1592);
or U9383 (N_9383,N_4837,N_4424);
and U9384 (N_9384,N_256,N_3524);
nand U9385 (N_9385,N_3172,N_1122);
and U9386 (N_9386,N_2762,N_2898);
and U9387 (N_9387,N_2929,N_3957);
or U9388 (N_9388,N_4627,N_4680);
or U9389 (N_9389,N_2807,N_2140);
xnor U9390 (N_9390,N_3924,N_3406);
xnor U9391 (N_9391,N_1573,N_4881);
nand U9392 (N_9392,N_2163,N_4584);
nand U9393 (N_9393,N_2970,N_1990);
or U9394 (N_9394,N_4481,N_916);
nand U9395 (N_9395,N_2718,N_986);
or U9396 (N_9396,N_2443,N_4129);
and U9397 (N_9397,N_2428,N_1481);
nor U9398 (N_9398,N_719,N_1124);
or U9399 (N_9399,N_1783,N_802);
and U9400 (N_9400,N_4878,N_1425);
or U9401 (N_9401,N_4669,N_758);
nor U9402 (N_9402,N_390,N_351);
nand U9403 (N_9403,N_689,N_942);
or U9404 (N_9404,N_1032,N_1734);
nor U9405 (N_9405,N_1273,N_4450);
xor U9406 (N_9406,N_240,N_3576);
and U9407 (N_9407,N_3715,N_2387);
nor U9408 (N_9408,N_2604,N_509);
and U9409 (N_9409,N_445,N_3603);
nor U9410 (N_9410,N_2221,N_1997);
nand U9411 (N_9411,N_4478,N_980);
or U9412 (N_9412,N_2538,N_4213);
nor U9413 (N_9413,N_2468,N_678);
and U9414 (N_9414,N_1606,N_323);
nor U9415 (N_9415,N_4225,N_2409);
and U9416 (N_9416,N_2911,N_3180);
xor U9417 (N_9417,N_171,N_1832);
nor U9418 (N_9418,N_292,N_1084);
or U9419 (N_9419,N_3426,N_3227);
nor U9420 (N_9420,N_1241,N_475);
and U9421 (N_9421,N_198,N_2131);
nand U9422 (N_9422,N_3082,N_1862);
nor U9423 (N_9423,N_3944,N_83);
nand U9424 (N_9424,N_2050,N_3486);
nor U9425 (N_9425,N_1674,N_1227);
nor U9426 (N_9426,N_4112,N_701);
nor U9427 (N_9427,N_1597,N_2584);
nor U9428 (N_9428,N_637,N_807);
nand U9429 (N_9429,N_2621,N_4576);
nand U9430 (N_9430,N_1964,N_824);
nand U9431 (N_9431,N_56,N_3368);
and U9432 (N_9432,N_133,N_1535);
xor U9433 (N_9433,N_2228,N_2968);
or U9434 (N_9434,N_4809,N_3642);
xor U9435 (N_9435,N_3264,N_387);
and U9436 (N_9436,N_4935,N_954);
or U9437 (N_9437,N_3079,N_1793);
or U9438 (N_9438,N_679,N_815);
or U9439 (N_9439,N_1187,N_4856);
and U9440 (N_9440,N_4429,N_1210);
or U9441 (N_9441,N_4133,N_2300);
or U9442 (N_9442,N_2161,N_568);
nand U9443 (N_9443,N_2759,N_765);
nand U9444 (N_9444,N_1454,N_653);
and U9445 (N_9445,N_1443,N_2878);
nand U9446 (N_9446,N_4199,N_4914);
nand U9447 (N_9447,N_4900,N_4505);
and U9448 (N_9448,N_2521,N_2248);
nor U9449 (N_9449,N_2649,N_3625);
nand U9450 (N_9450,N_4046,N_4983);
or U9451 (N_9451,N_1453,N_3243);
xnor U9452 (N_9452,N_358,N_3356);
nand U9453 (N_9453,N_4488,N_3903);
nor U9454 (N_9454,N_99,N_1419);
nand U9455 (N_9455,N_4330,N_1596);
xor U9456 (N_9456,N_1046,N_1331);
nand U9457 (N_9457,N_1253,N_4200);
xnor U9458 (N_9458,N_4279,N_3988);
or U9459 (N_9459,N_4971,N_951);
or U9460 (N_9460,N_3856,N_4653);
nand U9461 (N_9461,N_4954,N_2588);
and U9462 (N_9462,N_1395,N_4914);
or U9463 (N_9463,N_4786,N_1908);
and U9464 (N_9464,N_4178,N_873);
nand U9465 (N_9465,N_4068,N_4265);
and U9466 (N_9466,N_1842,N_2946);
nor U9467 (N_9467,N_2825,N_617);
xnor U9468 (N_9468,N_4280,N_4391);
xnor U9469 (N_9469,N_2638,N_590);
nand U9470 (N_9470,N_486,N_3288);
xor U9471 (N_9471,N_4633,N_2621);
nand U9472 (N_9472,N_4455,N_2607);
xnor U9473 (N_9473,N_614,N_935);
nand U9474 (N_9474,N_2018,N_4473);
and U9475 (N_9475,N_1788,N_4358);
xnor U9476 (N_9476,N_2098,N_3388);
and U9477 (N_9477,N_2210,N_262);
and U9478 (N_9478,N_2142,N_3711);
or U9479 (N_9479,N_3378,N_2402);
nor U9480 (N_9480,N_2591,N_3915);
nand U9481 (N_9481,N_2744,N_295);
xor U9482 (N_9482,N_3475,N_391);
nor U9483 (N_9483,N_3252,N_4901);
and U9484 (N_9484,N_3807,N_864);
and U9485 (N_9485,N_1421,N_2777);
xor U9486 (N_9486,N_2238,N_1347);
and U9487 (N_9487,N_1823,N_4821);
xnor U9488 (N_9488,N_4408,N_2357);
or U9489 (N_9489,N_244,N_1924);
and U9490 (N_9490,N_785,N_1268);
xor U9491 (N_9491,N_1843,N_4145);
or U9492 (N_9492,N_3234,N_3602);
nor U9493 (N_9493,N_3057,N_443);
nor U9494 (N_9494,N_2786,N_854);
nor U9495 (N_9495,N_1384,N_4917);
or U9496 (N_9496,N_4728,N_3836);
nand U9497 (N_9497,N_2222,N_1386);
and U9498 (N_9498,N_2290,N_3636);
nor U9499 (N_9499,N_4491,N_262);
nand U9500 (N_9500,N_4805,N_2823);
and U9501 (N_9501,N_1422,N_1550);
nor U9502 (N_9502,N_1065,N_1939);
or U9503 (N_9503,N_3656,N_877);
nor U9504 (N_9504,N_1752,N_3785);
nor U9505 (N_9505,N_2411,N_4887);
and U9506 (N_9506,N_157,N_515);
nand U9507 (N_9507,N_974,N_2762);
xor U9508 (N_9508,N_4779,N_906);
nor U9509 (N_9509,N_1693,N_3514);
nand U9510 (N_9510,N_2149,N_2983);
nor U9511 (N_9511,N_4419,N_3702);
nor U9512 (N_9512,N_1922,N_400);
and U9513 (N_9513,N_2600,N_4781);
and U9514 (N_9514,N_2683,N_508);
or U9515 (N_9515,N_4270,N_412);
and U9516 (N_9516,N_4202,N_1279);
nand U9517 (N_9517,N_444,N_2256);
or U9518 (N_9518,N_3273,N_1415);
nor U9519 (N_9519,N_712,N_4531);
or U9520 (N_9520,N_956,N_3981);
nor U9521 (N_9521,N_1298,N_1000);
nor U9522 (N_9522,N_3829,N_3209);
or U9523 (N_9523,N_140,N_410);
xor U9524 (N_9524,N_1372,N_1219);
nand U9525 (N_9525,N_4875,N_1691);
nor U9526 (N_9526,N_3757,N_4405);
or U9527 (N_9527,N_4079,N_1663);
or U9528 (N_9528,N_4295,N_3509);
xor U9529 (N_9529,N_4372,N_4930);
nand U9530 (N_9530,N_3682,N_3717);
nand U9531 (N_9531,N_4935,N_852);
or U9532 (N_9532,N_342,N_2290);
nor U9533 (N_9533,N_2454,N_1714);
xor U9534 (N_9534,N_3920,N_3321);
or U9535 (N_9535,N_1589,N_322);
nand U9536 (N_9536,N_188,N_2503);
nor U9537 (N_9537,N_1132,N_2853);
nand U9538 (N_9538,N_1002,N_1083);
xnor U9539 (N_9539,N_3662,N_1063);
nand U9540 (N_9540,N_3920,N_3045);
or U9541 (N_9541,N_643,N_2484);
or U9542 (N_9542,N_531,N_832);
or U9543 (N_9543,N_2842,N_1979);
and U9544 (N_9544,N_4477,N_448);
nor U9545 (N_9545,N_3484,N_2329);
xnor U9546 (N_9546,N_278,N_3876);
and U9547 (N_9547,N_3997,N_1504);
and U9548 (N_9548,N_4600,N_588);
xnor U9549 (N_9549,N_3168,N_2981);
nand U9550 (N_9550,N_2821,N_3141);
or U9551 (N_9551,N_2703,N_3570);
xor U9552 (N_9552,N_2300,N_2759);
and U9553 (N_9553,N_765,N_3702);
or U9554 (N_9554,N_4481,N_3870);
nor U9555 (N_9555,N_2765,N_3549);
or U9556 (N_9556,N_4660,N_239);
xnor U9557 (N_9557,N_3579,N_4756);
and U9558 (N_9558,N_4089,N_909);
or U9559 (N_9559,N_1720,N_1706);
nor U9560 (N_9560,N_2140,N_3024);
xor U9561 (N_9561,N_1305,N_2058);
and U9562 (N_9562,N_4328,N_688);
and U9563 (N_9563,N_1975,N_4156);
xnor U9564 (N_9564,N_359,N_2786);
or U9565 (N_9565,N_4072,N_2097);
nor U9566 (N_9566,N_4048,N_3788);
nand U9567 (N_9567,N_44,N_1863);
nand U9568 (N_9568,N_1110,N_2003);
nor U9569 (N_9569,N_2007,N_4131);
nor U9570 (N_9570,N_1272,N_3686);
nor U9571 (N_9571,N_2663,N_720);
xnor U9572 (N_9572,N_3190,N_3343);
nand U9573 (N_9573,N_1973,N_1894);
or U9574 (N_9574,N_303,N_2837);
nor U9575 (N_9575,N_4883,N_4059);
nor U9576 (N_9576,N_3006,N_1143);
xor U9577 (N_9577,N_3471,N_1709);
or U9578 (N_9578,N_1021,N_2105);
xnor U9579 (N_9579,N_2168,N_3777);
nor U9580 (N_9580,N_3745,N_2220);
and U9581 (N_9581,N_3746,N_1986);
or U9582 (N_9582,N_1787,N_3763);
xor U9583 (N_9583,N_4058,N_284);
nand U9584 (N_9584,N_4826,N_3688);
or U9585 (N_9585,N_979,N_3292);
nand U9586 (N_9586,N_2750,N_2043);
nor U9587 (N_9587,N_3349,N_4086);
or U9588 (N_9588,N_3273,N_2988);
and U9589 (N_9589,N_1097,N_1330);
nand U9590 (N_9590,N_553,N_2347);
or U9591 (N_9591,N_1656,N_3080);
or U9592 (N_9592,N_1754,N_4570);
and U9593 (N_9593,N_1502,N_3623);
and U9594 (N_9594,N_1572,N_1515);
and U9595 (N_9595,N_469,N_3287);
and U9596 (N_9596,N_4733,N_4966);
xor U9597 (N_9597,N_3138,N_4045);
and U9598 (N_9598,N_3295,N_3120);
nand U9599 (N_9599,N_1179,N_2082);
nand U9600 (N_9600,N_436,N_2834);
or U9601 (N_9601,N_3070,N_1142);
xor U9602 (N_9602,N_1988,N_4419);
nor U9603 (N_9603,N_1355,N_4809);
xor U9604 (N_9604,N_1182,N_1908);
or U9605 (N_9605,N_4368,N_2941);
nand U9606 (N_9606,N_1557,N_1052);
xnor U9607 (N_9607,N_336,N_2208);
and U9608 (N_9608,N_3920,N_2633);
and U9609 (N_9609,N_1488,N_3163);
nand U9610 (N_9610,N_4693,N_1246);
nor U9611 (N_9611,N_490,N_1505);
nor U9612 (N_9612,N_321,N_540);
and U9613 (N_9613,N_73,N_3294);
nor U9614 (N_9614,N_4933,N_4028);
or U9615 (N_9615,N_273,N_4503);
or U9616 (N_9616,N_2327,N_3223);
and U9617 (N_9617,N_3392,N_396);
and U9618 (N_9618,N_499,N_3449);
nand U9619 (N_9619,N_3937,N_2258);
nand U9620 (N_9620,N_4350,N_3204);
nand U9621 (N_9621,N_3700,N_3299);
nor U9622 (N_9622,N_699,N_3626);
nor U9623 (N_9623,N_576,N_957);
or U9624 (N_9624,N_4027,N_2197);
or U9625 (N_9625,N_1395,N_2390);
and U9626 (N_9626,N_101,N_4763);
or U9627 (N_9627,N_1398,N_4192);
or U9628 (N_9628,N_3032,N_4876);
and U9629 (N_9629,N_211,N_1152);
xor U9630 (N_9630,N_2244,N_1218);
nor U9631 (N_9631,N_4330,N_4582);
nand U9632 (N_9632,N_3531,N_1044);
nand U9633 (N_9633,N_393,N_2141);
nor U9634 (N_9634,N_2825,N_1213);
nand U9635 (N_9635,N_3591,N_1572);
and U9636 (N_9636,N_4284,N_1456);
nand U9637 (N_9637,N_187,N_1499);
nor U9638 (N_9638,N_3023,N_449);
or U9639 (N_9639,N_3303,N_654);
xor U9640 (N_9640,N_1316,N_3655);
nand U9641 (N_9641,N_4803,N_4684);
nor U9642 (N_9642,N_3726,N_3769);
xnor U9643 (N_9643,N_2567,N_985);
nand U9644 (N_9644,N_4736,N_695);
or U9645 (N_9645,N_4900,N_2845);
nor U9646 (N_9646,N_2384,N_3179);
xor U9647 (N_9647,N_3824,N_644);
nor U9648 (N_9648,N_3663,N_840);
xor U9649 (N_9649,N_1372,N_3364);
and U9650 (N_9650,N_2540,N_155);
and U9651 (N_9651,N_1574,N_4780);
nand U9652 (N_9652,N_2260,N_3563);
or U9653 (N_9653,N_3121,N_1151);
xor U9654 (N_9654,N_25,N_3866);
or U9655 (N_9655,N_3479,N_4510);
xor U9656 (N_9656,N_2985,N_3941);
or U9657 (N_9657,N_2855,N_4343);
xor U9658 (N_9658,N_2041,N_2078);
and U9659 (N_9659,N_2687,N_3639);
xor U9660 (N_9660,N_4464,N_4811);
or U9661 (N_9661,N_3952,N_1891);
nor U9662 (N_9662,N_745,N_4991);
nor U9663 (N_9663,N_438,N_446);
xnor U9664 (N_9664,N_1502,N_47);
xnor U9665 (N_9665,N_3150,N_1464);
xor U9666 (N_9666,N_2678,N_4641);
nand U9667 (N_9667,N_542,N_2945);
or U9668 (N_9668,N_2850,N_12);
nand U9669 (N_9669,N_2210,N_1955);
and U9670 (N_9670,N_1844,N_2959);
or U9671 (N_9671,N_2272,N_4040);
or U9672 (N_9672,N_1550,N_1065);
or U9673 (N_9673,N_4901,N_1312);
xor U9674 (N_9674,N_3067,N_4110);
xnor U9675 (N_9675,N_3787,N_1871);
or U9676 (N_9676,N_416,N_2479);
nand U9677 (N_9677,N_2801,N_2131);
xor U9678 (N_9678,N_4418,N_1134);
and U9679 (N_9679,N_2738,N_3941);
nand U9680 (N_9680,N_3095,N_274);
and U9681 (N_9681,N_840,N_1840);
and U9682 (N_9682,N_4015,N_2463);
or U9683 (N_9683,N_1206,N_1343);
nand U9684 (N_9684,N_2099,N_883);
nand U9685 (N_9685,N_1906,N_3696);
nor U9686 (N_9686,N_4130,N_1386);
nor U9687 (N_9687,N_1375,N_2516);
or U9688 (N_9688,N_702,N_3899);
xnor U9689 (N_9689,N_3300,N_1004);
nor U9690 (N_9690,N_1384,N_563);
nand U9691 (N_9691,N_669,N_2424);
or U9692 (N_9692,N_261,N_100);
xnor U9693 (N_9693,N_990,N_105);
nor U9694 (N_9694,N_2777,N_77);
xor U9695 (N_9695,N_12,N_2134);
and U9696 (N_9696,N_2620,N_4295);
or U9697 (N_9697,N_1317,N_2592);
nor U9698 (N_9698,N_4834,N_4412);
nand U9699 (N_9699,N_352,N_1337);
nand U9700 (N_9700,N_4540,N_2169);
nor U9701 (N_9701,N_4522,N_1526);
and U9702 (N_9702,N_1862,N_4243);
and U9703 (N_9703,N_3734,N_677);
and U9704 (N_9704,N_1993,N_2199);
xnor U9705 (N_9705,N_3694,N_3583);
and U9706 (N_9706,N_3071,N_2798);
xor U9707 (N_9707,N_3587,N_876);
and U9708 (N_9708,N_3567,N_1936);
and U9709 (N_9709,N_3725,N_4586);
xor U9710 (N_9710,N_2869,N_1914);
nand U9711 (N_9711,N_3012,N_4208);
nand U9712 (N_9712,N_517,N_3187);
xnor U9713 (N_9713,N_316,N_3091);
and U9714 (N_9714,N_3453,N_4868);
nor U9715 (N_9715,N_2444,N_90);
or U9716 (N_9716,N_682,N_3622);
and U9717 (N_9717,N_3701,N_4685);
xnor U9718 (N_9718,N_4087,N_3075);
or U9719 (N_9719,N_582,N_223);
nor U9720 (N_9720,N_4916,N_181);
nand U9721 (N_9721,N_309,N_2386);
or U9722 (N_9722,N_4899,N_2132);
nor U9723 (N_9723,N_27,N_3889);
or U9724 (N_9724,N_619,N_1349);
and U9725 (N_9725,N_1650,N_1051);
nor U9726 (N_9726,N_1669,N_3806);
nor U9727 (N_9727,N_2460,N_3705);
or U9728 (N_9728,N_3188,N_119);
nand U9729 (N_9729,N_635,N_2297);
and U9730 (N_9730,N_1933,N_1310);
or U9731 (N_9731,N_2767,N_988);
and U9732 (N_9732,N_3466,N_4645);
nor U9733 (N_9733,N_3323,N_1521);
nand U9734 (N_9734,N_911,N_3666);
nor U9735 (N_9735,N_2417,N_2971);
and U9736 (N_9736,N_685,N_2403);
nand U9737 (N_9737,N_1020,N_2457);
nor U9738 (N_9738,N_3767,N_1363);
nor U9739 (N_9739,N_2529,N_4626);
nor U9740 (N_9740,N_1804,N_2703);
xnor U9741 (N_9741,N_2215,N_4812);
xor U9742 (N_9742,N_4969,N_2081);
nor U9743 (N_9743,N_1862,N_4320);
and U9744 (N_9744,N_3214,N_4041);
or U9745 (N_9745,N_3744,N_2476);
xor U9746 (N_9746,N_2118,N_2199);
nand U9747 (N_9747,N_2875,N_1292);
nand U9748 (N_9748,N_4541,N_2136);
or U9749 (N_9749,N_1675,N_1397);
nand U9750 (N_9750,N_4159,N_4785);
and U9751 (N_9751,N_3215,N_1310);
and U9752 (N_9752,N_3284,N_1850);
and U9753 (N_9753,N_2378,N_722);
nand U9754 (N_9754,N_4489,N_3491);
and U9755 (N_9755,N_236,N_1083);
nand U9756 (N_9756,N_3947,N_2596);
nor U9757 (N_9757,N_3185,N_2161);
nand U9758 (N_9758,N_3900,N_2055);
and U9759 (N_9759,N_3414,N_3111);
nor U9760 (N_9760,N_4534,N_1976);
nand U9761 (N_9761,N_4447,N_4709);
xnor U9762 (N_9762,N_1397,N_1844);
nor U9763 (N_9763,N_2664,N_1955);
xor U9764 (N_9764,N_2489,N_4325);
xor U9765 (N_9765,N_4402,N_2097);
xnor U9766 (N_9766,N_3629,N_4571);
nor U9767 (N_9767,N_3404,N_1309);
or U9768 (N_9768,N_3306,N_1832);
and U9769 (N_9769,N_1101,N_4187);
xnor U9770 (N_9770,N_3415,N_2859);
and U9771 (N_9771,N_4575,N_3161);
nand U9772 (N_9772,N_2101,N_3762);
xnor U9773 (N_9773,N_2525,N_726);
nand U9774 (N_9774,N_4227,N_4086);
xor U9775 (N_9775,N_3671,N_287);
xor U9776 (N_9776,N_2057,N_4447);
nand U9777 (N_9777,N_2115,N_3861);
or U9778 (N_9778,N_1771,N_4837);
and U9779 (N_9779,N_4374,N_3960);
and U9780 (N_9780,N_2411,N_4001);
nand U9781 (N_9781,N_1603,N_3568);
nor U9782 (N_9782,N_2955,N_2969);
nand U9783 (N_9783,N_3705,N_3095);
or U9784 (N_9784,N_1920,N_4770);
and U9785 (N_9785,N_2840,N_1288);
nor U9786 (N_9786,N_164,N_2159);
or U9787 (N_9787,N_3948,N_3158);
xor U9788 (N_9788,N_3454,N_2766);
and U9789 (N_9789,N_1210,N_3880);
xnor U9790 (N_9790,N_2689,N_2620);
xnor U9791 (N_9791,N_282,N_4942);
nand U9792 (N_9792,N_4691,N_2140);
nor U9793 (N_9793,N_4715,N_528);
and U9794 (N_9794,N_1075,N_3262);
nor U9795 (N_9795,N_4258,N_284);
nor U9796 (N_9796,N_1050,N_654);
nor U9797 (N_9797,N_3290,N_306);
xor U9798 (N_9798,N_10,N_19);
nor U9799 (N_9799,N_2999,N_2876);
nand U9800 (N_9800,N_177,N_3709);
and U9801 (N_9801,N_4082,N_3828);
nand U9802 (N_9802,N_1299,N_1198);
nor U9803 (N_9803,N_254,N_2316);
nor U9804 (N_9804,N_3680,N_952);
nor U9805 (N_9805,N_2208,N_3306);
or U9806 (N_9806,N_4858,N_1042);
nand U9807 (N_9807,N_3084,N_1927);
and U9808 (N_9808,N_1078,N_2393);
and U9809 (N_9809,N_4190,N_4976);
xnor U9810 (N_9810,N_3805,N_579);
nor U9811 (N_9811,N_3168,N_1674);
nor U9812 (N_9812,N_415,N_2150);
nor U9813 (N_9813,N_3128,N_2790);
or U9814 (N_9814,N_675,N_4394);
nor U9815 (N_9815,N_3873,N_2868);
nor U9816 (N_9816,N_4263,N_186);
and U9817 (N_9817,N_1037,N_1679);
and U9818 (N_9818,N_1359,N_2009);
xnor U9819 (N_9819,N_116,N_1016);
and U9820 (N_9820,N_2813,N_2893);
and U9821 (N_9821,N_1627,N_1898);
and U9822 (N_9822,N_122,N_333);
nor U9823 (N_9823,N_641,N_3253);
or U9824 (N_9824,N_622,N_1076);
or U9825 (N_9825,N_2487,N_3229);
nor U9826 (N_9826,N_1951,N_1957);
and U9827 (N_9827,N_4556,N_4292);
nor U9828 (N_9828,N_124,N_1979);
and U9829 (N_9829,N_70,N_3706);
nand U9830 (N_9830,N_2467,N_3857);
and U9831 (N_9831,N_4682,N_2624);
nand U9832 (N_9832,N_112,N_2583);
or U9833 (N_9833,N_1077,N_119);
or U9834 (N_9834,N_805,N_1317);
nand U9835 (N_9835,N_821,N_1441);
xnor U9836 (N_9836,N_868,N_4044);
and U9837 (N_9837,N_2195,N_1173);
and U9838 (N_9838,N_1105,N_4958);
xor U9839 (N_9839,N_1339,N_1368);
nor U9840 (N_9840,N_1013,N_4295);
nand U9841 (N_9841,N_4513,N_1309);
nand U9842 (N_9842,N_3392,N_2390);
nand U9843 (N_9843,N_4361,N_743);
nand U9844 (N_9844,N_555,N_684);
xor U9845 (N_9845,N_651,N_2731);
xor U9846 (N_9846,N_4698,N_2338);
nand U9847 (N_9847,N_1071,N_991);
nor U9848 (N_9848,N_437,N_160);
xor U9849 (N_9849,N_3513,N_1828);
or U9850 (N_9850,N_2066,N_1955);
or U9851 (N_9851,N_3212,N_378);
or U9852 (N_9852,N_4272,N_3978);
nand U9853 (N_9853,N_3118,N_4765);
xnor U9854 (N_9854,N_1990,N_268);
xnor U9855 (N_9855,N_3574,N_2503);
nor U9856 (N_9856,N_1148,N_3903);
and U9857 (N_9857,N_1829,N_1620);
xor U9858 (N_9858,N_314,N_2657);
or U9859 (N_9859,N_460,N_3367);
xnor U9860 (N_9860,N_3232,N_1340);
xor U9861 (N_9861,N_983,N_2233);
and U9862 (N_9862,N_3411,N_2583);
xor U9863 (N_9863,N_1579,N_686);
nor U9864 (N_9864,N_2164,N_2284);
nand U9865 (N_9865,N_740,N_1506);
xor U9866 (N_9866,N_3634,N_3548);
xnor U9867 (N_9867,N_989,N_3564);
nor U9868 (N_9868,N_2431,N_3112);
and U9869 (N_9869,N_3698,N_2990);
nor U9870 (N_9870,N_1646,N_2036);
nor U9871 (N_9871,N_593,N_2486);
nand U9872 (N_9872,N_1254,N_3741);
nand U9873 (N_9873,N_2669,N_4521);
nand U9874 (N_9874,N_2582,N_3387);
nand U9875 (N_9875,N_3718,N_2067);
xor U9876 (N_9876,N_625,N_496);
nor U9877 (N_9877,N_4200,N_3125);
and U9878 (N_9878,N_1483,N_2795);
nand U9879 (N_9879,N_2134,N_3996);
nor U9880 (N_9880,N_4254,N_4401);
nor U9881 (N_9881,N_1784,N_3198);
xnor U9882 (N_9882,N_155,N_3742);
xor U9883 (N_9883,N_1583,N_311);
and U9884 (N_9884,N_1078,N_2331);
nand U9885 (N_9885,N_483,N_2588);
or U9886 (N_9886,N_743,N_4641);
and U9887 (N_9887,N_2575,N_2673);
and U9888 (N_9888,N_3398,N_1618);
nor U9889 (N_9889,N_2964,N_3367);
or U9890 (N_9890,N_3792,N_2080);
or U9891 (N_9891,N_1905,N_778);
or U9892 (N_9892,N_285,N_3197);
nor U9893 (N_9893,N_4287,N_4555);
nand U9894 (N_9894,N_3466,N_2306);
nand U9895 (N_9895,N_3728,N_625);
or U9896 (N_9896,N_1936,N_353);
nand U9897 (N_9897,N_1435,N_2930);
or U9898 (N_9898,N_354,N_2568);
and U9899 (N_9899,N_1065,N_4364);
or U9900 (N_9900,N_2952,N_2729);
xnor U9901 (N_9901,N_3294,N_2101);
nor U9902 (N_9902,N_1862,N_4104);
nor U9903 (N_9903,N_559,N_2603);
nor U9904 (N_9904,N_3470,N_4030);
or U9905 (N_9905,N_2135,N_3698);
nor U9906 (N_9906,N_3692,N_3465);
or U9907 (N_9907,N_1828,N_4378);
nor U9908 (N_9908,N_601,N_1704);
or U9909 (N_9909,N_4117,N_1703);
xor U9910 (N_9910,N_3215,N_4721);
nand U9911 (N_9911,N_2349,N_4380);
and U9912 (N_9912,N_3300,N_4458);
xnor U9913 (N_9913,N_3800,N_2931);
and U9914 (N_9914,N_2647,N_4087);
nand U9915 (N_9915,N_1898,N_1651);
and U9916 (N_9916,N_1431,N_1312);
or U9917 (N_9917,N_3052,N_4120);
nand U9918 (N_9918,N_2392,N_3649);
or U9919 (N_9919,N_3097,N_2558);
or U9920 (N_9920,N_4621,N_4516);
xor U9921 (N_9921,N_2416,N_1417);
and U9922 (N_9922,N_1223,N_973);
xnor U9923 (N_9923,N_2946,N_79);
nor U9924 (N_9924,N_3749,N_3389);
nor U9925 (N_9925,N_2372,N_1113);
nor U9926 (N_9926,N_2204,N_446);
or U9927 (N_9927,N_347,N_2016);
nand U9928 (N_9928,N_1958,N_1596);
nor U9929 (N_9929,N_4070,N_198);
nand U9930 (N_9930,N_3422,N_64);
xnor U9931 (N_9931,N_3911,N_4830);
nand U9932 (N_9932,N_4235,N_2215);
nand U9933 (N_9933,N_660,N_261);
and U9934 (N_9934,N_1543,N_753);
xor U9935 (N_9935,N_1732,N_4972);
and U9936 (N_9936,N_4227,N_2181);
nor U9937 (N_9937,N_1260,N_2815);
and U9938 (N_9938,N_2248,N_334);
or U9939 (N_9939,N_4186,N_1378);
nor U9940 (N_9940,N_2187,N_4425);
nor U9941 (N_9941,N_4041,N_1983);
xnor U9942 (N_9942,N_2739,N_4863);
nor U9943 (N_9943,N_3607,N_3905);
or U9944 (N_9944,N_274,N_2872);
nand U9945 (N_9945,N_4802,N_1045);
and U9946 (N_9946,N_811,N_4206);
or U9947 (N_9947,N_2389,N_898);
nor U9948 (N_9948,N_2499,N_3345);
nand U9949 (N_9949,N_1363,N_4744);
and U9950 (N_9950,N_4068,N_1706);
and U9951 (N_9951,N_1878,N_2605);
nand U9952 (N_9952,N_3358,N_2236);
xnor U9953 (N_9953,N_1755,N_2126);
xor U9954 (N_9954,N_580,N_96);
nand U9955 (N_9955,N_405,N_4345);
nor U9956 (N_9956,N_4187,N_3700);
or U9957 (N_9957,N_455,N_70);
xor U9958 (N_9958,N_3856,N_338);
nor U9959 (N_9959,N_2765,N_4783);
nor U9960 (N_9960,N_4719,N_1618);
and U9961 (N_9961,N_1582,N_4006);
and U9962 (N_9962,N_2145,N_1678);
nand U9963 (N_9963,N_3830,N_2620);
nor U9964 (N_9964,N_414,N_1608);
nand U9965 (N_9965,N_2457,N_2656);
nor U9966 (N_9966,N_3235,N_3216);
nand U9967 (N_9967,N_4167,N_3838);
xnor U9968 (N_9968,N_70,N_2733);
xnor U9969 (N_9969,N_1505,N_4081);
nand U9970 (N_9970,N_4190,N_3308);
nand U9971 (N_9971,N_3279,N_2876);
xnor U9972 (N_9972,N_2316,N_2944);
and U9973 (N_9973,N_1079,N_3314);
nor U9974 (N_9974,N_3962,N_2934);
nor U9975 (N_9975,N_3266,N_2085);
nand U9976 (N_9976,N_1728,N_3434);
nor U9977 (N_9977,N_2820,N_3824);
and U9978 (N_9978,N_1929,N_556);
nand U9979 (N_9979,N_1525,N_187);
nor U9980 (N_9980,N_4779,N_2669);
or U9981 (N_9981,N_1957,N_346);
xnor U9982 (N_9982,N_2834,N_1369);
nor U9983 (N_9983,N_306,N_3617);
and U9984 (N_9984,N_1815,N_1382);
or U9985 (N_9985,N_1893,N_1374);
nor U9986 (N_9986,N_716,N_3051);
nor U9987 (N_9987,N_2454,N_889);
nor U9988 (N_9988,N_4829,N_1677);
nor U9989 (N_9989,N_3217,N_35);
or U9990 (N_9990,N_459,N_243);
nor U9991 (N_9991,N_2352,N_3644);
and U9992 (N_9992,N_2617,N_1095);
nor U9993 (N_9993,N_846,N_1247);
or U9994 (N_9994,N_3150,N_2323);
xor U9995 (N_9995,N_3945,N_1385);
or U9996 (N_9996,N_4276,N_4237);
nand U9997 (N_9997,N_3969,N_2092);
xor U9998 (N_9998,N_1252,N_1059);
nor U9999 (N_9999,N_168,N_163);
and U10000 (N_10000,N_7974,N_6758);
and U10001 (N_10001,N_6086,N_9003);
nand U10002 (N_10002,N_7833,N_5771);
or U10003 (N_10003,N_8291,N_5088);
or U10004 (N_10004,N_5787,N_9563);
and U10005 (N_10005,N_7274,N_8538);
xor U10006 (N_10006,N_7103,N_7104);
or U10007 (N_10007,N_8822,N_7767);
or U10008 (N_10008,N_5079,N_6637);
or U10009 (N_10009,N_8287,N_9217);
nor U10010 (N_10010,N_5255,N_9363);
nand U10011 (N_10011,N_5448,N_7878);
nor U10012 (N_10012,N_9227,N_6652);
and U10013 (N_10013,N_9863,N_6610);
or U10014 (N_10014,N_8776,N_8999);
xnor U10015 (N_10015,N_6779,N_7025);
nand U10016 (N_10016,N_6916,N_8199);
nor U10017 (N_10017,N_6935,N_7150);
xor U10018 (N_10018,N_6231,N_9135);
nand U10019 (N_10019,N_5366,N_9359);
xor U10020 (N_10020,N_6100,N_9407);
or U10021 (N_10021,N_9914,N_8642);
nand U10022 (N_10022,N_5725,N_8553);
nand U10023 (N_10023,N_8187,N_7163);
and U10024 (N_10024,N_6039,N_5617);
and U10025 (N_10025,N_6495,N_8406);
nand U10026 (N_10026,N_8953,N_8340);
nand U10027 (N_10027,N_6256,N_9674);
or U10028 (N_10028,N_7648,N_7331);
nor U10029 (N_10029,N_7691,N_9970);
nor U10030 (N_10030,N_7529,N_9822);
nand U10031 (N_10031,N_7665,N_5230);
nand U10032 (N_10032,N_5963,N_9019);
nand U10033 (N_10033,N_9634,N_7569);
and U10034 (N_10034,N_8013,N_6529);
nand U10035 (N_10035,N_5349,N_7637);
or U10036 (N_10036,N_6463,N_6456);
nor U10037 (N_10037,N_7987,N_6931);
and U10038 (N_10038,N_5822,N_6295);
xnor U10039 (N_10039,N_5799,N_7587);
and U10040 (N_10040,N_6775,N_6627);
xor U10041 (N_10041,N_6405,N_9628);
xor U10042 (N_10042,N_8587,N_9740);
nor U10043 (N_10043,N_6820,N_5834);
and U10044 (N_10044,N_9859,N_7690);
nor U10045 (N_10045,N_6066,N_9259);
and U10046 (N_10046,N_6867,N_6869);
or U10047 (N_10047,N_9757,N_7593);
xor U10048 (N_10048,N_7774,N_6299);
nor U10049 (N_10049,N_9408,N_8629);
and U10050 (N_10050,N_7432,N_5999);
nor U10051 (N_10051,N_6265,N_9044);
or U10052 (N_10052,N_7280,N_8096);
and U10053 (N_10053,N_5836,N_7629);
or U10054 (N_10054,N_9930,N_5750);
or U10055 (N_10055,N_6785,N_6467);
nor U10056 (N_10056,N_7936,N_9738);
nor U10057 (N_10057,N_6719,N_8636);
nand U10058 (N_10058,N_6959,N_5876);
nor U10059 (N_10059,N_5428,N_8547);
nor U10060 (N_10060,N_9775,N_9643);
or U10061 (N_10061,N_9857,N_9815);
or U10062 (N_10062,N_9239,N_9426);
nor U10063 (N_10063,N_5134,N_5371);
xor U10064 (N_10064,N_5344,N_5036);
xor U10065 (N_10065,N_8328,N_9031);
nor U10066 (N_10066,N_9229,N_6502);
and U10067 (N_10067,N_8853,N_9152);
xnor U10068 (N_10068,N_8749,N_6626);
nand U10069 (N_10069,N_5003,N_5757);
and U10070 (N_10070,N_5130,N_7447);
or U10071 (N_10071,N_9734,N_5141);
and U10072 (N_10072,N_6648,N_8552);
xnor U10073 (N_10073,N_7430,N_5090);
or U10074 (N_10074,N_7760,N_7326);
xnor U10075 (N_10075,N_5866,N_6134);
and U10076 (N_10076,N_9209,N_7585);
nand U10077 (N_10077,N_6499,N_5156);
nor U10078 (N_10078,N_7316,N_7823);
nor U10079 (N_10079,N_9824,N_5826);
xor U10080 (N_10080,N_6001,N_9526);
xor U10081 (N_10081,N_7088,N_7337);
nor U10082 (N_10082,N_7887,N_5839);
and U10083 (N_10083,N_6702,N_6455);
or U10084 (N_10084,N_7941,N_6669);
or U10085 (N_10085,N_5780,N_8438);
xnor U10086 (N_10086,N_6382,N_8067);
xnor U10087 (N_10087,N_6107,N_8489);
and U10088 (N_10088,N_6907,N_5560);
or U10089 (N_10089,N_9186,N_6171);
and U10090 (N_10090,N_7804,N_7758);
nor U10091 (N_10091,N_9940,N_5621);
xnor U10092 (N_10092,N_5557,N_7141);
and U10093 (N_10093,N_7661,N_9184);
nand U10094 (N_10094,N_9461,N_6806);
nand U10095 (N_10095,N_9870,N_5018);
and U10096 (N_10096,N_8493,N_9877);
and U10097 (N_10097,N_9187,N_8167);
nor U10098 (N_10098,N_7342,N_9228);
or U10099 (N_10099,N_9385,N_6187);
xnor U10100 (N_10100,N_5360,N_6255);
nand U10101 (N_10101,N_5118,N_5584);
and U10102 (N_10102,N_9942,N_7858);
nand U10103 (N_10103,N_7543,N_8522);
xor U10104 (N_10104,N_5934,N_8481);
and U10105 (N_10105,N_9502,N_5631);
xnor U10106 (N_10106,N_8665,N_6164);
xor U10107 (N_10107,N_8325,N_8490);
nor U10108 (N_10108,N_7513,N_7492);
xor U10109 (N_10109,N_9320,N_7656);
nor U10110 (N_10110,N_5583,N_7605);
or U10111 (N_10111,N_8381,N_8673);
or U10112 (N_10112,N_8075,N_6248);
nand U10113 (N_10113,N_8689,N_9376);
and U10114 (N_10114,N_9979,N_6423);
nand U10115 (N_10115,N_6461,N_9021);
xnor U10116 (N_10116,N_7098,N_8919);
or U10117 (N_10117,N_5345,N_8379);
and U10118 (N_10118,N_9189,N_9934);
xnor U10119 (N_10119,N_7784,N_7195);
and U10120 (N_10120,N_8889,N_6366);
or U10121 (N_10121,N_8635,N_7654);
or U10122 (N_10122,N_7642,N_5127);
and U10123 (N_10123,N_6170,N_6061);
and U10124 (N_10124,N_7759,N_9590);
nor U10125 (N_10125,N_5745,N_8375);
and U10126 (N_10126,N_9527,N_5949);
nand U10127 (N_10127,N_8281,N_7478);
xnor U10128 (N_10128,N_7053,N_5146);
or U10129 (N_10129,N_6080,N_6359);
or U10130 (N_10130,N_5234,N_5388);
or U10131 (N_10131,N_5320,N_5927);
xor U10132 (N_10132,N_8781,N_8904);
xnor U10133 (N_10133,N_8404,N_5911);
or U10134 (N_10134,N_5660,N_6571);
nor U10135 (N_10135,N_5417,N_5887);
nor U10136 (N_10136,N_8832,N_5033);
xor U10137 (N_10137,N_9725,N_9507);
or U10138 (N_10138,N_9196,N_6215);
nor U10139 (N_10139,N_6432,N_7567);
nor U10140 (N_10140,N_5521,N_8345);
and U10141 (N_10141,N_5206,N_6951);
nand U10142 (N_10142,N_8194,N_8690);
and U10143 (N_10143,N_9467,N_7322);
xnor U10144 (N_10144,N_6832,N_6524);
or U10145 (N_10145,N_9396,N_7835);
or U10146 (N_10146,N_5465,N_9962);
nand U10147 (N_10147,N_8871,N_9872);
and U10148 (N_10148,N_7364,N_9112);
and U10149 (N_10149,N_9419,N_8606);
or U10150 (N_10150,N_6056,N_5095);
or U10151 (N_10151,N_9283,N_7323);
nor U10152 (N_10152,N_9749,N_5284);
nand U10153 (N_10153,N_8311,N_6106);
and U10154 (N_10154,N_8257,N_6605);
nand U10155 (N_10155,N_7057,N_5113);
xor U10156 (N_10156,N_8405,N_8136);
or U10157 (N_10157,N_9190,N_9456);
nor U10158 (N_10158,N_9572,N_9805);
or U10159 (N_10159,N_9398,N_7624);
or U10160 (N_10160,N_5019,N_6530);
nor U10161 (N_10161,N_5845,N_9618);
xor U10162 (N_10162,N_5274,N_6378);
nor U10163 (N_10163,N_7789,N_6546);
or U10164 (N_10164,N_8260,N_6857);
and U10165 (N_10165,N_6837,N_7837);
xor U10166 (N_10166,N_5442,N_6846);
nor U10167 (N_10167,N_8982,N_7501);
xor U10168 (N_10168,N_8693,N_6308);
or U10169 (N_10169,N_8223,N_6969);
and U10170 (N_10170,N_8903,N_5756);
nand U10171 (N_10171,N_7806,N_5155);
nand U10172 (N_10172,N_6263,N_7639);
xor U10173 (N_10173,N_9214,N_8019);
xor U10174 (N_10174,N_6173,N_9339);
or U10175 (N_10175,N_8495,N_5886);
nor U10176 (N_10176,N_6264,N_9620);
or U10177 (N_10177,N_6487,N_6884);
nand U10178 (N_10178,N_5053,N_7045);
nor U10179 (N_10179,N_8265,N_5636);
or U10180 (N_10180,N_8429,N_9171);
or U10181 (N_10181,N_9867,N_6576);
nand U10182 (N_10182,N_7657,N_7695);
nor U10183 (N_10183,N_6688,N_7776);
and U10184 (N_10184,N_8372,N_8051);
nor U10185 (N_10185,N_8302,N_6179);
nand U10186 (N_10186,N_7829,N_6595);
nand U10187 (N_10187,N_9163,N_5035);
xnor U10188 (N_10188,N_7590,N_6735);
and U10189 (N_10189,N_9841,N_6876);
nor U10190 (N_10190,N_7295,N_7237);
or U10191 (N_10191,N_8980,N_9838);
nand U10192 (N_10192,N_5433,N_5299);
or U10193 (N_10193,N_6518,N_6780);
xnor U10194 (N_10194,N_6193,N_9348);
and U10195 (N_10195,N_5768,N_8702);
or U10196 (N_10196,N_6982,N_8173);
nand U10197 (N_10197,N_8185,N_5312);
nand U10198 (N_10198,N_9501,N_6994);
xor U10199 (N_10199,N_6866,N_9933);
nand U10200 (N_10200,N_6352,N_6078);
and U10201 (N_10201,N_5806,N_5403);
xnor U10202 (N_10202,N_7007,N_5435);
nor U10203 (N_10203,N_6533,N_7959);
nand U10204 (N_10204,N_8143,N_8058);
nor U10205 (N_10205,N_7966,N_9974);
and U10206 (N_10206,N_6508,N_8261);
nor U10207 (N_10207,N_9847,N_8626);
nand U10208 (N_10208,N_7768,N_7166);
or U10209 (N_10209,N_7079,N_7292);
and U10210 (N_10210,N_6137,N_7105);
and U10211 (N_10211,N_8534,N_8551);
xnor U10212 (N_10212,N_8157,N_8681);
nand U10213 (N_10213,N_6678,N_8246);
nor U10214 (N_10214,N_6076,N_5577);
and U10215 (N_10215,N_5407,N_5050);
or U10216 (N_10216,N_6680,N_8488);
nand U10217 (N_10217,N_9213,N_7973);
and U10218 (N_10218,N_9913,N_8807);
nand U10219 (N_10219,N_8451,N_9335);
nand U10220 (N_10220,N_9002,N_9834);
nor U10221 (N_10221,N_6276,N_9635);
or U10222 (N_10222,N_5591,N_9980);
nand U10223 (N_10223,N_9731,N_8231);
nand U10224 (N_10224,N_9918,N_9420);
xor U10225 (N_10225,N_8559,N_7508);
nand U10226 (N_10226,N_7390,N_6438);
nand U10227 (N_10227,N_7728,N_8274);
or U10228 (N_10228,N_5147,N_5894);
and U10229 (N_10229,N_9140,N_9085);
xor U10230 (N_10230,N_5182,N_9515);
xor U10231 (N_10231,N_7557,N_6286);
and U10232 (N_10232,N_9036,N_9800);
nor U10233 (N_10233,N_7155,N_5165);
or U10234 (N_10234,N_5653,N_7922);
and U10235 (N_10235,N_8242,N_5792);
or U10236 (N_10236,N_9089,N_5703);
nor U10237 (N_10237,N_6828,N_5655);
nor U10238 (N_10238,N_8097,N_7377);
and U10239 (N_10239,N_5717,N_9772);
nand U10240 (N_10240,N_9964,N_7033);
nor U10241 (N_10241,N_5821,N_6506);
nor U10242 (N_10242,N_6548,N_9384);
nor U10243 (N_10243,N_8047,N_8384);
nand U10244 (N_10244,N_7477,N_8508);
or U10245 (N_10245,N_6048,N_9886);
nand U10246 (N_10246,N_9803,N_7903);
nand U10247 (N_10247,N_9144,N_9009);
and U10248 (N_10248,N_8332,N_9516);
and U10249 (N_10249,N_6676,N_9448);
or U10250 (N_10250,N_5023,N_7867);
nand U10251 (N_10251,N_7138,N_6617);
xnor U10252 (N_10252,N_8358,N_6363);
nand U10253 (N_10253,N_9078,N_7882);
or U10254 (N_10254,N_5900,N_8675);
or U10255 (N_10255,N_6253,N_8144);
or U10256 (N_10256,N_9433,N_7325);
nand U10257 (N_10257,N_5315,N_8149);
or U10258 (N_10258,N_9613,N_5455);
nor U10259 (N_10259,N_7625,N_8282);
and U10260 (N_10260,N_8401,N_7311);
nor U10261 (N_10261,N_7032,N_7533);
and U10262 (N_10262,N_5612,N_5695);
or U10263 (N_10263,N_5322,N_6872);
and U10264 (N_10264,N_9603,N_8370);
or U10265 (N_10265,N_5982,N_7180);
nor U10266 (N_10266,N_8373,N_6894);
nand U10267 (N_10267,N_6118,N_7121);
xor U10268 (N_10268,N_9959,N_7069);
xor U10269 (N_10269,N_9608,N_9538);
and U10270 (N_10270,N_8132,N_6975);
or U10271 (N_10271,N_5863,N_6609);
nand U10272 (N_10272,N_8813,N_8172);
xnor U10273 (N_10273,N_7741,N_6621);
nor U10274 (N_10274,N_7238,N_9948);
and U10275 (N_10275,N_6099,N_9733);
xor U10276 (N_10276,N_7128,N_5712);
or U10277 (N_10277,N_7821,N_9394);
xnor U10278 (N_10278,N_6447,N_6004);
or U10279 (N_10279,N_7608,N_5872);
xnor U10280 (N_10280,N_5766,N_7927);
or U10281 (N_10281,N_5161,N_6221);
xnor U10282 (N_10282,N_7798,N_8946);
or U10283 (N_10283,N_9016,N_8119);
nor U10284 (N_10284,N_6824,N_9779);
or U10285 (N_10285,N_5990,N_7114);
xnor U10286 (N_10286,N_9636,N_9529);
nor U10287 (N_10287,N_7341,N_5292);
nand U10288 (N_10288,N_7490,N_9550);
nand U10289 (N_10289,N_5646,N_7015);
nor U10290 (N_10290,N_9615,N_7000);
nand U10291 (N_10291,N_8494,N_8687);
nand U10292 (N_10292,N_7822,N_7439);
and U10293 (N_10293,N_9514,N_7431);
xnor U10294 (N_10294,N_8855,N_9377);
and U10295 (N_10295,N_6880,N_6055);
nor U10296 (N_10296,N_7947,N_7801);
or U10297 (N_10297,N_9505,N_5784);
or U10298 (N_10298,N_6968,N_5965);
nand U10299 (N_10299,N_8951,N_6732);
and U10300 (N_10300,N_9764,N_9937);
nand U10301 (N_10301,N_8485,N_6274);
xnor U10302 (N_10302,N_7363,N_8351);
nand U10303 (N_10303,N_8934,N_5150);
nand U10304 (N_10304,N_8976,N_5993);
or U10305 (N_10305,N_9640,N_9205);
and U10306 (N_10306,N_5499,N_9885);
nand U10307 (N_10307,N_7860,N_6802);
xnor U10308 (N_10308,N_6864,N_7827);
and U10309 (N_10309,N_9434,N_9273);
xor U10310 (N_10310,N_8471,N_8837);
and U10311 (N_10311,N_7350,N_5481);
nand U10312 (N_10312,N_7153,N_8441);
nor U10313 (N_10313,N_9455,N_9288);
nor U10314 (N_10314,N_5539,N_7064);
nor U10315 (N_10315,N_9825,N_8195);
xor U10316 (N_10316,N_6348,N_6521);
nand U10317 (N_10317,N_5825,N_7997);
xor U10318 (N_10318,N_9821,N_8222);
and U10319 (N_10319,N_9090,N_8997);
nand U10320 (N_10320,N_5446,N_7913);
and U10321 (N_10321,N_9369,N_7006);
nor U10322 (N_10322,N_9921,N_9292);
xor U10323 (N_10323,N_8483,N_6835);
or U10324 (N_10324,N_5045,N_8397);
or U10325 (N_10325,N_8700,N_7960);
and U10326 (N_10326,N_9837,N_6181);
or U10327 (N_10327,N_6769,N_6191);
nand U10328 (N_10328,N_8437,N_6199);
or U10329 (N_10329,N_6953,N_8521);
nand U10330 (N_10330,N_5697,N_7883);
xnor U10331 (N_10331,N_9416,N_5729);
nand U10332 (N_10332,N_6040,N_6765);
nor U10333 (N_10333,N_8634,N_6910);
nand U10334 (N_10334,N_9097,N_6756);
or U10335 (N_10335,N_8528,N_8150);
and U10336 (N_10336,N_7879,N_8304);
or U10337 (N_10337,N_7736,N_7825);
or U10338 (N_10338,N_9606,N_9030);
xnor U10339 (N_10339,N_5237,N_5008);
and U10340 (N_10340,N_5754,N_7761);
or U10341 (N_10341,N_9498,N_5589);
and U10342 (N_10342,N_8270,N_9994);
nor U10343 (N_10343,N_6511,N_5270);
nor U10344 (N_10344,N_5250,N_5992);
nor U10345 (N_10345,N_7715,N_7888);
nor U10346 (N_10346,N_9043,N_5313);
and U10347 (N_10347,N_8505,N_7034);
or U10348 (N_10348,N_8960,N_9765);
and U10349 (N_10349,N_5260,N_5289);
nor U10350 (N_10350,N_9565,N_7227);
xor U10351 (N_10351,N_8734,N_7132);
nand U10352 (N_10352,N_5476,N_8446);
xnor U10353 (N_10353,N_5281,N_8891);
and U10354 (N_10354,N_9793,N_9176);
nand U10355 (N_10355,N_8497,N_5651);
nand U10356 (N_10356,N_7159,N_8956);
nand U10357 (N_10357,N_5229,N_6887);
nand U10358 (N_10358,N_5807,N_8517);
nand U10359 (N_10359,N_5397,N_9074);
xor U10360 (N_10360,N_8879,N_7535);
nand U10361 (N_10361,N_6033,N_6836);
and U10362 (N_10362,N_5325,N_6358);
and U10363 (N_10363,N_5464,N_9548);
xor U10364 (N_10364,N_5994,N_6573);
or U10365 (N_10365,N_7359,N_9549);
nor U10366 (N_10366,N_6023,N_8276);
or U10367 (N_10367,N_9272,N_6068);
or U10368 (N_10368,N_7628,N_8778);
xor U10369 (N_10369,N_5548,N_6237);
or U10370 (N_10370,N_7582,N_8530);
and U10371 (N_10371,N_7392,N_7559);
nor U10372 (N_10372,N_7622,N_7551);
or U10373 (N_10373,N_5579,N_8558);
and U10374 (N_10374,N_6341,N_5030);
nand U10375 (N_10375,N_8326,N_7118);
nor U10376 (N_10376,N_6750,N_6752);
nand U10377 (N_10377,N_7001,N_8286);
nand U10378 (N_10378,N_9947,N_6766);
nand U10379 (N_10379,N_5162,N_7343);
nand U10380 (N_10380,N_9652,N_5073);
nand U10381 (N_10381,N_9892,N_8880);
or U10382 (N_10382,N_5974,N_9767);
nand U10383 (N_10383,N_6650,N_7215);
and U10384 (N_10384,N_9972,N_6158);
xnor U10385 (N_10385,N_9338,N_9445);
nand U10386 (N_10386,N_6559,N_8080);
xnor U10387 (N_10387,N_7734,N_8973);
xor U10388 (N_10388,N_5117,N_5779);
nor U10389 (N_10389,N_6611,N_7914);
and U10390 (N_10390,N_6585,N_7189);
and U10391 (N_10391,N_5996,N_8048);
and U10392 (N_10392,N_8992,N_6011);
nand U10393 (N_10393,N_6114,N_9497);
xnor U10394 (N_10394,N_7937,N_8457);
xnor U10395 (N_10395,N_6305,N_9059);
and U10396 (N_10396,N_9142,N_7328);
xnor U10397 (N_10397,N_5562,N_5930);
nand U10398 (N_10398,N_7996,N_8912);
xnor U10399 (N_10399,N_7740,N_8632);
xor U10400 (N_10400,N_6196,N_6480);
nand U10401 (N_10401,N_8869,N_7206);
or U10402 (N_10402,N_6042,N_7952);
nor U10403 (N_10403,N_5294,N_9291);
nand U10404 (N_10404,N_9629,N_8431);
or U10405 (N_10405,N_5473,N_5846);
or U10406 (N_10406,N_7772,N_8503);
nand U10407 (N_10407,N_9707,N_6225);
xor U10408 (N_10408,N_8677,N_7158);
nand U10409 (N_10409,N_9302,N_6550);
and U10410 (N_10410,N_9103,N_5673);
xor U10411 (N_10411,N_8474,N_9768);
nand U10412 (N_10412,N_6482,N_8804);
nand U10413 (N_10413,N_8268,N_8502);
nor U10414 (N_10414,N_7242,N_9324);
xor U10415 (N_10415,N_8874,N_9245);
nand U10416 (N_10416,N_9540,N_6861);
xnor U10417 (N_10417,N_9070,N_8083);
and U10418 (N_10418,N_8769,N_6051);
nor U10419 (N_10419,N_8181,N_8454);
xnor U10420 (N_10420,N_6371,N_8562);
or U10421 (N_10421,N_5550,N_7645);
and U10422 (N_10422,N_8383,N_8089);
and U10423 (N_10423,N_6177,N_6743);
or U10424 (N_10424,N_8314,N_9005);
and U10425 (N_10425,N_7961,N_9203);
xor U10426 (N_10426,N_7367,N_7757);
xnor U10427 (N_10427,N_9093,N_7256);
nor U10428 (N_10428,N_7503,N_7950);
nand U10429 (N_10429,N_5763,N_9286);
xor U10430 (N_10430,N_5995,N_9241);
nor U10431 (N_10431,N_5242,N_9588);
or U10432 (N_10432,N_7570,N_6381);
nor U10433 (N_10433,N_5416,N_5081);
nor U10434 (N_10434,N_6015,N_7687);
xor U10435 (N_10435,N_8971,N_6275);
or U10436 (N_10436,N_6596,N_5689);
or U10437 (N_10437,N_6726,N_7512);
and U10438 (N_10438,N_9164,N_5883);
nor U10439 (N_10439,N_8682,N_6847);
nor U10440 (N_10440,N_8026,N_9887);
nand U10441 (N_10441,N_5334,N_6470);
xor U10442 (N_10442,N_7245,N_9581);
nor U10443 (N_10443,N_7544,N_5520);
or U10444 (N_10444,N_8098,N_7095);
or U10445 (N_10445,N_9663,N_7677);
nor U10446 (N_10446,N_8447,N_9072);
nand U10447 (N_10447,N_6553,N_9534);
nand U10448 (N_10448,N_6665,N_6723);
xnor U10449 (N_10449,N_7838,N_8435);
nand U10450 (N_10450,N_5209,N_9423);
nand U10451 (N_10451,N_5188,N_5115);
nor U10452 (N_10452,N_7982,N_5778);
xor U10453 (N_10453,N_6297,N_9028);
xor U10454 (N_10454,N_5802,N_8106);
and U10455 (N_10455,N_8777,N_7616);
or U10456 (N_10456,N_5101,N_8610);
and U10457 (N_10457,N_7470,N_9531);
or U10458 (N_10458,N_5332,N_8408);
nand U10459 (N_10459,N_5148,N_7683);
and U10460 (N_10460,N_7404,N_7686);
xor U10461 (N_10461,N_5746,N_7719);
nand U10462 (N_10462,N_5311,N_5341);
and U10463 (N_10463,N_7260,N_9464);
xnor U10464 (N_10464,N_8719,N_8602);
nand U10465 (N_10465,N_7802,N_8409);
xnor U10466 (N_10466,N_5654,N_7055);
or U10467 (N_10467,N_8848,N_7234);
or U10468 (N_10468,N_8224,N_5109);
xnor U10469 (N_10469,N_5353,N_7580);
nor U10470 (N_10470,N_6844,N_7891);
nor U10471 (N_10471,N_6449,N_5827);
and U10472 (N_10472,N_7157,N_5172);
nor U10473 (N_10473,N_6019,N_9745);
xnor U10474 (N_10474,N_8327,N_5769);
and U10475 (N_10475,N_6580,N_9922);
xor U10476 (N_10476,N_5658,N_7892);
or U10477 (N_10477,N_8147,N_7408);
nor U10478 (N_10478,N_9218,N_7330);
nor U10479 (N_10479,N_8442,N_9829);
and U10480 (N_10480,N_7193,N_8053);
and U10481 (N_10481,N_6813,N_5421);
nand U10482 (N_10482,N_9404,N_6222);
nor U10483 (N_10483,N_8750,N_5533);
xor U10484 (N_10484,N_5216,N_7968);
and U10485 (N_10485,N_5126,N_8767);
nor U10486 (N_10486,N_9958,N_7612);
and U10487 (N_10487,N_6280,N_9309);
and U10488 (N_10488,N_9536,N_9794);
nand U10489 (N_10489,N_8228,N_7136);
xor U10490 (N_10490,N_7670,N_7395);
or U10491 (N_10491,N_8041,N_8998);
and U10492 (N_10492,N_9340,N_8329);
and U10493 (N_10493,N_9206,N_6725);
nand U10494 (N_10494,N_7518,N_9471);
or U10495 (N_10495,N_8239,N_6037);
or U10496 (N_10496,N_8872,N_7249);
or U10497 (N_10497,N_6227,N_8016);
nand U10498 (N_10498,N_7047,N_9799);
xor U10499 (N_10499,N_7797,N_9700);
xor U10500 (N_10500,N_5466,N_7170);
nand U10501 (N_10501,N_9417,N_6063);
nor U10502 (N_10502,N_9358,N_7201);
xnor U10503 (N_10503,N_8820,N_5701);
xnor U10504 (N_10504,N_5932,N_7284);
xor U10505 (N_10505,N_7881,N_7248);
and U10506 (N_10506,N_7306,N_5462);
nor U10507 (N_10507,N_7494,N_5541);
nand U10508 (N_10508,N_9224,N_7085);
xnor U10509 (N_10509,N_6346,N_9453);
xor U10510 (N_10510,N_5495,N_8943);
xnor U10511 (N_10511,N_6365,N_8006);
nand U10512 (N_10512,N_6013,N_9253);
or U10513 (N_10513,N_8433,N_8120);
nor U10514 (N_10514,N_9297,N_8557);
nand U10515 (N_10515,N_6411,N_7411);
or U10516 (N_10516,N_5441,N_9210);
nor U10517 (N_10517,N_6886,N_6116);
nor U10518 (N_10518,N_8407,N_9806);
and U10519 (N_10519,N_5678,N_6686);
xnor U10520 (N_10520,N_6510,N_5459);
or U10521 (N_10521,N_9180,N_9399);
nor U10522 (N_10522,N_6746,N_9879);
or U10523 (N_10523,N_9692,N_8655);
and U10524 (N_10524,N_6932,N_9126);
nor U10525 (N_10525,N_7907,N_5563);
and U10526 (N_10526,N_6172,N_6270);
or U10527 (N_10527,N_6337,N_7420);
and U10528 (N_10528,N_7409,N_7893);
or U10529 (N_10529,N_9390,N_9136);
nor U10530 (N_10530,N_8465,N_9177);
xnor U10531 (N_10531,N_7735,N_9484);
or U10532 (N_10532,N_9823,N_8940);
nor U10533 (N_10533,N_7145,N_5947);
or U10534 (N_10534,N_5937,N_7149);
nor U10535 (N_10535,N_8229,N_6552);
or U10536 (N_10536,N_7073,N_5601);
or U10537 (N_10537,N_7948,N_6323);
xor U10538 (N_10538,N_9315,N_9290);
nand U10539 (N_10539,N_7675,N_7147);
or U10540 (N_10540,N_5820,N_5240);
nor U10541 (N_10541,N_5159,N_5860);
xor U10542 (N_10542,N_6393,N_6103);
xnor U10543 (N_10543,N_7517,N_8808);
nor U10544 (N_10544,N_9657,N_6113);
nand U10545 (N_10545,N_8652,N_9850);
nor U10546 (N_10546,N_5896,N_7548);
or U10547 (N_10547,N_7969,N_7120);
and U10548 (N_10548,N_7198,N_5503);
nand U10549 (N_10549,N_5961,N_9744);
xnor U10550 (N_10550,N_7283,N_8631);
nor U10551 (N_10551,N_5200,N_6085);
or U10552 (N_10552,N_6408,N_8237);
or U10553 (N_10553,N_9623,N_9167);
or U10554 (N_10554,N_5110,N_7872);
nand U10555 (N_10555,N_9609,N_8391);
nor U10556 (N_10556,N_8550,N_7633);
nor U10557 (N_10557,N_9876,N_6531);
and U10558 (N_10558,N_5378,N_5080);
nor U10559 (N_10559,N_8110,N_9054);
and U10560 (N_10560,N_5828,N_6021);
xor U10561 (N_10561,N_9500,N_7671);
or U10562 (N_10562,N_5559,N_5668);
or U10563 (N_10563,N_7963,N_9884);
or U10564 (N_10564,N_8192,N_8064);
and U10565 (N_10565,N_8377,N_6140);
nor U10566 (N_10566,N_9704,N_5354);
and U10567 (N_10567,N_7851,N_7356);
and U10568 (N_10568,N_5984,N_6201);
xor U10569 (N_10569,N_5406,N_6706);
nor U10570 (N_10570,N_6223,N_7610);
nor U10571 (N_10571,N_6282,N_9797);
nand U10572 (N_10572,N_7641,N_6092);
xnor U10573 (N_10573,N_5552,N_8625);
nor U10574 (N_10574,N_7634,N_5263);
nor U10575 (N_10575,N_7462,N_5640);
nand U10576 (N_10576,N_7458,N_5967);
nor U10577 (N_10577,N_5933,N_9866);
or U10578 (N_10578,N_6684,N_7502);
and U10579 (N_10579,N_8323,N_6613);
nand U10580 (N_10580,N_5630,N_6934);
xor U10581 (N_10581,N_5191,N_9026);
nand U10582 (N_10582,N_6111,N_5207);
or U10583 (N_10583,N_8592,N_6948);
nand U10584 (N_10584,N_9013,N_5572);
nor U10585 (N_10585,N_5171,N_5913);
nor U10586 (N_10586,N_9910,N_6306);
nand U10587 (N_10587,N_6833,N_5878);
or U10588 (N_10588,N_5119,N_9695);
and U10589 (N_10589,N_7267,N_5456);
or U10590 (N_10590,N_6008,N_9475);
xnor U10591 (N_10591,N_9810,N_5838);
xnor U10592 (N_10592,N_6403,N_8151);
nor U10593 (N_10593,N_6696,N_8663);
or U10594 (N_10594,N_6168,N_8251);
or U10595 (N_10595,N_8201,N_8680);
and U10596 (N_10596,N_7398,N_5770);
nor U10597 (N_10597,N_8963,N_6230);
and U10598 (N_10598,N_6974,N_9559);
xor U10599 (N_10599,N_5422,N_8318);
xnor U10600 (N_10600,N_8217,N_7031);
and U10601 (N_10601,N_8841,N_8369);
nand U10602 (N_10602,N_5594,N_6047);
nand U10603 (N_10603,N_6908,N_8829);
and U10604 (N_10604,N_8601,N_8824);
or U10605 (N_10605,N_7063,N_7861);
xor U10606 (N_10606,N_8866,N_6468);
or U10607 (N_10607,N_8009,N_7839);
and U10608 (N_10608,N_9625,N_6988);
nor U10609 (N_10609,N_7667,N_5318);
nand U10610 (N_10610,N_5561,N_6738);
nor U10611 (N_10611,N_7171,N_5271);
nor U10612 (N_10612,N_5379,N_8588);
xor U10613 (N_10613,N_5835,N_8611);
or U10614 (N_10614,N_6919,N_8250);
nand U10615 (N_10615,N_8608,N_9983);
and U10616 (N_10616,N_8923,N_8654);
nand U10617 (N_10617,N_7305,N_5493);
and U10618 (N_10618,N_6731,N_6146);
or U10619 (N_10619,N_8938,N_6289);
or U10620 (N_10620,N_7358,N_8269);
and U10621 (N_10621,N_6410,N_5248);
or U10622 (N_10622,N_7995,N_7011);
nand U10623 (N_10623,N_9122,N_9686);
nand U10624 (N_10624,N_6477,N_5177);
or U10625 (N_10625,N_5393,N_8746);
or U10626 (N_10626,N_7599,N_5164);
or U10627 (N_10627,N_6602,N_5895);
nand U10628 (N_10628,N_5987,N_7885);
xor U10629 (N_10629,N_9508,N_8165);
or U10630 (N_10630,N_7540,N_7729);
nor U10631 (N_10631,N_9421,N_9499);
nor U10632 (N_10632,N_9127,N_5553);
nor U10633 (N_10633,N_6029,N_9631);
nand U10634 (N_10634,N_8958,N_6804);
nor U10635 (N_10635,N_6229,N_5513);
and U10636 (N_10636,N_5877,N_9888);
or U10637 (N_10637,N_7266,N_8374);
nor U10638 (N_10638,N_5269,N_5856);
nor U10639 (N_10639,N_8968,N_9792);
xor U10640 (N_10640,N_5751,N_7116);
xnor U10641 (N_10641,N_9746,N_9125);
xor U10642 (N_10642,N_7830,N_8209);
nor U10643 (N_10643,N_9951,N_7299);
or U10644 (N_10644,N_7181,N_9260);
and U10645 (N_10645,N_6053,N_7873);
or U10646 (N_10646,N_9969,N_6694);
xor U10647 (N_10647,N_9277,N_9612);
and U10648 (N_10648,N_7545,N_6882);
or U10649 (N_10649,N_7592,N_7056);
nand U10650 (N_10650,N_5068,N_9238);
or U10651 (N_10651,N_8007,N_5321);
nand U10652 (N_10652,N_7140,N_5525);
and U10653 (N_10653,N_5686,N_6888);
nand U10654 (N_10654,N_6890,N_7564);
nand U10655 (N_10655,N_9494,N_5058);
nor U10656 (N_10656,N_8427,N_6840);
nand U10657 (N_10657,N_6710,N_6671);
or U10658 (N_10658,N_5954,N_6770);
nand U10659 (N_10659,N_9162,N_9265);
or U10660 (N_10660,N_7090,N_6190);
xnor U10661 (N_10661,N_7749,N_7471);
and U10662 (N_10662,N_9672,N_8079);
xor U10663 (N_10663,N_8895,N_6334);
and U10664 (N_10664,N_8338,N_6670);
xor U10665 (N_10665,N_6634,N_6155);
nor U10666 (N_10666,N_5535,N_6912);
nor U10667 (N_10667,N_7617,N_7058);
and U10668 (N_10668,N_6587,N_9491);
or U10669 (N_10669,N_9520,N_5096);
and U10670 (N_10670,N_5343,N_8908);
nand U10671 (N_10671,N_5611,N_9485);
nand U10672 (N_10672,N_8892,N_8639);
or U10673 (N_10673,N_6683,N_8278);
xnor U10674 (N_10674,N_9955,N_7219);
xor U10675 (N_10675,N_5514,N_9010);
nand U10676 (N_10676,N_8806,N_6387);
nand U10677 (N_10677,N_9360,N_7745);
xor U10678 (N_10678,N_8619,N_7176);
xnor U10679 (N_10679,N_6472,N_8069);
nand U10680 (N_10680,N_6369,N_8031);
xnor U10681 (N_10681,N_7229,N_8786);
and U10682 (N_10682,N_5227,N_8259);
xor U10683 (N_10683,N_9688,N_8164);
and U10684 (N_10684,N_7609,N_7054);
nand U10685 (N_10685,N_8235,N_7327);
nor U10686 (N_10686,N_6333,N_5578);
and U10687 (N_10687,N_5972,N_6896);
or U10688 (N_10688,N_8439,N_7552);
xor U10689 (N_10689,N_9849,N_9923);
nand U10690 (N_10690,N_9134,N_6523);
nor U10691 (N_10691,N_7602,N_9194);
nor U10692 (N_10692,N_8411,N_6283);
or U10693 (N_10693,N_7753,N_7664);
xnor U10694 (N_10694,N_9967,N_7293);
or U10695 (N_10695,N_7106,N_5181);
nor U10696 (N_10696,N_5002,N_7926);
or U10697 (N_10697,N_5693,N_5483);
or U10698 (N_10698,N_6543,N_5885);
nor U10699 (N_10699,N_5254,N_9080);
xor U10700 (N_10700,N_5608,N_6385);
or U10701 (N_10701,N_5505,N_6067);
and U10702 (N_10702,N_6911,N_5065);
xnor U10703 (N_10703,N_5674,N_9680);
nor U10704 (N_10704,N_5265,N_9347);
nand U10705 (N_10705,N_7321,N_9346);
nor U10706 (N_10706,N_7130,N_6856);
xnor U10707 (N_10707,N_9029,N_8307);
xor U10708 (N_10708,N_8899,N_9430);
nor U10709 (N_10709,N_8003,N_8364);
and U10710 (N_10710,N_8115,N_8554);
nor U10711 (N_10711,N_7046,N_5194);
nand U10712 (N_10712,N_7221,N_7183);
xor U10713 (N_10713,N_9556,N_5623);
and U10714 (N_10714,N_7240,N_8486);
and U10715 (N_10715,N_8574,N_7199);
xor U10716 (N_10716,N_9833,N_5201);
or U10717 (N_10717,N_5006,N_8591);
nand U10718 (N_10718,N_9280,N_9483);
and U10719 (N_10719,N_6643,N_6703);
and U10720 (N_10720,N_5000,N_5272);
nand U10721 (N_10721,N_7191,N_5482);
and U10722 (N_10722,N_8094,N_9762);
or U10723 (N_10723,N_5011,N_7708);
xor U10724 (N_10724,N_9139,N_5875);
or U10725 (N_10725,N_5142,N_6441);
nand U10726 (N_10726,N_7226,N_8225);
nand U10727 (N_10727,N_5522,N_5593);
or U10728 (N_10728,N_5490,N_5833);
xor U10729 (N_10729,N_5173,N_7084);
xor U10730 (N_10730,N_6133,N_8355);
xor U10731 (N_10731,N_9869,N_5706);
nand U10732 (N_10732,N_7579,N_6522);
nand U10733 (N_10733,N_8666,N_8342);
or U10734 (N_10734,N_7701,N_7703);
nor U10735 (N_10735,N_8313,N_8950);
nand U10736 (N_10736,N_6761,N_5291);
and U10737 (N_10737,N_6630,N_6290);
or U10738 (N_10738,N_5056,N_9509);
or U10739 (N_10739,N_7110,N_6136);
xnor U10740 (N_10740,N_5868,N_6933);
or U10741 (N_10741,N_7676,N_9237);
nand U10742 (N_10742,N_7988,N_8346);
and U10743 (N_10743,N_7375,N_6414);
nor U10744 (N_10744,N_9719,N_6893);
nor U10745 (N_10745,N_9564,N_7435);
nor U10746 (N_10746,N_9294,N_7211);
and U10747 (N_10747,N_8529,N_9284);
xor U10748 (N_10748,N_7426,N_7832);
xnor U10749 (N_10749,N_7374,N_6207);
or U10750 (N_10750,N_6689,N_6267);
or U10751 (N_10751,N_5494,N_9215);
or U10752 (N_10752,N_8979,N_8341);
and U10753 (N_10753,N_6698,N_5547);
and U10754 (N_10754,N_5362,N_7889);
nand U10755 (N_10755,N_5492,N_5044);
and U10756 (N_10756,N_5186,N_7077);
nand U10757 (N_10757,N_5415,N_5970);
xor U10758 (N_10758,N_5960,N_8417);
nor U10759 (N_10759,N_7059,N_8117);
or U10760 (N_10760,N_8174,N_8159);
and U10761 (N_10761,N_8653,N_7291);
nor U10762 (N_10762,N_5222,N_7964);
nand U10763 (N_10763,N_9477,N_8216);
xnor U10764 (N_10764,N_7546,N_9600);
or U10765 (N_10765,N_9381,N_8024);
xor U10766 (N_10766,N_5694,N_9905);
and U10767 (N_10767,N_9802,N_8735);
and U10768 (N_10768,N_6161,N_8190);
xor U10769 (N_10769,N_7651,N_7065);
or U10770 (N_10770,N_7269,N_5498);
or U10771 (N_10771,N_5690,N_5040);
or U10772 (N_10772,N_8072,N_9157);
or U10773 (N_10773,N_6984,N_5290);
xor U10774 (N_10774,N_9890,N_5339);
or U10775 (N_10775,N_9698,N_8805);
xor U10776 (N_10776,N_6803,N_6081);
nand U10777 (N_10777,N_6955,N_9014);
and U10778 (N_10778,N_7812,N_8279);
nor U10779 (N_10779,N_8888,N_5267);
nor U10780 (N_10780,N_9932,N_7843);
nor U10781 (N_10781,N_5055,N_8842);
and U10782 (N_10782,N_5089,N_8772);
or U10783 (N_10783,N_8921,N_6773);
nor U10784 (N_10784,N_5316,N_9148);
xnor U10785 (N_10785,N_8111,N_7339);
nand U10786 (N_10786,N_5554,N_8322);
nand U10787 (N_10787,N_9844,N_6185);
or U10788 (N_10788,N_9048,N_8936);
and U10789 (N_10789,N_5942,N_6491);
xor U10790 (N_10790,N_9366,N_6335);
and U10791 (N_10791,N_7382,N_5220);
or U10792 (N_10792,N_9306,N_5097);
xnor U10793 (N_10793,N_7928,N_7288);
nor U10794 (N_10794,N_9269,N_5346);
nor U10795 (N_10795,N_6606,N_6395);
xnor U10796 (N_10796,N_5028,N_8944);
xor U10797 (N_10797,N_6917,N_7071);
xor U10798 (N_10798,N_6145,N_7902);
xor U10799 (N_10799,N_8445,N_7844);
and U10800 (N_10800,N_8422,N_8443);
xor U10801 (N_10801,N_7853,N_6629);
xnor U10802 (N_10802,N_8449,N_7134);
or U10803 (N_10803,N_8227,N_6300);
nand U10804 (N_10804,N_7272,N_9541);
nor U10805 (N_10805,N_5247,N_8603);
or U10806 (N_10806,N_8597,N_7932);
nand U10807 (N_10807,N_9687,N_8137);
nand U10808 (N_10808,N_5424,N_5037);
nand U10809 (N_10809,N_8742,N_9063);
or U10810 (N_10810,N_7521,N_6938);
xor U10811 (N_10811,N_9840,N_7584);
or U10812 (N_10812,N_8208,N_6728);
nand U10813 (N_10813,N_9479,N_7465);
nor U10814 (N_10814,N_7310,N_6625);
nand U10815 (N_10815,N_7520,N_8244);
xnor U10816 (N_10816,N_5093,N_5063);
nor U10817 (N_10817,N_5434,N_7528);
and U10818 (N_10818,N_6272,N_5862);
xnor U10819 (N_10819,N_7216,N_9248);
or U10820 (N_10820,N_5953,N_5582);
xor U10821 (N_10821,N_8604,N_8330);
nor U10822 (N_10822,N_9660,N_7886);
nand U10823 (N_10823,N_8175,N_5831);
nand U10824 (N_10824,N_8661,N_6928);
nor U10825 (N_10825,N_9756,N_6046);
or U10826 (N_10826,N_8044,N_9701);
xor U10827 (N_10827,N_6873,N_8063);
nor U10828 (N_10828,N_8162,N_9137);
or U10829 (N_10829,N_8650,N_8487);
xnor U10830 (N_10830,N_7067,N_5477);
nor U10831 (N_10831,N_5052,N_6924);
or U10832 (N_10832,N_8141,N_9780);
and U10833 (N_10833,N_6043,N_9153);
nand U10834 (N_10834,N_7192,N_8393);
and U10835 (N_10835,N_6160,N_6490);
nor U10836 (N_10836,N_5180,N_8519);
nand U10837 (N_10837,N_6097,N_6162);
nor U10838 (N_10838,N_5643,N_9920);
nand U10839 (N_10839,N_8036,N_6132);
and U10840 (N_10840,N_7365,N_9244);
nor U10841 (N_10841,N_6889,N_5516);
xnor U10842 (N_10842,N_7080,N_9630);
xor U10843 (N_10843,N_6848,N_8400);
nor U10844 (N_10844,N_7372,N_9651);
xor U10845 (N_10845,N_8523,N_8555);
nand U10846 (N_10846,N_9197,N_6149);
or U10847 (N_10847,N_7653,N_5604);
xor U10848 (N_10848,N_8696,N_9480);
or U10849 (N_10849,N_5975,N_8645);
nor U10850 (N_10850,N_5067,N_8844);
and U10851 (N_10851,N_9305,N_7682);
xor U10852 (N_10852,N_9262,N_7353);
and U10853 (N_10853,N_5061,N_9371);
nand U10854 (N_10854,N_8105,N_6729);
or U10855 (N_10855,N_7679,N_7135);
nor U10856 (N_10856,N_5426,N_5084);
xor U10857 (N_10857,N_8113,N_6685);
xor U10858 (N_10858,N_5021,N_6469);
or U10859 (N_10859,N_6878,N_5634);
xnor U10860 (N_10860,N_6435,N_6169);
or U10861 (N_10861,N_9518,N_6517);
or U10862 (N_10862,N_8040,N_8077);
nor U10863 (N_10863,N_6238,N_8630);
nand U10864 (N_10864,N_9223,N_8852);
or U10865 (N_10865,N_9092,N_7850);
or U10866 (N_10866,N_6936,N_7146);
xnor U10867 (N_10867,N_5370,N_8600);
or U10868 (N_10868,N_5785,N_9598);
and U10869 (N_10869,N_6567,N_5676);
and U10870 (N_10870,N_9897,N_8112);
xor U10871 (N_10871,N_5922,N_8576);
and U10872 (N_10872,N_9925,N_6921);
nand U10873 (N_10873,N_9336,N_8509);
nand U10874 (N_10874,N_6000,N_8656);
and U10875 (N_10875,N_8289,N_7852);
and U10876 (N_10876,N_8760,N_8308);
and U10877 (N_10877,N_8419,N_8926);
xnor U10878 (N_10878,N_6330,N_8705);
and U10879 (N_10879,N_9647,N_7710);
nand U10880 (N_10880,N_9008,N_6205);
xnor U10881 (N_10881,N_9355,N_8843);
xor U10882 (N_10882,N_5940,N_7125);
xnor U10883 (N_10883,N_7884,N_5212);
xor U10884 (N_10884,N_5112,N_9778);
nor U10885 (N_10885,N_7674,N_7258);
xor U10886 (N_10886,N_6370,N_6202);
and U10887 (N_10887,N_6210,N_6279);
and U10888 (N_10888,N_7029,N_7646);
nand U10889 (N_10889,N_6143,N_8275);
xor U10890 (N_10890,N_6581,N_9804);
xor U10891 (N_10891,N_6418,N_7618);
nand U10892 (N_10892,N_5374,N_6430);
or U10893 (N_10893,N_8352,N_5744);
or U10894 (N_10894,N_5054,N_9971);
and U10895 (N_10895,N_8299,N_5849);
nor U10896 (N_10896,N_7497,N_6568);
nor U10897 (N_10897,N_7532,N_6443);
and U10898 (N_10898,N_6871,N_5772);
xor U10899 (N_10899,N_6739,N_5440);
xnor U10900 (N_10900,N_6967,N_9105);
nor U10901 (N_10901,N_6232,N_6350);
and U10902 (N_10902,N_5264,N_6428);
and U10903 (N_10903,N_8563,N_9664);
and U10904 (N_10904,N_9521,N_9062);
and U10905 (N_10905,N_5257,N_8624);
nor U10906 (N_10906,N_5981,N_6302);
nor U10907 (N_10907,N_9595,N_8482);
and U10908 (N_10908,N_6117,N_9594);
or U10909 (N_10909,N_6918,N_5738);
nor U10910 (N_10910,N_5808,N_9911);
and U10911 (N_10911,N_9383,N_7601);
and U10912 (N_10912,N_9274,N_8986);
nor U10913 (N_10913,N_7595,N_7983);
xnor U10914 (N_10914,N_6964,N_7555);
and U10915 (N_10915,N_9577,N_8453);
or U10916 (N_10916,N_8584,N_9893);
xor U10917 (N_10917,N_8166,N_6925);
xor U10918 (N_10918,N_7900,N_7270);
xnor U10919 (N_10919,N_7771,N_7455);
xnor U10920 (N_10920,N_9201,N_6353);
nor U10921 (N_10921,N_7931,N_8205);
xor U10922 (N_10922,N_6233,N_7418);
xnor U10923 (N_10923,N_5453,N_8703);
or U10924 (N_10924,N_8021,N_9545);
nand U10925 (N_10925,N_9208,N_6478);
xor U10926 (N_10926,N_5991,N_8128);
xnor U10927 (N_10927,N_8233,N_8741);
or U10928 (N_10928,N_6445,N_9591);
and U10929 (N_10929,N_7172,N_8153);
xnor U10930 (N_10930,N_5210,N_6875);
nor U10931 (N_10931,N_5735,N_7352);
and U10932 (N_10932,N_8622,N_9868);
xnor U10933 (N_10933,N_6525,N_5952);
or U10934 (N_10934,N_5184,N_9333);
nor U10935 (N_10935,N_8609,N_7164);
or U10936 (N_10936,N_8220,N_8464);
nand U10937 (N_10937,N_7371,N_5605);
or U10938 (N_10938,N_8830,N_8595);
or U10939 (N_10939,N_8616,N_8102);
or U10940 (N_10940,N_5484,N_5420);
xor U10941 (N_10941,N_9064,N_9463);
or U10942 (N_10942,N_9936,N_9587);
or U10943 (N_10943,N_5504,N_6712);
and U10944 (N_10944,N_5925,N_8560);
xnor U10945 (N_10945,N_6488,N_5528);
and U10946 (N_10946,N_9535,N_5367);
nand U10947 (N_10947,N_7394,N_6744);
nor U10948 (N_10948,N_8817,N_5077);
and U10949 (N_10949,N_5679,N_9710);
nand U10950 (N_10950,N_9275,N_5278);
and U10951 (N_10951,N_5309,N_9506);
xor U10952 (N_10952,N_5549,N_6829);
nor U10953 (N_10953,N_7022,N_5998);
and U10954 (N_10954,N_6138,N_5085);
or U10955 (N_10955,N_6325,N_8737);
and U10956 (N_10956,N_5580,N_8967);
or U10957 (N_10957,N_6677,N_5700);
nand U10958 (N_10958,N_9356,N_8353);
nor U10959 (N_10959,N_6560,N_9115);
nor U10960 (N_10960,N_8785,N_5310);
and U10961 (N_10961,N_6105,N_8183);
and U10962 (N_10962,N_7005,N_7716);
nor U10963 (N_10963,N_8910,N_6947);
or U10964 (N_10964,N_8882,N_7698);
nand U10965 (N_10965,N_5412,N_7752);
and U10966 (N_10966,N_9730,N_7818);
nand U10967 (N_10967,N_9977,N_9826);
xor U10968 (N_10968,N_5672,N_6498);
or U10969 (N_10969,N_6790,N_7101);
or U10970 (N_10970,N_6635,N_8160);
nand U10971 (N_10971,N_8285,N_9342);
nor U10972 (N_10972,N_5585,N_8350);
or U10973 (N_10973,N_6681,N_9899);
or U10974 (N_10974,N_8213,N_8440);
xnor U10975 (N_10975,N_9007,N_9429);
or U10976 (N_10976,N_6653,N_9763);
nor U10977 (N_10977,N_7668,N_8761);
or U10978 (N_10978,N_5733,N_6396);
xnor U10979 (N_10979,N_6755,N_8462);
nor U10980 (N_10980,N_6311,N_5404);
xor U10981 (N_10981,N_6961,N_6906);
or U10982 (N_10982,N_5135,N_9326);
nor U10983 (N_10983,N_9332,N_7737);
nor U10984 (N_10984,N_7805,N_9051);
nor U10985 (N_10985,N_5394,N_6608);
nand U10986 (N_10986,N_7485,N_9432);
nand U10987 (N_10987,N_8473,N_7799);
nand U10988 (N_10988,N_6598,N_7415);
nor U10989 (N_10989,N_9551,N_5789);
xor U10990 (N_10990,N_9295,N_5602);
nand U10991 (N_10991,N_7702,N_7333);
nand U10992 (N_10992,N_5121,N_9102);
and U10993 (N_10993,N_8477,N_8002);
nand U10994 (N_10994,N_8130,N_8875);
nand U10995 (N_10995,N_9300,N_8188);
xor U10996 (N_10996,N_8402,N_8564);
nand U10997 (N_10997,N_6715,N_5558);
nand U10998 (N_10998,N_6827,N_8583);
nand U10999 (N_10999,N_9504,N_7264);
or U11000 (N_11000,N_7335,N_8023);
nand U11001 (N_11001,N_5091,N_5764);
and U11002 (N_11002,N_6386,N_8272);
or U11003 (N_11003,N_9992,N_5711);
xnor U11004 (N_11004,N_6556,N_6319);
nor U11005 (N_11005,N_6206,N_6816);
nand U11006 (N_11006,N_6194,N_9681);
nor U11007 (N_11007,N_7203,N_8030);
nor U11008 (N_11008,N_6554,N_6292);
nand U11009 (N_11009,N_9656,N_9146);
nor U11010 (N_11010,N_6183,N_9783);
and U11011 (N_11011,N_9685,N_9601);
nor U11012 (N_11012,N_6865,N_5074);
nor U11013 (N_11013,N_6249,N_9528);
nand U11014 (N_11014,N_5632,N_7401);
nand U11015 (N_11015,N_5128,N_5120);
xnor U11016 (N_11016,N_8389,N_5882);
nor U11017 (N_11017,N_5475,N_9706);
xnor U11018 (N_11018,N_9141,N_5474);
and U11019 (N_11019,N_8264,N_5610);
or U11020 (N_11020,N_8512,N_8531);
nor U11021 (N_11021,N_5245,N_8303);
nor U11022 (N_11022,N_7537,N_7783);
and U11023 (N_11023,N_6494,N_9293);
and U11024 (N_11024,N_6399,N_9711);
xnor U11025 (N_11025,N_5390,N_8828);
xor U11026 (N_11026,N_9462,N_8701);
or U11027 (N_11027,N_7684,N_9953);
or U11028 (N_11028,N_5741,N_9908);
nor U11029 (N_11029,N_8376,N_6425);
nand U11030 (N_11030,N_5641,N_8738);
nand U11031 (N_11031,N_6361,N_8460);
and U11032 (N_11032,N_6783,N_8978);
and U11033 (N_11033,N_8536,N_5256);
nor U11034 (N_11034,N_8197,N_6981);
and U11035 (N_11035,N_8796,N_9524);
nor U11036 (N_11036,N_6310,N_8514);
and U11037 (N_11037,N_5955,N_5613);
nand U11038 (N_11038,N_9204,N_8886);
nor U11039 (N_11039,N_5197,N_7989);
or U11040 (N_11040,N_6995,N_9296);
xnor U11041 (N_11041,N_8418,N_6620);
xor U11042 (N_11042,N_6858,N_5607);
nand U11043 (N_11043,N_6812,N_7165);
or U11044 (N_11044,N_8095,N_7875);
and U11045 (N_11045,N_7457,N_9226);
nor U11046 (N_11046,N_5943,N_5469);
or U11047 (N_11047,N_5626,N_8455);
or U11048 (N_11048,N_9391,N_7261);
nor U11049 (N_11049,N_8469,N_8775);
and U11050 (N_11050,N_8878,N_9316);
and U11051 (N_11051,N_9440,N_5670);
nor U11052 (N_11052,N_9329,N_8929);
nand U11053 (N_11053,N_5071,N_6999);
nand U11054 (N_11054,N_7796,N_7483);
xnor U11055 (N_11055,N_7013,N_5804);
nor U11056 (N_11056,N_7476,N_7689);
or U11057 (N_11057,N_9832,N_7459);
xnor U11058 (N_11058,N_9715,N_9965);
nor U11059 (N_11059,N_7589,N_7008);
and U11060 (N_11060,N_6412,N_5904);
xnor U11061 (N_11061,N_5166,N_6788);
or U11062 (N_11062,N_6859,N_9790);
xnor U11063 (N_11063,N_6407,N_9596);
and U11064 (N_11064,N_9104,N_9405);
nor U11065 (N_11065,N_5451,N_5823);
or U11066 (N_11066,N_7531,N_9076);
or U11067 (N_11067,N_7127,N_7506);
nor U11068 (N_11068,N_8994,N_8012);
xor U11069 (N_11069,N_7611,N_7636);
nand U11070 (N_11070,N_8920,N_6944);
or U11071 (N_11071,N_5231,N_7081);
or U11072 (N_11072,N_9121,N_6079);
nand U11073 (N_11073,N_6195,N_9853);
xnor U11074 (N_11074,N_7089,N_5573);
xor U11075 (N_11075,N_7845,N_7168);
and U11076 (N_11076,N_5567,N_8189);
and U11077 (N_11077,N_9212,N_7451);
nor U11078 (N_11078,N_9658,N_8107);
nand U11079 (N_11079,N_7803,N_9079);
or U11080 (N_11080,N_9427,N_7391);
nor U11081 (N_11081,N_5319,N_8784);
xor U11082 (N_11082,N_7631,N_8990);
or U11083 (N_11083,N_9413,N_7437);
xnor U11084 (N_11084,N_5151,N_6340);
or U11085 (N_11085,N_5556,N_8492);
nor U11086 (N_11086,N_9257,N_9459);
nand U11087 (N_11087,N_9954,N_7368);
or U11088 (N_11088,N_7309,N_8516);
and U11089 (N_11089,N_5512,N_7680);
and U11090 (N_11090,N_7924,N_6722);
nand U11091 (N_11091,N_7840,N_6440);
nor U11092 (N_11092,N_7866,N_5108);
nor U11093 (N_11093,N_8170,N_7479);
and U11094 (N_11094,N_6362,N_7586);
xnor U11095 (N_11095,N_7649,N_8360);
and U11096 (N_11096,N_9349,N_7444);
nor U11097 (N_11097,N_7072,N_8941);
and U11098 (N_11098,N_5901,N_5897);
nor U11099 (N_11099,N_8739,N_9641);
or U11100 (N_11100,N_9722,N_7916);
nor U11101 (N_11101,N_5944,N_7488);
or U11102 (N_11102,N_6591,N_7515);
xnor U11103 (N_11103,N_8823,N_6239);
or U11104 (N_11104,N_8633,N_9562);
nor U11105 (N_11105,N_8108,N_8078);
or U11106 (N_11106,N_7051,N_7188);
or U11107 (N_11107,N_6661,N_6516);
or U11108 (N_11108,N_9787,N_8877);
nor U11109 (N_11109,N_7810,N_7093);
or U11110 (N_11110,N_8838,N_8748);
nand U11111 (N_11111,N_8758,N_5198);
xnor U11112 (N_11112,N_8288,N_6586);
nand U11113 (N_11113,N_8779,N_9798);
nor U11114 (N_11114,N_6943,N_8945);
nand U11115 (N_11115,N_5639,N_7919);
nor U11116 (N_11116,N_8861,N_5487);
or U11117 (N_11117,N_9450,N_5929);
and U11118 (N_11118,N_5178,N_7207);
or U11119 (N_11119,N_8527,N_8436);
and U11120 (N_11120,N_8262,N_5902);
or U11121 (N_11121,N_9683,N_7857);
nor U11122 (N_11122,N_7493,N_6235);
or U11123 (N_11123,N_8709,N_8916);
nor U11124 (N_11124,N_6259,N_9159);
or U11125 (N_11125,N_5935,N_6368);
nor U11126 (N_11126,N_5699,N_5375);
and U11127 (N_11127,N_5980,N_8498);
nor U11128 (N_11128,N_8249,N_6668);
nor U11129 (N_11129,N_8366,N_8679);
and U11130 (N_11130,N_6003,N_7519);
and U11131 (N_11131,N_5129,N_9570);
nand U11132 (N_11132,N_5377,N_6713);
xor U11133 (N_11133,N_7985,N_7185);
nor U11134 (N_11134,N_5223,N_9978);
nand U11135 (N_11135,N_8623,N_6315);
and U11136 (N_11136,N_5565,N_6301);
nand U11137 (N_11137,N_5748,N_8207);
and U11138 (N_11138,N_8306,N_8018);
or U11139 (N_11139,N_5429,N_5638);
or U11140 (N_11140,N_8977,N_8005);
or U11141 (N_11141,N_5727,N_8954);
or U11142 (N_11142,N_9788,N_5486);
nand U11143 (N_11143,N_5072,N_9960);
nand U11144 (N_11144,N_5501,N_5819);
xor U11145 (N_11145,N_5102,N_5986);
or U11146 (N_11146,N_5905,N_5215);
nand U11147 (N_11147,N_7733,N_6091);
xnor U11148 (N_11148,N_8763,N_5163);
nand U11149 (N_11149,N_9250,N_8586);
xor U11150 (N_11150,N_6157,N_9247);
xnor U11151 (N_11151,N_9431,N_8388);
nand U11152 (N_11152,N_7315,N_9066);
nand U11153 (N_11153,N_5795,N_6096);
xor U11154 (N_11154,N_6791,N_8669);
nor U11155 (N_11155,N_7870,N_8684);
xnor U11156 (N_11156,N_5445,N_9473);
xnor U11157 (N_11157,N_7775,N_5480);
or U11158 (N_11158,N_8524,N_7406);
xnor U11159 (N_11159,N_5661,N_9777);
or U11160 (N_11160,N_7854,N_5871);
nand U11161 (N_11161,N_7868,N_8298);
or U11162 (N_11162,N_8788,N_5457);
nand U11163 (N_11163,N_6990,N_9258);
nor U11164 (N_11164,N_6807,N_7385);
or U11165 (N_11165,N_5261,N_8731);
nand U11166 (N_11166,N_6558,N_5304);
and U11167 (N_11167,N_7213,N_9774);
nor U11168 (N_11168,N_7824,N_7958);
nand U11169 (N_11169,N_8354,N_5488);
or U11170 (N_11170,N_7386,N_6753);
xnor U11171 (N_11171,N_5306,N_8670);
nand U11172 (N_11172,N_6397,N_8468);
or U11173 (N_11173,N_8925,N_8428);
or U11174 (N_11174,N_7376,N_8590);
xnor U11175 (N_11175,N_5997,N_5308);
xnor U11176 (N_11176,N_5782,N_7874);
or U11177 (N_11177,N_6018,N_9350);
nor U11178 (N_11178,N_9254,N_7730);
xnor U11179 (N_11179,N_5657,N_6002);
xor U11180 (N_11180,N_9626,N_6460);
and U11181 (N_11181,N_9334,N_7549);
xnor U11182 (N_11182,N_9593,N_5978);
nand U11183 (N_11183,N_9156,N_8127);
nor U11184 (N_11184,N_9082,N_6377);
and U11185 (N_11185,N_6006,N_6855);
nor U11186 (N_11186,N_6593,N_6150);
or U11187 (N_11187,N_6156,N_8685);
or U11188 (N_11188,N_6505,N_8901);
or U11189 (N_11189,N_6390,N_7414);
or U11190 (N_11190,N_7659,N_6258);
or U11191 (N_11191,N_9605,N_7097);
xor U11192 (N_11192,N_6064,N_5976);
nand U11193 (N_11193,N_8753,N_9219);
and U11194 (N_11194,N_5239,N_6320);
nand U11195 (N_11195,N_6088,N_5865);
xor U11196 (N_11196,N_9952,N_5707);
and U11197 (N_11197,N_8815,N_6175);
or U11198 (N_11198,N_6324,N_9523);
or U11199 (N_11199,N_7300,N_6849);
or U11200 (N_11200,N_6842,N_5625);
or U11201 (N_11201,N_9370,N_6163);
or U11202 (N_11202,N_6373,N_8202);
nand U11203 (N_11203,N_6900,N_9160);
nor U11204 (N_11204,N_5478,N_8793);
nand U11205 (N_11205,N_6561,N_7111);
nor U11206 (N_11206,N_6234,N_8114);
or U11207 (N_11207,N_5545,N_8762);
xnor U11208 (N_11208,N_5737,N_5629);
nor U11209 (N_11209,N_8266,N_7039);
and U11210 (N_11210,N_9182,N_8585);
and U11211 (N_11211,N_7247,N_5844);
or U11212 (N_11212,N_5324,N_7082);
nand U11213 (N_11213,N_6772,N_5758);
xor U11214 (N_11214,N_6862,N_8283);
nand U11215 (N_11215,N_5380,N_6787);
nor U11216 (N_11216,N_7018,N_7091);
or U11217 (N_11217,N_9496,N_5176);
or U11218 (N_11218,N_9776,N_6060);
and U11219 (N_11219,N_6314,N_9987);
nand U11220 (N_11220,N_8380,N_8335);
nor U11221 (N_11221,N_7856,N_9174);
or U11222 (N_11222,N_9813,N_7042);
or U11223 (N_11223,N_7290,N_6032);
nor U11224 (N_11224,N_5347,N_5287);
nand U11225 (N_11225,N_5253,N_7074);
or U11226 (N_11226,N_9319,N_9345);
and U11227 (N_11227,N_9444,N_7762);
or U11228 (N_11228,N_6538,N_6623);
or U11229 (N_11229,N_9990,N_9881);
nand U11230 (N_11230,N_7276,N_6444);
nand U11231 (N_11231,N_6940,N_9052);
and U11232 (N_11232,N_8812,N_8126);
and U11233 (N_11233,N_6400,N_7393);
or U11234 (N_11234,N_9155,N_6214);
or U11235 (N_11235,N_6479,N_9495);
nand U11236 (N_11236,N_7052,N_9827);
xnor U11237 (N_11237,N_7619,N_8996);
or U11238 (N_11238,N_5850,N_6212);
or U11239 (N_11239,N_8548,N_7196);
and U11240 (N_11240,N_6462,N_8723);
xor U11241 (N_11241,N_5923,N_5408);
and U11242 (N_11242,N_9287,N_9836);
nand U11243 (N_11243,N_8870,N_6417);
and U11244 (N_11244,N_7750,N_9845);
nand U11245 (N_11245,N_9661,N_5752);
or U11246 (N_11246,N_7133,N_6030);
xor U11247 (N_11247,N_7380,N_6655);
xor U11248 (N_11248,N_7984,N_6112);
or U11249 (N_11249,N_8706,N_5444);
nand U11250 (N_11250,N_6692,N_8392);
and U11251 (N_11251,N_9949,N_7939);
and U11252 (N_11252,N_7361,N_6998);
and U11253 (N_11253,N_5959,N_7436);
xor U11254 (N_11254,N_6811,N_6126);
or U11255 (N_11255,N_8410,N_5742);
xnor U11256 (N_11256,N_9754,N_7510);
or U11257 (N_11257,N_7562,N_8062);
or U11258 (N_11258,N_5598,N_9200);
nor U11259 (N_11259,N_6675,N_8090);
nor U11260 (N_11260,N_6716,N_6997);
nor U11261 (N_11261,N_5767,N_9808);
nand U11262 (N_11262,N_9438,N_6489);
or U11263 (N_11263,N_7971,N_6854);
xnor U11264 (N_11264,N_9023,N_9667);
or U11265 (N_11265,N_8218,N_9086);
nand U11266 (N_11266,N_6336,N_6589);
nand U11267 (N_11267,N_5411,N_5596);
nand U11268 (N_11268,N_8171,N_9188);
and U11269 (N_11269,N_7433,N_9489);
xor U11270 (N_11270,N_7566,N_6877);
and U11271 (N_11271,N_6800,N_7038);
nand U11272 (N_11272,N_7275,N_8061);
or U11273 (N_11273,N_8093,N_6392);
or U11274 (N_11274,N_9170,N_5203);
nor U11275 (N_11275,N_8054,N_8180);
or U11276 (N_11276,N_5798,N_5468);
xnor U11277 (N_11277,N_5765,N_7403);
or U11278 (N_11278,N_5285,N_8800);
nor U11279 (N_11279,N_9589,N_7746);
xor U11280 (N_11280,N_6691,N_9049);
nand U11281 (N_11281,N_6632,N_5732);
and U11282 (N_11282,N_6957,N_7078);
nand U11283 (N_11283,N_6142,N_8506);
nor U11284 (N_11284,N_6515,N_9622);
nor U11285 (N_11285,N_6823,N_5888);
nor U11286 (N_11286,N_6601,N_7027);
and U11287 (N_11287,N_6682,N_6597);
nor U11288 (N_11288,N_5774,N_5760);
or U11289 (N_11289,N_8847,N_9073);
and U11290 (N_11290,N_7846,N_6167);
or U11291 (N_11291,N_5106,N_6007);
nand U11292 (N_11292,N_8359,N_7405);
xnor U11293 (N_11293,N_6141,N_9891);
nand U11294 (N_11294,N_7222,N_5275);
or U11295 (N_11295,N_5816,N_8168);
and U11296 (N_11296,N_7632,N_9882);
nand U11297 (N_11297,N_5221,N_7239);
or U11298 (N_11298,N_6243,N_9791);
and U11299 (N_11299,N_8385,N_5258);
or U11300 (N_11300,N_7794,N_7456);
xnor U11301 (N_11301,N_7232,N_7788);
nor U11302 (N_11302,N_9517,N_8458);
or U11303 (N_11303,N_5696,N_6547);
or U11304 (N_11304,N_8637,N_9703);
xor U11305 (N_11305,N_8017,N_7956);
and U11306 (N_11306,N_8511,N_7820);
xor U11307 (N_11307,N_5331,N_6266);
or U11308 (N_11308,N_9567,N_7014);
or U11309 (N_11309,N_7443,N_6805);
nor U11310 (N_11310,N_7720,N_6254);
and U11311 (N_11311,N_6551,N_5447);
and U11312 (N_11312,N_6349,N_5460);
xor U11313 (N_11313,N_9225,N_9361);
or U11314 (N_11314,N_5170,N_8232);
nand U11315 (N_11315,N_6562,N_8991);
and U11316 (N_11316,N_9709,N_6125);
xnor U11317 (N_11317,N_7317,N_9119);
xor U11318 (N_11318,N_5401,N_5603);
or U11319 (N_11319,N_6904,N_7967);
and U11320 (N_11320,N_9705,N_6618);
nand U11321 (N_11321,N_5273,N_6277);
xnor U11322 (N_11322,N_7060,N_9638);
and U11323 (N_11323,N_6958,N_6036);
xnor U11324 (N_11324,N_6954,N_9442);
nand U11325 (N_11325,N_8211,N_8713);
or U11326 (N_11326,N_9065,N_5957);
xnor U11327 (N_11327,N_8390,N_6014);
nand U11328 (N_11328,N_6792,N_8027);
and U11329 (N_11329,N_5587,N_6572);
or U11330 (N_11330,N_5917,N_7413);
nand U11331 (N_11331,N_7604,N_8015);
nor U11332 (N_11332,N_9555,N_7373);
nor U11333 (N_11333,N_5698,N_6278);
xor U11334 (N_11334,N_5500,N_6375);
and U11335 (N_11335,N_9898,N_7092);
and U11336 (N_11336,N_5773,N_7912);
nor U11337 (N_11337,N_7650,N_6180);
and U11338 (N_11338,N_6437,N_7463);
nor U11339 (N_11339,N_8572,N_7152);
xnor U11340 (N_11340,N_9716,N_6492);
or U11341 (N_11341,N_5249,N_5259);
xor U11342 (N_11342,N_8520,N_6901);
xor U11343 (N_11343,N_5105,N_5137);
and U11344 (N_11344,N_9181,N_9091);
and U11345 (N_11345,N_7577,N_5470);
or U11346 (N_11346,N_7318,N_5298);
and U11347 (N_11347,N_5864,N_5919);
and U11348 (N_11348,N_8138,N_5858);
xnor U11349 (N_11349,N_9282,N_5908);
or U11350 (N_11350,N_5840,N_7976);
xnor U11351 (N_11351,N_5179,N_7786);
nand U11352 (N_11352,N_8928,N_6868);
nor U11353 (N_11353,N_7307,N_7596);
or U11354 (N_11354,N_8001,N_5609);
and U11355 (N_11355,N_5205,N_5114);
or U11356 (N_11356,N_9717,N_9428);
and U11357 (N_11357,N_8708,N_8747);
nor U11358 (N_11358,N_9592,N_9246);
or U11359 (N_11359,N_6717,N_8984);
nor U11360 (N_11360,N_7800,N_5138);
xnor U11361 (N_11361,N_5891,N_5125);
nor U11362 (N_11362,N_9721,N_8794);
xor U11363 (N_11363,N_5149,N_9476);
xnor U11364 (N_11364,N_7107,N_6763);
or U11365 (N_11365,N_5793,N_6899);
or U11366 (N_11366,N_5104,N_7688);
or U11367 (N_11367,N_5665,N_9735);
nand U11368 (N_11368,N_6131,N_7500);
xor U11369 (N_11369,N_6389,N_9327);
xor U11370 (N_11370,N_7707,N_7428);
nor U11371 (N_11371,N_7864,N_5351);
and U11372 (N_11372,N_5157,N_6767);
and U11373 (N_11373,N_6781,N_6992);
and U11374 (N_11374,N_5566,N_9809);
nand U11375 (N_11375,N_7565,N_9406);
or U11376 (N_11376,N_7319,N_5014);
or U11377 (N_11377,N_7934,N_5437);
nand U11378 (N_11378,N_9904,N_5815);
xor U11379 (N_11379,N_7726,N_9454);
nand U11380 (N_11380,N_9864,N_7217);
xnor U11381 (N_11381,N_7979,N_8707);
nor U11382 (N_11382,N_6182,N_7614);
nand U11383 (N_11383,N_8532,N_5659);
or U11384 (N_11384,N_5809,N_5461);
and U11385 (N_11385,N_9234,N_8177);
xnor U11386 (N_11386,N_6475,N_7491);
nand U11387 (N_11387,N_8902,N_7282);
nand U11388 (N_11388,N_9365,N_8339);
nor U11389 (N_11389,N_7351,N_7469);
and U11390 (N_11390,N_5024,N_6497);
nor U11391 (N_11391,N_7243,N_5425);
or U11392 (N_11392,N_7712,N_9058);
or U11393 (N_11393,N_5622,N_8556);
nand U11394 (N_11394,N_5527,N_9998);
nand U11395 (N_11395,N_8295,N_9198);
nand U11396 (N_11396,N_8964,N_7402);
xor U11397 (N_11397,N_9997,N_9989);
nand U11398 (N_11398,N_5174,N_5508);
or U11399 (N_11399,N_9578,N_6128);
or U11400 (N_11400,N_6045,N_9579);
or U11401 (N_11401,N_7975,N_6991);
nor U11402 (N_11402,N_6269,N_5086);
and U11403 (N_11403,N_7246,N_5357);
and U11404 (N_11404,N_8020,N_9095);
nand U11405 (N_11405,N_5590,N_8770);
nand U11406 (N_11406,N_7474,N_8876);
xor U11407 (N_11407,N_5794,N_7855);
nand U11408 (N_11408,N_6204,N_7486);
xnor U11409 (N_11409,N_8459,N_7621);
xor U11410 (N_11410,N_8254,N_8542);
nand U11411 (N_11411,N_7453,N_9314);
and U11412 (N_11412,N_9553,N_5731);
xnor U11413 (N_11413,N_6693,N_6704);
nand U11414 (N_11414,N_6262,N_8612);
or U11415 (N_11415,N_7739,N_5032);
nor U11416 (N_11416,N_8500,N_8972);
or U11417 (N_11417,N_7473,N_6687);
nor U11418 (N_11418,N_7424,N_8774);
and U11419 (N_11419,N_9632,N_9976);
xor U11420 (N_11420,N_9682,N_8163);
nor U11421 (N_11421,N_8688,N_7785);
and U11422 (N_11422,N_8363,N_9323);
and U11423 (N_11423,N_8641,N_5708);
nor U11424 (N_11424,N_5213,N_8139);
and U11425 (N_11425,N_5786,N_7421);
nand U11426 (N_11426,N_6273,N_7416);
or U11427 (N_11427,N_7265,N_6721);
or U11428 (N_11428,N_6070,N_5915);
nor U11429 (N_11429,N_5410,N_7200);
nand U11430 (N_11430,N_9166,N_7094);
xnor U11431 (N_11431,N_5098,N_5683);
and U11432 (N_11432,N_6926,N_8361);
xnor U11433 (N_11433,N_7588,N_6493);
nand U11434 (N_11434,N_8133,N_5702);
xnor U11435 (N_11435,N_7581,N_6351);
xor U11436 (N_11436,N_9917,N_8247);
and U11437 (N_11437,N_8988,N_6826);
nand U11438 (N_11438,N_6110,N_8818);
or U11439 (N_11439,N_6044,N_9642);
or U11440 (N_11440,N_5405,N_9614);
or U11441 (N_11441,N_5303,N_9673);
xor U11442 (N_11442,N_5392,N_6129);
and U11443 (N_11443,N_8961,N_6628);
nand U11444 (N_11444,N_5509,N_7329);
and U11445 (N_11445,N_8103,N_7542);
nor U11446 (N_11446,N_7017,N_7573);
xnor U11447 (N_11447,N_5133,N_7773);
xor U11448 (N_11448,N_8771,N_6818);
nand U11449 (N_11449,N_7754,N_9362);
nand U11450 (N_11450,N_6192,N_5193);
nor U11451 (N_11451,N_8344,N_6883);
and U11452 (N_11452,N_6966,N_7129);
and U11453 (N_11453,N_9943,N_5633);
and U11454 (N_11454,N_8898,N_5317);
nand U11455 (N_11455,N_9055,N_9771);
nand U11456 (N_11456,N_8082,N_7660);
and U11457 (N_11457,N_5070,N_9975);
or U11458 (N_11458,N_8387,N_5276);
nand U11459 (N_11459,N_9367,N_5906);
xor U11460 (N_11460,N_5715,N_6089);
nand U11461 (N_11461,N_9769,N_8412);
xor U11462 (N_11462,N_7273,N_5225);
nand U11463 (N_11463,N_7571,N_9143);
xnor U11464 (N_11464,N_9571,N_8578);
nand U11465 (N_11465,N_8491,N_8394);
xnor U11466 (N_11466,N_5238,N_5914);
nor U11467 (N_11467,N_6674,N_5047);
nand U11468 (N_11468,N_5062,N_9251);
nand U11469 (N_11469,N_8116,N_6640);
and U11470 (N_11470,N_7923,N_9785);
nor U11471 (N_11471,N_5592,N_5830);
nor U11472 (N_11472,N_5358,N_6496);
nand U11473 (N_11473,N_7259,N_9865);
nor U11474 (N_11474,N_8783,N_5619);
nor U11475 (N_11475,N_7438,N_6485);
xnor U11476 (N_11476,N_9281,N_9957);
xnor U11477 (N_11477,N_6768,N_8424);
xor U11478 (N_11478,N_6645,N_6049);
nor U11479 (N_11479,N_6419,N_5624);
or U11480 (N_11480,N_5647,N_8086);
or U11481 (N_11481,N_7004,N_5243);
or U11482 (N_11482,N_9113,N_8814);
nor U11483 (N_11483,N_6075,N_6839);
nor U11484 (N_11484,N_5568,N_7179);
and U11485 (N_11485,N_6144,N_9469);
nand U11486 (N_11486,N_7281,N_9094);
xnor U11487 (N_11487,N_5031,N_9544);
or U11488 (N_11488,N_5734,N_5295);
or U11489 (N_11489,N_5962,N_9222);
or U11490 (N_11490,N_5710,N_5348);
and U11491 (N_11491,N_5131,N_5662);
or U11492 (N_11492,N_5824,N_9490);
or U11493 (N_11493,N_5419,N_9724);
xnor U11494 (N_11494,N_8831,N_6022);
xor U11495 (N_11495,N_7037,N_9331);
and U11496 (N_11496,N_6034,N_6159);
nand U11497 (N_11497,N_9039,N_9830);
and U11498 (N_11498,N_8736,N_9539);
xnor U11499 (N_11499,N_6520,N_8129);
nor U11500 (N_11500,N_9183,N_8158);
nand U11501 (N_11501,N_9795,N_8425);
xor U11502 (N_11502,N_7673,N_5183);
nor U11503 (N_11503,N_9466,N_6313);
xnor U11504 (N_11504,N_9437,N_8757);
nand U11505 (N_11505,N_7780,N_6345);
or U11506 (N_11506,N_5924,N_6379);
xnor U11507 (N_11507,N_8743,N_5870);
xor U11508 (N_11508,N_9928,N_9099);
nor U11509 (N_11509,N_5739,N_9261);
nor U11510 (N_11510,N_9025,N_8245);
nor U11511 (N_11511,N_6476,N_7623);
xnor U11512 (N_11512,N_8135,N_8277);
nand U11513 (N_11513,N_6980,N_9554);
or U11514 (N_11514,N_9522,N_6287);
xor U11515 (N_11515,N_7766,N_5588);
or U11516 (N_11516,N_7400,N_8801);
nor U11517 (N_11517,N_5017,N_9669);
and U11518 (N_11518,N_7795,N_5228);
nand U11519 (N_11519,N_6987,N_5783);
nor U11520 (N_11520,N_6705,N_8605);
xnor U11521 (N_11521,N_9503,N_9655);
or U11522 (N_11522,N_9263,N_7880);
nand U11523 (N_11523,N_5926,N_5361);
and U11524 (N_11524,N_7254,N_9828);
and U11525 (N_11525,N_5600,N_7647);
or U11526 (N_11526,N_5543,N_5684);
nand U11527 (N_11527,N_9276,N_7849);
xor U11528 (N_11528,N_8499,N_5841);
xnor U11529 (N_11529,N_5323,N_9439);
nor U11530 (N_11530,N_5169,N_5132);
and U11531 (N_11531,N_9056,N_7727);
or U11532 (N_11532,N_5431,N_8014);
xor U11533 (N_11533,N_6431,N_8546);
nand U11534 (N_11534,N_5167,N_7509);
or U11535 (N_11535,N_7262,N_7162);
nand U11536 (N_11536,N_7523,N_8421);
or U11537 (N_11537,N_9902,N_5327);
or U11538 (N_11538,N_7672,N_7099);
nand U11539 (N_11539,N_6841,N_9624);
nor U11540 (N_11540,N_5012,N_9984);
or U11541 (N_11541,N_6152,N_7019);
xnor U11542 (N_11542,N_7449,N_7286);
or U11543 (N_11543,N_9446,N_6208);
and U11544 (N_11544,N_5945,N_5571);
xor U11545 (N_11545,N_9053,N_5817);
xor U11546 (N_11546,N_7225,N_5618);
xnor U11547 (N_11547,N_7556,N_5730);
and U11548 (N_11548,N_7263,N_7938);
xor U11549 (N_11549,N_9770,N_6240);
or U11550 (N_11550,N_5719,N_6376);
and U11551 (N_11551,N_7154,N_8240);
and U11552 (N_11552,N_6020,N_7711);
or U11553 (N_11553,N_9961,N_5721);
nor U11554 (N_11554,N_5413,N_5034);
or U11555 (N_11555,N_7942,N_5069);
nor U11556 (N_11556,N_6442,N_7536);
and U11557 (N_11557,N_7991,N_7847);
nand U11558 (N_11558,N_9945,N_8596);
xor U11559 (N_11559,N_7481,N_5314);
xnor U11560 (N_11560,N_5704,N_6261);
or U11561 (N_11561,N_5140,N_8140);
or U11562 (N_11562,N_5971,N_7250);
xnor U11563 (N_11563,N_5938,N_5869);
nor U11564 (N_11564,N_8386,N_7807);
nor U11565 (N_11565,N_6584,N_7294);
nor U11566 (N_11566,N_8348,N_9617);
and U11567 (N_11567,N_5293,N_7751);
nor U11568 (N_11568,N_8932,N_6331);
or U11569 (N_11569,N_5496,N_7904);
nor U11570 (N_11570,N_5139,N_9796);
nand U11571 (N_11571,N_9708,N_8154);
and U11572 (N_11572,N_8484,N_7550);
and U11573 (N_11573,N_9781,N_7113);
or U11574 (N_11574,N_6220,N_9328);
nor U11575 (N_11575,N_8305,N_9758);
nor U11576 (N_11576,N_6073,N_7700);
xnor U11577 (N_11577,N_7626,N_6466);
xnor U11578 (N_11578,N_8367,N_7522);
nand U11579 (N_11579,N_6575,N_8230);
nor U11580 (N_11580,N_9330,N_9919);
xor U11581 (N_11581,N_6574,N_6673);
or U11582 (N_11582,N_9000,N_6656);
xnor U11583 (N_11583,N_8463,N_8420);
xor U11584 (N_11584,N_7863,N_8927);
xnor U11585 (N_11585,N_8987,N_9493);
nor U11586 (N_11586,N_9533,N_8672);
nor U11587 (N_11587,N_7696,N_8196);
and U11588 (N_11588,N_8849,N_6978);
xnor U11589 (N_11589,N_9354,N_6742);
and U11590 (N_11590,N_9256,N_6612);
nand U11591 (N_11591,N_9101,N_5452);
nand U11592 (N_11592,N_8081,N_5762);
xnor U11593 (N_11593,N_8931,N_5656);
nand U11594 (N_11594,N_9050,N_8101);
nand U11595 (N_11595,N_8535,N_6245);
and U11596 (N_11596,N_6624,N_8887);
or U11597 (N_11597,N_9168,N_7086);
xnor U11598 (N_11598,N_5423,N_6219);
xnor U11599 (N_11599,N_6879,N_9621);
nor U11600 (N_11600,N_6642,N_8839);
or U11601 (N_11601,N_9889,N_7126);
or U11602 (N_11602,N_7954,N_6784);
nor U11603 (N_11603,N_7563,N_7186);
xor U11604 (N_11604,N_7949,N_5920);
xor U11605 (N_11605,N_5043,N_8317);
nand U11606 (N_11606,N_6660,N_5386);
and U11607 (N_11607,N_5087,N_8035);
or U11608 (N_11608,N_5979,N_6483);
and U11609 (N_11609,N_6213,N_6979);
nand U11610 (N_11610,N_6850,N_7906);
nor U11611 (N_11611,N_7040,N_7935);
nand U11612 (N_11612,N_7378,N_5187);
nand U11613 (N_11613,N_8674,N_5814);
nand U11614 (N_11614,N_5614,N_7235);
and U11615 (N_11615,N_9075,N_9132);
nand U11616 (N_11616,N_6795,N_9552);
nand U11617 (N_11617,N_8253,N_6542);
nor U11618 (N_11618,N_9883,N_8526);
or U11619 (N_11619,N_8975,N_7298);
or U11620 (N_11620,N_5519,N_8263);
nand U11621 (N_11621,N_7087,N_8671);
xnor U11622 (N_11622,N_6852,N_9123);
xor U11623 (N_11623,N_7576,N_8568);
nand U11624 (N_11624,N_5753,N_9131);
and U11625 (N_11625,N_6384,N_9015);
nand U11626 (N_11626,N_7379,N_5576);
and U11627 (N_11627,N_6357,N_6821);
or U11628 (N_11628,N_9916,N_9856);
xnor U11629 (N_11629,N_8219,N_9675);
and U11630 (N_11630,N_5776,N_6427);
nand U11631 (N_11631,N_9117,N_8985);
nand U11632 (N_11632,N_9006,N_7970);
and U11633 (N_11633,N_8011,N_9786);
nor U11634 (N_11634,N_7268,N_9894);
nand U11635 (N_11635,N_6293,N_7526);
nand U11636 (N_11636,N_7895,N_8566);
nor U11637 (N_11637,N_8543,N_8470);
nor U11638 (N_11638,N_9576,N_7210);
and U11639 (N_11639,N_6071,N_5847);
and U11640 (N_11640,N_7663,N_7397);
nand U11641 (N_11641,N_6659,N_6108);
and U11642 (N_11642,N_9267,N_9088);
nand U11643 (N_11643,N_6730,N_7920);
xor U11644 (N_11644,N_5418,N_8648);
nand U11645 (N_11645,N_9231,N_7347);
and U11646 (N_11646,N_5749,N_8657);
nor U11647 (N_11647,N_9034,N_7468);
nor U11648 (N_11648,N_5168,N_5009);
or U11649 (N_11649,N_8100,N_6993);
xnor U11650 (N_11650,N_8803,N_8280);
or U11651 (N_11651,N_5691,N_5969);
nor U11652 (N_11652,N_9318,N_5797);
nor U11653 (N_11653,N_9418,N_7446);
or U11654 (N_11654,N_9270,N_8396);
or U11655 (N_11655,N_9409,N_6851);
or U11656 (N_11656,N_7658,N_9568);
nand U11657 (N_11657,N_5338,N_7706);
nor U11658 (N_11658,N_5720,N_7301);
xor U11659 (N_11659,N_8942,N_9470);
nor U11660 (N_11660,N_6421,N_9236);
nand U11661 (N_11661,N_9924,N_7994);
or U11662 (N_11662,N_9637,N_6154);
xor U11663 (N_11663,N_6663,N_7482);
or U11664 (N_11664,N_5217,N_5154);
xnor U11665 (N_11665,N_5803,N_5985);
or U11666 (N_11666,N_6745,N_6622);
or U11667 (N_11667,N_6927,N_8008);
or U11668 (N_11668,N_5893,N_9907);
and U11669 (N_11669,N_6853,N_9926);
or U11670 (N_11670,N_8825,N_6565);
and U11671 (N_11671,N_9766,N_9639);
or U11672 (N_11672,N_5123,N_5297);
and U11673 (N_11673,N_5038,N_5854);
or U11674 (N_11674,N_9452,N_8756);
nor U11675 (N_11675,N_7253,N_7848);
nand U11676 (N_11676,N_7782,N_6870);
and U11677 (N_11677,N_9558,N_8959);
or U11678 (N_11678,N_9481,N_8922);
or U11679 (N_11679,N_6509,N_8827);
nand U11680 (N_11680,N_8667,N_7070);
nand U11681 (N_11681,N_8513,N_5642);
or U11682 (N_11682,N_8300,N_9666);
nor U11683 (N_11683,N_6364,N_6426);
nand U11684 (N_11684,N_7357,N_6226);
nand U11685 (N_11685,N_8252,N_6714);
nor U11686 (N_11686,N_9179,N_5244);
xor U11687 (N_11687,N_9077,N_8347);
or U11688 (N_11688,N_9150,N_6122);
xor U11689 (N_11689,N_5160,N_9586);
or U11690 (N_11690,N_9017,N_7061);
nor U11691 (N_11691,N_7747,N_7721);
xnor U11692 (N_11692,N_9644,N_7790);
nor U11693 (N_11693,N_6454,N_8607);
nand U11694 (N_11694,N_7425,N_7765);
nand U11695 (N_11695,N_6700,N_9138);
nor U11696 (N_11696,N_6799,N_7407);
or U11697 (N_11697,N_5892,N_5909);
or U11698 (N_11698,N_6709,N_6296);
nor U11699 (N_11699,N_7123,N_9584);
nor U11700 (N_11700,N_5628,N_6672);
nand U11701 (N_11701,N_7076,N_8034);
nor U11702 (N_11702,N_6218,N_5048);
or U11703 (N_11703,N_8695,N_9818);
xor U11704 (N_11704,N_5010,N_7472);
nand U11705 (N_11705,N_9388,N_5903);
or U11706 (N_11706,N_5775,N_9110);
and U11707 (N_11707,N_5083,N_6929);
and U11708 (N_11708,N_8255,N_5958);
nand U11709 (N_11709,N_8371,N_5524);
and U11710 (N_11710,N_5467,N_9543);
or U11711 (N_11711,N_8966,N_9874);
xor U11712 (N_11712,N_8065,N_8881);
xnor U11713 (N_11713,N_6176,N_9736);
or U11714 (N_11714,N_6500,N_9814);
nand U11715 (N_11715,N_9343,N_8937);
nand U11716 (N_11716,N_5391,N_5682);
xor U11717 (N_11717,N_7441,N_6439);
or U11718 (N_11718,N_6312,N_7869);
xnor U11719 (N_11719,N_5251,N_9325);
xor U11720 (N_11720,N_5333,N_8142);
nor U11721 (N_11721,N_5158,N_7214);
xnor U11722 (N_11722,N_9441,N_5219);
nand U11723 (N_11723,N_6535,N_6736);
xor U11724 (N_11724,N_8864,N_7681);
or U11725 (N_11725,N_6563,N_6284);
xor U11726 (N_11726,N_9530,N_9573);
and U11727 (N_11727,N_8074,N_7943);
nand U11728 (N_11728,N_5983,N_8337);
and U11729 (N_11729,N_9999,N_5368);
or U11730 (N_11730,N_6374,N_8710);
xnor U11731 (N_11731,N_6666,N_7144);
nor U11732 (N_11732,N_6059,N_8426);
nor U11733 (N_11733,N_9374,N_8184);
xnor U11734 (N_11734,N_9743,N_7423);
and U11735 (N_11735,N_9321,N_8983);
or U11736 (N_11736,N_9322,N_9723);
nor U11737 (N_11737,N_8155,N_6701);
nor U11738 (N_11738,N_7813,N_9702);
nor U11739 (N_11739,N_7024,N_6646);
nor U11740 (N_11740,N_7511,N_6986);
and U11741 (N_11741,N_6095,N_9585);
or U11742 (N_11742,N_6016,N_8214);
or U11743 (N_11743,N_9557,N_6281);
xnor U11744 (N_11744,N_5300,N_7036);
xor U11745 (N_11745,N_9653,N_9278);
and U11746 (N_11746,N_8152,N_5458);
and U11747 (N_11747,N_8084,N_9607);
xnor U11748 (N_11748,N_6189,N_6734);
and U11749 (N_11749,N_5025,N_5950);
nor U11750 (N_11750,N_6801,N_6241);
or U11751 (N_11751,N_7921,N_8722);
nand U11752 (N_11752,N_7119,N_8851);
and U11753 (N_11753,N_8798,N_7553);
nor U11754 (N_11754,N_7627,N_8575);
nor U11755 (N_11755,N_6074,N_9392);
xor U11756 (N_11756,N_7655,N_7396);
nand U11757 (N_11757,N_8507,N_8248);
xor U11758 (N_11758,N_6005,N_9216);
or U11759 (N_11759,N_6544,N_5373);
or U11760 (N_11760,N_5968,N_6017);
or U11761 (N_11761,N_7399,N_7467);
and U11762 (N_11762,N_6246,N_6094);
xor U11763 (N_11763,N_9173,N_9436);
nor U11764 (N_11764,N_5279,N_6503);
or U11765 (N_11765,N_5007,N_7828);
and U11766 (N_11766,N_6228,N_9120);
or U11767 (N_11767,N_8780,N_5941);
nor U11768 (N_11768,N_8448,N_5988);
or U11769 (N_11769,N_6406,N_8917);
xor U11770 (N_11770,N_5454,N_6422);
xnor U11771 (N_11771,N_8863,N_7541);
nand U11772 (N_11772,N_9760,N_9697);
and U11773 (N_11773,N_6098,N_7023);
or U11774 (N_11774,N_7615,N_7312);
nor U11775 (N_11775,N_8472,N_6458);
nor U11776 (N_11776,N_7910,N_5060);
nor U11777 (N_11777,N_6309,N_8540);
or U11778 (N_11778,N_5252,N_7381);
or U11779 (N_11779,N_6881,N_7946);
xor U11780 (N_11780,N_7743,N_9387);
nor U11781 (N_11781,N_7770,N_6087);
nand U11782 (N_11782,N_8712,N_5861);
or U11783 (N_11783,N_9789,N_8571);
or U11784 (N_11784,N_6450,N_6633);
and U11785 (N_11785,N_9207,N_7977);
xnor U11786 (N_11786,N_5511,N_8525);
xnor U11787 (N_11787,N_5409,N_6453);
xor U11788 (N_11788,N_8580,N_7422);
and U11789 (N_11789,N_6268,N_5001);
xnor U11790 (N_11790,N_7349,N_8028);
xor U11791 (N_11791,N_6026,N_6209);
or U11792 (N_11792,N_8759,N_9240);
nand U11793 (N_11793,N_9175,N_5143);
nand U11794 (N_11794,N_8179,N_8092);
nand U11795 (N_11795,N_9353,N_5329);
or U11796 (N_11796,N_6041,N_9100);
xnor U11797 (N_11797,N_8620,N_6257);
nor U11798 (N_11798,N_6317,N_8714);
or U11799 (N_11799,N_8939,N_8480);
xnor U11800 (N_11800,N_9966,N_8933);
and U11801 (N_11801,N_7124,N_6922);
xnor U11802 (N_11802,N_6874,N_6316);
xor U11803 (N_11803,N_6119,N_9755);
nand U11804 (N_11804,N_5491,N_6639);
or U11805 (N_11805,N_7277,N_6960);
nand U11806 (N_11806,N_9415,N_7834);
or U11807 (N_11807,N_5722,N_6557);
or U11808 (N_11808,N_7980,N_7208);
or U11809 (N_11809,N_9458,N_6942);
xnor U11810 (N_11810,N_7389,N_6347);
nor U11811 (N_11811,N_6541,N_5542);
or U11812 (N_11812,N_7713,N_9748);
or U11813 (N_11813,N_7955,N_8791);
nor U11814 (N_11814,N_9264,N_6989);
and U11815 (N_11815,N_7814,N_6035);
xor U11816 (N_11816,N_6540,N_9472);
xor U11817 (N_11817,N_5531,N_8729);
nand U11818 (N_11818,N_7999,N_8290);
nor U11819 (N_11819,N_9412,N_6012);
and U11820 (N_11820,N_6124,N_8221);
or U11821 (N_11821,N_5931,N_6288);
and U11822 (N_11822,N_9268,N_9906);
xnor U11823 (N_11823,N_9046,N_6830);
nand U11824 (N_11824,N_8273,N_5364);
xnor U11825 (N_11825,N_5136,N_9679);
and U11826 (N_11826,N_9022,N_6604);
xor U11827 (N_11827,N_8256,N_8732);
or U11828 (N_11828,N_7178,N_6062);
nor U11829 (N_11829,N_6976,N_9993);
nand U11830 (N_11830,N_6327,N_6200);
xor U11831 (N_11831,N_5581,N_9084);
nand U11832 (N_11832,N_6465,N_7338);
and U11833 (N_11833,N_9243,N_9750);
and U11834 (N_11834,N_6636,N_5020);
nand U11835 (N_11835,N_9255,N_8416);
and U11836 (N_11836,N_8085,N_6983);
nor U11837 (N_11837,N_9929,N_7096);
nor U11838 (N_11838,N_6583,N_8537);
and U11839 (N_11839,N_8799,N_5551);
nand U11840 (N_11840,N_9670,N_8816);
xor U11841 (N_11841,N_7174,N_9519);
nor U11842 (N_11842,N_5340,N_6372);
and U11843 (N_11843,N_9107,N_9761);
or U11844 (N_11844,N_5723,N_7911);
nand U11845 (N_11845,N_8382,N_6977);
nor U11846 (N_11846,N_8893,N_8234);
or U11847 (N_11847,N_5728,N_9024);
or U11848 (N_11848,N_6764,N_8475);
nand U11849 (N_11849,N_9938,N_6211);
nor U11850 (N_11850,N_6614,N_7662);
xnor U11851 (N_11851,N_9393,N_8423);
or U11852 (N_11852,N_6291,N_7755);
or U11853 (N_11853,N_7412,N_7050);
or U11854 (N_11854,N_9875,N_7148);
and U11855 (N_11855,N_5515,N_8811);
or U11856 (N_11856,N_6930,N_5526);
and U11857 (N_11857,N_7117,N_7815);
and U11858 (N_11858,N_5777,N_7297);
nand U11859 (N_11859,N_8850,N_5675);
nor U11860 (N_11860,N_5652,N_6197);
xor U11861 (N_11861,N_8726,N_9912);
nand U11862 (N_11862,N_6360,N_9193);
or U11863 (N_11863,N_9271,N_8949);
or U11864 (N_11864,N_6451,N_5736);
or U11865 (N_11865,N_7499,N_5355);
xnor U11866 (N_11866,N_6579,N_8627);
and U11867 (N_11867,N_6031,N_9252);
nand U11868 (N_11868,N_7871,N_7020);
xnor U11869 (N_11869,N_9468,N_9982);
nand U11870 (N_11870,N_8993,N_5153);
and U11871 (N_11871,N_8989,N_9447);
nor U11872 (N_11872,N_8567,N_7344);
nor U11873 (N_11873,N_5569,N_5211);
xor U11874 (N_11874,N_8206,N_9574);
xor U11875 (N_11875,N_8579,N_6507);
nand U11876 (N_11876,N_5190,N_5705);
nand U11877 (N_11877,N_5439,N_7704);
and U11878 (N_11878,N_6814,N_7231);
xnor U11879 (N_11879,N_7965,N_7591);
xnor U11880 (N_11880,N_7717,N_6549);
nor U11881 (N_11881,N_8907,N_5376);
or U11882 (N_11882,N_7876,N_6174);
and U11883 (N_11883,N_9616,N_6996);
and U11884 (N_11884,N_7410,N_8479);
nand U11885 (N_11885,N_5818,N_9510);
nand U11886 (N_11886,N_7909,N_7480);
nand U11887 (N_11887,N_9816,N_9451);
nand U11888 (N_11888,N_6242,N_8787);
nor U11889 (N_11889,N_6539,N_5718);
xor U11890 (N_11890,N_8178,N_8836);
xor U11891 (N_11891,N_9561,N_6754);
xnor U11892 (N_11892,N_7978,N_5218);
xnor U11893 (N_11893,N_5075,N_5544);
nor U11894 (N_11894,N_7484,N_6566);
nor U11895 (N_11895,N_9583,N_8452);
nand U11896 (N_11896,N_6760,N_5479);
or U11897 (N_11897,N_6537,N_6424);
and U11898 (N_11898,N_7940,N_7228);
nor U11899 (N_11899,N_5005,N_8915);
xor U11900 (N_11900,N_7304,N_8156);
and U11901 (N_11901,N_8518,N_6737);
nand U11902 (N_11902,N_7808,N_6224);
or U11903 (N_11903,N_7445,N_6130);
nand U11904 (N_11904,N_7944,N_9858);
nand U11905 (N_11905,N_6937,N_5681);
and U11906 (N_11906,N_6905,N_7244);
nor U11907 (N_11907,N_8810,N_6970);
xnor U11908 (N_11908,N_9202,N_8676);
nor U11909 (N_11909,N_7945,N_8621);
and U11910 (N_11910,N_7489,N_7575);
and U11911 (N_11911,N_6914,N_6398);
nand U11912 (N_11912,N_9737,N_5283);
and U11913 (N_11913,N_5843,N_9310);
or U11914 (N_11914,N_6473,N_6600);
nand U11915 (N_11915,N_9817,N_9963);
xor U11916 (N_11916,N_8594,N_5755);
and U11917 (N_11917,N_7278,N_7102);
nand U11918 (N_11918,N_5384,N_7644);
xnor U11919 (N_11919,N_7279,N_6651);
xnor U11920 (N_11920,N_6923,N_7998);
or U11921 (N_11921,N_8952,N_5387);
and U11922 (N_11922,N_9582,N_5677);
or U11923 (N_11923,N_8087,N_9575);
nor U11924 (N_11924,N_7161,N_8727);
nand U11925 (N_11925,N_8052,N_5246);
nor U11926 (N_11926,N_5144,N_8955);
and U11927 (N_11927,N_7962,N_6577);
or U11928 (N_11928,N_9511,N_8118);
and U11929 (N_11929,N_9373,N_8450);
or U11930 (N_11930,N_9386,N_8962);
nor U11931 (N_11931,N_9580,N_8122);
and U11932 (N_11932,N_6649,N_9492);
and U11933 (N_11933,N_6545,N_6057);
xor U11934 (N_11934,N_7369,N_8868);
or U11935 (N_11935,N_9646,N_5781);
and U11936 (N_11936,N_7109,N_7048);
xor U11937 (N_11937,N_6963,N_6394);
nor U11938 (N_11938,N_8768,N_9035);
and U11939 (N_11939,N_8766,N_5743);
nand U11940 (N_11940,N_6139,N_8840);
nor U11941 (N_11941,N_5262,N_7859);
and U11942 (N_11942,N_8478,N_5286);
xor U11943 (N_11943,N_9900,N_6501);
nor U11944 (N_11944,N_7972,N_9931);
or U11945 (N_11945,N_7697,N_9230);
and U11946 (N_11946,N_7841,N_9191);
xor U11947 (N_11947,N_9873,N_6404);
and U11948 (N_11948,N_7763,N_5438);
nor U11949 (N_11949,N_9645,N_7419);
and U11950 (N_11950,N_9759,N_7809);
xnor U11951 (N_11951,N_5107,N_9083);
xor U11952 (N_11952,N_6972,N_9011);
nand U11953 (N_11953,N_7475,N_7224);
nand U11954 (N_11954,N_7345,N_8076);
and U11955 (N_11955,N_8434,N_8618);
or U11956 (N_11956,N_6941,N_7516);
nor U11957 (N_11957,N_6564,N_5918);
nor U11958 (N_11958,N_6578,N_5336);
xnor U11959 (N_11959,N_8124,N_5185);
xor U11960 (N_11960,N_7434,N_8704);
or U11961 (N_11961,N_7925,N_6024);
or U11962 (N_11962,N_7460,N_5383);
xor U11963 (N_11963,N_7190,N_9478);
nand U11964 (N_11964,N_6619,N_7933);
xnor U11965 (N_11965,N_7640,N_7182);
or U11966 (N_11966,N_9040,N_8755);
xor U11967 (N_11967,N_8638,N_9696);
and U11968 (N_11968,N_8049,N_6794);
nand U11969 (N_11969,N_8969,N_8466);
or U11970 (N_11970,N_5916,N_9379);
nand U11971 (N_11971,N_7142,N_5195);
nand U11972 (N_11972,N_7561,N_6582);
xor U11973 (N_11973,N_9720,N_8057);
xor U11974 (N_11974,N_9684,N_6391);
nor U11975 (N_11975,N_6810,N_6796);
nor U11976 (N_11976,N_7062,N_9067);
xor U11977 (N_11977,N_8751,N_9752);
nand U11978 (N_11978,N_6798,N_7041);
nand U11979 (N_11979,N_8569,N_5051);
nor U11980 (N_11980,N_7898,N_8745);
nand U11981 (N_11981,N_5328,N_9425);
or U11982 (N_11982,N_7026,N_9659);
xor U11983 (N_11983,N_9512,N_6789);
and U11984 (N_11984,N_5489,N_6971);
nand U11985 (N_11985,N_9403,N_6603);
and U11986 (N_11986,N_8613,N_7450);
xnor U11987 (N_11987,N_7487,N_8970);
and U11988 (N_11988,N_6793,N_5026);
nor U11989 (N_11989,N_8146,N_9199);
and U11990 (N_11990,N_7534,N_5497);
nand U11991 (N_11991,N_7139,N_8066);
nand U11992 (N_11992,N_5791,N_7568);
xor U11993 (N_11993,N_7009,N_5414);
nor U11994 (N_11994,N_7212,N_6920);
xnor U11995 (N_11995,N_9151,N_7990);
or U11996 (N_11996,N_5449,N_8025);
nor U11997 (N_11997,N_5041,N_9165);
nand U11998 (N_11998,N_8716,N_7877);
nor U11999 (N_11999,N_9130,N_8911);
nor U12000 (N_12000,N_8792,N_5382);
nor U12001 (N_12001,N_8068,N_6895);
or U12002 (N_12002,N_5650,N_8885);
or U12003 (N_12003,N_9690,N_9784);
and U12004 (N_12004,N_5805,N_6083);
nor U12005 (N_12005,N_6065,N_7744);
xnor U12006 (N_12006,N_5637,N_7598);
and U12007 (N_12007,N_6965,N_8365);
nand U12008 (N_12008,N_6260,N_5369);
xor U12009 (N_12009,N_5396,N_5395);
nor U12010 (N_12010,N_8867,N_9400);
nand U12011 (N_12011,N_5472,N_8686);
xnor U12012 (N_12012,N_8790,N_6251);
nand U12013 (N_12013,N_5471,N_9694);
and U12014 (N_12014,N_6809,N_6786);
nor U12015 (N_12015,N_5226,N_6759);
nand U12016 (N_12016,N_8461,N_6825);
or U12017 (N_12017,N_9289,N_9699);
or U12018 (N_12018,N_7068,N_8715);
nand U12019 (N_12019,N_5301,N_6741);
or U12020 (N_12020,N_5837,N_6902);
nand U12021 (N_12021,N_9285,N_6664);
nor U12022 (N_12022,N_8698,N_8782);
xnor U12023 (N_12023,N_8145,N_8510);
xnor U12024 (N_12024,N_7756,N_6383);
nor U12025 (N_12025,N_6771,N_8821);
and U12026 (N_12026,N_8711,N_6148);
nand U12027 (N_12027,N_6641,N_5350);
or U12028 (N_12028,N_9732,N_7083);
nand U12029 (N_12029,N_8539,N_6570);
xnor U12030 (N_12030,N_9728,N_8203);
nor U12031 (N_12031,N_7177,N_9986);
nor U12032 (N_12032,N_6590,N_9861);
nor U12033 (N_12033,N_7255,N_7332);
and U12034 (N_12034,N_6774,N_7669);
xor U12035 (N_12035,N_6153,N_9739);
or U12036 (N_12036,N_8099,N_9662);
nand U12037 (N_12037,N_8593,N_6654);
nand U12038 (N_12038,N_9751,N_9650);
xor U12039 (N_12039,N_9071,N_9753);
nand U12040 (N_12040,N_6762,N_9474);
and U12041 (N_12041,N_7630,N_8615);
nor U12042 (N_12042,N_7296,N_7507);
nand U12043 (N_12043,N_9311,N_9402);
nand U12044 (N_12044,N_5342,N_6819);
nand U12045 (N_12045,N_9648,N_5671);
nand U12046 (N_12046,N_7194,N_6342);
or U12047 (N_12047,N_5027,N_8148);
xor U12048 (N_12048,N_6863,N_7160);
xor U12049 (N_12049,N_8981,N_6025);
nor U12050 (N_12050,N_8740,N_8301);
xor U12051 (N_12051,N_9597,N_9317);
and U12052 (N_12052,N_7666,N_9357);
xnor U12053 (N_12053,N_7524,N_6776);
nor U12054 (N_12054,N_5874,N_9862);
or U12055 (N_12055,N_7693,N_9482);
nor U12056 (N_12056,N_9235,N_5436);
nor U12057 (N_12057,N_8070,N_9627);
or U12058 (N_12058,N_8668,N_8900);
or U12059 (N_12059,N_7137,N_6058);
nand U12060 (N_12060,N_6151,N_9145);
or U12061 (N_12061,N_6536,N_8398);
xnor U12062 (N_12062,N_7917,N_9713);
nor U12063 (N_12063,N_7652,N_7635);
and U12064 (N_12064,N_8541,N_8544);
and U12065 (N_12065,N_8038,N_6298);
nand U12066 (N_12066,N_8043,N_6718);
xor U12067 (N_12067,N_8724,N_8212);
nor U12068 (N_12068,N_6415,N_8883);
nor U12069 (N_12069,N_5510,N_5022);
xnor U12070 (N_12070,N_7308,N_9727);
xor U12071 (N_12071,N_9422,N_5326);
nor U12072 (N_12072,N_7732,N_9211);
and U12073 (N_12073,N_5853,N_6504);
and U12074 (N_12074,N_6952,N_9465);
nor U12075 (N_12075,N_7370,N_9542);
nor U12076 (N_12076,N_6555,N_7030);
xnor U12077 (N_12077,N_8649,N_5851);
nand U12078 (N_12078,N_9801,N_9985);
xor U12079 (N_12079,N_8918,N_8121);
nor U12080 (N_12080,N_5192,N_5977);
nor U12081 (N_12081,N_5540,N_8644);
nor U12082 (N_12082,N_9037,N_6318);
and U12083 (N_12083,N_8924,N_9488);
and U12084 (N_12084,N_5443,N_9950);
xor U12085 (N_12085,N_7538,N_9649);
and U12086 (N_12086,N_5537,N_9042);
nand U12087 (N_12087,N_6203,N_5372);
xor U12088 (N_12088,N_5145,N_9116);
nor U12089 (N_12089,N_9192,N_8226);
nand U12090 (N_12090,N_8614,N_5687);
and U12091 (N_12091,N_6069,N_8765);
nor U12092 (N_12092,N_5859,N_6843);
nor U12093 (N_12093,N_5685,N_8331);
and U12094 (N_12094,N_7791,N_7442);
and U12095 (N_12095,N_7156,N_6433);
xnor U12096 (N_12096,N_5635,N_8856);
nor U12097 (N_12097,N_9375,N_6120);
xnor U12098 (N_12098,N_6860,N_9973);
or U12099 (N_12099,N_6471,N_7236);
nand U12100 (N_12100,N_7496,N_8362);
xor U12101 (N_12101,N_5092,N_6104);
or U12102 (N_12102,N_8193,N_8646);
nor U12103 (N_12103,N_9154,N_9602);
or U12104 (N_12104,N_6135,N_9038);
and U12105 (N_12105,N_5039,N_6028);
or U12106 (N_12106,N_9487,N_9301);
xor U12107 (N_12107,N_7498,N_6052);
xor U12108 (N_12108,N_9677,N_8884);
nand U12109 (N_12109,N_5627,N_7607);
nor U12110 (N_12110,N_8658,N_5049);
xor U12111 (N_12111,N_8640,N_7173);
nor U12112 (N_12112,N_6892,N_8186);
nand U12113 (N_12113,N_8271,N_6708);
and U12114 (N_12114,N_8721,N_8430);
nand U12115 (N_12115,N_7287,N_5973);
or U12116 (N_12116,N_5280,N_7597);
or U12117 (N_12117,N_7066,N_9395);
nor U12118 (N_12118,N_8060,N_6949);
or U12119 (N_12119,N_7100,N_8496);
and U12120 (N_12120,N_7685,N_7233);
nand U12121 (N_12121,N_9569,N_6484);
xor U12122 (N_12122,N_8859,N_8349);
nand U12123 (N_12123,N_9880,N_5645);
and U12124 (N_12124,N_6526,N_5570);
and U12125 (N_12125,N_6329,N_9712);
or U12126 (N_12126,N_5365,N_6343);
xnor U12127 (N_12127,N_9457,N_9449);
nand U12128 (N_12128,N_6027,N_9033);
nand U12129 (N_12129,N_9513,N_9249);
and U12130 (N_12130,N_9860,N_7197);
nand U12131 (N_12131,N_6592,N_6184);
or U12132 (N_12132,N_8456,N_8032);
xor U12133 (N_12133,N_6532,N_8833);
xor U12134 (N_12134,N_9935,N_7366);
and U12135 (N_12135,N_9308,N_9668);
or U12136 (N_12136,N_8071,N_5709);
nand U12137 (N_12137,N_6662,N_8191);
or U12138 (N_12138,N_8905,N_5352);
or U12139 (N_12139,N_8176,N_6448);
nor U12140 (N_12140,N_8930,N_9081);
nand U12141 (N_12141,N_9172,N_5574);
and U12142 (N_12142,N_8664,N_9096);
xor U12143 (N_12143,N_7383,N_8432);
and U12144 (N_12144,N_9001,N_8935);
or U12145 (N_12145,N_6294,N_6913);
xor U12146 (N_12146,N_8549,N_6903);
xnor U12147 (N_12147,N_7302,N_6946);
nand U12148 (N_12148,N_8691,N_7826);
nor U12149 (N_12149,N_6429,N_5518);
nand U12150 (N_12150,N_9835,N_8914);
xor U12151 (N_12151,N_8598,N_7204);
xnor U12152 (N_12152,N_5615,N_8809);
or U12153 (N_12153,N_9854,N_7748);
nand U12154 (N_12154,N_6402,N_7908);
xor U12155 (N_12155,N_7108,N_8570);
and U12156 (N_12156,N_5337,N_7324);
nand U12157 (N_12157,N_7606,N_8728);
or U12158 (N_12158,N_5307,N_5066);
or U12159 (N_12159,N_9389,N_6782);
xor U12160 (N_12160,N_5463,N_9741);
and U12161 (N_12161,N_7905,N_9981);
nor U12162 (N_12162,N_6332,N_7724);
nand U12163 (N_12163,N_8720,N_6101);
xor U12164 (N_12164,N_9220,N_5899);
and U12165 (N_12165,N_6077,N_9676);
xor U12166 (N_12166,N_7583,N_5680);
and U12167 (N_12167,N_5078,N_7603);
and U12168 (N_12168,N_6186,N_8651);
nand U12169 (N_12169,N_7314,N_6527);
nor U12170 (N_12170,N_9547,N_5288);
nor U12171 (N_12171,N_9946,N_6822);
nor U12172 (N_12172,N_5936,N_8617);
or U12173 (N_12173,N_9747,N_9460);
nand U12174 (N_12174,N_9304,N_7387);
nand U12175 (N_12175,N_6416,N_5175);
and U12176 (N_12176,N_7289,N_7594);
or U12177 (N_12177,N_5099,N_6891);
and U12178 (N_12178,N_5335,N_5100);
xor U12179 (N_12179,N_7464,N_8059);
xor U12180 (N_12180,N_5890,N_9811);
or U12181 (N_12181,N_5363,N_7793);
nor U12182 (N_12182,N_5948,N_8873);
nor U12183 (N_12183,N_9111,N_8909);
and U12184 (N_12184,N_7638,N_7714);
nor U12185 (N_12185,N_5029,N_7495);
nand U12186 (N_12186,N_5907,N_5564);
nand U12187 (N_12187,N_6102,N_9842);
nor U12188 (N_12188,N_5857,N_9279);
or U12189 (N_12189,N_5855,N_6147);
nor U12190 (N_12190,N_6973,N_9537);
and U12191 (N_12191,N_6304,N_7230);
or U12192 (N_12192,N_5004,N_8501);
nand U12193 (N_12193,N_7360,N_8659);
nor U12194 (N_12194,N_9831,N_8995);
nand U12195 (N_12195,N_8467,N_7112);
and U12196 (N_12196,N_9665,N_7334);
xor U12197 (N_12197,N_7957,N_9773);
and U12198 (N_12198,N_9018,N_7049);
and U12199 (N_12199,N_8320,N_5398);
nand U12200 (N_12200,N_7346,N_6321);
xor U12201 (N_12201,N_5796,N_5726);
or U12202 (N_12202,N_6690,N_5848);
xnor U12203 (N_12203,N_6127,N_9414);
xnor U12204 (N_12204,N_9878,N_9610);
nand U12205 (N_12205,N_5432,N_7336);
or U12206 (N_12206,N_8826,N_5204);
xor U12207 (N_12207,N_9108,N_6817);
and U12208 (N_12208,N_7348,N_6616);
or U12209 (N_12209,N_6748,N_9364);
nor U12210 (N_12210,N_7115,N_9337);
and U12211 (N_12211,N_5873,N_7452);
nand U12212 (N_12212,N_7354,N_7257);
and U12213 (N_12213,N_6354,N_7525);
and U12214 (N_12214,N_9061,N_7986);
nand U12215 (N_12215,N_8198,N_7012);
or U12216 (N_12216,N_8310,N_9307);
nor U12217 (N_12217,N_5989,N_8697);
xnor U12218 (N_12218,N_5586,N_7578);
nand U12219 (N_12219,N_9303,N_9047);
and U12220 (N_12220,N_8694,N_7643);
xnor U12221 (N_12221,N_9909,N_8039);
or U12222 (N_12222,N_8854,N_8414);
xor U12223 (N_12223,N_9996,N_6072);
xor U12224 (N_12224,N_9341,N_9118);
and U12225 (N_12225,N_6250,N_9532);
nor U12226 (N_12226,N_6236,N_7122);
xor U12227 (N_12227,N_6326,N_8744);
nand U12228 (N_12228,N_6244,N_7209);
nor U12229 (N_12229,N_7781,N_8444);
and U12230 (N_12230,N_7896,N_6050);
xor U12231 (N_12231,N_7303,N_8284);
and U12232 (N_12232,N_8647,N_5966);
or U12233 (N_12233,N_8628,N_7792);
nor U12234 (N_12234,N_7899,N_7340);
and U12235 (N_12235,N_5790,N_5714);
nor U12236 (N_12236,N_6647,N_9027);
xor U12237 (N_12237,N_8948,N_9129);
and U12238 (N_12238,N_5485,N_9819);
nor U12239 (N_12239,N_9693,N_9968);
or U12240 (N_12240,N_9939,N_9944);
or U12241 (N_12241,N_9045,N_6121);
nand U12242 (N_12242,N_6322,N_7044);
or U12243 (N_12243,N_6607,N_8725);
nor U12244 (N_12244,N_5663,N_8343);
nor U12245 (N_12245,N_9988,N_5939);
and U12246 (N_12246,N_5529,N_7384);
nand U12247 (N_12247,N_9298,N_9106);
nand U12248 (N_12248,N_8204,N_5881);
and U12249 (N_12249,N_5747,N_7547);
xnor U12250 (N_12250,N_9158,N_7723);
and U12251 (N_12251,N_7574,N_5507);
and U12252 (N_12252,N_6413,N_8316);
xor U12253 (N_12253,N_8678,N_7764);
nor U12254 (N_12254,N_6757,N_6962);
or U12255 (N_12255,N_9718,N_8533);
xor U12256 (N_12256,N_5669,N_5964);
and U12257 (N_12257,N_9726,N_5599);
or U12258 (N_12258,N_6165,N_6749);
nor U12259 (N_12259,N_7819,N_5082);
and U12260 (N_12260,N_6401,N_5517);
and U12261 (N_12261,N_5356,N_6644);
nor U12262 (N_12262,N_7021,N_7466);
xor U12263 (N_12263,N_8545,N_7678);
xor U12264 (N_12264,N_9169,N_8182);
nand U12265 (N_12265,N_9941,N_8692);
and U12266 (N_12266,N_6166,N_7817);
nand U12267 (N_12267,N_7016,N_9812);
xor U12268 (N_12268,N_8091,N_9195);
xnor U12269 (N_12269,N_5111,N_5103);
xor U12270 (N_12270,N_8504,N_9566);
xnor U12271 (N_12271,N_9068,N_6380);
and U12272 (N_12272,N_7929,N_6338);
nor U12273 (N_12273,N_6528,N_7699);
and U12274 (N_12274,N_5232,N_8894);
nor U12275 (N_12275,N_5196,N_9041);
nand U12276 (N_12276,N_8589,N_6109);
xnor U12277 (N_12277,N_9820,N_5889);
xnor U12278 (N_12278,N_5921,N_8050);
xnor U12279 (N_12279,N_8073,N_5801);
xor U12280 (N_12280,N_7169,N_5152);
nor U12281 (N_12281,N_7811,N_6123);
nand U12282 (N_12282,N_5644,N_6459);
xnor U12283 (N_12283,N_5951,N_7271);
or U12284 (N_12284,N_6420,N_5359);
or U12285 (N_12285,N_7429,N_7930);
nand U12286 (N_12286,N_8415,N_7220);
nand U12287 (N_12287,N_5042,N_6797);
or U12288 (N_12288,N_9855,N_8333);
xor U12289 (N_12289,N_8046,N_6724);
or U12290 (N_12290,N_8334,N_7560);
or U12291 (N_12291,N_9851,N_6285);
or U12292 (N_12292,N_8896,N_7779);
xor U12293 (N_12293,N_7992,N_9689);
xor U12294 (N_12294,N_6514,N_7742);
nor U12295 (N_12295,N_5381,N_6090);
nor U12296 (N_12296,N_6328,N_9782);
or U12297 (N_12297,N_8913,N_7918);
nand U12298 (N_12298,N_5530,N_9185);
nor U12299 (N_12299,N_5829,N_9133);
xor U12300 (N_12300,N_6486,N_5595);
nor U12301 (N_12301,N_5236,N_9411);
nor U12302 (N_12302,N_6252,N_6808);
and U12303 (N_12303,N_9397,N_8819);
xnor U12304 (N_12304,N_5620,N_8161);
xor U12305 (N_12305,N_6747,N_9057);
xnor U12306 (N_12306,N_7035,N_6657);
and U12307 (N_12307,N_7951,N_5277);
or U12308 (N_12308,N_6711,N_7251);
or U12309 (N_12309,N_6388,N_8292);
nor U12310 (N_12310,N_9124,N_7202);
or U12311 (N_12311,N_7865,N_8104);
xnor U12312 (N_12312,N_7010,N_9729);
xor U12313 (N_12313,N_7448,N_5879);
nand U12314 (N_12314,N_6355,N_5910);
nand U12315 (N_12315,N_5800,N_6815);
and U12316 (N_12316,N_9560,N_8368);
and U12317 (N_12317,N_5666,N_7504);
nor U12318 (N_12318,N_8088,N_6707);
and U12319 (N_12319,N_8336,N_5224);
and U12320 (N_12320,N_9221,N_5761);
nor U12321 (N_12321,N_5266,N_7778);
and U12322 (N_12322,N_9525,N_6534);
and U12323 (N_12323,N_6217,N_9114);
nor U12324 (N_12324,N_9927,N_9678);
xnor U12325 (N_12325,N_7816,N_8296);
nand U12326 (N_12326,N_8834,N_9671);
and U12327 (N_12327,N_6679,N_8399);
xor U12328 (N_12328,N_7440,N_6885);
or U12329 (N_12329,N_8561,N_6727);
nor U12330 (N_12330,N_8000,N_9178);
nor U12331 (N_12331,N_7718,N_8733);
or U12332 (N_12332,N_5664,N_8010);
xnor U12333 (N_12333,N_8906,N_7313);
xor U12334 (N_12334,N_8858,N_8321);
nand U12335 (N_12335,N_8315,N_7842);
nand U12336 (N_12336,N_5842,N_7953);
or U12337 (N_12337,N_5241,N_9599);
nor U12338 (N_12338,N_8413,N_7151);
or U12339 (N_12339,N_5716,N_9991);
nand U12340 (N_12340,N_5810,N_7777);
nor U12341 (N_12341,N_9344,N_9742);
or U12342 (N_12342,N_5076,N_7454);
or U12343 (N_12343,N_8974,N_5059);
or U12344 (N_12344,N_9161,N_8210);
xor U12345 (N_12345,N_7461,N_9368);
or U12346 (N_12346,N_5189,N_5385);
xor U12347 (N_12347,N_6631,N_5956);
or U12348 (N_12348,N_9546,N_8294);
and U12349 (N_12349,N_9312,N_9903);
xor U12350 (N_12350,N_5046,N_6446);
or U12351 (N_12351,N_7722,N_5688);
and U12352 (N_12352,N_6594,N_6452);
nor U12353 (N_12353,N_9611,N_7505);
and U12354 (N_12354,N_8565,N_8764);
xor U12355 (N_12355,N_8957,N_7388);
or U12356 (N_12356,N_6216,N_9895);
and U12357 (N_12357,N_6939,N_5013);
and U12358 (N_12358,N_8660,N_8846);
xor U12359 (N_12359,N_9435,N_7915);
or U12360 (N_12360,N_5124,N_7613);
nand U12361 (N_12361,N_7894,N_6599);
and U12362 (N_12362,N_8947,N_6845);
or U12363 (N_12363,N_9299,N_7320);
xor U12364 (N_12364,N_8056,N_8965);
or U12365 (N_12365,N_5523,N_8309);
nor U12366 (N_12366,N_8319,N_7043);
xnor U12367 (N_12367,N_5649,N_8236);
xnor U12368 (N_12368,N_5502,N_6344);
or U12369 (N_12369,N_7901,N_9352);
nor U12370 (N_12370,N_9378,N_6474);
or U12371 (N_12371,N_6898,N_6956);
and U12372 (N_12372,N_9060,N_6695);
nand U12373 (N_12373,N_7241,N_9147);
xor U12374 (N_12374,N_7355,N_8297);
xor U12375 (N_12375,N_7143,N_5898);
nor U12376 (N_12376,N_6638,N_7167);
xor U12377 (N_12377,N_7131,N_5305);
and U12378 (N_12378,N_6436,N_9995);
xor U12379 (N_12379,N_6897,N_6009);
or U12380 (N_12380,N_9109,N_6409);
nor U12381 (N_12381,N_8835,N_5928);
and U12382 (N_12382,N_5202,N_7285);
xnor U12383 (N_12383,N_9691,N_5214);
or U12384 (N_12384,N_5546,N_6481);
nor U12385 (N_12385,N_6667,N_5330);
nand U12386 (N_12386,N_9424,N_8699);
xor U12387 (N_12387,N_9807,N_8718);
nor U12388 (N_12388,N_5430,N_7558);
nand U12389 (N_12389,N_7003,N_8582);
or U12390 (N_12390,N_5616,N_5946);
nand U12391 (N_12391,N_7572,N_7738);
nor U12392 (N_12392,N_8395,N_6054);
or U12393 (N_12393,N_8860,N_6740);
nand U12394 (N_12394,N_6615,N_6777);
nand U12395 (N_12395,N_7600,N_5867);
xnor U12396 (N_12396,N_7692,N_9149);
and U12397 (N_12397,N_8324,N_8865);
nor U12398 (N_12398,N_6512,N_9714);
nor U12399 (N_12399,N_6588,N_9032);
xnor U12400 (N_12400,N_7252,N_8241);
nand U12401 (N_12401,N_8897,N_9604);
xnor U12402 (N_12402,N_5199,N_9901);
or U12403 (N_12403,N_7184,N_9486);
or U12404 (N_12404,N_9896,N_5912);
or U12405 (N_12405,N_5057,N_6339);
nand U12406 (N_12406,N_8037,N_7187);
nand U12407 (N_12407,N_6093,N_5713);
xnor U12408 (N_12408,N_6513,N_7725);
and U12409 (N_12409,N_5532,N_5648);
nand U12410 (N_12410,N_8730,N_8356);
nor U12411 (N_12411,N_6751,N_8029);
nand U12412 (N_12412,N_8293,N_7694);
nor U12413 (N_12413,N_7427,N_7890);
nand U12414 (N_12414,N_5852,N_6569);
or U12415 (N_12415,N_8802,N_9380);
and U12416 (N_12416,N_8717,N_5122);
nor U12417 (N_12417,N_7620,N_9619);
nor U12418 (N_12418,N_8109,N_7862);
xor U12419 (N_12419,N_6831,N_5884);
nand U12420 (N_12420,N_6915,N_5235);
xor U12421 (N_12421,N_8123,N_7028);
nand U12422 (N_12422,N_9654,N_6720);
xor U12423 (N_12423,N_8754,N_9843);
and U12424 (N_12424,N_9087,N_6303);
and U12425 (N_12425,N_5667,N_7709);
or U12426 (N_12426,N_7731,N_7836);
xor U12427 (N_12427,N_5399,N_9232);
or U12428 (N_12428,N_6084,N_8312);
and U12429 (N_12429,N_5538,N_8045);
xor U12430 (N_12430,N_8357,N_5296);
nand U12431 (N_12431,N_9266,N_8004);
and U12432 (N_12432,N_5064,N_8258);
nor U12433 (N_12433,N_8890,N_6271);
nor U12434 (N_12434,N_5740,N_8643);
xnor U12435 (N_12435,N_6247,N_7223);
nand U12436 (N_12436,N_5233,N_7175);
and U12437 (N_12437,N_5813,N_5402);
or U12438 (N_12438,N_6178,N_5389);
xor U12439 (N_12439,N_8131,N_8200);
or U12440 (N_12440,N_9313,N_5812);
nor U12441 (N_12441,N_5555,N_7530);
xnor U12442 (N_12442,N_8773,N_6198);
and U12443 (N_12443,N_8125,N_7218);
and U12444 (N_12444,N_7362,N_6834);
xnor U12445 (N_12445,N_8789,N_8378);
xnor U12446 (N_12446,N_8599,N_8267);
xor U12447 (N_12447,N_6838,N_9382);
xnor U12448 (N_12448,N_9372,N_5116);
or U12449 (N_12449,N_7993,N_8795);
nand U12450 (N_12450,N_5606,N_6457);
nor U12451 (N_12451,N_9069,N_5534);
nor U12452 (N_12452,N_5302,N_7539);
nand U12453 (N_12453,N_6950,N_9410);
nand U12454 (N_12454,N_5506,N_7075);
or U12455 (N_12455,N_8169,N_5759);
or U12456 (N_12456,N_9848,N_8238);
xnor U12457 (N_12457,N_9098,N_7002);
nand U12458 (N_12458,N_9846,N_7769);
nand U12459 (N_12459,N_9839,N_6519);
nor U12460 (N_12460,N_8215,N_8476);
nor U12461 (N_12461,N_5811,N_6307);
nor U12462 (N_12462,N_5832,N_5788);
nor U12463 (N_12463,N_8403,N_7514);
and U12464 (N_12464,N_8573,N_8577);
nand U12465 (N_12465,N_9852,N_8662);
nand U12466 (N_12466,N_8022,N_8862);
xnor U12467 (N_12467,N_5597,N_9351);
and U12468 (N_12468,N_6985,N_6699);
xor U12469 (N_12469,N_8515,N_9443);
and U12470 (N_12470,N_6658,N_8845);
or U12471 (N_12471,N_7705,N_6367);
and U12472 (N_12472,N_6356,N_9004);
xnor U12473 (N_12473,N_9128,N_6082);
nor U12474 (N_12474,N_8134,N_6778);
and U12475 (N_12475,N_8243,N_6945);
nor U12476 (N_12476,N_8797,N_8857);
nor U12477 (N_12477,N_7981,N_5450);
or U12478 (N_12478,N_8042,N_5400);
nor U12479 (N_12479,N_5536,N_5427);
or U12480 (N_12480,N_5208,N_9871);
xnor U12481 (N_12481,N_6115,N_9401);
or U12482 (N_12482,N_7831,N_7527);
or U12483 (N_12483,N_6909,N_9012);
xor U12484 (N_12484,N_7205,N_5724);
and U12485 (N_12485,N_6038,N_8055);
nand U12486 (N_12486,N_6188,N_9020);
nor U12487 (N_12487,N_7787,N_7417);
or U12488 (N_12488,N_9233,N_7554);
nor U12489 (N_12489,N_6464,N_5268);
or U12490 (N_12490,N_6697,N_9242);
nor U12491 (N_12491,N_8581,N_8752);
or U12492 (N_12492,N_5282,N_5094);
nand U12493 (N_12493,N_9915,N_7897);
and U12494 (N_12494,N_9956,N_6733);
and U12495 (N_12495,N_5015,N_5575);
xnor U12496 (N_12496,N_8683,N_5692);
or U12497 (N_12497,N_8033,N_9633);
and U12498 (N_12498,N_5880,N_5016);
or U12499 (N_12499,N_6010,N_6434);
nor U12500 (N_12500,N_5539,N_5049);
and U12501 (N_12501,N_5009,N_7019);
or U12502 (N_12502,N_9409,N_8091);
and U12503 (N_12503,N_7693,N_7588);
and U12504 (N_12504,N_6527,N_5548);
xor U12505 (N_12505,N_7702,N_9833);
nand U12506 (N_12506,N_8037,N_7885);
nor U12507 (N_12507,N_8871,N_8938);
nand U12508 (N_12508,N_5976,N_9844);
xnor U12509 (N_12509,N_8904,N_9369);
xor U12510 (N_12510,N_5079,N_5961);
nand U12511 (N_12511,N_8366,N_7274);
nor U12512 (N_12512,N_7855,N_8086);
and U12513 (N_12513,N_6864,N_5337);
xor U12514 (N_12514,N_8095,N_5166);
xor U12515 (N_12515,N_6979,N_9900);
nor U12516 (N_12516,N_5752,N_8488);
nand U12517 (N_12517,N_6893,N_7504);
nand U12518 (N_12518,N_5689,N_9124);
nand U12519 (N_12519,N_6329,N_9574);
xor U12520 (N_12520,N_8515,N_7306);
or U12521 (N_12521,N_5395,N_5702);
xnor U12522 (N_12522,N_9585,N_7923);
xor U12523 (N_12523,N_5658,N_8963);
and U12524 (N_12524,N_6304,N_7051);
xor U12525 (N_12525,N_7517,N_5581);
and U12526 (N_12526,N_5185,N_7114);
nor U12527 (N_12527,N_5927,N_8084);
nand U12528 (N_12528,N_7815,N_5568);
nor U12529 (N_12529,N_9350,N_9351);
nand U12530 (N_12530,N_9264,N_9434);
and U12531 (N_12531,N_8487,N_7777);
nand U12532 (N_12532,N_9983,N_6153);
nand U12533 (N_12533,N_5037,N_5774);
xor U12534 (N_12534,N_7671,N_5059);
nand U12535 (N_12535,N_5961,N_5258);
nand U12536 (N_12536,N_8721,N_7904);
nor U12537 (N_12537,N_5069,N_6650);
or U12538 (N_12538,N_8011,N_8086);
nor U12539 (N_12539,N_5648,N_9944);
nor U12540 (N_12540,N_6411,N_9947);
xnor U12541 (N_12541,N_9191,N_7671);
nand U12542 (N_12542,N_7059,N_9133);
nor U12543 (N_12543,N_6814,N_8023);
xnor U12544 (N_12544,N_7644,N_6473);
xnor U12545 (N_12545,N_9108,N_7005);
nand U12546 (N_12546,N_8225,N_5864);
nand U12547 (N_12547,N_8014,N_9620);
xor U12548 (N_12548,N_6289,N_8731);
nor U12549 (N_12549,N_6488,N_9923);
and U12550 (N_12550,N_5195,N_8309);
and U12551 (N_12551,N_9333,N_5432);
and U12552 (N_12552,N_9298,N_5235);
nor U12553 (N_12553,N_9537,N_6814);
and U12554 (N_12554,N_5425,N_5895);
or U12555 (N_12555,N_5947,N_7242);
or U12556 (N_12556,N_5643,N_5705);
nand U12557 (N_12557,N_6737,N_7561);
and U12558 (N_12558,N_9101,N_7953);
xnor U12559 (N_12559,N_8872,N_6628);
xnor U12560 (N_12560,N_5516,N_7558);
and U12561 (N_12561,N_8642,N_7779);
nand U12562 (N_12562,N_7234,N_8045);
nor U12563 (N_12563,N_8931,N_5798);
or U12564 (N_12564,N_6559,N_9575);
nand U12565 (N_12565,N_5292,N_8056);
nand U12566 (N_12566,N_5271,N_6612);
and U12567 (N_12567,N_5319,N_6266);
or U12568 (N_12568,N_6862,N_6804);
xor U12569 (N_12569,N_8268,N_5771);
nand U12570 (N_12570,N_7281,N_5471);
xnor U12571 (N_12571,N_5819,N_5721);
or U12572 (N_12572,N_7307,N_6763);
nand U12573 (N_12573,N_6323,N_5318);
or U12574 (N_12574,N_5353,N_9285);
and U12575 (N_12575,N_5012,N_8037);
xor U12576 (N_12576,N_8172,N_9046);
nor U12577 (N_12577,N_6565,N_9213);
and U12578 (N_12578,N_7374,N_5837);
or U12579 (N_12579,N_9183,N_6966);
nand U12580 (N_12580,N_7085,N_5150);
nor U12581 (N_12581,N_8601,N_5745);
or U12582 (N_12582,N_9055,N_9124);
and U12583 (N_12583,N_5645,N_6365);
nand U12584 (N_12584,N_6017,N_8387);
nand U12585 (N_12585,N_8435,N_5072);
xnor U12586 (N_12586,N_5508,N_5215);
or U12587 (N_12587,N_9138,N_9187);
nand U12588 (N_12588,N_5011,N_7810);
nor U12589 (N_12589,N_7529,N_7267);
xnor U12590 (N_12590,N_5009,N_8859);
nor U12591 (N_12591,N_9748,N_8004);
or U12592 (N_12592,N_6329,N_8584);
or U12593 (N_12593,N_7624,N_5371);
nand U12594 (N_12594,N_8455,N_8098);
nand U12595 (N_12595,N_8555,N_8000);
nor U12596 (N_12596,N_7728,N_7879);
nor U12597 (N_12597,N_8606,N_7461);
and U12598 (N_12598,N_9536,N_8077);
nand U12599 (N_12599,N_6013,N_9417);
or U12600 (N_12600,N_7991,N_7238);
xnor U12601 (N_12601,N_8414,N_5240);
nand U12602 (N_12602,N_6913,N_9607);
and U12603 (N_12603,N_9669,N_7010);
xnor U12604 (N_12604,N_8901,N_6051);
or U12605 (N_12605,N_6539,N_8145);
or U12606 (N_12606,N_7149,N_5253);
nor U12607 (N_12607,N_7094,N_6798);
nor U12608 (N_12608,N_7958,N_6119);
xnor U12609 (N_12609,N_9675,N_9221);
nor U12610 (N_12610,N_5573,N_7592);
xor U12611 (N_12611,N_5697,N_5563);
nand U12612 (N_12612,N_5384,N_5019);
nor U12613 (N_12613,N_6567,N_9171);
nor U12614 (N_12614,N_8276,N_5984);
and U12615 (N_12615,N_6058,N_6211);
or U12616 (N_12616,N_8677,N_8551);
nor U12617 (N_12617,N_9498,N_6462);
xor U12618 (N_12618,N_6426,N_5794);
nor U12619 (N_12619,N_7622,N_7477);
and U12620 (N_12620,N_5204,N_5985);
or U12621 (N_12621,N_9411,N_5358);
nor U12622 (N_12622,N_7145,N_5393);
and U12623 (N_12623,N_7516,N_9391);
nor U12624 (N_12624,N_6011,N_7143);
or U12625 (N_12625,N_5292,N_6145);
or U12626 (N_12626,N_5733,N_8551);
xnor U12627 (N_12627,N_6479,N_5545);
or U12628 (N_12628,N_8015,N_9282);
xnor U12629 (N_12629,N_6970,N_8171);
and U12630 (N_12630,N_8339,N_9860);
or U12631 (N_12631,N_5114,N_8979);
and U12632 (N_12632,N_8987,N_5187);
nand U12633 (N_12633,N_9584,N_7909);
or U12634 (N_12634,N_9393,N_8844);
or U12635 (N_12635,N_8923,N_9646);
and U12636 (N_12636,N_5104,N_5496);
nor U12637 (N_12637,N_8728,N_8242);
xnor U12638 (N_12638,N_5962,N_5747);
nand U12639 (N_12639,N_8923,N_7132);
xor U12640 (N_12640,N_6295,N_8211);
and U12641 (N_12641,N_8809,N_6579);
nand U12642 (N_12642,N_5201,N_8495);
nor U12643 (N_12643,N_5574,N_7045);
xor U12644 (N_12644,N_5127,N_8510);
xnor U12645 (N_12645,N_7492,N_5846);
nor U12646 (N_12646,N_6602,N_7520);
and U12647 (N_12647,N_9287,N_9954);
nor U12648 (N_12648,N_9495,N_9321);
or U12649 (N_12649,N_5711,N_5419);
nor U12650 (N_12650,N_9936,N_5064);
nor U12651 (N_12651,N_5178,N_5010);
or U12652 (N_12652,N_5641,N_8815);
or U12653 (N_12653,N_9591,N_7877);
nor U12654 (N_12654,N_7396,N_6784);
nor U12655 (N_12655,N_8413,N_9549);
and U12656 (N_12656,N_5113,N_6975);
and U12657 (N_12657,N_9138,N_8134);
nand U12658 (N_12658,N_7355,N_7130);
nand U12659 (N_12659,N_5243,N_8335);
or U12660 (N_12660,N_6876,N_8218);
nor U12661 (N_12661,N_6292,N_5076);
xnor U12662 (N_12662,N_6491,N_8123);
nor U12663 (N_12663,N_9605,N_8774);
and U12664 (N_12664,N_8147,N_5839);
xor U12665 (N_12665,N_5292,N_6661);
xnor U12666 (N_12666,N_9223,N_9026);
and U12667 (N_12667,N_9494,N_5057);
nand U12668 (N_12668,N_6361,N_6082);
and U12669 (N_12669,N_8386,N_8754);
xor U12670 (N_12670,N_6921,N_6469);
nor U12671 (N_12671,N_7589,N_8085);
or U12672 (N_12672,N_6888,N_6235);
and U12673 (N_12673,N_6878,N_9262);
xnor U12674 (N_12674,N_7452,N_8532);
xnor U12675 (N_12675,N_8373,N_8417);
nand U12676 (N_12676,N_6866,N_7382);
xnor U12677 (N_12677,N_7487,N_9702);
nor U12678 (N_12678,N_7426,N_6473);
or U12679 (N_12679,N_6292,N_8926);
nand U12680 (N_12680,N_9605,N_5542);
xnor U12681 (N_12681,N_6358,N_5908);
nor U12682 (N_12682,N_5083,N_9989);
nand U12683 (N_12683,N_9046,N_6257);
nand U12684 (N_12684,N_5524,N_9364);
xor U12685 (N_12685,N_5592,N_7287);
or U12686 (N_12686,N_8977,N_9292);
xor U12687 (N_12687,N_5298,N_7362);
or U12688 (N_12688,N_9459,N_5588);
or U12689 (N_12689,N_7723,N_6505);
or U12690 (N_12690,N_8724,N_8806);
nor U12691 (N_12691,N_9582,N_7717);
and U12692 (N_12692,N_9918,N_8111);
nor U12693 (N_12693,N_8975,N_9127);
xor U12694 (N_12694,N_9372,N_5471);
nand U12695 (N_12695,N_7257,N_7170);
and U12696 (N_12696,N_8720,N_8039);
and U12697 (N_12697,N_9470,N_8946);
or U12698 (N_12698,N_7301,N_9978);
xnor U12699 (N_12699,N_8104,N_6154);
xor U12700 (N_12700,N_9733,N_7859);
and U12701 (N_12701,N_6404,N_7564);
nand U12702 (N_12702,N_8106,N_8828);
nor U12703 (N_12703,N_9699,N_8441);
or U12704 (N_12704,N_9899,N_8587);
nand U12705 (N_12705,N_6228,N_6775);
or U12706 (N_12706,N_8044,N_8591);
nand U12707 (N_12707,N_8187,N_9236);
nor U12708 (N_12708,N_6099,N_6098);
nor U12709 (N_12709,N_5370,N_7502);
nor U12710 (N_12710,N_9958,N_6985);
xnor U12711 (N_12711,N_9168,N_5529);
xnor U12712 (N_12712,N_9666,N_5440);
nor U12713 (N_12713,N_9376,N_7424);
xor U12714 (N_12714,N_5101,N_9791);
nor U12715 (N_12715,N_8350,N_5237);
nand U12716 (N_12716,N_5833,N_5244);
nor U12717 (N_12717,N_6970,N_5118);
nor U12718 (N_12718,N_6131,N_9115);
nand U12719 (N_12719,N_7037,N_8858);
nor U12720 (N_12720,N_7169,N_9153);
and U12721 (N_12721,N_8386,N_6350);
nor U12722 (N_12722,N_7767,N_6156);
or U12723 (N_12723,N_5377,N_9427);
xnor U12724 (N_12724,N_8374,N_5621);
nand U12725 (N_12725,N_5431,N_8775);
xnor U12726 (N_12726,N_5637,N_9162);
nand U12727 (N_12727,N_9468,N_8141);
and U12728 (N_12728,N_9375,N_8619);
or U12729 (N_12729,N_9661,N_6523);
nor U12730 (N_12730,N_9464,N_7908);
nor U12731 (N_12731,N_6996,N_6314);
nand U12732 (N_12732,N_7822,N_5035);
and U12733 (N_12733,N_8074,N_6805);
xnor U12734 (N_12734,N_7500,N_7390);
nor U12735 (N_12735,N_9001,N_9389);
nor U12736 (N_12736,N_6405,N_5838);
or U12737 (N_12737,N_6671,N_6577);
and U12738 (N_12738,N_8196,N_5221);
xor U12739 (N_12739,N_8009,N_6883);
and U12740 (N_12740,N_7486,N_9715);
nor U12741 (N_12741,N_5485,N_5509);
or U12742 (N_12742,N_7455,N_5401);
nor U12743 (N_12743,N_6008,N_7328);
nand U12744 (N_12744,N_7593,N_5827);
nor U12745 (N_12745,N_7448,N_5040);
and U12746 (N_12746,N_5707,N_5172);
nand U12747 (N_12747,N_7454,N_5842);
nand U12748 (N_12748,N_6862,N_6653);
nand U12749 (N_12749,N_8692,N_5910);
xnor U12750 (N_12750,N_8565,N_9012);
and U12751 (N_12751,N_9333,N_6172);
xor U12752 (N_12752,N_5730,N_6304);
nor U12753 (N_12753,N_8782,N_9648);
nor U12754 (N_12754,N_8940,N_6715);
and U12755 (N_12755,N_6599,N_8904);
and U12756 (N_12756,N_8019,N_6654);
xnor U12757 (N_12757,N_5436,N_6213);
xor U12758 (N_12758,N_5543,N_6868);
nor U12759 (N_12759,N_9047,N_6044);
xor U12760 (N_12760,N_6953,N_9673);
nand U12761 (N_12761,N_8308,N_7866);
nand U12762 (N_12762,N_5017,N_6053);
nor U12763 (N_12763,N_9339,N_6487);
xor U12764 (N_12764,N_9030,N_7683);
xnor U12765 (N_12765,N_7296,N_5843);
nand U12766 (N_12766,N_8177,N_6665);
and U12767 (N_12767,N_8638,N_8182);
nor U12768 (N_12768,N_5858,N_8964);
nor U12769 (N_12769,N_9885,N_7641);
and U12770 (N_12770,N_8941,N_5704);
nor U12771 (N_12771,N_5208,N_5753);
nand U12772 (N_12772,N_7422,N_7310);
and U12773 (N_12773,N_5403,N_5581);
or U12774 (N_12774,N_7875,N_8523);
nor U12775 (N_12775,N_5010,N_6244);
or U12776 (N_12776,N_7436,N_8908);
or U12777 (N_12777,N_5316,N_7911);
and U12778 (N_12778,N_5496,N_8362);
nor U12779 (N_12779,N_5942,N_6068);
nand U12780 (N_12780,N_9708,N_9585);
nand U12781 (N_12781,N_7692,N_5208);
xor U12782 (N_12782,N_5786,N_7473);
and U12783 (N_12783,N_8339,N_8487);
or U12784 (N_12784,N_6454,N_5426);
nor U12785 (N_12785,N_5832,N_5409);
nand U12786 (N_12786,N_6325,N_6801);
nor U12787 (N_12787,N_6206,N_6058);
or U12788 (N_12788,N_6950,N_9405);
nor U12789 (N_12789,N_6709,N_7505);
or U12790 (N_12790,N_7478,N_6994);
and U12791 (N_12791,N_6684,N_5752);
xor U12792 (N_12792,N_5151,N_8212);
nor U12793 (N_12793,N_7220,N_6351);
and U12794 (N_12794,N_7521,N_7139);
xnor U12795 (N_12795,N_6388,N_8022);
and U12796 (N_12796,N_9890,N_5286);
xor U12797 (N_12797,N_9945,N_9911);
or U12798 (N_12798,N_6250,N_9265);
nor U12799 (N_12799,N_7391,N_7559);
and U12800 (N_12800,N_8739,N_9038);
nand U12801 (N_12801,N_6212,N_6659);
or U12802 (N_12802,N_9580,N_8114);
nor U12803 (N_12803,N_5690,N_8014);
or U12804 (N_12804,N_9183,N_5036);
xor U12805 (N_12805,N_5885,N_7650);
nor U12806 (N_12806,N_6815,N_9148);
nor U12807 (N_12807,N_9734,N_6659);
xor U12808 (N_12808,N_5200,N_7627);
xnor U12809 (N_12809,N_7690,N_6571);
nand U12810 (N_12810,N_7300,N_5217);
and U12811 (N_12811,N_6376,N_6544);
nand U12812 (N_12812,N_7194,N_7704);
or U12813 (N_12813,N_6590,N_6663);
nor U12814 (N_12814,N_5834,N_6407);
and U12815 (N_12815,N_5274,N_6233);
nand U12816 (N_12816,N_9242,N_6155);
or U12817 (N_12817,N_8678,N_5165);
nor U12818 (N_12818,N_8292,N_9653);
and U12819 (N_12819,N_8895,N_9968);
or U12820 (N_12820,N_8234,N_8543);
xor U12821 (N_12821,N_6409,N_7551);
nand U12822 (N_12822,N_9658,N_5696);
nand U12823 (N_12823,N_9318,N_6412);
nand U12824 (N_12824,N_7387,N_5492);
xnor U12825 (N_12825,N_7337,N_5763);
nand U12826 (N_12826,N_5595,N_5437);
nand U12827 (N_12827,N_6322,N_8895);
nor U12828 (N_12828,N_8542,N_8340);
xnor U12829 (N_12829,N_8079,N_9086);
nand U12830 (N_12830,N_5353,N_8426);
xor U12831 (N_12831,N_8008,N_8089);
nand U12832 (N_12832,N_9453,N_7413);
nor U12833 (N_12833,N_6035,N_5765);
xor U12834 (N_12834,N_7932,N_8786);
or U12835 (N_12835,N_8687,N_9169);
and U12836 (N_12836,N_7567,N_6849);
nor U12837 (N_12837,N_9686,N_9437);
nor U12838 (N_12838,N_7637,N_7229);
nand U12839 (N_12839,N_5981,N_8351);
xor U12840 (N_12840,N_6998,N_8630);
nor U12841 (N_12841,N_8825,N_5762);
and U12842 (N_12842,N_9421,N_7467);
and U12843 (N_12843,N_7592,N_9559);
and U12844 (N_12844,N_8365,N_9249);
nor U12845 (N_12845,N_9408,N_6827);
nor U12846 (N_12846,N_6604,N_7721);
or U12847 (N_12847,N_9553,N_6487);
nand U12848 (N_12848,N_9703,N_7091);
nor U12849 (N_12849,N_5636,N_5036);
or U12850 (N_12850,N_6495,N_8658);
nand U12851 (N_12851,N_8643,N_6442);
nor U12852 (N_12852,N_6436,N_7972);
or U12853 (N_12853,N_6201,N_5275);
and U12854 (N_12854,N_9496,N_8913);
and U12855 (N_12855,N_9596,N_7379);
xor U12856 (N_12856,N_6167,N_6424);
xor U12857 (N_12857,N_6318,N_5276);
nor U12858 (N_12858,N_6423,N_7552);
or U12859 (N_12859,N_7445,N_9632);
and U12860 (N_12860,N_6470,N_7764);
nand U12861 (N_12861,N_5121,N_8590);
nor U12862 (N_12862,N_7294,N_6880);
or U12863 (N_12863,N_6080,N_6101);
nand U12864 (N_12864,N_9154,N_6150);
or U12865 (N_12865,N_9093,N_8734);
nor U12866 (N_12866,N_8094,N_9843);
nor U12867 (N_12867,N_6535,N_6769);
nor U12868 (N_12868,N_6210,N_5086);
xor U12869 (N_12869,N_9301,N_5602);
nor U12870 (N_12870,N_8402,N_5808);
nor U12871 (N_12871,N_5204,N_6508);
nor U12872 (N_12872,N_8677,N_7523);
xor U12873 (N_12873,N_6613,N_7495);
nand U12874 (N_12874,N_8200,N_5683);
and U12875 (N_12875,N_8539,N_9540);
xnor U12876 (N_12876,N_6430,N_9907);
xnor U12877 (N_12877,N_5579,N_7012);
nand U12878 (N_12878,N_6821,N_5273);
and U12879 (N_12879,N_7399,N_7581);
xor U12880 (N_12880,N_9540,N_8801);
xor U12881 (N_12881,N_5699,N_5455);
nor U12882 (N_12882,N_7950,N_6195);
nor U12883 (N_12883,N_5497,N_8104);
nor U12884 (N_12884,N_5768,N_8554);
nor U12885 (N_12885,N_6787,N_9457);
nand U12886 (N_12886,N_8018,N_8038);
and U12887 (N_12887,N_5250,N_8912);
and U12888 (N_12888,N_7952,N_5177);
and U12889 (N_12889,N_8531,N_6985);
and U12890 (N_12890,N_9417,N_6485);
or U12891 (N_12891,N_6279,N_9530);
or U12892 (N_12892,N_8300,N_7939);
or U12893 (N_12893,N_5192,N_7287);
xor U12894 (N_12894,N_6165,N_8487);
or U12895 (N_12895,N_7705,N_7554);
or U12896 (N_12896,N_7382,N_9284);
nor U12897 (N_12897,N_9660,N_8463);
nand U12898 (N_12898,N_9615,N_5295);
nand U12899 (N_12899,N_7945,N_9593);
or U12900 (N_12900,N_8562,N_7311);
nor U12901 (N_12901,N_5185,N_7833);
or U12902 (N_12902,N_5464,N_6770);
xor U12903 (N_12903,N_8495,N_6463);
nor U12904 (N_12904,N_6018,N_7231);
xor U12905 (N_12905,N_5522,N_7790);
nor U12906 (N_12906,N_9017,N_6649);
xor U12907 (N_12907,N_6545,N_9566);
xnor U12908 (N_12908,N_8866,N_6158);
nand U12909 (N_12909,N_5451,N_5884);
or U12910 (N_12910,N_5620,N_7822);
xor U12911 (N_12911,N_9404,N_9066);
nor U12912 (N_12912,N_8969,N_9048);
nor U12913 (N_12913,N_9064,N_7616);
or U12914 (N_12914,N_9987,N_6396);
nor U12915 (N_12915,N_7503,N_5446);
or U12916 (N_12916,N_5392,N_9599);
or U12917 (N_12917,N_6273,N_8994);
xnor U12918 (N_12918,N_9688,N_5446);
or U12919 (N_12919,N_9566,N_8561);
and U12920 (N_12920,N_6368,N_8071);
nor U12921 (N_12921,N_9226,N_8599);
and U12922 (N_12922,N_5557,N_5638);
nor U12923 (N_12923,N_7969,N_9444);
or U12924 (N_12924,N_7235,N_8445);
or U12925 (N_12925,N_8657,N_8831);
xor U12926 (N_12926,N_8098,N_9376);
nand U12927 (N_12927,N_6068,N_9389);
xor U12928 (N_12928,N_5889,N_7514);
nand U12929 (N_12929,N_9677,N_5976);
nand U12930 (N_12930,N_9268,N_7559);
nor U12931 (N_12931,N_9947,N_6987);
xor U12932 (N_12932,N_8623,N_5158);
and U12933 (N_12933,N_6610,N_9081);
nor U12934 (N_12934,N_7866,N_7898);
nand U12935 (N_12935,N_7139,N_6219);
or U12936 (N_12936,N_8754,N_7814);
nor U12937 (N_12937,N_6467,N_7619);
xor U12938 (N_12938,N_9754,N_7060);
nand U12939 (N_12939,N_9037,N_8552);
and U12940 (N_12940,N_6746,N_6273);
nand U12941 (N_12941,N_8787,N_5596);
and U12942 (N_12942,N_8558,N_5094);
xor U12943 (N_12943,N_5451,N_7084);
nand U12944 (N_12944,N_8093,N_8608);
nand U12945 (N_12945,N_9213,N_9033);
xnor U12946 (N_12946,N_6882,N_8571);
nor U12947 (N_12947,N_7619,N_7169);
xnor U12948 (N_12948,N_6722,N_9943);
nand U12949 (N_12949,N_5236,N_7532);
xnor U12950 (N_12950,N_5181,N_8719);
or U12951 (N_12951,N_5523,N_6506);
and U12952 (N_12952,N_6307,N_6884);
nor U12953 (N_12953,N_6049,N_7880);
and U12954 (N_12954,N_9125,N_9515);
xor U12955 (N_12955,N_6270,N_7976);
xor U12956 (N_12956,N_5241,N_6866);
xor U12957 (N_12957,N_7175,N_7240);
or U12958 (N_12958,N_8665,N_6870);
or U12959 (N_12959,N_9114,N_5611);
and U12960 (N_12960,N_5244,N_8944);
or U12961 (N_12961,N_8297,N_5008);
and U12962 (N_12962,N_8613,N_6969);
nand U12963 (N_12963,N_9073,N_6890);
xor U12964 (N_12964,N_9931,N_6609);
nor U12965 (N_12965,N_8309,N_7124);
nand U12966 (N_12966,N_7641,N_5781);
xor U12967 (N_12967,N_8497,N_6367);
xor U12968 (N_12968,N_6315,N_6173);
xor U12969 (N_12969,N_5868,N_7588);
and U12970 (N_12970,N_8855,N_5733);
or U12971 (N_12971,N_9696,N_9119);
xor U12972 (N_12972,N_5634,N_9886);
xor U12973 (N_12973,N_6756,N_9446);
xor U12974 (N_12974,N_8246,N_5947);
and U12975 (N_12975,N_8970,N_8634);
or U12976 (N_12976,N_7120,N_9266);
nand U12977 (N_12977,N_5601,N_9616);
or U12978 (N_12978,N_9579,N_7136);
or U12979 (N_12979,N_9850,N_5981);
or U12980 (N_12980,N_7719,N_5040);
xnor U12981 (N_12981,N_5575,N_7408);
nor U12982 (N_12982,N_5580,N_9398);
or U12983 (N_12983,N_5475,N_5397);
nor U12984 (N_12984,N_5318,N_9017);
or U12985 (N_12985,N_8397,N_9119);
and U12986 (N_12986,N_7540,N_9132);
and U12987 (N_12987,N_7052,N_7890);
nor U12988 (N_12988,N_9361,N_9244);
and U12989 (N_12989,N_5164,N_5215);
or U12990 (N_12990,N_8600,N_7389);
nor U12991 (N_12991,N_8322,N_9466);
xor U12992 (N_12992,N_8576,N_6218);
or U12993 (N_12993,N_7395,N_5849);
nand U12994 (N_12994,N_9123,N_6342);
or U12995 (N_12995,N_8651,N_8885);
and U12996 (N_12996,N_9296,N_8747);
xor U12997 (N_12997,N_5432,N_8212);
nand U12998 (N_12998,N_8494,N_8746);
nor U12999 (N_12999,N_6551,N_5788);
nor U13000 (N_13000,N_8749,N_6269);
or U13001 (N_13001,N_8085,N_9970);
or U13002 (N_13002,N_9979,N_9376);
and U13003 (N_13003,N_7349,N_6817);
or U13004 (N_13004,N_5610,N_8630);
nand U13005 (N_13005,N_6391,N_8170);
or U13006 (N_13006,N_8095,N_6791);
nand U13007 (N_13007,N_6608,N_5494);
xnor U13008 (N_13008,N_9138,N_6681);
or U13009 (N_13009,N_8310,N_8764);
nand U13010 (N_13010,N_9792,N_8137);
xnor U13011 (N_13011,N_5628,N_9206);
and U13012 (N_13012,N_6501,N_7608);
nand U13013 (N_13013,N_9934,N_5771);
and U13014 (N_13014,N_8614,N_7021);
and U13015 (N_13015,N_7903,N_7757);
nor U13016 (N_13016,N_9289,N_7166);
or U13017 (N_13017,N_9454,N_8849);
nor U13018 (N_13018,N_7813,N_5327);
and U13019 (N_13019,N_5521,N_9973);
xnor U13020 (N_13020,N_5004,N_6503);
xnor U13021 (N_13021,N_9837,N_9418);
and U13022 (N_13022,N_8085,N_7059);
nand U13023 (N_13023,N_5174,N_7600);
nor U13024 (N_13024,N_8421,N_8603);
and U13025 (N_13025,N_9802,N_7506);
and U13026 (N_13026,N_9903,N_8811);
nand U13027 (N_13027,N_8923,N_8096);
or U13028 (N_13028,N_9096,N_6463);
nor U13029 (N_13029,N_7333,N_6937);
xnor U13030 (N_13030,N_9437,N_8660);
nand U13031 (N_13031,N_7737,N_7828);
nor U13032 (N_13032,N_8317,N_9854);
nor U13033 (N_13033,N_7922,N_7779);
or U13034 (N_13034,N_7630,N_9474);
nor U13035 (N_13035,N_9725,N_9496);
or U13036 (N_13036,N_9037,N_7116);
or U13037 (N_13037,N_8645,N_6119);
and U13038 (N_13038,N_9193,N_7499);
xor U13039 (N_13039,N_7314,N_5307);
and U13040 (N_13040,N_6521,N_8974);
or U13041 (N_13041,N_5510,N_7991);
nand U13042 (N_13042,N_9865,N_8894);
nor U13043 (N_13043,N_5590,N_7323);
nand U13044 (N_13044,N_5745,N_9817);
and U13045 (N_13045,N_9539,N_9821);
or U13046 (N_13046,N_6931,N_7803);
xnor U13047 (N_13047,N_8228,N_7133);
and U13048 (N_13048,N_9227,N_8838);
nor U13049 (N_13049,N_7283,N_6578);
nand U13050 (N_13050,N_6687,N_9613);
nand U13051 (N_13051,N_5432,N_7294);
and U13052 (N_13052,N_8653,N_5469);
nand U13053 (N_13053,N_5904,N_7947);
or U13054 (N_13054,N_8523,N_8106);
and U13055 (N_13055,N_9015,N_7057);
nand U13056 (N_13056,N_5526,N_5215);
nor U13057 (N_13057,N_6786,N_8394);
and U13058 (N_13058,N_5617,N_9762);
nor U13059 (N_13059,N_7022,N_5419);
nor U13060 (N_13060,N_5821,N_6550);
nand U13061 (N_13061,N_6423,N_5952);
nor U13062 (N_13062,N_5869,N_7403);
xor U13063 (N_13063,N_6997,N_9972);
xnor U13064 (N_13064,N_6331,N_5508);
or U13065 (N_13065,N_5197,N_8698);
or U13066 (N_13066,N_6364,N_6111);
or U13067 (N_13067,N_6826,N_5510);
nor U13068 (N_13068,N_5018,N_8756);
nor U13069 (N_13069,N_9648,N_8386);
and U13070 (N_13070,N_7181,N_5255);
nand U13071 (N_13071,N_7699,N_7012);
nor U13072 (N_13072,N_7346,N_5630);
and U13073 (N_13073,N_5072,N_8159);
xor U13074 (N_13074,N_9916,N_6958);
or U13075 (N_13075,N_9379,N_6335);
or U13076 (N_13076,N_9852,N_9312);
nor U13077 (N_13077,N_5187,N_9011);
nand U13078 (N_13078,N_5682,N_6850);
nor U13079 (N_13079,N_7318,N_5244);
xor U13080 (N_13080,N_7191,N_6906);
or U13081 (N_13081,N_8766,N_7737);
nor U13082 (N_13082,N_6886,N_5412);
and U13083 (N_13083,N_9530,N_7755);
or U13084 (N_13084,N_6277,N_6477);
and U13085 (N_13085,N_7378,N_5306);
xor U13086 (N_13086,N_8049,N_7002);
nor U13087 (N_13087,N_7849,N_5113);
nand U13088 (N_13088,N_5203,N_9076);
and U13089 (N_13089,N_7823,N_8035);
and U13090 (N_13090,N_8378,N_6415);
nand U13091 (N_13091,N_7577,N_6091);
or U13092 (N_13092,N_7708,N_7407);
and U13093 (N_13093,N_7052,N_5023);
and U13094 (N_13094,N_7827,N_6961);
xor U13095 (N_13095,N_6532,N_6933);
xnor U13096 (N_13096,N_8094,N_6638);
nor U13097 (N_13097,N_9031,N_9096);
and U13098 (N_13098,N_7919,N_9089);
nor U13099 (N_13099,N_7981,N_5979);
and U13100 (N_13100,N_8793,N_8291);
or U13101 (N_13101,N_8364,N_7448);
or U13102 (N_13102,N_5699,N_5008);
and U13103 (N_13103,N_9729,N_6381);
and U13104 (N_13104,N_7687,N_8955);
nand U13105 (N_13105,N_7348,N_6271);
or U13106 (N_13106,N_8209,N_7494);
or U13107 (N_13107,N_5451,N_8739);
nand U13108 (N_13108,N_5746,N_8789);
and U13109 (N_13109,N_9145,N_6957);
and U13110 (N_13110,N_9732,N_7827);
and U13111 (N_13111,N_5510,N_6484);
xor U13112 (N_13112,N_7198,N_7173);
or U13113 (N_13113,N_7661,N_8745);
nor U13114 (N_13114,N_5627,N_7469);
nor U13115 (N_13115,N_9277,N_8045);
nand U13116 (N_13116,N_8950,N_5954);
and U13117 (N_13117,N_9746,N_8995);
xnor U13118 (N_13118,N_8670,N_9389);
xnor U13119 (N_13119,N_5618,N_6028);
and U13120 (N_13120,N_6006,N_9293);
nand U13121 (N_13121,N_5776,N_8732);
and U13122 (N_13122,N_6484,N_9216);
nand U13123 (N_13123,N_7103,N_6455);
nand U13124 (N_13124,N_5659,N_6766);
nor U13125 (N_13125,N_6811,N_5575);
nand U13126 (N_13126,N_5380,N_8239);
xor U13127 (N_13127,N_9720,N_9548);
nor U13128 (N_13128,N_9343,N_7085);
xnor U13129 (N_13129,N_8681,N_6715);
xnor U13130 (N_13130,N_7730,N_7742);
or U13131 (N_13131,N_8245,N_7239);
nand U13132 (N_13132,N_5363,N_7744);
xor U13133 (N_13133,N_7374,N_5112);
or U13134 (N_13134,N_8210,N_9519);
and U13135 (N_13135,N_8294,N_9663);
nand U13136 (N_13136,N_5047,N_9163);
xor U13137 (N_13137,N_7322,N_5520);
or U13138 (N_13138,N_5574,N_6795);
or U13139 (N_13139,N_5809,N_6733);
nand U13140 (N_13140,N_7489,N_9883);
and U13141 (N_13141,N_7035,N_5782);
nor U13142 (N_13142,N_8295,N_9148);
xor U13143 (N_13143,N_5394,N_6005);
nor U13144 (N_13144,N_8111,N_8924);
and U13145 (N_13145,N_9439,N_5166);
xor U13146 (N_13146,N_6369,N_6382);
nand U13147 (N_13147,N_7856,N_6214);
and U13148 (N_13148,N_8442,N_9752);
or U13149 (N_13149,N_8720,N_5313);
and U13150 (N_13150,N_7308,N_5272);
nand U13151 (N_13151,N_8788,N_6258);
nor U13152 (N_13152,N_5983,N_5423);
or U13153 (N_13153,N_6841,N_5574);
xnor U13154 (N_13154,N_5685,N_6532);
xor U13155 (N_13155,N_6134,N_6315);
nand U13156 (N_13156,N_9967,N_8346);
nand U13157 (N_13157,N_7574,N_5554);
or U13158 (N_13158,N_5352,N_8189);
xnor U13159 (N_13159,N_5964,N_5713);
nand U13160 (N_13160,N_6834,N_9948);
and U13161 (N_13161,N_9995,N_8472);
or U13162 (N_13162,N_9450,N_9080);
or U13163 (N_13163,N_9792,N_6613);
nand U13164 (N_13164,N_5578,N_6001);
nand U13165 (N_13165,N_8076,N_5333);
and U13166 (N_13166,N_9390,N_9858);
nand U13167 (N_13167,N_5282,N_8765);
xnor U13168 (N_13168,N_8125,N_5346);
or U13169 (N_13169,N_5679,N_7911);
and U13170 (N_13170,N_8772,N_6892);
nor U13171 (N_13171,N_8451,N_6103);
or U13172 (N_13172,N_5747,N_5293);
and U13173 (N_13173,N_6112,N_7796);
nor U13174 (N_13174,N_5054,N_7797);
nand U13175 (N_13175,N_6223,N_8834);
nor U13176 (N_13176,N_8525,N_9192);
nand U13177 (N_13177,N_9959,N_9776);
nor U13178 (N_13178,N_8650,N_8970);
or U13179 (N_13179,N_5175,N_6143);
and U13180 (N_13180,N_6979,N_6112);
or U13181 (N_13181,N_7916,N_6654);
or U13182 (N_13182,N_5358,N_7860);
xnor U13183 (N_13183,N_5584,N_9908);
xnor U13184 (N_13184,N_5375,N_6618);
xor U13185 (N_13185,N_9457,N_8882);
nand U13186 (N_13186,N_9366,N_8042);
xor U13187 (N_13187,N_5196,N_6929);
nand U13188 (N_13188,N_6861,N_6752);
nand U13189 (N_13189,N_8279,N_8953);
and U13190 (N_13190,N_5994,N_9837);
or U13191 (N_13191,N_7097,N_5419);
or U13192 (N_13192,N_6901,N_7424);
nor U13193 (N_13193,N_7164,N_7117);
nor U13194 (N_13194,N_6261,N_8609);
or U13195 (N_13195,N_5747,N_8953);
and U13196 (N_13196,N_7401,N_6409);
nor U13197 (N_13197,N_8734,N_9721);
or U13198 (N_13198,N_5460,N_8948);
or U13199 (N_13199,N_9641,N_7814);
xnor U13200 (N_13200,N_5484,N_9055);
or U13201 (N_13201,N_7523,N_9421);
and U13202 (N_13202,N_6660,N_8892);
nand U13203 (N_13203,N_9326,N_6670);
nor U13204 (N_13204,N_7545,N_9158);
or U13205 (N_13205,N_8423,N_5485);
nor U13206 (N_13206,N_6400,N_7781);
nor U13207 (N_13207,N_6870,N_7449);
nand U13208 (N_13208,N_8340,N_7652);
or U13209 (N_13209,N_8131,N_8804);
and U13210 (N_13210,N_6964,N_6561);
nor U13211 (N_13211,N_6079,N_7383);
xor U13212 (N_13212,N_5771,N_6949);
xnor U13213 (N_13213,N_6079,N_8268);
or U13214 (N_13214,N_7335,N_6387);
and U13215 (N_13215,N_6523,N_5307);
and U13216 (N_13216,N_6842,N_8642);
and U13217 (N_13217,N_8037,N_9460);
or U13218 (N_13218,N_7865,N_6492);
xor U13219 (N_13219,N_6813,N_8846);
or U13220 (N_13220,N_5333,N_5155);
and U13221 (N_13221,N_5111,N_8210);
nand U13222 (N_13222,N_7089,N_8071);
nor U13223 (N_13223,N_5961,N_9875);
and U13224 (N_13224,N_5381,N_8844);
nand U13225 (N_13225,N_8871,N_8256);
and U13226 (N_13226,N_6964,N_8017);
nand U13227 (N_13227,N_8896,N_6879);
nor U13228 (N_13228,N_7220,N_9742);
nand U13229 (N_13229,N_9786,N_5701);
nand U13230 (N_13230,N_6954,N_9656);
nor U13231 (N_13231,N_7412,N_9870);
nor U13232 (N_13232,N_5589,N_9142);
and U13233 (N_13233,N_9210,N_9661);
nor U13234 (N_13234,N_9379,N_5500);
or U13235 (N_13235,N_7814,N_6299);
nor U13236 (N_13236,N_9011,N_8509);
xnor U13237 (N_13237,N_9127,N_9946);
xor U13238 (N_13238,N_6285,N_9997);
xnor U13239 (N_13239,N_6418,N_6767);
and U13240 (N_13240,N_8381,N_8613);
and U13241 (N_13241,N_7728,N_8451);
nor U13242 (N_13242,N_9772,N_7220);
xnor U13243 (N_13243,N_7027,N_6669);
or U13244 (N_13244,N_5552,N_9989);
nor U13245 (N_13245,N_6926,N_9670);
nor U13246 (N_13246,N_5387,N_7088);
and U13247 (N_13247,N_7634,N_9547);
and U13248 (N_13248,N_8200,N_7289);
nand U13249 (N_13249,N_8973,N_5654);
nand U13250 (N_13250,N_7610,N_7482);
and U13251 (N_13251,N_5979,N_8941);
xor U13252 (N_13252,N_6366,N_7116);
and U13253 (N_13253,N_6347,N_9406);
nand U13254 (N_13254,N_8886,N_6427);
and U13255 (N_13255,N_7159,N_5671);
and U13256 (N_13256,N_8079,N_8411);
or U13257 (N_13257,N_7242,N_6188);
and U13258 (N_13258,N_5279,N_8838);
and U13259 (N_13259,N_6880,N_5896);
nor U13260 (N_13260,N_9415,N_5463);
and U13261 (N_13261,N_5941,N_8257);
nor U13262 (N_13262,N_7743,N_8443);
nor U13263 (N_13263,N_8675,N_9358);
and U13264 (N_13264,N_9449,N_8779);
or U13265 (N_13265,N_5808,N_6465);
xnor U13266 (N_13266,N_8817,N_9811);
xor U13267 (N_13267,N_6841,N_7380);
or U13268 (N_13268,N_9233,N_7141);
or U13269 (N_13269,N_5502,N_5944);
and U13270 (N_13270,N_5635,N_7745);
nor U13271 (N_13271,N_8456,N_9686);
nor U13272 (N_13272,N_9340,N_8655);
xor U13273 (N_13273,N_6467,N_8897);
and U13274 (N_13274,N_5299,N_9162);
nor U13275 (N_13275,N_9360,N_6943);
or U13276 (N_13276,N_6825,N_8927);
nor U13277 (N_13277,N_9649,N_5113);
or U13278 (N_13278,N_9602,N_6394);
nand U13279 (N_13279,N_5117,N_7384);
nand U13280 (N_13280,N_5479,N_9249);
nor U13281 (N_13281,N_9291,N_9640);
nand U13282 (N_13282,N_9539,N_7640);
xor U13283 (N_13283,N_9763,N_9243);
and U13284 (N_13284,N_5471,N_6750);
or U13285 (N_13285,N_7553,N_9046);
or U13286 (N_13286,N_9665,N_5676);
or U13287 (N_13287,N_6923,N_6843);
nand U13288 (N_13288,N_6042,N_9861);
or U13289 (N_13289,N_6992,N_5805);
nor U13290 (N_13290,N_9102,N_6540);
or U13291 (N_13291,N_5411,N_8121);
xnor U13292 (N_13292,N_9949,N_5292);
xnor U13293 (N_13293,N_6575,N_7807);
xnor U13294 (N_13294,N_7998,N_8990);
nand U13295 (N_13295,N_6761,N_7257);
and U13296 (N_13296,N_5326,N_9579);
nor U13297 (N_13297,N_7879,N_5728);
nand U13298 (N_13298,N_7698,N_7884);
nand U13299 (N_13299,N_6464,N_8590);
or U13300 (N_13300,N_8493,N_5108);
xor U13301 (N_13301,N_7721,N_6767);
nor U13302 (N_13302,N_6756,N_5338);
nor U13303 (N_13303,N_8721,N_5137);
nand U13304 (N_13304,N_6060,N_8927);
nor U13305 (N_13305,N_8852,N_7361);
xnor U13306 (N_13306,N_5147,N_7079);
and U13307 (N_13307,N_9781,N_9979);
or U13308 (N_13308,N_6526,N_8976);
xnor U13309 (N_13309,N_5553,N_6533);
nand U13310 (N_13310,N_8252,N_5942);
nand U13311 (N_13311,N_6770,N_8860);
nor U13312 (N_13312,N_6238,N_7252);
nor U13313 (N_13313,N_8143,N_8440);
or U13314 (N_13314,N_8607,N_6956);
xnor U13315 (N_13315,N_6734,N_6476);
and U13316 (N_13316,N_6349,N_9806);
xnor U13317 (N_13317,N_6999,N_9880);
nand U13318 (N_13318,N_9682,N_7872);
nor U13319 (N_13319,N_5256,N_9863);
nand U13320 (N_13320,N_5096,N_6643);
xnor U13321 (N_13321,N_6576,N_6589);
xor U13322 (N_13322,N_7379,N_8622);
xnor U13323 (N_13323,N_8680,N_7422);
nand U13324 (N_13324,N_9852,N_6251);
nor U13325 (N_13325,N_8676,N_7565);
or U13326 (N_13326,N_5975,N_7647);
xnor U13327 (N_13327,N_9475,N_9501);
or U13328 (N_13328,N_5577,N_8066);
xor U13329 (N_13329,N_5407,N_7225);
and U13330 (N_13330,N_7042,N_7343);
and U13331 (N_13331,N_7597,N_9792);
xor U13332 (N_13332,N_7008,N_9122);
nand U13333 (N_13333,N_9382,N_5926);
and U13334 (N_13334,N_9642,N_7016);
xnor U13335 (N_13335,N_8842,N_9250);
nand U13336 (N_13336,N_8184,N_9194);
xnor U13337 (N_13337,N_7001,N_9415);
or U13338 (N_13338,N_5641,N_9138);
xnor U13339 (N_13339,N_8586,N_6586);
and U13340 (N_13340,N_6504,N_8582);
xor U13341 (N_13341,N_5063,N_6522);
or U13342 (N_13342,N_6326,N_8483);
nand U13343 (N_13343,N_5402,N_6427);
and U13344 (N_13344,N_8548,N_7146);
nand U13345 (N_13345,N_7338,N_7430);
and U13346 (N_13346,N_6050,N_8964);
or U13347 (N_13347,N_6558,N_7250);
nand U13348 (N_13348,N_5180,N_6944);
and U13349 (N_13349,N_6487,N_6668);
nand U13350 (N_13350,N_8237,N_6572);
nand U13351 (N_13351,N_9230,N_9448);
nand U13352 (N_13352,N_5873,N_5161);
or U13353 (N_13353,N_9369,N_8615);
or U13354 (N_13354,N_8929,N_9427);
nor U13355 (N_13355,N_5943,N_5809);
xor U13356 (N_13356,N_8203,N_5656);
nor U13357 (N_13357,N_5622,N_8387);
or U13358 (N_13358,N_8990,N_6712);
xor U13359 (N_13359,N_8597,N_9302);
nor U13360 (N_13360,N_6627,N_6894);
nand U13361 (N_13361,N_9433,N_5616);
xnor U13362 (N_13362,N_7357,N_6012);
or U13363 (N_13363,N_8710,N_8468);
nand U13364 (N_13364,N_9247,N_9762);
xnor U13365 (N_13365,N_9050,N_7045);
nand U13366 (N_13366,N_9085,N_5661);
or U13367 (N_13367,N_9357,N_7507);
nor U13368 (N_13368,N_9768,N_7765);
xnor U13369 (N_13369,N_8694,N_7161);
nand U13370 (N_13370,N_5725,N_5474);
nor U13371 (N_13371,N_7309,N_5416);
nor U13372 (N_13372,N_5999,N_9867);
nand U13373 (N_13373,N_7716,N_8115);
or U13374 (N_13374,N_8678,N_7487);
xor U13375 (N_13375,N_5915,N_8922);
and U13376 (N_13376,N_7896,N_7241);
xnor U13377 (N_13377,N_5922,N_9033);
or U13378 (N_13378,N_7569,N_8495);
or U13379 (N_13379,N_5901,N_9760);
nor U13380 (N_13380,N_7298,N_9776);
nor U13381 (N_13381,N_9715,N_6470);
xor U13382 (N_13382,N_9958,N_7954);
nor U13383 (N_13383,N_7907,N_6763);
nand U13384 (N_13384,N_5976,N_6504);
and U13385 (N_13385,N_7548,N_6043);
and U13386 (N_13386,N_5076,N_8301);
nor U13387 (N_13387,N_6583,N_6794);
xnor U13388 (N_13388,N_8369,N_7494);
or U13389 (N_13389,N_9779,N_7143);
nor U13390 (N_13390,N_5650,N_8583);
nand U13391 (N_13391,N_7300,N_8758);
xor U13392 (N_13392,N_6145,N_7483);
or U13393 (N_13393,N_7890,N_6891);
nand U13394 (N_13394,N_9515,N_6477);
xor U13395 (N_13395,N_8610,N_6814);
nand U13396 (N_13396,N_9156,N_6436);
xor U13397 (N_13397,N_9418,N_8123);
nor U13398 (N_13398,N_9744,N_7769);
nor U13399 (N_13399,N_9666,N_9650);
xor U13400 (N_13400,N_5795,N_9249);
nand U13401 (N_13401,N_8011,N_9279);
xor U13402 (N_13402,N_9327,N_7009);
nand U13403 (N_13403,N_5227,N_6899);
xor U13404 (N_13404,N_5471,N_9467);
nand U13405 (N_13405,N_5618,N_9615);
xor U13406 (N_13406,N_8239,N_7007);
or U13407 (N_13407,N_9388,N_8542);
nand U13408 (N_13408,N_5209,N_5884);
nand U13409 (N_13409,N_6846,N_5438);
and U13410 (N_13410,N_7642,N_7115);
xor U13411 (N_13411,N_9686,N_6233);
nor U13412 (N_13412,N_5247,N_8263);
xor U13413 (N_13413,N_6242,N_8184);
or U13414 (N_13414,N_8865,N_5561);
nor U13415 (N_13415,N_6862,N_6237);
or U13416 (N_13416,N_6710,N_6851);
or U13417 (N_13417,N_5762,N_8212);
nor U13418 (N_13418,N_5130,N_6612);
nand U13419 (N_13419,N_9459,N_7176);
nand U13420 (N_13420,N_7416,N_7009);
or U13421 (N_13421,N_5056,N_5260);
and U13422 (N_13422,N_9844,N_7245);
nand U13423 (N_13423,N_9486,N_7916);
nor U13424 (N_13424,N_8054,N_8339);
nand U13425 (N_13425,N_6601,N_5516);
or U13426 (N_13426,N_9209,N_6575);
xor U13427 (N_13427,N_7404,N_6629);
and U13428 (N_13428,N_5490,N_9993);
or U13429 (N_13429,N_5430,N_7114);
and U13430 (N_13430,N_6633,N_8709);
nand U13431 (N_13431,N_5458,N_7172);
nand U13432 (N_13432,N_9066,N_6138);
or U13433 (N_13433,N_5032,N_5204);
nor U13434 (N_13434,N_9099,N_9365);
and U13435 (N_13435,N_5532,N_9337);
and U13436 (N_13436,N_9575,N_9308);
nand U13437 (N_13437,N_8598,N_5939);
nor U13438 (N_13438,N_8825,N_8115);
nand U13439 (N_13439,N_7034,N_8363);
nor U13440 (N_13440,N_6285,N_8096);
nor U13441 (N_13441,N_8678,N_9529);
nand U13442 (N_13442,N_7223,N_5245);
nand U13443 (N_13443,N_6480,N_8452);
or U13444 (N_13444,N_8514,N_5044);
nand U13445 (N_13445,N_7447,N_8897);
xor U13446 (N_13446,N_8864,N_7824);
and U13447 (N_13447,N_7400,N_5868);
nor U13448 (N_13448,N_6472,N_5253);
or U13449 (N_13449,N_5119,N_9758);
and U13450 (N_13450,N_5148,N_6629);
or U13451 (N_13451,N_7935,N_7130);
nand U13452 (N_13452,N_6875,N_9699);
xor U13453 (N_13453,N_8695,N_9768);
nor U13454 (N_13454,N_8165,N_6678);
and U13455 (N_13455,N_6637,N_6572);
or U13456 (N_13456,N_8609,N_9204);
or U13457 (N_13457,N_6545,N_8539);
or U13458 (N_13458,N_7019,N_5869);
nor U13459 (N_13459,N_7053,N_6471);
and U13460 (N_13460,N_8396,N_8164);
nor U13461 (N_13461,N_7217,N_8280);
nand U13462 (N_13462,N_9223,N_9986);
nand U13463 (N_13463,N_5976,N_6712);
nand U13464 (N_13464,N_9918,N_5397);
and U13465 (N_13465,N_9172,N_6088);
nor U13466 (N_13466,N_8619,N_6998);
xor U13467 (N_13467,N_6218,N_6176);
nor U13468 (N_13468,N_8560,N_6542);
or U13469 (N_13469,N_9660,N_5414);
and U13470 (N_13470,N_9324,N_6562);
and U13471 (N_13471,N_7002,N_5303);
and U13472 (N_13472,N_6599,N_8282);
nand U13473 (N_13473,N_8538,N_6078);
or U13474 (N_13474,N_6796,N_5187);
nand U13475 (N_13475,N_7186,N_6372);
or U13476 (N_13476,N_8403,N_6649);
xnor U13477 (N_13477,N_5393,N_8889);
or U13478 (N_13478,N_9690,N_7693);
or U13479 (N_13479,N_8330,N_8095);
xnor U13480 (N_13480,N_6632,N_7682);
xnor U13481 (N_13481,N_6369,N_9139);
or U13482 (N_13482,N_8157,N_5001);
nand U13483 (N_13483,N_8543,N_8321);
xnor U13484 (N_13484,N_7136,N_7812);
or U13485 (N_13485,N_8230,N_5557);
nand U13486 (N_13486,N_7220,N_7439);
and U13487 (N_13487,N_9094,N_9450);
and U13488 (N_13488,N_6960,N_8433);
and U13489 (N_13489,N_7531,N_5992);
or U13490 (N_13490,N_9409,N_8089);
and U13491 (N_13491,N_9621,N_5050);
xor U13492 (N_13492,N_8829,N_5719);
or U13493 (N_13493,N_7214,N_5797);
xnor U13494 (N_13494,N_5172,N_5537);
and U13495 (N_13495,N_8828,N_6576);
nand U13496 (N_13496,N_7991,N_9357);
and U13497 (N_13497,N_8475,N_6521);
nor U13498 (N_13498,N_9342,N_8455);
nor U13499 (N_13499,N_9762,N_5766);
xor U13500 (N_13500,N_6382,N_5950);
nor U13501 (N_13501,N_5469,N_5900);
or U13502 (N_13502,N_5918,N_8069);
nor U13503 (N_13503,N_9296,N_9444);
nor U13504 (N_13504,N_5889,N_5491);
xor U13505 (N_13505,N_5841,N_9162);
nor U13506 (N_13506,N_8980,N_8235);
xor U13507 (N_13507,N_7559,N_7383);
nor U13508 (N_13508,N_5837,N_8367);
nand U13509 (N_13509,N_5666,N_7497);
or U13510 (N_13510,N_5396,N_7876);
nand U13511 (N_13511,N_5319,N_6844);
nand U13512 (N_13512,N_5503,N_8186);
nor U13513 (N_13513,N_7582,N_9433);
nand U13514 (N_13514,N_5435,N_9208);
or U13515 (N_13515,N_6629,N_8634);
nand U13516 (N_13516,N_6718,N_7988);
nor U13517 (N_13517,N_8173,N_8606);
xor U13518 (N_13518,N_8135,N_9621);
nand U13519 (N_13519,N_5775,N_9859);
nor U13520 (N_13520,N_8308,N_9878);
xor U13521 (N_13521,N_6253,N_7184);
and U13522 (N_13522,N_6257,N_7808);
nor U13523 (N_13523,N_5106,N_9425);
nand U13524 (N_13524,N_8424,N_6016);
and U13525 (N_13525,N_7919,N_5395);
nor U13526 (N_13526,N_5204,N_7106);
nor U13527 (N_13527,N_9039,N_9022);
nand U13528 (N_13528,N_7645,N_5448);
xor U13529 (N_13529,N_7623,N_7313);
or U13530 (N_13530,N_7644,N_7875);
nand U13531 (N_13531,N_8352,N_6585);
nand U13532 (N_13532,N_7579,N_5799);
or U13533 (N_13533,N_5119,N_7562);
nor U13534 (N_13534,N_5600,N_8504);
nor U13535 (N_13535,N_7347,N_8704);
xnor U13536 (N_13536,N_6105,N_8882);
and U13537 (N_13537,N_6581,N_7868);
and U13538 (N_13538,N_6612,N_5471);
and U13539 (N_13539,N_9895,N_8967);
nor U13540 (N_13540,N_7547,N_6001);
and U13541 (N_13541,N_6476,N_5331);
xnor U13542 (N_13542,N_7328,N_6437);
nor U13543 (N_13543,N_5432,N_5445);
and U13544 (N_13544,N_5989,N_7132);
xnor U13545 (N_13545,N_8562,N_8971);
xnor U13546 (N_13546,N_6364,N_5444);
xnor U13547 (N_13547,N_5129,N_7334);
or U13548 (N_13548,N_7946,N_9030);
and U13549 (N_13549,N_7556,N_8972);
nor U13550 (N_13550,N_8053,N_8210);
or U13551 (N_13551,N_9423,N_7180);
nand U13552 (N_13552,N_5915,N_6864);
nor U13553 (N_13553,N_9433,N_9933);
xnor U13554 (N_13554,N_5828,N_5105);
xor U13555 (N_13555,N_8565,N_5030);
xnor U13556 (N_13556,N_8273,N_8426);
and U13557 (N_13557,N_5205,N_9326);
nor U13558 (N_13558,N_7083,N_5277);
nor U13559 (N_13559,N_8625,N_8602);
xor U13560 (N_13560,N_8406,N_7715);
nor U13561 (N_13561,N_7756,N_9303);
xor U13562 (N_13562,N_9623,N_5804);
nand U13563 (N_13563,N_6119,N_6468);
nand U13564 (N_13564,N_6676,N_9989);
nand U13565 (N_13565,N_7871,N_8241);
nand U13566 (N_13566,N_5172,N_7736);
or U13567 (N_13567,N_8251,N_6239);
nand U13568 (N_13568,N_9828,N_7759);
and U13569 (N_13569,N_8160,N_5923);
and U13570 (N_13570,N_5990,N_8071);
xnor U13571 (N_13571,N_6328,N_8667);
and U13572 (N_13572,N_7539,N_5467);
or U13573 (N_13573,N_6639,N_6752);
or U13574 (N_13574,N_8070,N_9408);
or U13575 (N_13575,N_5865,N_8973);
or U13576 (N_13576,N_9307,N_8550);
and U13577 (N_13577,N_9781,N_8088);
nor U13578 (N_13578,N_5582,N_7043);
nand U13579 (N_13579,N_6751,N_5401);
xor U13580 (N_13580,N_8192,N_8436);
and U13581 (N_13581,N_6419,N_7602);
nor U13582 (N_13582,N_8022,N_9301);
xnor U13583 (N_13583,N_8964,N_7567);
or U13584 (N_13584,N_6953,N_6844);
and U13585 (N_13585,N_6553,N_6009);
xor U13586 (N_13586,N_7775,N_5125);
and U13587 (N_13587,N_5450,N_8131);
or U13588 (N_13588,N_6394,N_8568);
and U13589 (N_13589,N_5626,N_5024);
and U13590 (N_13590,N_6225,N_9766);
nand U13591 (N_13591,N_9985,N_7903);
xor U13592 (N_13592,N_7547,N_5248);
nand U13593 (N_13593,N_6007,N_7174);
nand U13594 (N_13594,N_7627,N_9534);
nor U13595 (N_13595,N_7903,N_6483);
xnor U13596 (N_13596,N_9600,N_5059);
and U13597 (N_13597,N_5003,N_9068);
or U13598 (N_13598,N_7096,N_7461);
or U13599 (N_13599,N_5950,N_9455);
xor U13600 (N_13600,N_5754,N_5916);
nor U13601 (N_13601,N_8586,N_8375);
and U13602 (N_13602,N_6283,N_6043);
nor U13603 (N_13603,N_5800,N_6894);
nand U13604 (N_13604,N_5597,N_8257);
nor U13605 (N_13605,N_7173,N_9372);
or U13606 (N_13606,N_6661,N_5817);
nand U13607 (N_13607,N_5637,N_5252);
nand U13608 (N_13608,N_6570,N_6330);
nor U13609 (N_13609,N_7946,N_9793);
nand U13610 (N_13610,N_6219,N_8076);
nor U13611 (N_13611,N_8173,N_6740);
and U13612 (N_13612,N_7027,N_8459);
and U13613 (N_13613,N_9513,N_5089);
nand U13614 (N_13614,N_6420,N_5202);
xor U13615 (N_13615,N_6442,N_6128);
nand U13616 (N_13616,N_8555,N_8489);
and U13617 (N_13617,N_6968,N_5669);
nand U13618 (N_13618,N_7995,N_9712);
or U13619 (N_13619,N_7041,N_8648);
or U13620 (N_13620,N_7143,N_8006);
nor U13621 (N_13621,N_7699,N_5083);
xnor U13622 (N_13622,N_9954,N_5204);
nand U13623 (N_13623,N_7119,N_5529);
xnor U13624 (N_13624,N_5918,N_6227);
nor U13625 (N_13625,N_6250,N_8391);
xor U13626 (N_13626,N_6955,N_9917);
and U13627 (N_13627,N_7602,N_5778);
and U13628 (N_13628,N_7900,N_6123);
xnor U13629 (N_13629,N_5114,N_5058);
and U13630 (N_13630,N_5877,N_6917);
nor U13631 (N_13631,N_6816,N_5071);
nand U13632 (N_13632,N_8232,N_6015);
xnor U13633 (N_13633,N_5168,N_6641);
xor U13634 (N_13634,N_6611,N_8412);
xnor U13635 (N_13635,N_6377,N_7330);
and U13636 (N_13636,N_6361,N_6244);
or U13637 (N_13637,N_8289,N_5663);
nor U13638 (N_13638,N_6647,N_7780);
nand U13639 (N_13639,N_9332,N_8084);
xor U13640 (N_13640,N_5109,N_6101);
xor U13641 (N_13641,N_6558,N_9582);
nor U13642 (N_13642,N_9049,N_6190);
or U13643 (N_13643,N_6688,N_5691);
and U13644 (N_13644,N_7695,N_6281);
nor U13645 (N_13645,N_5239,N_8032);
nand U13646 (N_13646,N_6509,N_5605);
nand U13647 (N_13647,N_5997,N_5514);
nand U13648 (N_13648,N_7391,N_6264);
or U13649 (N_13649,N_9221,N_5670);
xnor U13650 (N_13650,N_7082,N_9588);
nand U13651 (N_13651,N_8717,N_7342);
nand U13652 (N_13652,N_5717,N_6635);
and U13653 (N_13653,N_9485,N_7319);
xor U13654 (N_13654,N_6882,N_6839);
nor U13655 (N_13655,N_9151,N_6489);
nor U13656 (N_13656,N_6474,N_9206);
nor U13657 (N_13657,N_6799,N_6532);
xnor U13658 (N_13658,N_9838,N_7419);
xor U13659 (N_13659,N_8945,N_5274);
and U13660 (N_13660,N_7084,N_8139);
or U13661 (N_13661,N_6212,N_8835);
nand U13662 (N_13662,N_9631,N_9807);
nor U13663 (N_13663,N_8647,N_5797);
nand U13664 (N_13664,N_6368,N_5067);
nor U13665 (N_13665,N_7398,N_7713);
xnor U13666 (N_13666,N_9864,N_7152);
nor U13667 (N_13667,N_8253,N_5591);
xnor U13668 (N_13668,N_9191,N_7963);
and U13669 (N_13669,N_5230,N_7027);
and U13670 (N_13670,N_6703,N_8534);
xnor U13671 (N_13671,N_5234,N_8213);
nor U13672 (N_13672,N_7264,N_8237);
nor U13673 (N_13673,N_9559,N_5287);
or U13674 (N_13674,N_9151,N_9660);
nand U13675 (N_13675,N_7747,N_7399);
and U13676 (N_13676,N_7545,N_7490);
nand U13677 (N_13677,N_7915,N_8723);
and U13678 (N_13678,N_9892,N_8033);
nor U13679 (N_13679,N_8898,N_6772);
and U13680 (N_13680,N_9450,N_9293);
nand U13681 (N_13681,N_7103,N_8380);
and U13682 (N_13682,N_9034,N_7568);
and U13683 (N_13683,N_7654,N_8601);
nor U13684 (N_13684,N_6749,N_9221);
nand U13685 (N_13685,N_5169,N_9511);
nand U13686 (N_13686,N_9825,N_6671);
nor U13687 (N_13687,N_8299,N_8645);
nor U13688 (N_13688,N_8764,N_5193);
xnor U13689 (N_13689,N_7612,N_8852);
or U13690 (N_13690,N_5006,N_5846);
xor U13691 (N_13691,N_8919,N_9150);
nand U13692 (N_13692,N_5476,N_5576);
and U13693 (N_13693,N_8516,N_5789);
or U13694 (N_13694,N_9747,N_7960);
nand U13695 (N_13695,N_8463,N_7629);
nand U13696 (N_13696,N_8270,N_8334);
nor U13697 (N_13697,N_5604,N_5386);
xnor U13698 (N_13698,N_7707,N_6117);
nand U13699 (N_13699,N_9730,N_5865);
or U13700 (N_13700,N_7208,N_5408);
nand U13701 (N_13701,N_5806,N_8192);
nor U13702 (N_13702,N_5111,N_9137);
nor U13703 (N_13703,N_8455,N_9859);
and U13704 (N_13704,N_7063,N_9903);
and U13705 (N_13705,N_6321,N_9353);
nor U13706 (N_13706,N_6690,N_8655);
or U13707 (N_13707,N_5945,N_6935);
or U13708 (N_13708,N_9223,N_5138);
xnor U13709 (N_13709,N_6336,N_8261);
or U13710 (N_13710,N_7111,N_6231);
or U13711 (N_13711,N_6636,N_9664);
and U13712 (N_13712,N_6923,N_5257);
nand U13713 (N_13713,N_6084,N_5149);
xnor U13714 (N_13714,N_5724,N_6070);
nand U13715 (N_13715,N_5244,N_5566);
or U13716 (N_13716,N_7269,N_8011);
xor U13717 (N_13717,N_6421,N_8561);
nor U13718 (N_13718,N_8253,N_7759);
or U13719 (N_13719,N_7649,N_8049);
or U13720 (N_13720,N_9839,N_5465);
nor U13721 (N_13721,N_6494,N_9883);
nand U13722 (N_13722,N_9481,N_7233);
and U13723 (N_13723,N_5705,N_9153);
xnor U13724 (N_13724,N_6448,N_9319);
nor U13725 (N_13725,N_8612,N_9266);
nor U13726 (N_13726,N_7314,N_7838);
xor U13727 (N_13727,N_9024,N_7241);
xor U13728 (N_13728,N_7491,N_7440);
or U13729 (N_13729,N_6398,N_9682);
nand U13730 (N_13730,N_8124,N_7929);
nor U13731 (N_13731,N_5751,N_7466);
and U13732 (N_13732,N_9677,N_7330);
nor U13733 (N_13733,N_5712,N_9929);
xor U13734 (N_13734,N_5668,N_5136);
xor U13735 (N_13735,N_8236,N_9588);
and U13736 (N_13736,N_7366,N_6252);
or U13737 (N_13737,N_7513,N_8756);
or U13738 (N_13738,N_9929,N_9787);
xnor U13739 (N_13739,N_8263,N_5969);
and U13740 (N_13740,N_8179,N_6823);
and U13741 (N_13741,N_9422,N_7695);
nand U13742 (N_13742,N_5064,N_9136);
xor U13743 (N_13743,N_6890,N_5512);
xor U13744 (N_13744,N_9015,N_6058);
xnor U13745 (N_13745,N_5984,N_8009);
and U13746 (N_13746,N_6773,N_6946);
xnor U13747 (N_13747,N_7804,N_7745);
nor U13748 (N_13748,N_6899,N_7604);
nor U13749 (N_13749,N_9884,N_6916);
xor U13750 (N_13750,N_8178,N_7017);
or U13751 (N_13751,N_7837,N_5319);
nor U13752 (N_13752,N_8931,N_6411);
xnor U13753 (N_13753,N_7824,N_8967);
or U13754 (N_13754,N_6499,N_8101);
xnor U13755 (N_13755,N_7462,N_6717);
nand U13756 (N_13756,N_5974,N_5131);
nand U13757 (N_13757,N_6153,N_6447);
xor U13758 (N_13758,N_9813,N_5311);
or U13759 (N_13759,N_9550,N_6070);
or U13760 (N_13760,N_6314,N_5776);
and U13761 (N_13761,N_7243,N_5535);
or U13762 (N_13762,N_9656,N_7103);
nand U13763 (N_13763,N_9286,N_6078);
xor U13764 (N_13764,N_9835,N_8917);
nand U13765 (N_13765,N_6875,N_7406);
and U13766 (N_13766,N_9697,N_6798);
xor U13767 (N_13767,N_7368,N_7800);
or U13768 (N_13768,N_5528,N_8899);
xnor U13769 (N_13769,N_8047,N_9209);
nand U13770 (N_13770,N_9501,N_6349);
nor U13771 (N_13771,N_5882,N_9751);
and U13772 (N_13772,N_9892,N_5967);
or U13773 (N_13773,N_6665,N_6874);
or U13774 (N_13774,N_7852,N_5675);
xnor U13775 (N_13775,N_9368,N_5706);
xnor U13776 (N_13776,N_9298,N_7331);
or U13777 (N_13777,N_8362,N_7321);
nand U13778 (N_13778,N_9675,N_9534);
or U13779 (N_13779,N_6595,N_7566);
nand U13780 (N_13780,N_7760,N_6246);
and U13781 (N_13781,N_7884,N_6361);
and U13782 (N_13782,N_8759,N_7344);
nand U13783 (N_13783,N_6798,N_7238);
and U13784 (N_13784,N_6699,N_9858);
xnor U13785 (N_13785,N_7745,N_5220);
xor U13786 (N_13786,N_5504,N_7005);
nand U13787 (N_13787,N_6467,N_9625);
nor U13788 (N_13788,N_9005,N_8587);
nor U13789 (N_13789,N_7940,N_9230);
and U13790 (N_13790,N_8608,N_7503);
and U13791 (N_13791,N_5441,N_8562);
nor U13792 (N_13792,N_9487,N_5968);
and U13793 (N_13793,N_8840,N_5270);
nand U13794 (N_13794,N_6118,N_9828);
or U13795 (N_13795,N_8781,N_8405);
nor U13796 (N_13796,N_7772,N_6684);
xnor U13797 (N_13797,N_9238,N_6085);
or U13798 (N_13798,N_9983,N_7499);
nand U13799 (N_13799,N_5912,N_5652);
or U13800 (N_13800,N_6159,N_5603);
or U13801 (N_13801,N_5583,N_6142);
or U13802 (N_13802,N_6366,N_6590);
xor U13803 (N_13803,N_9987,N_5074);
nor U13804 (N_13804,N_5276,N_8956);
nor U13805 (N_13805,N_6253,N_6458);
or U13806 (N_13806,N_7405,N_7928);
or U13807 (N_13807,N_9501,N_8493);
and U13808 (N_13808,N_6708,N_8622);
xor U13809 (N_13809,N_8281,N_9830);
nand U13810 (N_13810,N_9716,N_8535);
or U13811 (N_13811,N_9423,N_5063);
xnor U13812 (N_13812,N_8682,N_9583);
or U13813 (N_13813,N_8587,N_7439);
nor U13814 (N_13814,N_9202,N_8065);
and U13815 (N_13815,N_9494,N_6720);
nor U13816 (N_13816,N_5559,N_7156);
nor U13817 (N_13817,N_5066,N_8987);
nand U13818 (N_13818,N_6986,N_5076);
or U13819 (N_13819,N_5147,N_5574);
xnor U13820 (N_13820,N_8806,N_8062);
xor U13821 (N_13821,N_9755,N_9472);
nor U13822 (N_13822,N_9508,N_6828);
or U13823 (N_13823,N_6737,N_9076);
and U13824 (N_13824,N_7966,N_5745);
and U13825 (N_13825,N_7703,N_9030);
nor U13826 (N_13826,N_9923,N_6408);
xor U13827 (N_13827,N_7408,N_7223);
and U13828 (N_13828,N_9610,N_8283);
nor U13829 (N_13829,N_9778,N_9891);
or U13830 (N_13830,N_7322,N_6840);
xor U13831 (N_13831,N_7620,N_9124);
nand U13832 (N_13832,N_6610,N_5421);
xor U13833 (N_13833,N_5319,N_5750);
or U13834 (N_13834,N_6014,N_6393);
or U13835 (N_13835,N_9923,N_6229);
xor U13836 (N_13836,N_7241,N_5057);
or U13837 (N_13837,N_5573,N_9018);
nor U13838 (N_13838,N_9810,N_8287);
nand U13839 (N_13839,N_6054,N_6125);
or U13840 (N_13840,N_7036,N_8207);
or U13841 (N_13841,N_7654,N_5818);
nor U13842 (N_13842,N_8683,N_7657);
nand U13843 (N_13843,N_7894,N_9220);
nand U13844 (N_13844,N_5111,N_9544);
nor U13845 (N_13845,N_6530,N_6986);
nand U13846 (N_13846,N_9720,N_6268);
xnor U13847 (N_13847,N_9230,N_6735);
and U13848 (N_13848,N_5906,N_8548);
nor U13849 (N_13849,N_7457,N_8349);
or U13850 (N_13850,N_6405,N_7267);
nor U13851 (N_13851,N_6860,N_5170);
nor U13852 (N_13852,N_9134,N_5528);
nand U13853 (N_13853,N_5989,N_5899);
or U13854 (N_13854,N_7822,N_5686);
nand U13855 (N_13855,N_6596,N_8403);
and U13856 (N_13856,N_6334,N_7237);
or U13857 (N_13857,N_6919,N_6365);
nor U13858 (N_13858,N_5311,N_6811);
xnor U13859 (N_13859,N_7533,N_7976);
and U13860 (N_13860,N_5984,N_5147);
or U13861 (N_13861,N_6690,N_6828);
nand U13862 (N_13862,N_6938,N_6817);
xnor U13863 (N_13863,N_8225,N_6676);
nor U13864 (N_13864,N_6422,N_8723);
xnor U13865 (N_13865,N_5787,N_6722);
and U13866 (N_13866,N_6017,N_9230);
or U13867 (N_13867,N_6338,N_6641);
nand U13868 (N_13868,N_8403,N_6561);
or U13869 (N_13869,N_7252,N_5468);
xnor U13870 (N_13870,N_6434,N_5164);
nor U13871 (N_13871,N_6627,N_5458);
nand U13872 (N_13872,N_9926,N_9788);
or U13873 (N_13873,N_7967,N_5407);
and U13874 (N_13874,N_8369,N_7552);
and U13875 (N_13875,N_8901,N_8323);
nand U13876 (N_13876,N_5817,N_8521);
xnor U13877 (N_13877,N_7249,N_8518);
nor U13878 (N_13878,N_9421,N_8846);
and U13879 (N_13879,N_9403,N_6932);
or U13880 (N_13880,N_6240,N_8649);
and U13881 (N_13881,N_9067,N_8282);
nand U13882 (N_13882,N_9942,N_8106);
and U13883 (N_13883,N_5542,N_8086);
nand U13884 (N_13884,N_5773,N_6231);
xor U13885 (N_13885,N_8393,N_6674);
and U13886 (N_13886,N_9011,N_8394);
nand U13887 (N_13887,N_9342,N_9926);
nand U13888 (N_13888,N_8603,N_6478);
and U13889 (N_13889,N_5191,N_5059);
nor U13890 (N_13890,N_7654,N_7497);
and U13891 (N_13891,N_6918,N_5851);
nand U13892 (N_13892,N_9918,N_9810);
nand U13893 (N_13893,N_7098,N_5442);
or U13894 (N_13894,N_5403,N_8556);
xor U13895 (N_13895,N_9294,N_5272);
nor U13896 (N_13896,N_8909,N_7918);
or U13897 (N_13897,N_8867,N_8293);
or U13898 (N_13898,N_6991,N_6996);
nor U13899 (N_13899,N_9571,N_7586);
nor U13900 (N_13900,N_8571,N_6022);
nand U13901 (N_13901,N_6961,N_9014);
or U13902 (N_13902,N_6582,N_8508);
or U13903 (N_13903,N_9636,N_8246);
or U13904 (N_13904,N_5267,N_7210);
and U13905 (N_13905,N_7550,N_8470);
xor U13906 (N_13906,N_5074,N_7404);
nor U13907 (N_13907,N_7256,N_5382);
or U13908 (N_13908,N_8112,N_7465);
or U13909 (N_13909,N_7143,N_8679);
or U13910 (N_13910,N_9414,N_7508);
or U13911 (N_13911,N_8400,N_9829);
or U13912 (N_13912,N_8871,N_9624);
and U13913 (N_13913,N_5978,N_8727);
nand U13914 (N_13914,N_6215,N_7948);
or U13915 (N_13915,N_9825,N_5310);
and U13916 (N_13916,N_7779,N_5213);
and U13917 (N_13917,N_8766,N_7161);
or U13918 (N_13918,N_8617,N_8728);
nor U13919 (N_13919,N_6113,N_8414);
and U13920 (N_13920,N_6779,N_9040);
and U13921 (N_13921,N_6030,N_8404);
xnor U13922 (N_13922,N_7242,N_8986);
nor U13923 (N_13923,N_5441,N_6091);
and U13924 (N_13924,N_6767,N_6207);
xor U13925 (N_13925,N_8034,N_6591);
nand U13926 (N_13926,N_9050,N_6593);
xor U13927 (N_13927,N_8685,N_6834);
nand U13928 (N_13928,N_9246,N_5488);
or U13929 (N_13929,N_8578,N_9718);
nor U13930 (N_13930,N_7142,N_5443);
and U13931 (N_13931,N_8085,N_8555);
nor U13932 (N_13932,N_7305,N_5961);
nand U13933 (N_13933,N_7861,N_9178);
nor U13934 (N_13934,N_8493,N_5215);
xor U13935 (N_13935,N_8176,N_8831);
nand U13936 (N_13936,N_6046,N_7547);
nor U13937 (N_13937,N_5447,N_7511);
or U13938 (N_13938,N_9258,N_5681);
nor U13939 (N_13939,N_8548,N_7649);
nand U13940 (N_13940,N_9927,N_7521);
xor U13941 (N_13941,N_5626,N_7245);
xnor U13942 (N_13942,N_8996,N_8637);
and U13943 (N_13943,N_7465,N_6317);
xnor U13944 (N_13944,N_5695,N_5117);
nor U13945 (N_13945,N_9360,N_5814);
and U13946 (N_13946,N_9932,N_6600);
or U13947 (N_13947,N_5780,N_5310);
or U13948 (N_13948,N_5794,N_9166);
xor U13949 (N_13949,N_5242,N_6486);
or U13950 (N_13950,N_8128,N_5041);
nand U13951 (N_13951,N_5731,N_9095);
and U13952 (N_13952,N_8624,N_8112);
and U13953 (N_13953,N_9060,N_6347);
nand U13954 (N_13954,N_9039,N_7595);
nor U13955 (N_13955,N_6340,N_5207);
nand U13956 (N_13956,N_7477,N_9284);
nand U13957 (N_13957,N_7374,N_8514);
and U13958 (N_13958,N_8308,N_6306);
and U13959 (N_13959,N_9764,N_9017);
xnor U13960 (N_13960,N_6457,N_5926);
nand U13961 (N_13961,N_6564,N_8504);
nand U13962 (N_13962,N_6805,N_6614);
or U13963 (N_13963,N_6730,N_5802);
xnor U13964 (N_13964,N_9465,N_5312);
or U13965 (N_13965,N_6160,N_6409);
and U13966 (N_13966,N_6662,N_7864);
nor U13967 (N_13967,N_8077,N_6321);
nor U13968 (N_13968,N_5204,N_8774);
xnor U13969 (N_13969,N_9416,N_5622);
nor U13970 (N_13970,N_9817,N_8632);
xor U13971 (N_13971,N_8713,N_5459);
and U13972 (N_13972,N_5123,N_6084);
nand U13973 (N_13973,N_9675,N_7851);
and U13974 (N_13974,N_6204,N_9165);
xor U13975 (N_13975,N_9071,N_8269);
nand U13976 (N_13976,N_8836,N_8680);
nor U13977 (N_13977,N_6548,N_6903);
xnor U13978 (N_13978,N_5118,N_9058);
nor U13979 (N_13979,N_8198,N_5745);
nor U13980 (N_13980,N_9562,N_6156);
nor U13981 (N_13981,N_7773,N_5003);
nand U13982 (N_13982,N_8001,N_6276);
or U13983 (N_13983,N_7990,N_9603);
nand U13984 (N_13984,N_7718,N_9665);
nand U13985 (N_13985,N_9571,N_8976);
and U13986 (N_13986,N_8890,N_7608);
and U13987 (N_13987,N_6950,N_9097);
or U13988 (N_13988,N_7331,N_5263);
nor U13989 (N_13989,N_6222,N_6646);
nor U13990 (N_13990,N_8230,N_9669);
nand U13991 (N_13991,N_8199,N_7202);
or U13992 (N_13992,N_8638,N_8692);
and U13993 (N_13993,N_8568,N_7801);
xor U13994 (N_13994,N_6072,N_7109);
or U13995 (N_13995,N_8170,N_8513);
and U13996 (N_13996,N_7223,N_9331);
nand U13997 (N_13997,N_5797,N_5882);
nor U13998 (N_13998,N_6815,N_6521);
nor U13999 (N_13999,N_9691,N_8874);
and U14000 (N_14000,N_9934,N_7203);
xnor U14001 (N_14001,N_6756,N_9719);
nand U14002 (N_14002,N_6818,N_8272);
xnor U14003 (N_14003,N_9192,N_8996);
or U14004 (N_14004,N_7070,N_8348);
nand U14005 (N_14005,N_5461,N_8820);
or U14006 (N_14006,N_8444,N_9079);
or U14007 (N_14007,N_6788,N_6713);
nand U14008 (N_14008,N_6766,N_6271);
nor U14009 (N_14009,N_5267,N_6385);
nand U14010 (N_14010,N_6409,N_5544);
and U14011 (N_14011,N_6391,N_8528);
and U14012 (N_14012,N_6302,N_9820);
xnor U14013 (N_14013,N_9865,N_5305);
xnor U14014 (N_14014,N_6688,N_7925);
or U14015 (N_14015,N_8110,N_7564);
or U14016 (N_14016,N_6372,N_5504);
nor U14017 (N_14017,N_5125,N_9445);
nor U14018 (N_14018,N_9203,N_9783);
or U14019 (N_14019,N_5993,N_5315);
xnor U14020 (N_14020,N_7428,N_7386);
nand U14021 (N_14021,N_6369,N_9766);
or U14022 (N_14022,N_5359,N_6857);
and U14023 (N_14023,N_8094,N_9548);
nor U14024 (N_14024,N_5437,N_6952);
and U14025 (N_14025,N_6330,N_5717);
and U14026 (N_14026,N_8320,N_6351);
nand U14027 (N_14027,N_6003,N_5033);
and U14028 (N_14028,N_6356,N_7415);
nand U14029 (N_14029,N_9886,N_8984);
xnor U14030 (N_14030,N_8023,N_5969);
and U14031 (N_14031,N_8513,N_7245);
nor U14032 (N_14032,N_6388,N_6608);
nor U14033 (N_14033,N_8717,N_5612);
xnor U14034 (N_14034,N_5945,N_6272);
xnor U14035 (N_14035,N_5383,N_7079);
nor U14036 (N_14036,N_5664,N_9332);
xor U14037 (N_14037,N_7094,N_5306);
xnor U14038 (N_14038,N_9288,N_5804);
xor U14039 (N_14039,N_6171,N_7247);
and U14040 (N_14040,N_6696,N_5454);
xnor U14041 (N_14041,N_7557,N_8195);
or U14042 (N_14042,N_8936,N_5478);
nor U14043 (N_14043,N_6018,N_8871);
or U14044 (N_14044,N_7929,N_6374);
and U14045 (N_14045,N_7215,N_6179);
xnor U14046 (N_14046,N_5849,N_5174);
and U14047 (N_14047,N_6727,N_9874);
nand U14048 (N_14048,N_7488,N_8286);
or U14049 (N_14049,N_5991,N_7365);
or U14050 (N_14050,N_6623,N_6865);
nand U14051 (N_14051,N_7479,N_8939);
nand U14052 (N_14052,N_9223,N_9878);
xor U14053 (N_14053,N_8068,N_6787);
or U14054 (N_14054,N_6806,N_8947);
nand U14055 (N_14055,N_7781,N_7006);
nand U14056 (N_14056,N_5198,N_8913);
or U14057 (N_14057,N_7565,N_9534);
nand U14058 (N_14058,N_8301,N_6084);
nor U14059 (N_14059,N_9999,N_5538);
or U14060 (N_14060,N_9942,N_7784);
nand U14061 (N_14061,N_8528,N_5579);
and U14062 (N_14062,N_6002,N_6486);
or U14063 (N_14063,N_9335,N_5571);
and U14064 (N_14064,N_6432,N_9142);
nand U14065 (N_14065,N_8147,N_5181);
nor U14066 (N_14066,N_6909,N_8913);
or U14067 (N_14067,N_6329,N_8320);
or U14068 (N_14068,N_9928,N_5038);
or U14069 (N_14069,N_5969,N_6192);
xor U14070 (N_14070,N_5163,N_6625);
or U14071 (N_14071,N_9078,N_8526);
xnor U14072 (N_14072,N_6529,N_7491);
nor U14073 (N_14073,N_9602,N_8238);
xor U14074 (N_14074,N_9292,N_8764);
nor U14075 (N_14075,N_8260,N_8786);
or U14076 (N_14076,N_5213,N_8468);
nor U14077 (N_14077,N_6180,N_5295);
or U14078 (N_14078,N_9317,N_8995);
nor U14079 (N_14079,N_6740,N_7164);
nand U14080 (N_14080,N_6348,N_8210);
nor U14081 (N_14081,N_6675,N_5293);
or U14082 (N_14082,N_7437,N_7970);
or U14083 (N_14083,N_5220,N_8028);
xnor U14084 (N_14084,N_8499,N_9194);
nor U14085 (N_14085,N_8489,N_6726);
nor U14086 (N_14086,N_8344,N_8275);
or U14087 (N_14087,N_6303,N_6719);
nor U14088 (N_14088,N_9953,N_9930);
xnor U14089 (N_14089,N_7233,N_9904);
xor U14090 (N_14090,N_8014,N_6248);
and U14091 (N_14091,N_6153,N_5437);
nor U14092 (N_14092,N_8331,N_6970);
nor U14093 (N_14093,N_6413,N_8983);
or U14094 (N_14094,N_9162,N_5755);
xnor U14095 (N_14095,N_5200,N_8852);
xnor U14096 (N_14096,N_7157,N_8050);
nand U14097 (N_14097,N_8400,N_9110);
nand U14098 (N_14098,N_6996,N_7971);
nor U14099 (N_14099,N_7451,N_8715);
or U14100 (N_14100,N_6011,N_9492);
xnor U14101 (N_14101,N_8695,N_5883);
xor U14102 (N_14102,N_7335,N_6513);
nand U14103 (N_14103,N_8046,N_9022);
or U14104 (N_14104,N_5988,N_7248);
xor U14105 (N_14105,N_8106,N_5609);
nand U14106 (N_14106,N_6571,N_5235);
and U14107 (N_14107,N_5198,N_8777);
xnor U14108 (N_14108,N_9773,N_7270);
and U14109 (N_14109,N_6218,N_7726);
nor U14110 (N_14110,N_9663,N_7870);
nor U14111 (N_14111,N_5741,N_8485);
xor U14112 (N_14112,N_9767,N_7893);
nand U14113 (N_14113,N_6694,N_6693);
nor U14114 (N_14114,N_7219,N_7988);
xor U14115 (N_14115,N_7681,N_6361);
xor U14116 (N_14116,N_9863,N_7503);
or U14117 (N_14117,N_9233,N_6519);
and U14118 (N_14118,N_5671,N_8503);
xor U14119 (N_14119,N_8427,N_5307);
nand U14120 (N_14120,N_7517,N_9164);
or U14121 (N_14121,N_7489,N_7938);
and U14122 (N_14122,N_6075,N_7221);
xor U14123 (N_14123,N_8623,N_9090);
nand U14124 (N_14124,N_8620,N_8946);
or U14125 (N_14125,N_9282,N_5183);
or U14126 (N_14126,N_6876,N_5374);
or U14127 (N_14127,N_8519,N_9959);
xor U14128 (N_14128,N_5818,N_8113);
and U14129 (N_14129,N_5208,N_9651);
or U14130 (N_14130,N_8038,N_8900);
nor U14131 (N_14131,N_9118,N_9293);
or U14132 (N_14132,N_7186,N_7441);
nand U14133 (N_14133,N_9801,N_6762);
nand U14134 (N_14134,N_9446,N_9247);
and U14135 (N_14135,N_8102,N_5787);
xnor U14136 (N_14136,N_5508,N_9512);
nand U14137 (N_14137,N_8507,N_5026);
nand U14138 (N_14138,N_8127,N_9426);
nand U14139 (N_14139,N_7242,N_5089);
xnor U14140 (N_14140,N_9183,N_8443);
xor U14141 (N_14141,N_9222,N_9388);
nand U14142 (N_14142,N_8408,N_6036);
or U14143 (N_14143,N_8858,N_9336);
nor U14144 (N_14144,N_9653,N_8192);
nand U14145 (N_14145,N_5032,N_6046);
or U14146 (N_14146,N_7558,N_6686);
and U14147 (N_14147,N_6781,N_7458);
xnor U14148 (N_14148,N_9140,N_5420);
xnor U14149 (N_14149,N_9315,N_8323);
nand U14150 (N_14150,N_7362,N_5060);
nor U14151 (N_14151,N_9829,N_5143);
nand U14152 (N_14152,N_6241,N_9392);
nor U14153 (N_14153,N_7240,N_9876);
nand U14154 (N_14154,N_5499,N_8811);
or U14155 (N_14155,N_7058,N_6229);
nor U14156 (N_14156,N_6042,N_7312);
nor U14157 (N_14157,N_7762,N_8924);
nor U14158 (N_14158,N_5384,N_8570);
nand U14159 (N_14159,N_6872,N_6661);
or U14160 (N_14160,N_9573,N_6950);
or U14161 (N_14161,N_8132,N_9464);
xnor U14162 (N_14162,N_6018,N_6410);
nand U14163 (N_14163,N_5989,N_7808);
and U14164 (N_14164,N_8291,N_7934);
nand U14165 (N_14165,N_6879,N_5448);
or U14166 (N_14166,N_8432,N_9547);
and U14167 (N_14167,N_9313,N_7225);
and U14168 (N_14168,N_6516,N_5912);
or U14169 (N_14169,N_6927,N_5462);
nor U14170 (N_14170,N_6366,N_7563);
nor U14171 (N_14171,N_6684,N_5292);
nand U14172 (N_14172,N_7706,N_6471);
and U14173 (N_14173,N_5344,N_9364);
nor U14174 (N_14174,N_7954,N_5114);
xnor U14175 (N_14175,N_5468,N_6152);
nand U14176 (N_14176,N_6095,N_5507);
xnor U14177 (N_14177,N_6043,N_6661);
nand U14178 (N_14178,N_8330,N_9170);
xnor U14179 (N_14179,N_5766,N_7504);
nor U14180 (N_14180,N_9628,N_8174);
and U14181 (N_14181,N_8596,N_8974);
or U14182 (N_14182,N_5382,N_6021);
xnor U14183 (N_14183,N_8514,N_8328);
nand U14184 (N_14184,N_7534,N_8195);
and U14185 (N_14185,N_5353,N_9829);
or U14186 (N_14186,N_9323,N_7032);
and U14187 (N_14187,N_8697,N_9834);
or U14188 (N_14188,N_9059,N_9549);
xor U14189 (N_14189,N_6484,N_9211);
or U14190 (N_14190,N_9713,N_6551);
or U14191 (N_14191,N_5338,N_8682);
nand U14192 (N_14192,N_6740,N_6108);
or U14193 (N_14193,N_8862,N_8918);
nand U14194 (N_14194,N_8175,N_5020);
nand U14195 (N_14195,N_5867,N_8731);
nand U14196 (N_14196,N_7333,N_5580);
and U14197 (N_14197,N_9006,N_7800);
or U14198 (N_14198,N_7245,N_9040);
or U14199 (N_14199,N_8510,N_7193);
or U14200 (N_14200,N_5229,N_5749);
nor U14201 (N_14201,N_7199,N_9675);
or U14202 (N_14202,N_7361,N_5311);
and U14203 (N_14203,N_8629,N_6531);
xor U14204 (N_14204,N_8806,N_6050);
and U14205 (N_14205,N_5251,N_7822);
nand U14206 (N_14206,N_8109,N_7880);
nand U14207 (N_14207,N_5095,N_9735);
xor U14208 (N_14208,N_8704,N_6419);
nand U14209 (N_14209,N_9446,N_9649);
nor U14210 (N_14210,N_8168,N_7599);
or U14211 (N_14211,N_8936,N_8240);
nand U14212 (N_14212,N_6466,N_6589);
nand U14213 (N_14213,N_6354,N_8829);
and U14214 (N_14214,N_6132,N_8421);
or U14215 (N_14215,N_9043,N_7235);
nor U14216 (N_14216,N_7556,N_8562);
nor U14217 (N_14217,N_6769,N_7924);
nor U14218 (N_14218,N_8149,N_9304);
nand U14219 (N_14219,N_5447,N_5655);
or U14220 (N_14220,N_6132,N_7631);
or U14221 (N_14221,N_9164,N_8563);
nand U14222 (N_14222,N_9106,N_8150);
and U14223 (N_14223,N_8657,N_9648);
xor U14224 (N_14224,N_7143,N_7360);
xnor U14225 (N_14225,N_9650,N_8247);
nor U14226 (N_14226,N_5551,N_9101);
or U14227 (N_14227,N_9253,N_8956);
nand U14228 (N_14228,N_9432,N_6744);
or U14229 (N_14229,N_7754,N_6616);
and U14230 (N_14230,N_8803,N_5045);
nand U14231 (N_14231,N_6049,N_8959);
or U14232 (N_14232,N_8412,N_9479);
and U14233 (N_14233,N_9743,N_9968);
or U14234 (N_14234,N_6817,N_8671);
or U14235 (N_14235,N_6444,N_7787);
nor U14236 (N_14236,N_7317,N_5877);
xnor U14237 (N_14237,N_8794,N_7883);
and U14238 (N_14238,N_5583,N_6084);
and U14239 (N_14239,N_6991,N_7475);
xnor U14240 (N_14240,N_8388,N_6080);
or U14241 (N_14241,N_6432,N_9591);
xor U14242 (N_14242,N_5975,N_6448);
nor U14243 (N_14243,N_6222,N_9621);
or U14244 (N_14244,N_7024,N_8960);
nand U14245 (N_14245,N_5789,N_6300);
or U14246 (N_14246,N_6686,N_9092);
and U14247 (N_14247,N_5958,N_6598);
xnor U14248 (N_14248,N_8872,N_5779);
nor U14249 (N_14249,N_7045,N_6566);
nor U14250 (N_14250,N_6536,N_8325);
or U14251 (N_14251,N_7178,N_8602);
xor U14252 (N_14252,N_5731,N_6987);
nand U14253 (N_14253,N_5463,N_7268);
xor U14254 (N_14254,N_6420,N_8185);
nand U14255 (N_14255,N_6427,N_9104);
or U14256 (N_14256,N_6011,N_8300);
xor U14257 (N_14257,N_7663,N_9014);
xnor U14258 (N_14258,N_8547,N_8091);
nand U14259 (N_14259,N_8763,N_9667);
xor U14260 (N_14260,N_8516,N_5540);
or U14261 (N_14261,N_5610,N_5057);
nand U14262 (N_14262,N_9882,N_8487);
nand U14263 (N_14263,N_7766,N_5132);
and U14264 (N_14264,N_9229,N_7781);
xnor U14265 (N_14265,N_9280,N_6413);
xor U14266 (N_14266,N_9182,N_5428);
nand U14267 (N_14267,N_9101,N_7414);
nand U14268 (N_14268,N_8612,N_5191);
and U14269 (N_14269,N_8016,N_9636);
and U14270 (N_14270,N_7040,N_5961);
or U14271 (N_14271,N_7422,N_7791);
and U14272 (N_14272,N_8100,N_7968);
xnor U14273 (N_14273,N_7061,N_6329);
or U14274 (N_14274,N_6201,N_7969);
and U14275 (N_14275,N_7544,N_8935);
xnor U14276 (N_14276,N_8735,N_5133);
xnor U14277 (N_14277,N_7141,N_7203);
nand U14278 (N_14278,N_9211,N_8375);
nor U14279 (N_14279,N_5923,N_9438);
nor U14280 (N_14280,N_6052,N_7851);
or U14281 (N_14281,N_5743,N_7159);
nand U14282 (N_14282,N_5012,N_6649);
nor U14283 (N_14283,N_8938,N_5973);
nor U14284 (N_14284,N_9576,N_6060);
nand U14285 (N_14285,N_6370,N_9115);
xnor U14286 (N_14286,N_7752,N_8882);
or U14287 (N_14287,N_9210,N_8244);
and U14288 (N_14288,N_5922,N_9870);
nor U14289 (N_14289,N_7958,N_5306);
and U14290 (N_14290,N_5084,N_7801);
nor U14291 (N_14291,N_6842,N_9631);
and U14292 (N_14292,N_9423,N_9290);
xor U14293 (N_14293,N_5714,N_6752);
nand U14294 (N_14294,N_5376,N_5692);
xnor U14295 (N_14295,N_5688,N_7373);
nor U14296 (N_14296,N_9283,N_8954);
nor U14297 (N_14297,N_6715,N_7832);
nand U14298 (N_14298,N_6744,N_5521);
or U14299 (N_14299,N_9990,N_5424);
nand U14300 (N_14300,N_7921,N_9772);
or U14301 (N_14301,N_5403,N_6403);
nand U14302 (N_14302,N_6541,N_6488);
or U14303 (N_14303,N_6883,N_8612);
nor U14304 (N_14304,N_9864,N_7517);
nor U14305 (N_14305,N_6263,N_9919);
xnor U14306 (N_14306,N_8823,N_6659);
or U14307 (N_14307,N_9197,N_5292);
or U14308 (N_14308,N_8750,N_8450);
or U14309 (N_14309,N_8630,N_9788);
nor U14310 (N_14310,N_8169,N_9141);
or U14311 (N_14311,N_6090,N_9783);
or U14312 (N_14312,N_8219,N_9567);
nand U14313 (N_14313,N_5106,N_6091);
and U14314 (N_14314,N_5700,N_5355);
xnor U14315 (N_14315,N_7713,N_5558);
xnor U14316 (N_14316,N_5616,N_7173);
xnor U14317 (N_14317,N_8733,N_5727);
nand U14318 (N_14318,N_7889,N_9369);
xnor U14319 (N_14319,N_6978,N_9878);
and U14320 (N_14320,N_7277,N_9700);
or U14321 (N_14321,N_7994,N_6736);
nor U14322 (N_14322,N_6711,N_7186);
nor U14323 (N_14323,N_9322,N_8880);
or U14324 (N_14324,N_9414,N_8212);
or U14325 (N_14325,N_8683,N_5706);
and U14326 (N_14326,N_9200,N_7262);
nor U14327 (N_14327,N_8294,N_6599);
nor U14328 (N_14328,N_8320,N_8515);
nor U14329 (N_14329,N_9143,N_6789);
xor U14330 (N_14330,N_7516,N_5808);
and U14331 (N_14331,N_9589,N_7494);
or U14332 (N_14332,N_9029,N_8179);
xnor U14333 (N_14333,N_8927,N_8897);
nor U14334 (N_14334,N_9377,N_5148);
or U14335 (N_14335,N_9994,N_9270);
nor U14336 (N_14336,N_6278,N_9076);
or U14337 (N_14337,N_8268,N_8919);
nand U14338 (N_14338,N_9776,N_7243);
nand U14339 (N_14339,N_8519,N_5289);
or U14340 (N_14340,N_7336,N_6522);
nor U14341 (N_14341,N_8986,N_6656);
or U14342 (N_14342,N_5053,N_5325);
or U14343 (N_14343,N_8402,N_6979);
nor U14344 (N_14344,N_5261,N_9657);
nor U14345 (N_14345,N_7409,N_6184);
nand U14346 (N_14346,N_9231,N_6969);
or U14347 (N_14347,N_6552,N_8952);
xor U14348 (N_14348,N_6755,N_9213);
or U14349 (N_14349,N_5320,N_6747);
and U14350 (N_14350,N_9146,N_8890);
and U14351 (N_14351,N_7706,N_7564);
nor U14352 (N_14352,N_8438,N_9477);
nand U14353 (N_14353,N_6656,N_8157);
xor U14354 (N_14354,N_6653,N_7835);
or U14355 (N_14355,N_7905,N_9176);
nor U14356 (N_14356,N_7481,N_7747);
xor U14357 (N_14357,N_5208,N_8802);
nor U14358 (N_14358,N_6351,N_8682);
xor U14359 (N_14359,N_9421,N_8624);
and U14360 (N_14360,N_8790,N_6905);
nand U14361 (N_14361,N_8577,N_9679);
xor U14362 (N_14362,N_6107,N_5048);
nor U14363 (N_14363,N_6843,N_8035);
nor U14364 (N_14364,N_8444,N_9694);
nand U14365 (N_14365,N_8587,N_7941);
nand U14366 (N_14366,N_9913,N_6415);
and U14367 (N_14367,N_6839,N_5684);
or U14368 (N_14368,N_9105,N_5174);
or U14369 (N_14369,N_6155,N_7751);
and U14370 (N_14370,N_9786,N_8049);
xnor U14371 (N_14371,N_8725,N_6786);
and U14372 (N_14372,N_8168,N_8259);
or U14373 (N_14373,N_5280,N_9636);
and U14374 (N_14374,N_8105,N_9624);
and U14375 (N_14375,N_8716,N_5434);
or U14376 (N_14376,N_9008,N_7593);
nand U14377 (N_14377,N_7522,N_5795);
nor U14378 (N_14378,N_5197,N_9203);
nand U14379 (N_14379,N_7187,N_9084);
nand U14380 (N_14380,N_9043,N_6965);
or U14381 (N_14381,N_9305,N_7362);
nand U14382 (N_14382,N_9063,N_5774);
nand U14383 (N_14383,N_9939,N_7474);
and U14384 (N_14384,N_5747,N_7854);
or U14385 (N_14385,N_6309,N_9315);
nand U14386 (N_14386,N_8246,N_7371);
nand U14387 (N_14387,N_7039,N_9319);
or U14388 (N_14388,N_5652,N_7067);
nor U14389 (N_14389,N_6197,N_9864);
or U14390 (N_14390,N_9713,N_8438);
xnor U14391 (N_14391,N_9819,N_5411);
nand U14392 (N_14392,N_8915,N_8008);
nor U14393 (N_14393,N_7182,N_9306);
nand U14394 (N_14394,N_9471,N_5485);
and U14395 (N_14395,N_6010,N_8821);
and U14396 (N_14396,N_8428,N_8923);
and U14397 (N_14397,N_9789,N_6834);
nand U14398 (N_14398,N_7269,N_7273);
xor U14399 (N_14399,N_6339,N_8758);
and U14400 (N_14400,N_9985,N_5413);
or U14401 (N_14401,N_9920,N_9075);
nor U14402 (N_14402,N_6186,N_9286);
and U14403 (N_14403,N_9204,N_9882);
nor U14404 (N_14404,N_8892,N_5162);
and U14405 (N_14405,N_5341,N_5687);
and U14406 (N_14406,N_9942,N_8541);
nand U14407 (N_14407,N_9734,N_5198);
xnor U14408 (N_14408,N_9055,N_9460);
nand U14409 (N_14409,N_6772,N_5350);
or U14410 (N_14410,N_6970,N_6954);
nor U14411 (N_14411,N_9675,N_6110);
and U14412 (N_14412,N_7953,N_9379);
nand U14413 (N_14413,N_7674,N_8974);
and U14414 (N_14414,N_6280,N_6931);
nor U14415 (N_14415,N_6763,N_5052);
and U14416 (N_14416,N_8199,N_8555);
xor U14417 (N_14417,N_5354,N_6628);
or U14418 (N_14418,N_6661,N_8704);
nand U14419 (N_14419,N_5826,N_9412);
and U14420 (N_14420,N_6178,N_6403);
or U14421 (N_14421,N_9168,N_7271);
nor U14422 (N_14422,N_9291,N_9144);
xor U14423 (N_14423,N_5777,N_9245);
xnor U14424 (N_14424,N_5401,N_7783);
xnor U14425 (N_14425,N_7295,N_9665);
nor U14426 (N_14426,N_9436,N_5809);
nor U14427 (N_14427,N_7751,N_5873);
xor U14428 (N_14428,N_8219,N_5040);
nand U14429 (N_14429,N_6975,N_5071);
and U14430 (N_14430,N_7389,N_8602);
nand U14431 (N_14431,N_6141,N_8531);
and U14432 (N_14432,N_6200,N_8534);
nand U14433 (N_14433,N_9299,N_7654);
or U14434 (N_14434,N_5166,N_7519);
nor U14435 (N_14435,N_7540,N_7184);
nor U14436 (N_14436,N_7549,N_9643);
or U14437 (N_14437,N_6051,N_6032);
and U14438 (N_14438,N_9668,N_8275);
and U14439 (N_14439,N_5504,N_8948);
and U14440 (N_14440,N_5654,N_5652);
nor U14441 (N_14441,N_5628,N_6034);
and U14442 (N_14442,N_5855,N_8755);
xor U14443 (N_14443,N_5579,N_8870);
xnor U14444 (N_14444,N_7098,N_8230);
nor U14445 (N_14445,N_8595,N_9577);
xnor U14446 (N_14446,N_7692,N_6179);
and U14447 (N_14447,N_9624,N_6657);
or U14448 (N_14448,N_5464,N_6274);
or U14449 (N_14449,N_7774,N_7952);
nor U14450 (N_14450,N_9625,N_9627);
nor U14451 (N_14451,N_7550,N_8816);
nor U14452 (N_14452,N_6481,N_5790);
nand U14453 (N_14453,N_7739,N_9130);
xor U14454 (N_14454,N_6486,N_8472);
nor U14455 (N_14455,N_6389,N_9729);
or U14456 (N_14456,N_7141,N_7300);
xnor U14457 (N_14457,N_7330,N_6152);
nand U14458 (N_14458,N_7131,N_9732);
and U14459 (N_14459,N_9830,N_5482);
nor U14460 (N_14460,N_5163,N_7691);
xor U14461 (N_14461,N_5108,N_5409);
or U14462 (N_14462,N_9188,N_7103);
xor U14463 (N_14463,N_5962,N_6677);
or U14464 (N_14464,N_5339,N_8937);
nor U14465 (N_14465,N_5733,N_9959);
and U14466 (N_14466,N_9324,N_9841);
or U14467 (N_14467,N_9840,N_9639);
nand U14468 (N_14468,N_5351,N_9703);
and U14469 (N_14469,N_5906,N_9656);
nand U14470 (N_14470,N_5110,N_9746);
and U14471 (N_14471,N_5809,N_9935);
nand U14472 (N_14472,N_8048,N_6918);
or U14473 (N_14473,N_9083,N_7903);
nand U14474 (N_14474,N_8397,N_5660);
nor U14475 (N_14475,N_6464,N_9777);
nor U14476 (N_14476,N_8728,N_7123);
nand U14477 (N_14477,N_6480,N_8654);
nand U14478 (N_14478,N_7905,N_6488);
or U14479 (N_14479,N_9468,N_5639);
nand U14480 (N_14480,N_7289,N_9647);
or U14481 (N_14481,N_7096,N_8023);
xnor U14482 (N_14482,N_8966,N_9956);
xor U14483 (N_14483,N_6322,N_9079);
nand U14484 (N_14484,N_7747,N_5811);
nor U14485 (N_14485,N_7067,N_9827);
xnor U14486 (N_14486,N_5286,N_6888);
nor U14487 (N_14487,N_7781,N_8660);
nand U14488 (N_14488,N_5860,N_8544);
or U14489 (N_14489,N_9175,N_8868);
or U14490 (N_14490,N_7765,N_8898);
or U14491 (N_14491,N_9037,N_7066);
nand U14492 (N_14492,N_7721,N_6098);
nor U14493 (N_14493,N_6403,N_6823);
nor U14494 (N_14494,N_8909,N_8461);
xnor U14495 (N_14495,N_5926,N_5332);
nor U14496 (N_14496,N_5992,N_8990);
or U14497 (N_14497,N_8423,N_8464);
or U14498 (N_14498,N_6710,N_9130);
nand U14499 (N_14499,N_7562,N_9826);
or U14500 (N_14500,N_9950,N_5114);
and U14501 (N_14501,N_9496,N_8276);
or U14502 (N_14502,N_6571,N_7599);
nor U14503 (N_14503,N_6284,N_5370);
and U14504 (N_14504,N_8237,N_9569);
or U14505 (N_14505,N_9676,N_5249);
and U14506 (N_14506,N_7877,N_5189);
or U14507 (N_14507,N_8850,N_9300);
nand U14508 (N_14508,N_5560,N_8130);
or U14509 (N_14509,N_5905,N_7485);
xnor U14510 (N_14510,N_9187,N_6193);
or U14511 (N_14511,N_6854,N_8067);
and U14512 (N_14512,N_9389,N_5071);
nand U14513 (N_14513,N_6316,N_8046);
or U14514 (N_14514,N_7630,N_7925);
or U14515 (N_14515,N_8073,N_9945);
or U14516 (N_14516,N_9422,N_9990);
xor U14517 (N_14517,N_7542,N_6461);
nor U14518 (N_14518,N_5866,N_7627);
and U14519 (N_14519,N_5294,N_5111);
and U14520 (N_14520,N_7269,N_8740);
and U14521 (N_14521,N_6933,N_9234);
xor U14522 (N_14522,N_6250,N_9715);
or U14523 (N_14523,N_7597,N_5044);
and U14524 (N_14524,N_8622,N_9890);
and U14525 (N_14525,N_5870,N_8336);
nand U14526 (N_14526,N_8836,N_5290);
nor U14527 (N_14527,N_7917,N_8508);
xnor U14528 (N_14528,N_8446,N_5116);
or U14529 (N_14529,N_6779,N_9429);
nand U14530 (N_14530,N_8467,N_5776);
xor U14531 (N_14531,N_6633,N_7819);
nand U14532 (N_14532,N_7141,N_8220);
xnor U14533 (N_14533,N_5521,N_8837);
nand U14534 (N_14534,N_5054,N_6553);
xor U14535 (N_14535,N_7268,N_5744);
nand U14536 (N_14536,N_9517,N_7407);
nand U14537 (N_14537,N_7186,N_7957);
nand U14538 (N_14538,N_6300,N_9003);
nand U14539 (N_14539,N_8941,N_8652);
nor U14540 (N_14540,N_9299,N_5693);
nor U14541 (N_14541,N_6747,N_5029);
nor U14542 (N_14542,N_6603,N_5938);
xnor U14543 (N_14543,N_6134,N_8660);
nor U14544 (N_14544,N_7405,N_6592);
and U14545 (N_14545,N_6821,N_9022);
xnor U14546 (N_14546,N_5790,N_6085);
and U14547 (N_14547,N_8586,N_9286);
nand U14548 (N_14548,N_8277,N_5694);
nor U14549 (N_14549,N_6408,N_9111);
or U14550 (N_14550,N_9215,N_6103);
xor U14551 (N_14551,N_5582,N_9217);
or U14552 (N_14552,N_9409,N_8706);
xor U14553 (N_14553,N_6469,N_9448);
or U14554 (N_14554,N_9284,N_6625);
and U14555 (N_14555,N_6781,N_5366);
nor U14556 (N_14556,N_7308,N_8368);
and U14557 (N_14557,N_8968,N_6602);
nand U14558 (N_14558,N_5565,N_8106);
nor U14559 (N_14559,N_8813,N_5053);
or U14560 (N_14560,N_8328,N_9667);
xnor U14561 (N_14561,N_7413,N_8348);
or U14562 (N_14562,N_6624,N_9630);
xnor U14563 (N_14563,N_7546,N_6436);
nand U14564 (N_14564,N_7250,N_9971);
nand U14565 (N_14565,N_8099,N_9259);
or U14566 (N_14566,N_9346,N_9610);
xnor U14567 (N_14567,N_9511,N_5977);
nand U14568 (N_14568,N_6729,N_7269);
nand U14569 (N_14569,N_7559,N_8894);
and U14570 (N_14570,N_5600,N_8636);
and U14571 (N_14571,N_8484,N_5520);
xor U14572 (N_14572,N_7989,N_9591);
xnor U14573 (N_14573,N_5987,N_5704);
nor U14574 (N_14574,N_5369,N_5573);
nor U14575 (N_14575,N_7466,N_7552);
nand U14576 (N_14576,N_9377,N_7500);
nor U14577 (N_14577,N_7766,N_7573);
xor U14578 (N_14578,N_8004,N_8382);
or U14579 (N_14579,N_9833,N_9035);
nand U14580 (N_14580,N_7073,N_6489);
xnor U14581 (N_14581,N_9884,N_8108);
nand U14582 (N_14582,N_5773,N_5462);
and U14583 (N_14583,N_6086,N_9897);
nor U14584 (N_14584,N_8693,N_9455);
nor U14585 (N_14585,N_6351,N_9400);
and U14586 (N_14586,N_9014,N_8192);
nand U14587 (N_14587,N_9106,N_8493);
xor U14588 (N_14588,N_9311,N_8822);
nand U14589 (N_14589,N_5184,N_6625);
nor U14590 (N_14590,N_6342,N_7677);
nor U14591 (N_14591,N_9762,N_6351);
nor U14592 (N_14592,N_6520,N_8551);
nand U14593 (N_14593,N_7417,N_8830);
or U14594 (N_14594,N_5288,N_5598);
nor U14595 (N_14595,N_5592,N_8761);
or U14596 (N_14596,N_6508,N_7885);
and U14597 (N_14597,N_9324,N_9620);
or U14598 (N_14598,N_7606,N_6722);
nand U14599 (N_14599,N_7990,N_7985);
xor U14600 (N_14600,N_7524,N_9144);
nor U14601 (N_14601,N_6526,N_6628);
and U14602 (N_14602,N_8009,N_6010);
nand U14603 (N_14603,N_5542,N_8938);
or U14604 (N_14604,N_6715,N_7831);
or U14605 (N_14605,N_9489,N_9514);
and U14606 (N_14606,N_5882,N_8644);
nor U14607 (N_14607,N_5890,N_9462);
xor U14608 (N_14608,N_9147,N_8924);
or U14609 (N_14609,N_9569,N_9534);
or U14610 (N_14610,N_7929,N_8017);
xor U14611 (N_14611,N_7654,N_7877);
xnor U14612 (N_14612,N_6304,N_6138);
xor U14613 (N_14613,N_5143,N_7999);
nor U14614 (N_14614,N_6635,N_9693);
nand U14615 (N_14615,N_5221,N_5093);
and U14616 (N_14616,N_6851,N_9515);
xnor U14617 (N_14617,N_8285,N_8782);
nor U14618 (N_14618,N_7528,N_5183);
nand U14619 (N_14619,N_6868,N_7038);
or U14620 (N_14620,N_9647,N_5626);
nand U14621 (N_14621,N_8492,N_5218);
and U14622 (N_14622,N_5614,N_6822);
nand U14623 (N_14623,N_9249,N_7808);
nor U14624 (N_14624,N_9864,N_9005);
and U14625 (N_14625,N_6827,N_7428);
and U14626 (N_14626,N_9921,N_6439);
nand U14627 (N_14627,N_5240,N_6651);
xor U14628 (N_14628,N_7272,N_5643);
nand U14629 (N_14629,N_6647,N_9644);
nand U14630 (N_14630,N_5257,N_5906);
or U14631 (N_14631,N_9697,N_7031);
and U14632 (N_14632,N_5119,N_8004);
or U14633 (N_14633,N_5074,N_6211);
nand U14634 (N_14634,N_6149,N_6275);
or U14635 (N_14635,N_6377,N_7645);
and U14636 (N_14636,N_8026,N_9913);
or U14637 (N_14637,N_8590,N_8634);
nand U14638 (N_14638,N_9942,N_5179);
xnor U14639 (N_14639,N_9559,N_9023);
nor U14640 (N_14640,N_5837,N_6613);
nand U14641 (N_14641,N_9523,N_9110);
nand U14642 (N_14642,N_9884,N_8558);
xor U14643 (N_14643,N_5285,N_9749);
and U14644 (N_14644,N_9355,N_7777);
and U14645 (N_14645,N_8205,N_6866);
and U14646 (N_14646,N_8115,N_5508);
and U14647 (N_14647,N_8393,N_9306);
nand U14648 (N_14648,N_6826,N_9534);
nand U14649 (N_14649,N_5786,N_6005);
nand U14650 (N_14650,N_9127,N_8891);
nand U14651 (N_14651,N_8085,N_7852);
and U14652 (N_14652,N_9402,N_6178);
xor U14653 (N_14653,N_5828,N_6819);
nor U14654 (N_14654,N_9942,N_8101);
and U14655 (N_14655,N_9738,N_7869);
or U14656 (N_14656,N_8006,N_7512);
nor U14657 (N_14657,N_8132,N_7034);
nand U14658 (N_14658,N_5579,N_5326);
xor U14659 (N_14659,N_7037,N_7234);
or U14660 (N_14660,N_9147,N_6158);
or U14661 (N_14661,N_5982,N_8883);
nand U14662 (N_14662,N_8421,N_5984);
and U14663 (N_14663,N_6529,N_9158);
nand U14664 (N_14664,N_5433,N_7128);
and U14665 (N_14665,N_9992,N_6410);
nand U14666 (N_14666,N_6354,N_9618);
nand U14667 (N_14667,N_6759,N_7486);
and U14668 (N_14668,N_7104,N_9202);
and U14669 (N_14669,N_8860,N_6486);
nor U14670 (N_14670,N_9368,N_7071);
and U14671 (N_14671,N_7808,N_7627);
or U14672 (N_14672,N_6606,N_6381);
xnor U14673 (N_14673,N_6595,N_8856);
and U14674 (N_14674,N_7885,N_7502);
nor U14675 (N_14675,N_5909,N_9568);
nor U14676 (N_14676,N_7991,N_5764);
nor U14677 (N_14677,N_5596,N_7906);
and U14678 (N_14678,N_6056,N_5375);
nor U14679 (N_14679,N_9194,N_8805);
nand U14680 (N_14680,N_9464,N_9790);
nor U14681 (N_14681,N_9999,N_5062);
nand U14682 (N_14682,N_7123,N_8805);
nand U14683 (N_14683,N_7576,N_9435);
nand U14684 (N_14684,N_5837,N_8917);
xor U14685 (N_14685,N_6087,N_7591);
xor U14686 (N_14686,N_7754,N_9372);
xnor U14687 (N_14687,N_9601,N_9189);
nor U14688 (N_14688,N_6819,N_8086);
nor U14689 (N_14689,N_5878,N_7668);
and U14690 (N_14690,N_6430,N_5740);
nor U14691 (N_14691,N_5267,N_5538);
nand U14692 (N_14692,N_7707,N_8069);
nor U14693 (N_14693,N_5075,N_5936);
and U14694 (N_14694,N_5225,N_6358);
xnor U14695 (N_14695,N_5789,N_9449);
and U14696 (N_14696,N_9380,N_5804);
and U14697 (N_14697,N_5412,N_8180);
or U14698 (N_14698,N_5145,N_7100);
nor U14699 (N_14699,N_9823,N_6237);
and U14700 (N_14700,N_5919,N_9602);
nand U14701 (N_14701,N_7779,N_7152);
or U14702 (N_14702,N_6373,N_5623);
xor U14703 (N_14703,N_7457,N_9215);
xnor U14704 (N_14704,N_9652,N_7116);
and U14705 (N_14705,N_6501,N_5737);
nand U14706 (N_14706,N_7480,N_8124);
and U14707 (N_14707,N_8491,N_5706);
xor U14708 (N_14708,N_5553,N_7793);
and U14709 (N_14709,N_6756,N_9341);
or U14710 (N_14710,N_5734,N_7914);
and U14711 (N_14711,N_5429,N_6671);
nand U14712 (N_14712,N_9360,N_7422);
and U14713 (N_14713,N_8459,N_8077);
xor U14714 (N_14714,N_5523,N_9310);
xnor U14715 (N_14715,N_9124,N_8930);
or U14716 (N_14716,N_9623,N_8151);
nand U14717 (N_14717,N_6864,N_5197);
nor U14718 (N_14718,N_5059,N_5545);
nand U14719 (N_14719,N_5544,N_8570);
xor U14720 (N_14720,N_8955,N_6694);
and U14721 (N_14721,N_8778,N_8315);
or U14722 (N_14722,N_9935,N_8423);
nand U14723 (N_14723,N_6161,N_5104);
and U14724 (N_14724,N_6701,N_9936);
and U14725 (N_14725,N_7666,N_6915);
and U14726 (N_14726,N_6791,N_9343);
and U14727 (N_14727,N_6026,N_8917);
nand U14728 (N_14728,N_6422,N_7379);
nand U14729 (N_14729,N_8922,N_8771);
or U14730 (N_14730,N_6798,N_6898);
xnor U14731 (N_14731,N_6263,N_8603);
or U14732 (N_14732,N_9539,N_9210);
xnor U14733 (N_14733,N_5628,N_7615);
xor U14734 (N_14734,N_9824,N_5320);
and U14735 (N_14735,N_8861,N_9289);
nor U14736 (N_14736,N_9958,N_6197);
or U14737 (N_14737,N_8412,N_9596);
or U14738 (N_14738,N_9968,N_8464);
nor U14739 (N_14739,N_6246,N_6196);
nand U14740 (N_14740,N_9500,N_6903);
nand U14741 (N_14741,N_5340,N_8765);
and U14742 (N_14742,N_7392,N_5942);
nand U14743 (N_14743,N_7281,N_9821);
nor U14744 (N_14744,N_6408,N_6949);
or U14745 (N_14745,N_7993,N_8050);
nor U14746 (N_14746,N_8545,N_9026);
xor U14747 (N_14747,N_8726,N_5117);
nor U14748 (N_14748,N_6017,N_9270);
nand U14749 (N_14749,N_6808,N_5498);
nand U14750 (N_14750,N_9665,N_6383);
nor U14751 (N_14751,N_7718,N_6683);
or U14752 (N_14752,N_9279,N_8083);
or U14753 (N_14753,N_9812,N_5464);
and U14754 (N_14754,N_6337,N_7160);
nor U14755 (N_14755,N_9180,N_6588);
and U14756 (N_14756,N_9468,N_8210);
and U14757 (N_14757,N_5968,N_6341);
or U14758 (N_14758,N_5789,N_9569);
xor U14759 (N_14759,N_9753,N_9489);
and U14760 (N_14760,N_8694,N_6176);
or U14761 (N_14761,N_6268,N_5051);
xor U14762 (N_14762,N_8598,N_7413);
nor U14763 (N_14763,N_7697,N_8589);
xor U14764 (N_14764,N_6404,N_8254);
and U14765 (N_14765,N_9116,N_7605);
or U14766 (N_14766,N_6826,N_6266);
xnor U14767 (N_14767,N_6375,N_6471);
and U14768 (N_14768,N_7047,N_8628);
or U14769 (N_14769,N_9744,N_6061);
nor U14770 (N_14770,N_6912,N_8623);
nand U14771 (N_14771,N_9238,N_8824);
nor U14772 (N_14772,N_9316,N_6387);
nor U14773 (N_14773,N_6052,N_6517);
nor U14774 (N_14774,N_6049,N_9138);
or U14775 (N_14775,N_6699,N_6596);
nor U14776 (N_14776,N_6889,N_5120);
and U14777 (N_14777,N_5554,N_8156);
nor U14778 (N_14778,N_9668,N_7891);
nor U14779 (N_14779,N_9356,N_7126);
xor U14780 (N_14780,N_8153,N_5368);
or U14781 (N_14781,N_7573,N_9285);
or U14782 (N_14782,N_9558,N_5900);
nand U14783 (N_14783,N_5961,N_7962);
nor U14784 (N_14784,N_6214,N_6123);
nand U14785 (N_14785,N_9347,N_5886);
nand U14786 (N_14786,N_9163,N_7080);
nor U14787 (N_14787,N_5944,N_6445);
nor U14788 (N_14788,N_6951,N_6554);
xor U14789 (N_14789,N_9001,N_7301);
and U14790 (N_14790,N_7145,N_7159);
nor U14791 (N_14791,N_9946,N_5197);
and U14792 (N_14792,N_8169,N_8553);
xor U14793 (N_14793,N_9231,N_6632);
nand U14794 (N_14794,N_9304,N_5812);
nand U14795 (N_14795,N_8636,N_8808);
and U14796 (N_14796,N_9980,N_9835);
and U14797 (N_14797,N_9960,N_5572);
xnor U14798 (N_14798,N_5913,N_6808);
or U14799 (N_14799,N_8778,N_8557);
nand U14800 (N_14800,N_8123,N_7273);
and U14801 (N_14801,N_5702,N_6438);
and U14802 (N_14802,N_5870,N_9444);
and U14803 (N_14803,N_8144,N_6049);
xor U14804 (N_14804,N_9243,N_5354);
or U14805 (N_14805,N_6420,N_9810);
nand U14806 (N_14806,N_9783,N_6621);
nor U14807 (N_14807,N_6332,N_6413);
nand U14808 (N_14808,N_5903,N_9956);
nor U14809 (N_14809,N_9709,N_9876);
or U14810 (N_14810,N_9011,N_5723);
nand U14811 (N_14811,N_8897,N_7634);
nand U14812 (N_14812,N_7621,N_9483);
or U14813 (N_14813,N_5835,N_7036);
and U14814 (N_14814,N_6041,N_6895);
or U14815 (N_14815,N_9490,N_5347);
or U14816 (N_14816,N_7957,N_6294);
and U14817 (N_14817,N_8047,N_7812);
nor U14818 (N_14818,N_9824,N_7422);
and U14819 (N_14819,N_8778,N_5174);
xnor U14820 (N_14820,N_8788,N_5669);
nor U14821 (N_14821,N_5261,N_5361);
nor U14822 (N_14822,N_8302,N_8090);
nor U14823 (N_14823,N_8615,N_5513);
and U14824 (N_14824,N_9471,N_5181);
nor U14825 (N_14825,N_5375,N_7707);
or U14826 (N_14826,N_8883,N_9942);
nand U14827 (N_14827,N_9546,N_7265);
xor U14828 (N_14828,N_7703,N_6224);
nand U14829 (N_14829,N_6370,N_7015);
and U14830 (N_14830,N_5737,N_6749);
nand U14831 (N_14831,N_7172,N_9703);
or U14832 (N_14832,N_8822,N_8438);
xor U14833 (N_14833,N_7022,N_6710);
nand U14834 (N_14834,N_9196,N_9624);
nor U14835 (N_14835,N_9960,N_8901);
nor U14836 (N_14836,N_7145,N_5800);
or U14837 (N_14837,N_6638,N_6426);
or U14838 (N_14838,N_9436,N_6187);
nand U14839 (N_14839,N_6866,N_9047);
or U14840 (N_14840,N_7590,N_7651);
and U14841 (N_14841,N_6472,N_7428);
xor U14842 (N_14842,N_6550,N_8789);
or U14843 (N_14843,N_5087,N_8093);
nor U14844 (N_14844,N_5125,N_5702);
nand U14845 (N_14845,N_8669,N_8766);
nand U14846 (N_14846,N_5433,N_9176);
and U14847 (N_14847,N_8684,N_7126);
nor U14848 (N_14848,N_8992,N_9140);
xnor U14849 (N_14849,N_5083,N_7304);
or U14850 (N_14850,N_6307,N_7042);
nand U14851 (N_14851,N_5212,N_5857);
or U14852 (N_14852,N_6555,N_5159);
xnor U14853 (N_14853,N_6848,N_5689);
and U14854 (N_14854,N_8744,N_5956);
nor U14855 (N_14855,N_7138,N_9425);
and U14856 (N_14856,N_7113,N_7517);
xor U14857 (N_14857,N_7265,N_9510);
and U14858 (N_14858,N_5206,N_7052);
nand U14859 (N_14859,N_6071,N_6228);
nor U14860 (N_14860,N_5015,N_8892);
and U14861 (N_14861,N_5725,N_5245);
or U14862 (N_14862,N_6712,N_7155);
or U14863 (N_14863,N_6622,N_8614);
nand U14864 (N_14864,N_8028,N_6887);
and U14865 (N_14865,N_7724,N_9810);
and U14866 (N_14866,N_7092,N_5617);
xor U14867 (N_14867,N_5005,N_8160);
xnor U14868 (N_14868,N_8109,N_6516);
nor U14869 (N_14869,N_5148,N_6655);
or U14870 (N_14870,N_9281,N_8229);
xor U14871 (N_14871,N_6659,N_9257);
xnor U14872 (N_14872,N_6969,N_7597);
nor U14873 (N_14873,N_8534,N_8304);
nand U14874 (N_14874,N_6916,N_7219);
nand U14875 (N_14875,N_7915,N_6954);
xnor U14876 (N_14876,N_8097,N_5460);
nor U14877 (N_14877,N_7910,N_6336);
nand U14878 (N_14878,N_9518,N_8003);
nor U14879 (N_14879,N_6718,N_9031);
xor U14880 (N_14880,N_5937,N_5827);
xnor U14881 (N_14881,N_8482,N_7940);
or U14882 (N_14882,N_5073,N_9924);
xor U14883 (N_14883,N_7633,N_5630);
or U14884 (N_14884,N_5619,N_7886);
xor U14885 (N_14885,N_7646,N_5889);
and U14886 (N_14886,N_5277,N_6738);
nand U14887 (N_14887,N_6848,N_8922);
xnor U14888 (N_14888,N_9251,N_7616);
nor U14889 (N_14889,N_9044,N_9550);
xor U14890 (N_14890,N_8972,N_9714);
nand U14891 (N_14891,N_7563,N_7913);
and U14892 (N_14892,N_8804,N_9220);
nor U14893 (N_14893,N_7754,N_8031);
xnor U14894 (N_14894,N_7701,N_9804);
or U14895 (N_14895,N_6546,N_6032);
xnor U14896 (N_14896,N_9230,N_8396);
nor U14897 (N_14897,N_7923,N_5609);
xnor U14898 (N_14898,N_9013,N_9371);
and U14899 (N_14899,N_8045,N_5865);
and U14900 (N_14900,N_8869,N_9677);
or U14901 (N_14901,N_7921,N_5975);
xnor U14902 (N_14902,N_8531,N_5179);
and U14903 (N_14903,N_8718,N_7397);
nand U14904 (N_14904,N_7065,N_5233);
xor U14905 (N_14905,N_5277,N_8874);
xor U14906 (N_14906,N_8833,N_8898);
nand U14907 (N_14907,N_5631,N_7386);
nand U14908 (N_14908,N_6609,N_7103);
nand U14909 (N_14909,N_6219,N_9732);
xnor U14910 (N_14910,N_7020,N_5137);
nor U14911 (N_14911,N_9028,N_7335);
or U14912 (N_14912,N_8048,N_9544);
and U14913 (N_14913,N_9529,N_5493);
xor U14914 (N_14914,N_8720,N_5657);
or U14915 (N_14915,N_5443,N_6616);
nand U14916 (N_14916,N_6435,N_7373);
nand U14917 (N_14917,N_6416,N_9692);
and U14918 (N_14918,N_6678,N_7981);
xnor U14919 (N_14919,N_8569,N_9640);
or U14920 (N_14920,N_5473,N_8521);
xnor U14921 (N_14921,N_8237,N_8372);
and U14922 (N_14922,N_5636,N_7843);
and U14923 (N_14923,N_8271,N_9021);
xor U14924 (N_14924,N_9926,N_6370);
nor U14925 (N_14925,N_9441,N_5121);
nor U14926 (N_14926,N_8416,N_7138);
and U14927 (N_14927,N_5703,N_8006);
nor U14928 (N_14928,N_6743,N_6307);
or U14929 (N_14929,N_6938,N_7699);
nand U14930 (N_14930,N_6485,N_7931);
and U14931 (N_14931,N_7747,N_5520);
nor U14932 (N_14932,N_6656,N_7961);
and U14933 (N_14933,N_9791,N_6433);
xnor U14934 (N_14934,N_9527,N_6730);
or U14935 (N_14935,N_7721,N_5611);
nand U14936 (N_14936,N_6242,N_8140);
nand U14937 (N_14937,N_8528,N_7057);
nor U14938 (N_14938,N_7606,N_6051);
nand U14939 (N_14939,N_9614,N_9717);
nor U14940 (N_14940,N_7860,N_8224);
xnor U14941 (N_14941,N_6022,N_8171);
or U14942 (N_14942,N_5547,N_5150);
and U14943 (N_14943,N_9719,N_5816);
and U14944 (N_14944,N_5822,N_7769);
nor U14945 (N_14945,N_8106,N_5604);
nor U14946 (N_14946,N_6904,N_8390);
nor U14947 (N_14947,N_7206,N_5646);
xor U14948 (N_14948,N_8575,N_7855);
nand U14949 (N_14949,N_6163,N_6937);
nand U14950 (N_14950,N_8468,N_7850);
nand U14951 (N_14951,N_7580,N_7784);
and U14952 (N_14952,N_6878,N_9421);
nor U14953 (N_14953,N_6843,N_9570);
or U14954 (N_14954,N_7469,N_7151);
or U14955 (N_14955,N_9864,N_7878);
and U14956 (N_14956,N_7026,N_5472);
or U14957 (N_14957,N_5433,N_7728);
xnor U14958 (N_14958,N_6301,N_5226);
xor U14959 (N_14959,N_5411,N_5405);
and U14960 (N_14960,N_9625,N_9667);
or U14961 (N_14961,N_7917,N_5991);
nor U14962 (N_14962,N_9939,N_7612);
or U14963 (N_14963,N_8018,N_7078);
nor U14964 (N_14964,N_9462,N_5220);
xor U14965 (N_14965,N_7984,N_5018);
xnor U14966 (N_14966,N_5212,N_7849);
or U14967 (N_14967,N_7452,N_8083);
nor U14968 (N_14968,N_8323,N_6120);
and U14969 (N_14969,N_7186,N_6575);
nand U14970 (N_14970,N_9793,N_7898);
xnor U14971 (N_14971,N_6956,N_7692);
or U14972 (N_14972,N_9900,N_6883);
nand U14973 (N_14973,N_8061,N_7923);
or U14974 (N_14974,N_5210,N_6963);
xor U14975 (N_14975,N_7750,N_8741);
nand U14976 (N_14976,N_5293,N_6709);
nand U14977 (N_14977,N_5233,N_9354);
and U14978 (N_14978,N_8590,N_6687);
xnor U14979 (N_14979,N_5748,N_7847);
or U14980 (N_14980,N_5836,N_5630);
nor U14981 (N_14981,N_9480,N_6626);
or U14982 (N_14982,N_8634,N_8413);
or U14983 (N_14983,N_6626,N_8095);
nor U14984 (N_14984,N_8071,N_5700);
nand U14985 (N_14985,N_6860,N_8498);
nor U14986 (N_14986,N_5261,N_6035);
or U14987 (N_14987,N_6161,N_7706);
nor U14988 (N_14988,N_7247,N_5260);
xnor U14989 (N_14989,N_6308,N_8278);
and U14990 (N_14990,N_7048,N_5256);
xor U14991 (N_14991,N_5922,N_5640);
xor U14992 (N_14992,N_7089,N_5941);
nand U14993 (N_14993,N_7957,N_6839);
xor U14994 (N_14994,N_9968,N_9194);
nor U14995 (N_14995,N_9856,N_5857);
and U14996 (N_14996,N_8999,N_9827);
or U14997 (N_14997,N_5260,N_5376);
nand U14998 (N_14998,N_8245,N_7191);
nor U14999 (N_14999,N_6433,N_7021);
or U15000 (N_15000,N_10906,N_14145);
xor U15001 (N_15001,N_12355,N_13264);
or U15002 (N_15002,N_14189,N_13132);
or U15003 (N_15003,N_13871,N_11078);
nor U15004 (N_15004,N_11917,N_13350);
and U15005 (N_15005,N_14679,N_12359);
nor U15006 (N_15006,N_14912,N_10744);
nor U15007 (N_15007,N_13488,N_13353);
or U15008 (N_15008,N_11308,N_12361);
xnor U15009 (N_15009,N_14453,N_13303);
and U15010 (N_15010,N_13276,N_14202);
nand U15011 (N_15011,N_13222,N_10391);
nand U15012 (N_15012,N_13467,N_13472);
nor U15013 (N_15013,N_13852,N_11574);
xnor U15014 (N_15014,N_10904,N_11492);
xor U15015 (N_15015,N_13363,N_13967);
and U15016 (N_15016,N_13802,N_13249);
or U15017 (N_15017,N_11581,N_10644);
or U15018 (N_15018,N_10717,N_10945);
nor U15019 (N_15019,N_13692,N_14007);
nor U15020 (N_15020,N_13855,N_10829);
or U15021 (N_15021,N_12810,N_14770);
and U15022 (N_15022,N_12216,N_13922);
xor U15023 (N_15023,N_13447,N_12177);
nand U15024 (N_15024,N_12090,N_11448);
xor U15025 (N_15025,N_10460,N_12271);
or U15026 (N_15026,N_14265,N_10121);
or U15027 (N_15027,N_14290,N_10014);
nor U15028 (N_15028,N_12579,N_10055);
and U15029 (N_15029,N_14363,N_14199);
nand U15030 (N_15030,N_14087,N_11591);
or U15031 (N_15031,N_10238,N_13816);
nor U15032 (N_15032,N_10349,N_11199);
or U15033 (N_15033,N_11541,N_11179);
or U15034 (N_15034,N_11182,N_13448);
and U15035 (N_15035,N_11024,N_13574);
xor U15036 (N_15036,N_14262,N_11374);
nor U15037 (N_15037,N_12136,N_14218);
nand U15038 (N_15038,N_13780,N_10513);
nor U15039 (N_15039,N_14157,N_10506);
nor U15040 (N_15040,N_14201,N_11515);
xor U15041 (N_15041,N_14236,N_10366);
xnor U15042 (N_15042,N_13212,N_10448);
xnor U15043 (N_15043,N_13845,N_11465);
or U15044 (N_15044,N_13422,N_12161);
nor U15045 (N_15045,N_12829,N_11631);
nand U15046 (N_15046,N_11955,N_12235);
or U15047 (N_15047,N_11503,N_12566);
and U15048 (N_15048,N_11552,N_13801);
nor U15049 (N_15049,N_11178,N_11248);
xnor U15050 (N_15050,N_13201,N_11212);
nand U15051 (N_15051,N_13951,N_12528);
xor U15052 (N_15052,N_12595,N_13044);
and U15053 (N_15053,N_11932,N_11081);
nor U15054 (N_15054,N_14254,N_13256);
and U15055 (N_15055,N_11243,N_12378);
xor U15056 (N_15056,N_10043,N_14962);
nor U15057 (N_15057,N_12201,N_13195);
nand U15058 (N_15058,N_14360,N_12236);
xnor U15059 (N_15059,N_10673,N_10364);
or U15060 (N_15060,N_11305,N_12521);
xor U15061 (N_15061,N_12312,N_12739);
or U15062 (N_15062,N_11033,N_13618);
and U15063 (N_15063,N_10503,N_10462);
or U15064 (N_15064,N_13300,N_10346);
and U15065 (N_15065,N_10425,N_11923);
nor U15066 (N_15066,N_14424,N_11766);
xnor U15067 (N_15067,N_11071,N_12200);
nor U15068 (N_15068,N_11003,N_12217);
nand U15069 (N_15069,N_10843,N_13073);
xor U15070 (N_15070,N_10167,N_11519);
xnor U15071 (N_15071,N_11018,N_11043);
xor U15072 (N_15072,N_12910,N_13068);
xor U15073 (N_15073,N_14818,N_13035);
nor U15074 (N_15074,N_10698,N_10863);
nor U15075 (N_15075,N_13748,N_12133);
and U15076 (N_15076,N_11440,N_12655);
nor U15077 (N_15077,N_14474,N_12961);
and U15078 (N_15078,N_14824,N_10041);
nor U15079 (N_15079,N_12466,N_13888);
or U15080 (N_15080,N_12852,N_11936);
nor U15081 (N_15081,N_12730,N_13808);
and U15082 (N_15082,N_13456,N_12727);
xnor U15083 (N_15083,N_13483,N_12827);
nand U15084 (N_15084,N_14647,N_14162);
xnor U15085 (N_15085,N_13439,N_13588);
xor U15086 (N_15086,N_13108,N_12875);
nor U15087 (N_15087,N_12454,N_14657);
nor U15088 (N_15088,N_12295,N_14811);
and U15089 (N_15089,N_10988,N_12652);
and U15090 (N_15090,N_10684,N_13309);
or U15091 (N_15091,N_12221,N_12174);
nand U15092 (N_15092,N_10216,N_11136);
xnor U15093 (N_15093,N_11262,N_14552);
nand U15094 (N_15094,N_11066,N_13160);
and U15095 (N_15095,N_11909,N_13968);
nand U15096 (N_15096,N_12607,N_11617);
and U15097 (N_15097,N_10679,N_12823);
xnor U15098 (N_15098,N_10831,N_10812);
xor U15099 (N_15099,N_10617,N_12463);
and U15100 (N_15100,N_10686,N_11446);
xor U15101 (N_15101,N_13873,N_10849);
xnor U15102 (N_15102,N_12125,N_11569);
nand U15103 (N_15103,N_13513,N_14547);
and U15104 (N_15104,N_12694,N_11694);
or U15105 (N_15105,N_10984,N_12198);
nand U15106 (N_15106,N_10955,N_13462);
and U15107 (N_15107,N_13174,N_11566);
nor U15108 (N_15108,N_11313,N_12564);
nand U15109 (N_15109,N_14367,N_11925);
nor U15110 (N_15110,N_13479,N_11233);
and U15111 (N_15111,N_13928,N_14689);
nor U15112 (N_15112,N_11323,N_11473);
nand U15113 (N_15113,N_12879,N_10193);
xnor U15114 (N_15114,N_11482,N_13964);
or U15115 (N_15115,N_11603,N_11301);
or U15116 (N_15116,N_14816,N_14815);
nand U15117 (N_15117,N_13323,N_14739);
xnor U15118 (N_15118,N_12003,N_12542);
and U15119 (N_15119,N_11501,N_12726);
and U15120 (N_15120,N_10806,N_10642);
nand U15121 (N_15121,N_12797,N_10900);
and U15122 (N_15122,N_13321,N_11629);
nand U15123 (N_15123,N_12949,N_12316);
xnor U15124 (N_15124,N_10212,N_12212);
xor U15125 (N_15125,N_10790,N_12213);
xnor U15126 (N_15126,N_13616,N_12620);
nor U15127 (N_15127,N_14943,N_14208);
and U15128 (N_15128,N_11389,N_10763);
xnor U15129 (N_15129,N_13787,N_13807);
and U15130 (N_15130,N_13476,N_12258);
nand U15131 (N_15131,N_13115,N_12414);
nor U15132 (N_15132,N_12379,N_13356);
xor U15133 (N_15133,N_12028,N_11572);
nor U15134 (N_15134,N_13361,N_11823);
nor U15135 (N_15135,N_11284,N_11056);
or U15136 (N_15136,N_12168,N_13082);
nor U15137 (N_15137,N_10409,N_10809);
nor U15138 (N_15138,N_12900,N_12390);
nand U15139 (N_15139,N_12979,N_14089);
and U15140 (N_15140,N_10682,N_13484);
and U15141 (N_15141,N_10530,N_12822);
nand U15142 (N_15142,N_12269,N_14873);
or U15143 (N_15143,N_12496,N_13952);
or U15144 (N_15144,N_13294,N_10241);
and U15145 (N_15145,N_11029,N_14871);
and U15146 (N_15146,N_14836,N_12101);
nor U15147 (N_15147,N_10217,N_14413);
xor U15148 (N_15148,N_11757,N_14005);
or U15149 (N_15149,N_12464,N_12742);
and U15150 (N_15150,N_11759,N_14538);
and U15151 (N_15151,N_13750,N_13796);
nor U15152 (N_15152,N_10493,N_12479);
nor U15153 (N_15153,N_10836,N_10243);
nor U15154 (N_15154,N_10404,N_13665);
xor U15155 (N_15155,N_12530,N_11824);
nor U15156 (N_15156,N_13494,N_14350);
and U15157 (N_15157,N_14707,N_14083);
or U15158 (N_15158,N_12184,N_11135);
nand U15159 (N_15159,N_12056,N_13288);
nor U15160 (N_15160,N_10034,N_14206);
xor U15161 (N_15161,N_13349,N_13176);
xor U15162 (N_15162,N_13271,N_11838);
or U15163 (N_15163,N_11228,N_12292);
nand U15164 (N_15164,N_11525,N_11847);
nand U15165 (N_15165,N_10279,N_14584);
nand U15166 (N_15166,N_12305,N_12684);
nor U15167 (N_15167,N_13755,N_10368);
nor U15168 (N_15168,N_13630,N_13345);
nor U15169 (N_15169,N_11609,N_12369);
and U15170 (N_15170,N_14765,N_10050);
or U15171 (N_15171,N_13708,N_13614);
nand U15172 (N_15172,N_12938,N_12882);
nor U15173 (N_15173,N_10875,N_12318);
xor U15174 (N_15174,N_14263,N_13219);
and U15175 (N_15175,N_14428,N_10467);
or U15176 (N_15176,N_14183,N_12724);
nand U15177 (N_15177,N_12105,N_10278);
xor U15178 (N_15178,N_11297,N_11467);
or U15179 (N_15179,N_13088,N_10886);
or U15180 (N_15180,N_13703,N_13338);
and U15181 (N_15181,N_12605,N_13604);
or U15182 (N_15182,N_14196,N_10242);
or U15183 (N_15183,N_14421,N_10736);
or U15184 (N_15184,N_12300,N_10520);
and U15185 (N_15185,N_12476,N_14127);
xor U15186 (N_15186,N_12130,N_12923);
nor U15187 (N_15187,N_11662,N_13835);
nand U15188 (N_15188,N_11736,N_11578);
nand U15189 (N_15189,N_14193,N_12232);
xor U15190 (N_15190,N_14370,N_12188);
nand U15191 (N_15191,N_13105,N_12919);
or U15192 (N_15192,N_12218,N_11557);
and U15193 (N_15193,N_12254,N_14135);
nor U15194 (N_15194,N_13072,N_12612);
nand U15195 (N_15195,N_12935,N_14351);
nand U15196 (N_15196,N_14927,N_13122);
xnor U15197 (N_15197,N_12012,N_13840);
nand U15198 (N_15198,N_12229,N_14275);
nand U15199 (N_15199,N_13999,N_14148);
nand U15200 (N_15200,N_10224,N_12341);
and U15201 (N_15201,N_13490,N_10463);
and U15202 (N_15202,N_14492,N_13150);
nor U15203 (N_15203,N_10525,N_10942);
or U15204 (N_15204,N_13648,N_14706);
xnor U15205 (N_15205,N_12976,N_14016);
nor U15206 (N_15206,N_11967,N_13365);
xnor U15207 (N_15207,N_10997,N_13799);
and U15208 (N_15208,N_11762,N_14156);
or U15209 (N_15209,N_11677,N_14524);
and U15210 (N_15210,N_11359,N_12909);
nor U15211 (N_15211,N_11741,N_11845);
nand U15212 (N_15212,N_14408,N_11663);
xnor U15213 (N_15213,N_11969,N_13442);
and U15214 (N_15214,N_13981,N_14956);
nor U15215 (N_15215,N_11983,N_10813);
nor U15216 (N_15216,N_14153,N_12145);
or U15217 (N_15217,N_11386,N_13400);
nand U15218 (N_15218,N_14881,N_10962);
nor U15219 (N_15219,N_11979,N_14397);
xnor U15220 (N_15220,N_10202,N_10350);
nor U15221 (N_15221,N_11045,N_12363);
nand U15222 (N_15222,N_11690,N_13501);
and U15223 (N_15223,N_12782,N_14844);
nand U15224 (N_15224,N_11257,N_11192);
nor U15225 (N_15225,N_14061,N_11089);
or U15226 (N_15226,N_14745,N_13929);
nor U15227 (N_15227,N_11711,N_12665);
xor U15228 (N_15228,N_14638,N_12748);
nand U15229 (N_15229,N_14551,N_13909);
or U15230 (N_15230,N_14581,N_12706);
and U15231 (N_15231,N_10189,N_14555);
nor U15232 (N_15232,N_10626,N_14800);
or U15233 (N_15233,N_14920,N_13992);
nor U15234 (N_15234,N_10606,N_14597);
nand U15235 (N_15235,N_14170,N_13744);
and U15236 (N_15236,N_14674,N_11851);
xnor U15237 (N_15237,N_14839,N_13553);
and U15238 (N_15238,N_12862,N_12131);
nand U15239 (N_15239,N_13587,N_12962);
nor U15240 (N_15240,N_14308,N_13403);
nor U15241 (N_15241,N_13585,N_10000);
nor U15242 (N_15242,N_10133,N_12601);
or U15243 (N_15243,N_14591,N_10758);
nand U15244 (N_15244,N_10430,N_10411);
xnor U15245 (N_15245,N_11250,N_11122);
and U15246 (N_15246,N_12769,N_14966);
nor U15247 (N_15247,N_14009,N_14435);
and U15248 (N_15248,N_11328,N_12166);
and U15249 (N_15249,N_14728,N_10010);
and U15250 (N_15250,N_14166,N_12786);
nor U15251 (N_15251,N_12425,N_13084);
xor U15252 (N_15252,N_14971,N_12745);
and U15253 (N_15253,N_12076,N_10447);
nor U15254 (N_15254,N_13916,N_11221);
or U15255 (N_15255,N_13385,N_10885);
nor U15256 (N_15256,N_10678,N_13600);
xnor U15257 (N_15257,N_14338,N_12273);
xnor U15258 (N_15258,N_13743,N_13079);
nor U15259 (N_15259,N_11709,N_13012);
or U15260 (N_15260,N_12465,N_12907);
xnor U15261 (N_15261,N_10687,N_14282);
nand U15262 (N_15262,N_13567,N_12847);
and U15263 (N_15263,N_10001,N_12195);
and U15264 (N_15264,N_11937,N_10372);
and U15265 (N_15265,N_14169,N_11527);
nor U15266 (N_15266,N_10514,N_10970);
nand U15267 (N_15267,N_14255,N_10799);
and U15268 (N_15268,N_14964,N_14138);
xor U15269 (N_15269,N_10239,N_13949);
and U15270 (N_15270,N_14493,N_10966);
nand U15271 (N_15271,N_12828,N_14081);
xnor U15272 (N_15272,N_14215,N_10180);
xnor U15273 (N_15273,N_10648,N_10097);
xor U15274 (N_15274,N_10311,N_10027);
or U15275 (N_15275,N_10754,N_14194);
and U15276 (N_15276,N_12324,N_12659);
xor U15277 (N_15277,N_14102,N_10316);
nor U15278 (N_15278,N_13507,N_14411);
nor U15279 (N_15279,N_14395,N_13039);
nand U15280 (N_15280,N_10594,N_11201);
or U15281 (N_15281,N_14496,N_10414);
and U15282 (N_15282,N_11831,N_13113);
and U15283 (N_15283,N_13404,N_11115);
or U15284 (N_15284,N_13629,N_10558);
nor U15285 (N_15285,N_11790,N_12830);
and U15286 (N_15286,N_10492,N_10473);
and U15287 (N_15287,N_10570,N_14082);
nor U15288 (N_15288,N_14313,N_13701);
nor U15289 (N_15289,N_12973,N_13924);
nand U15290 (N_15290,N_13517,N_13671);
or U15291 (N_15291,N_11700,N_11502);
xnor U15292 (N_15292,N_13684,N_11614);
xnor U15293 (N_15293,N_13340,N_11131);
or U15294 (N_15294,N_10441,N_12833);
xnor U15295 (N_15295,N_14374,N_12880);
and U15296 (N_15296,N_10047,N_10561);
nor U15297 (N_15297,N_12768,N_11140);
or U15298 (N_15298,N_12146,N_10168);
nand U15299 (N_15299,N_11746,N_10619);
nor U15300 (N_15300,N_13912,N_10928);
xnor U15301 (N_15301,N_12332,N_13454);
nor U15302 (N_15302,N_11317,N_12557);
and U15303 (N_15303,N_12908,N_13654);
nand U15304 (N_15304,N_11375,N_11994);
or U15305 (N_15305,N_12123,N_13142);
nor U15306 (N_15306,N_13984,N_12013);
and U15307 (N_15307,N_10177,N_12721);
nand U15308 (N_15308,N_11723,N_13866);
nor U15309 (N_15309,N_12328,N_14857);
xor U15310 (N_15310,N_11849,N_10490);
xor U15311 (N_15311,N_11940,N_12443);
or U15312 (N_15312,N_14781,N_14326);
or U15313 (N_15313,N_13825,N_12290);
nor U15314 (N_15314,N_11283,N_11725);
xor U15315 (N_15315,N_14810,N_14304);
nor U15316 (N_15316,N_11894,N_12794);
or U15317 (N_15317,N_10085,N_13137);
or U15318 (N_15318,N_12365,N_10737);
nand U15319 (N_15319,N_13861,N_12686);
nand U15320 (N_15320,N_13184,N_14832);
and U15321 (N_15321,N_13257,N_10280);
nand U15322 (N_15322,N_13192,N_13465);
nand U15323 (N_15323,N_14510,N_12920);
nor U15324 (N_15324,N_10868,N_10780);
nand U15325 (N_15325,N_10537,N_12696);
nor U15326 (N_15326,N_13579,N_14334);
and U15327 (N_15327,N_11927,N_12209);
and U15328 (N_15328,N_11092,N_14669);
xor U15329 (N_15329,N_13186,N_13894);
nor U15330 (N_15330,N_10021,N_11431);
xor U15331 (N_15331,N_13458,N_10127);
xnor U15332 (N_15332,N_14149,N_12106);
or U15333 (N_15333,N_12197,N_10884);
and U15334 (N_15334,N_13591,N_11883);
nand U15335 (N_15335,N_14192,N_13489);
or U15336 (N_15336,N_10516,N_13175);
xor U15337 (N_15337,N_14921,N_14767);
or U15338 (N_15338,N_11010,N_13738);
xor U15339 (N_15339,N_13895,N_11447);
nand U15340 (N_15340,N_11854,N_10547);
or U15341 (N_15341,N_12912,N_13634);
xor U15342 (N_15342,N_12052,N_10795);
nor U15343 (N_15343,N_13480,N_11890);
and U15344 (N_15344,N_12819,N_10774);
and U15345 (N_15345,N_11806,N_14348);
nor U15346 (N_15346,N_14385,N_10089);
nand U15347 (N_15347,N_12152,N_10924);
or U15348 (N_15348,N_11480,N_12417);
nand U15349 (N_15349,N_13767,N_13390);
nand U15350 (N_15350,N_10339,N_12301);
nand U15351 (N_15351,N_11127,N_10670);
and U15352 (N_15352,N_12362,N_13182);
xor U15353 (N_15353,N_11751,N_11015);
and U15354 (N_15354,N_12395,N_12821);
or U15355 (N_15355,N_14834,N_14572);
nor U15356 (N_15356,N_11347,N_13948);
or U15357 (N_15357,N_11827,N_14251);
or U15358 (N_15358,N_13341,N_12594);
or U15359 (N_15359,N_14177,N_11175);
nand U15360 (N_15360,N_14349,N_11442);
or U15361 (N_15361,N_13104,N_10272);
and U15362 (N_15362,N_14429,N_14048);
xor U15363 (N_15363,N_13236,N_11429);
and U15364 (N_15364,N_12474,N_12538);
nand U15365 (N_15365,N_14633,N_14827);
xnor U15366 (N_15366,N_10011,N_14682);
nor U15367 (N_15367,N_10161,N_12715);
and U15368 (N_15368,N_10325,N_10173);
xor U15369 (N_15369,N_13497,N_10740);
nor U15370 (N_15370,N_14627,N_11765);
or U15371 (N_15371,N_10559,N_14112);
or U15372 (N_15372,N_12311,N_14204);
nor U15373 (N_15373,N_10521,N_10484);
nand U15374 (N_15374,N_14143,N_13689);
or U15375 (N_15375,N_12906,N_10752);
nand U15376 (N_15376,N_11195,N_11848);
and U15377 (N_15377,N_11781,N_11906);
or U15378 (N_15378,N_11684,N_10295);
or U15379 (N_15379,N_11732,N_11764);
or U15380 (N_15380,N_11640,N_11914);
or U15381 (N_15381,N_14527,N_13387);
and U15382 (N_15382,N_10528,N_10823);
and U15383 (N_15383,N_10319,N_13204);
or U15384 (N_15384,N_11035,N_14136);
nor U15385 (N_15385,N_11106,N_13890);
or U15386 (N_15386,N_11880,N_14354);
and U15387 (N_15387,N_13089,N_13183);
nand U15388 (N_15388,N_12658,N_12791);
nor U15389 (N_15389,N_11793,N_13324);
nand U15390 (N_15390,N_12939,N_10902);
and U15391 (N_15391,N_10661,N_10363);
nor U15392 (N_15392,N_11084,N_10361);
and U15393 (N_15393,N_10292,N_12243);
xnor U15394 (N_15394,N_14771,N_11961);
xor U15395 (N_15395,N_13557,N_12593);
or U15396 (N_15396,N_11722,N_14986);
nor U15397 (N_15397,N_13749,N_13788);
and U15398 (N_15398,N_14219,N_12038);
and U15399 (N_15399,N_12616,N_13413);
or U15400 (N_15400,N_11338,N_10927);
nand U15401 (N_15401,N_13207,N_14992);
and U15402 (N_15402,N_13884,N_10342);
and U15403 (N_15403,N_14903,N_12484);
or U15404 (N_15404,N_10287,N_13058);
nor U15405 (N_15405,N_13487,N_14649);
nor U15406 (N_15406,N_11796,N_10304);
nor U15407 (N_15407,N_11051,N_14936);
and U15408 (N_15408,N_14783,N_10200);
and U15409 (N_15409,N_12965,N_13011);
or U15410 (N_15410,N_14715,N_12568);
nand U15411 (N_15411,N_11786,N_11679);
and U15412 (N_15412,N_13540,N_14681);
or U15413 (N_15413,N_14457,N_10921);
xnor U15414 (N_15414,N_14002,N_10699);
nor U15415 (N_15415,N_13102,N_10785);
or U15416 (N_15416,N_13197,N_10922);
nand U15417 (N_15417,N_13793,N_13357);
or U15418 (N_15418,N_10851,N_10871);
nor U15419 (N_15419,N_11871,N_14644);
nand U15420 (N_15420,N_11256,N_11820);
and U15421 (N_15421,N_10604,N_10195);
and U15422 (N_15422,N_12119,N_14646);
and U15423 (N_15423,N_13606,N_14359);
or U15424 (N_15424,N_14299,N_10635);
nor U15425 (N_15425,N_14888,N_10783);
or U15426 (N_15426,N_11637,N_14481);
and U15427 (N_15427,N_13459,N_14032);
xnor U15428 (N_15428,N_12440,N_14065);
xnor U15429 (N_15429,N_14507,N_14747);
and U15430 (N_15430,N_11471,N_10386);
xnor U15431 (N_15431,N_12732,N_14115);
or U15432 (N_15432,N_10053,N_13921);
nand U15433 (N_15433,N_13584,N_11430);
nand U15434 (N_15434,N_13243,N_13312);
nor U15435 (N_15435,N_12241,N_14182);
or U15436 (N_15436,N_14529,N_10844);
nor U15437 (N_15437,N_14698,N_12661);
xor U15438 (N_15438,N_14173,N_11358);
nor U15439 (N_15439,N_10543,N_13461);
nor U15440 (N_15440,N_11996,N_10963);
and U15441 (N_15441,N_10383,N_12980);
nand U15442 (N_15442,N_10247,N_12222);
and U15443 (N_15443,N_14697,N_10246);
or U15444 (N_15444,N_10826,N_12750);
nand U15445 (N_15445,N_13359,N_14238);
and U15446 (N_15446,N_11718,N_12406);
nand U15447 (N_15447,N_12477,N_12924);
nor U15448 (N_15448,N_12807,N_13676);
and U15449 (N_15449,N_13158,N_10791);
nand U15450 (N_15450,N_11382,N_14101);
xor U15451 (N_15451,N_11544,N_14981);
xor U15452 (N_15452,N_13352,N_10240);
nand U15453 (N_15453,N_13966,N_10190);
nand U15454 (N_15454,N_11340,N_12124);
nor U15455 (N_15455,N_10887,N_10554);
and U15456 (N_15456,N_11329,N_11858);
and U15457 (N_15457,N_10802,N_11835);
or U15458 (N_15458,N_13171,N_10058);
or U15459 (N_15459,N_14642,N_10038);
xnor U15460 (N_15460,N_10627,N_14412);
nand U15461 (N_15461,N_14191,N_13177);
or U15462 (N_15462,N_14073,N_13469);
and U15463 (N_15463,N_10095,N_14756);
and U15464 (N_15464,N_14893,N_13499);
nand U15465 (N_15465,N_11993,N_14663);
nand U15466 (N_15466,N_10105,N_12878);
nand U15467 (N_15467,N_14445,N_10158);
nor U15468 (N_15468,N_10067,N_14417);
or U15469 (N_15469,N_10110,N_10301);
nand U15470 (N_15470,N_13609,N_13358);
nand U15471 (N_15471,N_14444,N_11885);
xor U15472 (N_15472,N_11379,N_14155);
nor U15473 (N_15473,N_13481,N_14603);
and U15474 (N_15474,N_10612,N_13640);
or U15475 (N_15475,N_11142,N_11656);
or U15476 (N_15476,N_11697,N_12237);
and U15477 (N_15477,N_12481,N_12741);
nand U15478 (N_15478,N_13935,N_14303);
and U15479 (N_15479,N_12784,N_14108);
and U15480 (N_15480,N_14675,N_11702);
and U15481 (N_15481,N_10035,N_14693);
nand U15482 (N_15482,N_10719,N_12572);
nor U15483 (N_15483,N_14383,N_10793);
and U15484 (N_15484,N_11779,N_14586);
nand U15485 (N_15485,N_14117,N_11335);
or U15486 (N_15486,N_10798,N_14643);
or U15487 (N_15487,N_13687,N_14621);
nand U15488 (N_15488,N_12422,N_13826);
or U15489 (N_15489,N_12480,N_10639);
nor U15490 (N_15490,N_14128,N_11657);
or U15491 (N_15491,N_12449,N_13166);
xnor U15492 (N_15492,N_11683,N_12508);
and U15493 (N_15493,N_12259,N_10445);
or U15494 (N_15494,N_12921,N_11494);
or U15495 (N_15495,N_10471,N_12155);
and U15496 (N_15496,N_11411,N_11238);
and U15497 (N_15497,N_12128,N_12646);
nor U15498 (N_15498,N_11783,N_10428);
or U15499 (N_15499,N_10290,N_12864);
or U15500 (N_15500,N_10006,N_11975);
or U15501 (N_15501,N_10563,N_11419);
nand U15502 (N_15502,N_12245,N_10941);
xnor U15503 (N_15503,N_10817,N_10076);
nor U15504 (N_15504,N_12497,N_10766);
nand U15505 (N_15505,N_12242,N_11346);
xnor U15506 (N_15506,N_10897,N_14568);
or U15507 (N_15507,N_10435,N_10636);
or U15508 (N_15508,N_13643,N_12096);
xnor U15509 (N_15509,N_13524,N_10165);
nand U15510 (N_15510,N_14754,N_10781);
nand U15511 (N_15511,N_10548,N_11349);
xnor U15512 (N_15512,N_10257,N_11082);
or U15513 (N_15513,N_13777,N_12954);
and U15514 (N_15514,N_14989,N_14625);
and U15515 (N_15515,N_12970,N_11154);
nor U15516 (N_15516,N_11956,N_13934);
nand U15517 (N_15517,N_10801,N_10653);
nand U15518 (N_15518,N_12825,N_10936);
and U15519 (N_15519,N_12413,N_12298);
xnor U15520 (N_15520,N_12898,N_13004);
and U15521 (N_15521,N_11073,N_14999);
nand U15522 (N_15522,N_14732,N_14592);
and U15523 (N_15523,N_11461,N_14000);
nor U15524 (N_15524,N_10078,N_11166);
or U15525 (N_15525,N_12635,N_14260);
and U15526 (N_15526,N_11675,N_12215);
nand U15527 (N_15527,N_13010,N_14123);
or U15528 (N_15528,N_11987,N_12446);
xnor U15529 (N_15529,N_11701,N_11385);
xnor U15530 (N_15530,N_10423,N_14289);
and U15531 (N_15531,N_11990,N_10703);
and U15532 (N_15532,N_14242,N_12792);
or U15533 (N_15533,N_12343,N_13814);
nor U15534 (N_15534,N_10042,N_12083);
nand U15535 (N_15535,N_12147,N_14057);
or U15536 (N_15536,N_14974,N_11132);
nand U15537 (N_15537,N_12053,N_11337);
or U15538 (N_15538,N_13371,N_11576);
and U15539 (N_15539,N_10651,N_12276);
nand U15540 (N_15540,N_14062,N_10859);
nand U15541 (N_15541,N_12151,N_14580);
or U15542 (N_15542,N_12253,N_14840);
nor U15543 (N_15543,N_12093,N_12338);
or U15544 (N_15544,N_12571,N_13080);
and U15545 (N_15545,N_13774,N_13215);
nand U15546 (N_15546,N_14332,N_12026);
nand U15547 (N_15547,N_13725,N_14051);
nor U15548 (N_15548,N_12210,N_11815);
xor U15549 (N_15549,N_11981,N_10305);
and U15550 (N_15550,N_14034,N_11560);
and U15551 (N_15551,N_11713,N_11211);
nand U15552 (N_15552,N_13147,N_10535);
nand U15553 (N_15553,N_13063,N_13263);
nor U15554 (N_15554,N_12148,N_10134);
xnor U15555 (N_15555,N_12088,N_13529);
or U15556 (N_15556,N_13210,N_12214);
nand U15557 (N_15557,N_11753,N_11546);
nand U15558 (N_15558,N_13598,N_10899);
and U15559 (N_15559,N_12224,N_12097);
and U15560 (N_15560,N_11724,N_10118);
and U15561 (N_15561,N_13728,N_11356);
nand U15562 (N_15562,N_14498,N_14550);
xor U15563 (N_15563,N_10162,N_12339);
or U15564 (N_15564,N_10958,N_14656);
or U15565 (N_15565,N_11760,N_13887);
and U15566 (N_15566,N_14323,N_14264);
nor U15567 (N_15567,N_13317,N_14132);
nand U15568 (N_15568,N_14226,N_14978);
and U15569 (N_15569,N_11226,N_13029);
xor U15570 (N_15570,N_13478,N_12626);
or U15571 (N_15571,N_11320,N_14184);
xnor U15572 (N_15572,N_10087,N_13635);
or U15573 (N_15573,N_14468,N_13958);
or U15574 (N_15574,N_10037,N_12439);
nor U15575 (N_15575,N_12040,N_10720);
xnor U15576 (N_15576,N_10775,N_10715);
xor U15577 (N_15577,N_10427,N_14768);
and U15578 (N_15578,N_11628,N_10967);
nor U15579 (N_15579,N_10013,N_12380);
nand U15580 (N_15580,N_12675,N_13696);
or U15581 (N_15581,N_14654,N_11960);
and U15582 (N_15582,N_10233,N_14594);
nor U15583 (N_15583,N_10968,N_13034);
nor U15584 (N_15584,N_12649,N_10633);
nand U15585 (N_15585,N_14353,N_13839);
and U15586 (N_15586,N_11523,N_13759);
nand U15587 (N_15587,N_13971,N_12883);
or U15588 (N_15588,N_12377,N_10874);
or U15589 (N_15589,N_11528,N_11920);
xnor U15590 (N_15590,N_12118,N_11506);
nor U15591 (N_15591,N_11155,N_14700);
nor U15592 (N_15592,N_11934,N_10100);
nand U15593 (N_15593,N_10263,N_14516);
and U15594 (N_15594,N_13970,N_14316);
xnor U15595 (N_15595,N_14628,N_12325);
nor U15596 (N_15596,N_10996,N_13070);
or U15597 (N_15597,N_10230,N_10847);
or U15598 (N_15598,N_11946,N_13700);
nor U15599 (N_15599,N_14528,N_10620);
nor U15600 (N_15600,N_10972,N_13407);
nand U15601 (N_15601,N_11548,N_12374);
or U15602 (N_15602,N_11439,N_13525);
nor U15603 (N_15603,N_13143,N_12057);
and U15604 (N_15604,N_14787,N_10568);
xnor U15605 (N_15605,N_11627,N_12738);
xnor U15606 (N_15606,N_12717,N_14632);
nand U15607 (N_15607,N_13721,N_12336);
xnor U15608 (N_15608,N_11468,N_12447);
xor U15609 (N_15609,N_12872,N_11377);
or U15610 (N_15610,N_13938,N_12710);
or U15611 (N_15611,N_10674,N_13085);
and U15612 (N_15612,N_14786,N_11837);
nor U15613 (N_15613,N_10145,N_12171);
or U15614 (N_15614,N_11067,N_12795);
xor U15615 (N_15615,N_11952,N_12238);
nor U15616 (N_15616,N_10213,N_10950);
and U15617 (N_15617,N_13240,N_11857);
nor U15618 (N_15618,N_11315,N_12922);
nor U15619 (N_15619,N_14648,N_13593);
and U15620 (N_15620,N_12399,N_14917);
xnor U15621 (N_15621,N_12297,N_10557);
or U15622 (N_15622,N_13601,N_13663);
or U15623 (N_15623,N_11869,N_11383);
nor U15624 (N_15624,N_10546,N_10975);
and U15625 (N_15625,N_14293,N_10392);
and U15626 (N_15626,N_12805,N_10671);
nand U15627 (N_15627,N_12843,N_12000);
nand U15628 (N_15628,N_11687,N_13699);
and U15629 (N_15629,N_12204,N_12504);
and U15630 (N_15630,N_12811,N_10778);
xnor U15631 (N_15631,N_11394,N_12031);
xor U15632 (N_15632,N_11710,N_13377);
nor U15633 (N_15633,N_13094,N_14110);
nand U15634 (N_15634,N_11717,N_10397);
or U15635 (N_15635,N_12002,N_13910);
or U15636 (N_15636,N_13415,N_10150);
or U15637 (N_15637,N_10419,N_14812);
nand U15638 (N_15638,N_10692,N_11597);
nand U15639 (N_15639,N_13009,N_13973);
xor U15640 (N_15640,N_13021,N_12746);
and U15641 (N_15641,N_10070,N_10009);
xor U15642 (N_15642,N_13847,N_10059);
nor U15643 (N_15643,N_14533,N_13715);
xor U15644 (N_15644,N_14738,N_14852);
nor U15645 (N_15645,N_11738,N_13675);
nand U15646 (N_15646,N_13440,N_14608);
and U15647 (N_15647,N_14158,N_14735);
xor U15648 (N_15648,N_11062,N_11039);
or U15649 (N_15649,N_12434,N_12189);
nor U15650 (N_15650,N_11417,N_10379);
or U15651 (N_15651,N_10846,N_14405);
or U15652 (N_15652,N_11636,N_10616);
nand U15653 (N_15653,N_10415,N_11976);
xor U15654 (N_15654,N_10882,N_10825);
nand U15655 (N_15655,N_11034,N_11624);
nand U15656 (N_15656,N_14879,N_10951);
xor U15657 (N_15657,N_12691,N_12841);
nor U15658 (N_15658,N_14250,N_12019);
xnor U15659 (N_15659,N_12859,N_11074);
nand U15660 (N_15660,N_10273,N_12021);
or U15661 (N_15661,N_10560,N_11241);
xor U15662 (N_15662,N_13162,N_10191);
or U15663 (N_15663,N_14241,N_12580);
nand U15664 (N_15664,N_10459,N_11754);
nand U15665 (N_15665,N_12942,N_14858);
or U15666 (N_15666,N_12456,N_12788);
nor U15667 (N_15667,N_10948,N_11150);
nand U15668 (N_15668,N_12643,N_14458);
nand U15669 (N_15669,N_11203,N_11745);
or U15670 (N_15670,N_14662,N_11183);
or U15671 (N_15671,N_10889,N_11189);
and U15672 (N_15672,N_13293,N_10971);
or U15673 (N_15673,N_10529,N_10615);
nand U15674 (N_15674,N_12230,N_12153);
or U15675 (N_15675,N_11404,N_12445);
nor U15676 (N_15676,N_12858,N_11194);
or U15677 (N_15677,N_10590,N_14300);
nand U15678 (N_15678,N_13679,N_14666);
or U15679 (N_15679,N_12629,N_13368);
or U15680 (N_15680,N_13898,N_13899);
xnor U15681 (N_15681,N_10505,N_13541);
nand U15682 (N_15682,N_14919,N_11643);
nand U15683 (N_15683,N_10929,N_11100);
nand U15684 (N_15684,N_14079,N_14331);
nor U15685 (N_15685,N_14536,N_13412);
nand U15686 (N_15686,N_10113,N_12438);
xor U15687 (N_15687,N_11870,N_13512);
xor U15688 (N_15688,N_14604,N_11850);
xnor U15689 (N_15689,N_12084,N_14965);
nand U15690 (N_15690,N_14972,N_12396);
or U15691 (N_15691,N_10987,N_13056);
and U15692 (N_15692,N_13235,N_14957);
nor U15693 (N_15693,N_14758,N_11910);
nor U15694 (N_15694,N_12719,N_14111);
nand U15695 (N_15695,N_13437,N_10282);
and U15696 (N_15696,N_14691,N_10574);
or U15697 (N_15697,N_13069,N_14025);
nor U15698 (N_15698,N_11282,N_12711);
and U15699 (N_15699,N_10876,N_12589);
nand U15700 (N_15700,N_10629,N_12482);
nor U15701 (N_15701,N_11978,N_14785);
or U15702 (N_15702,N_12172,N_10194);
and U15703 (N_15703,N_13896,N_13803);
and U15704 (N_15704,N_11777,N_14952);
or U15705 (N_15705,N_12955,N_13398);
nor U15706 (N_15706,N_10373,N_10375);
xnor U15707 (N_15707,N_12192,N_10412);
and U15708 (N_15708,N_12205,N_10750);
or U15709 (N_15709,N_10957,N_13552);
or U15710 (N_15710,N_13582,N_10656);
or U15711 (N_15711,N_10318,N_14731);
xor U15712 (N_15712,N_13662,N_14994);
or U15713 (N_15713,N_13279,N_11532);
or U15714 (N_15714,N_14797,N_13875);
xor U15715 (N_15715,N_12611,N_12035);
and U15716 (N_15716,N_14658,N_11930);
nor U15717 (N_15717,N_11639,N_12877);
nor U15718 (N_15718,N_13308,N_11227);
nand U15719 (N_15719,N_11343,N_13831);
nand U15720 (N_15720,N_13315,N_12881);
xor U15721 (N_15721,N_10838,N_13003);
and U15722 (N_15722,N_10710,N_12432);
nand U15723 (N_15723,N_10980,N_12707);
xnor U15724 (N_15724,N_11086,N_14274);
nand U15725 (N_15725,N_11863,N_14748);
or U15726 (N_15726,N_10856,N_11428);
nor U15727 (N_15727,N_13110,N_12448);
and U15728 (N_15728,N_11096,N_12770);
xor U15729 (N_15729,N_13561,N_11866);
nand U15730 (N_15730,N_11915,N_10345);
or U15731 (N_15731,N_10367,N_14861);
or U15732 (N_15732,N_13532,N_14546);
or U15733 (N_15733,N_11840,N_12137);
or U15734 (N_15734,N_11991,N_13881);
nor U15735 (N_15735,N_12832,N_12624);
and U15736 (N_15736,N_12613,N_10439);
nand U15737 (N_15737,N_11445,N_10072);
xnor U15738 (N_15738,N_11079,N_14344);
and U15739 (N_15739,N_13025,N_12461);
and U15740 (N_15740,N_12299,N_14814);
or U15741 (N_15741,N_10998,N_14945);
and U15742 (N_15742,N_13452,N_12160);
nand U15743 (N_15743,N_10683,N_13097);
and U15744 (N_15744,N_11644,N_13865);
or U15745 (N_15745,N_14120,N_14947);
or U15746 (N_15746,N_11206,N_14831);
nor U15747 (N_15747,N_11369,N_14228);
and U15748 (N_15748,N_10944,N_14257);
nand U15749 (N_15749,N_12081,N_13711);
nor U15750 (N_15750,N_11699,N_14479);
nand U15751 (N_15751,N_10203,N_10135);
nand U15752 (N_15752,N_11138,N_10508);
nor U15753 (N_15753,N_13445,N_11002);
nand U15754 (N_15754,N_14433,N_10075);
xor U15755 (N_15755,N_13941,N_13455);
nand U15756 (N_15756,N_13957,N_12491);
xnor U15757 (N_15757,N_10283,N_14342);
xnor U15758 (N_15758,N_11125,N_11505);
nor U15759 (N_15759,N_13274,N_12266);
xnor U15760 (N_15760,N_11128,N_14460);
nor U15761 (N_15761,N_13314,N_11792);
or U15762 (N_15762,N_11452,N_12455);
and U15763 (N_15763,N_11453,N_11069);
nor U15764 (N_15764,N_10265,N_12185);
xor U15765 (N_15765,N_10923,N_13794);
and U15766 (N_15766,N_10486,N_13946);
nor U15767 (N_15767,N_12565,N_13266);
or U15768 (N_15768,N_12499,N_11704);
and U15769 (N_15769,N_12757,N_10622);
or U15770 (N_15770,N_10991,N_14172);
or U15771 (N_15771,N_14877,N_10236);
and U15772 (N_15772,N_14004,N_12469);
nor U15773 (N_15773,N_10694,N_12384);
nand U15774 (N_15774,N_13800,N_14140);
and U15775 (N_15775,N_14100,N_13224);
xnor U15776 (N_15776,N_11742,N_11844);
nand U15777 (N_15777,N_12061,N_14845);
nor U15778 (N_15778,N_10136,N_11667);
nand U15779 (N_15779,N_11876,N_13053);
and U15780 (N_15780,N_10148,N_10274);
and U15781 (N_15781,N_11625,N_12072);
xor U15782 (N_15782,N_12423,N_13795);
and U15783 (N_15783,N_14673,N_11152);
and U15784 (N_15784,N_10621,N_14341);
xnor U15785 (N_15785,N_14931,N_14709);
and U15786 (N_15786,N_10911,N_13037);
nand U15787 (N_15787,N_12554,N_14454);
nand U15788 (N_15788,N_10759,N_12257);
or U15789 (N_15789,N_11273,N_12493);
and U15790 (N_15790,N_14161,N_13366);
nor U15791 (N_15791,N_14564,N_14295);
and U15792 (N_15792,N_13617,N_10920);
nor U15793 (N_15793,N_10469,N_12010);
nor U15794 (N_15794,N_13813,N_12492);
or U15795 (N_15795,N_11357,N_12358);
xnor U15796 (N_15796,N_13599,N_12536);
or U15797 (N_15797,N_14554,N_14488);
nor U15798 (N_15798,N_12039,N_14776);
nor U15799 (N_15799,N_10748,N_12885);
xor U15800 (N_15800,N_11618,N_10725);
nor U15801 (N_15801,N_12489,N_11951);
nor U15802 (N_15802,N_11209,N_10051);
or U15803 (N_15803,N_14216,N_11292);
xnor U15804 (N_15804,N_10015,N_14330);
or U15805 (N_15805,N_11537,N_14078);
and U15806 (N_15806,N_10816,N_10057);
nand U15807 (N_15807,N_12085,N_12591);
nor U15808 (N_15808,N_11496,N_10454);
nor U15809 (N_15809,N_14514,N_12582);
nor U15810 (N_15810,N_10219,N_10611);
nor U15811 (N_15811,N_12462,N_11865);
nand U15812 (N_15812,N_14317,N_13510);
or U15813 (N_15813,N_12260,N_10131);
and U15814 (N_15814,N_12633,N_13431);
nand U15815 (N_15815,N_14381,N_10400);
xor U15816 (N_15816,N_11005,N_11311);
or U15817 (N_15817,N_13397,N_13059);
and U15818 (N_15818,N_11488,N_11299);
or U15819 (N_15819,N_13140,N_11401);
nand U15820 (N_15820,N_14487,N_11318);
nor U15821 (N_15821,N_12737,N_14513);
xnor U15822 (N_15822,N_12866,N_10007);
and U15823 (N_15823,N_10179,N_14180);
nor U15824 (N_15824,N_10672,N_11798);
and U15825 (N_15825,N_11326,N_11810);
or U15826 (N_15826,N_12428,N_11822);
xnor U15827 (N_15827,N_11545,N_10153);
nand U15828 (N_15828,N_13057,N_13710);
nor U15829 (N_15829,N_11156,N_13181);
and U15830 (N_15830,N_10183,N_10637);
nand U15831 (N_15831,N_11682,N_11716);
or U15832 (N_15832,N_12558,N_14906);
xor U15833 (N_15833,N_13031,N_11509);
nand U15834 (N_15834,N_11950,N_10867);
or U15835 (N_15835,N_12848,N_11588);
and U15836 (N_15836,N_12330,N_13066);
and U15837 (N_15837,N_14243,N_14799);
xnor U15838 (N_15838,N_11734,N_11265);
nand U15839 (N_15839,N_13045,N_14419);
xnor U15840 (N_15840,N_12779,N_12886);
nor U15841 (N_15841,N_13492,N_12731);
and U15842 (N_15842,N_14168,N_13533);
and U15843 (N_15843,N_14637,N_12958);
nor U15844 (N_15844,N_10204,N_12756);
or U15845 (N_15845,N_13014,N_14859);
nand U15846 (N_15846,N_10092,N_13449);
and U15847 (N_15847,N_10466,N_14235);
and U15848 (N_15848,N_12346,N_11108);
nor U15849 (N_15849,N_12680,N_11407);
xor U15850 (N_15850,N_14280,N_13534);
xor U15851 (N_15851,N_11648,N_13071);
nor U15852 (N_15852,N_14064,N_11269);
and U15853 (N_15853,N_12323,N_13612);
nand U15854 (N_15854,N_10512,N_14509);
xnor U15855 (N_15855,N_11376,N_12223);
or U15856 (N_15856,N_13017,N_11342);
nand U15857 (N_15857,N_10693,N_12936);
and U15858 (N_15858,N_11737,N_13307);
nand U15859 (N_15859,N_14519,N_13809);
nand U15860 (N_15860,N_13155,N_10640);
and U15861 (N_15861,N_12501,N_12808);
and U15862 (N_15862,N_12641,N_11772);
and U15863 (N_15863,N_10313,N_12861);
nand U15864 (N_15864,N_12321,N_13421);
or U15865 (N_15865,N_14500,N_11164);
xnor U15866 (N_15866,N_11512,N_12351);
nand U15867 (N_15867,N_11372,N_11595);
nor U15868 (N_15868,N_12024,N_11860);
or U15869 (N_15869,N_11049,N_10108);
xnor U15870 (N_15870,N_12623,N_11938);
nor U15871 (N_15871,N_12903,N_10123);
or U15872 (N_15872,N_13720,N_11707);
and U15873 (N_15873,N_13372,N_13985);
and U15874 (N_15874,N_12388,N_13874);
nand U15875 (N_15875,N_13548,N_12679);
nand U15876 (N_15876,N_10437,N_11593);
and U15877 (N_15877,N_14436,N_11332);
and U15878 (N_15878,N_11911,N_13000);
xnor U15879 (N_15879,N_12687,N_11813);
nor U15880 (N_15880,N_10949,N_14596);
or U15881 (N_15881,N_10999,N_13139);
xnor U15882 (N_15882,N_13217,N_11821);
nor U15883 (N_15883,N_13920,N_10883);
nor U15884 (N_15884,N_11113,N_14725);
xnor U15885 (N_15885,N_12834,N_14285);
xor U15886 (N_15886,N_11180,N_11373);
nand U15887 (N_15887,N_13621,N_12754);
or U15888 (N_15888,N_12163,N_13653);
nand U15889 (N_15889,N_12869,N_11903);
nor U15890 (N_15890,N_10285,N_11599);
nor U15891 (N_15891,N_14817,N_13337);
nand U15892 (N_15892,N_12437,N_10631);
xor U15893 (N_15893,N_10119,N_13535);
nand U15894 (N_15894,N_10138,N_11016);
or U15895 (N_15895,N_14499,N_11829);
xnor U15896 (N_15896,N_12514,N_12682);
nand U15897 (N_15897,N_13060,N_11068);
xor U15898 (N_15898,N_11493,N_12519);
or U15899 (N_15899,N_10174,N_13905);
xnor U15900 (N_15900,N_10807,N_10355);
nor U15901 (N_15901,N_11196,N_11888);
nand U15902 (N_15902,N_14655,N_12068);
xor U15903 (N_15903,N_13515,N_13163);
and U15904 (N_15904,N_11030,N_10267);
nor U15905 (N_15905,N_13117,N_14187);
nand U15906 (N_15906,N_11752,N_12141);
xnor U15907 (N_15907,N_10111,N_11513);
and U15908 (N_15908,N_13528,N_11893);
xor U15909 (N_15909,N_13570,N_13622);
nand U15910 (N_15910,N_13281,N_14949);
nor U15911 (N_15911,N_10542,N_11695);
nor U15912 (N_15912,N_13446,N_12734);
nor U15913 (N_15913,N_11058,N_14891);
xor U15914 (N_15914,N_14146,N_11834);
xnor U15915 (N_15915,N_12075,N_12333);
or U15916 (N_15916,N_10256,N_12814);
xnor U15917 (N_15917,N_13736,N_12700);
and U15918 (N_15918,N_11054,N_13019);
nand U15919 (N_15919,N_10171,N_11928);
or U15920 (N_15920,N_10276,N_11875);
nor U15921 (N_15921,N_11187,N_13200);
and U15922 (N_15922,N_11004,N_14807);
or U15923 (N_15923,N_11899,N_11678);
xor U15924 (N_15924,N_12103,N_12452);
nor U15925 (N_15925,N_10390,N_13730);
or U15926 (N_15926,N_12352,N_14415);
or U15927 (N_15927,N_13638,N_11986);
xnor U15928 (N_15928,N_10550,N_13907);
xor U15929 (N_15929,N_10733,N_12289);
and U15930 (N_15930,N_11395,N_12529);
or U15931 (N_15931,N_13597,N_13950);
nand U15932 (N_15932,N_14314,N_11954);
nor U15933 (N_15933,N_10073,N_13869);
xnor U15934 (N_15934,N_10956,N_10461);
nand U15935 (N_15935,N_10449,N_11579);
nand U15936 (N_15936,N_14296,N_11247);
xnor U15937 (N_15937,N_12901,N_12376);
or U15938 (N_15938,N_10077,N_12348);
nor U15939 (N_15939,N_10048,N_12050);
nor U15940 (N_15940,N_10327,N_12347);
nand U15941 (N_15941,N_13328,N_13061);
nand U15942 (N_15942,N_10248,N_11499);
nor U15943 (N_15943,N_10416,N_12018);
xnor U15944 (N_15944,N_11162,N_12510);
or U15945 (N_15945,N_10478,N_14185);
and U15946 (N_15946,N_11077,N_13571);
xor U15947 (N_15947,N_10741,N_14230);
xor U15948 (N_15948,N_12426,N_10343);
and U15949 (N_15949,N_10739,N_13466);
or U15950 (N_15950,N_14640,N_10464);
and U15951 (N_15951,N_12062,N_12014);
nor U15952 (N_15952,N_11139,N_13849);
nor U15953 (N_15953,N_11564,N_14573);
xnor U15954 (N_15954,N_11561,N_14298);
and U15955 (N_15955,N_14634,N_14097);
or U15956 (N_15956,N_10796,N_11259);
xnor U15957 (N_15957,N_13172,N_11726);
and U15958 (N_15958,N_12033,N_13735);
and U15959 (N_15959,N_13560,N_11366);
and U15960 (N_15960,N_12891,N_13428);
xor U15961 (N_15961,N_12280,N_14720);
and U15962 (N_15962,N_14661,N_11571);
xnor U15963 (N_15963,N_13901,N_14522);
xor U15964 (N_15964,N_12537,N_10562);
or U15965 (N_15965,N_13230,N_14848);
or U15966 (N_15966,N_10096,N_11497);
or U15967 (N_15967,N_14382,N_13116);
nand U15968 (N_15968,N_13620,N_13779);
and U15969 (N_15969,N_13250,N_13267);
xnor U15970 (N_15970,N_14629,N_10519);
nor U15971 (N_15971,N_12409,N_12573);
nor U15972 (N_15972,N_10378,N_11486);
xnor U15973 (N_15973,N_13168,N_11800);
nand U15974 (N_15974,N_12401,N_14392);
nand U15975 (N_15975,N_13619,N_13225);
or U15976 (N_15976,N_10020,N_14865);
nand U15977 (N_15977,N_10456,N_12020);
and U15978 (N_15978,N_13193,N_10531);
xor U15979 (N_15979,N_12337,N_13536);
or U15980 (N_15980,N_11279,N_14880);
xnor U15981 (N_15981,N_12925,N_12047);
or U15982 (N_15982,N_13124,N_12945);
and U15983 (N_15983,N_11378,N_14038);
nor U15984 (N_15984,N_14616,N_10056);
nand U15985 (N_15985,N_14377,N_12071);
and U15986 (N_15986,N_11296,N_11968);
xor U15987 (N_15987,N_10603,N_14266);
or U15988 (N_15988,N_10939,N_11391);
and U15989 (N_15989,N_13564,N_14589);
nand U15990 (N_15990,N_10255,N_13238);
and U15991 (N_15991,N_13027,N_11230);
xor U15992 (N_15992,N_10054,N_11105);
nand U15993 (N_15993,N_10788,N_10235);
or U15994 (N_15994,N_10994,N_12004);
xor U15995 (N_15995,N_11997,N_13976);
or U15996 (N_15996,N_14389,N_11526);
and U15997 (N_15997,N_11149,N_10181);
xor U15998 (N_15998,N_13953,N_12650);
or U15999 (N_15999,N_12785,N_14641);
or U16000 (N_16000,N_12304,N_13295);
xnor U16001 (N_16001,N_11485,N_13008);
or U16002 (N_16002,N_13979,N_13423);
xor U16003 (N_16003,N_10857,N_10877);
nand U16004 (N_16004,N_11520,N_10046);
nand U16005 (N_16005,N_10730,N_12142);
xor U16006 (N_16006,N_13740,N_12826);
and U16007 (N_16007,N_13106,N_14139);
and U16008 (N_16008,N_11188,N_11170);
nand U16009 (N_16009,N_13278,N_14121);
or U16010 (N_16010,N_10182,N_14680);
and U16011 (N_16011,N_13453,N_11130);
and U16012 (N_16012,N_13062,N_13298);
nand U16013 (N_16013,N_11325,N_11381);
or U16014 (N_16014,N_12385,N_14600);
and U16015 (N_16015,N_13889,N_12735);
or U16016 (N_16016,N_13820,N_13944);
or U16017 (N_16017,N_13165,N_13304);
and U16018 (N_16018,N_12639,N_14951);
nand U16019 (N_16019,N_12640,N_13433);
or U16020 (N_16020,N_12603,N_13426);
or U16021 (N_16021,N_10841,N_10399);
nor U16022 (N_16022,N_13789,N_10533);
nand U16023 (N_16023,N_14477,N_10424);
xnor U16024 (N_16024,N_13556,N_13126);
nor U16025 (N_16025,N_11652,N_10628);
xnor U16026 (N_16026,N_11642,N_14475);
nand U16027 (N_16027,N_12345,N_14885);
nor U16028 (N_16028,N_11441,N_14752);
and U16029 (N_16029,N_12366,N_11898);
xnor U16030 (N_16030,N_10352,N_13677);
or U16031 (N_16031,N_14526,N_14924);
nand U16032 (N_16032,N_10332,N_12315);
or U16033 (N_16033,N_14821,N_13939);
xnor U16034 (N_16034,N_10602,N_13539);
nor U16035 (N_16035,N_14150,N_10083);
xor U16036 (N_16036,N_10310,N_14766);
xnor U16037 (N_16037,N_10870,N_12723);
xor U16038 (N_16038,N_11514,N_14804);
nor U16039 (N_16039,N_11733,N_10691);
or U16040 (N_16040,N_12410,N_14067);
and U16041 (N_16041,N_13589,N_12458);
xor U16042 (N_16042,N_11245,N_10701);
or U16043 (N_16043,N_14036,N_14447);
nor U16044 (N_16044,N_14823,N_11334);
nand U16045 (N_16045,N_10860,N_11586);
nor U16046 (N_16046,N_14122,N_12392);
nor U16047 (N_16047,N_14606,N_14937);
or U16048 (N_16048,N_10407,N_12575);
nand U16049 (N_16049,N_12386,N_11980);
and U16050 (N_16050,N_10580,N_11653);
xnor U16051 (N_16051,N_14559,N_11641);
xnor U16052 (N_16052,N_12851,N_12471);
nor U16053 (N_16053,N_14926,N_11879);
or U16054 (N_16054,N_10275,N_10226);
nand U16055 (N_16055,N_14694,N_10160);
or U16056 (N_16056,N_13531,N_12803);
nand U16057 (N_16057,N_14843,N_13668);
or U16058 (N_16058,N_14229,N_14472);
nand U16059 (N_16059,N_13783,N_13297);
and U16060 (N_16060,N_12060,N_14188);
or U16061 (N_16061,N_10347,N_12653);
nand U16062 (N_16062,N_10575,N_14151);
nor U16063 (N_16063,N_12634,N_10488);
or U16064 (N_16064,N_12435,N_14403);
nand U16065 (N_16065,N_13508,N_11234);
nand U16066 (N_16066,N_13299,N_12543);
nand U16067 (N_16067,N_12520,N_11276);
nor U16068 (N_16068,N_12279,N_12621);
nor U16069 (N_16069,N_14059,N_10593);
or U16070 (N_16070,N_10676,N_13130);
xnor U16071 (N_16071,N_12569,N_14798);
nor U16072 (N_16072,N_12806,N_13797);
and U16073 (N_16073,N_10175,N_10592);
or U16074 (N_16074,N_14029,N_14609);
or U16075 (N_16075,N_14761,N_10494);
and U16076 (N_16076,N_11836,N_11884);
nand U16077 (N_16077,N_14449,N_10953);
nand U16078 (N_16078,N_10544,N_10306);
or U16079 (N_16079,N_14897,N_13669);
or U16080 (N_16080,N_11563,N_13006);
and U16081 (N_16081,N_12996,N_14104);
nor U16082 (N_16082,N_10128,N_14207);
or U16083 (N_16083,N_11882,N_12561);
or U16084 (N_16084,N_12158,N_14311);
nand U16085 (N_16085,N_13255,N_10742);
nand U16086 (N_16086,N_10895,N_10309);
or U16087 (N_16087,N_13925,N_11143);
and U16088 (N_16088,N_10094,N_10081);
nor U16089 (N_16089,N_10808,N_12609);
and U16090 (N_16090,N_10293,N_11536);
xor U16091 (N_16091,N_10782,N_11137);
nand U16092 (N_16092,N_12801,N_11466);
xor U16093 (N_16093,N_12525,N_10385);
nor U16094 (N_16094,N_13218,N_14301);
nand U16095 (N_16095,N_14327,N_10432);
xor U16096 (N_16096,N_11287,N_13690);
and U16097 (N_16097,N_12842,N_10747);
nand U16098 (N_16098,N_13573,N_13773);
xor U16099 (N_16099,N_14910,N_11531);
or U16100 (N_16100,N_10982,N_13563);
or U16101 (N_16101,N_12283,N_12670);
nor U16102 (N_16102,N_11926,N_13087);
xnor U16103 (N_16103,N_14446,N_13262);
or U16104 (N_16104,N_13493,N_13133);
nand U16105 (N_16105,N_14329,N_11237);
or U16106 (N_16106,N_10406,N_14719);
or U16107 (N_16107,N_14595,N_12937);
nor U16108 (N_16108,N_13882,N_10380);
and U16109 (N_16109,N_14176,N_10401);
nor U16110 (N_16110,N_10538,N_11778);
nand U16111 (N_16111,N_13416,N_10858);
nor U16112 (N_16112,N_12357,N_11963);
nor U16113 (N_16113,N_13167,N_11312);
nand U16114 (N_16114,N_10680,N_13918);
nor U16115 (N_16115,N_10779,N_11959);
or U16116 (N_16116,N_11254,N_13382);
xnor U16117 (N_16117,N_14729,N_10101);
nor U16118 (N_16118,N_12303,N_14925);
nor U16119 (N_16119,N_12460,N_10036);
nand U16120 (N_16120,N_11826,N_12943);
xnor U16121 (N_16121,N_10685,N_13732);
nand U16122 (N_16122,N_13833,N_13926);
nand U16123 (N_16123,N_14269,N_11685);
and U16124 (N_16124,N_12115,N_12587);
nor U16125 (N_16125,N_11556,N_11632);
xnor U16126 (N_16126,N_11612,N_13914);
and U16127 (N_16127,N_13693,N_14982);
and U16128 (N_16128,N_12157,N_13991);
and U16129 (N_16129,N_11281,N_12991);
nand U16130 (N_16130,N_10709,N_14757);
or U16131 (N_16131,N_14410,N_10600);
and U16132 (N_16132,N_14443,N_11387);
and U16133 (N_16133,N_11805,N_14601);
xor U16134 (N_16134,N_12132,N_13613);
nor U16135 (N_16135,N_13296,N_14114);
nor U16136 (N_16136,N_12576,N_14835);
and U16137 (N_16137,N_11145,N_14459);
xnor U16138 (N_16138,N_14325,N_12989);
and U16139 (N_16139,N_14740,N_13569);
and U16140 (N_16140,N_12186,N_11775);
or U16141 (N_16141,N_11331,N_12889);
nor U16142 (N_16142,N_10308,N_13090);
nand U16143 (N_16143,N_13734,N_12846);
or U16144 (N_16144,N_13223,N_14660);
and U16145 (N_16145,N_11592,N_13527);
nor U16146 (N_16146,N_14464,N_14670);
xnor U16147 (N_16147,N_10475,N_11457);
or U16148 (N_16148,N_12988,N_14019);
and U16149 (N_16149,N_13791,N_10220);
xor U16150 (N_16150,N_14688,N_11931);
xnor U16151 (N_16151,N_12331,N_14530);
or U16152 (N_16152,N_10159,N_14239);
and U16153 (N_16153,N_11205,N_14441);
and U16154 (N_16154,N_12483,N_11622);
or U16155 (N_16155,N_10655,N_12472);
or U16156 (N_16156,N_13936,N_11436);
nand U16157 (N_16157,N_10704,N_13369);
xnor U16158 (N_16158,N_13503,N_11289);
or U16159 (N_16159,N_12857,N_12764);
nor U16160 (N_16160,N_14022,N_12540);
or U16161 (N_16161,N_10943,N_13798);
and U16162 (N_16162,N_13649,N_10223);
xnor U16163 (N_16163,N_13784,N_11294);
nor U16164 (N_16164,N_11479,N_13853);
nor U16165 (N_16165,N_11921,N_12373);
or U16166 (N_16166,N_14651,N_10052);
or U16167 (N_16167,N_14793,N_10244);
xor U16168 (N_16168,N_10068,N_10259);
xnor U16169 (N_16169,N_13209,N_10032);
and U16170 (N_16170,N_11355,N_10197);
nand U16171 (N_16171,N_13688,N_13754);
xnor U16172 (N_16172,N_14092,N_12356);
nand U16173 (N_16173,N_13830,N_13870);
or U16174 (N_16174,N_14099,N_11521);
xor U16175 (N_16175,N_14696,N_12725);
nor U16176 (N_16176,N_13729,N_10572);
nor U16177 (N_16177,N_10487,N_13208);
nor U16178 (N_16178,N_12894,N_11437);
xor U16179 (N_16179,N_11615,N_12329);
or U16180 (N_16180,N_10890,N_11819);
and U16181 (N_16181,N_14872,N_12926);
nor U16182 (N_16182,N_12981,N_14461);
nor U16183 (N_16183,N_12802,N_11897);
xor U16184 (N_16184,N_12840,N_12505);
and U16185 (N_16185,N_10623,N_13468);
and U16186 (N_16186,N_14261,N_11825);
and U16187 (N_16187,N_12495,N_14125);
nor U16188 (N_16188,N_14268,N_10403);
nand U16189 (N_16189,N_12485,N_12233);
or U16190 (N_16190,N_12058,N_11354);
or U16191 (N_16191,N_11669,N_11060);
nor U16192 (N_16192,N_12503,N_12098);
xnor U16193 (N_16193,N_11567,N_13120);
xnor U16194 (N_16194,N_14234,N_13393);
and U16195 (N_16195,N_11244,N_11795);
nor U16196 (N_16196,N_12393,N_11168);
xor U16197 (N_16197,N_11696,N_11310);
xor U16198 (N_16198,N_10502,N_12631);
nand U16199 (N_16199,N_11539,N_12023);
xor U16200 (N_16200,N_14463,N_13667);
xor U16201 (N_16201,N_13151,N_11027);
nand U16202 (N_16202,N_14306,N_14043);
and U16203 (N_16203,N_13496,N_13125);
nor U16204 (N_16204,N_11889,N_11213);
nand U16205 (N_16205,N_11423,N_14556);
nor U16206 (N_16206,N_13680,N_14066);
nand U16207 (N_16207,N_13064,N_10063);
nor U16208 (N_16208,N_12638,N_11444);
xor U16209 (N_16209,N_10979,N_13547);
or U16210 (N_16210,N_12690,N_10567);
or U16211 (N_16211,N_14539,N_10277);
nor U16212 (N_16212,N_14340,N_10232);
xor U16213 (N_16213,N_11224,N_14820);
nor U16214 (N_16214,N_13386,N_13962);
and U16215 (N_16215,N_10086,N_11507);
nor U16216 (N_16216,N_11802,N_12100);
or U16217 (N_16217,N_11094,N_11197);
nor U16218 (N_16218,N_11602,N_10252);
xnor U16219 (N_16219,N_12117,N_13318);
or U16220 (N_16220,N_14014,N_11965);
xor U16221 (N_16221,N_10064,N_14749);
or U16222 (N_16222,N_13112,N_13227);
or U16223 (N_16223,N_10333,N_11422);
or U16224 (N_16224,N_10632,N_13965);
nand U16225 (N_16225,N_11134,N_11972);
nor U16226 (N_16226,N_13883,N_14789);
and U16227 (N_16227,N_10792,N_13419);
or U16228 (N_16228,N_14723,N_13655);
or U16229 (N_16229,N_10227,N_10231);
nand U16230 (N_16230,N_14940,N_12585);
or U16231 (N_16231,N_10610,N_13644);
xnor U16232 (N_16232,N_12122,N_13682);
nand U16233 (N_16233,N_11459,N_11400);
and U16234 (N_16234,N_11014,N_11408);
or U16235 (N_16235,N_11235,N_13253);
nor U16236 (N_16236,N_12507,N_14561);
nand U16237 (N_16237,N_13435,N_10029);
or U16238 (N_16238,N_11585,N_11116);
xnor U16239 (N_16239,N_13498,N_12067);
or U16240 (N_16240,N_10854,N_14495);
nor U16241 (N_16241,N_11719,N_11231);
xnor U16242 (N_16242,N_14171,N_10800);
or U16243 (N_16243,N_12915,N_10296);
nor U16244 (N_16244,N_11604,N_12897);
xor U16245 (N_16245,N_12709,N_12034);
and U16246 (N_16246,N_11905,N_10088);
or U16247 (N_16247,N_10861,N_11705);
nor U16248 (N_16248,N_10869,N_13378);
nand U16249 (N_16249,N_11856,N_13129);
nand U16250 (N_16250,N_12683,N_13289);
nand U16251 (N_16251,N_11655,N_11842);
nor U16252 (N_16252,N_12267,N_12457);
and U16253 (N_16253,N_14364,N_12517);
xor U16254 (N_16254,N_11198,N_14055);
or U16255 (N_16255,N_13258,N_11962);
or U16256 (N_16256,N_11973,N_12660);
and U16257 (N_16257,N_14506,N_11420);
nor U16258 (N_16258,N_14086,N_14746);
xor U16259 (N_16259,N_12154,N_14432);
nor U16260 (N_16260,N_10124,N_11090);
nor U16261 (N_16261,N_12265,N_12953);
nand U16262 (N_16262,N_11945,N_14685);
xnor U16263 (N_16263,N_11491,N_10727);
nor U16264 (N_16264,N_12225,N_11415);
or U16265 (N_16265,N_13241,N_12950);
or U16266 (N_16266,N_12839,N_11255);
xor U16267 (N_16267,N_10154,N_11739);
nor U16268 (N_16268,N_12553,N_11553);
nor U16269 (N_16269,N_14769,N_14154);
and U16270 (N_16270,N_13565,N_14612);
and U16271 (N_16271,N_10977,N_12429);
nand U16272 (N_16272,N_12688,N_10660);
or U16273 (N_16273,N_14837,N_12932);
or U16274 (N_16274,N_13360,N_12191);
xor U16275 (N_16275,N_11833,N_14137);
nor U16276 (N_16276,N_12636,N_14467);
and U16277 (N_16277,N_11791,N_13367);
nor U16278 (N_16278,N_12007,N_11598);
and U16279 (N_16279,N_11044,N_14144);
or U16280 (N_16280,N_13942,N_12112);
nand U16281 (N_16281,N_13650,N_11904);
and U16282 (N_16282,N_10142,N_14221);
xor U16283 (N_16283,N_10961,N_10211);
xor U16284 (N_16284,N_11728,N_13311);
or U16285 (N_16285,N_14979,N_13331);
xnor U16286 (N_16286,N_11661,N_12420);
nor U16287 (N_16287,N_14212,N_12203);
xnor U16288 (N_16288,N_14473,N_10192);
xnor U16289 (N_16289,N_11691,N_10837);
and U16290 (N_16290,N_13792,N_13810);
or U16291 (N_16291,N_10613,N_14901);
and U16292 (N_16292,N_14470,N_13877);
and U16293 (N_16293,N_12246,N_11000);
nor U16294 (N_16294,N_11748,N_11664);
and U16295 (N_16295,N_13376,N_13495);
and U16296 (N_16296,N_14355,N_10446);
or U16297 (N_16297,N_13660,N_10176);
or U16298 (N_16298,N_11686,N_14915);
and U16299 (N_16299,N_11804,N_13641);
nand U16300 (N_16300,N_10323,N_14876);
and U16301 (N_16301,N_13118,N_10199);
or U16302 (N_16302,N_13320,N_10288);
nand U16303 (N_16303,N_13389,N_10152);
nand U16304 (N_16304,N_13194,N_11022);
or U16305 (N_16305,N_10433,N_14855);
xnor U16306 (N_16306,N_10125,N_10578);
nand U16307 (N_16307,N_14324,N_14012);
or U16308 (N_16308,N_10738,N_10706);
and U16309 (N_16309,N_13763,N_10990);
or U16310 (N_16310,N_12086,N_10398);
and U16311 (N_16311,N_14365,N_13575);
xor U16312 (N_16312,N_12059,N_13811);
or U16313 (N_16313,N_10444,N_12933);
xor U16314 (N_16314,N_11173,N_11474);
nand U16315 (N_16315,N_11708,N_10824);
or U16316 (N_16316,N_12678,N_12383);
or U16317 (N_16317,N_13164,N_14404);
nand U16318 (N_16318,N_13245,N_11216);
and U16319 (N_16319,N_12983,N_13306);
and U16320 (N_16320,N_14718,N_12397);
or U16321 (N_16321,N_13065,N_13911);
xor U16322 (N_16322,N_14060,N_14409);
or U16323 (N_16323,N_12733,N_14883);
nor U16324 (N_16324,N_14319,N_11475);
nand U16325 (N_16325,N_13568,N_10916);
xor U16326 (N_16326,N_13746,N_10713);
xor U16327 (N_16327,N_14898,N_14948);
nor U16328 (N_16328,N_13745,N_14448);
nor U16329 (N_16329,N_14849,N_11665);
xor U16330 (N_16330,N_12896,N_11402);
xnor U16331 (N_16331,N_14482,N_10501);
or U16332 (N_16332,N_10420,N_11427);
or U16333 (N_16333,N_14866,N_14088);
and U16334 (N_16334,N_13960,N_10479);
or U16335 (N_16335,N_13402,N_10155);
xor U16336 (N_16336,N_13502,N_10405);
nand U16337 (N_16337,N_10209,N_12544);
and U16338 (N_16338,N_12535,N_10582);
or U16339 (N_16339,N_14548,N_11580);
and U16340 (N_16340,N_14610,N_10819);
and U16341 (N_16341,N_13523,N_11646);
or U16342 (N_16342,N_14543,N_14023);
nand U16343 (N_16343,N_13685,N_11478);
nand U16344 (N_16344,N_12867,N_14024);
nand U16345 (N_16345,N_10509,N_11469);
and U16346 (N_16346,N_11341,N_14279);
xnor U16347 (N_16347,N_13406,N_11021);
nand U16348 (N_16348,N_12956,N_12911);
xor U16349 (N_16349,N_10555,N_10474);
nand U16350 (N_16350,N_12751,N_14096);
nor U16351 (N_16351,N_13290,N_14934);
nor U16352 (N_16352,N_14420,N_10044);
or U16353 (N_16353,N_11414,N_14366);
nand U16354 (N_16354,N_10028,N_12545);
xor U16355 (N_16355,N_13157,N_11489);
or U16356 (N_16356,N_13545,N_12716);
xnor U16357 (N_16357,N_10726,N_11403);
and U16358 (N_16358,N_10893,N_12403);
nor U16359 (N_16359,N_10751,N_12288);
or U16360 (N_16360,N_14093,N_14762);
and U16361 (N_16361,N_11161,N_13764);
and U16362 (N_16362,N_10126,N_13259);
and U16363 (N_16363,N_11438,N_14504);
nand U16364 (N_16364,N_12977,N_11610);
or U16365 (N_16365,N_13554,N_11295);
and U16366 (N_16366,N_10431,N_14195);
or U16367 (N_16367,N_10888,N_11370);
or U16368 (N_16368,N_10909,N_11464);
and U16369 (N_16369,N_13731,N_10360);
nor U16370 (N_16370,N_10818,N_12398);
xor U16371 (N_16371,N_12548,N_14683);
nand U16372 (N_16372,N_10331,N_14676);
nor U16373 (N_16373,N_12313,N_14650);
and U16374 (N_16374,N_10321,N_10839);
nand U16375 (N_16375,N_12767,N_11172);
nor U16376 (N_16376,N_13443,N_14535);
nand U16377 (N_16377,N_12065,N_10880);
xor U16378 (N_16378,N_14283,N_11758);
nor U16379 (N_16379,N_14759,N_14391);
or U16380 (N_16380,N_11053,N_12306);
nor U16381 (N_16381,N_12644,N_10115);
or U16382 (N_16382,N_10917,N_11939);
or U16383 (N_16383,N_11147,N_10524);
xnor U16384 (N_16384,N_10566,N_14015);
or U16385 (N_16385,N_14968,N_10526);
nand U16386 (N_16386,N_13837,N_11190);
nand U16387 (N_16387,N_12560,N_12982);
and U16388 (N_16388,N_10591,N_14011);
and U16389 (N_16389,N_10185,N_11111);
xor U16390 (N_16390,N_12984,N_13189);
and U16391 (N_16391,N_12800,N_11755);
xnor U16392 (N_16392,N_12628,N_12701);
and U16393 (N_16393,N_10237,N_14540);
nor U16394 (N_16394,N_14950,N_13576);
and U16395 (N_16395,N_12831,N_13766);
or U16396 (N_16396,N_10156,N_13969);
xnor U16397 (N_16397,N_10551,N_14018);
or U16398 (N_16398,N_12844,N_14567);
nor U16399 (N_16399,N_12102,N_10534);
nor U16400 (N_16400,N_12450,N_14181);
nor U16401 (N_16401,N_14245,N_13007);
nor U16402 (N_16402,N_11654,N_10499);
nand U16403 (N_16403,N_13785,N_10584);
or U16404 (N_16404,N_11570,N_14455);
nor U16405 (N_16405,N_14031,N_10952);
or U16406 (N_16406,N_14288,N_10587);
or U16407 (N_16407,N_12220,N_11744);
or U16408 (N_16408,N_12776,N_12656);
nand U16409 (N_16409,N_14006,N_12563);
nand U16410 (N_16410,N_13959,N_14862);
nand U16411 (N_16411,N_11504,N_10297);
xor U16412 (N_16412,N_13843,N_11251);
xor U16413 (N_16413,N_14959,N_13776);
nor U16414 (N_16414,N_13409,N_14993);
nor U16415 (N_16415,N_10896,N_11853);
or U16416 (N_16416,N_11995,N_11828);
xnor U16417 (N_16417,N_11789,N_12527);
nand U16418 (N_16418,N_11083,N_14491);
nor U16419 (N_16419,N_11547,N_14886);
or U16420 (N_16420,N_14549,N_11093);
xnor U16421 (N_16421,N_14602,N_11330);
nand U16422 (N_16422,N_14095,N_10810);
xnor U16423 (N_16423,N_12193,N_10348);
nand U16424 (N_16424,N_10497,N_12780);
nor U16425 (N_16425,N_13229,N_10903);
nand U16426 (N_16426,N_12677,N_10541);
xor U16427 (N_16427,N_14570,N_13408);
or U16428 (N_16428,N_11788,N_12562);
or U16429 (N_16429,N_12159,N_14109);
and U16430 (N_16430,N_13451,N_11538);
xnor U16431 (N_16431,N_12960,N_11872);
nor U16432 (N_16432,N_10576,N_14864);
or U16433 (N_16433,N_12574,N_13354);
nand U16434 (N_16434,N_10908,N_12632);
or U16435 (N_16435,N_14727,N_14343);
xor U16436 (N_16436,N_11117,N_14328);
or U16437 (N_16437,N_14320,N_12534);
nor U16438 (N_16438,N_10834,N_14863);
and U16439 (N_16439,N_12120,N_11151);
and U16440 (N_16440,N_13154,N_13526);
nor U16441 (N_16441,N_10344,N_14294);
nor U16442 (N_16442,N_14778,N_11316);
and U16443 (N_16443,N_12091,N_11012);
nand U16444 (N_16444,N_11363,N_11202);
nand U16445 (N_16445,N_14819,N_10830);
and U16446 (N_16446,N_10753,N_12865);
xnor U16447 (N_16447,N_13790,N_10976);
xnor U16448 (N_16448,N_13625,N_14130);
xor U16449 (N_16449,N_10978,N_11351);
and U16450 (N_16450,N_10732,N_11109);
nor U16451 (N_16451,N_14041,N_13963);
or U16452 (N_16452,N_13956,N_10228);
xor U16453 (N_16453,N_11638,N_14544);
xor U16454 (N_16454,N_14369,N_13590);
or U16455 (N_16455,N_12793,N_13156);
and U16456 (N_16456,N_12586,N_13047);
or U16457 (N_16457,N_12695,N_10539);
nand U16458 (N_16458,N_10764,N_13188);
nand U16459 (N_16459,N_13859,N_10761);
xnor U16460 (N_16460,N_13915,N_12262);
or U16461 (N_16461,N_14987,N_10442);
nand U16462 (N_16462,N_10695,N_10708);
or U16463 (N_16463,N_10184,N_10312);
xnor U16464 (N_16464,N_10066,N_12856);
or U16465 (N_16465,N_11680,N_14875);
xnor U16466 (N_16466,N_12645,N_11040);
and U16467 (N_16467,N_11481,N_13520);
and U16468 (N_16468,N_13460,N_13141);
and U16469 (N_16469,N_12533,N_12854);
or U16470 (N_16470,N_12190,N_10268);
nand U16471 (N_16471,N_11816,N_14874);
xor U16472 (N_16472,N_11929,N_10716);
nor U16473 (N_16473,N_11763,N_12176);
and U16474 (N_16474,N_10515,N_14476);
or U16475 (N_16475,N_10330,N_10690);
and U16476 (N_16476,N_10522,N_12113);
and U16477 (N_16477,N_12837,N_14039);
or U16478 (N_16478,N_12813,N_14380);
nand U16479 (N_16479,N_12444,N_14483);
xor U16480 (N_16480,N_11454,N_14017);
nor U16481 (N_16481,N_12905,N_12308);
xnor U16482 (N_16482,N_10892,N_14198);
or U16483 (N_16483,N_10322,N_11535);
nand U16484 (N_16484,N_11006,N_10840);
and U16485 (N_16485,N_14297,N_10178);
and U16486 (N_16486,N_14386,N_12964);
or U16487 (N_16487,N_13310,N_10583);
and U16488 (N_16488,N_13247,N_10595);
nand U16489 (N_16489,N_13067,N_10382);
nor U16490 (N_16490,N_12532,N_13348);
and U16491 (N_16491,N_13486,N_10767);
or U16492 (N_16492,N_11362,N_10850);
or U16493 (N_16493,N_14422,N_11740);
nand U16494 (N_16494,N_10828,N_11322);
nor U16495 (N_16495,N_13893,N_10881);
or U16496 (N_16496,N_13681,N_13239);
nor U16497 (N_16497,N_14227,N_14532);
xnor U16498 (N_16498,N_11596,N_12708);
nor U16499 (N_16499,N_12663,N_10688);
nand U16500 (N_16500,N_12073,N_11749);
nand U16501 (N_16501,N_13761,N_14072);
and U16502 (N_16502,N_12281,N_12761);
nand U16503 (N_16503,N_11818,N_11456);
nand U16504 (N_16504,N_11970,N_10381);
or U16505 (N_16505,N_12617,N_11729);
or U16506 (N_16506,N_11046,N_14008);
and U16507 (N_16507,N_10030,N_12931);
nand U16508 (N_16508,N_14887,N_14163);
nand U16509 (N_16509,N_13605,N_14830);
xor U16510 (N_16510,N_11530,N_13326);
nor U16511 (N_16511,N_11191,N_13429);
or U16512 (N_16512,N_11055,N_12884);
nor U16513 (N_16513,N_10107,N_14790);
and U16514 (N_16514,N_13906,N_10164);
nand U16515 (N_16515,N_13580,N_12622);
xnor U16516 (N_16516,N_11036,N_13937);
or U16517 (N_16517,N_13511,N_12408);
nor U16518 (N_16518,N_10757,N_10930);
or U16519 (N_16519,N_12836,N_13891);
or U16520 (N_16520,N_10351,N_12001);
xnor U16521 (N_16521,N_10413,N_14167);
and U16522 (N_16522,N_12017,N_11103);
nor U16523 (N_16523,N_10933,N_14040);
nor U16524 (N_16524,N_14997,N_11119);
and U16525 (N_16525,N_11064,N_12129);
or U16526 (N_16526,N_10630,N_14635);
and U16527 (N_16527,N_13020,N_14484);
nand U16528 (N_16528,N_12614,N_13330);
and U16529 (N_16529,N_11533,N_14741);
nand U16530 (N_16530,N_13032,N_10724);
and U16531 (N_16531,N_10298,N_12064);
xor U16532 (N_16532,N_14587,N_14152);
nor U16533 (N_16533,N_11384,N_14717);
and U16534 (N_16534,N_14502,N_14588);
and U16535 (N_16535,N_14736,N_11999);
nor U16536 (N_16536,N_14684,N_11495);
nor U16537 (N_16537,N_13450,N_11133);
nand U16538 (N_16538,N_14841,N_11193);
and U16539 (N_16539,N_13336,N_10141);
nand U16540 (N_16540,N_11409,N_10359);
and U16541 (N_16541,N_10371,N_10146);
or U16542 (N_16542,N_14703,N_11406);
nor U16543 (N_16543,N_13562,N_12986);
nor U16544 (N_16544,N_11666,N_14253);
and U16545 (N_16545,N_13603,N_11091);
nand U16546 (N_16546,N_14652,N_12488);
xnor U16547 (N_16547,N_11171,N_13737);
xor U16548 (N_16548,N_10912,N_10315);
or U16549 (N_16549,N_11258,N_14116);
or U16550 (N_16550,N_11268,N_12143);
or U16551 (N_16551,N_14760,N_11065);
nand U16552 (N_16552,N_11573,N_11126);
nor U16553 (N_16553,N_12307,N_14985);
and U16554 (N_16554,N_10130,N_14955);
nor U16555 (N_16555,N_11360,N_12673);
xor U16556 (N_16556,N_10071,N_14292);
xor U16557 (N_16557,N_14743,N_10498);
and U16558 (N_16558,N_14677,N_13980);
xor U16559 (N_16559,N_14938,N_14734);
nor U16560 (N_16560,N_12913,N_10470);
nor U16561 (N_16561,N_12405,N_12676);
and U16562 (N_16562,N_12340,N_13632);
nor U16563 (N_16563,N_13997,N_11037);
and U16564 (N_16564,N_10144,N_11260);
nor U16565 (N_16565,N_11712,N_10601);
and U16566 (N_16566,N_13724,N_11924);
xnor U16567 (N_16567,N_13099,N_11964);
nor U16568 (N_16568,N_11670,N_10649);
and U16569 (N_16569,N_12968,N_12011);
and U16570 (N_16570,N_14105,N_10084);
xor U16571 (N_16571,N_12255,N_13316);
xnor U16572 (N_16572,N_14231,N_11540);
xnor U16573 (N_16573,N_12182,N_14850);
and U16574 (N_16574,N_10540,N_12244);
xnor U16575 (N_16575,N_10002,N_12995);
nor U16576 (N_16576,N_13658,N_13747);
xor U16577 (N_16577,N_10762,N_13391);
nand U16578 (N_16578,N_10109,N_14309);
nand U16579 (N_16579,N_14346,N_11052);
and U16580 (N_16580,N_14889,N_12772);
or U16581 (N_16581,N_13135,N_12089);
and U16582 (N_16582,N_10033,N_10573);
and U16583 (N_16583,N_13631,N_12674);
nand U16584 (N_16584,N_14991,N_12809);
or U16585 (N_16585,N_11477,N_13581);
xor U16586 (N_16586,N_13765,N_14557);
nor U16587 (N_16587,N_13904,N_11575);
xnor U16588 (N_16588,N_11611,N_11941);
xnor U16589 (N_16589,N_11594,N_14575);
xor U16590 (N_16590,N_14699,N_14809);
or U16591 (N_16591,N_13179,N_10718);
nand U16592 (N_16592,N_14399,N_13867);
and U16593 (N_16593,N_14258,N_11463);
nor U16594 (N_16594,N_14954,N_10862);
nand U16595 (N_16595,N_10852,N_12116);
and U16596 (N_16596,N_13824,N_14437);
nand U16597 (N_16597,N_10017,N_12284);
nand U16598 (N_16598,N_10507,N_13286);
nand U16599 (N_16599,N_12498,N_10172);
nand U16600 (N_16600,N_13978,N_10336);
nor U16601 (N_16601,N_13723,N_14545);
xor U16602 (N_16602,N_14944,N_10170);
and U16603 (N_16603,N_11868,N_12364);
and U16604 (N_16604,N_11799,N_14271);
or U16605 (N_16605,N_12375,N_12916);
xnor U16606 (N_16606,N_12969,N_13931);
xnor U16607 (N_16607,N_11862,N_10596);
nor U16608 (N_16608,N_14751,N_12598);
xor U16609 (N_16609,N_14990,N_13639);
nand U16610 (N_16610,N_10329,N_12799);
and U16611 (N_16611,N_10954,N_11076);
or U16612 (N_16612,N_13273,N_12957);
xnor U16613 (N_16613,N_12664,N_13260);
and U16614 (N_16614,N_11977,N_13231);
nand U16615 (N_16615,N_10205,N_13769);
nand U16616 (N_16616,N_14133,N_14624);
or U16617 (N_16617,N_14003,N_13806);
and U16618 (N_16618,N_14932,N_13885);
or U16619 (N_16619,N_12774,N_11219);
xor U16620 (N_16620,N_11774,N_13647);
and U16621 (N_16621,N_14084,N_11843);
and U16622 (N_16622,N_12490,N_11508);
and U16623 (N_16623,N_13111,N_13504);
nand U16624 (N_16624,N_11350,N_10776);
nor U16625 (N_16625,N_12899,N_11013);
or U16626 (N_16626,N_10702,N_11649);
or U16627 (N_16627,N_12109,N_11953);
or U16628 (N_16628,N_13558,N_12180);
xnor U16629 (N_16629,N_11339,N_11767);
nor U16630 (N_16630,N_10210,N_10932);
nand U16631 (N_16631,N_10151,N_13583);
and U16632 (N_16632,N_11410,N_14576);
or U16633 (N_16633,N_10465,N_12418);
nor U16634 (N_16634,N_10722,N_10989);
nand U16635 (N_16635,N_12293,N_10477);
xnor U16636 (N_16636,N_13477,N_14425);
nor U16637 (N_16637,N_13301,N_11776);
or U16638 (N_16638,N_12657,N_14233);
nor U16639 (N_16639,N_13917,N_11088);
or U16640 (N_16640,N_14623,N_12282);
nand U16641 (N_16641,N_14895,N_10320);
and U16642 (N_16642,N_11944,N_12718);
nand U16643 (N_16643,N_12506,N_12419);
xnor U16644 (N_16644,N_14702,N_11555);
or U16645 (N_16645,N_14668,N_10946);
xor U16646 (N_16646,N_12685,N_14232);
and U16647 (N_16647,N_13474,N_10910);
or U16648 (N_16648,N_13694,N_14795);
xnor U16649 (N_16649,N_14090,N_11303);
xor U16650 (N_16650,N_10098,N_14165);
nand U16651 (N_16651,N_14659,N_10545);
or U16652 (N_16652,N_10689,N_10657);
or U16653 (N_16653,N_14248,N_13961);
or U16654 (N_16654,N_14518,N_13645);
nand U16655 (N_16655,N_14237,N_14434);
nor U16656 (N_16656,N_10607,N_13818);
xnor U16657 (N_16657,N_11803,N_10250);
or U16658 (N_16658,N_12335,N_11157);
xor U16659 (N_16659,N_13213,N_13343);
or U16660 (N_16660,N_11181,N_10370);
nand U16661 (N_16661,N_13138,N_11274);
nor U16662 (N_16662,N_10489,N_11948);
nor U16663 (N_16663,N_10597,N_12387);
xor U16664 (N_16664,N_13272,N_13506);
xor U16665 (N_16665,N_13858,N_12893);
nand U16666 (N_16666,N_13292,N_13040);
nand U16667 (N_16667,N_13268,N_12699);
and U16668 (N_16668,N_10581,N_10207);
xor U16669 (N_16669,N_12798,N_10833);
or U16670 (N_16670,N_13848,N_11266);
and U16671 (N_16671,N_13674,N_12697);
xor U16672 (N_16672,N_14851,N_13051);
nor U16673 (N_16673,N_13420,N_14001);
nand U16674 (N_16674,N_14050,N_11896);
nand U16675 (N_16675,N_13153,N_14774);
nand U16676 (N_16676,N_13834,N_11542);
and U16677 (N_16677,N_14256,N_12442);
and U16678 (N_16678,N_14063,N_13838);
or U16679 (N_16679,N_12974,N_14142);
or U16680 (N_16680,N_12863,N_10008);
nor U16681 (N_16681,N_12150,N_14358);
and U16682 (N_16682,N_12183,N_14744);
nor U16683 (N_16683,N_13399,N_12549);
or U16684 (N_16684,N_11773,N_14710);
xor U16685 (N_16685,N_10934,N_14911);
and U16686 (N_16686,N_14521,N_11524);
xnor U16687 (N_16687,N_12753,N_11001);
and U16688 (N_16688,N_10654,N_13551);
nand U16689 (N_16689,N_11368,N_11750);
nand U16690 (N_16690,N_12275,N_13475);
xnor U16691 (N_16691,N_11619,N_13379);
nor U16692 (N_16692,N_14558,N_12291);
and U16693 (N_16693,N_14505,N_11476);
and U16694 (N_16694,N_12032,N_14942);
nor U16695 (N_16695,N_14914,N_11998);
and U16696 (N_16696,N_12344,N_11144);
and U16697 (N_16697,N_10564,N_11184);
nor U16698 (N_16698,N_11107,N_12016);
xnor U16699 (N_16699,N_11321,N_13989);
and U16700 (N_16700,N_14755,N_10697);
and U16701 (N_16701,N_10901,N_11041);
nand U16702 (N_16702,N_13216,N_13702);
and U16703 (N_16703,N_12602,N_11761);
and U16704 (N_16704,N_13718,N_12381);
nor U16705 (N_16705,N_14352,N_11405);
xnor U16706 (N_16706,N_14794,N_14805);
and U16707 (N_16707,N_11692,N_12771);
nand U16708 (N_16708,N_11285,N_10845);
or U16709 (N_16709,N_10729,N_11371);
and U16710 (N_16710,N_13760,N_12411);
and U16711 (N_16711,N_11608,N_12371);
nor U16712 (N_16712,N_14828,N_11118);
or U16713 (N_16713,N_12394,N_10438);
and U16714 (N_16714,N_10786,N_14773);
or U16715 (N_16715,N_10485,N_14013);
xor U16716 (N_16716,N_10510,N_11688);
nand U16717 (N_16717,N_12226,N_14049);
nand U16718 (N_16718,N_12592,N_12360);
and U16719 (N_16719,N_13405,N_13642);
or U16720 (N_16720,N_10132,N_14988);
nor U16721 (N_16721,N_13096,N_11892);
xor U16722 (N_16722,N_10362,N_13636);
xor U16723 (N_16723,N_10820,N_13577);
or U16724 (N_16724,N_12319,N_11449);
nand U16725 (N_16725,N_13441,N_14969);
or U16726 (N_16726,N_11210,N_12713);
nor U16727 (N_16727,N_11551,N_13844);
nor U16728 (N_16728,N_10365,N_14440);
nor U16729 (N_16729,N_14973,N_13093);
and U16730 (N_16730,N_13457,N_12045);
nor U16731 (N_16731,N_11559,N_10114);
and U16732 (N_16732,N_14336,N_14884);
or U16733 (N_16733,N_13485,N_10434);
nor U16734 (N_16734,N_13624,N_14984);
xnor U16735 (N_16735,N_10005,N_14742);
xor U16736 (N_16736,N_13322,N_11177);
or U16737 (N_16737,N_12625,N_10281);
nor U16738 (N_16738,N_14186,N_10082);
xor U16739 (N_16739,N_10643,N_13325);
xnor U16740 (N_16740,N_14402,N_12619);
nor U16741 (N_16741,N_13611,N_11026);
nand U16742 (N_16742,N_10245,N_10500);
xor U16743 (N_16743,N_11098,N_14414);
nor U16744 (N_16744,N_13464,N_12567);
or U16745 (N_16745,N_10755,N_11881);
or U16746 (N_16746,N_12941,N_12667);
nor U16747 (N_16747,N_13954,N_11743);
and U16748 (N_16748,N_13972,N_10873);
xnor U16749 (N_16749,N_12583,N_11807);
nor U16750 (N_16750,N_10026,N_11309);
and U16751 (N_16751,N_11267,N_10771);
nor U16752 (N_16752,N_10734,N_14622);
nor U16753 (N_16753,N_12722,N_13860);
or U16754 (N_16754,N_11306,N_13042);
and U16755 (N_16755,N_14598,N_10140);
nor U16756 (N_16756,N_12985,N_10358);
and U16757 (N_16757,N_13714,N_14489);
nand U16758 (N_16758,N_12074,N_10451);
nand U16759 (N_16759,N_14578,N_14469);
and U16760 (N_16760,N_14825,N_14933);
or U16761 (N_16761,N_13977,N_12978);
nor U16762 (N_16762,N_11989,N_13344);
and U16763 (N_16763,N_12287,N_14501);
or U16764 (N_16764,N_12642,N_12494);
xor U16765 (N_16765,N_13854,N_13862);
nor U16766 (N_16766,N_10417,N_12789);
or U16767 (N_16767,N_12515,N_11623);
xor U16768 (N_16768,N_14802,N_11353);
nor U16769 (N_16769,N_12990,N_10797);
nor U16770 (N_16770,N_13152,N_14996);
nor U16771 (N_16771,N_12600,N_10937);
xor U16772 (N_16772,N_11947,N_12322);
nand U16773 (N_16773,N_12853,N_12412);
or U16774 (N_16774,N_14721,N_14225);
or U16775 (N_16775,N_12121,N_10700);
nand U16776 (N_16776,N_11846,N_13043);
xnor U16777 (N_16777,N_14614,N_13782);
and U16778 (N_16778,N_12743,N_12518);
and U16779 (N_16779,N_13908,N_14124);
or U16780 (N_16780,N_14456,N_13879);
xor U16781 (N_16781,N_13327,N_13005);
nand U16782 (N_16782,N_12648,N_10112);
and U16783 (N_16783,N_13892,N_13550);
nor U16784 (N_16784,N_12314,N_11397);
nand U16785 (N_16785,N_13052,N_14775);
or U16786 (N_16786,N_13242,N_10832);
or U16787 (N_16787,N_11167,N_14430);
and U16788 (N_16788,N_11048,N_10353);
xnor U16789 (N_16789,N_11500,N_11413);
or U16790 (N_16790,N_11886,N_13903);
nand U16791 (N_16791,N_14210,N_13566);
or U16792 (N_16792,N_11398,N_13762);
nand U16793 (N_16793,N_14690,N_14856);
xor U16794 (N_16794,N_10589,N_13091);
xor U16795 (N_16795,N_12162,N_11797);
xor U16796 (N_16796,N_13221,N_12599);
nor U16797 (N_16797,N_12577,N_10731);
nand U16798 (N_16798,N_14784,N_10677);
xnor U16799 (N_16799,N_10139,N_10872);
and U16800 (N_16800,N_10986,N_14714);
or U16801 (N_16801,N_14803,N_14272);
or U16802 (N_16802,N_12870,N_13434);
nand U16803 (N_16803,N_11163,N_13727);
nand U16804 (N_16804,N_14118,N_12169);
nand U16805 (N_16805,N_12512,N_13902);
or U16806 (N_16806,N_10675,N_13751);
nor U16807 (N_16807,N_12127,N_13880);
xor U16808 (N_16808,N_10269,N_14267);
xnor U16809 (N_16809,N_10208,N_14427);
nand U16810 (N_16810,N_10588,N_13717);
nand U16811 (N_16811,N_13438,N_12552);
nor U16812 (N_16812,N_14033,N_11443);
xor U16813 (N_16813,N_14928,N_10225);
nor U16814 (N_16814,N_14252,N_10981);
or U16815 (N_16815,N_11714,N_12698);
and U16816 (N_16816,N_11794,N_14590);
or U16817 (N_16817,N_10264,N_13522);
or U16818 (N_16818,N_11208,N_14503);
or U16819 (N_16819,N_10328,N_11698);
xor U16820 (N_16820,N_12604,N_10768);
and U16821 (N_16821,N_14074,N_11220);
or U16822 (N_16822,N_12758,N_12581);
nand U16823 (N_16823,N_13518,N_10402);
and U16824 (N_16824,N_13335,N_14113);
and U16825 (N_16825,N_13786,N_14217);
and U16826 (N_16826,N_14822,N_14220);
or U16827 (N_16827,N_12104,N_14042);
xnor U16828 (N_16828,N_12175,N_13804);
xor U16829 (N_16829,N_11817,N_14337);
and U16830 (N_16830,N_14808,N_12672);
nor U16831 (N_16831,N_11460,N_14026);
xor U16832 (N_16832,N_10914,N_14480);
and U16833 (N_16833,N_10721,N_10453);
and U16834 (N_16834,N_14639,N_13897);
nand U16835 (N_16835,N_14777,N_10898);
and U16836 (N_16836,N_13280,N_12618);
or U16837 (N_16837,N_14451,N_13661);
xnor U16838 (N_16838,N_12868,N_10117);
xnor U16839 (N_16839,N_14585,N_13756);
nand U16840 (N_16840,N_11159,N_12547);
xor U16841 (N_16841,N_12051,N_14868);
or U16842 (N_16842,N_14224,N_13829);
nor U16843 (N_16843,N_10335,N_12555);
xnor U16844 (N_16844,N_12108,N_12888);
or U16845 (N_16845,N_10452,N_13362);
xor U16846 (N_16846,N_10326,N_13704);
xor U16847 (N_16847,N_12342,N_13996);
and U16848 (N_16848,N_14708,N_11992);
nand U16849 (N_16849,N_11510,N_12704);
nand U16850 (N_16850,N_14687,N_10149);
and U16851 (N_16851,N_13036,N_10712);
and U16852 (N_16852,N_10918,N_12747);
or U16853 (N_16853,N_12773,N_10018);
nand U16854 (N_16854,N_13248,N_10369);
xor U16855 (N_16855,N_14276,N_12740);
xor U16856 (N_16856,N_11668,N_11650);
or U16857 (N_16857,N_14052,N_13095);
nand U16858 (N_16858,N_14508,N_13199);
xor U16859 (N_16859,N_12080,N_10915);
or U16860 (N_16860,N_12134,N_13055);
xor U16861 (N_16861,N_13836,N_10440);
or U16862 (N_16862,N_14534,N_12556);
xnor U16863 (N_16863,N_10201,N_14333);
nand U16864 (N_16864,N_11681,N_10188);
nand U16865 (N_16865,N_12729,N_13974);
xnor U16866 (N_16866,N_14497,N_12370);
or U16867 (N_16867,N_12107,N_11756);
nor U16868 (N_16868,N_13815,N_10556);
nand U16869 (N_16869,N_14287,N_14418);
xnor U16870 (N_16870,N_13572,N_12516);
or U16871 (N_16871,N_14909,N_11518);
or U16872 (N_16872,N_10532,N_11239);
or U16873 (N_16873,N_11099,N_13339);
nand U16874 (N_16874,N_14579,N_13313);
nor U16875 (N_16875,N_14068,N_10012);
nand U16876 (N_16876,N_13842,N_13473);
and U16877 (N_16877,N_11511,N_14209);
xor U16878 (N_16878,N_13594,N_14244);
nor U16879 (N_16879,N_13013,N_13947);
nand U16880 (N_16880,N_10106,N_12372);
and U16881 (N_16881,N_10647,N_14716);
xor U16882 (N_16882,N_12951,N_11232);
xnor U16883 (N_16883,N_13305,N_11943);
nand U16884 (N_16884,N_11589,N_10879);
or U16885 (N_16885,N_10045,N_14605);
nor U16886 (N_16886,N_12904,N_13214);
or U16887 (N_16887,N_10302,N_13234);
and U16888 (N_16888,N_14134,N_12918);
nor U16889 (N_16889,N_11584,N_10866);
nor U16890 (N_16890,N_13395,N_10356);
and U16891 (N_16891,N_14961,N_10553);
xnor U16892 (N_16892,N_10669,N_10284);
and U16893 (N_16893,N_14813,N_11590);
or U16894 (N_16894,N_12860,N_12441);
xor U16895 (N_16895,N_14203,N_13270);
or U16896 (N_16896,N_14958,N_12855);
nand U16897 (N_16897,N_13592,N_11207);
nand U16898 (N_16898,N_14726,N_13509);
xor U16899 (N_16899,N_14953,N_13394);
xnor U16900 (N_16900,N_13482,N_11176);
nor U16901 (N_16901,N_11587,N_12138);
and U16902 (N_16902,N_11922,N_14321);
xor U16903 (N_16903,N_11780,N_10234);
nor U16904 (N_16904,N_14704,N_13282);
xor U16905 (N_16905,N_14712,N_10634);
nand U16906 (N_16906,N_12415,N_12027);
and U16907 (N_16907,N_14929,N_13265);
nor U16908 (N_16908,N_13775,N_10261);
and U16909 (N_16909,N_12666,N_14010);
or U16910 (N_16910,N_12353,N_12777);
xor U16911 (N_16911,N_11424,N_12092);
nor U16912 (N_16912,N_14106,N_11647);
xor U16913 (N_16913,N_10641,N_14398);
or U16914 (N_16914,N_10458,N_12967);
nor U16915 (N_16915,N_10625,N_13075);
nand U16916 (N_16916,N_11365,N_12095);
xor U16917 (N_16917,N_14174,N_14379);
xnor U16918 (N_16918,N_12082,N_13516);
nor U16919 (N_16919,N_12714,N_10116);
or U16920 (N_16920,N_13549,N_13430);
or U16921 (N_16921,N_14636,N_14388);
or U16922 (N_16922,N_12453,N_12278);
and U16923 (N_16923,N_10396,N_10472);
xor U16924 (N_16924,N_13048,N_13121);
and U16925 (N_16925,N_12702,N_12992);
nand U16926 (N_16926,N_13805,N_14896);
xnor U16927 (N_16927,N_10418,N_12404);
xnor U16928 (N_16928,N_14376,N_14537);
nand U16929 (N_16929,N_13722,N_11223);
and U16930 (N_16930,N_11225,N_12264);
nor U16931 (N_16931,N_13863,N_13246);
and U16932 (N_16932,N_11577,N_11988);
nor U16933 (N_16933,N_10480,N_13076);
nand U16934 (N_16934,N_10659,N_14772);
xnor U16935 (N_16935,N_11859,N_12421);
and U16936 (N_16936,N_14613,N_12077);
and U16937 (N_16937,N_14562,N_13602);
nand U16938 (N_16938,N_14091,N_12144);
nor U16939 (N_16939,N_12430,N_14779);
and U16940 (N_16940,N_11901,N_11319);
xor U16941 (N_16941,N_13709,N_12744);
xnor U16942 (N_16942,N_14322,N_12327);
nor U16943 (N_16943,N_13145,N_10579);
xor U16944 (N_16944,N_13146,N_12940);
xnor U16945 (N_16945,N_13134,N_10822);
and U16946 (N_16946,N_12927,N_14486);
or U16947 (N_16947,N_12975,N_13673);
or U16948 (N_16948,N_12248,N_14730);
xor U16949 (N_16949,N_11727,N_10122);
nand U16950 (N_16950,N_14980,N_14305);
nor U16951 (N_16951,N_12005,N_14763);
nor U16952 (N_16952,N_14842,N_10266);
xnor U16953 (N_16953,N_13202,N_12042);
nand U16954 (N_16954,N_11633,N_12367);
nor U16955 (N_16955,N_11348,N_12778);
nor U16956 (N_16956,N_10334,N_10147);
xor U16957 (N_16957,N_13626,N_13332);
nor U16958 (N_16958,N_12804,N_11958);
and U16959 (N_16959,N_11063,N_13664);
nand U16960 (N_16960,N_14020,N_14878);
or U16961 (N_16961,N_11160,N_14963);
nor U16962 (N_16962,N_10387,N_14737);
nand U16963 (N_16963,N_11120,N_11085);
or U16964 (N_16964,N_13252,N_10395);
nand U16965 (N_16965,N_12227,N_14806);
nand U16966 (N_16966,N_14222,N_12334);
nor U16967 (N_16967,N_13041,N_12427);
nand U16968 (N_16968,N_11605,N_14983);
or U16969 (N_16969,N_10947,N_14394);
nor U16970 (N_16970,N_11070,N_12310);
nor U16971 (N_16971,N_11985,N_10303);
or U16972 (N_16972,N_11916,N_14531);
xor U16973 (N_16973,N_10664,N_14829);
nand U16974 (N_16974,N_13244,N_10060);
or U16975 (N_16975,N_10668,N_13945);
nor U16976 (N_16976,N_13190,N_13251);
xor U16977 (N_16977,N_13757,N_12681);
nor U16978 (N_16978,N_11291,N_14672);
nor U16979 (N_16979,N_11432,N_11364);
and U16980 (N_16980,N_11784,N_10853);
and U16981 (N_16981,N_13375,N_13851);
nand U16982 (N_16982,N_10586,N_14291);
or U16983 (N_16983,N_14560,N_13823);
nor U16984 (N_16984,N_14908,N_12475);
or U16985 (N_16985,N_10711,N_11102);
xor U16986 (N_16986,N_14302,N_11782);
nor U16987 (N_16987,N_14695,N_14273);
nand U16988 (N_16988,N_14246,N_13414);
or U16989 (N_16989,N_12006,N_10667);
and U16990 (N_16990,N_10024,N_11498);
and U16991 (N_16991,N_13046,N_14035);
and U16992 (N_16992,N_11490,N_10805);
xor U16993 (N_16993,N_11080,N_13919);
and U16994 (N_16994,N_11689,N_11361);
nand U16995 (N_16995,N_10681,N_14869);
nand U16996 (N_16996,N_13283,N_12522);
nor U16997 (N_16997,N_14021,N_10549);
nor U16998 (N_16998,N_10665,N_13876);
and U16999 (N_16999,N_13886,N_12531);
xor U17000 (N_17000,N_10864,N_12820);
or U17001 (N_17001,N_13771,N_11148);
xnor U17002 (N_17002,N_12194,N_11307);
and U17003 (N_17003,N_10756,N_13038);
nand U17004 (N_17004,N_10569,N_13608);
or U17005 (N_17005,N_13436,N_13100);
nor U17006 (N_17006,N_12140,N_12054);
nand U17007 (N_17007,N_10787,N_10965);
and U17008 (N_17008,N_13275,N_10705);
nand U17009 (N_17009,N_12871,N_14027);
nand U17010 (N_17010,N_13726,N_10777);
xnor U17011 (N_17011,N_13220,N_13841);
nor U17012 (N_17012,N_12294,N_11809);
nand U17013 (N_17013,N_14724,N_10300);
and U17014 (N_17014,N_13868,N_12368);
nand U17015 (N_17015,N_11607,N_11217);
xnor U17016 (N_17016,N_10062,N_13697);
nor U17017 (N_17017,N_14147,N_10609);
nor U17018 (N_17018,N_12928,N_10662);
nor U17019 (N_17019,N_10960,N_14653);
xor U17020 (N_17020,N_11008,N_14764);
nor U17021 (N_17021,N_12873,N_10377);
nand U17022 (N_17022,N_12070,N_14058);
xor U17023 (N_17023,N_14045,N_10357);
and U17024 (N_17024,N_13530,N_11458);
and U17025 (N_17025,N_10974,N_11047);
nand U17026 (N_17026,N_13555,N_14339);
and U17027 (N_17027,N_12087,N_13196);
xor U17028 (N_17028,N_11451,N_10605);
nor U17029 (N_17029,N_11158,N_12228);
or U17030 (N_17030,N_10254,N_13666);
or U17031 (N_17031,N_11484,N_11123);
xnor U17032 (N_17032,N_12752,N_11253);
xnor U17033 (N_17033,N_10198,N_13444);
nor U17034 (N_17034,N_11873,N_14667);
nor U17035 (N_17035,N_12400,N_10973);
nor U17036 (N_17036,N_11286,N_10258);
or U17037 (N_17037,N_11416,N_10476);
and U17038 (N_17038,N_12890,N_13846);
xor U17039 (N_17039,N_12588,N_13169);
nand U17040 (N_17040,N_11517,N_13024);
xnor U17041 (N_17041,N_11600,N_14375);
and U17042 (N_17042,N_13030,N_11771);
xor U17043 (N_17043,N_14423,N_14249);
nor U17044 (N_17044,N_12139,N_10746);
or U17045 (N_17045,N_10215,N_14611);
nand U17046 (N_17046,N_14200,N_11215);
and U17047 (N_17047,N_10340,N_10650);
and U17048 (N_17048,N_13623,N_12156);
or U17049 (N_17049,N_13417,N_11087);
and U17050 (N_17050,N_14077,N_10614);
xnor U17051 (N_17051,N_13742,N_12173);
nand U17052 (N_17052,N_10253,N_14582);
and U17053 (N_17053,N_10743,N_11396);
xor U17054 (N_17054,N_14713,N_12268);
nand U17055 (N_17055,N_11236,N_14853);
nand U17056 (N_17056,N_10769,N_11891);
xor U17057 (N_17057,N_14523,N_12584);
xor U17058 (N_17058,N_13713,N_11032);
or U17059 (N_17059,N_13411,N_13302);
and U17060 (N_17060,N_12043,N_12326);
xnor U17061 (N_17061,N_14583,N_14577);
or U17062 (N_17062,N_11277,N_14565);
or U17063 (N_17063,N_14037,N_13628);
nand U17064 (N_17064,N_14452,N_10855);
and U17065 (N_17065,N_12952,N_12211);
nor U17066 (N_17066,N_14284,N_11104);
nand U17067 (N_17067,N_14047,N_13955);
nor U17068 (N_17068,N_14044,N_11300);
xor U17069 (N_17069,N_14916,N_11252);
nand U17070 (N_17070,N_14722,N_10811);
nor U17071 (N_17071,N_12114,N_11174);
nor U17072 (N_17072,N_13987,N_13559);
nand U17073 (N_17073,N_11543,N_12263);
and U17074 (N_17074,N_14190,N_10652);
xnor U17075 (N_17075,N_13705,N_10022);
nor U17076 (N_17076,N_11984,N_13514);
xor U17077 (N_17077,N_13144,N_12239);
and U17078 (N_17078,N_14515,N_14085);
or U17079 (N_17079,N_11038,N_11185);
xor U17080 (N_17080,N_12850,N_14599);
xnor U17081 (N_17081,N_14617,N_12627);
or U17082 (N_17082,N_14922,N_14307);
nor U17083 (N_17083,N_10938,N_11433);
and U17084 (N_17084,N_10270,N_14247);
nor U17085 (N_17085,N_10093,N_12187);
and U17086 (N_17086,N_10495,N_14711);
nor U17087 (N_17087,N_14970,N_14941);
nand U17088 (N_17088,N_14478,N_11218);
xnor U17089 (N_17089,N_14053,N_11110);
and U17090 (N_17090,N_12760,N_13127);
nor U17091 (N_17091,N_10992,N_11832);
and U17092 (N_17092,N_11841,N_10374);
nand U17093 (N_17093,N_14401,N_11487);
or U17094 (N_17094,N_11568,N_10157);
and U17095 (N_17095,N_10935,N_11367);
nor U17096 (N_17096,N_14356,N_10251);
and U17097 (N_17097,N_13373,N_13986);
or U17098 (N_17098,N_12286,N_13706);
nor U17099 (N_17099,N_12500,N_12247);
or U17100 (N_17100,N_14975,N_10025);
nor U17101 (N_17101,N_11434,N_11333);
nor U17102 (N_17102,N_13544,N_10585);
or U17103 (N_17103,N_11616,N_12972);
and U17104 (N_17104,N_12078,N_13226);
and U17105 (N_17105,N_11101,N_11672);
or U17106 (N_17106,N_10169,N_11028);
nor U17107 (N_17107,N_13114,N_12720);
and U17108 (N_17108,N_11290,N_14671);
xnor U17109 (N_17109,N_13287,N_12149);
xor U17110 (N_17110,N_12914,N_11352);
nor U17111 (N_17111,N_12712,N_13388);
and U17112 (N_17112,N_13657,N_13983);
xor U17113 (N_17113,N_14069,N_13180);
nand U17114 (N_17114,N_12824,N_10421);
or U17115 (N_17115,N_14618,N_14645);
and U17116 (N_17116,N_12249,N_13491);
or U17117 (N_17117,N_12815,N_13319);
nand U17118 (N_17118,N_12887,N_10483);
or U17119 (N_17119,N_12207,N_10307);
and U17120 (N_17120,N_14780,N_11900);
nor U17121 (N_17121,N_12987,N_13203);
or U17122 (N_17122,N_10436,N_11075);
or U17123 (N_17123,N_12513,N_12179);
xnor U17124 (N_17124,N_12015,N_13028);
nand U17125 (N_17125,N_11418,N_13392);
nand U17126 (N_17126,N_11272,N_12524);
or U17127 (N_17127,N_12487,N_14462);
nor U17128 (N_17128,N_14054,N_12993);
nor U17129 (N_17129,N_13856,N_11785);
or U17130 (N_17130,N_11801,N_10222);
or U17131 (N_17131,N_13401,N_11874);
nand U17132 (N_17132,N_13607,N_10186);
xor U17133 (N_17133,N_12781,N_10163);
xor U17134 (N_17134,N_14223,N_12590);
nor U17135 (N_17135,N_10624,N_14030);
nand U17136 (N_17136,N_10518,N_10294);
or U17137 (N_17137,N_13148,N_14960);
xor U17138 (N_17138,N_11426,N_13342);
or U17139 (N_17139,N_11720,N_10814);
and U17140 (N_17140,N_12022,N_11913);
nor U17141 (N_17141,N_14178,N_11186);
xnor U17142 (N_17142,N_14791,N_10993);
xor U17143 (N_17143,N_10552,N_14393);
xnor U17144 (N_17144,N_10049,N_11676);
and U17145 (N_17145,N_14913,N_14071);
xor U17146 (N_17146,N_10426,N_13817);
xor U17147 (N_17147,N_14439,N_11735);
and U17148 (N_17148,N_10389,N_12668);
nor U17149 (N_17149,N_11314,N_10658);
nand U17150 (N_17150,N_10443,N_11703);
and U17151 (N_17151,N_13329,N_11942);
xnor U17152 (N_17152,N_14075,N_10707);
or U17153 (N_17153,N_12029,N_10645);
xnor U17154 (N_17154,N_13637,N_11327);
nand U17155 (N_17155,N_13083,N_10523);
nand U17156 (N_17156,N_14615,N_11249);
nand U17157 (N_17157,N_12196,N_13092);
nor U17158 (N_17158,N_10393,N_12934);
nand U17159 (N_17159,N_11529,N_12391);
and U17160 (N_17160,N_12963,N_10749);
nor U17161 (N_17161,N_12539,N_12929);
nor U17162 (N_17162,N_13812,N_13768);
xor U17163 (N_17163,N_14801,N_13119);
xor U17164 (N_17164,N_12424,N_13380);
nor U17165 (N_17165,N_11706,N_13269);
nor U17166 (N_17166,N_13772,N_12998);
and U17167 (N_17167,N_12596,N_13538);
xnor U17168 (N_17168,N_11072,N_10039);
or U17169 (N_17169,N_12749,N_13016);
nor U17170 (N_17170,N_11933,N_14213);
and U17171 (N_17171,N_13521,N_11388);
nor U17172 (N_17172,N_10196,N_14553);
nand U17173 (N_17173,N_11912,N_13659);
or U17174 (N_17174,N_10065,N_11918);
or U17175 (N_17175,N_11450,N_12812);
or U17176 (N_17176,N_13827,N_10638);
nand U17177 (N_17177,N_11165,N_14918);
xor U17178 (N_17178,N_11050,N_11895);
xnor U17179 (N_17179,N_13346,N_12689);
and U17180 (N_17180,N_14847,N_12459);
or U17181 (N_17181,N_14792,N_14197);
xor U17182 (N_17182,N_12252,N_12272);
nand U17183 (N_17183,N_11031,N_11620);
nor U17184 (N_17184,N_13261,N_14892);
nor U17185 (N_17185,N_11097,N_12849);
nand U17186 (N_17186,N_13081,N_14976);
nor U17187 (N_17187,N_14574,N_12966);
or U17188 (N_17188,N_13733,N_11887);
and U17189 (N_17189,N_11153,N_12630);
or U17190 (N_17190,N_10770,N_14902);
and U17191 (N_17191,N_10384,N_14240);
xor U17192 (N_17192,N_14870,N_11298);
xnor U17193 (N_17193,N_10061,N_10827);
nor U17194 (N_17194,N_10457,N_13646);
nand U17195 (N_17195,N_12526,N_12765);
or U17196 (N_17196,N_12796,N_11582);
and U17197 (N_17197,N_11516,N_12790);
and U17198 (N_17198,N_11562,N_14387);
nor U17199 (N_17199,N_14368,N_14923);
nand U17200 (N_17200,N_12451,N_13683);
and U17201 (N_17201,N_10337,N_13719);
xor U17202 (N_17202,N_13995,N_11462);
or U17203 (N_17203,N_11336,N_10728);
and U17204 (N_17204,N_11345,N_14318);
and U17205 (N_17205,N_11659,N_13712);
nand U17206 (N_17206,N_13656,N_12066);
and U17207 (N_17207,N_12037,N_10835);
nor U17208 (N_17208,N_11019,N_11169);
xor U17209 (N_17209,N_10143,N_10765);
nor U17210 (N_17210,N_12206,N_10598);
nor U17211 (N_17211,N_10187,N_12251);
and U17212 (N_17212,N_11549,N_12069);
nor U17213 (N_17213,N_14867,N_14826);
or U17214 (N_17214,N_14907,N_11671);
xnor U17215 (N_17215,N_13198,N_11861);
nand U17216 (N_17216,N_10214,N_13864);
nor U17217 (N_17217,N_10491,N_10959);
and U17218 (N_17218,N_13149,N_13098);
or U17219 (N_17219,N_11264,N_12164);
or U17220 (N_17220,N_11645,N_10842);
or U17221 (N_17221,N_13872,N_11730);
and U17222 (N_17222,N_12610,N_12099);
or U17223 (N_17223,N_11658,N_12178);
nor U17224 (N_17224,N_13988,N_12838);
nor U17225 (N_17225,N_10985,N_12570);
or U17226 (N_17226,N_13543,N_11278);
and U17227 (N_17227,N_13652,N_14935);
or U17228 (N_17228,N_10080,N_13463);
xor U17229 (N_17229,N_12546,N_13716);
or U17230 (N_17230,N_14998,N_12523);
nor U17231 (N_17231,N_13900,N_11902);
or U17232 (N_17232,N_13001,N_13933);
xor U17233 (N_17233,N_12309,N_10249);
or U17234 (N_17234,N_14407,N_14525);
xnor U17235 (N_17235,N_13237,N_13101);
or U17236 (N_17236,N_10286,N_13633);
or U17237 (N_17237,N_12787,N_13206);
nor U17238 (N_17238,N_11660,N_13178);
nor U17239 (N_17239,N_14076,N_13500);
nor U17240 (N_17240,N_10723,N_12320);
nor U17241 (N_17241,N_12766,N_13131);
nor U17242 (N_17242,N_11982,N_14733);
and U17243 (N_17243,N_12502,N_10735);
nand U17244 (N_17244,N_13930,N_11059);
nor U17245 (N_17245,N_14860,N_10773);
or U17246 (N_17246,N_11747,N_14520);
xor U17247 (N_17247,N_14905,N_13828);
or U17248 (N_17248,N_13819,N_12917);
or U17249 (N_17249,N_10341,N_11324);
nor U17250 (N_17250,N_14205,N_10291);
nor U17251 (N_17251,N_11839,N_12008);
or U17252 (N_17252,N_12079,N_11304);
xor U17253 (N_17253,N_10031,N_14164);
or U17254 (N_17254,N_11693,N_14384);
xnor U17255 (N_17255,N_10314,N_13347);
xnor U17256 (N_17256,N_13015,N_14750);
xnor U17257 (N_17257,N_14159,N_10794);
nor U17258 (N_17258,N_12902,N_13878);
and U17259 (N_17259,N_10784,N_13383);
or U17260 (N_17260,N_14438,N_14175);
and U17261 (N_17261,N_11770,N_10504);
nand U17262 (N_17262,N_11830,N_14426);
and U17263 (N_17263,N_11392,N_13128);
or U17264 (N_17264,N_12044,N_14465);
and U17265 (N_17265,N_10772,N_14701);
and U17266 (N_17266,N_13470,N_12433);
xor U17267 (N_17267,N_11204,N_10919);
and U17268 (N_17268,N_11852,N_14357);
xnor U17269 (N_17269,N_11141,N_13107);
or U17270 (N_17270,N_14259,N_10878);
and U17271 (N_17271,N_10074,N_13686);
and U17272 (N_17272,N_11261,N_13205);
or U17273 (N_17273,N_11380,N_12181);
and U17274 (N_17274,N_11812,N_12055);
nand U17275 (N_17275,N_11200,N_12946);
nor U17276 (N_17276,N_14967,N_11949);
and U17277 (N_17277,N_14361,N_14665);
or U17278 (N_17278,N_11393,N_12407);
nor U17279 (N_17279,N_12959,N_14512);
xor U17280 (N_17280,N_12705,N_10599);
nand U17281 (N_17281,N_10527,N_14854);
xnor U17282 (N_17282,N_12219,N_13739);
nand U17283 (N_17283,N_11390,N_11768);
and U17284 (N_17284,N_12947,N_12994);
xnor U17285 (N_17285,N_13821,N_12930);
and U17286 (N_17286,N_12202,N_11550);
or U17287 (N_17287,N_14485,N_14894);
nor U17288 (N_17288,N_10696,N_11626);
nand U17289 (N_17289,N_11057,N_14838);
or U17290 (N_17290,N_10964,N_11011);
or U17291 (N_17291,N_12126,N_12662);
and U17292 (N_17292,N_13054,N_12615);
xnor U17293 (N_17293,N_12637,N_12692);
nand U17294 (N_17294,N_10745,N_11222);
xnor U17295 (N_17295,N_14416,N_10894);
nor U17296 (N_17296,N_12048,N_11399);
nor U17297 (N_17297,N_10926,N_10865);
or U17298 (N_17298,N_14119,N_11674);
nand U17299 (N_17299,N_13578,N_14899);
or U17300 (N_17300,N_12285,N_11651);
or U17301 (N_17301,N_11009,N_11017);
or U17302 (N_17302,N_13161,N_10129);
or U17303 (N_17303,N_13374,N_10496);
or U17304 (N_17304,N_12693,N_13351);
or U17305 (N_17305,N_10565,N_12302);
xnor U17306 (N_17306,N_13173,N_12036);
and U17307 (N_17307,N_13672,N_11935);
and U17308 (N_17308,N_14335,N_12167);
nor U17309 (N_17309,N_11855,N_14753);
xor U17310 (N_17310,N_13707,N_10803);
nor U17311 (N_17311,N_13651,N_10079);
and U17312 (N_17312,N_14569,N_14890);
and U17313 (N_17313,N_12608,N_14056);
nor U17314 (N_17314,N_14141,N_12317);
and U17315 (N_17315,N_13670,N_13850);
nand U17316 (N_17316,N_12402,N_13615);
or U17317 (N_17317,N_11470,N_14278);
or U17318 (N_17318,N_13078,N_11270);
nor U17319 (N_17319,N_14098,N_13678);
nand U17320 (N_17320,N_10931,N_13627);
and U17321 (N_17321,N_11240,N_14946);
and U17322 (N_17322,N_10450,N_14345);
or U17323 (N_17323,N_12382,N_12046);
nor U17324 (N_17324,N_12277,N_13758);
nor U17325 (N_17325,N_14995,N_11246);
xor U17326 (N_17326,N_10289,N_12971);
nand U17327 (N_17327,N_10666,N_10925);
and U17328 (N_17328,N_12478,N_14678);
nand U17329 (N_17329,N_10913,N_12470);
or U17330 (N_17330,N_11634,N_13832);
xnor U17331 (N_17331,N_11630,N_12256);
or U17332 (N_17332,N_12170,N_11293);
or U17333 (N_17333,N_11112,N_14930);
nand U17334 (N_17334,N_10905,N_12835);
nor U17335 (N_17335,N_12783,N_13022);
or U17336 (N_17336,N_12009,N_12876);
nand U17337 (N_17337,N_14686,N_14131);
and U17338 (N_17338,N_11877,N_11957);
and U17339 (N_17339,N_10376,N_11095);
or U17340 (N_17340,N_13546,N_13185);
and U17341 (N_17341,N_10016,N_10804);
nor U17342 (N_17342,N_13994,N_11455);
nor U17343 (N_17343,N_11121,N_14904);
and U17344 (N_17344,N_14566,N_12892);
xnor U17345 (N_17345,N_13778,N_10338);
xor U17346 (N_17346,N_12063,N_14788);
nand U17347 (N_17347,N_14103,N_13982);
xnor U17348 (N_17348,N_13410,N_13170);
xnor U17349 (N_17349,N_12759,N_14977);
or U17350 (N_17350,N_14541,N_14619);
nor U17351 (N_17351,N_14846,N_14511);
nor U17352 (N_17352,N_12671,N_13425);
xnor U17353 (N_17353,N_12597,N_13364);
or U17354 (N_17354,N_11421,N_11601);
and U17355 (N_17355,N_10995,N_11864);
or U17356 (N_17356,N_10299,N_12165);
nand U17357 (N_17357,N_13233,N_11715);
or U17358 (N_17358,N_13033,N_13471);
nor U17359 (N_17359,N_10019,N_13232);
nor U17360 (N_17360,N_12234,N_11271);
or U17361 (N_17361,N_12551,N_13691);
or U17362 (N_17362,N_14315,N_12274);
or U17363 (N_17363,N_14626,N_12030);
nor U17364 (N_17364,N_12250,N_12389);
xor U17365 (N_17365,N_12669,N_12997);
nor U17366 (N_17366,N_11974,N_12468);
xnor U17367 (N_17367,N_10040,N_11020);
nand U17368 (N_17368,N_11114,N_13291);
or U17369 (N_17369,N_13998,N_14542);
nand U17370 (N_17370,N_10103,N_10090);
or U17371 (N_17371,N_12349,N_10166);
xor U17372 (N_17372,N_10517,N_14211);
or U17373 (N_17373,N_10394,N_12775);
or U17374 (N_17374,N_13418,N_13943);
nand U17375 (N_17375,N_13018,N_13781);
and U17376 (N_17376,N_12816,N_12578);
xor U17377 (N_17377,N_11412,N_11129);
nor U17378 (N_17378,N_13228,N_13586);
or U17379 (N_17379,N_12550,N_14900);
or U17380 (N_17380,N_10468,N_10104);
nor U17381 (N_17381,N_10577,N_13940);
and U17382 (N_17382,N_10714,N_12354);
nand U17383 (N_17383,N_13333,N_10789);
nand U17384 (N_17384,N_13187,N_13396);
xor U17385 (N_17385,N_14372,N_14450);
and U17386 (N_17386,N_14094,N_10262);
nand U17387 (N_17387,N_10940,N_11814);
and U17388 (N_17388,N_10120,N_11124);
nor U17389 (N_17389,N_13537,N_13254);
nand U17390 (N_17390,N_13023,N_11769);
nor U17391 (N_17391,N_12416,N_14939);
nor U17392 (N_17392,N_13990,N_13596);
and U17393 (N_17393,N_12651,N_14466);
nand U17394 (N_17394,N_10317,N_13610);
nand U17395 (N_17395,N_10760,N_10324);
xnor U17396 (N_17396,N_12135,N_12703);
nor U17397 (N_17397,N_10271,N_12948);
nor U17398 (N_17398,N_10618,N_10388);
xnor U17399 (N_17399,N_12111,N_14126);
nand U17400 (N_17400,N_13077,N_11146);
nand U17401 (N_17401,N_13427,N_10003);
nor U17402 (N_17402,N_13975,N_13109);
nand U17403 (N_17403,N_14882,N_14406);
and U17404 (N_17404,N_11919,N_12728);
xor U17405 (N_17405,N_13519,N_14362);
nor U17406 (N_17406,N_12845,N_10260);
or U17407 (N_17407,N_11583,N_10608);
xor U17408 (N_17408,N_14400,N_14490);
nand U17409 (N_17409,N_14371,N_12350);
or U17410 (N_17410,N_14563,N_13927);
xor U17411 (N_17411,N_11025,N_11867);
nor U17412 (N_17412,N_11558,N_13103);
or U17413 (N_17413,N_12654,N_11288);
or U17414 (N_17414,N_13822,N_14281);
and U17415 (N_17415,N_13932,N_13913);
xor U17416 (N_17416,N_13086,N_14277);
or U17417 (N_17417,N_10907,N_11302);
and U17418 (N_17418,N_12431,N_13752);
or U17419 (N_17419,N_12261,N_14378);
and U17420 (N_17420,N_13334,N_14442);
nor U17421 (N_17421,N_13277,N_14631);
xor U17422 (N_17422,N_13595,N_13381);
nand U17423 (N_17423,N_10408,N_14070);
nand U17424 (N_17424,N_12944,N_13384);
or U17425 (N_17425,N_14028,N_12762);
xnor U17426 (N_17426,N_10983,N_11263);
or U17427 (N_17427,N_13049,N_11042);
xnor U17428 (N_17428,N_13370,N_11878);
nor U17429 (N_17429,N_11811,N_10422);
and U17430 (N_17430,N_12736,N_12895);
and U17431 (N_17431,N_10646,N_12240);
or U17432 (N_17432,N_13753,N_14494);
nor U17433 (N_17433,N_13857,N_11787);
xor U17434 (N_17434,N_12999,N_12208);
and U17435 (N_17435,N_14080,N_11534);
xor U17436 (N_17436,N_11731,N_12296);
and U17437 (N_17437,N_13698,N_10091);
or U17438 (N_17438,N_11023,N_14312);
nor U17439 (N_17439,N_10815,N_14607);
nand U17440 (N_17440,N_12874,N_11007);
nand U17441 (N_17441,N_14620,N_12647);
or U17442 (N_17442,N_14214,N_12041);
xor U17443 (N_17443,N_12817,N_14396);
nor U17444 (N_17444,N_10229,N_11280);
nor U17445 (N_17445,N_13993,N_11214);
and U17446 (N_17446,N_11808,N_13026);
xnor U17447 (N_17447,N_14705,N_11907);
nor U17448 (N_17448,N_14571,N_10004);
and U17449 (N_17449,N_13770,N_12436);
and U17450 (N_17450,N_12559,N_11522);
nand U17451 (N_17451,N_13123,N_13505);
or U17452 (N_17452,N_13002,N_12755);
xor U17453 (N_17453,N_11971,N_11344);
or U17454 (N_17454,N_13284,N_11275);
xor U17455 (N_17455,N_10536,N_13050);
nor U17456 (N_17456,N_10023,N_10571);
and U17457 (N_17457,N_10206,N_10218);
and U17458 (N_17458,N_11061,N_14593);
nor U17459 (N_17459,N_12049,N_12467);
nand U17460 (N_17460,N_11908,N_10891);
nor U17461 (N_17461,N_12541,N_14630);
and U17462 (N_17462,N_11229,N_13355);
nor U17463 (N_17463,N_13191,N_13542);
xnor U17464 (N_17464,N_10429,N_12511);
xor U17465 (N_17465,N_11435,N_14160);
and U17466 (N_17466,N_13695,N_12473);
nor U17467 (N_17467,N_13074,N_14373);
or U17468 (N_17468,N_14179,N_14664);
nand U17469 (N_17469,N_13923,N_10482);
or U17470 (N_17470,N_14692,N_14270);
nand U17471 (N_17471,N_13211,N_12818);
and U17472 (N_17472,N_14833,N_14107);
or U17473 (N_17473,N_10481,N_11483);
nor U17474 (N_17474,N_10969,N_13424);
or U17475 (N_17475,N_10221,N_14310);
and U17476 (N_17476,N_11635,N_13285);
xor U17477 (N_17477,N_10663,N_10511);
or U17478 (N_17478,N_12231,N_12199);
xnor U17479 (N_17479,N_11966,N_12094);
nand U17480 (N_17480,N_11472,N_13741);
or U17481 (N_17481,N_11721,N_12486);
or U17482 (N_17482,N_10455,N_14796);
or U17483 (N_17483,N_11554,N_10099);
and U17484 (N_17484,N_11621,N_10410);
nor U17485 (N_17485,N_12509,N_10821);
and U17486 (N_17486,N_11606,N_11425);
or U17487 (N_17487,N_12763,N_10069);
or U17488 (N_17488,N_14046,N_14517);
nand U17489 (N_17489,N_14782,N_14347);
nor U17490 (N_17490,N_10354,N_12110);
xor U17491 (N_17491,N_10102,N_11613);
nand U17492 (N_17492,N_13136,N_14129);
nor U17493 (N_17493,N_12025,N_14471);
and U17494 (N_17494,N_10137,N_14431);
nand U17495 (N_17495,N_14390,N_11673);
and U17496 (N_17496,N_11565,N_10848);
and U17497 (N_17497,N_14286,N_12270);
nor U17498 (N_17498,N_13159,N_11242);
and U17499 (N_17499,N_12606,N_13432);
or U17500 (N_17500,N_13968,N_14301);
and U17501 (N_17501,N_13805,N_12252);
xnor U17502 (N_17502,N_14193,N_12124);
nor U17503 (N_17503,N_13193,N_12641);
nor U17504 (N_17504,N_14860,N_11198);
xor U17505 (N_17505,N_12903,N_10074);
xnor U17506 (N_17506,N_12244,N_10074);
nand U17507 (N_17507,N_14922,N_13340);
or U17508 (N_17508,N_13319,N_13759);
nand U17509 (N_17509,N_10245,N_11251);
and U17510 (N_17510,N_10975,N_11863);
nor U17511 (N_17511,N_13168,N_14454);
nor U17512 (N_17512,N_11367,N_12183);
nand U17513 (N_17513,N_12782,N_13469);
nand U17514 (N_17514,N_10797,N_13061);
nor U17515 (N_17515,N_13577,N_12995);
nand U17516 (N_17516,N_10087,N_12491);
nand U17517 (N_17517,N_14983,N_10335);
or U17518 (N_17518,N_12939,N_10553);
xor U17519 (N_17519,N_11313,N_12386);
xnor U17520 (N_17520,N_11342,N_10391);
nor U17521 (N_17521,N_11660,N_13494);
and U17522 (N_17522,N_12240,N_12984);
or U17523 (N_17523,N_11054,N_11279);
or U17524 (N_17524,N_14516,N_11609);
nor U17525 (N_17525,N_13249,N_13751);
and U17526 (N_17526,N_14584,N_11770);
nand U17527 (N_17527,N_12102,N_13479);
xnor U17528 (N_17528,N_13462,N_11248);
xnor U17529 (N_17529,N_14138,N_10249);
and U17530 (N_17530,N_13387,N_10494);
nand U17531 (N_17531,N_12316,N_12288);
xor U17532 (N_17532,N_14653,N_14216);
nor U17533 (N_17533,N_11577,N_12110);
or U17534 (N_17534,N_12766,N_12616);
xnor U17535 (N_17535,N_12422,N_12482);
nor U17536 (N_17536,N_13232,N_12192);
nand U17537 (N_17537,N_14722,N_12759);
and U17538 (N_17538,N_10183,N_12745);
xnor U17539 (N_17539,N_12853,N_11356);
nor U17540 (N_17540,N_13091,N_12748);
nor U17541 (N_17541,N_11366,N_14606);
nand U17542 (N_17542,N_13244,N_13687);
and U17543 (N_17543,N_13117,N_10764);
and U17544 (N_17544,N_10832,N_14805);
and U17545 (N_17545,N_10589,N_11171);
xor U17546 (N_17546,N_13917,N_12570);
xnor U17547 (N_17547,N_12869,N_11709);
nor U17548 (N_17548,N_12969,N_12484);
xnor U17549 (N_17549,N_10225,N_12052);
xor U17550 (N_17550,N_12642,N_12152);
nand U17551 (N_17551,N_13610,N_10044);
or U17552 (N_17552,N_14894,N_13114);
or U17553 (N_17553,N_11925,N_11504);
nand U17554 (N_17554,N_14498,N_12636);
nor U17555 (N_17555,N_11153,N_14219);
nor U17556 (N_17556,N_12055,N_13311);
or U17557 (N_17557,N_14765,N_11324);
nand U17558 (N_17558,N_10776,N_14392);
nor U17559 (N_17559,N_12614,N_11814);
or U17560 (N_17560,N_11814,N_10172);
nor U17561 (N_17561,N_11521,N_14848);
nand U17562 (N_17562,N_10121,N_12973);
xnor U17563 (N_17563,N_13598,N_12652);
nor U17564 (N_17564,N_13782,N_10724);
and U17565 (N_17565,N_10212,N_10341);
nor U17566 (N_17566,N_13376,N_12135);
nor U17567 (N_17567,N_14560,N_14637);
xor U17568 (N_17568,N_14099,N_10364);
xor U17569 (N_17569,N_13511,N_14782);
and U17570 (N_17570,N_10288,N_13150);
nor U17571 (N_17571,N_13381,N_12440);
or U17572 (N_17572,N_12413,N_14832);
and U17573 (N_17573,N_12543,N_10488);
xnor U17574 (N_17574,N_12325,N_10620);
or U17575 (N_17575,N_12345,N_14075);
and U17576 (N_17576,N_11683,N_10274);
or U17577 (N_17577,N_13248,N_14373);
and U17578 (N_17578,N_13253,N_10747);
xor U17579 (N_17579,N_14209,N_11927);
and U17580 (N_17580,N_12047,N_12852);
nand U17581 (N_17581,N_11396,N_11770);
xor U17582 (N_17582,N_14896,N_14763);
xor U17583 (N_17583,N_12197,N_10046);
and U17584 (N_17584,N_10696,N_10442);
nor U17585 (N_17585,N_10413,N_13318);
nand U17586 (N_17586,N_14129,N_10703);
or U17587 (N_17587,N_12323,N_10913);
nand U17588 (N_17588,N_13425,N_14646);
xnor U17589 (N_17589,N_14499,N_14989);
and U17590 (N_17590,N_13640,N_14714);
nor U17591 (N_17591,N_13576,N_11047);
and U17592 (N_17592,N_12614,N_14735);
and U17593 (N_17593,N_10210,N_12195);
xor U17594 (N_17594,N_12091,N_11756);
nand U17595 (N_17595,N_10396,N_11460);
and U17596 (N_17596,N_12369,N_12354);
and U17597 (N_17597,N_11598,N_14858);
or U17598 (N_17598,N_11694,N_10354);
xnor U17599 (N_17599,N_12487,N_12651);
xor U17600 (N_17600,N_13844,N_14346);
nand U17601 (N_17601,N_11636,N_13024);
and U17602 (N_17602,N_13548,N_13533);
and U17603 (N_17603,N_13214,N_13132);
and U17604 (N_17604,N_10897,N_10058);
or U17605 (N_17605,N_14389,N_13292);
xnor U17606 (N_17606,N_13553,N_14980);
xor U17607 (N_17607,N_11557,N_12596);
nand U17608 (N_17608,N_14908,N_13834);
nor U17609 (N_17609,N_10599,N_14196);
xnor U17610 (N_17610,N_12080,N_12702);
nor U17611 (N_17611,N_12604,N_12080);
xnor U17612 (N_17612,N_12053,N_10592);
nand U17613 (N_17613,N_12373,N_14446);
nand U17614 (N_17614,N_13753,N_13639);
nand U17615 (N_17615,N_11191,N_13121);
and U17616 (N_17616,N_12633,N_14528);
or U17617 (N_17617,N_11697,N_10998);
nor U17618 (N_17618,N_10005,N_14391);
nor U17619 (N_17619,N_11279,N_13683);
or U17620 (N_17620,N_12801,N_11679);
nor U17621 (N_17621,N_13365,N_13802);
and U17622 (N_17622,N_12860,N_10577);
nand U17623 (N_17623,N_12703,N_10616);
nand U17624 (N_17624,N_12507,N_12051);
nand U17625 (N_17625,N_10846,N_10087);
and U17626 (N_17626,N_13304,N_10591);
nand U17627 (N_17627,N_13409,N_12424);
nor U17628 (N_17628,N_13431,N_13570);
xor U17629 (N_17629,N_12777,N_14911);
and U17630 (N_17630,N_10120,N_11183);
xnor U17631 (N_17631,N_10717,N_12776);
xor U17632 (N_17632,N_11999,N_11363);
or U17633 (N_17633,N_12434,N_12951);
xor U17634 (N_17634,N_14911,N_13887);
nor U17635 (N_17635,N_12019,N_12358);
nor U17636 (N_17636,N_11578,N_14055);
xnor U17637 (N_17637,N_12489,N_14957);
or U17638 (N_17638,N_12175,N_10126);
or U17639 (N_17639,N_11795,N_12781);
or U17640 (N_17640,N_11961,N_12116);
and U17641 (N_17641,N_14247,N_11403);
and U17642 (N_17642,N_10786,N_13356);
and U17643 (N_17643,N_10599,N_12021);
nor U17644 (N_17644,N_11428,N_11861);
and U17645 (N_17645,N_13426,N_10973);
nor U17646 (N_17646,N_12141,N_14104);
or U17647 (N_17647,N_11952,N_12455);
and U17648 (N_17648,N_14254,N_12867);
and U17649 (N_17649,N_14437,N_11641);
or U17650 (N_17650,N_13584,N_12216);
xor U17651 (N_17651,N_13042,N_10231);
and U17652 (N_17652,N_13202,N_12613);
nand U17653 (N_17653,N_14951,N_12175);
nand U17654 (N_17654,N_12667,N_10862);
nand U17655 (N_17655,N_13388,N_10098);
or U17656 (N_17656,N_10536,N_14592);
nor U17657 (N_17657,N_14368,N_14162);
xnor U17658 (N_17658,N_14091,N_13053);
xor U17659 (N_17659,N_11318,N_12751);
or U17660 (N_17660,N_11019,N_13455);
xnor U17661 (N_17661,N_12676,N_12167);
xor U17662 (N_17662,N_13960,N_10457);
and U17663 (N_17663,N_14597,N_14442);
xnor U17664 (N_17664,N_10328,N_13132);
or U17665 (N_17665,N_10234,N_13926);
and U17666 (N_17666,N_11071,N_12959);
nand U17667 (N_17667,N_11350,N_10919);
xnor U17668 (N_17668,N_13295,N_10376);
or U17669 (N_17669,N_14696,N_11632);
and U17670 (N_17670,N_13082,N_13325);
and U17671 (N_17671,N_11569,N_14367);
and U17672 (N_17672,N_13317,N_10713);
or U17673 (N_17673,N_11910,N_13841);
or U17674 (N_17674,N_10893,N_11889);
xor U17675 (N_17675,N_11278,N_12394);
nor U17676 (N_17676,N_14530,N_14565);
nor U17677 (N_17677,N_11166,N_11079);
or U17678 (N_17678,N_14092,N_14686);
or U17679 (N_17679,N_14610,N_13926);
nor U17680 (N_17680,N_11297,N_13811);
and U17681 (N_17681,N_12100,N_11015);
nand U17682 (N_17682,N_13065,N_13849);
nor U17683 (N_17683,N_12228,N_12791);
xnor U17684 (N_17684,N_10086,N_13829);
nor U17685 (N_17685,N_11751,N_10122);
xnor U17686 (N_17686,N_12679,N_12081);
nand U17687 (N_17687,N_14469,N_12576);
or U17688 (N_17688,N_12449,N_14875);
xor U17689 (N_17689,N_10313,N_12208);
and U17690 (N_17690,N_11216,N_10858);
nand U17691 (N_17691,N_13668,N_10212);
xor U17692 (N_17692,N_11519,N_13460);
or U17693 (N_17693,N_11536,N_14833);
nor U17694 (N_17694,N_14262,N_10969);
or U17695 (N_17695,N_14273,N_13424);
nor U17696 (N_17696,N_10753,N_13762);
or U17697 (N_17697,N_11416,N_11044);
or U17698 (N_17698,N_14624,N_12744);
or U17699 (N_17699,N_10486,N_12251);
nor U17700 (N_17700,N_12563,N_14778);
nor U17701 (N_17701,N_10968,N_12038);
nand U17702 (N_17702,N_10509,N_10375);
xor U17703 (N_17703,N_13183,N_14537);
nand U17704 (N_17704,N_13944,N_11529);
nor U17705 (N_17705,N_11606,N_13643);
nand U17706 (N_17706,N_13150,N_10921);
nand U17707 (N_17707,N_12801,N_10319);
xor U17708 (N_17708,N_10856,N_12217);
nand U17709 (N_17709,N_11821,N_13239);
nor U17710 (N_17710,N_11527,N_11463);
nand U17711 (N_17711,N_14218,N_10824);
and U17712 (N_17712,N_10749,N_10366);
or U17713 (N_17713,N_14730,N_10962);
xnor U17714 (N_17714,N_13175,N_12408);
nand U17715 (N_17715,N_14580,N_12779);
nand U17716 (N_17716,N_12094,N_11551);
nand U17717 (N_17717,N_13993,N_14427);
xnor U17718 (N_17718,N_10239,N_10806);
nand U17719 (N_17719,N_12751,N_13534);
and U17720 (N_17720,N_10002,N_11143);
and U17721 (N_17721,N_12794,N_14441);
or U17722 (N_17722,N_14601,N_10617);
nor U17723 (N_17723,N_12022,N_12298);
nand U17724 (N_17724,N_13657,N_11824);
and U17725 (N_17725,N_13668,N_10164);
or U17726 (N_17726,N_11537,N_11984);
xor U17727 (N_17727,N_10629,N_13496);
nor U17728 (N_17728,N_14753,N_10739);
nor U17729 (N_17729,N_11743,N_14386);
and U17730 (N_17730,N_11303,N_13876);
xnor U17731 (N_17731,N_14503,N_14793);
xor U17732 (N_17732,N_13508,N_13109);
nor U17733 (N_17733,N_14384,N_11757);
or U17734 (N_17734,N_11890,N_14931);
or U17735 (N_17735,N_11229,N_14893);
and U17736 (N_17736,N_13433,N_14654);
or U17737 (N_17737,N_13183,N_14771);
xor U17738 (N_17738,N_13146,N_11601);
and U17739 (N_17739,N_14774,N_14438);
and U17740 (N_17740,N_11312,N_12867);
xnor U17741 (N_17741,N_14528,N_11944);
nor U17742 (N_17742,N_10730,N_14932);
nor U17743 (N_17743,N_11804,N_12276);
and U17744 (N_17744,N_12836,N_10143);
or U17745 (N_17745,N_13233,N_14046);
and U17746 (N_17746,N_14888,N_11801);
nand U17747 (N_17747,N_10047,N_12841);
xnor U17748 (N_17748,N_11221,N_11365);
nor U17749 (N_17749,N_11822,N_14968);
xor U17750 (N_17750,N_11629,N_14256);
or U17751 (N_17751,N_10565,N_12447);
nand U17752 (N_17752,N_10723,N_10608);
nand U17753 (N_17753,N_14449,N_13188);
or U17754 (N_17754,N_12419,N_11161);
nand U17755 (N_17755,N_13766,N_12400);
xnor U17756 (N_17756,N_13363,N_12575);
or U17757 (N_17757,N_12579,N_14802);
and U17758 (N_17758,N_10529,N_11728);
nor U17759 (N_17759,N_13823,N_10715);
and U17760 (N_17760,N_12438,N_13717);
nor U17761 (N_17761,N_11818,N_13084);
and U17762 (N_17762,N_13005,N_13102);
nand U17763 (N_17763,N_12543,N_11004);
xor U17764 (N_17764,N_11573,N_10485);
and U17765 (N_17765,N_13418,N_14184);
and U17766 (N_17766,N_12532,N_11173);
nand U17767 (N_17767,N_10315,N_12124);
or U17768 (N_17768,N_10523,N_11338);
or U17769 (N_17769,N_11495,N_12846);
and U17770 (N_17770,N_11296,N_11482);
or U17771 (N_17771,N_12094,N_11416);
nor U17772 (N_17772,N_14654,N_10970);
or U17773 (N_17773,N_14151,N_14375);
nor U17774 (N_17774,N_12047,N_14479);
xor U17775 (N_17775,N_11817,N_11909);
and U17776 (N_17776,N_14380,N_13344);
or U17777 (N_17777,N_11895,N_11590);
nor U17778 (N_17778,N_14784,N_13094);
nand U17779 (N_17779,N_14637,N_13900);
or U17780 (N_17780,N_13181,N_12186);
xor U17781 (N_17781,N_10979,N_11032);
nor U17782 (N_17782,N_10370,N_11728);
nor U17783 (N_17783,N_10318,N_13241);
nor U17784 (N_17784,N_12343,N_13176);
nand U17785 (N_17785,N_11572,N_11273);
and U17786 (N_17786,N_10748,N_10967);
nor U17787 (N_17787,N_13795,N_13270);
nor U17788 (N_17788,N_13965,N_11627);
nor U17789 (N_17789,N_14384,N_10694);
nand U17790 (N_17790,N_12078,N_12690);
nor U17791 (N_17791,N_14360,N_10389);
xor U17792 (N_17792,N_11027,N_11464);
nor U17793 (N_17793,N_10357,N_11667);
and U17794 (N_17794,N_10766,N_13396);
or U17795 (N_17795,N_13573,N_11424);
or U17796 (N_17796,N_14823,N_13169);
and U17797 (N_17797,N_13664,N_11717);
xnor U17798 (N_17798,N_13650,N_13977);
and U17799 (N_17799,N_13292,N_11284);
xnor U17800 (N_17800,N_12212,N_10971);
nor U17801 (N_17801,N_10553,N_13859);
and U17802 (N_17802,N_12146,N_13835);
or U17803 (N_17803,N_11206,N_11741);
and U17804 (N_17804,N_10441,N_12111);
nand U17805 (N_17805,N_12235,N_12791);
or U17806 (N_17806,N_10467,N_14904);
and U17807 (N_17807,N_13611,N_11165);
nor U17808 (N_17808,N_10911,N_12081);
or U17809 (N_17809,N_10668,N_12795);
xor U17810 (N_17810,N_14314,N_10541);
and U17811 (N_17811,N_14773,N_11657);
nor U17812 (N_17812,N_11648,N_14566);
nand U17813 (N_17813,N_14432,N_12414);
nor U17814 (N_17814,N_12744,N_14814);
or U17815 (N_17815,N_10751,N_14401);
and U17816 (N_17816,N_12790,N_12114);
or U17817 (N_17817,N_11892,N_13599);
or U17818 (N_17818,N_12461,N_13141);
nor U17819 (N_17819,N_13842,N_10685);
nor U17820 (N_17820,N_11928,N_12179);
and U17821 (N_17821,N_11700,N_13897);
xnor U17822 (N_17822,N_11943,N_11666);
and U17823 (N_17823,N_13513,N_11705);
or U17824 (N_17824,N_13662,N_12703);
xor U17825 (N_17825,N_10552,N_12948);
xor U17826 (N_17826,N_14124,N_10932);
xor U17827 (N_17827,N_11577,N_14694);
nor U17828 (N_17828,N_10196,N_13615);
nand U17829 (N_17829,N_12950,N_14628);
xor U17830 (N_17830,N_10622,N_12566);
or U17831 (N_17831,N_10721,N_11280);
nand U17832 (N_17832,N_10587,N_11628);
and U17833 (N_17833,N_10860,N_12597);
xor U17834 (N_17834,N_12151,N_11989);
xnor U17835 (N_17835,N_13838,N_12823);
and U17836 (N_17836,N_11777,N_12349);
and U17837 (N_17837,N_12837,N_13752);
nor U17838 (N_17838,N_12907,N_10038);
nand U17839 (N_17839,N_13434,N_12326);
nor U17840 (N_17840,N_11951,N_11765);
nor U17841 (N_17841,N_14040,N_14592);
nor U17842 (N_17842,N_12466,N_14982);
and U17843 (N_17843,N_14761,N_12362);
xor U17844 (N_17844,N_13753,N_10865);
nand U17845 (N_17845,N_10830,N_12997);
nor U17846 (N_17846,N_14786,N_13735);
xnor U17847 (N_17847,N_13175,N_11827);
nand U17848 (N_17848,N_12265,N_12280);
nand U17849 (N_17849,N_13165,N_14081);
and U17850 (N_17850,N_14490,N_12380);
xnor U17851 (N_17851,N_11635,N_11733);
nor U17852 (N_17852,N_13951,N_10065);
nand U17853 (N_17853,N_11438,N_12743);
or U17854 (N_17854,N_13461,N_11511);
nand U17855 (N_17855,N_12754,N_14624);
or U17856 (N_17856,N_10429,N_14455);
nor U17857 (N_17857,N_13771,N_10245);
and U17858 (N_17858,N_14870,N_10905);
and U17859 (N_17859,N_13731,N_12678);
nor U17860 (N_17860,N_11628,N_10371);
or U17861 (N_17861,N_10730,N_11526);
nand U17862 (N_17862,N_13299,N_10684);
nor U17863 (N_17863,N_10391,N_10465);
xor U17864 (N_17864,N_13183,N_14610);
or U17865 (N_17865,N_13664,N_11594);
xnor U17866 (N_17866,N_10557,N_10277);
xnor U17867 (N_17867,N_10162,N_10565);
xor U17868 (N_17868,N_14280,N_12179);
or U17869 (N_17869,N_10687,N_10337);
xor U17870 (N_17870,N_14824,N_13233);
and U17871 (N_17871,N_10485,N_13651);
or U17872 (N_17872,N_13929,N_10410);
and U17873 (N_17873,N_11673,N_14261);
and U17874 (N_17874,N_12932,N_14926);
and U17875 (N_17875,N_13198,N_12714);
nor U17876 (N_17876,N_13703,N_13495);
or U17877 (N_17877,N_12852,N_14421);
nor U17878 (N_17878,N_10106,N_13194);
or U17879 (N_17879,N_13169,N_11055);
and U17880 (N_17880,N_14342,N_10181);
nor U17881 (N_17881,N_12415,N_13306);
and U17882 (N_17882,N_14372,N_11541);
or U17883 (N_17883,N_11573,N_12722);
nand U17884 (N_17884,N_10462,N_12469);
and U17885 (N_17885,N_11546,N_11760);
and U17886 (N_17886,N_14266,N_14406);
and U17887 (N_17887,N_11840,N_13656);
xor U17888 (N_17888,N_10063,N_13321);
or U17889 (N_17889,N_11740,N_13112);
and U17890 (N_17890,N_14062,N_10313);
nand U17891 (N_17891,N_14157,N_12733);
nor U17892 (N_17892,N_13983,N_11115);
nand U17893 (N_17893,N_13419,N_12282);
xnor U17894 (N_17894,N_12041,N_13406);
nand U17895 (N_17895,N_10126,N_10003);
xnor U17896 (N_17896,N_14907,N_11770);
xor U17897 (N_17897,N_10833,N_10429);
or U17898 (N_17898,N_14640,N_14490);
and U17899 (N_17899,N_10654,N_14933);
nor U17900 (N_17900,N_11841,N_11375);
and U17901 (N_17901,N_14151,N_11401);
nand U17902 (N_17902,N_11853,N_14099);
xnor U17903 (N_17903,N_10182,N_13612);
nand U17904 (N_17904,N_14860,N_12607);
and U17905 (N_17905,N_12160,N_13295);
xnor U17906 (N_17906,N_14494,N_14831);
nor U17907 (N_17907,N_12709,N_12328);
nor U17908 (N_17908,N_13666,N_12692);
or U17909 (N_17909,N_12269,N_10749);
or U17910 (N_17910,N_10716,N_11945);
xnor U17911 (N_17911,N_12231,N_14617);
xnor U17912 (N_17912,N_11192,N_12176);
and U17913 (N_17913,N_14261,N_11811);
or U17914 (N_17914,N_10376,N_14110);
and U17915 (N_17915,N_14001,N_13437);
xnor U17916 (N_17916,N_10583,N_10058);
xor U17917 (N_17917,N_12878,N_12489);
and U17918 (N_17918,N_14155,N_14861);
and U17919 (N_17919,N_10656,N_14907);
or U17920 (N_17920,N_14927,N_14068);
and U17921 (N_17921,N_14048,N_14756);
xor U17922 (N_17922,N_13716,N_12560);
nor U17923 (N_17923,N_10167,N_13314);
nor U17924 (N_17924,N_13855,N_14023);
nand U17925 (N_17925,N_10197,N_11614);
nor U17926 (N_17926,N_14540,N_12268);
or U17927 (N_17927,N_13530,N_14616);
nand U17928 (N_17928,N_11618,N_12826);
nand U17929 (N_17929,N_12893,N_11656);
nor U17930 (N_17930,N_11941,N_11506);
xnor U17931 (N_17931,N_10637,N_10468);
nand U17932 (N_17932,N_12655,N_10080);
or U17933 (N_17933,N_14145,N_13063);
and U17934 (N_17934,N_14875,N_10052);
or U17935 (N_17935,N_12606,N_13973);
xor U17936 (N_17936,N_14720,N_10510);
or U17937 (N_17937,N_11721,N_10049);
xnor U17938 (N_17938,N_13293,N_10178);
or U17939 (N_17939,N_13829,N_10113);
nor U17940 (N_17940,N_12545,N_13364);
and U17941 (N_17941,N_10785,N_10839);
or U17942 (N_17942,N_14764,N_14664);
nand U17943 (N_17943,N_11804,N_14487);
or U17944 (N_17944,N_10630,N_12681);
xor U17945 (N_17945,N_13471,N_14665);
xnor U17946 (N_17946,N_12565,N_13483);
or U17947 (N_17947,N_13203,N_13834);
and U17948 (N_17948,N_12281,N_12684);
xnor U17949 (N_17949,N_11810,N_11284);
and U17950 (N_17950,N_14007,N_10243);
nor U17951 (N_17951,N_13492,N_12103);
or U17952 (N_17952,N_13063,N_11375);
or U17953 (N_17953,N_12892,N_10768);
nor U17954 (N_17954,N_12622,N_10125);
nor U17955 (N_17955,N_14665,N_13774);
xor U17956 (N_17956,N_11738,N_12818);
or U17957 (N_17957,N_11689,N_13154);
or U17958 (N_17958,N_13370,N_13840);
and U17959 (N_17959,N_10314,N_10559);
nand U17960 (N_17960,N_13371,N_13530);
nand U17961 (N_17961,N_13321,N_14654);
nand U17962 (N_17962,N_10847,N_13035);
nor U17963 (N_17963,N_14435,N_10800);
or U17964 (N_17964,N_14957,N_13524);
or U17965 (N_17965,N_12150,N_13957);
xnor U17966 (N_17966,N_13668,N_14820);
xor U17967 (N_17967,N_14852,N_11960);
xnor U17968 (N_17968,N_11815,N_12185);
and U17969 (N_17969,N_11433,N_10848);
xnor U17970 (N_17970,N_13318,N_10786);
or U17971 (N_17971,N_10971,N_10694);
nand U17972 (N_17972,N_14413,N_13365);
or U17973 (N_17973,N_10529,N_13736);
or U17974 (N_17974,N_14166,N_13199);
and U17975 (N_17975,N_11761,N_14680);
nand U17976 (N_17976,N_14968,N_13424);
or U17977 (N_17977,N_14216,N_11235);
nor U17978 (N_17978,N_11286,N_10282);
nor U17979 (N_17979,N_10801,N_13398);
and U17980 (N_17980,N_13897,N_11279);
and U17981 (N_17981,N_13951,N_11846);
nor U17982 (N_17982,N_10428,N_13155);
xor U17983 (N_17983,N_12128,N_10116);
xnor U17984 (N_17984,N_12970,N_11807);
xor U17985 (N_17985,N_12131,N_13403);
and U17986 (N_17986,N_11309,N_13239);
xor U17987 (N_17987,N_10247,N_14815);
and U17988 (N_17988,N_10753,N_12405);
xor U17989 (N_17989,N_11381,N_13561);
and U17990 (N_17990,N_12268,N_12309);
nand U17991 (N_17991,N_14994,N_13020);
and U17992 (N_17992,N_10824,N_12773);
and U17993 (N_17993,N_11037,N_11147);
and U17994 (N_17994,N_12232,N_12356);
or U17995 (N_17995,N_10125,N_10036);
nor U17996 (N_17996,N_11956,N_10769);
nand U17997 (N_17997,N_10756,N_10349);
nor U17998 (N_17998,N_12707,N_13966);
xnor U17999 (N_17999,N_10266,N_13606);
xor U18000 (N_18000,N_14888,N_11639);
nor U18001 (N_18001,N_13603,N_13846);
xor U18002 (N_18002,N_14335,N_12686);
xor U18003 (N_18003,N_11182,N_11125);
nor U18004 (N_18004,N_11421,N_14685);
and U18005 (N_18005,N_11071,N_10693);
nor U18006 (N_18006,N_11715,N_14813);
and U18007 (N_18007,N_10790,N_11721);
xor U18008 (N_18008,N_10284,N_10803);
xnor U18009 (N_18009,N_14961,N_11803);
and U18010 (N_18010,N_13751,N_14889);
or U18011 (N_18011,N_13743,N_10445);
nand U18012 (N_18012,N_14071,N_12533);
or U18013 (N_18013,N_10792,N_10249);
nor U18014 (N_18014,N_11826,N_14923);
nor U18015 (N_18015,N_14973,N_13263);
xnor U18016 (N_18016,N_10026,N_13337);
xor U18017 (N_18017,N_10414,N_10552);
and U18018 (N_18018,N_14518,N_11437);
xnor U18019 (N_18019,N_13133,N_13632);
or U18020 (N_18020,N_10948,N_10839);
xor U18021 (N_18021,N_12547,N_14836);
nor U18022 (N_18022,N_14251,N_13826);
nor U18023 (N_18023,N_11440,N_11962);
and U18024 (N_18024,N_14714,N_14413);
xor U18025 (N_18025,N_11116,N_12128);
nor U18026 (N_18026,N_10039,N_10830);
and U18027 (N_18027,N_11147,N_13869);
nand U18028 (N_18028,N_12892,N_13150);
xnor U18029 (N_18029,N_11362,N_10373);
and U18030 (N_18030,N_13928,N_13297);
nor U18031 (N_18031,N_13751,N_10701);
and U18032 (N_18032,N_10285,N_10974);
nand U18033 (N_18033,N_12264,N_13026);
and U18034 (N_18034,N_11954,N_10340);
xor U18035 (N_18035,N_12986,N_10439);
nor U18036 (N_18036,N_14772,N_10293);
xor U18037 (N_18037,N_12372,N_14077);
xnor U18038 (N_18038,N_13976,N_14427);
or U18039 (N_18039,N_12351,N_12231);
nand U18040 (N_18040,N_14195,N_11803);
and U18041 (N_18041,N_13412,N_13914);
xnor U18042 (N_18042,N_10397,N_11863);
xnor U18043 (N_18043,N_11758,N_12788);
nand U18044 (N_18044,N_11766,N_12163);
and U18045 (N_18045,N_13730,N_13429);
xnor U18046 (N_18046,N_14044,N_14470);
or U18047 (N_18047,N_14700,N_11613);
or U18048 (N_18048,N_14727,N_14283);
xnor U18049 (N_18049,N_12085,N_13321);
nor U18050 (N_18050,N_13735,N_12774);
xnor U18051 (N_18051,N_10775,N_10771);
and U18052 (N_18052,N_13349,N_13704);
nand U18053 (N_18053,N_10560,N_13182);
xnor U18054 (N_18054,N_12585,N_14788);
nand U18055 (N_18055,N_12032,N_12636);
xor U18056 (N_18056,N_14885,N_10264);
nand U18057 (N_18057,N_12189,N_14074);
xnor U18058 (N_18058,N_14187,N_11362);
and U18059 (N_18059,N_10272,N_12881);
xor U18060 (N_18060,N_10468,N_12869);
and U18061 (N_18061,N_13679,N_14398);
or U18062 (N_18062,N_13497,N_12677);
nand U18063 (N_18063,N_14728,N_14308);
and U18064 (N_18064,N_12458,N_12375);
or U18065 (N_18065,N_12612,N_14958);
or U18066 (N_18066,N_10874,N_10133);
or U18067 (N_18067,N_10334,N_12498);
xor U18068 (N_18068,N_10224,N_14458);
xnor U18069 (N_18069,N_12077,N_12276);
or U18070 (N_18070,N_11851,N_12940);
or U18071 (N_18071,N_13549,N_10875);
or U18072 (N_18072,N_13856,N_12127);
nand U18073 (N_18073,N_11039,N_13524);
and U18074 (N_18074,N_12492,N_10750);
nand U18075 (N_18075,N_13589,N_12347);
xnor U18076 (N_18076,N_13408,N_12647);
or U18077 (N_18077,N_10850,N_12447);
xor U18078 (N_18078,N_12408,N_13879);
or U18079 (N_18079,N_10367,N_13279);
xnor U18080 (N_18080,N_12367,N_11047);
and U18081 (N_18081,N_13974,N_13627);
and U18082 (N_18082,N_10620,N_13186);
xnor U18083 (N_18083,N_11875,N_10934);
nand U18084 (N_18084,N_14596,N_13374);
and U18085 (N_18085,N_12488,N_10936);
nand U18086 (N_18086,N_14934,N_12741);
and U18087 (N_18087,N_13440,N_14066);
and U18088 (N_18088,N_11794,N_13347);
and U18089 (N_18089,N_14009,N_14906);
or U18090 (N_18090,N_12895,N_14533);
and U18091 (N_18091,N_11152,N_14109);
xor U18092 (N_18092,N_10566,N_13720);
nand U18093 (N_18093,N_10554,N_14908);
nand U18094 (N_18094,N_13206,N_14487);
nand U18095 (N_18095,N_12644,N_14665);
nor U18096 (N_18096,N_10549,N_12317);
or U18097 (N_18097,N_14735,N_11731);
nand U18098 (N_18098,N_13012,N_12337);
and U18099 (N_18099,N_12567,N_12628);
xor U18100 (N_18100,N_11240,N_11527);
and U18101 (N_18101,N_10169,N_10999);
nor U18102 (N_18102,N_12543,N_12878);
or U18103 (N_18103,N_11755,N_11388);
xnor U18104 (N_18104,N_12127,N_14200);
and U18105 (N_18105,N_10406,N_13071);
nor U18106 (N_18106,N_13392,N_12942);
or U18107 (N_18107,N_11742,N_12075);
and U18108 (N_18108,N_12089,N_14041);
nor U18109 (N_18109,N_12265,N_10948);
or U18110 (N_18110,N_10454,N_10475);
or U18111 (N_18111,N_10299,N_10297);
or U18112 (N_18112,N_13837,N_11022);
or U18113 (N_18113,N_10444,N_14851);
nand U18114 (N_18114,N_10912,N_13770);
xor U18115 (N_18115,N_13797,N_10162);
nand U18116 (N_18116,N_12484,N_14635);
or U18117 (N_18117,N_11874,N_11610);
and U18118 (N_18118,N_13127,N_12128);
xor U18119 (N_18119,N_12806,N_11714);
or U18120 (N_18120,N_13826,N_14809);
and U18121 (N_18121,N_11570,N_10333);
or U18122 (N_18122,N_14838,N_10010);
or U18123 (N_18123,N_12834,N_10029);
or U18124 (N_18124,N_12363,N_13928);
nand U18125 (N_18125,N_13828,N_10775);
nor U18126 (N_18126,N_14943,N_14795);
and U18127 (N_18127,N_10914,N_14497);
and U18128 (N_18128,N_13126,N_11011);
nor U18129 (N_18129,N_13347,N_12990);
nand U18130 (N_18130,N_13578,N_14966);
nor U18131 (N_18131,N_14347,N_13009);
or U18132 (N_18132,N_11535,N_14834);
or U18133 (N_18133,N_11430,N_12664);
nor U18134 (N_18134,N_13009,N_12020);
nor U18135 (N_18135,N_11394,N_14005);
nand U18136 (N_18136,N_12418,N_11054);
xnor U18137 (N_18137,N_11868,N_11960);
nor U18138 (N_18138,N_10733,N_12246);
xnor U18139 (N_18139,N_11522,N_12481);
xnor U18140 (N_18140,N_13715,N_13757);
or U18141 (N_18141,N_14027,N_11790);
xnor U18142 (N_18142,N_11440,N_11954);
or U18143 (N_18143,N_14055,N_11950);
nand U18144 (N_18144,N_13249,N_10800);
and U18145 (N_18145,N_14116,N_11909);
nand U18146 (N_18146,N_10153,N_14701);
and U18147 (N_18147,N_14217,N_13249);
nand U18148 (N_18148,N_10830,N_14120);
xnor U18149 (N_18149,N_13056,N_14876);
nand U18150 (N_18150,N_14462,N_10222);
xor U18151 (N_18151,N_13856,N_13974);
nand U18152 (N_18152,N_10484,N_10879);
xnor U18153 (N_18153,N_13114,N_12508);
nor U18154 (N_18154,N_14762,N_13852);
and U18155 (N_18155,N_11995,N_11804);
nor U18156 (N_18156,N_14257,N_10846);
xnor U18157 (N_18157,N_10731,N_11348);
nor U18158 (N_18158,N_10674,N_12537);
nand U18159 (N_18159,N_11401,N_13078);
and U18160 (N_18160,N_13158,N_10489);
xor U18161 (N_18161,N_14105,N_11246);
and U18162 (N_18162,N_10956,N_10490);
or U18163 (N_18163,N_10146,N_12235);
and U18164 (N_18164,N_10171,N_11063);
and U18165 (N_18165,N_13331,N_10978);
nand U18166 (N_18166,N_13519,N_13648);
nor U18167 (N_18167,N_12643,N_10850);
nor U18168 (N_18168,N_11810,N_12408);
nor U18169 (N_18169,N_10911,N_14415);
and U18170 (N_18170,N_14684,N_12864);
or U18171 (N_18171,N_13645,N_14962);
and U18172 (N_18172,N_10550,N_11533);
xor U18173 (N_18173,N_11882,N_11985);
nor U18174 (N_18174,N_10092,N_11980);
xor U18175 (N_18175,N_14814,N_12435);
nand U18176 (N_18176,N_11189,N_12854);
nand U18177 (N_18177,N_14040,N_10027);
nor U18178 (N_18178,N_11584,N_10828);
nand U18179 (N_18179,N_13141,N_14072);
or U18180 (N_18180,N_14647,N_12764);
nand U18181 (N_18181,N_10951,N_14253);
xnor U18182 (N_18182,N_10159,N_11956);
and U18183 (N_18183,N_10254,N_12288);
xor U18184 (N_18184,N_10414,N_14457);
nor U18185 (N_18185,N_13690,N_10966);
and U18186 (N_18186,N_14220,N_12007);
or U18187 (N_18187,N_13758,N_11371);
or U18188 (N_18188,N_14827,N_11990);
xor U18189 (N_18189,N_13431,N_11179);
nor U18190 (N_18190,N_11098,N_14180);
and U18191 (N_18191,N_12942,N_12637);
xor U18192 (N_18192,N_13610,N_11513);
nand U18193 (N_18193,N_12163,N_13676);
or U18194 (N_18194,N_13855,N_10232);
xor U18195 (N_18195,N_11100,N_13165);
and U18196 (N_18196,N_13618,N_13610);
and U18197 (N_18197,N_10647,N_13007);
nand U18198 (N_18198,N_14613,N_14305);
and U18199 (N_18199,N_12889,N_14544);
nor U18200 (N_18200,N_13630,N_14805);
nand U18201 (N_18201,N_12974,N_13156);
nor U18202 (N_18202,N_11613,N_12034);
or U18203 (N_18203,N_13298,N_12241);
nor U18204 (N_18204,N_12169,N_14234);
and U18205 (N_18205,N_14460,N_13474);
nor U18206 (N_18206,N_14119,N_11310);
nor U18207 (N_18207,N_12292,N_10933);
nand U18208 (N_18208,N_14174,N_14302);
xnor U18209 (N_18209,N_12973,N_10881);
or U18210 (N_18210,N_11354,N_14606);
nor U18211 (N_18211,N_11987,N_14860);
or U18212 (N_18212,N_10895,N_14248);
nor U18213 (N_18213,N_10197,N_12078);
or U18214 (N_18214,N_11496,N_14882);
or U18215 (N_18215,N_13816,N_14161);
and U18216 (N_18216,N_12623,N_13243);
and U18217 (N_18217,N_13097,N_13523);
and U18218 (N_18218,N_13149,N_12392);
nand U18219 (N_18219,N_11661,N_10168);
and U18220 (N_18220,N_14997,N_11826);
nor U18221 (N_18221,N_12509,N_10678);
nor U18222 (N_18222,N_10775,N_14911);
nand U18223 (N_18223,N_12535,N_11893);
xor U18224 (N_18224,N_12678,N_11142);
xor U18225 (N_18225,N_13548,N_11696);
xor U18226 (N_18226,N_10690,N_10644);
nor U18227 (N_18227,N_10059,N_12084);
or U18228 (N_18228,N_11176,N_13949);
or U18229 (N_18229,N_11118,N_12539);
and U18230 (N_18230,N_13628,N_11349);
and U18231 (N_18231,N_12937,N_13962);
xnor U18232 (N_18232,N_13595,N_14224);
nor U18233 (N_18233,N_12183,N_12968);
nand U18234 (N_18234,N_11359,N_10302);
nor U18235 (N_18235,N_14714,N_13110);
and U18236 (N_18236,N_14996,N_14385);
or U18237 (N_18237,N_10077,N_14533);
and U18238 (N_18238,N_12620,N_11120);
nand U18239 (N_18239,N_12263,N_11999);
nand U18240 (N_18240,N_14626,N_13048);
nor U18241 (N_18241,N_14967,N_11720);
xnor U18242 (N_18242,N_13011,N_13155);
or U18243 (N_18243,N_10987,N_13377);
nand U18244 (N_18244,N_12102,N_13274);
nor U18245 (N_18245,N_10054,N_14465);
nor U18246 (N_18246,N_10366,N_13434);
and U18247 (N_18247,N_13334,N_10050);
nand U18248 (N_18248,N_14372,N_11874);
nand U18249 (N_18249,N_10056,N_12313);
or U18250 (N_18250,N_12007,N_10856);
or U18251 (N_18251,N_12596,N_13801);
nor U18252 (N_18252,N_11540,N_13181);
nor U18253 (N_18253,N_12731,N_14941);
xor U18254 (N_18254,N_12273,N_14788);
nor U18255 (N_18255,N_10157,N_14241);
or U18256 (N_18256,N_12500,N_13344);
nand U18257 (N_18257,N_11508,N_10662);
nor U18258 (N_18258,N_11388,N_10717);
or U18259 (N_18259,N_12982,N_12285);
xor U18260 (N_18260,N_14408,N_10735);
xor U18261 (N_18261,N_13441,N_14654);
xor U18262 (N_18262,N_11817,N_12538);
and U18263 (N_18263,N_11299,N_10928);
nor U18264 (N_18264,N_14410,N_11065);
or U18265 (N_18265,N_10433,N_14612);
nor U18266 (N_18266,N_10416,N_14668);
xor U18267 (N_18267,N_13806,N_11051);
or U18268 (N_18268,N_12793,N_14999);
and U18269 (N_18269,N_11057,N_14486);
nor U18270 (N_18270,N_13237,N_10638);
and U18271 (N_18271,N_13153,N_14969);
nand U18272 (N_18272,N_10572,N_12734);
nand U18273 (N_18273,N_10032,N_13068);
or U18274 (N_18274,N_11394,N_12097);
and U18275 (N_18275,N_12174,N_10858);
or U18276 (N_18276,N_12074,N_10302);
nor U18277 (N_18277,N_14745,N_14594);
xor U18278 (N_18278,N_11285,N_12500);
xor U18279 (N_18279,N_14731,N_14279);
or U18280 (N_18280,N_14036,N_10677);
xnor U18281 (N_18281,N_12807,N_10202);
nor U18282 (N_18282,N_11099,N_10207);
xnor U18283 (N_18283,N_13038,N_11049);
nand U18284 (N_18284,N_13420,N_10360);
and U18285 (N_18285,N_13260,N_10589);
and U18286 (N_18286,N_11275,N_12804);
nand U18287 (N_18287,N_12149,N_11699);
nor U18288 (N_18288,N_10598,N_10343);
and U18289 (N_18289,N_12410,N_12163);
nand U18290 (N_18290,N_11432,N_12335);
nor U18291 (N_18291,N_11545,N_13079);
nor U18292 (N_18292,N_14134,N_14506);
xnor U18293 (N_18293,N_12191,N_11623);
and U18294 (N_18294,N_12273,N_14820);
and U18295 (N_18295,N_14133,N_14166);
or U18296 (N_18296,N_12842,N_12379);
nor U18297 (N_18297,N_10063,N_14447);
and U18298 (N_18298,N_10497,N_14227);
and U18299 (N_18299,N_13460,N_11564);
or U18300 (N_18300,N_10236,N_12450);
nor U18301 (N_18301,N_14373,N_12490);
or U18302 (N_18302,N_12725,N_13284);
nor U18303 (N_18303,N_14811,N_10501);
or U18304 (N_18304,N_14598,N_13098);
or U18305 (N_18305,N_11169,N_11905);
xnor U18306 (N_18306,N_14613,N_11566);
nor U18307 (N_18307,N_11680,N_10922);
nor U18308 (N_18308,N_14141,N_11261);
nand U18309 (N_18309,N_12713,N_13592);
nand U18310 (N_18310,N_11397,N_13994);
or U18311 (N_18311,N_10520,N_12439);
nor U18312 (N_18312,N_14326,N_13438);
or U18313 (N_18313,N_13108,N_10113);
nor U18314 (N_18314,N_13973,N_14572);
nand U18315 (N_18315,N_14649,N_10793);
and U18316 (N_18316,N_13681,N_13994);
nand U18317 (N_18317,N_13461,N_12227);
nand U18318 (N_18318,N_12513,N_11146);
xnor U18319 (N_18319,N_14684,N_11999);
nor U18320 (N_18320,N_12872,N_10617);
or U18321 (N_18321,N_10432,N_10779);
or U18322 (N_18322,N_12274,N_12025);
nor U18323 (N_18323,N_11256,N_11996);
xnor U18324 (N_18324,N_11831,N_12957);
and U18325 (N_18325,N_12445,N_14492);
nor U18326 (N_18326,N_12517,N_13906);
nor U18327 (N_18327,N_12184,N_10214);
nor U18328 (N_18328,N_14095,N_10602);
and U18329 (N_18329,N_10736,N_11035);
nand U18330 (N_18330,N_12787,N_10886);
xor U18331 (N_18331,N_12065,N_11158);
and U18332 (N_18332,N_14202,N_11712);
nand U18333 (N_18333,N_14419,N_13947);
xor U18334 (N_18334,N_10643,N_12599);
nand U18335 (N_18335,N_12962,N_13339);
and U18336 (N_18336,N_12550,N_12089);
or U18337 (N_18337,N_13065,N_14710);
and U18338 (N_18338,N_13840,N_12036);
or U18339 (N_18339,N_12366,N_10939);
nand U18340 (N_18340,N_13283,N_12042);
xnor U18341 (N_18341,N_11157,N_14903);
xor U18342 (N_18342,N_11751,N_10218);
xnor U18343 (N_18343,N_11979,N_14683);
nor U18344 (N_18344,N_10032,N_10990);
and U18345 (N_18345,N_14626,N_10018);
or U18346 (N_18346,N_12283,N_14561);
xnor U18347 (N_18347,N_12068,N_11670);
xor U18348 (N_18348,N_12917,N_10063);
xnor U18349 (N_18349,N_13647,N_14393);
nor U18350 (N_18350,N_13399,N_11224);
xnor U18351 (N_18351,N_11133,N_12256);
and U18352 (N_18352,N_13681,N_13933);
xor U18353 (N_18353,N_14327,N_13595);
or U18354 (N_18354,N_10277,N_10245);
xnor U18355 (N_18355,N_13707,N_12409);
and U18356 (N_18356,N_11622,N_13933);
and U18357 (N_18357,N_10617,N_10840);
nand U18358 (N_18358,N_13837,N_10692);
and U18359 (N_18359,N_11331,N_10821);
nor U18360 (N_18360,N_12519,N_10791);
nor U18361 (N_18361,N_13314,N_10839);
nand U18362 (N_18362,N_11733,N_12909);
nor U18363 (N_18363,N_13569,N_10503);
or U18364 (N_18364,N_14827,N_10670);
or U18365 (N_18365,N_14720,N_12807);
or U18366 (N_18366,N_13028,N_13696);
nor U18367 (N_18367,N_13652,N_11561);
nor U18368 (N_18368,N_11065,N_14941);
nand U18369 (N_18369,N_14430,N_10285);
nand U18370 (N_18370,N_12033,N_10647);
or U18371 (N_18371,N_12454,N_10293);
or U18372 (N_18372,N_12265,N_11008);
nor U18373 (N_18373,N_14764,N_12081);
nand U18374 (N_18374,N_14454,N_13787);
or U18375 (N_18375,N_13280,N_10527);
or U18376 (N_18376,N_10509,N_13450);
or U18377 (N_18377,N_10834,N_12598);
nand U18378 (N_18378,N_13890,N_10531);
xnor U18379 (N_18379,N_12435,N_12051);
or U18380 (N_18380,N_11869,N_11253);
nand U18381 (N_18381,N_11250,N_13808);
and U18382 (N_18382,N_13232,N_12255);
or U18383 (N_18383,N_11158,N_10390);
and U18384 (N_18384,N_13789,N_10696);
nand U18385 (N_18385,N_13223,N_10366);
or U18386 (N_18386,N_11065,N_11212);
nand U18387 (N_18387,N_10617,N_14459);
nor U18388 (N_18388,N_12113,N_12175);
and U18389 (N_18389,N_11287,N_13606);
xnor U18390 (N_18390,N_13742,N_14944);
and U18391 (N_18391,N_14072,N_12636);
nor U18392 (N_18392,N_13156,N_10357);
nor U18393 (N_18393,N_11933,N_12119);
nand U18394 (N_18394,N_12012,N_11937);
nor U18395 (N_18395,N_10121,N_13564);
or U18396 (N_18396,N_10879,N_13809);
or U18397 (N_18397,N_14350,N_10861);
and U18398 (N_18398,N_12969,N_14196);
or U18399 (N_18399,N_14443,N_14800);
nand U18400 (N_18400,N_14709,N_12378);
nor U18401 (N_18401,N_12354,N_11591);
nand U18402 (N_18402,N_12256,N_13804);
xnor U18403 (N_18403,N_14140,N_10625);
nor U18404 (N_18404,N_11572,N_13313);
nand U18405 (N_18405,N_12194,N_10049);
and U18406 (N_18406,N_10413,N_14142);
and U18407 (N_18407,N_12388,N_10260);
and U18408 (N_18408,N_13221,N_12612);
xnor U18409 (N_18409,N_12437,N_12721);
and U18410 (N_18410,N_11010,N_11570);
or U18411 (N_18411,N_10974,N_14074);
nand U18412 (N_18412,N_12743,N_11968);
or U18413 (N_18413,N_10950,N_11656);
and U18414 (N_18414,N_13027,N_13053);
nor U18415 (N_18415,N_13418,N_10040);
nor U18416 (N_18416,N_13930,N_13185);
xor U18417 (N_18417,N_12576,N_13463);
nor U18418 (N_18418,N_13822,N_14963);
xnor U18419 (N_18419,N_13918,N_14440);
xor U18420 (N_18420,N_13684,N_13563);
nor U18421 (N_18421,N_13188,N_12460);
and U18422 (N_18422,N_12194,N_12609);
nand U18423 (N_18423,N_11940,N_14375);
nor U18424 (N_18424,N_10048,N_11039);
nand U18425 (N_18425,N_13371,N_14642);
nand U18426 (N_18426,N_10560,N_14467);
xor U18427 (N_18427,N_12761,N_13751);
nor U18428 (N_18428,N_11799,N_12338);
xnor U18429 (N_18429,N_13715,N_13143);
nor U18430 (N_18430,N_11667,N_10633);
or U18431 (N_18431,N_12881,N_10659);
nand U18432 (N_18432,N_10432,N_11609);
or U18433 (N_18433,N_12708,N_14592);
or U18434 (N_18434,N_13604,N_10643);
nand U18435 (N_18435,N_10113,N_14343);
or U18436 (N_18436,N_10216,N_10680);
xnor U18437 (N_18437,N_10263,N_10483);
or U18438 (N_18438,N_13024,N_11373);
xor U18439 (N_18439,N_11545,N_14747);
or U18440 (N_18440,N_11949,N_13785);
xor U18441 (N_18441,N_10622,N_12670);
xnor U18442 (N_18442,N_13994,N_14669);
or U18443 (N_18443,N_11047,N_11267);
nor U18444 (N_18444,N_12923,N_12506);
and U18445 (N_18445,N_12687,N_10180);
or U18446 (N_18446,N_10532,N_12125);
or U18447 (N_18447,N_10113,N_11003);
and U18448 (N_18448,N_13058,N_14906);
and U18449 (N_18449,N_11396,N_10257);
nor U18450 (N_18450,N_11858,N_10241);
nor U18451 (N_18451,N_12407,N_11515);
and U18452 (N_18452,N_12983,N_10263);
nor U18453 (N_18453,N_12875,N_13046);
nand U18454 (N_18454,N_12628,N_14841);
nand U18455 (N_18455,N_10036,N_11690);
and U18456 (N_18456,N_14999,N_13599);
nor U18457 (N_18457,N_14468,N_12876);
or U18458 (N_18458,N_12614,N_13631);
xnor U18459 (N_18459,N_12208,N_10555);
or U18460 (N_18460,N_11143,N_14515);
nor U18461 (N_18461,N_14072,N_12125);
and U18462 (N_18462,N_11738,N_11155);
and U18463 (N_18463,N_14992,N_11093);
nand U18464 (N_18464,N_11500,N_14245);
nor U18465 (N_18465,N_14247,N_13748);
nand U18466 (N_18466,N_13023,N_14484);
or U18467 (N_18467,N_14621,N_14285);
or U18468 (N_18468,N_13284,N_12456);
xnor U18469 (N_18469,N_11009,N_14583);
nor U18470 (N_18470,N_12853,N_10383);
or U18471 (N_18471,N_11651,N_14267);
nand U18472 (N_18472,N_12153,N_10489);
nand U18473 (N_18473,N_12874,N_10744);
nand U18474 (N_18474,N_11164,N_13297);
xor U18475 (N_18475,N_13211,N_11439);
or U18476 (N_18476,N_10524,N_10189);
xnor U18477 (N_18477,N_10255,N_10721);
nand U18478 (N_18478,N_13712,N_10370);
or U18479 (N_18479,N_11711,N_12051);
nor U18480 (N_18480,N_14999,N_11036);
xnor U18481 (N_18481,N_14155,N_14270);
nor U18482 (N_18482,N_14703,N_12510);
and U18483 (N_18483,N_14765,N_11071);
xor U18484 (N_18484,N_13181,N_11036);
nor U18485 (N_18485,N_11180,N_10081);
and U18486 (N_18486,N_12368,N_13164);
xnor U18487 (N_18487,N_13408,N_10833);
nor U18488 (N_18488,N_13614,N_13640);
nor U18489 (N_18489,N_12287,N_12740);
and U18490 (N_18490,N_12173,N_14626);
xor U18491 (N_18491,N_13065,N_12954);
nor U18492 (N_18492,N_11636,N_12385);
nor U18493 (N_18493,N_12257,N_11084);
and U18494 (N_18494,N_14899,N_10256);
nand U18495 (N_18495,N_12839,N_14335);
and U18496 (N_18496,N_10627,N_10995);
nand U18497 (N_18497,N_13759,N_14040);
nand U18498 (N_18498,N_10013,N_14265);
xnor U18499 (N_18499,N_14655,N_10296);
and U18500 (N_18500,N_11840,N_10769);
and U18501 (N_18501,N_13506,N_10280);
and U18502 (N_18502,N_11799,N_10303);
xnor U18503 (N_18503,N_11511,N_13037);
xnor U18504 (N_18504,N_13411,N_11849);
or U18505 (N_18505,N_10792,N_10056);
nor U18506 (N_18506,N_11091,N_12845);
or U18507 (N_18507,N_14278,N_12304);
and U18508 (N_18508,N_14207,N_11701);
or U18509 (N_18509,N_14817,N_12172);
and U18510 (N_18510,N_10819,N_13395);
and U18511 (N_18511,N_11794,N_12448);
nor U18512 (N_18512,N_10138,N_12090);
nor U18513 (N_18513,N_14996,N_11281);
or U18514 (N_18514,N_13074,N_12113);
or U18515 (N_18515,N_11850,N_14088);
nand U18516 (N_18516,N_12880,N_10517);
nor U18517 (N_18517,N_12545,N_10546);
or U18518 (N_18518,N_13232,N_11473);
and U18519 (N_18519,N_10627,N_10844);
and U18520 (N_18520,N_10660,N_11524);
and U18521 (N_18521,N_10404,N_10633);
nand U18522 (N_18522,N_12797,N_14050);
nor U18523 (N_18523,N_11426,N_10742);
xor U18524 (N_18524,N_11773,N_12845);
xnor U18525 (N_18525,N_10959,N_10359);
or U18526 (N_18526,N_14430,N_13095);
or U18527 (N_18527,N_12306,N_10428);
nor U18528 (N_18528,N_11312,N_14263);
nor U18529 (N_18529,N_10901,N_10521);
or U18530 (N_18530,N_13964,N_11557);
nor U18531 (N_18531,N_12204,N_10624);
or U18532 (N_18532,N_14108,N_14458);
or U18533 (N_18533,N_10945,N_12765);
xor U18534 (N_18534,N_10203,N_13885);
and U18535 (N_18535,N_13517,N_10143);
and U18536 (N_18536,N_14444,N_12954);
xor U18537 (N_18537,N_11956,N_13171);
and U18538 (N_18538,N_11297,N_12603);
nor U18539 (N_18539,N_12255,N_14173);
xor U18540 (N_18540,N_10738,N_11290);
and U18541 (N_18541,N_14863,N_14182);
nand U18542 (N_18542,N_11756,N_13219);
nand U18543 (N_18543,N_12294,N_12998);
nor U18544 (N_18544,N_14255,N_13180);
or U18545 (N_18545,N_12915,N_14607);
nor U18546 (N_18546,N_13571,N_14795);
or U18547 (N_18547,N_11213,N_14717);
xor U18548 (N_18548,N_10152,N_10730);
or U18549 (N_18549,N_14608,N_11179);
and U18550 (N_18550,N_13584,N_12788);
and U18551 (N_18551,N_13314,N_13268);
xnor U18552 (N_18552,N_13139,N_14681);
nor U18553 (N_18553,N_12166,N_11643);
nor U18554 (N_18554,N_11892,N_14641);
nor U18555 (N_18555,N_14348,N_11739);
nand U18556 (N_18556,N_11647,N_10354);
xor U18557 (N_18557,N_14399,N_10744);
xor U18558 (N_18558,N_14654,N_14857);
and U18559 (N_18559,N_12809,N_14893);
or U18560 (N_18560,N_14151,N_11675);
nor U18561 (N_18561,N_12495,N_12703);
nor U18562 (N_18562,N_10272,N_11797);
nor U18563 (N_18563,N_11515,N_13394);
nand U18564 (N_18564,N_11763,N_12194);
and U18565 (N_18565,N_12730,N_12181);
nand U18566 (N_18566,N_13104,N_11824);
or U18567 (N_18567,N_13370,N_10289);
xor U18568 (N_18568,N_10530,N_12237);
xnor U18569 (N_18569,N_11836,N_10199);
nor U18570 (N_18570,N_14471,N_11776);
xor U18571 (N_18571,N_14351,N_10714);
nor U18572 (N_18572,N_12950,N_14730);
nand U18573 (N_18573,N_11315,N_10162);
and U18574 (N_18574,N_14653,N_11172);
xor U18575 (N_18575,N_14965,N_12939);
nor U18576 (N_18576,N_13443,N_13127);
nand U18577 (N_18577,N_12190,N_14890);
nor U18578 (N_18578,N_13191,N_11884);
nor U18579 (N_18579,N_12815,N_13549);
xor U18580 (N_18580,N_10270,N_10137);
nand U18581 (N_18581,N_13995,N_14970);
xnor U18582 (N_18582,N_10595,N_13108);
xnor U18583 (N_18583,N_12951,N_14954);
and U18584 (N_18584,N_12778,N_12676);
and U18585 (N_18585,N_14594,N_13645);
or U18586 (N_18586,N_10643,N_10537);
xnor U18587 (N_18587,N_13949,N_14362);
nor U18588 (N_18588,N_12106,N_12335);
nor U18589 (N_18589,N_13493,N_13924);
nor U18590 (N_18590,N_12267,N_11138);
nor U18591 (N_18591,N_14814,N_14195);
nor U18592 (N_18592,N_10034,N_13789);
or U18593 (N_18593,N_12323,N_10350);
and U18594 (N_18594,N_10292,N_11417);
nand U18595 (N_18595,N_13671,N_14005);
xor U18596 (N_18596,N_13768,N_12177);
and U18597 (N_18597,N_13585,N_11496);
nor U18598 (N_18598,N_13948,N_13554);
or U18599 (N_18599,N_13123,N_11870);
nor U18600 (N_18600,N_13511,N_13344);
and U18601 (N_18601,N_13758,N_14180);
xnor U18602 (N_18602,N_14721,N_14398);
nor U18603 (N_18603,N_13021,N_10094);
nor U18604 (N_18604,N_11449,N_13779);
nor U18605 (N_18605,N_10924,N_14386);
nand U18606 (N_18606,N_12871,N_13148);
nand U18607 (N_18607,N_10600,N_12435);
or U18608 (N_18608,N_11010,N_10738);
and U18609 (N_18609,N_11971,N_12709);
nor U18610 (N_18610,N_10455,N_12670);
nand U18611 (N_18611,N_11309,N_14580);
and U18612 (N_18612,N_14864,N_11739);
and U18613 (N_18613,N_12127,N_10267);
nand U18614 (N_18614,N_10365,N_11371);
or U18615 (N_18615,N_14285,N_10632);
or U18616 (N_18616,N_14769,N_12517);
and U18617 (N_18617,N_10567,N_13073);
and U18618 (N_18618,N_11447,N_13127);
nand U18619 (N_18619,N_13455,N_13683);
and U18620 (N_18620,N_10171,N_13545);
nor U18621 (N_18621,N_10452,N_12387);
nand U18622 (N_18622,N_13290,N_13065);
or U18623 (N_18623,N_10938,N_13959);
nand U18624 (N_18624,N_12435,N_11315);
and U18625 (N_18625,N_11453,N_10346);
nor U18626 (N_18626,N_14652,N_14829);
xnor U18627 (N_18627,N_10437,N_11332);
nor U18628 (N_18628,N_14526,N_10009);
or U18629 (N_18629,N_12937,N_14405);
xnor U18630 (N_18630,N_12553,N_11530);
xnor U18631 (N_18631,N_14484,N_11431);
nand U18632 (N_18632,N_13786,N_12971);
nor U18633 (N_18633,N_10583,N_12925);
xor U18634 (N_18634,N_10643,N_12462);
and U18635 (N_18635,N_12665,N_14327);
nor U18636 (N_18636,N_13474,N_10621);
xor U18637 (N_18637,N_12989,N_11251);
nor U18638 (N_18638,N_14903,N_11635);
nand U18639 (N_18639,N_10010,N_14796);
or U18640 (N_18640,N_13857,N_11415);
and U18641 (N_18641,N_14240,N_12715);
xor U18642 (N_18642,N_13610,N_13289);
nand U18643 (N_18643,N_10036,N_10531);
nor U18644 (N_18644,N_12172,N_14984);
or U18645 (N_18645,N_11247,N_14075);
xnor U18646 (N_18646,N_11670,N_12472);
nand U18647 (N_18647,N_11039,N_13309);
nand U18648 (N_18648,N_12020,N_12183);
nor U18649 (N_18649,N_12410,N_11778);
and U18650 (N_18650,N_10639,N_11138);
and U18651 (N_18651,N_12269,N_12523);
nor U18652 (N_18652,N_13089,N_10890);
nor U18653 (N_18653,N_11383,N_14132);
nand U18654 (N_18654,N_10640,N_14028);
nor U18655 (N_18655,N_12277,N_14865);
xnor U18656 (N_18656,N_13868,N_13277);
xor U18657 (N_18657,N_14870,N_14756);
and U18658 (N_18658,N_10877,N_10114);
nand U18659 (N_18659,N_14922,N_11516);
xor U18660 (N_18660,N_14734,N_14281);
and U18661 (N_18661,N_11259,N_14259);
and U18662 (N_18662,N_11947,N_10271);
xor U18663 (N_18663,N_13310,N_14442);
nor U18664 (N_18664,N_13673,N_12913);
nand U18665 (N_18665,N_13138,N_12048);
and U18666 (N_18666,N_14073,N_10584);
and U18667 (N_18667,N_10401,N_12975);
nor U18668 (N_18668,N_14538,N_12989);
xor U18669 (N_18669,N_11768,N_11870);
nor U18670 (N_18670,N_13497,N_11261);
or U18671 (N_18671,N_11809,N_12202);
or U18672 (N_18672,N_12113,N_10631);
and U18673 (N_18673,N_11257,N_13526);
nand U18674 (N_18674,N_13242,N_11341);
nor U18675 (N_18675,N_12022,N_14320);
xnor U18676 (N_18676,N_12265,N_11596);
nand U18677 (N_18677,N_12831,N_12039);
nor U18678 (N_18678,N_10775,N_14837);
nor U18679 (N_18679,N_11110,N_11426);
and U18680 (N_18680,N_14962,N_11758);
or U18681 (N_18681,N_13298,N_12982);
nand U18682 (N_18682,N_12670,N_13545);
and U18683 (N_18683,N_14773,N_11662);
or U18684 (N_18684,N_12102,N_10967);
nand U18685 (N_18685,N_14714,N_14156);
and U18686 (N_18686,N_12609,N_10967);
nor U18687 (N_18687,N_12844,N_12173);
nand U18688 (N_18688,N_14926,N_10387);
nand U18689 (N_18689,N_10012,N_10236);
nor U18690 (N_18690,N_14650,N_14793);
nand U18691 (N_18691,N_12288,N_10120);
and U18692 (N_18692,N_10984,N_13177);
nand U18693 (N_18693,N_11860,N_12956);
nor U18694 (N_18694,N_12453,N_14296);
and U18695 (N_18695,N_13491,N_11505);
nand U18696 (N_18696,N_14538,N_10675);
nand U18697 (N_18697,N_14575,N_11536);
nor U18698 (N_18698,N_10177,N_14369);
nand U18699 (N_18699,N_13048,N_13125);
nand U18700 (N_18700,N_13966,N_14561);
nor U18701 (N_18701,N_13999,N_13653);
nor U18702 (N_18702,N_10446,N_10576);
nand U18703 (N_18703,N_10634,N_14106);
nand U18704 (N_18704,N_10705,N_11650);
and U18705 (N_18705,N_11591,N_12865);
or U18706 (N_18706,N_12097,N_10239);
and U18707 (N_18707,N_14010,N_10681);
and U18708 (N_18708,N_10449,N_11390);
and U18709 (N_18709,N_14984,N_13060);
nor U18710 (N_18710,N_10761,N_13213);
nand U18711 (N_18711,N_12828,N_10531);
xor U18712 (N_18712,N_11933,N_11117);
nor U18713 (N_18713,N_14902,N_10150);
nand U18714 (N_18714,N_14366,N_11639);
nor U18715 (N_18715,N_12109,N_13962);
and U18716 (N_18716,N_11650,N_12993);
and U18717 (N_18717,N_11027,N_13414);
nor U18718 (N_18718,N_14421,N_10804);
xor U18719 (N_18719,N_11733,N_14287);
or U18720 (N_18720,N_10997,N_14964);
nor U18721 (N_18721,N_14163,N_12911);
xnor U18722 (N_18722,N_10584,N_10588);
or U18723 (N_18723,N_12263,N_11257);
xor U18724 (N_18724,N_11266,N_12526);
or U18725 (N_18725,N_13259,N_10171);
nor U18726 (N_18726,N_12736,N_11433);
xor U18727 (N_18727,N_14250,N_14132);
nand U18728 (N_18728,N_14450,N_14389);
and U18729 (N_18729,N_10426,N_11088);
or U18730 (N_18730,N_14213,N_13060);
nand U18731 (N_18731,N_13495,N_10220);
nor U18732 (N_18732,N_14954,N_12021);
nor U18733 (N_18733,N_10067,N_13177);
and U18734 (N_18734,N_12074,N_12452);
and U18735 (N_18735,N_10876,N_14235);
xor U18736 (N_18736,N_12769,N_11079);
nor U18737 (N_18737,N_13544,N_11242);
nand U18738 (N_18738,N_14141,N_10440);
nor U18739 (N_18739,N_14268,N_14819);
and U18740 (N_18740,N_11755,N_13275);
or U18741 (N_18741,N_10614,N_11827);
xnor U18742 (N_18742,N_10189,N_12313);
or U18743 (N_18743,N_14566,N_11148);
nor U18744 (N_18744,N_10779,N_11804);
and U18745 (N_18745,N_12369,N_12232);
nor U18746 (N_18746,N_14914,N_10672);
nand U18747 (N_18747,N_10920,N_13016);
or U18748 (N_18748,N_10097,N_13969);
or U18749 (N_18749,N_12771,N_10457);
and U18750 (N_18750,N_12750,N_14568);
xor U18751 (N_18751,N_10923,N_14899);
nor U18752 (N_18752,N_11029,N_13297);
xnor U18753 (N_18753,N_13619,N_14325);
and U18754 (N_18754,N_11810,N_13411);
and U18755 (N_18755,N_10724,N_10548);
nand U18756 (N_18756,N_13085,N_14405);
and U18757 (N_18757,N_12830,N_14308);
nand U18758 (N_18758,N_12795,N_14805);
xnor U18759 (N_18759,N_13604,N_10607);
nand U18760 (N_18760,N_10261,N_13768);
and U18761 (N_18761,N_14749,N_13977);
nand U18762 (N_18762,N_13914,N_14990);
or U18763 (N_18763,N_10003,N_11119);
nor U18764 (N_18764,N_10468,N_14084);
nor U18765 (N_18765,N_13275,N_12419);
and U18766 (N_18766,N_10048,N_12480);
or U18767 (N_18767,N_13621,N_10881);
or U18768 (N_18768,N_10676,N_10624);
and U18769 (N_18769,N_11005,N_14775);
xnor U18770 (N_18770,N_10944,N_10085);
xnor U18771 (N_18771,N_11604,N_12257);
and U18772 (N_18772,N_10042,N_12117);
or U18773 (N_18773,N_11313,N_14200);
or U18774 (N_18774,N_12912,N_10341);
nand U18775 (N_18775,N_12274,N_14408);
nor U18776 (N_18776,N_13805,N_12942);
nor U18777 (N_18777,N_10924,N_13805);
xor U18778 (N_18778,N_12792,N_11973);
xor U18779 (N_18779,N_13500,N_10555);
nand U18780 (N_18780,N_13180,N_10905);
and U18781 (N_18781,N_12584,N_13529);
or U18782 (N_18782,N_12430,N_14445);
nand U18783 (N_18783,N_12796,N_12482);
and U18784 (N_18784,N_12984,N_12879);
and U18785 (N_18785,N_11051,N_11552);
nor U18786 (N_18786,N_12188,N_14186);
nand U18787 (N_18787,N_12557,N_14722);
nand U18788 (N_18788,N_14562,N_10832);
nor U18789 (N_18789,N_13103,N_12390);
and U18790 (N_18790,N_10023,N_10661);
or U18791 (N_18791,N_12592,N_11345);
nand U18792 (N_18792,N_13810,N_11690);
nand U18793 (N_18793,N_11777,N_13074);
nor U18794 (N_18794,N_13982,N_10107);
or U18795 (N_18795,N_12068,N_13449);
and U18796 (N_18796,N_13568,N_10421);
nor U18797 (N_18797,N_11354,N_11014);
and U18798 (N_18798,N_11036,N_13841);
nor U18799 (N_18799,N_14347,N_13526);
or U18800 (N_18800,N_14779,N_11423);
and U18801 (N_18801,N_13549,N_14973);
or U18802 (N_18802,N_12468,N_14965);
and U18803 (N_18803,N_11466,N_13651);
nand U18804 (N_18804,N_12606,N_10341);
nand U18805 (N_18805,N_14194,N_12723);
xor U18806 (N_18806,N_12527,N_10224);
nand U18807 (N_18807,N_13037,N_10479);
nor U18808 (N_18808,N_14744,N_11280);
or U18809 (N_18809,N_10338,N_10165);
xnor U18810 (N_18810,N_10300,N_11043);
nand U18811 (N_18811,N_11341,N_12903);
nor U18812 (N_18812,N_11560,N_10247);
or U18813 (N_18813,N_14687,N_13658);
or U18814 (N_18814,N_10162,N_14420);
and U18815 (N_18815,N_11199,N_11072);
and U18816 (N_18816,N_11416,N_14825);
and U18817 (N_18817,N_10052,N_10733);
and U18818 (N_18818,N_14776,N_12958);
nor U18819 (N_18819,N_11975,N_14135);
or U18820 (N_18820,N_10234,N_13862);
and U18821 (N_18821,N_11255,N_13288);
xor U18822 (N_18822,N_10094,N_13549);
and U18823 (N_18823,N_13325,N_10548);
nand U18824 (N_18824,N_10776,N_13157);
and U18825 (N_18825,N_10548,N_10715);
and U18826 (N_18826,N_13676,N_12653);
nor U18827 (N_18827,N_10116,N_12905);
and U18828 (N_18828,N_14000,N_14396);
xnor U18829 (N_18829,N_12106,N_14517);
nand U18830 (N_18830,N_13704,N_14775);
or U18831 (N_18831,N_12550,N_14571);
nor U18832 (N_18832,N_14745,N_10159);
and U18833 (N_18833,N_14097,N_12218);
xnor U18834 (N_18834,N_13940,N_14432);
nand U18835 (N_18835,N_11652,N_11953);
nand U18836 (N_18836,N_12007,N_12928);
nand U18837 (N_18837,N_12523,N_12372);
or U18838 (N_18838,N_13111,N_10081);
nor U18839 (N_18839,N_10173,N_12381);
nor U18840 (N_18840,N_10920,N_10905);
xor U18841 (N_18841,N_13690,N_14970);
nor U18842 (N_18842,N_10256,N_10539);
xnor U18843 (N_18843,N_13471,N_11243);
or U18844 (N_18844,N_14383,N_10154);
nor U18845 (N_18845,N_10390,N_13761);
and U18846 (N_18846,N_11219,N_14819);
or U18847 (N_18847,N_10834,N_12223);
xor U18848 (N_18848,N_10086,N_11720);
xor U18849 (N_18849,N_12366,N_12995);
xnor U18850 (N_18850,N_10224,N_14460);
or U18851 (N_18851,N_13056,N_14873);
xnor U18852 (N_18852,N_14141,N_11075);
nand U18853 (N_18853,N_12532,N_10035);
and U18854 (N_18854,N_10819,N_10004);
xnor U18855 (N_18855,N_10974,N_14542);
nand U18856 (N_18856,N_14343,N_11526);
xnor U18857 (N_18857,N_10265,N_14231);
and U18858 (N_18858,N_14283,N_14747);
xor U18859 (N_18859,N_14179,N_12857);
xnor U18860 (N_18860,N_11306,N_13775);
nand U18861 (N_18861,N_11252,N_10006);
and U18862 (N_18862,N_12029,N_13823);
xor U18863 (N_18863,N_14388,N_12775);
nor U18864 (N_18864,N_12992,N_11966);
xnor U18865 (N_18865,N_14622,N_14388);
nor U18866 (N_18866,N_13188,N_10242);
nand U18867 (N_18867,N_14045,N_11405);
nor U18868 (N_18868,N_10654,N_13772);
nor U18869 (N_18869,N_14593,N_11337);
nand U18870 (N_18870,N_14817,N_13274);
or U18871 (N_18871,N_10564,N_12899);
nand U18872 (N_18872,N_12551,N_12382);
and U18873 (N_18873,N_10221,N_10433);
nor U18874 (N_18874,N_11971,N_14451);
or U18875 (N_18875,N_11439,N_13711);
nand U18876 (N_18876,N_12421,N_11435);
nor U18877 (N_18877,N_11834,N_12114);
nand U18878 (N_18878,N_11494,N_11013);
or U18879 (N_18879,N_11349,N_11429);
and U18880 (N_18880,N_10092,N_11061);
nor U18881 (N_18881,N_12466,N_13499);
nor U18882 (N_18882,N_10091,N_13098);
nor U18883 (N_18883,N_14602,N_13278);
xor U18884 (N_18884,N_10811,N_12210);
or U18885 (N_18885,N_13956,N_12459);
and U18886 (N_18886,N_12314,N_13934);
or U18887 (N_18887,N_12507,N_14768);
xnor U18888 (N_18888,N_12291,N_11190);
nor U18889 (N_18889,N_11852,N_10477);
or U18890 (N_18890,N_11501,N_12964);
xnor U18891 (N_18891,N_11838,N_11088);
nand U18892 (N_18892,N_11160,N_14336);
nand U18893 (N_18893,N_13191,N_14656);
or U18894 (N_18894,N_14262,N_13962);
or U18895 (N_18895,N_11156,N_10751);
or U18896 (N_18896,N_11993,N_12371);
nor U18897 (N_18897,N_14307,N_13186);
and U18898 (N_18898,N_13728,N_10183);
xor U18899 (N_18899,N_10946,N_10939);
and U18900 (N_18900,N_11861,N_12438);
xnor U18901 (N_18901,N_14511,N_14290);
nor U18902 (N_18902,N_14824,N_12519);
nand U18903 (N_18903,N_10261,N_10860);
and U18904 (N_18904,N_13920,N_11242);
nor U18905 (N_18905,N_10521,N_13271);
xnor U18906 (N_18906,N_10596,N_10910);
nand U18907 (N_18907,N_10877,N_12523);
nor U18908 (N_18908,N_12483,N_12305);
nor U18909 (N_18909,N_12504,N_10623);
nor U18910 (N_18910,N_14918,N_11179);
xnor U18911 (N_18911,N_11299,N_12879);
nand U18912 (N_18912,N_13957,N_12246);
xor U18913 (N_18913,N_13855,N_10189);
xor U18914 (N_18914,N_12431,N_14154);
nor U18915 (N_18915,N_12221,N_10885);
nor U18916 (N_18916,N_14717,N_12201);
or U18917 (N_18917,N_12105,N_14039);
and U18918 (N_18918,N_12438,N_11578);
nand U18919 (N_18919,N_10297,N_13903);
nand U18920 (N_18920,N_14121,N_10745);
or U18921 (N_18921,N_14071,N_11685);
nor U18922 (N_18922,N_10528,N_14753);
xor U18923 (N_18923,N_11261,N_13392);
xnor U18924 (N_18924,N_12544,N_10776);
nor U18925 (N_18925,N_10374,N_14277);
or U18926 (N_18926,N_14852,N_14124);
and U18927 (N_18927,N_13568,N_11230);
nand U18928 (N_18928,N_10903,N_14733);
xnor U18929 (N_18929,N_10799,N_11167);
or U18930 (N_18930,N_11592,N_10987);
nor U18931 (N_18931,N_13718,N_11912);
and U18932 (N_18932,N_14841,N_12317);
nand U18933 (N_18933,N_12457,N_13097);
and U18934 (N_18934,N_13045,N_10324);
nand U18935 (N_18935,N_13103,N_13154);
nor U18936 (N_18936,N_10663,N_11413);
xor U18937 (N_18937,N_14165,N_13693);
and U18938 (N_18938,N_12700,N_10185);
xnor U18939 (N_18939,N_14012,N_10937);
nor U18940 (N_18940,N_13892,N_14167);
nor U18941 (N_18941,N_10138,N_12271);
xnor U18942 (N_18942,N_12388,N_13022);
xnor U18943 (N_18943,N_10035,N_13463);
nor U18944 (N_18944,N_13129,N_11466);
or U18945 (N_18945,N_14705,N_11459);
xor U18946 (N_18946,N_10592,N_14139);
and U18947 (N_18947,N_10813,N_14764);
xnor U18948 (N_18948,N_11803,N_12105);
nor U18949 (N_18949,N_12898,N_14113);
nor U18950 (N_18950,N_14122,N_13970);
or U18951 (N_18951,N_14008,N_10712);
xnor U18952 (N_18952,N_14428,N_10107);
nor U18953 (N_18953,N_11788,N_14695);
or U18954 (N_18954,N_13734,N_11674);
xor U18955 (N_18955,N_10009,N_11394);
nor U18956 (N_18956,N_13136,N_10165);
and U18957 (N_18957,N_12926,N_11756);
nor U18958 (N_18958,N_14861,N_12553);
nand U18959 (N_18959,N_14899,N_11338);
and U18960 (N_18960,N_11484,N_13817);
nand U18961 (N_18961,N_14193,N_11893);
nand U18962 (N_18962,N_14272,N_11951);
and U18963 (N_18963,N_13176,N_14783);
and U18964 (N_18964,N_10743,N_14108);
or U18965 (N_18965,N_12780,N_14196);
nand U18966 (N_18966,N_14800,N_13859);
xor U18967 (N_18967,N_11825,N_12360);
and U18968 (N_18968,N_13605,N_12560);
nand U18969 (N_18969,N_14976,N_14113);
nand U18970 (N_18970,N_11228,N_14563);
and U18971 (N_18971,N_14654,N_13752);
nand U18972 (N_18972,N_13055,N_14034);
nand U18973 (N_18973,N_11501,N_13016);
or U18974 (N_18974,N_10717,N_13112);
nor U18975 (N_18975,N_14822,N_11762);
nor U18976 (N_18976,N_14722,N_13068);
or U18977 (N_18977,N_14785,N_14052);
and U18978 (N_18978,N_11648,N_12494);
nand U18979 (N_18979,N_14664,N_13612);
nand U18980 (N_18980,N_12572,N_12190);
xnor U18981 (N_18981,N_11256,N_11841);
xnor U18982 (N_18982,N_10568,N_12231);
nand U18983 (N_18983,N_10472,N_13578);
nand U18984 (N_18984,N_12366,N_13795);
nand U18985 (N_18985,N_10652,N_14328);
and U18986 (N_18986,N_13632,N_10198);
or U18987 (N_18987,N_10712,N_12711);
and U18988 (N_18988,N_13082,N_11704);
and U18989 (N_18989,N_10071,N_11524);
nand U18990 (N_18990,N_10748,N_14493);
nand U18991 (N_18991,N_12819,N_12290);
nor U18992 (N_18992,N_10621,N_10000);
and U18993 (N_18993,N_12502,N_11417);
xor U18994 (N_18994,N_14635,N_12795);
and U18995 (N_18995,N_14436,N_13316);
xor U18996 (N_18996,N_14288,N_14075);
nand U18997 (N_18997,N_10845,N_12730);
nor U18998 (N_18998,N_14263,N_12742);
and U18999 (N_18999,N_11624,N_11472);
or U19000 (N_19000,N_11573,N_14177);
nor U19001 (N_19001,N_12219,N_12132);
nor U19002 (N_19002,N_12160,N_13042);
and U19003 (N_19003,N_14698,N_10960);
nand U19004 (N_19004,N_11014,N_11105);
or U19005 (N_19005,N_12577,N_13944);
nor U19006 (N_19006,N_10012,N_13795);
and U19007 (N_19007,N_10702,N_12276);
and U19008 (N_19008,N_14848,N_14194);
xor U19009 (N_19009,N_13674,N_13795);
nor U19010 (N_19010,N_14684,N_14811);
nor U19011 (N_19011,N_12974,N_10031);
xor U19012 (N_19012,N_11997,N_14784);
nand U19013 (N_19013,N_12827,N_13918);
xnor U19014 (N_19014,N_11696,N_11298);
and U19015 (N_19015,N_11406,N_12053);
nand U19016 (N_19016,N_10273,N_11070);
and U19017 (N_19017,N_14195,N_11997);
or U19018 (N_19018,N_13747,N_13634);
and U19019 (N_19019,N_11420,N_14204);
xnor U19020 (N_19020,N_11522,N_11729);
xor U19021 (N_19021,N_13534,N_12128);
or U19022 (N_19022,N_13611,N_12335);
and U19023 (N_19023,N_10857,N_13818);
nor U19024 (N_19024,N_14468,N_13730);
nand U19025 (N_19025,N_11225,N_13203);
and U19026 (N_19026,N_11495,N_13525);
and U19027 (N_19027,N_14044,N_14179);
nand U19028 (N_19028,N_13583,N_13922);
or U19029 (N_19029,N_13113,N_12342);
or U19030 (N_19030,N_14332,N_11034);
and U19031 (N_19031,N_12823,N_13903);
xor U19032 (N_19032,N_11502,N_13433);
nand U19033 (N_19033,N_13543,N_14168);
xnor U19034 (N_19034,N_13607,N_14002);
nand U19035 (N_19035,N_12656,N_11193);
or U19036 (N_19036,N_13737,N_11568);
nand U19037 (N_19037,N_11343,N_10228);
nand U19038 (N_19038,N_12925,N_11721);
xor U19039 (N_19039,N_11128,N_14121);
nand U19040 (N_19040,N_14769,N_14694);
or U19041 (N_19041,N_11181,N_11238);
and U19042 (N_19042,N_11383,N_11713);
nand U19043 (N_19043,N_10212,N_13239);
nor U19044 (N_19044,N_10452,N_11254);
nor U19045 (N_19045,N_11416,N_11608);
xor U19046 (N_19046,N_14731,N_10874);
and U19047 (N_19047,N_13390,N_12168);
or U19048 (N_19048,N_10834,N_10236);
xnor U19049 (N_19049,N_13168,N_10269);
nand U19050 (N_19050,N_10360,N_12215);
and U19051 (N_19051,N_11905,N_14459);
nor U19052 (N_19052,N_13751,N_14010);
nand U19053 (N_19053,N_13474,N_13730);
or U19054 (N_19054,N_14742,N_13924);
and U19055 (N_19055,N_10339,N_10627);
xor U19056 (N_19056,N_14222,N_13900);
or U19057 (N_19057,N_12172,N_12163);
nand U19058 (N_19058,N_14434,N_14090);
nor U19059 (N_19059,N_10253,N_12733);
nor U19060 (N_19060,N_11474,N_11531);
xor U19061 (N_19061,N_14679,N_14087);
nor U19062 (N_19062,N_10253,N_12528);
nor U19063 (N_19063,N_12347,N_12295);
and U19064 (N_19064,N_11117,N_13005);
or U19065 (N_19065,N_12247,N_13295);
or U19066 (N_19066,N_10592,N_12577);
nand U19067 (N_19067,N_11011,N_11476);
or U19068 (N_19068,N_11232,N_14230);
nor U19069 (N_19069,N_12729,N_11097);
xor U19070 (N_19070,N_10195,N_11542);
nor U19071 (N_19071,N_11429,N_14939);
xor U19072 (N_19072,N_10962,N_14221);
xor U19073 (N_19073,N_13343,N_10109);
or U19074 (N_19074,N_11661,N_12909);
and U19075 (N_19075,N_14343,N_13299);
nor U19076 (N_19076,N_13626,N_11250);
xnor U19077 (N_19077,N_14421,N_12178);
nand U19078 (N_19078,N_14690,N_12775);
and U19079 (N_19079,N_12743,N_11889);
or U19080 (N_19080,N_11167,N_14432);
nand U19081 (N_19081,N_12352,N_13394);
nand U19082 (N_19082,N_11426,N_11506);
and U19083 (N_19083,N_11879,N_14649);
xnor U19084 (N_19084,N_11289,N_13308);
nand U19085 (N_19085,N_12602,N_11770);
and U19086 (N_19086,N_10263,N_14470);
nor U19087 (N_19087,N_12660,N_13603);
xor U19088 (N_19088,N_10967,N_10727);
or U19089 (N_19089,N_11696,N_11795);
or U19090 (N_19090,N_14058,N_11491);
nor U19091 (N_19091,N_14432,N_13345);
nand U19092 (N_19092,N_14393,N_13390);
xor U19093 (N_19093,N_10608,N_11556);
nor U19094 (N_19094,N_11237,N_11400);
or U19095 (N_19095,N_13605,N_13407);
or U19096 (N_19096,N_14541,N_13588);
or U19097 (N_19097,N_11455,N_14504);
xor U19098 (N_19098,N_11735,N_14419);
or U19099 (N_19099,N_12040,N_12395);
nor U19100 (N_19100,N_10086,N_12104);
and U19101 (N_19101,N_10787,N_14405);
and U19102 (N_19102,N_13212,N_11883);
xnor U19103 (N_19103,N_12439,N_11433);
xnor U19104 (N_19104,N_13907,N_14071);
xor U19105 (N_19105,N_10204,N_10757);
and U19106 (N_19106,N_12215,N_10466);
or U19107 (N_19107,N_13627,N_11206);
or U19108 (N_19108,N_14109,N_11904);
nor U19109 (N_19109,N_12653,N_11933);
xnor U19110 (N_19110,N_10279,N_14781);
nand U19111 (N_19111,N_14872,N_11191);
or U19112 (N_19112,N_14949,N_13747);
and U19113 (N_19113,N_14402,N_12041);
xnor U19114 (N_19114,N_12707,N_10499);
or U19115 (N_19115,N_14058,N_10976);
and U19116 (N_19116,N_10121,N_10147);
or U19117 (N_19117,N_10403,N_13273);
xnor U19118 (N_19118,N_13523,N_14644);
xor U19119 (N_19119,N_12421,N_10423);
nand U19120 (N_19120,N_12425,N_12829);
nand U19121 (N_19121,N_13210,N_10473);
xnor U19122 (N_19122,N_10371,N_14666);
and U19123 (N_19123,N_10655,N_11638);
nand U19124 (N_19124,N_13822,N_12719);
and U19125 (N_19125,N_14033,N_14975);
xnor U19126 (N_19126,N_13582,N_11896);
nor U19127 (N_19127,N_11270,N_13902);
xor U19128 (N_19128,N_14069,N_12924);
and U19129 (N_19129,N_14378,N_14882);
and U19130 (N_19130,N_11029,N_13073);
and U19131 (N_19131,N_11946,N_11027);
xor U19132 (N_19132,N_10420,N_14303);
nand U19133 (N_19133,N_10632,N_10807);
nor U19134 (N_19134,N_11405,N_14131);
and U19135 (N_19135,N_12300,N_11306);
nand U19136 (N_19136,N_11160,N_12798);
xor U19137 (N_19137,N_14307,N_11099);
and U19138 (N_19138,N_10709,N_13359);
nand U19139 (N_19139,N_13831,N_14598);
or U19140 (N_19140,N_10088,N_13364);
xnor U19141 (N_19141,N_12392,N_14515);
nor U19142 (N_19142,N_10562,N_11787);
nand U19143 (N_19143,N_12387,N_10508);
xor U19144 (N_19144,N_11950,N_13928);
nand U19145 (N_19145,N_11939,N_12437);
and U19146 (N_19146,N_10035,N_12003);
nand U19147 (N_19147,N_10698,N_12502);
or U19148 (N_19148,N_13813,N_12683);
and U19149 (N_19149,N_12945,N_12321);
xor U19150 (N_19150,N_14188,N_10777);
nor U19151 (N_19151,N_12175,N_13626);
nor U19152 (N_19152,N_12126,N_14739);
and U19153 (N_19153,N_12496,N_14534);
or U19154 (N_19154,N_12608,N_14701);
or U19155 (N_19155,N_14165,N_13232);
nor U19156 (N_19156,N_11484,N_11003);
and U19157 (N_19157,N_14961,N_11508);
nor U19158 (N_19158,N_13964,N_10895);
or U19159 (N_19159,N_12399,N_12727);
nor U19160 (N_19160,N_13066,N_12479);
xnor U19161 (N_19161,N_12405,N_14192);
nor U19162 (N_19162,N_14735,N_14736);
and U19163 (N_19163,N_12069,N_12183);
and U19164 (N_19164,N_13785,N_13193);
or U19165 (N_19165,N_11647,N_12418);
nor U19166 (N_19166,N_11725,N_13692);
nand U19167 (N_19167,N_10175,N_14449);
nor U19168 (N_19168,N_10621,N_14290);
nand U19169 (N_19169,N_10688,N_12342);
nand U19170 (N_19170,N_14709,N_13183);
nand U19171 (N_19171,N_13446,N_13344);
or U19172 (N_19172,N_10685,N_13169);
xor U19173 (N_19173,N_14182,N_14728);
or U19174 (N_19174,N_13001,N_11485);
or U19175 (N_19175,N_14904,N_11144);
nor U19176 (N_19176,N_14202,N_13548);
and U19177 (N_19177,N_12344,N_11509);
and U19178 (N_19178,N_11097,N_13660);
and U19179 (N_19179,N_14842,N_12185);
or U19180 (N_19180,N_13684,N_14386);
nand U19181 (N_19181,N_11488,N_13781);
nor U19182 (N_19182,N_14144,N_11103);
and U19183 (N_19183,N_14378,N_13369);
or U19184 (N_19184,N_11884,N_12161);
nand U19185 (N_19185,N_11036,N_12420);
xnor U19186 (N_19186,N_13031,N_11014);
and U19187 (N_19187,N_11170,N_12199);
nand U19188 (N_19188,N_14653,N_14528);
or U19189 (N_19189,N_12568,N_14357);
xnor U19190 (N_19190,N_14794,N_14074);
or U19191 (N_19191,N_10453,N_11214);
or U19192 (N_19192,N_14477,N_11790);
nor U19193 (N_19193,N_10314,N_12541);
and U19194 (N_19194,N_14483,N_12403);
nand U19195 (N_19195,N_12514,N_11739);
or U19196 (N_19196,N_11370,N_12631);
nor U19197 (N_19197,N_14964,N_10324);
xor U19198 (N_19198,N_14150,N_14285);
and U19199 (N_19199,N_12652,N_10378);
nand U19200 (N_19200,N_10352,N_12699);
nand U19201 (N_19201,N_10980,N_10616);
xnor U19202 (N_19202,N_10905,N_10658);
or U19203 (N_19203,N_14191,N_10727);
or U19204 (N_19204,N_12354,N_14908);
xor U19205 (N_19205,N_11505,N_12255);
and U19206 (N_19206,N_13511,N_10633);
nand U19207 (N_19207,N_11241,N_12145);
nor U19208 (N_19208,N_11027,N_14453);
and U19209 (N_19209,N_10608,N_14067);
xnor U19210 (N_19210,N_14416,N_12834);
nand U19211 (N_19211,N_13620,N_12683);
or U19212 (N_19212,N_14858,N_13515);
nor U19213 (N_19213,N_10479,N_14194);
xor U19214 (N_19214,N_12346,N_13761);
xnor U19215 (N_19215,N_11148,N_12388);
and U19216 (N_19216,N_12044,N_13968);
and U19217 (N_19217,N_10610,N_14956);
nand U19218 (N_19218,N_14798,N_11996);
nor U19219 (N_19219,N_11914,N_10535);
xnor U19220 (N_19220,N_12323,N_13172);
or U19221 (N_19221,N_12031,N_10801);
nand U19222 (N_19222,N_11248,N_14810);
nor U19223 (N_19223,N_14570,N_12298);
nand U19224 (N_19224,N_12287,N_14490);
nand U19225 (N_19225,N_13920,N_11437);
and U19226 (N_19226,N_13333,N_12315);
nand U19227 (N_19227,N_11580,N_10100);
and U19228 (N_19228,N_12963,N_11055);
or U19229 (N_19229,N_11019,N_13100);
or U19230 (N_19230,N_11607,N_14232);
nand U19231 (N_19231,N_13234,N_12187);
or U19232 (N_19232,N_10212,N_11992);
xnor U19233 (N_19233,N_13499,N_13304);
xor U19234 (N_19234,N_11912,N_14644);
nand U19235 (N_19235,N_13660,N_11159);
and U19236 (N_19236,N_11559,N_12587);
and U19237 (N_19237,N_14461,N_10838);
nor U19238 (N_19238,N_10362,N_13170);
nand U19239 (N_19239,N_12073,N_11275);
and U19240 (N_19240,N_13125,N_13085);
nor U19241 (N_19241,N_13279,N_12615);
and U19242 (N_19242,N_14599,N_14644);
nand U19243 (N_19243,N_12856,N_11259);
nand U19244 (N_19244,N_12607,N_12031);
and U19245 (N_19245,N_11020,N_13908);
and U19246 (N_19246,N_14532,N_14799);
or U19247 (N_19247,N_13461,N_11513);
nand U19248 (N_19248,N_14364,N_12386);
nand U19249 (N_19249,N_13761,N_12665);
and U19250 (N_19250,N_14531,N_14490);
xnor U19251 (N_19251,N_10464,N_13215);
nor U19252 (N_19252,N_13619,N_11474);
nor U19253 (N_19253,N_10370,N_12882);
nor U19254 (N_19254,N_14523,N_10831);
nand U19255 (N_19255,N_14188,N_14227);
or U19256 (N_19256,N_12080,N_12897);
and U19257 (N_19257,N_13673,N_14474);
nand U19258 (N_19258,N_12630,N_12318);
nand U19259 (N_19259,N_12668,N_13159);
nand U19260 (N_19260,N_13307,N_11078);
and U19261 (N_19261,N_14096,N_12273);
xor U19262 (N_19262,N_10550,N_13646);
nor U19263 (N_19263,N_11226,N_11978);
or U19264 (N_19264,N_11185,N_11785);
xnor U19265 (N_19265,N_12787,N_13591);
xor U19266 (N_19266,N_14703,N_13264);
and U19267 (N_19267,N_14871,N_14163);
nand U19268 (N_19268,N_13768,N_10926);
or U19269 (N_19269,N_10592,N_10748);
or U19270 (N_19270,N_11226,N_13814);
and U19271 (N_19271,N_12951,N_14283);
xnor U19272 (N_19272,N_10804,N_13050);
nor U19273 (N_19273,N_13829,N_11853);
nor U19274 (N_19274,N_11756,N_12310);
and U19275 (N_19275,N_10734,N_10323);
and U19276 (N_19276,N_10639,N_13477);
nor U19277 (N_19277,N_11152,N_11466);
nand U19278 (N_19278,N_14201,N_11938);
nor U19279 (N_19279,N_11741,N_11558);
nor U19280 (N_19280,N_11667,N_10758);
xnor U19281 (N_19281,N_11890,N_14499);
or U19282 (N_19282,N_11229,N_14959);
and U19283 (N_19283,N_10572,N_13777);
nor U19284 (N_19284,N_14095,N_13975);
or U19285 (N_19285,N_13712,N_13976);
and U19286 (N_19286,N_11701,N_13594);
nor U19287 (N_19287,N_13549,N_13370);
and U19288 (N_19288,N_13879,N_11167);
xor U19289 (N_19289,N_12600,N_10830);
nor U19290 (N_19290,N_11001,N_13747);
and U19291 (N_19291,N_11658,N_12355);
xor U19292 (N_19292,N_14608,N_13193);
nand U19293 (N_19293,N_11341,N_13736);
nand U19294 (N_19294,N_13351,N_12017);
and U19295 (N_19295,N_14752,N_10096);
nand U19296 (N_19296,N_10388,N_11100);
xnor U19297 (N_19297,N_13241,N_14935);
nand U19298 (N_19298,N_11286,N_11845);
and U19299 (N_19299,N_13132,N_12440);
or U19300 (N_19300,N_14776,N_11839);
nand U19301 (N_19301,N_12703,N_10314);
nand U19302 (N_19302,N_12130,N_10144);
nor U19303 (N_19303,N_13923,N_12331);
or U19304 (N_19304,N_14041,N_14476);
nand U19305 (N_19305,N_12685,N_11900);
nand U19306 (N_19306,N_11034,N_12142);
nand U19307 (N_19307,N_10406,N_11076);
nand U19308 (N_19308,N_11995,N_10138);
nor U19309 (N_19309,N_14516,N_14375);
or U19310 (N_19310,N_13129,N_10071);
xnor U19311 (N_19311,N_14966,N_12678);
nor U19312 (N_19312,N_12875,N_14849);
xor U19313 (N_19313,N_14427,N_10768);
and U19314 (N_19314,N_10592,N_10785);
nor U19315 (N_19315,N_10746,N_13698);
nand U19316 (N_19316,N_11458,N_11967);
or U19317 (N_19317,N_11321,N_12858);
nor U19318 (N_19318,N_10123,N_14094);
nor U19319 (N_19319,N_12822,N_12341);
nand U19320 (N_19320,N_14261,N_10066);
xor U19321 (N_19321,N_10711,N_14583);
xor U19322 (N_19322,N_10781,N_12819);
nor U19323 (N_19323,N_10732,N_10752);
or U19324 (N_19324,N_11485,N_11504);
and U19325 (N_19325,N_14683,N_13711);
nand U19326 (N_19326,N_13273,N_13798);
nand U19327 (N_19327,N_10743,N_13100);
nor U19328 (N_19328,N_13518,N_12860);
nor U19329 (N_19329,N_12846,N_12259);
nand U19330 (N_19330,N_12199,N_11747);
xor U19331 (N_19331,N_13153,N_11437);
and U19332 (N_19332,N_13020,N_12043);
or U19333 (N_19333,N_14854,N_14117);
or U19334 (N_19334,N_11273,N_11462);
or U19335 (N_19335,N_12981,N_12485);
or U19336 (N_19336,N_12199,N_13274);
and U19337 (N_19337,N_14159,N_11399);
and U19338 (N_19338,N_10717,N_14015);
nor U19339 (N_19339,N_11045,N_10411);
xor U19340 (N_19340,N_11123,N_10735);
nor U19341 (N_19341,N_12375,N_13219);
and U19342 (N_19342,N_11555,N_14186);
and U19343 (N_19343,N_14301,N_13311);
nand U19344 (N_19344,N_10392,N_12768);
xor U19345 (N_19345,N_14235,N_14283);
nand U19346 (N_19346,N_12695,N_14425);
or U19347 (N_19347,N_11617,N_10334);
nand U19348 (N_19348,N_10021,N_10751);
or U19349 (N_19349,N_14596,N_10043);
nand U19350 (N_19350,N_13815,N_13916);
and U19351 (N_19351,N_10071,N_11197);
and U19352 (N_19352,N_12355,N_10888);
xnor U19353 (N_19353,N_14926,N_11690);
nand U19354 (N_19354,N_14247,N_12595);
or U19355 (N_19355,N_10656,N_12709);
nand U19356 (N_19356,N_11184,N_13124);
or U19357 (N_19357,N_12726,N_11534);
nor U19358 (N_19358,N_11835,N_13194);
nor U19359 (N_19359,N_10426,N_12664);
nand U19360 (N_19360,N_13275,N_13537);
and U19361 (N_19361,N_13705,N_10957);
and U19362 (N_19362,N_10961,N_14991);
xor U19363 (N_19363,N_14605,N_13964);
or U19364 (N_19364,N_11500,N_13394);
nand U19365 (N_19365,N_12629,N_13413);
and U19366 (N_19366,N_13457,N_14863);
or U19367 (N_19367,N_11992,N_14155);
or U19368 (N_19368,N_12893,N_13486);
or U19369 (N_19369,N_11710,N_10992);
or U19370 (N_19370,N_11918,N_10217);
nor U19371 (N_19371,N_11322,N_14089);
and U19372 (N_19372,N_12155,N_12829);
nand U19373 (N_19373,N_10911,N_12672);
xor U19374 (N_19374,N_14188,N_12863);
nor U19375 (N_19375,N_13517,N_12646);
nand U19376 (N_19376,N_11526,N_11823);
and U19377 (N_19377,N_13765,N_10587);
or U19378 (N_19378,N_12137,N_11433);
nand U19379 (N_19379,N_12593,N_13207);
and U19380 (N_19380,N_12563,N_10760);
nor U19381 (N_19381,N_13788,N_11465);
nor U19382 (N_19382,N_14985,N_13457);
and U19383 (N_19383,N_11354,N_13203);
and U19384 (N_19384,N_14613,N_11820);
and U19385 (N_19385,N_14522,N_13632);
and U19386 (N_19386,N_14641,N_13983);
nor U19387 (N_19387,N_13223,N_14548);
nand U19388 (N_19388,N_11350,N_14557);
nand U19389 (N_19389,N_13204,N_11956);
nand U19390 (N_19390,N_13112,N_14311);
or U19391 (N_19391,N_11627,N_12545);
and U19392 (N_19392,N_12975,N_11008);
and U19393 (N_19393,N_14136,N_11998);
nand U19394 (N_19394,N_14040,N_13769);
nand U19395 (N_19395,N_13006,N_13641);
and U19396 (N_19396,N_10151,N_14859);
nand U19397 (N_19397,N_11558,N_10086);
or U19398 (N_19398,N_12871,N_13678);
nand U19399 (N_19399,N_12058,N_10852);
xor U19400 (N_19400,N_12295,N_11583);
and U19401 (N_19401,N_13434,N_10956);
nand U19402 (N_19402,N_12628,N_14228);
nor U19403 (N_19403,N_13996,N_10436);
nor U19404 (N_19404,N_11739,N_13661);
and U19405 (N_19405,N_11649,N_12634);
nor U19406 (N_19406,N_13786,N_13220);
and U19407 (N_19407,N_12731,N_14566);
and U19408 (N_19408,N_10303,N_14350);
xor U19409 (N_19409,N_12747,N_12895);
or U19410 (N_19410,N_10479,N_14223);
or U19411 (N_19411,N_12501,N_10181);
nor U19412 (N_19412,N_12968,N_12500);
nor U19413 (N_19413,N_10223,N_10663);
and U19414 (N_19414,N_13675,N_12539);
xnor U19415 (N_19415,N_11880,N_13353);
nor U19416 (N_19416,N_12760,N_13263);
and U19417 (N_19417,N_11040,N_12707);
or U19418 (N_19418,N_10070,N_14966);
xnor U19419 (N_19419,N_10452,N_13817);
or U19420 (N_19420,N_12670,N_11779);
or U19421 (N_19421,N_14662,N_13499);
nand U19422 (N_19422,N_11550,N_12144);
or U19423 (N_19423,N_14563,N_10519);
nor U19424 (N_19424,N_10310,N_14842);
nor U19425 (N_19425,N_14599,N_10712);
xnor U19426 (N_19426,N_14118,N_13795);
nor U19427 (N_19427,N_12758,N_12087);
nor U19428 (N_19428,N_14000,N_13006);
xor U19429 (N_19429,N_11528,N_12695);
nor U19430 (N_19430,N_14509,N_11543);
nor U19431 (N_19431,N_10401,N_13390);
and U19432 (N_19432,N_10096,N_10508);
and U19433 (N_19433,N_10395,N_10122);
or U19434 (N_19434,N_12943,N_14200);
and U19435 (N_19435,N_10104,N_14976);
and U19436 (N_19436,N_14759,N_14727);
nor U19437 (N_19437,N_12038,N_13494);
and U19438 (N_19438,N_12045,N_13071);
or U19439 (N_19439,N_13338,N_12628);
xnor U19440 (N_19440,N_13503,N_14254);
nor U19441 (N_19441,N_14967,N_12156);
xor U19442 (N_19442,N_13832,N_12441);
nor U19443 (N_19443,N_14978,N_11003);
nand U19444 (N_19444,N_10076,N_13036);
and U19445 (N_19445,N_13305,N_10486);
nand U19446 (N_19446,N_13973,N_14740);
xnor U19447 (N_19447,N_12939,N_12385);
or U19448 (N_19448,N_11318,N_10966);
nor U19449 (N_19449,N_12814,N_10846);
or U19450 (N_19450,N_13411,N_13103);
nor U19451 (N_19451,N_10305,N_12956);
or U19452 (N_19452,N_10484,N_13281);
xnor U19453 (N_19453,N_11984,N_13406);
or U19454 (N_19454,N_10120,N_14309);
and U19455 (N_19455,N_13725,N_10000);
nand U19456 (N_19456,N_10404,N_14012);
xnor U19457 (N_19457,N_10458,N_10109);
nand U19458 (N_19458,N_10894,N_13958);
and U19459 (N_19459,N_14757,N_14059);
xor U19460 (N_19460,N_13782,N_10638);
xor U19461 (N_19461,N_14072,N_14112);
xnor U19462 (N_19462,N_14294,N_10723);
xor U19463 (N_19463,N_12850,N_11542);
xnor U19464 (N_19464,N_13808,N_13370);
or U19465 (N_19465,N_14042,N_11735);
nand U19466 (N_19466,N_10750,N_10873);
xor U19467 (N_19467,N_14523,N_14104);
nand U19468 (N_19468,N_13982,N_12365);
xnor U19469 (N_19469,N_13051,N_13265);
or U19470 (N_19470,N_10688,N_14878);
nor U19471 (N_19471,N_11461,N_10604);
nor U19472 (N_19472,N_10016,N_12716);
and U19473 (N_19473,N_10784,N_12372);
nand U19474 (N_19474,N_13723,N_11003);
nor U19475 (N_19475,N_10751,N_11659);
or U19476 (N_19476,N_11349,N_11037);
or U19477 (N_19477,N_13787,N_14724);
or U19478 (N_19478,N_13845,N_11215);
nand U19479 (N_19479,N_12990,N_14589);
nor U19480 (N_19480,N_10589,N_12548);
nand U19481 (N_19481,N_11981,N_13132);
nand U19482 (N_19482,N_11600,N_13438);
nand U19483 (N_19483,N_13872,N_13602);
nor U19484 (N_19484,N_13314,N_12495);
nor U19485 (N_19485,N_11320,N_12006);
xnor U19486 (N_19486,N_14724,N_10105);
nor U19487 (N_19487,N_13261,N_11163);
nor U19488 (N_19488,N_11133,N_11541);
nand U19489 (N_19489,N_10919,N_13622);
nor U19490 (N_19490,N_14229,N_12258);
or U19491 (N_19491,N_14103,N_13750);
nor U19492 (N_19492,N_13516,N_14829);
xnor U19493 (N_19493,N_11854,N_14053);
nor U19494 (N_19494,N_13939,N_12227);
nor U19495 (N_19495,N_12406,N_10133);
and U19496 (N_19496,N_12529,N_14209);
or U19497 (N_19497,N_13173,N_14822);
or U19498 (N_19498,N_14031,N_11418);
or U19499 (N_19499,N_14292,N_13077);
nand U19500 (N_19500,N_14183,N_13269);
nor U19501 (N_19501,N_11142,N_11014);
xnor U19502 (N_19502,N_11754,N_11231);
nor U19503 (N_19503,N_12117,N_10394);
nor U19504 (N_19504,N_14675,N_11640);
xnor U19505 (N_19505,N_13702,N_11772);
and U19506 (N_19506,N_12408,N_14299);
nor U19507 (N_19507,N_12206,N_11797);
nor U19508 (N_19508,N_13442,N_12247);
xor U19509 (N_19509,N_10817,N_12920);
xor U19510 (N_19510,N_13566,N_13334);
nor U19511 (N_19511,N_11264,N_13993);
nor U19512 (N_19512,N_13535,N_12539);
xnor U19513 (N_19513,N_10672,N_10535);
xnor U19514 (N_19514,N_13532,N_14092);
and U19515 (N_19515,N_10398,N_13901);
and U19516 (N_19516,N_14815,N_11274);
nor U19517 (N_19517,N_11067,N_10467);
xor U19518 (N_19518,N_14415,N_12779);
and U19519 (N_19519,N_13036,N_11686);
nand U19520 (N_19520,N_14464,N_14001);
nand U19521 (N_19521,N_14002,N_14032);
or U19522 (N_19522,N_13193,N_12004);
and U19523 (N_19523,N_14044,N_13031);
nor U19524 (N_19524,N_11358,N_12720);
nor U19525 (N_19525,N_10082,N_11569);
nand U19526 (N_19526,N_13915,N_12426);
and U19527 (N_19527,N_11055,N_14025);
nand U19528 (N_19528,N_11272,N_14410);
nand U19529 (N_19529,N_14718,N_11153);
xor U19530 (N_19530,N_14327,N_10242);
nand U19531 (N_19531,N_14548,N_14995);
nor U19532 (N_19532,N_12186,N_10466);
and U19533 (N_19533,N_14770,N_14976);
nor U19534 (N_19534,N_13914,N_13982);
nand U19535 (N_19535,N_11114,N_10326);
and U19536 (N_19536,N_10134,N_13374);
or U19537 (N_19537,N_14608,N_14763);
xor U19538 (N_19538,N_10665,N_10142);
and U19539 (N_19539,N_11388,N_12844);
xnor U19540 (N_19540,N_14535,N_10343);
and U19541 (N_19541,N_13393,N_10139);
nor U19542 (N_19542,N_13106,N_12738);
nor U19543 (N_19543,N_12935,N_10194);
nand U19544 (N_19544,N_11028,N_14999);
nor U19545 (N_19545,N_13822,N_14747);
nand U19546 (N_19546,N_13563,N_12529);
nor U19547 (N_19547,N_12776,N_13958);
or U19548 (N_19548,N_10074,N_11394);
and U19549 (N_19549,N_12652,N_13222);
nor U19550 (N_19550,N_13554,N_11141);
xnor U19551 (N_19551,N_11476,N_10321);
nand U19552 (N_19552,N_12417,N_12992);
xor U19553 (N_19553,N_12209,N_13703);
xor U19554 (N_19554,N_10376,N_10833);
xnor U19555 (N_19555,N_14218,N_13310);
nor U19556 (N_19556,N_13555,N_14792);
nor U19557 (N_19557,N_14984,N_10988);
nor U19558 (N_19558,N_13027,N_10523);
nor U19559 (N_19559,N_10611,N_14648);
nor U19560 (N_19560,N_13629,N_12194);
xor U19561 (N_19561,N_12500,N_13839);
nor U19562 (N_19562,N_12460,N_11506);
nor U19563 (N_19563,N_14799,N_12615);
or U19564 (N_19564,N_11364,N_10798);
nor U19565 (N_19565,N_12449,N_14522);
and U19566 (N_19566,N_13639,N_14405);
or U19567 (N_19567,N_11376,N_13623);
xnor U19568 (N_19568,N_13589,N_11290);
and U19569 (N_19569,N_10356,N_12281);
and U19570 (N_19570,N_11315,N_13331);
or U19571 (N_19571,N_13004,N_11522);
and U19572 (N_19572,N_10972,N_11952);
or U19573 (N_19573,N_13444,N_12518);
nor U19574 (N_19574,N_10450,N_10482);
and U19575 (N_19575,N_12660,N_14849);
or U19576 (N_19576,N_13650,N_14740);
or U19577 (N_19577,N_14573,N_10542);
and U19578 (N_19578,N_14623,N_10048);
nand U19579 (N_19579,N_11523,N_10913);
nand U19580 (N_19580,N_12422,N_14696);
nor U19581 (N_19581,N_10491,N_13770);
and U19582 (N_19582,N_12632,N_14822);
xnor U19583 (N_19583,N_14206,N_10519);
or U19584 (N_19584,N_10043,N_12539);
nand U19585 (N_19585,N_14524,N_10262);
xnor U19586 (N_19586,N_14985,N_11231);
xor U19587 (N_19587,N_10774,N_13208);
nor U19588 (N_19588,N_14178,N_12066);
or U19589 (N_19589,N_14159,N_12018);
or U19590 (N_19590,N_12062,N_11396);
xnor U19591 (N_19591,N_14987,N_10742);
or U19592 (N_19592,N_11104,N_10339);
or U19593 (N_19593,N_11512,N_11457);
nand U19594 (N_19594,N_12586,N_12443);
nor U19595 (N_19595,N_13834,N_13297);
xor U19596 (N_19596,N_11571,N_10180);
nor U19597 (N_19597,N_13324,N_12278);
xnor U19598 (N_19598,N_13976,N_10444);
nand U19599 (N_19599,N_13235,N_10417);
or U19600 (N_19600,N_11468,N_10338);
or U19601 (N_19601,N_12029,N_11867);
nor U19602 (N_19602,N_13526,N_12600);
and U19603 (N_19603,N_11052,N_14603);
nor U19604 (N_19604,N_11882,N_13123);
nor U19605 (N_19605,N_13788,N_14767);
and U19606 (N_19606,N_14796,N_10708);
nand U19607 (N_19607,N_11881,N_14121);
and U19608 (N_19608,N_12546,N_12531);
nor U19609 (N_19609,N_14675,N_14140);
nor U19610 (N_19610,N_12651,N_11065);
xor U19611 (N_19611,N_10833,N_12062);
nand U19612 (N_19612,N_11743,N_10125);
xnor U19613 (N_19613,N_11443,N_12635);
and U19614 (N_19614,N_11185,N_13648);
or U19615 (N_19615,N_13432,N_14732);
xnor U19616 (N_19616,N_12728,N_14085);
xor U19617 (N_19617,N_11031,N_13945);
or U19618 (N_19618,N_11535,N_10299);
or U19619 (N_19619,N_10839,N_13166);
or U19620 (N_19620,N_10291,N_11060);
nand U19621 (N_19621,N_11449,N_13690);
nand U19622 (N_19622,N_12979,N_14922);
and U19623 (N_19623,N_13894,N_10040);
or U19624 (N_19624,N_10707,N_11566);
nand U19625 (N_19625,N_11758,N_14448);
xnor U19626 (N_19626,N_12340,N_14456);
and U19627 (N_19627,N_11992,N_12717);
or U19628 (N_19628,N_14590,N_14601);
and U19629 (N_19629,N_11810,N_11432);
nor U19630 (N_19630,N_13450,N_12782);
xor U19631 (N_19631,N_11560,N_12294);
nor U19632 (N_19632,N_12518,N_10690);
nand U19633 (N_19633,N_13570,N_10130);
nand U19634 (N_19634,N_10221,N_11998);
nand U19635 (N_19635,N_10569,N_12348);
xnor U19636 (N_19636,N_14114,N_13911);
or U19637 (N_19637,N_10743,N_12219);
nand U19638 (N_19638,N_12478,N_14077);
nand U19639 (N_19639,N_11442,N_13453);
nand U19640 (N_19640,N_10962,N_13513);
and U19641 (N_19641,N_10775,N_10643);
xor U19642 (N_19642,N_14613,N_12615);
and U19643 (N_19643,N_11649,N_11529);
or U19644 (N_19644,N_12278,N_12125);
nor U19645 (N_19645,N_12135,N_11304);
and U19646 (N_19646,N_10447,N_12709);
nand U19647 (N_19647,N_14875,N_13152);
nand U19648 (N_19648,N_12281,N_13558);
nor U19649 (N_19649,N_11487,N_13938);
or U19650 (N_19650,N_14445,N_13806);
xnor U19651 (N_19651,N_14209,N_14686);
nor U19652 (N_19652,N_10893,N_14051);
xor U19653 (N_19653,N_10550,N_13572);
or U19654 (N_19654,N_14632,N_11202);
or U19655 (N_19655,N_12060,N_10754);
and U19656 (N_19656,N_12706,N_12623);
or U19657 (N_19657,N_12513,N_11350);
nor U19658 (N_19658,N_10326,N_13195);
and U19659 (N_19659,N_14146,N_12190);
nor U19660 (N_19660,N_11477,N_14172);
nand U19661 (N_19661,N_11726,N_10859);
nor U19662 (N_19662,N_12120,N_11323);
and U19663 (N_19663,N_13077,N_10600);
xor U19664 (N_19664,N_10960,N_12973);
or U19665 (N_19665,N_11208,N_11945);
nand U19666 (N_19666,N_12457,N_10199);
and U19667 (N_19667,N_12881,N_14947);
xor U19668 (N_19668,N_14958,N_10350);
or U19669 (N_19669,N_12032,N_11341);
or U19670 (N_19670,N_13175,N_13833);
and U19671 (N_19671,N_12306,N_11011);
xnor U19672 (N_19672,N_10670,N_12067);
and U19673 (N_19673,N_13210,N_13185);
and U19674 (N_19674,N_10276,N_13074);
xor U19675 (N_19675,N_11482,N_10371);
or U19676 (N_19676,N_14170,N_14919);
and U19677 (N_19677,N_10281,N_11506);
and U19678 (N_19678,N_13467,N_12505);
nand U19679 (N_19679,N_10100,N_10859);
or U19680 (N_19680,N_12334,N_14825);
or U19681 (N_19681,N_10292,N_11540);
or U19682 (N_19682,N_13346,N_11138);
nand U19683 (N_19683,N_13199,N_13943);
or U19684 (N_19684,N_12884,N_12863);
nor U19685 (N_19685,N_10849,N_13559);
or U19686 (N_19686,N_13335,N_13686);
xor U19687 (N_19687,N_12357,N_14704);
nor U19688 (N_19688,N_13602,N_12943);
or U19689 (N_19689,N_13946,N_10742);
nor U19690 (N_19690,N_13565,N_10254);
nand U19691 (N_19691,N_13818,N_13228);
and U19692 (N_19692,N_14197,N_12399);
xor U19693 (N_19693,N_11865,N_10369);
xor U19694 (N_19694,N_10340,N_11950);
nand U19695 (N_19695,N_14096,N_14488);
nand U19696 (N_19696,N_12059,N_11429);
and U19697 (N_19697,N_14590,N_11689);
xnor U19698 (N_19698,N_12951,N_13515);
xor U19699 (N_19699,N_12491,N_10653);
and U19700 (N_19700,N_12070,N_11422);
xor U19701 (N_19701,N_13289,N_13481);
xor U19702 (N_19702,N_11100,N_10421);
and U19703 (N_19703,N_10305,N_13329);
xnor U19704 (N_19704,N_14231,N_10036);
xor U19705 (N_19705,N_14691,N_14346);
xnor U19706 (N_19706,N_14406,N_10298);
xor U19707 (N_19707,N_14200,N_12895);
nand U19708 (N_19708,N_11174,N_12161);
nand U19709 (N_19709,N_10719,N_14732);
nand U19710 (N_19710,N_10548,N_14530);
or U19711 (N_19711,N_12870,N_13408);
and U19712 (N_19712,N_10752,N_14154);
and U19713 (N_19713,N_10613,N_10773);
nor U19714 (N_19714,N_10303,N_12398);
nand U19715 (N_19715,N_12283,N_13266);
nand U19716 (N_19716,N_10566,N_14079);
xor U19717 (N_19717,N_12797,N_12966);
xor U19718 (N_19718,N_13424,N_11861);
or U19719 (N_19719,N_12665,N_12783);
xnor U19720 (N_19720,N_14643,N_12023);
and U19721 (N_19721,N_10635,N_13038);
nand U19722 (N_19722,N_11026,N_10473);
or U19723 (N_19723,N_13964,N_13087);
xnor U19724 (N_19724,N_10356,N_10542);
and U19725 (N_19725,N_13941,N_13755);
or U19726 (N_19726,N_14595,N_12169);
and U19727 (N_19727,N_14947,N_10467);
xor U19728 (N_19728,N_14931,N_10591);
xor U19729 (N_19729,N_14959,N_11183);
nor U19730 (N_19730,N_10991,N_10484);
xnor U19731 (N_19731,N_13794,N_11412);
or U19732 (N_19732,N_14212,N_13055);
xor U19733 (N_19733,N_11192,N_10145);
nand U19734 (N_19734,N_11492,N_13903);
or U19735 (N_19735,N_14729,N_13246);
nor U19736 (N_19736,N_14616,N_13241);
nand U19737 (N_19737,N_11109,N_14408);
nor U19738 (N_19738,N_12163,N_11261);
xor U19739 (N_19739,N_12759,N_14081);
or U19740 (N_19740,N_14304,N_11582);
nor U19741 (N_19741,N_14029,N_11127);
nor U19742 (N_19742,N_14308,N_11336);
or U19743 (N_19743,N_12963,N_13343);
and U19744 (N_19744,N_12310,N_14379);
xor U19745 (N_19745,N_11462,N_11911);
or U19746 (N_19746,N_13948,N_12639);
xor U19747 (N_19747,N_12989,N_12801);
xor U19748 (N_19748,N_11172,N_12399);
or U19749 (N_19749,N_10269,N_11151);
nor U19750 (N_19750,N_14531,N_11621);
nor U19751 (N_19751,N_12735,N_14719);
nand U19752 (N_19752,N_13597,N_12946);
or U19753 (N_19753,N_13203,N_13265);
nand U19754 (N_19754,N_11056,N_14068);
xor U19755 (N_19755,N_14463,N_13700);
and U19756 (N_19756,N_10044,N_14102);
nand U19757 (N_19757,N_13536,N_10290);
nand U19758 (N_19758,N_12842,N_11547);
xnor U19759 (N_19759,N_11017,N_10612);
and U19760 (N_19760,N_12328,N_13570);
xnor U19761 (N_19761,N_12727,N_12808);
xnor U19762 (N_19762,N_11279,N_11152);
or U19763 (N_19763,N_11164,N_12130);
nand U19764 (N_19764,N_10839,N_14118);
nor U19765 (N_19765,N_11522,N_10947);
nand U19766 (N_19766,N_10851,N_12144);
and U19767 (N_19767,N_14935,N_11397);
nor U19768 (N_19768,N_13813,N_11848);
xnor U19769 (N_19769,N_10156,N_14985);
nor U19770 (N_19770,N_11772,N_10308);
nand U19771 (N_19771,N_12118,N_13768);
nor U19772 (N_19772,N_14118,N_14923);
nor U19773 (N_19773,N_11537,N_12801);
and U19774 (N_19774,N_11920,N_13175);
and U19775 (N_19775,N_10153,N_14065);
nand U19776 (N_19776,N_14346,N_11234);
nand U19777 (N_19777,N_10192,N_12934);
nor U19778 (N_19778,N_14030,N_12917);
nor U19779 (N_19779,N_10712,N_13138);
and U19780 (N_19780,N_12049,N_13189);
xnor U19781 (N_19781,N_13292,N_13834);
and U19782 (N_19782,N_13511,N_10026);
or U19783 (N_19783,N_10524,N_12311);
nor U19784 (N_19784,N_10964,N_14310);
xor U19785 (N_19785,N_10419,N_10151);
nor U19786 (N_19786,N_11701,N_13459);
and U19787 (N_19787,N_12344,N_13282);
or U19788 (N_19788,N_11750,N_10920);
nand U19789 (N_19789,N_12480,N_12401);
nor U19790 (N_19790,N_13124,N_14467);
xnor U19791 (N_19791,N_11443,N_14812);
nand U19792 (N_19792,N_12911,N_12901);
nand U19793 (N_19793,N_10707,N_11239);
xor U19794 (N_19794,N_10933,N_11791);
and U19795 (N_19795,N_11970,N_12418);
or U19796 (N_19796,N_10315,N_13441);
and U19797 (N_19797,N_11779,N_14453);
nand U19798 (N_19798,N_13224,N_14577);
xnor U19799 (N_19799,N_14992,N_14468);
or U19800 (N_19800,N_10634,N_12550);
nor U19801 (N_19801,N_14965,N_14014);
nor U19802 (N_19802,N_14699,N_10791);
nand U19803 (N_19803,N_10656,N_13053);
nor U19804 (N_19804,N_12416,N_10721);
or U19805 (N_19805,N_10167,N_14384);
and U19806 (N_19806,N_13428,N_14185);
and U19807 (N_19807,N_10762,N_10296);
nor U19808 (N_19808,N_11075,N_13574);
nor U19809 (N_19809,N_14680,N_13986);
and U19810 (N_19810,N_14984,N_10111);
or U19811 (N_19811,N_10223,N_13216);
and U19812 (N_19812,N_11638,N_10646);
nand U19813 (N_19813,N_14928,N_13153);
nor U19814 (N_19814,N_13796,N_14901);
and U19815 (N_19815,N_12713,N_10644);
and U19816 (N_19816,N_12829,N_11874);
nor U19817 (N_19817,N_11265,N_14947);
nand U19818 (N_19818,N_12559,N_10102);
nor U19819 (N_19819,N_12388,N_11914);
xor U19820 (N_19820,N_13117,N_10659);
and U19821 (N_19821,N_11901,N_10580);
and U19822 (N_19822,N_10384,N_13704);
xor U19823 (N_19823,N_14552,N_14829);
xor U19824 (N_19824,N_10458,N_13724);
xor U19825 (N_19825,N_14028,N_10273);
or U19826 (N_19826,N_11943,N_10107);
and U19827 (N_19827,N_13549,N_10972);
nand U19828 (N_19828,N_14305,N_11373);
xnor U19829 (N_19829,N_12107,N_11493);
nor U19830 (N_19830,N_13098,N_10710);
or U19831 (N_19831,N_14529,N_10436);
nor U19832 (N_19832,N_10564,N_11978);
or U19833 (N_19833,N_14159,N_14809);
and U19834 (N_19834,N_11120,N_11043);
or U19835 (N_19835,N_14814,N_11620);
xor U19836 (N_19836,N_12845,N_14213);
and U19837 (N_19837,N_10301,N_13690);
and U19838 (N_19838,N_13772,N_10032);
xor U19839 (N_19839,N_12748,N_14491);
and U19840 (N_19840,N_11981,N_13090);
xnor U19841 (N_19841,N_11679,N_14734);
and U19842 (N_19842,N_12703,N_12132);
xor U19843 (N_19843,N_13086,N_12065);
nor U19844 (N_19844,N_12315,N_12788);
nor U19845 (N_19845,N_10203,N_11757);
or U19846 (N_19846,N_12616,N_10127);
or U19847 (N_19847,N_14320,N_10921);
nand U19848 (N_19848,N_10282,N_11460);
nor U19849 (N_19849,N_10389,N_10576);
and U19850 (N_19850,N_13728,N_14781);
and U19851 (N_19851,N_13118,N_10386);
xor U19852 (N_19852,N_14508,N_10192);
nor U19853 (N_19853,N_14025,N_13474);
nor U19854 (N_19854,N_10488,N_10371);
or U19855 (N_19855,N_14311,N_11213);
and U19856 (N_19856,N_12723,N_12821);
nor U19857 (N_19857,N_11578,N_14905);
nor U19858 (N_19858,N_13310,N_10498);
or U19859 (N_19859,N_14231,N_11186);
nor U19860 (N_19860,N_12501,N_12816);
or U19861 (N_19861,N_13596,N_13790);
and U19862 (N_19862,N_13628,N_13852);
nor U19863 (N_19863,N_11120,N_10570);
and U19864 (N_19864,N_11971,N_13239);
nor U19865 (N_19865,N_11440,N_14841);
and U19866 (N_19866,N_12733,N_14711);
nor U19867 (N_19867,N_13653,N_11071);
and U19868 (N_19868,N_13684,N_10402);
nand U19869 (N_19869,N_12516,N_14207);
or U19870 (N_19870,N_13424,N_10290);
or U19871 (N_19871,N_12587,N_14060);
xnor U19872 (N_19872,N_13852,N_11706);
xnor U19873 (N_19873,N_11242,N_11580);
nand U19874 (N_19874,N_13647,N_14684);
nor U19875 (N_19875,N_12707,N_12785);
and U19876 (N_19876,N_13484,N_12900);
and U19877 (N_19877,N_12654,N_14525);
and U19878 (N_19878,N_11725,N_11589);
or U19879 (N_19879,N_12812,N_14189);
and U19880 (N_19880,N_12163,N_14737);
and U19881 (N_19881,N_11486,N_13760);
xnor U19882 (N_19882,N_12496,N_11664);
nor U19883 (N_19883,N_12604,N_14181);
nor U19884 (N_19884,N_12893,N_11168);
nor U19885 (N_19885,N_13241,N_10475);
and U19886 (N_19886,N_12549,N_13316);
and U19887 (N_19887,N_14141,N_12760);
or U19888 (N_19888,N_12775,N_14896);
xnor U19889 (N_19889,N_13021,N_12353);
and U19890 (N_19890,N_13460,N_10725);
and U19891 (N_19891,N_14978,N_10620);
xnor U19892 (N_19892,N_13035,N_10794);
or U19893 (N_19893,N_13285,N_10963);
or U19894 (N_19894,N_14074,N_11727);
nand U19895 (N_19895,N_12614,N_12029);
nor U19896 (N_19896,N_12611,N_14107);
nor U19897 (N_19897,N_13748,N_11661);
or U19898 (N_19898,N_14774,N_12992);
nor U19899 (N_19899,N_14904,N_14093);
nand U19900 (N_19900,N_10213,N_12769);
and U19901 (N_19901,N_13947,N_13209);
and U19902 (N_19902,N_13967,N_14037);
or U19903 (N_19903,N_14440,N_11593);
nor U19904 (N_19904,N_11017,N_13819);
or U19905 (N_19905,N_13538,N_12188);
xnor U19906 (N_19906,N_13599,N_14101);
and U19907 (N_19907,N_14597,N_14586);
nand U19908 (N_19908,N_12014,N_11970);
and U19909 (N_19909,N_14357,N_13569);
nor U19910 (N_19910,N_14134,N_14030);
nor U19911 (N_19911,N_13779,N_12902);
and U19912 (N_19912,N_10951,N_11956);
and U19913 (N_19913,N_12389,N_11799);
nor U19914 (N_19914,N_13571,N_10560);
and U19915 (N_19915,N_10998,N_14330);
or U19916 (N_19916,N_14903,N_13514);
and U19917 (N_19917,N_14243,N_14792);
nand U19918 (N_19918,N_11034,N_10215);
or U19919 (N_19919,N_12535,N_10828);
or U19920 (N_19920,N_11929,N_11518);
xor U19921 (N_19921,N_13641,N_12112);
or U19922 (N_19922,N_10101,N_10406);
and U19923 (N_19923,N_12063,N_14112);
nand U19924 (N_19924,N_12211,N_12883);
xor U19925 (N_19925,N_13552,N_13345);
nand U19926 (N_19926,N_13167,N_12994);
nand U19927 (N_19927,N_12839,N_11820);
nand U19928 (N_19928,N_14521,N_11797);
xor U19929 (N_19929,N_10692,N_13403);
xnor U19930 (N_19930,N_14320,N_10402);
nor U19931 (N_19931,N_11031,N_12077);
or U19932 (N_19932,N_12950,N_10906);
or U19933 (N_19933,N_13177,N_14034);
nor U19934 (N_19934,N_10323,N_10328);
or U19935 (N_19935,N_11253,N_10791);
nand U19936 (N_19936,N_13667,N_14671);
nand U19937 (N_19937,N_13585,N_10902);
nand U19938 (N_19938,N_12483,N_12782);
and U19939 (N_19939,N_11035,N_11041);
nand U19940 (N_19940,N_12748,N_12001);
or U19941 (N_19941,N_14327,N_12448);
and U19942 (N_19942,N_13415,N_11223);
or U19943 (N_19943,N_14017,N_11883);
nand U19944 (N_19944,N_14452,N_13763);
nand U19945 (N_19945,N_14041,N_12379);
or U19946 (N_19946,N_13785,N_13183);
and U19947 (N_19947,N_11623,N_11944);
xor U19948 (N_19948,N_14158,N_12465);
or U19949 (N_19949,N_14714,N_11630);
nand U19950 (N_19950,N_13287,N_14676);
xor U19951 (N_19951,N_12432,N_10251);
xor U19952 (N_19952,N_13088,N_11996);
xor U19953 (N_19953,N_10977,N_12064);
nand U19954 (N_19954,N_12774,N_13906);
nor U19955 (N_19955,N_11510,N_10772);
nor U19956 (N_19956,N_13586,N_13481);
and U19957 (N_19957,N_14132,N_14161);
nand U19958 (N_19958,N_12590,N_14778);
or U19959 (N_19959,N_10338,N_13467);
nor U19960 (N_19960,N_14053,N_10102);
nor U19961 (N_19961,N_10949,N_11615);
and U19962 (N_19962,N_12005,N_13579);
nand U19963 (N_19963,N_11912,N_10197);
or U19964 (N_19964,N_14894,N_10317);
or U19965 (N_19965,N_13286,N_10366);
xnor U19966 (N_19966,N_14953,N_10766);
nor U19967 (N_19967,N_11566,N_11146);
xor U19968 (N_19968,N_11252,N_13676);
nand U19969 (N_19969,N_12897,N_10690);
xor U19970 (N_19970,N_11752,N_13080);
or U19971 (N_19971,N_13191,N_14413);
or U19972 (N_19972,N_13040,N_13515);
nand U19973 (N_19973,N_13885,N_14760);
nor U19974 (N_19974,N_14518,N_10012);
xor U19975 (N_19975,N_14037,N_13506);
nor U19976 (N_19976,N_14816,N_13007);
xnor U19977 (N_19977,N_10348,N_12250);
nor U19978 (N_19978,N_13108,N_14297);
or U19979 (N_19979,N_12821,N_12921);
and U19980 (N_19980,N_14276,N_11789);
and U19981 (N_19981,N_10793,N_11519);
nor U19982 (N_19982,N_12291,N_10243);
nand U19983 (N_19983,N_12912,N_13839);
or U19984 (N_19984,N_14159,N_11258);
nor U19985 (N_19985,N_10124,N_14599);
xor U19986 (N_19986,N_10293,N_11365);
nor U19987 (N_19987,N_14977,N_11415);
nand U19988 (N_19988,N_10001,N_11349);
nor U19989 (N_19989,N_14558,N_13583);
and U19990 (N_19990,N_11596,N_12869);
and U19991 (N_19991,N_10277,N_14376);
nand U19992 (N_19992,N_11355,N_10962);
nor U19993 (N_19993,N_11193,N_12884);
or U19994 (N_19994,N_12504,N_12766);
xnor U19995 (N_19995,N_12970,N_12149);
or U19996 (N_19996,N_12507,N_10859);
or U19997 (N_19997,N_10430,N_14110);
nor U19998 (N_19998,N_13053,N_12782);
and U19999 (N_19999,N_14427,N_10611);
and U20000 (N_20000,N_18439,N_18091);
and U20001 (N_20001,N_16460,N_17265);
or U20002 (N_20002,N_18841,N_16624);
nand U20003 (N_20003,N_19194,N_19575);
or U20004 (N_20004,N_16740,N_18805);
or U20005 (N_20005,N_16509,N_19445);
or U20006 (N_20006,N_19301,N_16614);
nand U20007 (N_20007,N_17300,N_19437);
nor U20008 (N_20008,N_18318,N_17459);
and U20009 (N_20009,N_16407,N_17177);
and U20010 (N_20010,N_15883,N_18932);
xnor U20011 (N_20011,N_16666,N_16898);
nor U20012 (N_20012,N_18814,N_18126);
and U20013 (N_20013,N_17677,N_18326);
nor U20014 (N_20014,N_15246,N_16559);
and U20015 (N_20015,N_16987,N_15845);
xnor U20016 (N_20016,N_15904,N_15214);
xor U20017 (N_20017,N_16020,N_15457);
nor U20018 (N_20018,N_19834,N_16231);
and U20019 (N_20019,N_19990,N_17663);
and U20020 (N_20020,N_18302,N_18227);
nor U20021 (N_20021,N_19610,N_16662);
and U20022 (N_20022,N_16786,N_19162);
or U20023 (N_20023,N_15344,N_19775);
xnor U20024 (N_20024,N_18834,N_15512);
or U20025 (N_20025,N_16441,N_16355);
nor U20026 (N_20026,N_15728,N_18324);
or U20027 (N_20027,N_18109,N_15442);
and U20028 (N_20028,N_16124,N_15239);
nand U20029 (N_20029,N_16145,N_19612);
xor U20030 (N_20030,N_17378,N_15188);
or U20031 (N_20031,N_15645,N_19022);
and U20032 (N_20032,N_16332,N_17056);
xnor U20033 (N_20033,N_16429,N_18680);
nor U20034 (N_20034,N_18849,N_18512);
nand U20035 (N_20035,N_18080,N_17541);
xnor U20036 (N_20036,N_16387,N_16750);
and U20037 (N_20037,N_18392,N_19439);
nand U20038 (N_20038,N_15293,N_17024);
xor U20039 (N_20039,N_18278,N_18463);
or U20040 (N_20040,N_16983,N_19178);
nor U20041 (N_20041,N_15200,N_17255);
xnor U20042 (N_20042,N_17767,N_16045);
nand U20043 (N_20043,N_16270,N_18937);
and U20044 (N_20044,N_16405,N_15921);
nor U20045 (N_20045,N_17866,N_18233);
or U20046 (N_20046,N_15872,N_17421);
or U20047 (N_20047,N_19520,N_19877);
or U20048 (N_20048,N_17293,N_17888);
nor U20049 (N_20049,N_16287,N_19205);
or U20050 (N_20050,N_16591,N_16594);
or U20051 (N_20051,N_19589,N_17340);
nor U20052 (N_20052,N_18986,N_17568);
nand U20053 (N_20053,N_16217,N_16223);
nand U20054 (N_20054,N_18583,N_18017);
nor U20055 (N_20055,N_19550,N_15716);
or U20056 (N_20056,N_17280,N_16367);
xnor U20057 (N_20057,N_18601,N_18428);
xor U20058 (N_20058,N_19149,N_16615);
nor U20059 (N_20059,N_15877,N_17157);
nor U20060 (N_20060,N_17604,N_17722);
and U20061 (N_20061,N_19536,N_16069);
nor U20062 (N_20062,N_18070,N_17458);
xor U20063 (N_20063,N_15220,N_16916);
nand U20064 (N_20064,N_17987,N_19161);
nand U20065 (N_20065,N_17811,N_17558);
nand U20066 (N_20066,N_16753,N_18709);
nor U20067 (N_20067,N_16400,N_18329);
or U20068 (N_20068,N_18801,N_17017);
or U20069 (N_20069,N_15788,N_18315);
xnor U20070 (N_20070,N_16076,N_16868);
and U20071 (N_20071,N_16764,N_16086);
nor U20072 (N_20072,N_19266,N_19286);
and U20073 (N_20073,N_17451,N_19939);
and U20074 (N_20074,N_17662,N_16189);
xor U20075 (N_20075,N_19521,N_16665);
nand U20076 (N_20076,N_15097,N_16580);
or U20077 (N_20077,N_19700,N_15211);
nand U20078 (N_20078,N_15042,N_18090);
nand U20079 (N_20079,N_18536,N_19725);
xor U20080 (N_20080,N_19416,N_16745);
and U20081 (N_20081,N_18177,N_16159);
nand U20082 (N_20082,N_19780,N_18187);
and U20083 (N_20083,N_18589,N_17509);
or U20084 (N_20084,N_18872,N_16238);
and U20085 (N_20085,N_19310,N_16893);
nor U20086 (N_20086,N_18060,N_19261);
xnor U20087 (N_20087,N_16727,N_15977);
nand U20088 (N_20088,N_18573,N_15894);
and U20089 (N_20089,N_18864,N_19446);
nand U20090 (N_20090,N_19914,N_15186);
or U20091 (N_20091,N_15460,N_18621);
nor U20092 (N_20092,N_17788,N_17230);
and U20093 (N_20093,N_18896,N_19692);
or U20094 (N_20094,N_18487,N_16852);
xnor U20095 (N_20095,N_16411,N_19240);
nand U20096 (N_20096,N_15229,N_16891);
nand U20097 (N_20097,N_18241,N_17332);
nand U20098 (N_20098,N_16982,N_18391);
nor U20099 (N_20099,N_15178,N_15858);
nand U20100 (N_20100,N_15676,N_18414);
xnor U20101 (N_20101,N_17596,N_17759);
or U20102 (N_20102,N_17914,N_18173);
and U20103 (N_20103,N_18730,N_16483);
or U20104 (N_20104,N_18618,N_18997);
or U20105 (N_20105,N_17494,N_15011);
nor U20106 (N_20106,N_15114,N_17189);
nand U20107 (N_20107,N_18887,N_16515);
and U20108 (N_20108,N_18321,N_17175);
xnor U20109 (N_20109,N_17702,N_17506);
xor U20110 (N_20110,N_15451,N_15016);
or U20111 (N_20111,N_19385,N_15455);
or U20112 (N_20112,N_18852,N_19702);
or U20113 (N_20113,N_17426,N_18687);
and U20114 (N_20114,N_15181,N_16451);
and U20115 (N_20115,N_16251,N_16301);
xnor U20116 (N_20116,N_17098,N_19994);
nor U20117 (N_20117,N_15829,N_18440);
or U20118 (N_20118,N_16535,N_19985);
nand U20119 (N_20119,N_16129,N_15822);
xnor U20120 (N_20120,N_19010,N_16314);
or U20121 (N_20121,N_17093,N_16830);
or U20122 (N_20122,N_17769,N_18015);
xor U20123 (N_20123,N_15435,N_19360);
or U20124 (N_20124,N_15499,N_18389);
or U20125 (N_20125,N_17739,N_15237);
and U20126 (N_20126,N_17385,N_15218);
and U20127 (N_20127,N_19840,N_16130);
xnor U20128 (N_20128,N_17149,N_18783);
and U20129 (N_20129,N_19561,N_18368);
and U20130 (N_20130,N_18556,N_17998);
xor U20131 (N_20131,N_16005,N_19603);
xnor U20132 (N_20132,N_17354,N_16965);
nor U20133 (N_20133,N_16345,N_16219);
or U20134 (N_20134,N_16437,N_15621);
nand U20135 (N_20135,N_16257,N_17926);
nor U20136 (N_20136,N_15545,N_19324);
and U20137 (N_20137,N_15202,N_17855);
xor U20138 (N_20138,N_17617,N_16225);
nor U20139 (N_20139,N_19498,N_17441);
or U20140 (N_20140,N_17873,N_16139);
nand U20141 (N_20141,N_18279,N_16310);
nand U20142 (N_20142,N_15539,N_19951);
xor U20143 (N_20143,N_18599,N_17348);
xor U20144 (N_20144,N_15837,N_15167);
or U20145 (N_20145,N_18271,N_18784);
or U20146 (N_20146,N_15007,N_16178);
nand U20147 (N_20147,N_16403,N_16165);
and U20148 (N_20148,N_19027,N_16508);
or U20149 (N_20149,N_15027,N_15698);
and U20150 (N_20150,N_18811,N_16705);
xnor U20151 (N_20151,N_16929,N_18584);
nor U20152 (N_20152,N_19225,N_17133);
xnor U20153 (N_20153,N_17813,N_18336);
nand U20154 (N_20154,N_16681,N_19584);
xor U20155 (N_20155,N_15169,N_16833);
xnor U20156 (N_20156,N_19433,N_15009);
nor U20157 (N_20157,N_19228,N_17766);
or U20158 (N_20158,N_19312,N_19798);
nand U20159 (N_20159,N_19136,N_19763);
and U20160 (N_20160,N_18421,N_19978);
or U20161 (N_20161,N_19676,N_19703);
xor U20162 (N_20162,N_18685,N_18266);
xnor U20163 (N_20163,N_17642,N_15475);
and U20164 (N_20164,N_16099,N_16192);
xnor U20165 (N_20165,N_18275,N_16391);
and U20166 (N_20166,N_16643,N_18384);
nor U20167 (N_20167,N_17307,N_18224);
and U20168 (N_20168,N_15331,N_15652);
nor U20169 (N_20169,N_16561,N_18410);
nand U20170 (N_20170,N_16773,N_16708);
and U20171 (N_20171,N_18980,N_15930);
and U20172 (N_20172,N_16686,N_17960);
nor U20173 (N_20173,N_18359,N_17867);
and U20174 (N_20174,N_17762,N_19921);
or U20175 (N_20175,N_15774,N_19256);
xnor U20176 (N_20176,N_15775,N_16731);
or U20177 (N_20177,N_16656,N_18218);
or U20178 (N_20178,N_15340,N_16055);
or U20179 (N_20179,N_19835,N_18020);
nor U20180 (N_20180,N_15074,N_16679);
nand U20181 (N_20181,N_17887,N_19146);
or U20182 (N_20182,N_15642,N_18299);
and U20183 (N_20183,N_18395,N_16562);
and U20184 (N_20184,N_18148,N_18375);
and U20185 (N_20185,N_16133,N_16867);
xor U20186 (N_20186,N_19335,N_16973);
nand U20187 (N_20187,N_16938,N_16966);
nor U20188 (N_20188,N_19338,N_17893);
nor U20189 (N_20189,N_15908,N_15917);
nand U20190 (N_20190,N_19899,N_15313);
and U20191 (N_20191,N_18047,N_15315);
and U20192 (N_20192,N_19747,N_19783);
or U20193 (N_20193,N_17163,N_18050);
xnor U20194 (N_20194,N_17972,N_17609);
and U20195 (N_20195,N_18602,N_16034);
and U20196 (N_20196,N_17550,N_19483);
and U20197 (N_20197,N_19327,N_16854);
xnor U20198 (N_20198,N_18298,N_18721);
xnor U20199 (N_20199,N_17949,N_17969);
nor U20200 (N_20200,N_16101,N_15948);
or U20201 (N_20201,N_15969,N_18360);
xor U20202 (N_20202,N_19341,N_16632);
and U20203 (N_20203,N_15907,N_17288);
nand U20204 (N_20204,N_19611,N_18429);
nand U20205 (N_20205,N_15725,N_16644);
xnor U20206 (N_20206,N_19343,N_19267);
or U20207 (N_20207,N_19428,N_19894);
and U20208 (N_20208,N_19631,N_19373);
and U20209 (N_20209,N_19019,N_17401);
or U20210 (N_20210,N_16790,N_15497);
xnor U20211 (N_20211,N_15528,N_18972);
nand U20212 (N_20212,N_16774,N_15143);
and U20213 (N_20213,N_17925,N_17437);
nor U20214 (N_20214,N_15436,N_19245);
and U20215 (N_20215,N_18962,N_15098);
nor U20216 (N_20216,N_18288,N_17194);
or U20217 (N_20217,N_15556,N_15132);
nand U20218 (N_20218,N_19505,N_18403);
nor U20219 (N_20219,N_18055,N_16956);
xnor U20220 (N_20220,N_17695,N_15933);
nand U20221 (N_20221,N_15940,N_16673);
nor U20222 (N_20222,N_15941,N_15189);
xor U20223 (N_20223,N_19082,N_15047);
xnor U20224 (N_20224,N_17368,N_19793);
and U20225 (N_20225,N_19500,N_18434);
or U20226 (N_20226,N_18374,N_15006);
nor U20227 (N_20227,N_17383,N_17874);
xnor U20228 (N_20228,N_17329,N_15136);
nor U20229 (N_20229,N_17886,N_16357);
nand U20230 (N_20230,N_19784,N_18955);
nand U20231 (N_20231,N_16970,N_18470);
and U20232 (N_20232,N_16649,N_17755);
nand U20233 (N_20233,N_18994,N_18307);
and U20234 (N_20234,N_18917,N_15892);
nand U20235 (N_20235,N_15374,N_15013);
or U20236 (N_20236,N_17222,N_19996);
or U20237 (N_20237,N_16992,N_19815);
nand U20238 (N_20238,N_19912,N_16877);
nor U20239 (N_20239,N_15334,N_16195);
xor U20240 (N_20240,N_17190,N_15778);
xnor U20241 (N_20241,N_17211,N_16904);
nor U20242 (N_20242,N_16486,N_15381);
and U20243 (N_20243,N_18675,N_16366);
or U20244 (N_20244,N_18873,N_16191);
nor U20245 (N_20245,N_15626,N_15974);
nor U20246 (N_20246,N_17948,N_16828);
and U20247 (N_20247,N_17823,N_17658);
or U20248 (N_20248,N_15665,N_19002);
or U20249 (N_20249,N_17266,N_16894);
nand U20250 (N_20250,N_15723,N_19845);
or U20251 (N_20251,N_17899,N_16393);
or U20252 (N_20252,N_18198,N_18041);
nor U20253 (N_20253,N_19903,N_17796);
and U20254 (N_20254,N_19318,N_15059);
xnor U20255 (N_20255,N_19348,N_16272);
and U20256 (N_20256,N_15543,N_17725);
xnor U20257 (N_20257,N_15316,N_15719);
or U20258 (N_20258,N_17560,N_15663);
xnor U20259 (N_20259,N_15889,N_19544);
nor U20260 (N_20260,N_15477,N_19976);
and U20261 (N_20261,N_16853,N_19907);
nand U20262 (N_20262,N_17598,N_16637);
nor U20263 (N_20263,N_16876,N_19089);
nand U20264 (N_20264,N_17352,N_16621);
xnor U20265 (N_20265,N_16744,N_17913);
or U20266 (N_20266,N_17894,N_16839);
nor U20267 (N_20267,N_15309,N_19151);
nand U20268 (N_20268,N_18567,N_18492);
and U20269 (N_20269,N_15343,N_19797);
and U20270 (N_20270,N_15292,N_16638);
or U20271 (N_20271,N_15996,N_15876);
xnor U20272 (N_20272,N_17216,N_19191);
nand U20273 (N_20273,N_17828,N_18740);
or U20274 (N_20274,N_19470,N_18978);
nand U20275 (N_20275,N_15773,N_18503);
nand U20276 (N_20276,N_16430,N_18232);
and U20277 (N_20277,N_16019,N_16013);
or U20278 (N_20278,N_15993,N_17798);
nor U20279 (N_20279,N_15681,N_16211);
nor U20280 (N_20280,N_15958,N_19760);
xor U20281 (N_20281,N_17636,N_19268);
or U20282 (N_20282,N_19135,N_18798);
nor U20283 (N_20283,N_17433,N_18136);
xnor U20284 (N_20284,N_19102,N_15113);
xnor U20285 (N_20285,N_16748,N_18682);
xor U20286 (N_20286,N_18130,N_17967);
and U20287 (N_20287,N_18040,N_16556);
nand U20288 (N_20288,N_16131,N_19396);
nand U20289 (N_20289,N_17158,N_15414);
and U20290 (N_20290,N_16824,N_16382);
xor U20291 (N_20291,N_16497,N_15732);
nand U20292 (N_20292,N_19790,N_16942);
or U20293 (N_20293,N_18982,N_17167);
nand U20294 (N_20294,N_18386,N_16514);
or U20295 (N_20295,N_18046,N_17736);
or U20296 (N_20296,N_15540,N_17993);
or U20297 (N_20297,N_15857,N_17308);
xnor U20298 (N_20298,N_16140,N_15932);
or U20299 (N_20299,N_18444,N_15995);
or U20300 (N_20300,N_18546,N_16995);
nor U20301 (N_20301,N_15817,N_15861);
nor U20302 (N_20302,N_16613,N_15588);
and U20303 (N_20303,N_16125,N_19965);
xnor U20304 (N_20304,N_18427,N_17109);
or U20305 (N_20305,N_18231,N_15741);
or U20306 (N_20306,N_17675,N_19946);
xnor U20307 (N_20307,N_15280,N_15730);
and U20308 (N_20308,N_15312,N_17192);
and U20309 (N_20309,N_18537,N_15464);
nor U20310 (N_20310,N_19252,N_17810);
nand U20311 (N_20311,N_15580,N_15804);
nand U20312 (N_20312,N_19863,N_17072);
xor U20313 (N_20313,N_19473,N_16421);
xnor U20314 (N_20314,N_17427,N_16531);
xor U20315 (N_20315,N_18971,N_19956);
or U20316 (N_20316,N_18825,N_15498);
xnor U20317 (N_20317,N_19992,N_16915);
nand U20318 (N_20318,N_19600,N_16447);
and U20319 (N_20319,N_19525,N_17720);
or U20320 (N_20320,N_18312,N_19805);
and U20321 (N_20321,N_16245,N_19697);
or U20322 (N_20322,N_15036,N_19031);
xnor U20323 (N_20323,N_18480,N_16385);
or U20324 (N_20324,N_18793,N_19055);
or U20325 (N_20325,N_17703,N_19534);
nand U20326 (N_20326,N_17172,N_17452);
or U20327 (N_20327,N_17398,N_19636);
or U20328 (N_20328,N_16470,N_17424);
nor U20329 (N_20329,N_15207,N_18471);
and U20330 (N_20330,N_19645,N_15926);
nand U20331 (N_20331,N_15350,N_16431);
nand U20332 (N_20332,N_15501,N_18133);
or U20333 (N_20333,N_19113,N_19140);
nand U20334 (N_20334,N_16517,N_17145);
nor U20335 (N_20335,N_15997,N_19734);
and U20336 (N_20336,N_17325,N_19443);
nand U20337 (N_20337,N_16048,N_15938);
or U20338 (N_20338,N_16454,N_18308);
nor U20339 (N_20339,N_16793,N_16742);
nor U20340 (N_20340,N_18727,N_19842);
and U20341 (N_20341,N_16949,N_19867);
or U20342 (N_20342,N_15001,N_16906);
or U20343 (N_20343,N_17814,N_15251);
nor U20344 (N_20344,N_19238,N_19208);
xnor U20345 (N_20345,N_15506,N_18807);
xnor U20346 (N_20346,N_18089,N_16701);
or U20347 (N_20347,N_15401,N_16127);
or U20348 (N_20348,N_17328,N_17513);
or U20349 (N_20349,N_17333,N_19761);
and U20350 (N_20350,N_17182,N_16694);
xor U20351 (N_20351,N_18373,N_19599);
nor U20352 (N_20352,N_18472,N_15939);
and U20353 (N_20353,N_15361,N_16611);
and U20354 (N_20354,N_18426,N_19316);
nor U20355 (N_20355,N_17330,N_16897);
nor U20356 (N_20356,N_16081,N_17771);
and U20357 (N_20357,N_19107,N_16475);
or U20358 (N_20358,N_18767,N_16880);
xor U20359 (N_20359,N_17953,N_15777);
nor U20360 (N_20360,N_17344,N_16683);
nand U20361 (N_20361,N_16575,N_18711);
and U20362 (N_20362,N_19386,N_18792);
xnor U20363 (N_20363,N_16714,N_15602);
xnor U20364 (N_20364,N_16888,N_15609);
and U20365 (N_20365,N_18816,N_17464);
and U20366 (N_20366,N_15409,N_17497);
xor U20367 (N_20367,N_15250,N_17876);
nor U20368 (N_20368,N_19742,N_16602);
nand U20369 (N_20369,N_19651,N_16106);
xnor U20370 (N_20370,N_16709,N_15577);
or U20371 (N_20371,N_18839,N_16100);
nand U20372 (N_20372,N_18992,N_17865);
xor U20373 (N_20373,N_16379,N_16491);
or U20374 (N_20374,N_16703,N_17089);
nand U20375 (N_20375,N_19481,N_17460);
or U20376 (N_20376,N_18249,N_18129);
nand U20377 (N_20377,N_15647,N_16592);
xnor U20378 (N_20378,N_17225,N_15934);
nand U20379 (N_20379,N_18975,N_18750);
or U20380 (N_20380,N_19756,N_18703);
nor U20381 (N_20381,N_15884,N_16255);
and U20382 (N_20382,N_19024,N_17779);
nand U20383 (N_20383,N_19961,N_15418);
xnor U20384 (N_20384,N_17065,N_18757);
xnor U20385 (N_20385,N_19421,N_15541);
or U20386 (N_20386,N_15023,N_19011);
xnor U20387 (N_20387,N_19998,N_19401);
nor U20388 (N_20388,N_19478,N_15240);
xor U20389 (N_20389,N_19900,N_16619);
nand U20390 (N_20390,N_16699,N_19145);
and U20391 (N_20391,N_15650,N_15266);
nor U20392 (N_20392,N_16248,N_16678);
and U20393 (N_20393,N_16801,N_15763);
nor U20394 (N_20394,N_19803,N_19617);
or U20395 (N_20395,N_18388,N_19451);
and U20396 (N_20396,N_15289,N_19736);
or U20397 (N_20397,N_16845,N_17066);
nand U20398 (N_20398,N_19079,N_16826);
or U20399 (N_20399,N_18137,N_15641);
nor U20400 (N_20400,N_17327,N_15620);
nor U20401 (N_20401,N_15784,N_18998);
and U20402 (N_20402,N_17461,N_18406);
nor U20403 (N_20403,N_17060,N_19352);
nor U20404 (N_20404,N_15893,N_15086);
or U20405 (N_20405,N_17534,N_17439);
nor U20406 (N_20406,N_16882,N_17900);
and U20407 (N_20407,N_16031,N_15310);
xnor U20408 (N_20408,N_15514,N_19185);
xnor U20409 (N_20409,N_18624,N_19229);
nor U20410 (N_20410,N_16374,N_17188);
nand U20411 (N_20411,N_19657,N_16754);
or U20412 (N_20412,N_19259,N_18003);
xor U20413 (N_20413,N_17585,N_18035);
or U20414 (N_20414,N_18422,N_18533);
nor U20415 (N_20415,N_18781,N_19785);
xnor U20416 (N_20416,N_17369,N_15991);
and U20417 (N_20417,N_18666,N_18030);
xor U20418 (N_20418,N_18604,N_18735);
or U20419 (N_20419,N_15349,N_19576);
or U20420 (N_20420,N_16163,N_18945);
or U20421 (N_20421,N_17517,N_15112);
nor U20422 (N_20422,N_17927,N_19494);
nand U20423 (N_20423,N_16693,N_19850);
nand U20424 (N_20424,N_16655,N_16291);
nand U20425 (N_20425,N_18715,N_18548);
nor U20426 (N_20426,N_15819,N_18119);
nor U20427 (N_20427,N_16767,N_19271);
nand U20428 (N_20428,N_17870,N_15749);
xnor U20429 (N_20429,N_15824,N_18493);
and U20430 (N_20430,N_17890,N_18963);
xnor U20431 (N_20431,N_16293,N_15582);
and U20432 (N_20432,N_17081,N_18954);
nor U20433 (N_20433,N_18303,N_19980);
nand U20434 (N_20434,N_18262,N_16654);
xor U20435 (N_20435,N_19744,N_19937);
nand U20436 (N_20436,N_16971,N_17103);
or U20437 (N_20437,N_15664,N_19226);
xor U20438 (N_20438,N_18154,N_19332);
or U20439 (N_20439,N_15172,N_15760);
nand U20440 (N_20440,N_17976,N_17033);
or U20441 (N_20441,N_15886,N_18613);
nor U20442 (N_20442,N_18322,N_16011);
nor U20443 (N_20443,N_16532,N_18018);
nor U20444 (N_20444,N_19776,N_18762);
xor U20445 (N_20445,N_15233,N_16462);
or U20446 (N_20446,N_18333,N_17481);
nor U20447 (N_20447,N_19731,N_17078);
xnor U20448 (N_20448,N_19526,N_16817);
or U20449 (N_20449,N_17819,N_15102);
nand U20450 (N_20450,N_17723,N_15568);
nand U20451 (N_20451,N_17709,N_16490);
nand U20452 (N_20452,N_15300,N_16577);
nor U20453 (N_20453,N_16813,N_19732);
nor U20454 (N_20454,N_17850,N_15511);
nand U20455 (N_20455,N_19876,N_19699);
nor U20456 (N_20456,N_17244,N_17715);
xnor U20457 (N_20457,N_18032,N_15285);
and U20458 (N_20458,N_18092,N_19025);
and U20459 (N_20459,N_16972,N_16485);
xor U20460 (N_20460,N_18836,N_16242);
or U20461 (N_20461,N_16737,N_15944);
or U20462 (N_20462,N_16797,N_17734);
nor U20463 (N_20463,N_18698,N_19183);
xor U20464 (N_20464,N_15885,N_17841);
or U20465 (N_20465,N_19224,N_15306);
nor U20466 (N_20466,N_15177,N_18436);
and U20467 (N_20467,N_17220,N_19195);
and U20468 (N_20468,N_16534,N_15038);
xnor U20469 (N_20469,N_15619,N_19581);
xnor U20470 (N_20470,N_16056,N_16675);
nand U20471 (N_20471,N_19688,N_19647);
nand U20472 (N_20472,N_18327,N_16118);
or U20473 (N_20473,N_15254,N_15744);
or U20474 (N_20474,N_18382,N_16598);
xor U20475 (N_20475,N_18116,N_16202);
nand U20476 (N_20476,N_18842,N_19853);
or U20477 (N_20477,N_15551,N_16981);
or U20478 (N_20478,N_19673,N_17986);
nand U20479 (N_20479,N_15679,N_19328);
nor U20480 (N_20480,N_15058,N_16563);
or U20481 (N_20481,N_19197,N_18710);
nand U20482 (N_20482,N_16337,N_17203);
xor U20483 (N_20483,N_17286,N_16024);
or U20484 (N_20484,N_18891,N_17834);
and U20485 (N_20485,N_19051,N_19317);
nand U20486 (N_20486,N_15605,N_16176);
nor U20487 (N_20487,N_17510,N_19114);
nand U20488 (N_20488,N_17666,N_19460);
xnor U20489 (N_20489,N_15649,N_18534);
nand U20490 (N_20490,N_19144,N_17571);
xor U20491 (N_20491,N_15219,N_18876);
and U20492 (N_20492,N_15373,N_16885);
nand U20493 (N_20493,N_18587,N_17667);
nor U20494 (N_20494,N_17895,N_15794);
xor U20495 (N_20495,N_16073,N_19242);
nor U20496 (N_20496,N_16639,N_16997);
nand U20497 (N_20497,N_18242,N_16871);
nand U20498 (N_20498,N_16484,N_17345);
nand U20499 (N_20499,N_15928,N_17240);
nor U20500 (N_20500,N_16103,N_19908);
nor U20501 (N_20501,N_16554,N_18027);
and U20502 (N_20502,N_16346,N_16586);
xor U20503 (N_20503,N_15524,N_19806);
nand U20504 (N_20504,N_16779,N_17444);
xor U20505 (N_20505,N_19694,N_18598);
xnor U20506 (N_20506,N_17012,N_19564);
xor U20507 (N_20507,N_17320,N_17941);
nand U20508 (N_20508,N_17489,N_15715);
or U20509 (N_20509,N_17282,N_16229);
xnor U20510 (N_20510,N_18006,N_19442);
nand U20511 (N_20511,N_16803,N_17136);
nand U20512 (N_20512,N_18419,N_19538);
or U20513 (N_20513,N_17978,N_16695);
or U20514 (N_20514,N_16620,N_16725);
xor U20515 (N_20515,N_17100,N_16110);
and U20516 (N_20516,N_18699,N_18771);
nand U20517 (N_20517,N_18810,N_17799);
nor U20518 (N_20518,N_16224,N_17974);
nor U20519 (N_20519,N_19549,N_15028);
nor U20520 (N_20520,N_19201,N_18756);
nor U20521 (N_20521,N_18616,N_16664);
or U20522 (N_20522,N_17782,N_15459);
and U20523 (N_20523,N_15117,N_19983);
xor U20524 (N_20524,N_18052,N_15421);
nor U20525 (N_20525,N_15426,N_16896);
xor U20526 (N_20526,N_17933,N_18269);
nand U20527 (N_20527,N_17097,N_19378);
or U20528 (N_20528,N_19875,N_15610);
or U20529 (N_20529,N_18076,N_18667);
or U20530 (N_20530,N_18549,N_16089);
or U20531 (N_20531,N_16404,N_16246);
and U20532 (N_20532,N_18600,N_15687);
nand U20533 (N_20533,N_19816,N_18889);
or U20534 (N_20534,N_16213,N_15868);
nor U20535 (N_20535,N_18733,N_16849);
nor U20536 (N_20536,N_17829,N_15005);
or U20537 (N_20537,N_17035,N_17334);
xor U20538 (N_20538,N_19362,N_16571);
nand U20539 (N_20539,N_16600,N_17871);
nor U20540 (N_20540,N_19609,N_17215);
or U20541 (N_20541,N_17655,N_15276);
xor U20542 (N_20542,N_18305,N_17085);
and U20543 (N_20543,N_17797,N_16342);
or U20544 (N_20544,N_15428,N_18902);
nor U20545 (N_20545,N_18831,N_17673);
nor U20546 (N_20546,N_18246,N_17685);
nor U20547 (N_20547,N_18862,N_18936);
nand U20548 (N_20548,N_17698,N_17456);
or U20549 (N_20549,N_15430,N_15927);
nand U20550 (N_20550,N_18704,N_18916);
xor U20551 (N_20551,N_17906,N_16996);
xnor U20552 (N_20552,N_18656,N_15734);
xor U20553 (N_20553,N_15816,N_16667);
or U20554 (N_20554,N_19787,N_19585);
nor U20555 (N_20555,N_19374,N_16260);
nand U20556 (N_20556,N_15077,N_17746);
nor U20557 (N_20557,N_16609,N_15859);
and U20558 (N_20558,N_19833,N_16785);
or U20559 (N_20559,N_16668,N_17069);
and U20560 (N_20560,N_17486,N_17859);
xor U20561 (N_20561,N_16459,N_19906);
nor U20562 (N_20562,N_19003,N_16477);
or U20563 (N_20563,N_16834,N_16147);
nor U20564 (N_20564,N_18164,N_15213);
nand U20565 (N_20565,N_17338,N_19772);
nand U20566 (N_20566,N_19913,N_17749);
xor U20567 (N_20567,N_18474,N_15532);
or U20568 (N_20568,N_18668,N_18201);
xnor U20569 (N_20569,N_18568,N_18181);
and U20570 (N_20570,N_19206,N_15767);
nand U20571 (N_20571,N_16151,N_15277);
nor U20572 (N_20572,N_19757,N_16295);
nor U20573 (N_20573,N_18499,N_16170);
and U20574 (N_20574,N_15203,N_17405);
or U20575 (N_20575,N_19765,N_19471);
or U20576 (N_20576,N_18505,N_18960);
or U20577 (N_20577,N_16095,N_19711);
xnor U20578 (N_20578,N_15891,N_17030);
xnor U20579 (N_20579,N_19495,N_15454);
xnor U20580 (N_20580,N_17579,N_17693);
or U20581 (N_20581,N_15412,N_16861);
and U20582 (N_20582,N_15090,N_15107);
and U20583 (N_20583,N_19417,N_17943);
or U20584 (N_20584,N_19094,N_18462);
nand U20585 (N_20585,N_15092,N_17968);
nor U20586 (N_20586,N_19217,N_15466);
nor U20587 (N_20587,N_17731,N_18310);
or U20588 (N_20588,N_19943,N_15273);
and U20589 (N_20589,N_18100,N_19364);
nand U20590 (N_20590,N_17138,N_17839);
or U20591 (N_20591,N_15558,N_18078);
nand U20592 (N_20592,N_19159,N_15615);
nand U20593 (N_20593,N_15397,N_16901);
xor U20594 (N_20594,N_16576,N_17966);
or U20595 (N_20595,N_18478,N_17463);
and U20596 (N_20596,N_16492,N_15699);
xnor U20597 (N_20597,N_16263,N_18029);
nand U20598 (N_20598,N_15998,N_19810);
xnor U20599 (N_20599,N_18654,N_15231);
and U20600 (N_20600,N_19047,N_17751);
nand U20601 (N_20601,N_15981,N_16372);
nor U20602 (N_20602,N_17279,N_16927);
or U20603 (N_20603,N_16209,N_16313);
or U20604 (N_20604,N_15400,N_16062);
and U20605 (N_20605,N_19213,N_17540);
and U20606 (N_20606,N_18104,N_16503);
or U20607 (N_20607,N_17742,N_19628);
and U20608 (N_20608,N_18605,N_19970);
or U20609 (N_20609,N_18926,N_18061);
nand U20610 (N_20610,N_18496,N_19289);
and U20611 (N_20611,N_18005,N_16236);
nor U20612 (N_20612,N_19361,N_15278);
and U20613 (N_20613,N_18208,N_16302);
or U20614 (N_20614,N_15882,N_16286);
xnor U20615 (N_20615,N_17611,N_18168);
and U20616 (N_20616,N_17745,N_18511);
nand U20617 (N_20617,N_19447,N_15030);
xnor U20618 (N_20618,N_17932,N_15425);
nor U20619 (N_20619,N_18644,N_18135);
xnor U20620 (N_20620,N_15127,N_18959);
or U20621 (N_20621,N_19095,N_18967);
and U20622 (N_20622,N_18753,N_17010);
or U20623 (N_20623,N_15362,N_17246);
or U20624 (N_20624,N_19302,N_17519);
xor U20625 (N_20625,N_17111,N_17707);
nand U20626 (N_20626,N_15324,N_16855);
nor U20627 (N_20627,N_17638,N_15584);
or U20628 (N_20628,N_17312,N_16757);
and U20629 (N_20629,N_16889,N_15356);
or U20630 (N_20630,N_19368,N_16746);
and U20631 (N_20631,N_17945,N_17047);
xnor U20632 (N_20632,N_16415,N_17530);
nand U20633 (N_20633,N_18267,N_19061);
and U20634 (N_20634,N_19357,N_17438);
nand U20635 (N_20635,N_17400,N_18313);
nor U20636 (N_20636,N_19618,N_18014);
xnor U20637 (N_20637,N_19370,N_15875);
or U20638 (N_20638,N_18466,N_15458);
nor U20639 (N_20639,N_15470,N_18590);
or U20640 (N_20640,N_15546,N_19038);
xnor U20641 (N_20641,N_16325,N_17962);
nand U20642 (N_20642,N_15881,N_15085);
and U20643 (N_20643,N_19988,N_16296);
nor U20644 (N_20644,N_17275,N_18769);
nand U20645 (N_20645,N_15351,N_15299);
and U20646 (N_20646,N_16340,N_15929);
and U20647 (N_20647,N_18996,N_17818);
or U20648 (N_20648,N_15746,N_17479);
nor U20649 (N_20649,N_19037,N_19555);
nor U20650 (N_20650,N_19701,N_15740);
nor U20651 (N_20651,N_16277,N_17415);
or U20652 (N_20652,N_16890,N_15795);
and U20653 (N_20653,N_18099,N_18525);
nand U20654 (N_20654,N_15726,N_15429);
or U20655 (N_20655,N_16818,N_19233);
and U20656 (N_20656,N_15637,N_15046);
or U20657 (N_20657,N_16409,N_16783);
nand U20658 (N_20658,N_16537,N_19488);
and U20659 (N_20659,N_16440,N_15624);
xnor U20660 (N_20660,N_17599,N_17951);
nand U20661 (N_20661,N_19604,N_17794);
nand U20662 (N_20662,N_17614,N_15660);
nand U20663 (N_20663,N_16608,N_19587);
nand U20664 (N_20664,N_16669,N_15108);
nand U20665 (N_20665,N_16528,N_15737);
nand U20666 (N_20666,N_18460,N_16321);
nor U20667 (N_20667,N_17692,N_19935);
nor U20668 (N_20668,N_16541,N_17919);
nor U20669 (N_20669,N_18287,N_17276);
or U20670 (N_20670,N_15919,N_16749);
nor U20671 (N_20671,N_19689,N_19333);
xor U20672 (N_20672,N_19232,N_17262);
and U20673 (N_20673,N_16928,N_19847);
nand U20674 (N_20674,N_16707,N_19573);
nand U20675 (N_20675,N_16692,N_19663);
nand U20676 (N_20676,N_17815,N_16523);
or U20677 (N_20677,N_16227,N_19690);
or U20678 (N_20678,N_19231,N_15603);
xnor U20679 (N_20679,N_15835,N_19565);
or U20680 (N_20680,N_16597,N_17995);
xnor U20681 (N_20681,N_19795,N_16025);
nor U20682 (N_20682,N_16544,N_18057);
xnor U20683 (N_20683,N_17733,N_16820);
and U20684 (N_20684,N_15887,N_15371);
xnor U20685 (N_20685,N_15096,N_19448);
xor U20686 (N_20686,N_15208,N_17184);
and U20687 (N_20687,N_15825,N_16250);
nand U20688 (N_20688,N_15983,N_19786);
nand U20689 (N_20689,N_17689,N_19743);
xor U20690 (N_20690,N_17591,N_16502);
or U20691 (N_20691,N_15682,N_16173);
nor U20692 (N_20692,N_19295,N_16653);
xnor U20693 (N_20693,N_17981,N_19671);
or U20694 (N_20694,N_18485,N_18108);
xnor U20695 (N_20695,N_15326,N_17587);
nor U20696 (N_20696,N_16569,N_19595);
nand U20697 (N_20697,N_15444,N_19043);
nor U20698 (N_20698,N_16606,N_15192);
or U20699 (N_20699,N_16042,N_17039);
and U20700 (N_20700,N_17659,N_17198);
xnor U20701 (N_20701,N_18362,N_18648);
or U20702 (N_20702,N_17862,N_17935);
nand U20703 (N_20703,N_19296,N_15297);
or U20704 (N_20704,N_17653,N_16950);
nor U20705 (N_20705,N_15869,N_15537);
and U20706 (N_20706,N_16874,N_17840);
and U20707 (N_20707,N_15531,N_15149);
xor U20708 (N_20708,N_16706,N_16892);
nor U20709 (N_20709,N_18068,N_15901);
or U20710 (N_20710,N_17973,N_18942);
nand U20711 (N_20711,N_18664,N_18416);
xnor U20712 (N_20712,N_18433,N_15375);
or U20713 (N_20713,N_17690,N_15792);
and U20714 (N_20714,N_17143,N_19129);
nor U20715 (N_20715,N_19406,N_19727);
nor U20716 (N_20716,N_18625,N_17507);
and U20717 (N_20717,N_19932,N_15187);
or U20718 (N_20718,N_17958,N_16581);
xnor U20719 (N_20719,N_17337,N_16550);
nor U20720 (N_20720,N_16612,N_16276);
xnor U20721 (N_20721,N_19234,N_19602);
nand U20722 (N_20722,N_15492,N_18199);
nand U20723 (N_20723,N_16789,N_18910);
xor U20724 (N_20724,N_15508,N_16064);
or U20725 (N_20725,N_19502,N_15713);
or U20726 (N_20726,N_16262,N_18274);
nand U20727 (N_20727,N_17173,N_15643);
xnor U20728 (N_20728,N_19822,N_16338);
xnor U20729 (N_20729,N_17036,N_16827);
xor U20730 (N_20730,N_19394,N_15843);
nand U20731 (N_20731,N_15705,N_18919);
or U20732 (N_20732,N_15076,N_19029);
nor U20733 (N_20733,N_16001,N_16121);
and U20734 (N_20734,N_19836,N_16658);
and U20735 (N_20735,N_19843,N_19838);
nor U20736 (N_20736,N_19160,N_17055);
and U20737 (N_20737,N_16909,N_18947);
nand U20738 (N_20738,N_19096,N_16822);
xnor U20739 (N_20739,N_17744,N_18044);
or U20740 (N_20740,N_15377,N_18171);
or U20741 (N_20741,N_15286,N_17038);
xnor U20742 (N_20742,N_19175,N_15406);
or U20743 (N_20743,N_16741,N_17061);
and U20744 (N_20744,N_18170,N_18900);
nand U20745 (N_20745,N_17555,N_16526);
or U20746 (N_20746,N_15384,N_16419);
nor U20747 (N_20747,N_16525,N_15606);
or U20748 (N_20748,N_19280,N_15798);
xor U20749 (N_20749,N_18342,N_19883);
or U20750 (N_20750,N_16132,N_17016);
nand U20751 (N_20751,N_15680,N_18167);
nor U20752 (N_20752,N_17005,N_15507);
nor U20753 (N_20753,N_19030,N_15393);
nand U20754 (N_20754,N_16960,N_16098);
nor U20755 (N_20755,N_15693,N_18530);
nand U20756 (N_20756,N_17059,N_18476);
or U20757 (N_20757,N_19080,N_17117);
nand U20758 (N_20758,N_15831,N_16030);
xor U20759 (N_20759,N_17860,N_15402);
or U20760 (N_20760,N_18929,N_19730);
nand U20761 (N_20761,N_15139,N_19487);
nand U20762 (N_20762,N_17128,N_18351);
nand U20763 (N_20763,N_15724,N_17397);
nand U20764 (N_20764,N_19659,N_17801);
and U20765 (N_20765,N_19720,N_16146);
nand U20766 (N_20766,N_17525,N_18036);
or U20767 (N_20767,N_19199,N_18746);
nor U20768 (N_20768,N_17372,N_17000);
and U20769 (N_20769,N_16386,N_17727);
and U20770 (N_20770,N_18669,N_15048);
or U20771 (N_20771,N_17436,N_19666);
and U20772 (N_20772,N_19110,N_19832);
nand U20773 (N_20773,N_18454,N_17272);
nand U20774 (N_20774,N_17411,N_15962);
nand U20775 (N_20775,N_17916,N_19915);
nand U20776 (N_20776,N_18120,N_16218);
nor U20777 (N_20777,N_16150,N_18033);
nor U20778 (N_20778,N_18131,N_18204);
nand U20779 (N_20779,N_19898,N_19143);
or U20780 (N_20780,N_19336,N_18335);
or U20781 (N_20781,N_19590,N_16584);
or U20782 (N_20782,N_19453,N_15554);
nor U20783 (N_20783,N_17704,N_17857);
nand U20784 (N_20784,N_17045,N_17168);
or U20785 (N_20785,N_16539,N_16676);
xor U20786 (N_20786,N_18059,N_16540);
and U20787 (N_20787,N_18286,N_15052);
nand U20788 (N_20788,N_19737,N_15700);
nor U20789 (N_20789,N_19684,N_17310);
xnor U20790 (N_20790,N_15559,N_17237);
nor U20791 (N_20791,N_17880,N_17249);
nand U20792 (N_20792,N_15572,N_18450);
or U20793 (N_20793,N_15612,N_17546);
nor U20794 (N_20794,N_15201,N_15979);
nand U20795 (N_20795,N_19808,N_15931);
or U20796 (N_20796,N_15971,N_15216);
and U20797 (N_20797,N_16593,N_19804);
or U20798 (N_20798,N_18398,N_17567);
and U20799 (N_20799,N_19739,N_19895);
or U20800 (N_20800,N_19969,N_15469);
or U20801 (N_20801,N_19411,N_16353);
and U20802 (N_20802,N_15345,N_17793);
or U20803 (N_20803,N_15493,N_16905);
nor U20804 (N_20804,N_17795,N_16009);
and U20805 (N_20805,N_18285,N_19427);
xnor U20806 (N_20806,N_18211,N_17197);
and U20807 (N_20807,N_16388,N_18854);
and U20808 (N_20808,N_16206,N_15039);
and U20809 (N_20809,N_18585,N_19254);
or U20810 (N_20810,N_17646,N_18357);
xnor U20811 (N_20811,N_17153,N_15026);
and U20812 (N_20812,N_19053,N_19342);
and U20813 (N_20813,N_16261,N_19365);
or U20814 (N_20814,N_19260,N_16816);
nor U20815 (N_20815,N_16128,N_15376);
and U20816 (N_20816,N_17139,N_15812);
nor U20817 (N_20817,N_18330,N_15411);
and U20818 (N_20818,N_16384,N_16334);
nor U20819 (N_20819,N_17592,N_19817);
nand U20820 (N_20820,N_16237,N_15259);
or U20821 (N_20821,N_19968,N_17301);
or U20822 (N_20822,N_17622,N_19290);
nor U20823 (N_20823,N_19771,N_18064);
or U20824 (N_20824,N_19436,N_18518);
nor U20825 (N_20825,N_18341,N_18446);
nand U20826 (N_20826,N_17569,N_15710);
or U20827 (N_20827,N_15709,N_18457);
xnor U20828 (N_20828,N_17440,N_17947);
and U20829 (N_20829,N_18317,N_17606);
nor U20830 (N_20830,N_18066,N_17410);
and U20831 (N_20831,N_18255,N_19305);
and U20832 (N_20832,N_15335,N_15410);
nor U20833 (N_20833,N_19860,N_16157);
and U20834 (N_20834,N_19465,N_16186);
and U20835 (N_20835,N_19118,N_17075);
nor U20836 (N_20836,N_18692,N_17367);
nand U20837 (N_20837,N_17543,N_18366);
nor U20838 (N_20838,N_19548,N_17195);
nand U20839 (N_20839,N_16142,N_16416);
nand U20840 (N_20840,N_18220,N_15191);
and U20841 (N_20841,N_15281,N_16884);
nor U20842 (N_20842,N_15772,N_16914);
nand U20843 (N_20843,N_16510,N_18153);
nand U20844 (N_20844,N_18352,N_15855);
and U20845 (N_20845,N_17011,N_19456);
xor U20846 (N_20846,N_16476,N_18340);
nor U20847 (N_20847,N_17843,N_17711);
nand U20848 (N_20848,N_18244,N_15935);
and U20849 (N_20849,N_19614,N_17226);
nor U20850 (N_20850,N_19750,N_16271);
or U20851 (N_20851,N_19677,N_19670);
nand U20852 (N_20852,N_19973,N_15164);
or U20853 (N_20853,N_15803,N_15298);
nand U20854 (N_20854,N_17008,N_19464);
nor U20855 (N_20855,N_17902,N_18316);
nor U20856 (N_20856,N_18989,N_17849);
or U20857 (N_20857,N_19251,N_15583);
nor U20858 (N_20858,N_18633,N_18797);
nand U20859 (N_20859,N_17468,N_15911);
or U20860 (N_20860,N_15209,N_19613);
or U20861 (N_20861,N_16724,N_16631);
or U20862 (N_20862,N_17386,N_15702);
nand U20863 (N_20863,N_17465,N_16059);
nand U20864 (N_20864,N_15014,N_15838);
and U20865 (N_20865,N_15629,N_16087);
nand U20866 (N_20866,N_19008,N_19605);
and U20867 (N_20867,N_18110,N_19041);
nand U20868 (N_20868,N_18679,N_16138);
nor U20869 (N_20869,N_15764,N_19753);
xnor U20870 (N_20870,N_17505,N_15145);
nor U20871 (N_20871,N_19920,N_15770);
nor U20872 (N_20872,N_15153,N_15867);
xnor U20873 (N_20873,N_16336,N_18974);
nor U20874 (N_20874,N_17476,N_16616);
or U20875 (N_20875,N_16072,N_15851);
nand U20876 (N_20876,N_15171,N_16281);
nand U20877 (N_20877,N_15850,N_18361);
nor U20878 (N_20878,N_19050,N_16696);
nor U20879 (N_20879,N_15756,N_18742);
xor U20880 (N_20880,N_16425,N_16094);
and U20881 (N_20881,N_17561,N_16595);
nand U20882 (N_20882,N_18385,N_15561);
nor U20883 (N_20883,N_17936,N_19405);
xor U20884 (N_20884,N_18237,N_17922);
or U20885 (N_20885,N_15332,N_19244);
xor U20886 (N_20886,N_18866,N_16582);
nand U20887 (N_20887,N_15105,N_16015);
and U20888 (N_20888,N_17652,N_18780);
nand U20889 (N_20889,N_19952,N_18012);
or U20890 (N_20890,N_16318,N_19532);
or U20891 (N_20891,N_18449,N_17648);
xor U20892 (N_20892,N_16863,N_17965);
xnor U20893 (N_20893,N_18420,N_16784);
nand U20894 (N_20894,N_19644,N_17726);
nand U20895 (N_20895,N_18265,N_15352);
nor U20896 (N_20896,N_19667,N_18961);
or U20897 (N_20897,N_17324,N_17480);
nand U20898 (N_20898,N_17772,N_17522);
nand U20899 (N_20899,N_17908,N_19919);
xor U20900 (N_20900,N_18951,N_19620);
or U20901 (N_20901,N_17346,N_18297);
nor U20902 (N_20902,N_19705,N_17108);
nor U20903 (N_20903,N_17825,N_17891);
and U20904 (N_20904,N_18159,N_18545);
and U20905 (N_20905,N_19979,N_18779);
nor U20906 (N_20906,N_17484,N_15302);
nand U20907 (N_20907,N_15657,N_19941);
nand U20908 (N_20908,N_19767,N_19070);
nor U20909 (N_20909,N_15574,N_17706);
nand U20910 (N_20910,N_15057,N_16881);
xnor U20911 (N_20911,N_16633,N_15786);
nor U20912 (N_20912,N_19375,N_18097);
nand U20913 (N_20913,N_19577,N_15982);
xor U20914 (N_20914,N_18555,N_17542);
or U20915 (N_20915,N_17299,N_19347);
and U20916 (N_20916,N_18659,N_17326);
or U20917 (N_20917,N_19075,N_19187);
xnor U20918 (N_20918,N_17204,N_17730);
and U20919 (N_20919,N_19766,N_17305);
xor U20920 (N_20920,N_17676,N_17347);
nand U20921 (N_20921,N_17878,N_18435);
xor U20922 (N_20922,N_16677,N_15184);
or U20923 (N_20923,N_17228,N_17178);
nand U20924 (N_20924,N_19936,N_18183);
and U20925 (N_20925,N_17950,N_16290);
or U20926 (N_20926,N_17107,N_18023);
nand U20927 (N_20927,N_15062,N_16053);
xnor U20928 (N_20928,N_15810,N_15467);
xnor U20929 (N_20929,N_19852,N_17083);
xor U20930 (N_20930,N_15368,N_16572);
and U20931 (N_20931,N_16371,N_15592);
nand U20932 (N_20932,N_17132,N_15391);
xor U20933 (N_20933,N_18898,N_16162);
or U20934 (N_20934,N_19056,N_18765);
nor U20935 (N_20935,N_19891,N_19128);
and U20936 (N_20936,N_16368,N_19948);
and U20937 (N_20937,N_18999,N_16917);
nor U20938 (N_20938,N_17122,N_19821);
nor U20939 (N_20939,N_17738,N_17625);
and U20940 (N_20940,N_19349,N_15210);
nor U20941 (N_20941,N_17454,N_19438);
and U20942 (N_20942,N_17708,N_17123);
xor U20943 (N_20943,N_19596,N_15070);
or U20944 (N_20944,N_19518,N_17623);
and U20945 (N_20945,N_17193,N_16604);
xnor U20946 (N_20946,N_16443,N_17116);
or U20947 (N_20947,N_18320,N_17448);
nor U20948 (N_20948,N_16549,N_15972);
nor U20949 (N_20949,N_19454,N_16560);
and U20950 (N_20950,N_15789,N_19642);
and U20951 (N_20951,N_17836,N_17898);
and U20952 (N_20952,N_19630,N_15833);
xor U20953 (N_20953,N_16456,N_17851);
nand U20954 (N_20954,N_19309,N_16734);
and U20955 (N_20955,N_17660,N_18123);
nor U20956 (N_20956,N_18072,N_18940);
xnor U20957 (N_20957,N_15055,N_15061);
or U20958 (N_20958,N_18132,N_16858);
xnor U20959 (N_20959,N_16570,N_16518);
and U20960 (N_20960,N_18339,N_17776);
nand U20961 (N_20961,N_15658,N_18531);
nor U20962 (N_20962,N_19653,N_17402);
or U20963 (N_20963,N_17027,N_15757);
and U20964 (N_20964,N_19303,N_15328);
or U20965 (N_20965,N_17651,N_15964);
xor U20966 (N_20966,N_15476,N_18828);
xnor U20967 (N_20967,N_18920,N_15383);
and U20968 (N_20968,N_18693,N_15245);
xnor U20969 (N_20969,N_16946,N_18906);
and U20970 (N_20970,N_15914,N_17556);
nor U20971 (N_20971,N_18886,N_16990);
and U20972 (N_20972,N_16810,N_18651);
nand U20973 (N_20973,N_19048,N_15567);
nand U20974 (N_20974,N_16364,N_18370);
xor U20975 (N_20975,N_15708,N_16991);
xnor U20976 (N_20976,N_15790,N_19426);
xor U20977 (N_20977,N_17774,N_17952);
nor U20978 (N_20978,N_17626,N_15758);
nand U20979 (N_20979,N_17712,N_19392);
nor U20980 (N_20980,N_16689,N_19918);
or U20981 (N_20981,N_19017,N_18868);
nor U20982 (N_20982,N_19291,N_17180);
nor U20983 (N_20983,N_17236,N_19497);
nand U20984 (N_20984,N_16037,N_15762);
nor U20985 (N_20985,N_18411,N_18881);
nor U20986 (N_20986,N_16046,N_15044);
and U20987 (N_20987,N_18197,N_18282);
xor U20988 (N_20988,N_17187,N_15793);
nor U20989 (N_20989,N_15294,N_19219);
nor U20990 (N_20990,N_17688,N_17763);
nand U20991 (N_20991,N_19212,N_16066);
nand U20992 (N_20992,N_17885,N_18107);
nor U20993 (N_20993,N_17531,N_17446);
nand U20994 (N_20994,N_16835,N_18645);
xor U20995 (N_20995,N_18387,N_19627);
and U20996 (N_20996,N_19759,N_15846);
nand U20997 (N_20997,N_15267,N_16018);
nor U20998 (N_20998,N_16326,N_15727);
nand U20999 (N_20999,N_16463,N_17800);
xnor U21000 (N_21000,N_19415,N_16910);
or U21001 (N_21001,N_17232,N_17588);
nand U21002 (N_21002,N_17713,N_15395);
nand U21003 (N_21003,N_16732,N_17503);
or U21004 (N_21004,N_17580,N_17491);
or U21005 (N_21005,N_19372,N_16210);
nand U21006 (N_21006,N_15538,N_16418);
xor U21007 (N_21007,N_15142,N_17607);
and U21008 (N_21008,N_16070,N_18196);
nand U21009 (N_21009,N_18912,N_19966);
nor U21010 (N_21010,N_17250,N_17238);
or U21011 (N_21011,N_17627,N_19297);
nand U21012 (N_21012,N_16723,N_17413);
nand U21013 (N_21013,N_17234,N_16021);
nand U21014 (N_21014,N_19886,N_18939);
nand U21015 (N_21015,N_16718,N_17041);
nor U21016 (N_21016,N_17938,N_18914);
or U21017 (N_21017,N_16035,N_17257);
and U21018 (N_21018,N_18280,N_15182);
xnor U21019 (N_21019,N_17724,N_16052);
nand U21020 (N_21020,N_19059,N_15367);
nor U21021 (N_21021,N_15295,N_15378);
xnor U21022 (N_21022,N_19639,N_17789);
and U21023 (N_21023,N_15639,N_17373);
or U21024 (N_21024,N_18835,N_16446);
nand U21025 (N_21025,N_19393,N_19323);
and U21026 (N_21026,N_18344,N_16169);
xor U21027 (N_21027,N_17760,N_16630);
nor U21028 (N_21028,N_17042,N_18381);
and U21029 (N_21029,N_16324,N_15064);
xnor U21030 (N_21030,N_15865,N_15329);
nor U21031 (N_21031,N_19064,N_16349);
and U21032 (N_21032,N_16711,N_15318);
nor U21033 (N_21033,N_18490,N_18162);
nand U21034 (N_21034,N_17179,N_19999);
nor U21035 (N_21035,N_18179,N_17705);
nor U21036 (N_21036,N_17697,N_16113);
and U21037 (N_21037,N_16243,N_17665);
nor U21038 (N_21038,N_19529,N_17768);
and U21039 (N_21039,N_15151,N_15513);
and U21040 (N_21040,N_16622,N_18642);
nand U21041 (N_21041,N_16722,N_17006);
xnor U21042 (N_21042,N_16760,N_19198);
nor U21043 (N_21043,N_16012,N_16900);
and U21044 (N_21044,N_16264,N_18706);
or U21045 (N_21045,N_19130,N_19930);
xor U21046 (N_21046,N_19958,N_16212);
or U21047 (N_21047,N_15902,N_17121);
and U21048 (N_21048,N_18383,N_17174);
xor U21049 (N_21049,N_18111,N_18056);
nor U21050 (N_21050,N_15405,N_15380);
nand U21051 (N_21051,N_16752,N_18944);
and U21052 (N_21052,N_17394,N_18705);
xnor U21053 (N_21053,N_19479,N_19165);
xnor U21054 (N_21054,N_15776,N_18437);
xnor U21055 (N_21055,N_15194,N_18295);
xnor U21056 (N_21056,N_18402,N_18824);
and U21057 (N_21057,N_18028,N_17271);
or U21058 (N_21058,N_18369,N_18062);
nand U21059 (N_21059,N_15141,N_15104);
or U21060 (N_21060,N_16322,N_19861);
nor U21061 (N_21061,N_18763,N_19910);
nor U21062 (N_21062,N_19265,N_16886);
nor U21063 (N_21063,N_17316,N_15479);
xnor U21064 (N_21064,N_16823,N_15478);
xor U21065 (N_21065,N_18915,N_17090);
xor U21066 (N_21066,N_16547,N_19006);
and U21067 (N_21067,N_16105,N_15088);
and U21068 (N_21068,N_19081,N_19109);
nand U21069 (N_21069,N_17863,N_16078);
or U21070 (N_21070,N_17761,N_17502);
and U21071 (N_21071,N_17537,N_19329);
nand U21072 (N_21072,N_19121,N_15706);
nor U21073 (N_21073,N_16908,N_17528);
xor U21074 (N_21074,N_15950,N_16039);
nor U21075 (N_21075,N_19905,N_18212);
or U21076 (N_21076,N_18843,N_16362);
nand U21077 (N_21077,N_17086,N_19073);
or U21078 (N_21078,N_15272,N_17608);
nor U21079 (N_21079,N_18833,N_18442);
and U21080 (N_21080,N_17837,N_16214);
nand U21081 (N_21081,N_17803,N_15811);
or U21082 (N_21082,N_18950,N_15446);
xor U21083 (N_21083,N_19885,N_15238);
or U21084 (N_21084,N_16375,N_15021);
xor U21085 (N_21085,N_17339,N_16381);
nand U21086 (N_21086,N_16455,N_18063);
xor U21087 (N_21087,N_16599,N_17970);
xnor U21088 (N_21088,N_17988,N_15110);
and U21089 (N_21089,N_19377,N_19880);
nor U21090 (N_21090,N_16516,N_17374);
xor U21091 (N_21091,N_17296,N_15976);
xor U21092 (N_21092,N_16435,N_19698);
nand U21093 (N_21093,N_16027,N_16155);
and U21094 (N_21094,N_17817,N_15832);
or U21095 (N_21095,N_16873,N_15228);
nand U21096 (N_21096,N_16496,N_19754);
or U21097 (N_21097,N_19770,N_16065);
nor U21098 (N_21098,N_15510,N_16821);
or U21099 (N_21099,N_19574,N_15308);
or U21100 (N_21100,N_18334,N_15456);
nor U21101 (N_21101,N_17696,N_18445);
and U21102 (N_21102,N_19170,N_19546);
xor U21103 (N_21103,N_19597,N_18860);
nor U21104 (N_21104,N_18338,N_17716);
and U21105 (N_21105,N_15152,N_17420);
xor U21106 (N_21106,N_19264,N_15206);
and U21107 (N_21107,N_15170,N_19862);
and U21108 (N_21108,N_18800,N_18289);
xor U21109 (N_21109,N_16268,N_18899);
xnor U21110 (N_21110,N_16500,N_17247);
and U21111 (N_21111,N_16096,N_19299);
nor U21112 (N_21112,N_17210,N_17872);
nand U21113 (N_21113,N_19026,N_17213);
nand U21114 (N_21114,N_19132,N_19512);
xor U21115 (N_21115,N_18676,N_15327);
and U21116 (N_21116,N_16265,N_16674);
xnor U21117 (N_21117,N_19678,N_17923);
xor U21118 (N_21118,N_18488,N_18734);
xor U21119 (N_21119,N_19344,N_16623);
or U21120 (N_21120,N_15394,N_19182);
or U21121 (N_21121,N_16398,N_19586);
nand U21122 (N_21122,N_15423,N_17826);
or U21123 (N_21123,N_18702,N_16047);
nand U21124 (N_21124,N_17212,N_18787);
nand U21125 (N_21125,N_18118,N_15566);
xor U21126 (N_21126,N_17001,N_17714);
and U21127 (N_21127,N_17672,N_17419);
xnor U21128 (N_21128,N_17242,N_16003);
nand U21129 (N_21129,N_18678,N_15270);
and U21130 (N_21130,N_17500,N_16625);
and U21131 (N_21131,N_18752,N_15951);
nand U21132 (N_21132,N_19940,N_17079);
nor U21133 (N_21133,N_17842,N_18713);
nand U21134 (N_21134,N_15284,N_17934);
and U21135 (N_21135,N_16799,N_19960);
nor U21136 (N_21136,N_17956,N_17382);
nand U21137 (N_21137,N_15553,N_19506);
and U21138 (N_21138,N_18239,N_16829);
or U21139 (N_21139,N_18686,N_15146);
xnor U21140 (N_21140,N_16453,N_15366);
or U21141 (N_21141,N_19661,N_17377);
and U21142 (N_21142,N_16370,N_18557);
nand U21143 (N_21143,N_16628,N_18586);
nand U21144 (N_21144,N_17013,N_15488);
nor U21145 (N_21145,N_18976,N_18102);
nor U21146 (N_21146,N_15536,N_18479);
nor U21147 (N_21147,N_19707,N_19713);
nand U21148 (N_21148,N_18142,N_18701);
nor U21149 (N_21149,N_17134,N_17643);
nand U21150 (N_21150,N_16298,N_16352);
xor U21151 (N_21151,N_18815,N_18263);
and U21152 (N_21152,N_15504,N_17946);
and U21153 (N_21153,N_17838,N_18670);
and U21154 (N_21154,N_18356,N_16235);
or U21155 (N_21155,N_16838,N_16720);
and U21156 (N_21156,N_15897,N_19963);
or U21157 (N_21157,N_15848,N_19870);
or U21158 (N_21158,N_16998,N_17539);
nor U21159 (N_21159,N_15432,N_19346);
and U21160 (N_21160,N_17735,N_15805);
nor U21161 (N_21161,N_15520,N_19382);
and U21162 (N_21162,N_18731,N_18822);
xnor U21163 (N_21163,N_19841,N_19236);
and U21164 (N_21164,N_16331,N_15382);
xnor U21165 (N_21165,N_18026,N_17883);
and U21166 (N_21166,N_18202,N_18172);
nor U21167 (N_21167,N_17057,N_15747);
and U21168 (N_21168,N_17159,N_19545);
and U21169 (N_21169,N_15012,N_19715);
and U21170 (N_21170,N_15255,N_17475);
xor U21171 (N_21171,N_15782,N_19100);
nand U21172 (N_21172,N_19562,N_18694);
nand U21173 (N_21173,N_17527,N_19712);
xor U21174 (N_21174,N_18819,N_18838);
nand U21175 (N_21175,N_16957,N_16199);
nand U21176 (N_21176,N_19274,N_18988);
nand U21177 (N_21177,N_17091,N_18277);
nor U21178 (N_21178,N_17219,N_19311);
and U21179 (N_21179,N_17051,N_16989);
xnor U21180 (N_21180,N_19028,N_16524);
or U21181 (N_21181,N_17613,N_18409);
xor U21182 (N_21182,N_18461,N_18081);
nor U21183 (N_21183,N_19091,N_18526);
nand U21184 (N_21184,N_19381,N_15234);
or U21185 (N_21185,N_15339,N_17102);
xor U21186 (N_21186,N_17515,N_15037);
xor U21187 (N_21187,N_16427,N_18851);
nand U21188 (N_21188,N_18058,N_17127);
or U21189 (N_21189,N_16079,N_15515);
xnor U21190 (N_21190,N_16354,N_18455);
or U21191 (N_21191,N_15490,N_16935);
nor U21192 (N_21192,N_19066,N_19933);
nand U21193 (N_21193,N_16794,N_17251);
and U21194 (N_21194,N_19084,N_18022);
nand U21195 (N_21195,N_17674,N_15195);
xnor U21196 (N_21196,N_15392,N_19890);
and U21197 (N_21197,N_18661,N_15671);
and U21198 (N_21198,N_16311,N_18161);
xnor U21199 (N_21199,N_18773,N_19239);
nand U21200 (N_21200,N_18911,N_15735);
and U21201 (N_21201,N_16553,N_17565);
nor U21202 (N_21202,N_16952,N_16002);
xnor U21203 (N_21203,N_18404,N_19137);
or U21204 (N_21204,N_16135,N_18565);
nand U21205 (N_21205,N_18749,N_19740);
nand U21206 (N_21206,N_19938,N_15826);
xor U21207 (N_21207,N_19656,N_18964);
and U21208 (N_21208,N_17131,N_16975);
or U21209 (N_21209,N_17892,N_16167);
and U21210 (N_21210,N_18348,N_17363);
xor U21211 (N_21211,N_15365,N_19412);
xor U21212 (N_21212,N_18372,N_17183);
xor U21213 (N_21213,N_17231,N_19977);
nor U21214 (N_21214,N_17554,N_16610);
xor U21215 (N_21215,N_19430,N_19764);
nand U21216 (N_21216,N_19691,N_17985);
nor U21217 (N_21217,N_15176,N_16494);
nor U21218 (N_21218,N_15472,N_18623);
or U21219 (N_21219,N_16068,N_19354);
xnor U21220 (N_21220,N_17430,N_16626);
and U21221 (N_21221,N_19625,N_17270);
nand U21222 (N_21222,N_19509,N_19955);
or U21223 (N_21223,N_17963,N_18875);
xnor U21224 (N_21224,N_19158,N_19517);
nor U21225 (N_21225,N_19560,N_16179);
xnor U21226 (N_21226,N_19917,N_18222);
nor U21227 (N_21227,N_18580,N_16426);
nor U21228 (N_21228,N_15369,N_15502);
xnor U21229 (N_21229,N_16306,N_15957);
xor U21230 (N_21230,N_17488,N_15447);
nand U21231 (N_21231,N_18821,N_16014);
xnor U21232 (N_21232,N_19716,N_18147);
nor U21233 (N_21233,N_17644,N_18923);
nor U21234 (N_21234,N_15720,N_17171);
nor U21235 (N_21235,N_16197,N_16006);
and U21236 (N_21236,N_16819,N_15634);
and U21237 (N_21237,N_16444,N_17147);
nand U21238 (N_21238,N_18144,N_17557);
xor U21239 (N_21239,N_17990,N_18504);
xnor U21240 (N_21240,N_16288,N_15900);
and U21241 (N_21241,N_16254,N_18399);
xnor U21242 (N_21242,N_17245,N_18379);
and U21243 (N_21243,N_15990,N_17791);
and U21244 (N_21244,N_15873,N_15158);
nor U21245 (N_21245,N_19045,N_16259);
and U21246 (N_21246,N_15185,N_18182);
nand U21247 (N_21247,N_15890,N_15906);
xor U21248 (N_21248,N_17524,N_18252);
xor U21249 (N_21249,N_16029,N_15963);
nor U21250 (N_21250,N_15051,N_18160);
nor U21251 (N_21251,N_19123,N_17105);
nor U21252 (N_21252,N_16943,N_16993);
or U21253 (N_21253,N_19601,N_19060);
xor U21254 (N_21254,N_15841,N_17808);
xnor U21255 (N_21255,N_16543,N_15967);
nand U21256 (N_21256,N_17277,N_17112);
nand U21257 (N_21257,N_15560,N_17822);
nor U21258 (N_21258,N_15388,N_18578);
xnor U21259 (N_21259,N_17869,N_18804);
nor U21260 (N_21260,N_16401,N_18684);
nor U21261 (N_21261,N_19662,N_17861);
or U21262 (N_21262,N_19869,N_17832);
and U21263 (N_21263,N_17656,N_18949);
xnor U21264 (N_21264,N_18464,N_19925);
or U21265 (N_21265,N_15692,N_16410);
nor U21266 (N_21266,N_16565,N_15148);
and U21267 (N_21267,N_17621,N_18013);
or U21268 (N_21268,N_18002,N_16883);
nand U21269 (N_21269,N_16954,N_17050);
and U21270 (N_21270,N_16487,N_19071);
or U21271 (N_21271,N_18577,N_17589);
xor U21272 (N_21272,N_17026,N_18631);
and U21273 (N_21273,N_19665,N_19475);
nand U21274 (N_21274,N_15087,N_17356);
xor U21275 (N_21275,N_19489,N_19049);
nor U21276 (N_21276,N_16640,N_16887);
nand U21277 (N_21277,N_15320,N_15296);
nor U21278 (N_21278,N_19083,N_15083);
and U21279 (N_21279,N_19227,N_19813);
nand U21280 (N_21280,N_17146,N_17717);
and U21281 (N_21281,N_15261,N_17370);
nand U21282 (N_21282,N_19463,N_18737);
xnor U21283 (N_21283,N_18726,N_15440);
nor U21284 (N_21284,N_18331,N_15779);
xor U21285 (N_21285,N_18079,N_15674);
and U21286 (N_21286,N_19111,N_18139);
nor U21287 (N_21287,N_17504,N_19398);
nand U21288 (N_21288,N_16617,N_15279);
nor U21289 (N_21289,N_19246,N_19477);
nand U21290 (N_21290,N_17021,N_19390);
xnor U21291 (N_21291,N_17897,N_19638);
or U21292 (N_21292,N_17106,N_18652);
xor U21293 (N_21293,N_17432,N_19674);
or U21294 (N_21294,N_16061,N_15094);
nand U21295 (N_21295,N_15031,N_17743);
or U21296 (N_21296,N_16520,N_16865);
nor U21297 (N_21297,N_15787,N_15630);
or U21298 (N_21298,N_17267,N_19559);
nor U21299 (N_21299,N_15862,N_19307);
nand U21300 (N_21300,N_15965,N_17492);
xor U21301 (N_21301,N_16860,N_18650);
nand U21302 (N_21302,N_15598,N_16895);
nand U21303 (N_21303,N_18969,N_19326);
nor U21304 (N_21304,N_18755,N_16751);
nor U21305 (N_21305,N_17845,N_17076);
nand U21306 (N_21306,N_15936,N_18093);
xnor U21307 (N_21307,N_19413,N_17364);
or U21308 (N_21308,N_18879,N_16471);
nand U21309 (N_21309,N_15644,N_16428);
nor U21310 (N_21310,N_19552,N_18459);
and U21311 (N_21311,N_16762,N_19826);
and U21312 (N_21312,N_16465,N_19220);
and U21313 (N_21313,N_16988,N_17306);
xnor U21314 (N_21314,N_15667,N_15427);
and U21315 (N_21315,N_19112,N_19655);
and U21316 (N_21316,N_19991,N_18739);
xor U21317 (N_21317,N_15527,N_18632);
nand U21318 (N_21318,N_17331,N_17162);
xnor U21319 (N_21319,N_18408,N_19424);
nand U21320 (N_21320,N_15703,N_19777);
and U21321 (N_21321,N_18516,N_17053);
nand U21322 (N_21322,N_17062,N_18660);
and U21323 (N_21323,N_19557,N_16041);
nor U21324 (N_21324,N_19641,N_16728);
and U21325 (N_21325,N_17905,N_15487);
or U21326 (N_21326,N_18931,N_18152);
nand U21327 (N_21327,N_18809,N_15874);
and U21328 (N_21328,N_16792,N_15484);
or U21329 (N_21329,N_17140,N_19598);
nor U21330 (N_21330,N_15662,N_15670);
and U21331 (N_21331,N_19419,N_18500);
xor U21332 (N_21332,N_19062,N_17343);
nor U21333 (N_21333,N_17322,N_18572);
or U21334 (N_21334,N_18547,N_17319);
or U21335 (N_21335,N_16837,N_17875);
nor U21336 (N_21336,N_19404,N_16682);
and U21337 (N_21337,N_16327,N_19300);
xor U21338 (N_21338,N_15587,N_19476);
nor U21339 (N_21339,N_18354,N_15697);
nand U21340 (N_21340,N_18745,N_15093);
nand U21341 (N_21341,N_18688,N_18210);
and U21342 (N_21342,N_15823,N_15690);
or U21343 (N_21343,N_18643,N_15197);
nor U21344 (N_21344,N_19987,N_15398);
nand U21345 (N_21345,N_17291,N_19928);
xnor U21346 (N_21346,N_18893,N_16278);
xnor U21347 (N_21347,N_19554,N_18475);
and U21348 (N_21348,N_17287,N_16870);
xor U21349 (N_21349,N_17223,N_18626);
and U21350 (N_21350,N_19423,N_15611);
nor U21351 (N_21351,N_16232,N_16596);
and U21352 (N_21352,N_17691,N_16329);
nand U21353 (N_21353,N_17208,N_17928);
xnor U21354 (N_21354,N_18048,N_18979);
nor U21355 (N_21355,N_17961,N_17046);
xnor U21356 (N_21356,N_17252,N_18603);
and U21357 (N_21357,N_15123,N_18456);
and U21358 (N_21358,N_16985,N_17816);
nand U21359 (N_21359,N_19431,N_16962);
or U21360 (N_21360,N_15248,N_19492);
and U21361 (N_21361,N_15818,N_15174);
or U21362 (N_21362,N_16527,N_15827);
nor U21363 (N_21363,N_16542,N_15750);
nand U21364 (N_21364,N_16747,N_15830);
nor U21365 (N_21365,N_18867,N_16396);
or U21366 (N_21366,N_16168,N_18535);
nand U21367 (N_21367,N_16160,N_15771);
nand U21368 (N_21368,N_18214,N_18407);
nand U21369 (N_21369,N_16161,N_19658);
nand U21370 (N_21370,N_18443,N_17074);
nor U21371 (N_21371,N_17721,N_15548);
xnor U21372 (N_21372,N_18826,N_15937);
xnor U21373 (N_21373,N_15125,N_17431);
nand U21374 (N_21374,N_16933,N_19216);
nor U21375 (N_21375,N_17478,N_18847);
or U21376 (N_21376,N_16299,N_15168);
and U21377 (N_21377,N_16108,N_19582);
xnor U21378 (N_21378,N_18658,N_18248);
or U21379 (N_21379,N_17466,N_19457);
nand U21380 (N_21380,N_17748,N_19942);
or U21381 (N_21381,N_17728,N_18225);
nand U21382 (N_21382,N_19356,N_18859);
or U21383 (N_21383,N_19455,N_17350);
xor U21384 (N_21384,N_17657,N_17572);
nand U21385 (N_21385,N_17518,N_17285);
nor U21386 (N_21386,N_18345,N_18935);
or U21387 (N_21387,N_19482,N_18273);
nor U21388 (N_21388,N_17918,N_17209);
or U21389 (N_21389,N_16420,N_15480);
nand U21390 (N_21390,N_17470,N_15474);
or U21391 (N_21391,N_17686,N_15111);
nor U21392 (N_21392,N_18744,N_18261);
or U21393 (N_21393,N_15041,N_15040);
nand U21394 (N_21394,N_19643,N_16738);
and U21395 (N_21395,N_17989,N_15032);
nand U21396 (N_21396,N_19117,N_18441);
and U21397 (N_21397,N_15232,N_18077);
nand U21398 (N_21398,N_17284,N_18901);
or U21399 (N_21399,N_19253,N_19751);
and U21400 (N_21400,N_18928,N_16083);
nor U21401 (N_21401,N_17741,N_18857);
xor U21402 (N_21402,N_16713,N_17064);
nor U21403 (N_21403,N_16568,N_18105);
nor U21404 (N_21404,N_15230,N_15165);
and U21405 (N_21405,N_15473,N_16077);
xor U21406 (N_21406,N_16802,N_18965);
xor U21407 (N_21407,N_18597,N_16805);
or U21408 (N_21408,N_16253,N_16798);
and U21409 (N_21409,N_17590,N_18913);
or U21410 (N_21410,N_15147,N_15523);
xnor U21411 (N_21411,N_19503,N_19504);
nand U21412 (N_21412,N_18722,N_19005);
and U21413 (N_21413,N_16369,N_15043);
or U21414 (N_21414,N_16207,N_18883);
nor U21415 (N_21415,N_19142,N_17578);
and U21416 (N_21416,N_18538,N_15575);
nor U21417 (N_21417,N_16196,N_19119);
or U21418 (N_21418,N_18243,N_18363);
or U21419 (N_21419,N_16434,N_17283);
nand U21420 (N_21420,N_16228,N_15416);
or U21421 (N_21421,N_17389,N_17485);
nor U21422 (N_21422,N_19801,N_18808);
or U21423 (N_21423,N_15342,N_19434);
xor U21424 (N_21424,N_19547,N_18069);
nand U21425 (N_21425,N_18021,N_17551);
xor U21426 (N_21426,N_18481,N_16770);
or U21427 (N_21427,N_18397,N_15241);
nand U21428 (N_21428,N_19133,N_19722);
or U21429 (N_21429,N_16472,N_16847);
nor U21430 (N_21430,N_16383,N_19539);
xor U21431 (N_21431,N_15748,N_15797);
xor U21432 (N_21432,N_16948,N_17490);
and U21433 (N_21433,N_16220,N_15212);
xor U21434 (N_21434,N_19422,N_17221);
xnor U21435 (N_21435,N_18235,N_18612);
nand U21436 (N_21436,N_15571,N_15390);
nand U21437 (N_21437,N_19126,N_16663);
nand U21438 (N_21438,N_18390,N_19139);
nor U21439 (N_21439,N_16499,N_16573);
nand U21440 (N_21440,N_15399,N_16378);
or U21441 (N_21441,N_15271,N_15060);
or U21442 (N_21442,N_15301,N_15355);
or U21443 (N_21443,N_18596,N_18073);
nor U21444 (N_21444,N_17907,N_18510);
nand U21445 (N_21445,N_18973,N_17254);
or U21446 (N_21446,N_17114,N_16092);
xnor U21447 (N_21447,N_18482,N_18724);
xor U21448 (N_21448,N_16181,N_17428);
and U21449 (N_21449,N_16182,N_15307);
nor U21450 (N_21450,N_19949,N_19533);
xor U21451 (N_21451,N_16922,N_16402);
nand U21452 (N_21452,N_18067,N_19535);
xor U21453 (N_21453,N_18522,N_16468);
xnor U21454 (N_21454,N_19458,N_17511);
nor U21455 (N_21455,N_17422,N_15604);
nor U21456 (N_21456,N_15947,N_16567);
nand U21457 (N_21457,N_19389,N_18907);
and U21458 (N_21458,N_15095,N_18957);
nand U21459 (N_21459,N_19902,N_15221);
and U21460 (N_21460,N_18870,N_18646);
and U21461 (N_21461,N_15529,N_17835);
nor U21462 (N_21462,N_17028,N_15552);
or U21463 (N_21463,N_15264,N_15054);
nand U21464 (N_21464,N_19169,N_18521);
xnor U21465 (N_21465,N_15955,N_19974);
xnor U21466 (N_21466,N_15909,N_16961);
and U21467 (N_21467,N_18848,N_16279);
or U21468 (N_21468,N_17833,N_17233);
and U21469 (N_21469,N_19429,N_15678);
and U21470 (N_21470,N_16171,N_18125);
nand U21471 (N_21471,N_19207,N_18452);
nand U21472 (N_21472,N_16448,N_15683);
and U21473 (N_21473,N_17462,N_17942);
xnor U21474 (N_21474,N_19258,N_18494);
xor U21475 (N_21475,N_17018,N_18649);
nand U21476 (N_21476,N_18219,N_15694);
and U21477 (N_21477,N_16519,N_15888);
xor U21478 (N_21478,N_17297,N_16452);
nand U21479 (N_21479,N_18314,N_19995);
nor U21480 (N_21480,N_15357,N_16050);
nand U21481 (N_21481,N_19320,N_18608);
nand U21482 (N_21482,N_15791,N_18465);
xnor U21483 (N_21483,N_18788,N_15988);
and U21484 (N_21484,N_18008,N_16761);
nand U21485 (N_21485,N_16634,N_15871);
and U21486 (N_21486,N_15618,N_19632);
nand U21487 (N_21487,N_18284,N_18882);
nor U21488 (N_21488,N_19115,N_18941);
and U21489 (N_21489,N_18892,N_15765);
nor U21490 (N_21490,N_17070,N_17635);
nor U21491 (N_21491,N_15607,N_16869);
or U21492 (N_21492,N_15712,N_15923);
xor U21493 (N_21493,N_18451,N_18863);
and U21494 (N_21494,N_16304,N_19018);
nand U21495 (N_21495,N_16256,N_15675);
nor U21496 (N_21496,N_19292,N_16315);
xor U21497 (N_21497,N_19104,N_16344);
nor U21498 (N_21498,N_19148,N_15091);
and U21499 (N_21499,N_19052,N_19723);
or U21500 (N_21500,N_19054,N_15224);
nand U21501 (N_21501,N_17785,N_19331);
or U21502 (N_21502,N_15780,N_15072);
and U21503 (N_21503,N_16931,N_16049);
or U21504 (N_21504,N_16208,N_16697);
nor U21505 (N_21505,N_19748,N_15864);
or U21506 (N_21506,N_16234,N_18257);
nor U21507 (N_21507,N_17700,N_17483);
nor U21508 (N_21508,N_19397,N_15880);
nor U21509 (N_21509,N_19745,N_17514);
nand U21510 (N_21510,N_17009,N_16831);
or U21511 (N_21511,N_18885,N_17259);
nand U21512 (N_21512,N_19069,N_17831);
and U21513 (N_21513,N_18581,N_15024);
or U21514 (N_21514,N_19646,N_18151);
xor U21515 (N_21515,N_15745,N_19351);
xnor U21516 (N_21516,N_16530,N_17031);
nor U21517 (N_21517,N_17901,N_17732);
and U21518 (N_21518,N_16548,N_17467);
nand U21519 (N_21519,N_17740,N_18874);
nand U21520 (N_21520,N_19531,N_18946);
and U21521 (N_21521,N_17624,N_18924);
xnor U21522 (N_21522,N_18268,N_15570);
or U21523 (N_21523,N_19773,N_18758);
xor U21524 (N_21524,N_19592,N_15236);
and U21525 (N_21525,N_16482,N_17616);
and U21526 (N_21526,N_15045,N_15956);
nand U21527 (N_21527,N_15999,N_16363);
or U21528 (N_21528,N_16319,N_17639);
nand U21529 (N_21529,N_18837,N_18146);
nor U21530 (N_21530,N_16166,N_19866);
or U21531 (N_21531,N_19221,N_19849);
and U21532 (N_21532,N_16642,N_18897);
xor U21533 (N_21533,N_18968,N_15106);
nor U21534 (N_21534,N_18186,N_19953);
and U21535 (N_21535,N_17992,N_17274);
nand U21536 (N_21536,N_17166,N_18869);
nand U21537 (N_21537,N_16601,N_18425);
nor U21538 (N_21538,N_17559,N_19486);
xor U21539 (N_21539,N_17200,N_16307);
and U21540 (N_21540,N_18938,N_15379);
nand U21541 (N_21541,N_17224,N_15879);
xnor U21542 (N_21542,N_15813,N_18542);
or U21543 (N_21543,N_15262,N_17381);
nor U21544 (N_21544,N_16968,N_18663);
and U21545 (N_21545,N_18349,N_15364);
or U21546 (N_21546,N_15954,N_19516);
xor U21547 (N_21547,N_17125,N_15595);
or U21548 (N_21548,N_16249,N_19944);
or U21549 (N_21549,N_18430,N_15330);
or U21550 (N_21550,N_18088,N_15150);
or U21551 (N_21551,N_16438,N_17737);
nor U21552 (N_21552,N_19124,N_16408);
nand U21553 (N_21553,N_17392,N_18630);
nor U21554 (N_21554,N_19524,N_15321);
nand U21555 (N_21555,N_19270,N_16719);
nor U21556 (N_21556,N_15834,N_17920);
and U21557 (N_21557,N_17160,N_19881);
xor U21558 (N_21558,N_15180,N_17054);
or U21559 (N_21559,N_16716,N_19752);
and U21560 (N_21560,N_17583,N_19672);
nor U21561 (N_21561,N_19782,N_18174);
or U21562 (N_21562,N_18311,N_15980);
or U21563 (N_21563,N_17600,N_17562);
nor U21564 (N_21564,N_18365,N_19074);
and U21565 (N_21565,N_17844,N_17205);
or U21566 (N_21566,N_19391,N_15438);
and U21567 (N_21567,N_17820,N_17679);
nor U21568 (N_21568,N_16183,N_19166);
nor U21569 (N_21569,N_16102,N_19924);
and U21570 (N_21570,N_16574,N_19092);
or U21571 (N_21571,N_16397,N_16377);
nand U21572 (N_21572,N_16051,N_19285);
nand U21573 (N_21573,N_18323,N_19811);
and U21574 (N_21574,N_15576,N_19758);
nor U21575 (N_21575,N_18995,N_15116);
and U21576 (N_21576,N_15323,N_16781);
or U21577 (N_21577,N_16921,N_18551);
xnor U21578 (N_21578,N_15852,N_19093);
and U21579 (N_21579,N_16134,N_15534);
nand U21580 (N_21580,N_18228,N_19945);
and U21581 (N_21581,N_19799,N_16657);
nor U21582 (N_21582,N_19339,N_15025);
xor U21583 (N_21583,N_17575,N_17315);
and U21584 (N_21584,N_19085,N_19068);
and U21585 (N_21585,N_15562,N_19624);
nor U21586 (N_21586,N_18209,N_19626);
and U21587 (N_21587,N_18853,N_19848);
and U21588 (N_21588,N_18415,N_17780);
and U21589 (N_21589,N_19313,N_19828);
nor U21590 (N_21590,N_15718,N_18840);
nand U21591 (N_21591,N_17994,N_15783);
and U21592 (N_21592,N_19490,N_18918);
xor U21593 (N_21593,N_17302,N_18570);
and U21594 (N_21594,N_15053,N_19366);
and U21595 (N_21595,N_16844,N_16953);
xor U21596 (N_21596,N_18607,N_18226);
xor U21597 (N_21597,N_16074,N_18343);
or U21598 (N_21598,N_16672,N_15222);
or U21599 (N_21599,N_17384,N_19916);
or U21600 (N_21600,N_18592,N_18380);
or U21601 (N_21601,N_16766,N_19281);
nand U21602 (N_21602,N_19272,N_18635);
or U21603 (N_21603,N_19044,N_16038);
and U21604 (N_21604,N_19733,N_18970);
or U21605 (N_21605,N_19035,N_15420);
and U21606 (N_21606,N_15461,N_18640);
nor U21607 (N_21607,N_17099,N_17487);
nor U21608 (N_21608,N_19057,N_16414);
and U21609 (N_21609,N_15761,N_17477);
nor U21610 (N_21610,N_19021,N_16060);
nor U21611 (N_21611,N_15437,N_18743);
xnor U21612 (N_21612,N_19680,N_15896);
and U21613 (N_21613,N_17806,N_18143);
xnor U21614 (N_21614,N_19293,N_19131);
nor U21615 (N_21615,N_16112,N_17142);
nor U21616 (N_21616,N_15101,N_17169);
and U21617 (N_21617,N_19794,N_16843);
xnor U21618 (N_21618,N_18367,N_16305);
and U21619 (N_21619,N_18594,N_17501);
nand U21620 (N_21620,N_17002,N_16376);
or U21621 (N_21621,N_17982,N_16645);
nand U21622 (N_21622,N_15622,N_19322);
nand U21623 (N_21623,N_18127,N_15863);
or U21624 (N_21624,N_15445,N_17680);
and U21625 (N_21625,N_17612,N_19214);
nand U21626 (N_21626,N_19156,N_17882);
xor U21627 (N_21627,N_19287,N_15079);
xor U21628 (N_21628,N_15217,N_18776);
nand U21629 (N_21629,N_19485,N_16566);
xnor U21630 (N_21630,N_16450,N_19192);
xor U21631 (N_21631,N_19184,N_16439);
and U21632 (N_21632,N_19257,N_18673);
and U21633 (N_21633,N_15163,N_17298);
nand U21634 (N_21634,N_17295,N_15739);
xnor U21635 (N_21635,N_16862,N_18515);
or U21636 (N_21636,N_17423,N_17586);
xor U21637 (N_21637,N_18042,N_16123);
xnor U21638 (N_21638,N_16955,N_15903);
or U21639 (N_21639,N_18672,N_17729);
and U21640 (N_21640,N_16684,N_19097);
and U21641 (N_21641,N_19190,N_17827);
xor U21642 (N_21642,N_18794,N_15625);
xnor U21643 (N_21643,N_18053,N_19623);
or U21644 (N_21644,N_16648,N_18150);
or U21645 (N_21645,N_16959,N_17455);
and U21646 (N_21646,N_19755,N_17784);
or U21647 (N_21647,N_17493,N_17647);
nor U21648 (N_21648,N_19134,N_18813);
nor U21649 (N_21649,N_15119,N_16924);
nand U21650 (N_21650,N_17025,N_15542);
nor U21651 (N_21651,N_18728,N_17362);
nand U21652 (N_21652,N_16758,N_19523);
nand U21653 (N_21653,N_17268,N_19315);
nor U21654 (N_21654,N_17087,N_18328);
nor U21655 (N_21655,N_19634,N_16323);
and U21656 (N_21656,N_19829,N_15878);
or U21657 (N_21657,N_18984,N_16994);
nand U21658 (N_21658,N_15268,N_19802);
xnor U21659 (N_21659,N_19825,N_19686);
or U21660 (N_21660,N_19283,N_15578);
and U21661 (N_21661,N_16587,N_18820);
nor U21662 (N_21662,N_15828,N_16423);
xnor U21663 (N_21663,N_16174,N_19345);
nand U21664 (N_21664,N_15129,N_19566);
or U21665 (N_21665,N_17573,N_15656);
nand U21666 (N_21666,N_18207,N_19420);
or U21667 (N_21667,N_19950,N_17669);
nor U21668 (N_21668,N_17661,N_19141);
or U21669 (N_21669,N_17148,N_17576);
or U21670 (N_21670,N_15573,N_18377);
xnor U21671 (N_21671,N_16091,N_17264);
nor U21672 (N_21672,N_19153,N_17395);
and U21673 (N_21673,N_15815,N_18655);
xnor U21674 (N_21674,N_16911,N_18413);
nor U21675 (N_21675,N_18785,N_19282);
xor U21676 (N_21676,N_15569,N_19078);
xnor U21677 (N_21677,N_15631,N_16007);
or U21678 (N_21678,N_18458,N_17853);
or U21679 (N_21679,N_19685,N_16504);
or U21680 (N_21680,N_16111,N_15601);
or U21681 (N_21681,N_18453,N_19844);
or U21682 (N_21682,N_18865,N_18117);
nor U21683 (N_21683,N_17077,N_18786);
and U21684 (N_21684,N_15555,N_16193);
and U21685 (N_21685,N_17218,N_16273);
or U21686 (N_21686,N_19591,N_18948);
nand U21687 (N_21687,N_19823,N_18141);
nor U21688 (N_21688,N_18134,N_17879);
or U21689 (N_21689,N_15987,N_19868);
xor U21690 (N_21690,N_19294,N_15844);
xor U21691 (N_21691,N_19679,N_15736);
and U21692 (N_21692,N_17538,N_19934);
xor U21693 (N_21693,N_17022,N_18038);
nor U21694 (N_21694,N_19334,N_16700);
or U21695 (N_21695,N_16685,N_15500);
xor U21696 (N_21696,N_17032,N_17498);
or U21697 (N_21697,N_17126,N_18844);
and U21698 (N_21698,N_17884,N_19687);
xnor U21699 (N_21699,N_15448,N_18582);
or U21700 (N_21700,N_16137,N_19654);
and U21701 (N_21701,N_19202,N_17848);
nor U21702 (N_21702,N_19180,N_19400);
nor U21703 (N_21703,N_15269,N_16356);
nand U21704 (N_21704,N_19892,N_17019);
xor U21705 (N_21705,N_15544,N_17778);
or U21706 (N_21706,N_18283,N_16449);
and U21707 (N_21707,N_16650,N_16389);
nor U21708 (N_21708,N_19696,N_18595);
nor U21709 (N_21709,N_18114,N_19846);
nand U21710 (N_21710,N_18523,N_19728);
and U21711 (N_21711,N_17904,N_16280);
xnor U21712 (N_21712,N_18799,N_17095);
xor U21713 (N_21713,N_16864,N_18497);
and U21714 (N_21714,N_19493,N_18707);
and U21715 (N_21715,N_16788,N_19033);
and U21716 (N_21716,N_16085,N_16840);
nor U21717 (N_21717,N_18544,N_16671);
nor U21718 (N_21718,N_16977,N_18732);
and U21719 (N_21719,N_16216,N_19409);
nand U21720 (N_21720,N_17710,N_19594);
or U21721 (N_21721,N_18818,N_16175);
and U21722 (N_21722,N_16698,N_16008);
or U21723 (N_21723,N_19893,N_17073);
xnor U21724 (N_21724,N_18720,N_18007);
and U21725 (N_21725,N_18217,N_18184);
nor U21726 (N_21726,N_19818,N_16919);
xor U21727 (N_21727,N_18527,N_16687);
nor U21728 (N_21728,N_16777,N_16308);
xnor U21729 (N_21729,N_16180,N_17243);
nor U21730 (N_21730,N_17037,N_17858);
and U21731 (N_21731,N_19358,N_15066);
nor U21732 (N_21732,N_18221,N_16347);
nand U21733 (N_21733,N_16875,N_19388);
nor U21734 (N_21734,N_18622,N_15325);
nand U21735 (N_21735,N_18823,N_16004);
nand U21736 (N_21736,N_15075,N_16284);
xor U21737 (N_21737,N_17323,N_18981);
nor U21738 (N_21738,N_16775,N_15337);
nand U21739 (N_21739,N_19543,N_18541);
or U21740 (N_21740,N_17176,N_15018);
and U21741 (N_21741,N_18309,N_17495);
and U21742 (N_21742,N_18802,N_18290);
nand U21743 (N_21743,N_19127,N_16022);
xor U21744 (N_21744,N_16067,N_18564);
nor U21745 (N_21745,N_18952,N_17141);
nor U21746 (N_21746,N_17975,N_16691);
and U21747 (N_21747,N_15711,N_18216);
xnor U21748 (N_21748,N_15029,N_15496);
nor U21749 (N_21749,N_15314,N_16558);
and U21750 (N_21750,N_15452,N_16702);
nand U21751 (N_21751,N_17821,N_17764);
nor U21752 (N_21752,N_18895,N_18259);
or U21753 (N_21753,N_18803,N_15985);
nor U21754 (N_21754,N_19383,N_18795);
and U21755 (N_21755,N_17067,N_16148);
xnor U21756 (N_21756,N_15441,N_16505);
or U21757 (N_21757,N_18296,N_19032);
or U21758 (N_21758,N_17650,N_16918);
xor U21759 (N_21759,N_16551,N_16963);
xnor U21760 (N_21760,N_19218,N_15942);
and U21761 (N_21761,N_18095,N_15449);
and U21762 (N_21762,N_17682,N_18691);
xor U21763 (N_21763,N_17615,N_19152);
xnor U21764 (N_21764,N_17552,N_19579);
nor U21765 (N_21765,N_16778,N_18540);
nor U21766 (N_21766,N_15199,N_17292);
nor U21767 (N_21767,N_19607,N_16800);
nor U21768 (N_21768,N_15549,N_17896);
and U21769 (N_21769,N_18747,N_17361);
xnor U21770 (N_21770,N_17412,N_19410);
nor U21771 (N_21771,N_18636,N_19551);
nor U21772 (N_21772,N_17584,N_17191);
nand U21773 (N_21773,N_16605,N_17854);
nand U21774 (N_21774,N_15751,N_15049);
xnor U21775 (N_21775,N_15020,N_19250);
or U21776 (N_21776,N_15223,N_19856);
or U21777 (N_21777,N_15155,N_15385);
and U21778 (N_21778,N_19865,N_17129);
nand U21779 (N_21779,N_16341,N_15920);
or U21780 (N_21780,N_15235,N_18738);
nor U21781 (N_21781,N_18376,N_17628);
nor U21782 (N_21782,N_19036,N_15137);
nand U21783 (N_21783,N_15204,N_19718);
nand U21784 (N_21784,N_15465,N_16478);
and U21785 (N_21785,N_16226,N_19168);
or U21786 (N_21786,N_17472,N_18729);
nor U21787 (N_21787,N_17846,N_17217);
nand U21788 (N_21788,N_15731,N_18832);
xor U21789 (N_21789,N_18156,N_15358);
and U21790 (N_21790,N_18291,N_15752);
or U21791 (N_21791,N_19762,N_17447);
nor U21792 (N_21792,N_15646,N_17375);
xor U21793 (N_21793,N_18764,N_16923);
or U21794 (N_21794,N_15082,N_15821);
xor U21795 (N_21795,N_15685,N_19669);
nand U21796 (N_21796,N_15175,N_19414);
and U21797 (N_21797,N_19395,N_17407);
or U21798 (N_21798,N_16335,N_15138);
nor U21799 (N_21799,N_19729,N_16071);
and U21800 (N_21800,N_16285,N_15372);
nor U21801 (N_21801,N_19530,N_19507);
nor U21802 (N_21802,N_15491,N_16629);
nand U21803 (N_21803,N_15959,N_18158);
xor U21804 (N_21804,N_16651,N_17852);
nor U21805 (N_21805,N_18103,N_15003);
xor U21806 (N_21806,N_19606,N_15019);
xor U21807 (N_21807,N_18106,N_18213);
or U21808 (N_21808,N_17577,N_15922);
xor U21809 (N_21809,N_17040,N_17909);
nand U21810 (N_21810,N_15975,N_19090);
or U21811 (N_21811,N_17553,N_15433);
xnor U21812 (N_21812,N_15257,N_17520);
xor U21813 (N_21813,N_16926,N_15518);
or U21814 (N_21814,N_16704,N_18122);
nand U21815 (N_21815,N_15597,N_18514);
and U21816 (N_21816,N_16899,N_19379);
and U21817 (N_21817,N_17921,N_15840);
and U21818 (N_21818,N_15596,N_19211);
nand U21819 (N_21819,N_17161,N_18084);
nor U21820 (N_21820,N_16097,N_19558);
and U21821 (N_21821,N_18716,N_19174);
or U21822 (N_21822,N_18180,N_16330);
nand U21823 (N_21823,N_17889,N_15769);
xor U21824 (N_21824,N_19467,N_19563);
or U21825 (N_21825,N_18011,N_15159);
nand U21826 (N_21826,N_16557,N_17807);
nor U21827 (N_21827,N_16841,N_15099);
or U21828 (N_21828,N_16185,N_15839);
nor U21829 (N_21829,N_19363,N_16688);
nor U21830 (N_21830,N_19172,N_19682);
nand U21831 (N_21831,N_15002,N_19807);
or U21832 (N_21832,N_18401,N_18019);
or U21833 (N_21833,N_17964,N_18304);
nand U21834 (N_21834,N_15590,N_15729);
xnor U21835 (N_21835,N_17910,N_19660);
nor U21836 (N_21836,N_19714,N_19872);
nand U21837 (N_21837,N_19230,N_17545);
or U21838 (N_21838,N_17406,N_17787);
nor U21839 (N_21839,N_16258,N_16289);
nor U21840 (N_21840,N_16842,N_19441);
or U21841 (N_21841,N_15847,N_15994);
and U21842 (N_21842,N_19929,N_17357);
and U21843 (N_21843,N_19982,N_19468);
and U21844 (N_21844,N_17101,N_15669);
xnor U21845 (N_21845,N_19077,N_16660);
nand U21846 (N_21846,N_16424,N_19425);
or U21847 (N_21847,N_15443,N_15162);
nor U21848 (N_21848,N_19652,N_16032);
and U21849 (N_21849,N_18412,N_17336);
xor U21850 (N_21850,N_15056,N_19076);
xnor U21851 (N_21851,N_19556,N_15389);
or U21852 (N_21852,N_17959,N_15439);
nor U21853 (N_21853,N_17151,N_15564);
xnor U21854 (N_21854,N_18049,N_15579);
nand U21855 (N_21855,N_15485,N_19067);
nand U21856 (N_21856,N_18074,N_15157);
nor U21857 (N_21857,N_15263,N_19593);
nand U21858 (N_21858,N_19122,N_17790);
xnor U21859 (N_21859,N_19157,N_15802);
and U21860 (N_21860,N_17206,N_18230);
xor U21861 (N_21861,N_15608,N_18075);
nand U21862 (N_21862,N_17435,N_15768);
and U21863 (N_21863,N_19440,N_18203);
xnor U21864 (N_21864,N_16269,N_16154);
nor U21865 (N_21865,N_18507,N_17227);
nand U21866 (N_21866,N_18484,N_15486);
nand U21867 (N_21867,N_18806,N_16772);
and U21868 (N_21868,N_19964,N_19196);
nand U21869 (N_21869,N_17620,N_19541);
nor U21870 (N_21870,N_16809,N_19854);
nor U21871 (N_21871,N_17533,N_16122);
and U21872 (N_21872,N_19911,N_15910);
and U21873 (N_21873,N_17135,N_16093);
nand U21874 (N_21874,N_15422,N_17630);
and U21875 (N_21875,N_15616,N_15526);
xor U21876 (N_21876,N_17443,N_16856);
xnor U21877 (N_21877,N_16857,N_18647);
or U21878 (N_21878,N_18543,N_15161);
and U21879 (N_21879,N_19186,N_19116);
nand U21880 (N_21880,N_16458,N_18519);
nand U21881 (N_21881,N_16866,N_18045);
and U21882 (N_21882,N_18539,N_18477);
xnor U21883 (N_21883,N_18695,N_19353);
xor U21884 (N_21884,N_17115,N_18966);
or U21885 (N_21885,N_19830,N_19355);
nand U21886 (N_21886,N_16365,N_17523);
or U21887 (N_21887,N_17110,N_15353);
and U21888 (N_21888,N_18985,N_15134);
or U21889 (N_21889,N_16521,N_15992);
and U21890 (N_21890,N_16080,N_17118);
nand U21891 (N_21891,N_17281,N_17349);
nor U21892 (N_21892,N_19350,N_17154);
xnor U21893 (N_21893,N_19619,N_18486);
or U21894 (N_21894,N_17775,N_18163);
or U21895 (N_21895,N_17939,N_19120);
and U21896 (N_21896,N_17619,N_19098);
nand U21897 (N_21897,N_17812,N_18192);
or U21898 (N_21898,N_18637,N_15346);
and U21899 (N_21899,N_18696,N_18293);
nand U21900 (N_21900,N_18689,N_18054);
and U21901 (N_21901,N_17773,N_15970);
nand U21902 (N_21902,N_19150,N_15519);
nand U21903 (N_21903,N_18353,N_19962);
and U21904 (N_21904,N_19864,N_18394);
nand U21905 (N_21905,N_15015,N_17512);
nand U21906 (N_21906,N_17358,N_16545);
and U21907 (N_21907,N_19046,N_15348);
nand U21908 (N_21908,N_17445,N_17387);
or U21909 (N_21909,N_16974,N_16394);
xor U21910 (N_21910,N_18524,N_15648);
and U21911 (N_21911,N_16153,N_15463);
nor U21912 (N_21912,N_19837,N_18448);
or U21913 (N_21913,N_18638,N_19480);
or U21914 (N_21914,N_16316,N_19721);
xor U21915 (N_21915,N_17564,N_15516);
xnor U21916 (N_21916,N_17181,N_18796);
xor U21917 (N_21917,N_15004,N_16126);
and U21918 (N_21918,N_15968,N_17664);
and U21919 (N_21919,N_15205,N_17088);
nor U21920 (N_21920,N_19462,N_18858);
nand U21921 (N_21921,N_18121,N_18554);
nor U21922 (N_21922,N_15126,N_16769);
or U21923 (N_21923,N_19989,N_16172);
nand U21924 (N_21924,N_19515,N_15415);
or U21925 (N_21925,N_17566,N_15483);
or U21926 (N_21926,N_15586,N_17278);
xor U21927 (N_21927,N_18337,N_16215);
nand U21928 (N_21928,N_16969,N_19537);
or U21929 (N_21929,N_19399,N_15989);
nor U21930 (N_21930,N_15265,N_19781);
xor U21931 (N_21931,N_19273,N_19769);
xor U21932 (N_21932,N_17391,N_18861);
or U21933 (N_21933,N_17408,N_19927);
nor U21934 (N_21934,N_17015,N_18956);
nor U21935 (N_21935,N_17260,N_16417);
nand U21936 (N_21936,N_19695,N_17120);
and U21937 (N_21937,N_17678,N_16590);
nand U21938 (N_21938,N_15796,N_18772);
nand U21939 (N_21939,N_19501,N_19878);
nor U21940 (N_21940,N_18176,N_17365);
or U21941 (N_21941,N_17104,N_19681);
nor U21942 (N_21942,N_19926,N_17804);
nand U21943 (N_21943,N_16156,N_18629);
and U21944 (N_21944,N_16755,N_19222);
or U21945 (N_21945,N_17318,N_15503);
nand U21946 (N_21946,N_19519,N_18124);
or U21947 (N_21947,N_18155,N_19210);
and U21948 (N_21948,N_18393,N_15193);
nand U21949 (N_21949,N_15118,N_19163);
or U21950 (N_21950,N_17605,N_18690);
nor U21951 (N_21951,N_17508,N_19387);
xor U21952 (N_21952,N_17469,N_16057);
nand U21953 (N_21953,N_16980,N_19499);
nand U21954 (N_21954,N_15275,N_15946);
nor U21955 (N_21955,N_17758,N_17954);
nand U21956 (N_21956,N_17453,N_19724);
xnor U21957 (N_21957,N_15133,N_15659);
or U21958 (N_21958,N_18489,N_16221);
or U21959 (N_21959,N_19588,N_18418);
xnor U21960 (N_21960,N_16480,N_15419);
xor U21961 (N_21961,N_16017,N_15638);
nor U21962 (N_21962,N_15290,N_15370);
nand U21963 (N_21963,N_16589,N_18094);
and U21964 (N_21964,N_19247,N_15258);
and U21965 (N_21965,N_19615,N_18884);
xor U21966 (N_21966,N_17429,N_17457);
and U21967 (N_21967,N_19858,N_15227);
xnor U21968 (N_21968,N_17399,N_16607);
nor U21969 (N_21969,N_17856,N_19710);
xnor U21970 (N_21970,N_17450,N_18943);
or U21971 (N_21971,N_19088,N_15431);
or U21972 (N_21972,N_15585,N_18719);
nor U21973 (N_21973,N_16964,N_19664);
nor U21974 (N_21974,N_19540,N_19738);
and U21975 (N_21975,N_15521,N_18417);
xor U21976 (N_21976,N_15100,N_18748);
xor U21977 (N_21977,N_18653,N_18782);
nand U21978 (N_21978,N_18830,N_15733);
nand U21979 (N_21979,N_18086,N_16204);
nand U21980 (N_21980,N_16925,N_15898);
or U21981 (N_21981,N_15684,N_18247);
xnor U21982 (N_21982,N_15636,N_19248);
nor U21983 (N_21983,N_17971,N_16726);
xor U21984 (N_21984,N_15124,N_15978);
nand U21985 (N_21985,N_19275,N_18550);
nand U21986 (N_21986,N_17229,N_17549);
xor U21987 (N_21987,N_15131,N_15870);
nor U21988 (N_21988,N_18983,N_18469);
nor U21989 (N_21989,N_16044,N_19779);
and U21990 (N_21990,N_18085,N_19888);
or U21991 (N_21991,N_17532,N_17261);
xor U21992 (N_21992,N_17601,N_18101);
or U21993 (N_21993,N_15599,N_16282);
nand U21994 (N_21994,N_16951,N_16188);
nor U21995 (N_21995,N_15766,N_16555);
or U21996 (N_21996,N_16436,N_16390);
or U21997 (N_21997,N_18178,N_16023);
nand U21998 (N_21998,N_19004,N_18903);
nor U21999 (N_21999,N_18251,N_16058);
xor U22000 (N_22000,N_19800,N_15918);
or U22001 (N_22001,N_19000,N_15721);
xnor U22002 (N_22002,N_15413,N_18909);
and U22003 (N_22003,N_17273,N_19774);
or U22004 (N_22004,N_19384,N_16075);
xor U22005 (N_22005,N_19569,N_16399);
or U22006 (N_22006,N_17595,N_17380);
nand U22007 (N_22007,N_18513,N_16536);
nor U22008 (N_22008,N_16636,N_18082);
nor U22009 (N_22009,N_15654,N_19884);
and U22010 (N_22010,N_16670,N_16392);
nor U22011 (N_22011,N_19874,N_15842);
xor U22012 (N_22012,N_19402,N_15215);
xor U22013 (N_22013,N_16141,N_19193);
nand U22014 (N_22014,N_18588,N_19971);
nand U22015 (N_22015,N_15632,N_15363);
xnor U22016 (N_22016,N_18083,N_15450);
nor U22017 (N_22017,N_16546,N_15179);
xnor U22018 (N_22018,N_15359,N_19432);
or U22019 (N_22019,N_15925,N_19571);
nor U22020 (N_22020,N_18396,N_16635);
nand U22021 (N_22021,N_18509,N_18904);
nand U22022 (N_22022,N_17113,N_15000);
and U22023 (N_22023,N_18272,N_17996);
and U22024 (N_22024,N_19778,N_16380);
and U22025 (N_22025,N_15722,N_16585);
and U22026 (N_22026,N_16292,N_16320);
and U22027 (N_22027,N_15225,N_17637);
nand U22028 (N_22028,N_16787,N_16489);
nor U22029 (N_22029,N_18657,N_15482);
and U22030 (N_22030,N_17930,N_17924);
or U22031 (N_22031,N_17289,N_15613);
nand U22032 (N_22032,N_16680,N_15853);
and U22033 (N_22033,N_18736,N_18281);
nand U22034 (N_22034,N_16976,N_15144);
nor U22035 (N_22035,N_16350,N_15961);
xnor U22036 (N_22036,N_17434,N_19304);
nor U22037 (N_22037,N_18627,N_18166);
xor U22038 (N_22038,N_16240,N_19635);
nor U22039 (N_22039,N_17786,N_16479);
or U22040 (N_22040,N_15695,N_16239);
or U22041 (N_22041,N_17640,N_18760);
nor U22042 (N_22042,N_16984,N_19746);
and U22043 (N_22043,N_15354,N_16647);
and U22044 (N_22044,N_19749,N_19188);
nor U22045 (N_22045,N_18215,N_16947);
xnor U22046 (N_22046,N_16043,N_19262);
or U22047 (N_22047,N_18113,N_18775);
xnor U22048 (N_22048,N_17049,N_19171);
xor U22049 (N_22049,N_15689,N_15672);
nor U22050 (N_22050,N_16361,N_17185);
xor U22051 (N_22051,N_19491,N_15120);
nor U22052 (N_22052,N_19466,N_17403);
nand U22053 (N_22053,N_15288,N_16806);
and U22054 (N_22054,N_16457,N_16851);
xor U22055 (N_22055,N_15404,N_17355);
xor U22056 (N_22056,N_16578,N_15424);
nand U22057 (N_22057,N_19179,N_18258);
nand U22058 (N_22058,N_19007,N_16198);
and U22059 (N_22059,N_17341,N_16190);
nor U22060 (N_22060,N_18364,N_17940);
xor U22061 (N_22061,N_17629,N_19319);
or U22062 (N_22062,N_16177,N_16194);
xnor U22063 (N_22063,N_19014,N_18639);
nor U22064 (N_22064,N_19189,N_16825);
nor U22065 (N_22065,N_19959,N_15593);
and U22066 (N_22066,N_18610,N_19768);
or U22067 (N_22067,N_18930,N_19717);
nand U22068 (N_22068,N_19173,N_19101);
nor U22069 (N_22069,N_17983,N_16506);
and U22070 (N_22070,N_17670,N_15628);
nand U22071 (N_22071,N_15103,N_17955);
xor U22072 (N_22072,N_16771,N_19553);
or U22073 (N_22073,N_17999,N_16878);
nand U22074 (N_22074,N_16618,N_15156);
nor U22075 (N_22075,N_18561,N_18617);
or U22076 (N_22076,N_18987,N_19528);
xnor U22077 (N_22077,N_17535,N_17196);
nor U22078 (N_22078,N_18200,N_16297);
nor U22079 (N_22079,N_17526,N_15035);
or U22080 (N_22080,N_15801,N_19719);
nor U22081 (N_22081,N_16090,N_18620);
nand U22082 (N_22082,N_15808,N_18234);
xor U22083 (N_22083,N_15068,N_17824);
nor U22084 (N_22084,N_16359,N_17376);
xnor U22085 (N_22085,N_19306,N_18671);
nor U22086 (N_22086,N_19882,N_15173);
xnor U22087 (N_22087,N_15945,N_15408);
or U22088 (N_22088,N_17043,N_18495);
and U22089 (N_22089,N_19622,N_19508);
or U22090 (N_22090,N_17912,N_18347);
nand U22091 (N_22091,N_19177,N_17164);
xnor U22092 (N_22092,N_16945,N_18378);
and U22093 (N_22093,N_18681,N_16136);
nor U22094 (N_22094,N_16300,N_16815);
and U22095 (N_22095,N_17248,N_16343);
and U22096 (N_22096,N_18276,N_19367);
nor U22097 (N_22097,N_18009,N_17529);
or U22098 (N_22098,N_17003,N_19527);
xor U22099 (N_22099,N_18039,N_16149);
xor U22100 (N_22100,N_17096,N_16913);
xnor U22101 (N_22101,N_18405,N_16944);
xor U22102 (N_22102,N_16978,N_18774);
or U22103 (N_22103,N_18400,N_16120);
nand U22104 (N_22104,N_15759,N_15655);
nand U22105 (N_22105,N_15291,N_17931);
xor U22106 (N_22106,N_19277,N_17977);
nand U22107 (N_22107,N_19278,N_15360);
nand U22108 (N_22108,N_18096,N_18846);
xor U22109 (N_22109,N_19469,N_19909);
and U22110 (N_22110,N_18087,N_16912);
or U22111 (N_22111,N_19967,N_18034);
nand U22112 (N_22112,N_19851,N_17020);
nand U22113 (N_22113,N_19459,N_15984);
or U22114 (N_22114,N_17048,N_17303);
nor U22115 (N_22115,N_19235,N_15799);
nand U22116 (N_22116,N_15895,N_16461);
nor U22117 (N_22117,N_17396,N_18140);
xnor U22118 (N_22118,N_19408,N_19147);
or U22119 (N_22119,N_18431,N_18683);
and U22120 (N_22120,N_19981,N_15836);
nor U22121 (N_22121,N_18236,N_17304);
nand U22122 (N_22122,N_18473,N_16303);
and U22123 (N_22123,N_17980,N_19371);
xnor U22124 (N_22124,N_15495,N_19789);
nor U22125 (N_22125,N_16266,N_19857);
or U22126 (N_22126,N_17809,N_18024);
xnor U22127 (N_22127,N_18517,N_15666);
xnor U22128 (N_22128,N_16814,N_15453);
xor U22129 (N_22129,N_18294,N_18761);
xnor U22130 (N_22130,N_17290,N_19675);
nand U22131 (N_22131,N_17687,N_15081);
nand U22132 (N_22132,N_18890,N_15073);
nor U22133 (N_22133,N_19889,N_18700);
xor U22134 (N_22134,N_18609,N_19276);
and U22135 (N_22135,N_15034,N_16274);
and U22136 (N_22136,N_19896,N_18812);
nor U22137 (N_22137,N_15614,N_18606);
and U22138 (N_22138,N_16000,N_19741);
and U22139 (N_22139,N_17633,N_18790);
and U22140 (N_22140,N_15533,N_16782);
and U22141 (N_22141,N_19106,N_16406);
and U22142 (N_22142,N_19376,N_16187);
nand U22143 (N_22143,N_17979,N_15050);
nand U22144 (N_22144,N_15591,N_15905);
and U22145 (N_22145,N_19704,N_18149);
or U22146 (N_22146,N_16205,N_15434);
xor U22147 (N_22147,N_15283,N_15960);
nand U22148 (N_22148,N_17474,N_19472);
and U22149 (N_22149,N_15915,N_17570);
nor U22150 (N_22150,N_16144,N_19325);
nand U22151 (N_22151,N_18245,N_19855);
and U22152 (N_22152,N_15913,N_19058);
or U22153 (N_22153,N_16493,N_16026);
nand U22154 (N_22154,N_18977,N_19820);
nor U22155 (N_22155,N_18855,N_18933);
nor U22156 (N_22156,N_19016,N_18990);
nor U22157 (N_22157,N_17654,N_16203);
xor U22158 (N_22158,N_16902,N_18717);
or U22159 (N_22159,N_16360,N_19200);
or U22160 (N_22160,N_15785,N_16373);
xor U22161 (N_22161,N_16848,N_19249);
and U22162 (N_22162,N_15154,N_15338);
nor U22163 (N_22163,N_19237,N_17155);
xor U22164 (N_22164,N_15282,N_19649);
or U22165 (N_22165,N_19735,N_19461);
nand U22166 (N_22166,N_18128,N_15860);
xor U22167 (N_22167,N_17694,N_15953);
and U22168 (N_22168,N_18845,N_18817);
and U22169 (N_22169,N_17830,N_17805);
and U22170 (N_22170,N_17770,N_16939);
or U22171 (N_22171,N_17496,N_18506);
and U22172 (N_22172,N_18043,N_17416);
xnor U22173 (N_22173,N_19012,N_15274);
nor U22174 (N_22174,N_17360,N_17202);
or U22175 (N_22175,N_17393,N_17781);
or U22176 (N_22176,N_19640,N_15668);
and U22177 (N_22177,N_15322,N_19809);
nand U22178 (N_22178,N_18468,N_19337);
or U22179 (N_22179,N_18190,N_18193);
nand U22180 (N_22180,N_18615,N_19871);
and U22181 (N_22181,N_15912,N_17317);
or U22182 (N_22182,N_18641,N_18065);
or U22183 (N_22183,N_17130,N_17668);
nand U22184 (N_22184,N_18628,N_15916);
nor U22185 (N_22185,N_17597,N_17235);
or U22186 (N_22186,N_19708,N_15807);
nand U22187 (N_22187,N_19621,N_17957);
or U22188 (N_22188,N_15304,N_19203);
nand U22189 (N_22189,N_18718,N_17903);
nor U22190 (N_22190,N_18270,N_16184);
or U22191 (N_22191,N_17753,N_18256);
xor U22192 (N_22192,N_17034,N_19403);
nor U22193 (N_22193,N_15249,N_18350);
nor U22194 (N_22194,N_15417,N_16275);
and U22195 (N_22195,N_15814,N_16116);
or U22196 (N_22196,N_15067,N_15319);
nor U22197 (N_22197,N_18905,N_18553);
nand U22198 (N_22198,N_15247,N_17258);
and U22199 (N_22199,N_19449,N_17516);
and U22200 (N_22200,N_19215,N_16028);
nand U22201 (N_22201,N_15627,N_15305);
xnor U22202 (N_22202,N_18563,N_19887);
nor U22203 (N_22203,N_18438,N_18958);
nor U22204 (N_22204,N_16317,N_16715);
or U22205 (N_22205,N_16941,N_16780);
xnor U22206 (N_22206,N_15069,N_18194);
or U22207 (N_22207,N_17353,N_19063);
or U22208 (N_22208,N_15243,N_17754);
nand U22209 (N_22209,N_18560,N_18878);
xnor U22210 (N_22210,N_16538,N_19993);
nand U22211 (N_22211,N_17917,N_17253);
nand U22212 (N_22212,N_15661,N_15522);
and U22213 (N_22213,N_17574,N_16796);
and U22214 (N_22214,N_19065,N_15677);
nor U22215 (N_22215,N_17269,N_16879);
and U22216 (N_22216,N_16054,N_19241);
xnor U22217 (N_22217,N_19931,N_16807);
or U22218 (N_22218,N_18191,N_17186);
xnor U22219 (N_22219,N_16690,N_17632);
xor U22220 (N_22220,N_15135,N_16859);
or U22221 (N_22221,N_18708,N_15589);
xnor U22222 (N_22222,N_19450,N_18558);
or U22223 (N_22223,N_19452,N_16512);
nor U22224 (N_22224,N_16474,N_15078);
xnor U22225 (N_22225,N_18325,N_16768);
nand U22226 (N_22226,N_16412,N_15242);
nor U22227 (N_22227,N_19176,N_18827);
xnor U22228 (N_22228,N_17641,N_17752);
and U22229 (N_22229,N_16934,N_19167);
xnor U22230 (N_22230,N_19648,N_16513);
nor U22231 (N_22231,N_19827,N_18112);
or U22232 (N_22232,N_18223,N_19957);
or U22233 (N_22233,N_18185,N_16333);
nand U22234 (N_22234,N_18508,N_19819);
nor U22235 (N_22235,N_19709,N_18993);
nand U22236 (N_22236,N_18037,N_15547);
or U22237 (N_22237,N_15253,N_16115);
and U22238 (N_22238,N_17521,N_15633);
nor U22239 (N_22239,N_19567,N_16358);
xor U22240 (N_22240,N_16756,N_18447);
xor U22241 (N_22241,N_15336,N_18674);
nand U22242 (N_22242,N_19511,N_17080);
and U22243 (N_22243,N_18925,N_19629);
or U22244 (N_22244,N_19020,N_19314);
nand U22245 (N_22245,N_15717,N_15806);
nor U22246 (N_22246,N_16641,N_18953);
nor U22247 (N_22247,N_15517,N_17881);
and U22248 (N_22248,N_18789,N_16082);
xor U22249 (N_22249,N_19108,N_18138);
and U22250 (N_22250,N_17581,N_16936);
or U22251 (N_22251,N_16395,N_15287);
and U22252 (N_22252,N_15949,N_15198);
and U22253 (N_22253,N_19788,N_16564);
or U22254 (N_22254,N_18778,N_19072);
nand U22255 (N_22255,N_15714,N_19181);
nor U22256 (N_22256,N_15973,N_15089);
and U22257 (N_22257,N_16464,N_19726);
nand U22258 (N_22258,N_16646,N_15396);
and U22259 (N_22259,N_16759,N_18205);
or U22260 (N_22260,N_19042,N_18206);
nor U22261 (N_22261,N_19407,N_17864);
and U22262 (N_22262,N_17044,N_17294);
nor U22263 (N_22263,N_17563,N_18254);
xor U22264 (N_22264,N_19321,N_19284);
or U22265 (N_22265,N_17092,N_17084);
xor U22266 (N_22266,N_16143,N_16507);
and U22267 (N_22267,N_19279,N_18991);
and U22268 (N_22268,N_17757,N_16312);
and U22269 (N_22269,N_18071,N_18016);
and U22270 (N_22270,N_15952,N_18576);
xor U22271 (N_22271,N_19954,N_16158);
nand U22272 (N_22272,N_15743,N_17877);
xor U22273 (N_22273,N_19570,N_15704);
and U22274 (N_22274,N_17618,N_18922);
or U22275 (N_22275,N_17371,N_19087);
and U22276 (N_22276,N_19513,N_18759);
nor U22277 (N_22277,N_15403,N_17201);
or U22278 (N_22278,N_15462,N_17094);
or U22279 (N_22279,N_16940,N_17718);
nand U22280 (N_22280,N_16733,N_15753);
xor U22281 (N_22281,N_17499,N_17366);
or U22282 (N_22282,N_19369,N_19155);
or U22283 (N_22283,N_17911,N_16488);
or U22284 (N_22284,N_16522,N_15252);
nor U22285 (N_22285,N_19792,N_15809);
xor U22286 (N_22286,N_19859,N_18665);
nor U22287 (N_22287,N_16339,N_18238);
and U22288 (N_22288,N_18574,N_15820);
nor U22289 (N_22289,N_16659,N_17256);
nor U22290 (N_22290,N_16473,N_19298);
or U22291 (N_22291,N_19474,N_18491);
nand U22292 (N_22292,N_19001,N_15617);
nor U22293 (N_22293,N_15742,N_19514);
and U22294 (N_22294,N_16735,N_16872);
and U22295 (N_22295,N_17929,N_17471);
or U22296 (N_22296,N_18025,N_19330);
nor U22297 (N_22297,N_19542,N_16088);
or U22298 (N_22298,N_18571,N_19873);
nand U22299 (N_22299,N_18004,N_18051);
nor U22300 (N_22300,N_19154,N_15550);
xor U22301 (N_22301,N_19359,N_15651);
and U22302 (N_22302,N_19340,N_18165);
or U22303 (N_22303,N_18260,N_18371);
nor U22304 (N_22304,N_15481,N_18000);
xor U22305 (N_22305,N_15691,N_17342);
nand U22306 (N_22306,N_15640,N_16533);
nand U22307 (N_22307,N_15115,N_19986);
and U22308 (N_22308,N_16721,N_17388);
and U22309 (N_22309,N_16201,N_19580);
and U22310 (N_22310,N_15260,N_18634);
nand U22311 (N_22311,N_17156,N_19308);
xnor U22312 (N_22312,N_16351,N_18766);
nor U22313 (N_22313,N_16603,N_15317);
and U22314 (N_22314,N_17747,N_18927);
nor U22315 (N_22315,N_17547,N_18829);
nor U22316 (N_22316,N_17602,N_17548);
nor U22317 (N_22317,N_16999,N_16107);
nand U22318 (N_22318,N_17417,N_15183);
or U22319 (N_22319,N_18532,N_15563);
nand U22320 (N_22320,N_15121,N_18188);
or U22321 (N_22321,N_19204,N_18880);
nor U22322 (N_22322,N_16309,N_15557);
nor U22323 (N_22323,N_16016,N_15800);
nor U22324 (N_22324,N_16481,N_19578);
and U22325 (N_22325,N_18483,N_18253);
or U22326 (N_22326,N_17649,N_16230);
nand U22327 (N_22327,N_19444,N_15525);
nand U22328 (N_22328,N_16294,N_17207);
and U22329 (N_22329,N_19839,N_16811);
or U22330 (N_22330,N_15084,N_17414);
nor U22331 (N_22331,N_19831,N_19814);
or U22332 (N_22332,N_19706,N_15065);
nand U22333 (N_22333,N_15196,N_18306);
xnor U22334 (N_22334,N_19223,N_15226);
nand U22335 (N_22335,N_15738,N_15489);
or U22336 (N_22336,N_16850,N_18877);
or U22337 (N_22337,N_18358,N_18175);
nand U22338 (N_22338,N_17449,N_15986);
and U22339 (N_22339,N_18611,N_16846);
and U22340 (N_22340,N_16920,N_18292);
nor U22341 (N_22341,N_18791,N_18614);
nand U22342 (N_22342,N_18529,N_17379);
nand U22343 (N_22343,N_18501,N_15109);
xor U22344 (N_22344,N_19099,N_15673);
or U22345 (N_22345,N_17802,N_17582);
nor U22346 (N_22346,N_15600,N_17756);
nand U22347 (N_22347,N_16730,N_19693);
and U22348 (N_22348,N_15311,N_17610);
xor U22349 (N_22349,N_18934,N_18229);
xnor U22350 (N_22350,N_17137,N_16729);
nand U22351 (N_22351,N_17473,N_17390);
and U22352 (N_22352,N_15535,N_18562);
nand U22353 (N_22353,N_17991,N_18768);
and U22354 (N_22354,N_16795,N_16958);
or U22355 (N_22355,N_19583,N_19138);
xor U22356 (N_22356,N_18001,N_16328);
or U22357 (N_22357,N_16588,N_18770);
or U22358 (N_22358,N_16986,N_19263);
or U22359 (N_22359,N_17004,N_18301);
nor U22360 (N_22360,N_19947,N_18741);
nand U22361 (N_22361,N_18157,N_19484);
nand U22362 (N_22362,N_17063,N_16763);
xor U22363 (N_22363,N_15017,N_17536);
nor U22364 (N_22364,N_19243,N_15244);
xor U22365 (N_22365,N_17684,N_16765);
nor U22366 (N_22366,N_18552,N_16084);
nand U22367 (N_22367,N_17701,N_18921);
or U22368 (N_22368,N_16804,N_19824);
nand U22369 (N_22369,N_18569,N_16152);
nor U22370 (N_22370,N_15707,N_19418);
nor U22371 (N_22371,N_17335,N_16661);
nand U22372 (N_22372,N_19812,N_15849);
nor U22373 (N_22373,N_16836,N_16200);
nand U22374 (N_22374,N_17309,N_18593);
or U22375 (N_22375,N_15581,N_17937);
nand U22376 (N_22376,N_19791,N_19435);
xnor U22377 (N_22377,N_17313,N_18528);
xnor U22378 (N_22378,N_15022,N_15943);
xnor U22379 (N_22379,N_19125,N_18250);
and U22380 (N_22380,N_16114,N_15856);
nor U22381 (N_22381,N_17014,N_18145);
and U22382 (N_22382,N_17603,N_19103);
nand U22383 (N_22383,N_18423,N_16467);
and U22384 (N_22384,N_15166,N_18723);
and U22385 (N_22385,N_18712,N_18240);
nand U22386 (N_22386,N_18424,N_18619);
nor U22387 (N_22387,N_15010,N_15754);
xnor U22388 (N_22388,N_17765,N_15140);
nand U22389 (N_22389,N_17199,N_17029);
nand U22390 (N_22390,N_15505,N_19923);
xnor U22391 (N_22391,N_18467,N_18662);
nand U22392 (N_22392,N_16104,N_17944);
or U22393 (N_22393,N_19897,N_18498);
xor U22394 (N_22394,N_18332,N_17750);
and U22395 (N_22395,N_15387,N_17783);
nand U22396 (N_22396,N_16252,N_16442);
xnor U22397 (N_22397,N_17984,N_17052);
nor U22398 (N_22398,N_18697,N_18908);
and U22399 (N_22399,N_17058,N_18677);
nor U22400 (N_22400,N_19522,N_18714);
nand U22401 (N_22401,N_19013,N_15509);
nand U22402 (N_22402,N_17915,N_16010);
or U22403 (N_22403,N_18115,N_19650);
nand U22404 (N_22404,N_18850,N_17409);
or U22405 (N_22405,N_16808,N_16432);
or U22406 (N_22406,N_17418,N_16247);
nand U22407 (N_22407,N_19922,N_17792);
nor U22408 (N_22408,N_16119,N_16233);
xnor U22409 (N_22409,N_17263,N_15341);
xor U22410 (N_22410,N_15755,N_18725);
and U22411 (N_22411,N_16930,N_18319);
xor U22412 (N_22412,N_17359,N_18189);
nand U22413 (N_22413,N_19616,N_16937);
nor U22414 (N_22414,N_17351,N_17082);
and U22415 (N_22415,N_15303,N_19904);
or U22416 (N_22416,N_16907,N_19288);
and U22417 (N_22417,N_16109,N_15256);
and U22418 (N_22418,N_19796,N_15530);
nand U22419 (N_22419,N_16433,N_16812);
and U22420 (N_22420,N_17544,N_19015);
nor U22421 (N_22421,N_19572,N_15594);
xnor U22422 (N_22422,N_17847,N_15468);
nand U22423 (N_22423,N_16552,N_15063);
nand U22424 (N_22424,N_19034,N_17239);
xnor U22425 (N_22425,N_17124,N_18346);
or U22426 (N_22426,N_18432,N_19380);
nor U22427 (N_22427,N_15854,N_16501);
nand U22428 (N_22428,N_18098,N_18591);
nor U22429 (N_22429,N_18894,N_18754);
nor U22430 (N_22430,N_15071,N_17404);
xnor U22431 (N_22431,N_17442,N_16832);
nor U22432 (N_22432,N_15866,N_19975);
and U22433 (N_22433,N_16063,N_18751);
nand U22434 (N_22434,N_15653,N_15635);
or U22435 (N_22435,N_17068,N_17314);
nor U22436 (N_22436,N_15494,N_18871);
or U22437 (N_22437,N_19023,N_16498);
or U22438 (N_22438,N_17482,N_17007);
or U22439 (N_22439,N_18856,N_17214);
and U22440 (N_22440,N_17321,N_15347);
nor U22441 (N_22441,N_19608,N_16739);
xnor U22442 (N_22442,N_19984,N_16267);
nor U22443 (N_22443,N_15899,N_15128);
nand U22444 (N_22444,N_15130,N_16117);
or U22445 (N_22445,N_16627,N_18300);
nand U22446 (N_22446,N_18579,N_18010);
nor U22447 (N_22447,N_18566,N_15080);
xor U22448 (N_22448,N_17683,N_16903);
or U22449 (N_22449,N_19164,N_19496);
xnor U22450 (N_22450,N_17593,N_16348);
nand U22451 (N_22451,N_19255,N_15688);
nor U22452 (N_22452,N_15686,N_15471);
or U22453 (N_22453,N_18559,N_19269);
xor U22454 (N_22454,N_16445,N_16511);
or U22455 (N_22455,N_17997,N_18264);
xor U22456 (N_22456,N_16776,N_17634);
or U22457 (N_22457,N_17119,N_17719);
or U22458 (N_22458,N_17777,N_16495);
nor U22459 (N_22459,N_19683,N_15008);
and U22460 (N_22460,N_16422,N_18195);
nand U22461 (N_22461,N_15333,N_16469);
nor U22462 (N_22462,N_19568,N_16712);
or U22463 (N_22463,N_19997,N_18502);
nand U22464 (N_22464,N_17311,N_17165);
and U22465 (N_22465,N_15190,N_16710);
nor U22466 (N_22466,N_18520,N_19086);
xor U22467 (N_22467,N_15122,N_19039);
and U22468 (N_22468,N_19668,N_19105);
xor U22469 (N_22469,N_17631,N_19510);
or U22470 (N_22470,N_17425,N_16736);
nand U22471 (N_22471,N_15966,N_17241);
nor U22472 (N_22472,N_17170,N_17150);
or U22473 (N_22473,N_15407,N_17594);
xnor U22474 (N_22474,N_19637,N_15781);
xnor U22475 (N_22475,N_16652,N_19633);
or U22476 (N_22476,N_19009,N_15565);
and U22477 (N_22477,N_18031,N_18355);
nor U22478 (N_22478,N_18888,N_17144);
or U22479 (N_22479,N_16164,N_16033);
xor U22480 (N_22480,N_18575,N_15696);
and U22481 (N_22481,N_16791,N_16466);
or U22482 (N_22482,N_19879,N_16717);
xnor U22483 (N_22483,N_17681,N_16529);
nand U22484 (N_22484,N_16222,N_15623);
nand U22485 (N_22485,N_17152,N_16036);
or U22486 (N_22486,N_15160,N_16579);
nand U22487 (N_22487,N_16743,N_16583);
nand U22488 (N_22488,N_15924,N_16413);
xor U22489 (N_22489,N_18777,N_19901);
nor U22490 (N_22490,N_18169,N_19972);
nand U22491 (N_22491,N_16979,N_17645);
xnor U22492 (N_22492,N_16040,N_17023);
nand U22493 (N_22493,N_17868,N_16967);
or U22494 (N_22494,N_17671,N_15701);
or U22495 (N_22495,N_17071,N_17699);
nand U22496 (N_22496,N_15033,N_15386);
nor U22497 (N_22497,N_16283,N_16932);
or U22498 (N_22498,N_19040,N_16244);
xnor U22499 (N_22499,N_16241,N_19209);
and U22500 (N_22500,N_15573,N_19572);
or U22501 (N_22501,N_17213,N_18864);
nand U22502 (N_22502,N_19752,N_16085);
xor U22503 (N_22503,N_17541,N_19851);
nor U22504 (N_22504,N_18850,N_15922);
xor U22505 (N_22505,N_15638,N_15883);
xor U22506 (N_22506,N_18407,N_19694);
xor U22507 (N_22507,N_17603,N_15536);
or U22508 (N_22508,N_18061,N_18103);
nand U22509 (N_22509,N_15405,N_19926);
and U22510 (N_22510,N_17934,N_18375);
nor U22511 (N_22511,N_17177,N_15430);
or U22512 (N_22512,N_15667,N_19349);
nand U22513 (N_22513,N_16011,N_19125);
nor U22514 (N_22514,N_17695,N_16919);
nor U22515 (N_22515,N_17002,N_16048);
nor U22516 (N_22516,N_17623,N_16648);
xnor U22517 (N_22517,N_16809,N_17712);
or U22518 (N_22518,N_19160,N_17151);
xnor U22519 (N_22519,N_18172,N_18118);
or U22520 (N_22520,N_17101,N_17061);
or U22521 (N_22521,N_17790,N_15330);
nor U22522 (N_22522,N_17903,N_15596);
and U22523 (N_22523,N_18159,N_15656);
or U22524 (N_22524,N_15244,N_19874);
and U22525 (N_22525,N_16043,N_18035);
xor U22526 (N_22526,N_18870,N_19556);
and U22527 (N_22527,N_19140,N_17920);
and U22528 (N_22528,N_16542,N_16587);
xor U22529 (N_22529,N_15911,N_15440);
xor U22530 (N_22530,N_16425,N_18278);
nor U22531 (N_22531,N_18444,N_16595);
or U22532 (N_22532,N_15653,N_16481);
or U22533 (N_22533,N_18200,N_19610);
or U22534 (N_22534,N_18596,N_17767);
xor U22535 (N_22535,N_18823,N_19232);
nor U22536 (N_22536,N_17357,N_18109);
and U22537 (N_22537,N_15551,N_18939);
and U22538 (N_22538,N_19711,N_16149);
xnor U22539 (N_22539,N_19803,N_15461);
nor U22540 (N_22540,N_15826,N_18173);
xor U22541 (N_22541,N_19709,N_19578);
xor U22542 (N_22542,N_19644,N_17993);
nor U22543 (N_22543,N_18840,N_15020);
and U22544 (N_22544,N_18403,N_15750);
and U22545 (N_22545,N_19117,N_17027);
nand U22546 (N_22546,N_15968,N_15573);
or U22547 (N_22547,N_17942,N_18245);
or U22548 (N_22548,N_15296,N_15467);
nor U22549 (N_22549,N_16881,N_18087);
or U22550 (N_22550,N_18104,N_17413);
nor U22551 (N_22551,N_17156,N_17647);
nor U22552 (N_22552,N_17216,N_18118);
xnor U22553 (N_22553,N_17085,N_15687);
xnor U22554 (N_22554,N_17538,N_19202);
nand U22555 (N_22555,N_15499,N_16805);
xnor U22556 (N_22556,N_15545,N_16662);
nor U22557 (N_22557,N_18024,N_18317);
nand U22558 (N_22558,N_17386,N_15707);
and U22559 (N_22559,N_19176,N_19544);
or U22560 (N_22560,N_19569,N_18027);
and U22561 (N_22561,N_17494,N_15926);
and U22562 (N_22562,N_18578,N_19250);
nor U22563 (N_22563,N_15870,N_17521);
xor U22564 (N_22564,N_18227,N_15586);
or U22565 (N_22565,N_19969,N_16377);
and U22566 (N_22566,N_15740,N_18472);
nor U22567 (N_22567,N_15485,N_15147);
nand U22568 (N_22568,N_18259,N_17967);
nand U22569 (N_22569,N_17347,N_15634);
and U22570 (N_22570,N_17499,N_19735);
xnor U22571 (N_22571,N_16914,N_15833);
and U22572 (N_22572,N_17384,N_15640);
nand U22573 (N_22573,N_17207,N_15362);
nor U22574 (N_22574,N_15365,N_15190);
or U22575 (N_22575,N_17412,N_16425);
or U22576 (N_22576,N_18735,N_15556);
or U22577 (N_22577,N_15107,N_18938);
and U22578 (N_22578,N_16242,N_19231);
or U22579 (N_22579,N_16500,N_19362);
and U22580 (N_22580,N_19366,N_15960);
xor U22581 (N_22581,N_19032,N_15368);
nor U22582 (N_22582,N_18683,N_19279);
nand U22583 (N_22583,N_15461,N_19830);
xnor U22584 (N_22584,N_15965,N_19348);
xor U22585 (N_22585,N_18057,N_19760);
nor U22586 (N_22586,N_16189,N_18760);
xor U22587 (N_22587,N_17037,N_15376);
or U22588 (N_22588,N_18929,N_16493);
xnor U22589 (N_22589,N_15808,N_17255);
or U22590 (N_22590,N_18763,N_17508);
xnor U22591 (N_22591,N_19971,N_15522);
nand U22592 (N_22592,N_17909,N_15356);
and U22593 (N_22593,N_17319,N_16062);
and U22594 (N_22594,N_17254,N_19411);
nor U22595 (N_22595,N_16794,N_19015);
or U22596 (N_22596,N_17619,N_17291);
nand U22597 (N_22597,N_19427,N_19859);
xnor U22598 (N_22598,N_16278,N_16422);
xnor U22599 (N_22599,N_19572,N_17435);
nand U22600 (N_22600,N_16264,N_18389);
nand U22601 (N_22601,N_19996,N_16128);
nor U22602 (N_22602,N_18392,N_17556);
and U22603 (N_22603,N_18789,N_18177);
nand U22604 (N_22604,N_18606,N_17518);
nand U22605 (N_22605,N_19032,N_16404);
or U22606 (N_22606,N_15106,N_18794);
or U22607 (N_22607,N_15176,N_19951);
or U22608 (N_22608,N_15675,N_16425);
or U22609 (N_22609,N_17939,N_16907);
nor U22610 (N_22610,N_16728,N_17507);
and U22611 (N_22611,N_19112,N_19423);
or U22612 (N_22612,N_19773,N_16203);
xor U22613 (N_22613,N_17074,N_18838);
nor U22614 (N_22614,N_15118,N_18635);
or U22615 (N_22615,N_15463,N_19223);
nor U22616 (N_22616,N_17804,N_15227);
or U22617 (N_22617,N_15790,N_18802);
and U22618 (N_22618,N_15464,N_17774);
or U22619 (N_22619,N_17546,N_18585);
and U22620 (N_22620,N_19203,N_16048);
nand U22621 (N_22621,N_17710,N_18360);
xor U22622 (N_22622,N_19663,N_18615);
or U22623 (N_22623,N_18290,N_19134);
nand U22624 (N_22624,N_15087,N_18062);
xnor U22625 (N_22625,N_16803,N_17179);
or U22626 (N_22626,N_19766,N_17663);
xor U22627 (N_22627,N_19461,N_18971);
nor U22628 (N_22628,N_18899,N_17528);
and U22629 (N_22629,N_16220,N_17942);
or U22630 (N_22630,N_18190,N_18597);
xnor U22631 (N_22631,N_19386,N_18923);
nand U22632 (N_22632,N_19786,N_18881);
or U22633 (N_22633,N_18380,N_15744);
and U22634 (N_22634,N_16538,N_18337);
and U22635 (N_22635,N_16982,N_19622);
or U22636 (N_22636,N_17987,N_18712);
xnor U22637 (N_22637,N_18908,N_18669);
nor U22638 (N_22638,N_15067,N_16446);
nand U22639 (N_22639,N_15464,N_17569);
and U22640 (N_22640,N_18707,N_18722);
xor U22641 (N_22641,N_19624,N_15516);
and U22642 (N_22642,N_18029,N_19127);
or U22643 (N_22643,N_18077,N_18862);
and U22644 (N_22644,N_18222,N_17723);
nand U22645 (N_22645,N_16153,N_19314);
xnor U22646 (N_22646,N_16751,N_16784);
or U22647 (N_22647,N_16452,N_16603);
nand U22648 (N_22648,N_19436,N_17403);
and U22649 (N_22649,N_17186,N_16315);
nor U22650 (N_22650,N_16233,N_19305);
xnor U22651 (N_22651,N_19877,N_19596);
and U22652 (N_22652,N_15708,N_17475);
or U22653 (N_22653,N_19430,N_18739);
nor U22654 (N_22654,N_17238,N_16304);
nand U22655 (N_22655,N_16508,N_16973);
nand U22656 (N_22656,N_15404,N_17055);
xor U22657 (N_22657,N_18635,N_17606);
xor U22658 (N_22658,N_16058,N_15413);
or U22659 (N_22659,N_15476,N_15414);
nand U22660 (N_22660,N_19205,N_19843);
or U22661 (N_22661,N_15319,N_17089);
nand U22662 (N_22662,N_15096,N_19321);
and U22663 (N_22663,N_16326,N_15410);
nand U22664 (N_22664,N_18585,N_19154);
and U22665 (N_22665,N_19781,N_16161);
or U22666 (N_22666,N_19341,N_15443);
xnor U22667 (N_22667,N_15083,N_18180);
nand U22668 (N_22668,N_16819,N_16256);
and U22669 (N_22669,N_19785,N_19520);
xor U22670 (N_22670,N_19279,N_19082);
and U22671 (N_22671,N_15888,N_17874);
or U22672 (N_22672,N_19458,N_19449);
or U22673 (N_22673,N_15041,N_16432);
nor U22674 (N_22674,N_17125,N_16148);
xnor U22675 (N_22675,N_16751,N_18427);
nor U22676 (N_22676,N_19047,N_16201);
xor U22677 (N_22677,N_19543,N_19146);
or U22678 (N_22678,N_19816,N_16322);
xor U22679 (N_22679,N_15359,N_15724);
xor U22680 (N_22680,N_19160,N_16633);
or U22681 (N_22681,N_18948,N_16932);
xor U22682 (N_22682,N_16646,N_18363);
xnor U22683 (N_22683,N_15164,N_15223);
or U22684 (N_22684,N_17167,N_16562);
xor U22685 (N_22685,N_19776,N_15268);
nand U22686 (N_22686,N_16965,N_16274);
nand U22687 (N_22687,N_18598,N_19747);
and U22688 (N_22688,N_19245,N_17959);
nand U22689 (N_22689,N_15732,N_16965);
nor U22690 (N_22690,N_15339,N_19441);
and U22691 (N_22691,N_16852,N_17079);
or U22692 (N_22692,N_15798,N_17550);
and U22693 (N_22693,N_19861,N_17452);
or U22694 (N_22694,N_16686,N_15720);
nand U22695 (N_22695,N_19384,N_18810);
or U22696 (N_22696,N_18956,N_15826);
nand U22697 (N_22697,N_17097,N_15591);
nand U22698 (N_22698,N_15923,N_17236);
xor U22699 (N_22699,N_15988,N_17580);
nand U22700 (N_22700,N_18443,N_17287);
or U22701 (N_22701,N_18470,N_15841);
nand U22702 (N_22702,N_16632,N_15305);
nor U22703 (N_22703,N_19950,N_18555);
and U22704 (N_22704,N_18040,N_19805);
nand U22705 (N_22705,N_19110,N_19114);
nand U22706 (N_22706,N_15481,N_15803);
or U22707 (N_22707,N_18122,N_15193);
xnor U22708 (N_22708,N_16078,N_15569);
and U22709 (N_22709,N_17899,N_16401);
and U22710 (N_22710,N_17024,N_18737);
xnor U22711 (N_22711,N_15727,N_15484);
and U22712 (N_22712,N_18125,N_15919);
and U22713 (N_22713,N_18887,N_16234);
xnor U22714 (N_22714,N_17170,N_19507);
or U22715 (N_22715,N_17463,N_15287);
nor U22716 (N_22716,N_17219,N_18720);
and U22717 (N_22717,N_19789,N_17788);
or U22718 (N_22718,N_19933,N_17394);
nand U22719 (N_22719,N_16355,N_18295);
xnor U22720 (N_22720,N_18597,N_15661);
and U22721 (N_22721,N_18994,N_17947);
nor U22722 (N_22722,N_18529,N_16856);
xor U22723 (N_22723,N_16030,N_19072);
nor U22724 (N_22724,N_15844,N_18625);
nand U22725 (N_22725,N_19267,N_17116);
or U22726 (N_22726,N_15269,N_17240);
or U22727 (N_22727,N_18233,N_18025);
and U22728 (N_22728,N_17479,N_15371);
xor U22729 (N_22729,N_18308,N_19516);
xnor U22730 (N_22730,N_17121,N_15372);
nor U22731 (N_22731,N_16539,N_19878);
or U22732 (N_22732,N_18073,N_18193);
nand U22733 (N_22733,N_17425,N_16793);
or U22734 (N_22734,N_18801,N_17765);
or U22735 (N_22735,N_16671,N_18366);
nor U22736 (N_22736,N_19179,N_18391);
or U22737 (N_22737,N_16556,N_18559);
nand U22738 (N_22738,N_17205,N_16620);
nand U22739 (N_22739,N_19061,N_19570);
and U22740 (N_22740,N_19804,N_19818);
nand U22741 (N_22741,N_15021,N_15707);
nand U22742 (N_22742,N_19581,N_17672);
and U22743 (N_22743,N_15517,N_17126);
xor U22744 (N_22744,N_16543,N_16741);
and U22745 (N_22745,N_15747,N_18217);
nand U22746 (N_22746,N_16641,N_16091);
xor U22747 (N_22747,N_15576,N_19137);
and U22748 (N_22748,N_15217,N_16079);
nand U22749 (N_22749,N_19443,N_19790);
nand U22750 (N_22750,N_18048,N_18267);
nor U22751 (N_22751,N_19787,N_18244);
nor U22752 (N_22752,N_17159,N_19131);
nand U22753 (N_22753,N_18539,N_16647);
nor U22754 (N_22754,N_17088,N_16471);
xnor U22755 (N_22755,N_15608,N_15604);
nor U22756 (N_22756,N_17843,N_18729);
and U22757 (N_22757,N_19728,N_15298);
xor U22758 (N_22758,N_17170,N_15773);
xnor U22759 (N_22759,N_16323,N_18718);
xor U22760 (N_22760,N_17207,N_17122);
xnor U22761 (N_22761,N_17949,N_18331);
nand U22762 (N_22762,N_17703,N_17585);
and U22763 (N_22763,N_15912,N_17390);
or U22764 (N_22764,N_17851,N_19718);
and U22765 (N_22765,N_17530,N_19563);
nand U22766 (N_22766,N_17333,N_15666);
xnor U22767 (N_22767,N_16915,N_19026);
and U22768 (N_22768,N_16044,N_15712);
nor U22769 (N_22769,N_19112,N_16874);
nor U22770 (N_22770,N_18841,N_19049);
xor U22771 (N_22771,N_18166,N_18698);
and U22772 (N_22772,N_15795,N_19539);
xnor U22773 (N_22773,N_18896,N_17636);
nor U22774 (N_22774,N_18769,N_16337);
and U22775 (N_22775,N_19383,N_19064);
nor U22776 (N_22776,N_15701,N_18572);
xnor U22777 (N_22777,N_16075,N_17382);
or U22778 (N_22778,N_19608,N_17887);
and U22779 (N_22779,N_19701,N_15019);
and U22780 (N_22780,N_19783,N_19336);
nand U22781 (N_22781,N_18029,N_18198);
or U22782 (N_22782,N_15719,N_15068);
or U22783 (N_22783,N_17871,N_18133);
or U22784 (N_22784,N_17472,N_17206);
nor U22785 (N_22785,N_19828,N_15152);
nand U22786 (N_22786,N_18371,N_18626);
and U22787 (N_22787,N_15892,N_18770);
or U22788 (N_22788,N_15618,N_19755);
or U22789 (N_22789,N_15916,N_18295);
or U22790 (N_22790,N_15977,N_17643);
nand U22791 (N_22791,N_18762,N_19138);
or U22792 (N_22792,N_17639,N_15037);
nand U22793 (N_22793,N_18828,N_18537);
or U22794 (N_22794,N_17024,N_16172);
nand U22795 (N_22795,N_15084,N_19521);
nor U22796 (N_22796,N_16498,N_15164);
or U22797 (N_22797,N_16729,N_19668);
and U22798 (N_22798,N_17609,N_16889);
xnor U22799 (N_22799,N_18081,N_17505);
nand U22800 (N_22800,N_18382,N_15970);
or U22801 (N_22801,N_18908,N_15242);
nor U22802 (N_22802,N_15779,N_16492);
xor U22803 (N_22803,N_17563,N_19589);
and U22804 (N_22804,N_15699,N_15949);
nand U22805 (N_22805,N_16138,N_16508);
nor U22806 (N_22806,N_16006,N_18185);
or U22807 (N_22807,N_18012,N_15764);
or U22808 (N_22808,N_16344,N_19186);
xor U22809 (N_22809,N_19218,N_15283);
nor U22810 (N_22810,N_17884,N_15079);
nand U22811 (N_22811,N_17687,N_17319);
xnor U22812 (N_22812,N_15186,N_16147);
or U22813 (N_22813,N_15830,N_15193);
nor U22814 (N_22814,N_17349,N_16734);
and U22815 (N_22815,N_16248,N_19003);
xnor U22816 (N_22816,N_17038,N_18633);
nor U22817 (N_22817,N_16386,N_19385);
nor U22818 (N_22818,N_19975,N_16728);
xor U22819 (N_22819,N_18762,N_16772);
xor U22820 (N_22820,N_16991,N_17604);
xnor U22821 (N_22821,N_18434,N_19243);
and U22822 (N_22822,N_17519,N_19116);
xnor U22823 (N_22823,N_19027,N_19930);
xnor U22824 (N_22824,N_17577,N_17116);
nand U22825 (N_22825,N_15579,N_19923);
nor U22826 (N_22826,N_18226,N_17858);
or U22827 (N_22827,N_15186,N_15486);
nor U22828 (N_22828,N_16783,N_19112);
xnor U22829 (N_22829,N_19529,N_15347);
or U22830 (N_22830,N_18017,N_16607);
or U22831 (N_22831,N_17238,N_15901);
nand U22832 (N_22832,N_15525,N_15815);
nand U22833 (N_22833,N_19180,N_19134);
nor U22834 (N_22834,N_15846,N_19424);
nand U22835 (N_22835,N_18110,N_18340);
and U22836 (N_22836,N_16452,N_19876);
and U22837 (N_22837,N_18349,N_16715);
or U22838 (N_22838,N_19584,N_15436);
nand U22839 (N_22839,N_19569,N_16425);
or U22840 (N_22840,N_19741,N_19516);
and U22841 (N_22841,N_16935,N_17133);
and U22842 (N_22842,N_19809,N_19039);
or U22843 (N_22843,N_17343,N_18684);
or U22844 (N_22844,N_17466,N_19883);
nand U22845 (N_22845,N_16350,N_16057);
nor U22846 (N_22846,N_19897,N_18638);
and U22847 (N_22847,N_17720,N_15129);
or U22848 (N_22848,N_18915,N_18231);
and U22849 (N_22849,N_19778,N_17502);
or U22850 (N_22850,N_19360,N_15638);
nor U22851 (N_22851,N_19340,N_17071);
nor U22852 (N_22852,N_19714,N_19779);
nand U22853 (N_22853,N_17764,N_15565);
nand U22854 (N_22854,N_19858,N_15769);
and U22855 (N_22855,N_16770,N_16474);
and U22856 (N_22856,N_17959,N_18731);
xnor U22857 (N_22857,N_17431,N_18884);
xnor U22858 (N_22858,N_16883,N_15551);
nand U22859 (N_22859,N_17685,N_18762);
nand U22860 (N_22860,N_15167,N_18592);
nand U22861 (N_22861,N_18146,N_15055);
nand U22862 (N_22862,N_15985,N_15878);
nor U22863 (N_22863,N_15987,N_19016);
and U22864 (N_22864,N_16134,N_16558);
xnor U22865 (N_22865,N_17016,N_18762);
and U22866 (N_22866,N_15020,N_16789);
and U22867 (N_22867,N_19505,N_16093);
or U22868 (N_22868,N_15895,N_15443);
nor U22869 (N_22869,N_17387,N_15042);
xor U22870 (N_22870,N_19206,N_19666);
or U22871 (N_22871,N_17227,N_19541);
xor U22872 (N_22872,N_19624,N_17906);
nor U22873 (N_22873,N_16628,N_18512);
nand U22874 (N_22874,N_19641,N_19298);
nand U22875 (N_22875,N_19939,N_15772);
nor U22876 (N_22876,N_15975,N_15660);
nor U22877 (N_22877,N_16775,N_17878);
or U22878 (N_22878,N_19524,N_17957);
and U22879 (N_22879,N_18000,N_18582);
nand U22880 (N_22880,N_15445,N_19500);
nand U22881 (N_22881,N_19362,N_15056);
and U22882 (N_22882,N_19165,N_15396);
nor U22883 (N_22883,N_16049,N_18042);
xor U22884 (N_22884,N_15808,N_17356);
or U22885 (N_22885,N_15192,N_16638);
nand U22886 (N_22886,N_18404,N_18622);
or U22887 (N_22887,N_18633,N_15807);
xor U22888 (N_22888,N_18790,N_15235);
and U22889 (N_22889,N_15540,N_18948);
nor U22890 (N_22890,N_17113,N_19852);
and U22891 (N_22891,N_19559,N_18774);
and U22892 (N_22892,N_16340,N_17826);
nand U22893 (N_22893,N_18215,N_16061);
or U22894 (N_22894,N_17240,N_18016);
xnor U22895 (N_22895,N_16082,N_17912);
xnor U22896 (N_22896,N_15633,N_19962);
nor U22897 (N_22897,N_19865,N_19066);
nand U22898 (N_22898,N_17519,N_16183);
nor U22899 (N_22899,N_16130,N_18621);
nand U22900 (N_22900,N_17970,N_15366);
and U22901 (N_22901,N_16590,N_19416);
and U22902 (N_22902,N_19656,N_18460);
and U22903 (N_22903,N_15234,N_18196);
nand U22904 (N_22904,N_19837,N_18409);
or U22905 (N_22905,N_17473,N_16119);
and U22906 (N_22906,N_16879,N_15894);
and U22907 (N_22907,N_19147,N_16282);
xnor U22908 (N_22908,N_15447,N_17275);
and U22909 (N_22909,N_15139,N_16377);
nor U22910 (N_22910,N_19361,N_15964);
nor U22911 (N_22911,N_18671,N_15161);
xnor U22912 (N_22912,N_19581,N_17392);
nor U22913 (N_22913,N_17646,N_15502);
and U22914 (N_22914,N_17958,N_15121);
or U22915 (N_22915,N_18367,N_17761);
nor U22916 (N_22916,N_16807,N_15936);
xor U22917 (N_22917,N_16302,N_18023);
and U22918 (N_22918,N_17688,N_16366);
xor U22919 (N_22919,N_15712,N_15365);
or U22920 (N_22920,N_16223,N_16648);
nor U22921 (N_22921,N_18573,N_15540);
or U22922 (N_22922,N_18007,N_15074);
nand U22923 (N_22923,N_17016,N_19732);
xnor U22924 (N_22924,N_18484,N_18299);
and U22925 (N_22925,N_18677,N_15725);
nor U22926 (N_22926,N_18012,N_19341);
nor U22927 (N_22927,N_18394,N_18701);
or U22928 (N_22928,N_16060,N_17837);
xnor U22929 (N_22929,N_15801,N_17938);
or U22930 (N_22930,N_15119,N_15629);
and U22931 (N_22931,N_18604,N_16618);
xor U22932 (N_22932,N_17820,N_16446);
xor U22933 (N_22933,N_15602,N_16008);
nor U22934 (N_22934,N_16641,N_15532);
and U22935 (N_22935,N_17892,N_18205);
and U22936 (N_22936,N_19305,N_19570);
nor U22937 (N_22937,N_16774,N_16231);
or U22938 (N_22938,N_19764,N_18553);
and U22939 (N_22939,N_15755,N_18659);
and U22940 (N_22940,N_16281,N_18358);
xnor U22941 (N_22941,N_15324,N_19543);
and U22942 (N_22942,N_15403,N_15186);
or U22943 (N_22943,N_15244,N_17393);
or U22944 (N_22944,N_18879,N_16746);
or U22945 (N_22945,N_17735,N_17311);
or U22946 (N_22946,N_19491,N_19048);
xor U22947 (N_22947,N_17363,N_19758);
or U22948 (N_22948,N_15429,N_18219);
xor U22949 (N_22949,N_18513,N_17285);
xor U22950 (N_22950,N_15626,N_17908);
or U22951 (N_22951,N_19419,N_15648);
nor U22952 (N_22952,N_18589,N_19452);
nor U22953 (N_22953,N_17546,N_15532);
nor U22954 (N_22954,N_15692,N_17712);
or U22955 (N_22955,N_19675,N_15347);
nor U22956 (N_22956,N_19225,N_18591);
nor U22957 (N_22957,N_16176,N_18033);
nand U22958 (N_22958,N_15948,N_17467);
xor U22959 (N_22959,N_16434,N_19573);
and U22960 (N_22960,N_16159,N_17999);
or U22961 (N_22961,N_15070,N_19116);
nor U22962 (N_22962,N_18217,N_17599);
nand U22963 (N_22963,N_18700,N_19965);
and U22964 (N_22964,N_17576,N_18730);
or U22965 (N_22965,N_18525,N_18938);
nor U22966 (N_22966,N_15828,N_17301);
nor U22967 (N_22967,N_17257,N_17715);
and U22968 (N_22968,N_16812,N_18636);
and U22969 (N_22969,N_19528,N_19326);
and U22970 (N_22970,N_17951,N_18374);
nand U22971 (N_22971,N_19096,N_17591);
or U22972 (N_22972,N_15874,N_17365);
nor U22973 (N_22973,N_19525,N_16570);
nand U22974 (N_22974,N_17259,N_16649);
or U22975 (N_22975,N_15876,N_18792);
and U22976 (N_22976,N_17347,N_19132);
nand U22977 (N_22977,N_17034,N_17945);
or U22978 (N_22978,N_16142,N_15412);
nand U22979 (N_22979,N_15915,N_17855);
and U22980 (N_22980,N_19984,N_18264);
nand U22981 (N_22981,N_19921,N_15565);
xor U22982 (N_22982,N_19898,N_15066);
nor U22983 (N_22983,N_17334,N_17765);
or U22984 (N_22984,N_18705,N_19527);
xnor U22985 (N_22985,N_17371,N_16358);
and U22986 (N_22986,N_19286,N_19539);
or U22987 (N_22987,N_19416,N_17650);
nor U22988 (N_22988,N_15255,N_17047);
or U22989 (N_22989,N_19032,N_16323);
or U22990 (N_22990,N_17068,N_18330);
xnor U22991 (N_22991,N_15407,N_17147);
nand U22992 (N_22992,N_19882,N_15835);
or U22993 (N_22993,N_19735,N_17517);
nor U22994 (N_22994,N_15011,N_17302);
and U22995 (N_22995,N_15289,N_16047);
nand U22996 (N_22996,N_16176,N_19465);
or U22997 (N_22997,N_17805,N_19279);
xnor U22998 (N_22998,N_18153,N_19733);
nor U22999 (N_22999,N_17607,N_16715);
nor U23000 (N_23000,N_15083,N_16950);
or U23001 (N_23001,N_18775,N_15496);
nand U23002 (N_23002,N_18482,N_18594);
or U23003 (N_23003,N_19172,N_19173);
nand U23004 (N_23004,N_15376,N_17479);
or U23005 (N_23005,N_17397,N_18575);
nand U23006 (N_23006,N_17896,N_15154);
or U23007 (N_23007,N_16645,N_17354);
xor U23008 (N_23008,N_15922,N_17297);
nand U23009 (N_23009,N_15013,N_16867);
nor U23010 (N_23010,N_19130,N_15267);
and U23011 (N_23011,N_15351,N_17950);
and U23012 (N_23012,N_19327,N_15067);
or U23013 (N_23013,N_16755,N_16722);
or U23014 (N_23014,N_19162,N_17837);
nor U23015 (N_23015,N_19138,N_19757);
xor U23016 (N_23016,N_19310,N_19908);
nor U23017 (N_23017,N_18725,N_18038);
or U23018 (N_23018,N_18037,N_15106);
and U23019 (N_23019,N_16840,N_17315);
nand U23020 (N_23020,N_15829,N_17875);
and U23021 (N_23021,N_19591,N_16721);
or U23022 (N_23022,N_17279,N_15116);
xnor U23023 (N_23023,N_16244,N_18119);
nor U23024 (N_23024,N_15815,N_18184);
nor U23025 (N_23025,N_17475,N_18060);
or U23026 (N_23026,N_15188,N_17029);
or U23027 (N_23027,N_18426,N_17837);
and U23028 (N_23028,N_18886,N_18683);
nor U23029 (N_23029,N_19743,N_17600);
or U23030 (N_23030,N_18069,N_19889);
nand U23031 (N_23031,N_19111,N_19933);
nor U23032 (N_23032,N_17436,N_15186);
nand U23033 (N_23033,N_19050,N_18967);
nand U23034 (N_23034,N_19953,N_17674);
xnor U23035 (N_23035,N_18110,N_15899);
nor U23036 (N_23036,N_19506,N_17385);
xor U23037 (N_23037,N_17655,N_15292);
and U23038 (N_23038,N_15607,N_18457);
nor U23039 (N_23039,N_18634,N_16759);
xnor U23040 (N_23040,N_15052,N_19517);
and U23041 (N_23041,N_15582,N_17577);
nand U23042 (N_23042,N_15858,N_19432);
xnor U23043 (N_23043,N_16247,N_18871);
nor U23044 (N_23044,N_16037,N_15137);
or U23045 (N_23045,N_16121,N_18607);
and U23046 (N_23046,N_17748,N_15752);
or U23047 (N_23047,N_16051,N_17113);
or U23048 (N_23048,N_16390,N_19843);
nand U23049 (N_23049,N_17072,N_18357);
nand U23050 (N_23050,N_16592,N_15223);
and U23051 (N_23051,N_18997,N_19123);
nand U23052 (N_23052,N_18687,N_17421);
or U23053 (N_23053,N_18708,N_15292);
xor U23054 (N_23054,N_17724,N_15540);
nor U23055 (N_23055,N_19650,N_17613);
xor U23056 (N_23056,N_17658,N_19403);
xor U23057 (N_23057,N_19626,N_17027);
nand U23058 (N_23058,N_17841,N_18882);
nor U23059 (N_23059,N_15116,N_15220);
nor U23060 (N_23060,N_18395,N_19529);
nand U23061 (N_23061,N_19460,N_18291);
nand U23062 (N_23062,N_16271,N_15518);
xnor U23063 (N_23063,N_15324,N_18111);
and U23064 (N_23064,N_18823,N_16600);
and U23065 (N_23065,N_18771,N_15146);
nand U23066 (N_23066,N_15775,N_18552);
nand U23067 (N_23067,N_17521,N_18827);
xor U23068 (N_23068,N_15376,N_19046);
and U23069 (N_23069,N_17959,N_19848);
and U23070 (N_23070,N_18697,N_18825);
and U23071 (N_23071,N_19709,N_16100);
and U23072 (N_23072,N_15855,N_16294);
nor U23073 (N_23073,N_17544,N_18897);
xnor U23074 (N_23074,N_19945,N_15068);
xor U23075 (N_23075,N_17977,N_16386);
or U23076 (N_23076,N_17207,N_19579);
or U23077 (N_23077,N_19407,N_15079);
and U23078 (N_23078,N_17296,N_18277);
xor U23079 (N_23079,N_16226,N_18577);
xor U23080 (N_23080,N_18896,N_17223);
nor U23081 (N_23081,N_19292,N_17838);
or U23082 (N_23082,N_16068,N_17700);
xnor U23083 (N_23083,N_16095,N_16616);
xnor U23084 (N_23084,N_16162,N_17510);
or U23085 (N_23085,N_16380,N_19833);
nand U23086 (N_23086,N_16798,N_19429);
nand U23087 (N_23087,N_17161,N_17618);
xor U23088 (N_23088,N_16766,N_19107);
nand U23089 (N_23089,N_18737,N_16761);
and U23090 (N_23090,N_18263,N_18751);
xor U23091 (N_23091,N_18816,N_15722);
and U23092 (N_23092,N_19811,N_17169);
xnor U23093 (N_23093,N_16898,N_17372);
or U23094 (N_23094,N_18067,N_17453);
and U23095 (N_23095,N_19506,N_16737);
or U23096 (N_23096,N_19366,N_19272);
xnor U23097 (N_23097,N_16528,N_16320);
nor U23098 (N_23098,N_17715,N_16650);
xnor U23099 (N_23099,N_19240,N_17851);
nor U23100 (N_23100,N_18262,N_19430);
xor U23101 (N_23101,N_18031,N_17902);
nand U23102 (N_23102,N_19946,N_17574);
nor U23103 (N_23103,N_19871,N_17414);
xor U23104 (N_23104,N_17031,N_15496);
xor U23105 (N_23105,N_18714,N_18370);
and U23106 (N_23106,N_18758,N_16405);
or U23107 (N_23107,N_18476,N_16708);
nor U23108 (N_23108,N_18354,N_17104);
or U23109 (N_23109,N_15915,N_18894);
nor U23110 (N_23110,N_16162,N_17543);
xor U23111 (N_23111,N_15839,N_19124);
and U23112 (N_23112,N_17193,N_19223);
xor U23113 (N_23113,N_17100,N_15222);
xnor U23114 (N_23114,N_18894,N_15024);
or U23115 (N_23115,N_16883,N_17308);
nor U23116 (N_23116,N_16274,N_16203);
and U23117 (N_23117,N_18111,N_15520);
nand U23118 (N_23118,N_18610,N_16477);
or U23119 (N_23119,N_17529,N_17132);
and U23120 (N_23120,N_19970,N_15210);
and U23121 (N_23121,N_17163,N_16196);
xnor U23122 (N_23122,N_16660,N_15730);
and U23123 (N_23123,N_15198,N_16405);
nand U23124 (N_23124,N_16740,N_18947);
or U23125 (N_23125,N_19425,N_18174);
nand U23126 (N_23126,N_16501,N_16728);
nand U23127 (N_23127,N_19870,N_17814);
nor U23128 (N_23128,N_18376,N_16747);
xnor U23129 (N_23129,N_15151,N_16517);
and U23130 (N_23130,N_16648,N_15758);
xnor U23131 (N_23131,N_15089,N_17008);
nand U23132 (N_23132,N_15130,N_16661);
xor U23133 (N_23133,N_16423,N_17319);
nor U23134 (N_23134,N_18827,N_17200);
nand U23135 (N_23135,N_16174,N_15156);
or U23136 (N_23136,N_16280,N_19715);
and U23137 (N_23137,N_17645,N_15472);
nand U23138 (N_23138,N_19170,N_17932);
xnor U23139 (N_23139,N_17592,N_18556);
nor U23140 (N_23140,N_18288,N_19856);
xor U23141 (N_23141,N_17566,N_17967);
or U23142 (N_23142,N_15952,N_16230);
nor U23143 (N_23143,N_17015,N_17752);
or U23144 (N_23144,N_15864,N_18753);
and U23145 (N_23145,N_16215,N_18017);
nor U23146 (N_23146,N_15880,N_18768);
xnor U23147 (N_23147,N_19405,N_17045);
and U23148 (N_23148,N_16821,N_16191);
nand U23149 (N_23149,N_19719,N_17486);
or U23150 (N_23150,N_15601,N_15311);
nor U23151 (N_23151,N_19880,N_15603);
or U23152 (N_23152,N_16238,N_15262);
nor U23153 (N_23153,N_16945,N_19264);
and U23154 (N_23154,N_17726,N_16199);
nor U23155 (N_23155,N_16018,N_17294);
nand U23156 (N_23156,N_15878,N_19982);
or U23157 (N_23157,N_17288,N_16691);
nand U23158 (N_23158,N_17306,N_17122);
and U23159 (N_23159,N_18528,N_17630);
or U23160 (N_23160,N_19019,N_15949);
and U23161 (N_23161,N_18491,N_17605);
and U23162 (N_23162,N_16783,N_18061);
nor U23163 (N_23163,N_15175,N_15591);
nor U23164 (N_23164,N_16300,N_19934);
nor U23165 (N_23165,N_16221,N_18983);
and U23166 (N_23166,N_19544,N_16709);
nor U23167 (N_23167,N_17588,N_18450);
nor U23168 (N_23168,N_18484,N_19403);
nor U23169 (N_23169,N_16125,N_19858);
nor U23170 (N_23170,N_15387,N_15475);
and U23171 (N_23171,N_15044,N_19208);
and U23172 (N_23172,N_17853,N_19504);
or U23173 (N_23173,N_19462,N_17168);
nor U23174 (N_23174,N_17021,N_16348);
nand U23175 (N_23175,N_17516,N_16952);
and U23176 (N_23176,N_18992,N_19575);
or U23177 (N_23177,N_19306,N_17181);
nand U23178 (N_23178,N_17791,N_19858);
nand U23179 (N_23179,N_19281,N_17753);
nor U23180 (N_23180,N_17358,N_19214);
and U23181 (N_23181,N_19544,N_16076);
xnor U23182 (N_23182,N_19374,N_19689);
nor U23183 (N_23183,N_16561,N_19867);
nor U23184 (N_23184,N_17004,N_18259);
xnor U23185 (N_23185,N_16632,N_18447);
nand U23186 (N_23186,N_15027,N_19636);
nor U23187 (N_23187,N_19576,N_18903);
nor U23188 (N_23188,N_19915,N_15599);
xor U23189 (N_23189,N_16723,N_16042);
nor U23190 (N_23190,N_15942,N_17642);
or U23191 (N_23191,N_18346,N_17169);
and U23192 (N_23192,N_19868,N_18131);
nand U23193 (N_23193,N_19586,N_15819);
xor U23194 (N_23194,N_15832,N_16525);
or U23195 (N_23195,N_15326,N_15936);
or U23196 (N_23196,N_18705,N_16045);
xnor U23197 (N_23197,N_15683,N_19465);
and U23198 (N_23198,N_18748,N_18703);
nand U23199 (N_23199,N_16726,N_19722);
xnor U23200 (N_23200,N_18984,N_16769);
or U23201 (N_23201,N_17850,N_15128);
nand U23202 (N_23202,N_16895,N_16648);
xnor U23203 (N_23203,N_15407,N_18401);
nor U23204 (N_23204,N_19932,N_19936);
or U23205 (N_23205,N_16200,N_17854);
nor U23206 (N_23206,N_19554,N_18063);
xnor U23207 (N_23207,N_15580,N_17139);
nor U23208 (N_23208,N_18168,N_17900);
nand U23209 (N_23209,N_19116,N_19981);
and U23210 (N_23210,N_16125,N_16610);
and U23211 (N_23211,N_19344,N_17294);
xor U23212 (N_23212,N_15924,N_16572);
nand U23213 (N_23213,N_19041,N_19670);
or U23214 (N_23214,N_16879,N_19848);
nor U23215 (N_23215,N_15987,N_16162);
nor U23216 (N_23216,N_18741,N_15105);
xor U23217 (N_23217,N_18157,N_18646);
and U23218 (N_23218,N_18262,N_16863);
nand U23219 (N_23219,N_17719,N_17002);
or U23220 (N_23220,N_15848,N_16993);
and U23221 (N_23221,N_16486,N_19717);
nor U23222 (N_23222,N_15579,N_17899);
nor U23223 (N_23223,N_18267,N_18976);
xnor U23224 (N_23224,N_16599,N_16010);
nor U23225 (N_23225,N_17502,N_15130);
or U23226 (N_23226,N_18593,N_18985);
and U23227 (N_23227,N_18774,N_17234);
and U23228 (N_23228,N_17736,N_19056);
or U23229 (N_23229,N_15909,N_18615);
xnor U23230 (N_23230,N_17366,N_17942);
nand U23231 (N_23231,N_17114,N_19865);
xnor U23232 (N_23232,N_17711,N_18918);
xor U23233 (N_23233,N_18964,N_16612);
nor U23234 (N_23234,N_15801,N_19908);
nor U23235 (N_23235,N_18642,N_15507);
or U23236 (N_23236,N_15544,N_17091);
or U23237 (N_23237,N_19347,N_18552);
xnor U23238 (N_23238,N_18024,N_19830);
or U23239 (N_23239,N_15916,N_18717);
and U23240 (N_23240,N_19790,N_15136);
nand U23241 (N_23241,N_18566,N_18588);
nand U23242 (N_23242,N_17918,N_17313);
nor U23243 (N_23243,N_17847,N_19938);
or U23244 (N_23244,N_15286,N_16263);
or U23245 (N_23245,N_16639,N_16579);
xor U23246 (N_23246,N_15326,N_17975);
nand U23247 (N_23247,N_18074,N_16066);
nand U23248 (N_23248,N_17611,N_16212);
xor U23249 (N_23249,N_16301,N_17483);
xnor U23250 (N_23250,N_16164,N_19165);
nand U23251 (N_23251,N_17826,N_19839);
nand U23252 (N_23252,N_19508,N_16150);
and U23253 (N_23253,N_19362,N_19172);
xnor U23254 (N_23254,N_19363,N_19652);
nand U23255 (N_23255,N_16027,N_19099);
and U23256 (N_23256,N_17297,N_16733);
xor U23257 (N_23257,N_15066,N_17685);
xnor U23258 (N_23258,N_19214,N_15750);
and U23259 (N_23259,N_18693,N_19315);
xor U23260 (N_23260,N_17879,N_18526);
nor U23261 (N_23261,N_17373,N_16302);
or U23262 (N_23262,N_16529,N_17151);
nand U23263 (N_23263,N_16052,N_16200);
nor U23264 (N_23264,N_19761,N_19483);
nor U23265 (N_23265,N_18837,N_19953);
xnor U23266 (N_23266,N_18643,N_18240);
or U23267 (N_23267,N_15671,N_16768);
and U23268 (N_23268,N_17856,N_18510);
nor U23269 (N_23269,N_18413,N_16458);
xor U23270 (N_23270,N_17577,N_19281);
or U23271 (N_23271,N_17806,N_15054);
or U23272 (N_23272,N_18315,N_19979);
and U23273 (N_23273,N_17467,N_16074);
and U23274 (N_23274,N_16284,N_15341);
xnor U23275 (N_23275,N_17313,N_17712);
nand U23276 (N_23276,N_17305,N_15166);
nor U23277 (N_23277,N_16353,N_16424);
nand U23278 (N_23278,N_18700,N_17893);
nand U23279 (N_23279,N_18225,N_15712);
and U23280 (N_23280,N_19139,N_18265);
and U23281 (N_23281,N_16308,N_16291);
and U23282 (N_23282,N_18097,N_18855);
nand U23283 (N_23283,N_16580,N_16711);
or U23284 (N_23284,N_17608,N_18478);
nor U23285 (N_23285,N_17808,N_16546);
xnor U23286 (N_23286,N_18307,N_19942);
or U23287 (N_23287,N_15847,N_15792);
nand U23288 (N_23288,N_19094,N_18975);
nand U23289 (N_23289,N_16679,N_16033);
nor U23290 (N_23290,N_16029,N_16660);
or U23291 (N_23291,N_17718,N_16365);
xnor U23292 (N_23292,N_18576,N_15535);
xnor U23293 (N_23293,N_19294,N_18474);
nand U23294 (N_23294,N_15962,N_18772);
or U23295 (N_23295,N_18092,N_16271);
nor U23296 (N_23296,N_17890,N_18510);
or U23297 (N_23297,N_19997,N_15264);
xnor U23298 (N_23298,N_16737,N_19684);
or U23299 (N_23299,N_18752,N_19941);
and U23300 (N_23300,N_17474,N_17351);
xor U23301 (N_23301,N_18507,N_15462);
or U23302 (N_23302,N_16199,N_18355);
nor U23303 (N_23303,N_18358,N_15714);
or U23304 (N_23304,N_18388,N_16204);
nor U23305 (N_23305,N_18526,N_15803);
nor U23306 (N_23306,N_18503,N_17145);
and U23307 (N_23307,N_17594,N_15302);
nand U23308 (N_23308,N_16059,N_15751);
xnor U23309 (N_23309,N_16002,N_19221);
or U23310 (N_23310,N_15719,N_15664);
xor U23311 (N_23311,N_15491,N_16418);
nor U23312 (N_23312,N_16470,N_16057);
nor U23313 (N_23313,N_18956,N_16430);
nand U23314 (N_23314,N_18318,N_18143);
or U23315 (N_23315,N_19530,N_16710);
nor U23316 (N_23316,N_19130,N_15644);
or U23317 (N_23317,N_16404,N_19382);
nor U23318 (N_23318,N_18418,N_18193);
xnor U23319 (N_23319,N_17279,N_15092);
nor U23320 (N_23320,N_19980,N_19853);
nor U23321 (N_23321,N_19483,N_19085);
or U23322 (N_23322,N_17646,N_16311);
nor U23323 (N_23323,N_19041,N_15599);
nand U23324 (N_23324,N_15552,N_17079);
or U23325 (N_23325,N_18123,N_19773);
and U23326 (N_23326,N_18314,N_15286);
xor U23327 (N_23327,N_16437,N_16079);
nor U23328 (N_23328,N_19167,N_15513);
or U23329 (N_23329,N_15486,N_18446);
nand U23330 (N_23330,N_17352,N_16604);
nor U23331 (N_23331,N_19624,N_18204);
xor U23332 (N_23332,N_15091,N_15314);
nor U23333 (N_23333,N_16720,N_15458);
xor U23334 (N_23334,N_18177,N_19746);
nor U23335 (N_23335,N_16673,N_18973);
nand U23336 (N_23336,N_19732,N_15009);
or U23337 (N_23337,N_17522,N_16105);
and U23338 (N_23338,N_16264,N_19840);
xor U23339 (N_23339,N_16060,N_15012);
nand U23340 (N_23340,N_18544,N_18176);
nand U23341 (N_23341,N_17430,N_16670);
or U23342 (N_23342,N_18588,N_19912);
xnor U23343 (N_23343,N_17397,N_16822);
or U23344 (N_23344,N_16048,N_16283);
nor U23345 (N_23345,N_17499,N_17386);
nand U23346 (N_23346,N_17278,N_17121);
nor U23347 (N_23347,N_18875,N_16577);
and U23348 (N_23348,N_17483,N_19321);
and U23349 (N_23349,N_18592,N_18803);
or U23350 (N_23350,N_17204,N_16369);
nor U23351 (N_23351,N_18838,N_16596);
xnor U23352 (N_23352,N_16202,N_19626);
nand U23353 (N_23353,N_15154,N_18672);
xor U23354 (N_23354,N_17064,N_18088);
nor U23355 (N_23355,N_17633,N_18781);
xnor U23356 (N_23356,N_19715,N_15677);
or U23357 (N_23357,N_16981,N_18595);
or U23358 (N_23358,N_17312,N_19324);
or U23359 (N_23359,N_19724,N_17252);
nand U23360 (N_23360,N_16494,N_18114);
nand U23361 (N_23361,N_19382,N_19050);
nor U23362 (N_23362,N_19962,N_17663);
or U23363 (N_23363,N_15941,N_16796);
and U23364 (N_23364,N_15814,N_16486);
nor U23365 (N_23365,N_18499,N_19641);
and U23366 (N_23366,N_15554,N_16768);
and U23367 (N_23367,N_17232,N_17277);
nor U23368 (N_23368,N_19595,N_15378);
or U23369 (N_23369,N_19893,N_15630);
xnor U23370 (N_23370,N_16125,N_17551);
or U23371 (N_23371,N_15386,N_16236);
nand U23372 (N_23372,N_18658,N_18871);
xnor U23373 (N_23373,N_18335,N_18343);
nor U23374 (N_23374,N_15858,N_18578);
nand U23375 (N_23375,N_16161,N_19312);
nand U23376 (N_23376,N_19518,N_16683);
or U23377 (N_23377,N_19153,N_17421);
xor U23378 (N_23378,N_18256,N_19164);
or U23379 (N_23379,N_16244,N_16945);
and U23380 (N_23380,N_19279,N_17327);
nor U23381 (N_23381,N_19508,N_17180);
or U23382 (N_23382,N_17213,N_19240);
and U23383 (N_23383,N_17210,N_15929);
nor U23384 (N_23384,N_19407,N_18741);
xor U23385 (N_23385,N_18479,N_19928);
or U23386 (N_23386,N_17099,N_19707);
nor U23387 (N_23387,N_15647,N_18308);
nand U23388 (N_23388,N_18122,N_16440);
and U23389 (N_23389,N_15199,N_17158);
xnor U23390 (N_23390,N_19136,N_17069);
nor U23391 (N_23391,N_16281,N_15189);
nand U23392 (N_23392,N_18032,N_18980);
nand U23393 (N_23393,N_16824,N_16179);
or U23394 (N_23394,N_19992,N_15576);
and U23395 (N_23395,N_15858,N_18711);
xnor U23396 (N_23396,N_18434,N_19635);
nor U23397 (N_23397,N_16558,N_15150);
xor U23398 (N_23398,N_15359,N_18046);
or U23399 (N_23399,N_16401,N_17702);
or U23400 (N_23400,N_17380,N_17812);
or U23401 (N_23401,N_19200,N_15291);
xnor U23402 (N_23402,N_19013,N_19151);
nor U23403 (N_23403,N_15020,N_18655);
nand U23404 (N_23404,N_15410,N_15222);
and U23405 (N_23405,N_19908,N_19095);
xnor U23406 (N_23406,N_15394,N_17553);
xor U23407 (N_23407,N_19443,N_15209);
nor U23408 (N_23408,N_19104,N_16885);
nor U23409 (N_23409,N_19125,N_17876);
xnor U23410 (N_23410,N_18903,N_18438);
xnor U23411 (N_23411,N_16886,N_17394);
or U23412 (N_23412,N_15801,N_17774);
or U23413 (N_23413,N_18144,N_16099);
and U23414 (N_23414,N_16140,N_19511);
nand U23415 (N_23415,N_15433,N_18508);
nor U23416 (N_23416,N_16831,N_19491);
xor U23417 (N_23417,N_18873,N_15394);
nor U23418 (N_23418,N_18906,N_17754);
nor U23419 (N_23419,N_15818,N_19914);
xor U23420 (N_23420,N_16376,N_19242);
nor U23421 (N_23421,N_18698,N_17830);
or U23422 (N_23422,N_18869,N_18707);
or U23423 (N_23423,N_16142,N_18993);
and U23424 (N_23424,N_15277,N_18336);
nand U23425 (N_23425,N_18113,N_17296);
or U23426 (N_23426,N_17697,N_16664);
or U23427 (N_23427,N_18294,N_15109);
nand U23428 (N_23428,N_16778,N_15450);
and U23429 (N_23429,N_15370,N_16512);
nand U23430 (N_23430,N_18608,N_15445);
nor U23431 (N_23431,N_15480,N_19347);
nor U23432 (N_23432,N_15922,N_17210);
xnor U23433 (N_23433,N_17433,N_17188);
nand U23434 (N_23434,N_16593,N_16088);
xor U23435 (N_23435,N_16126,N_15782);
xnor U23436 (N_23436,N_19092,N_17332);
xor U23437 (N_23437,N_18202,N_15261);
nor U23438 (N_23438,N_15661,N_15904);
nand U23439 (N_23439,N_16067,N_17901);
nand U23440 (N_23440,N_18590,N_17060);
and U23441 (N_23441,N_17184,N_15641);
and U23442 (N_23442,N_15379,N_16499);
and U23443 (N_23443,N_15599,N_16134);
or U23444 (N_23444,N_18780,N_19583);
nand U23445 (N_23445,N_17282,N_18978);
nand U23446 (N_23446,N_18029,N_19718);
or U23447 (N_23447,N_19678,N_18701);
or U23448 (N_23448,N_15605,N_17646);
nor U23449 (N_23449,N_15999,N_18929);
nand U23450 (N_23450,N_16007,N_16469);
or U23451 (N_23451,N_17779,N_17081);
xor U23452 (N_23452,N_19332,N_15480);
nand U23453 (N_23453,N_19716,N_19143);
nand U23454 (N_23454,N_19912,N_18613);
and U23455 (N_23455,N_17900,N_17452);
xnor U23456 (N_23456,N_15778,N_17891);
or U23457 (N_23457,N_17557,N_19459);
nand U23458 (N_23458,N_18601,N_15530);
nor U23459 (N_23459,N_18593,N_17883);
nor U23460 (N_23460,N_15186,N_17215);
xnor U23461 (N_23461,N_17732,N_18146);
nor U23462 (N_23462,N_16689,N_17445);
and U23463 (N_23463,N_16986,N_18848);
nand U23464 (N_23464,N_15242,N_16530);
and U23465 (N_23465,N_18211,N_16815);
and U23466 (N_23466,N_15758,N_18244);
nand U23467 (N_23467,N_18634,N_16702);
nor U23468 (N_23468,N_16799,N_17529);
xnor U23469 (N_23469,N_15056,N_15740);
nor U23470 (N_23470,N_18183,N_19450);
or U23471 (N_23471,N_18407,N_15612);
or U23472 (N_23472,N_16084,N_19680);
or U23473 (N_23473,N_17252,N_17036);
nand U23474 (N_23474,N_17002,N_17038);
nand U23475 (N_23475,N_18557,N_18372);
nand U23476 (N_23476,N_15645,N_15302);
xnor U23477 (N_23477,N_16299,N_19444);
or U23478 (N_23478,N_19933,N_17413);
nor U23479 (N_23479,N_18644,N_16213);
xor U23480 (N_23480,N_15008,N_17413);
nand U23481 (N_23481,N_16867,N_18502);
nand U23482 (N_23482,N_18310,N_15375);
nor U23483 (N_23483,N_18155,N_15324);
or U23484 (N_23484,N_18573,N_16022);
nor U23485 (N_23485,N_16200,N_18990);
or U23486 (N_23486,N_15161,N_15763);
nor U23487 (N_23487,N_15911,N_17181);
or U23488 (N_23488,N_16773,N_18790);
and U23489 (N_23489,N_19922,N_15629);
xor U23490 (N_23490,N_18659,N_16551);
xnor U23491 (N_23491,N_15551,N_19472);
xnor U23492 (N_23492,N_15362,N_15493);
or U23493 (N_23493,N_18237,N_15398);
or U23494 (N_23494,N_19752,N_17262);
nor U23495 (N_23495,N_19940,N_18351);
or U23496 (N_23496,N_16903,N_19654);
or U23497 (N_23497,N_17686,N_19584);
xnor U23498 (N_23498,N_19076,N_19464);
nand U23499 (N_23499,N_19037,N_19754);
nor U23500 (N_23500,N_18360,N_17878);
and U23501 (N_23501,N_19977,N_19937);
nor U23502 (N_23502,N_19874,N_18608);
nand U23503 (N_23503,N_15184,N_18023);
nor U23504 (N_23504,N_18524,N_17980);
or U23505 (N_23505,N_18900,N_16565);
xnor U23506 (N_23506,N_17923,N_19026);
xnor U23507 (N_23507,N_16688,N_15110);
or U23508 (N_23508,N_18991,N_17413);
or U23509 (N_23509,N_15782,N_15673);
or U23510 (N_23510,N_17304,N_17971);
or U23511 (N_23511,N_17052,N_19165);
nand U23512 (N_23512,N_17155,N_16714);
nand U23513 (N_23513,N_17583,N_17075);
and U23514 (N_23514,N_18858,N_15366);
or U23515 (N_23515,N_16190,N_17003);
nand U23516 (N_23516,N_16567,N_16110);
xor U23517 (N_23517,N_16484,N_19876);
and U23518 (N_23518,N_17392,N_17370);
xnor U23519 (N_23519,N_16861,N_17669);
xor U23520 (N_23520,N_16795,N_19537);
nor U23521 (N_23521,N_16167,N_18137);
nand U23522 (N_23522,N_17957,N_15218);
nand U23523 (N_23523,N_15406,N_19810);
and U23524 (N_23524,N_18041,N_18018);
or U23525 (N_23525,N_18742,N_17702);
or U23526 (N_23526,N_17889,N_17599);
and U23527 (N_23527,N_18892,N_16013);
xor U23528 (N_23528,N_19439,N_19094);
and U23529 (N_23529,N_19078,N_18865);
nor U23530 (N_23530,N_19865,N_17415);
and U23531 (N_23531,N_15752,N_16363);
xor U23532 (N_23532,N_18887,N_19992);
nand U23533 (N_23533,N_18395,N_15426);
or U23534 (N_23534,N_15824,N_19057);
and U23535 (N_23535,N_18250,N_15424);
or U23536 (N_23536,N_16526,N_15636);
and U23537 (N_23537,N_15544,N_19427);
xnor U23538 (N_23538,N_15892,N_19098);
xor U23539 (N_23539,N_16737,N_17603);
nor U23540 (N_23540,N_15228,N_19396);
and U23541 (N_23541,N_19606,N_15436);
nor U23542 (N_23542,N_18173,N_18017);
and U23543 (N_23543,N_17294,N_16099);
or U23544 (N_23544,N_18128,N_15807);
and U23545 (N_23545,N_19260,N_18747);
nand U23546 (N_23546,N_16130,N_19791);
nor U23547 (N_23547,N_15608,N_19902);
nand U23548 (N_23548,N_19044,N_18258);
nand U23549 (N_23549,N_17429,N_18252);
and U23550 (N_23550,N_18900,N_16725);
nand U23551 (N_23551,N_17357,N_19528);
and U23552 (N_23552,N_18558,N_18256);
nand U23553 (N_23553,N_16129,N_17826);
nand U23554 (N_23554,N_18366,N_17261);
nand U23555 (N_23555,N_17327,N_16202);
or U23556 (N_23556,N_17892,N_18636);
or U23557 (N_23557,N_18169,N_19330);
xor U23558 (N_23558,N_18079,N_18267);
or U23559 (N_23559,N_17336,N_15361);
and U23560 (N_23560,N_15374,N_16558);
xnor U23561 (N_23561,N_19891,N_17566);
nor U23562 (N_23562,N_17634,N_18177);
xnor U23563 (N_23563,N_18018,N_15723);
or U23564 (N_23564,N_15734,N_16979);
and U23565 (N_23565,N_17707,N_15010);
or U23566 (N_23566,N_19818,N_15393);
or U23567 (N_23567,N_16372,N_19850);
or U23568 (N_23568,N_16197,N_19087);
nor U23569 (N_23569,N_15555,N_15559);
or U23570 (N_23570,N_18500,N_17979);
or U23571 (N_23571,N_18209,N_19634);
or U23572 (N_23572,N_17886,N_18126);
nor U23573 (N_23573,N_15384,N_18406);
nor U23574 (N_23574,N_17302,N_16835);
or U23575 (N_23575,N_17459,N_19477);
xor U23576 (N_23576,N_19639,N_15823);
and U23577 (N_23577,N_17119,N_19874);
and U23578 (N_23578,N_16944,N_15761);
xor U23579 (N_23579,N_16399,N_18607);
or U23580 (N_23580,N_17924,N_18989);
and U23581 (N_23581,N_17380,N_15854);
nand U23582 (N_23582,N_19724,N_16682);
nor U23583 (N_23583,N_15760,N_18883);
xnor U23584 (N_23584,N_16642,N_18931);
nor U23585 (N_23585,N_17984,N_15113);
and U23586 (N_23586,N_16504,N_16694);
and U23587 (N_23587,N_15935,N_19828);
or U23588 (N_23588,N_19729,N_18775);
or U23589 (N_23589,N_15194,N_15093);
and U23590 (N_23590,N_16579,N_17463);
and U23591 (N_23591,N_18451,N_16398);
nand U23592 (N_23592,N_19785,N_18383);
and U23593 (N_23593,N_15091,N_15624);
or U23594 (N_23594,N_15033,N_18160);
nand U23595 (N_23595,N_17557,N_16869);
and U23596 (N_23596,N_17709,N_15699);
nor U23597 (N_23597,N_18597,N_18359);
and U23598 (N_23598,N_17103,N_16266);
nand U23599 (N_23599,N_17615,N_17252);
nor U23600 (N_23600,N_16283,N_17073);
or U23601 (N_23601,N_19198,N_19582);
nand U23602 (N_23602,N_15809,N_15091);
or U23603 (N_23603,N_16204,N_17312);
xor U23604 (N_23604,N_17014,N_17669);
nand U23605 (N_23605,N_19050,N_18085);
and U23606 (N_23606,N_19123,N_15180);
nand U23607 (N_23607,N_19800,N_19455);
xnor U23608 (N_23608,N_18557,N_15765);
nand U23609 (N_23609,N_18312,N_19959);
nand U23610 (N_23610,N_19433,N_15339);
nor U23611 (N_23611,N_17705,N_19222);
nand U23612 (N_23612,N_18062,N_16015);
and U23613 (N_23613,N_16472,N_16519);
xnor U23614 (N_23614,N_17045,N_15186);
xnor U23615 (N_23615,N_19271,N_18461);
nand U23616 (N_23616,N_16613,N_17941);
nand U23617 (N_23617,N_17292,N_16274);
and U23618 (N_23618,N_19167,N_18027);
nor U23619 (N_23619,N_15797,N_16886);
nand U23620 (N_23620,N_15041,N_19524);
xnor U23621 (N_23621,N_17438,N_15026);
and U23622 (N_23622,N_19733,N_16042);
nor U23623 (N_23623,N_15483,N_19875);
and U23624 (N_23624,N_15756,N_19062);
and U23625 (N_23625,N_16798,N_15811);
and U23626 (N_23626,N_16632,N_16101);
nor U23627 (N_23627,N_16211,N_15246);
and U23628 (N_23628,N_19336,N_19967);
and U23629 (N_23629,N_19032,N_16450);
and U23630 (N_23630,N_15842,N_15640);
nand U23631 (N_23631,N_18983,N_19543);
nand U23632 (N_23632,N_17879,N_18129);
nor U23633 (N_23633,N_18441,N_18251);
and U23634 (N_23634,N_15509,N_18868);
and U23635 (N_23635,N_15879,N_17954);
and U23636 (N_23636,N_15925,N_17221);
and U23637 (N_23637,N_17341,N_19009);
or U23638 (N_23638,N_18912,N_15724);
nand U23639 (N_23639,N_15655,N_17688);
xor U23640 (N_23640,N_18563,N_17743);
or U23641 (N_23641,N_15672,N_19218);
nand U23642 (N_23642,N_15282,N_17567);
and U23643 (N_23643,N_15262,N_17134);
nand U23644 (N_23644,N_16963,N_15274);
and U23645 (N_23645,N_15934,N_19951);
nor U23646 (N_23646,N_17915,N_18923);
and U23647 (N_23647,N_18928,N_17717);
nand U23648 (N_23648,N_19530,N_19225);
or U23649 (N_23649,N_16570,N_19610);
and U23650 (N_23650,N_18382,N_19275);
nand U23651 (N_23651,N_16332,N_19546);
or U23652 (N_23652,N_17224,N_17727);
nand U23653 (N_23653,N_16432,N_17839);
xor U23654 (N_23654,N_17739,N_19454);
and U23655 (N_23655,N_18897,N_18058);
or U23656 (N_23656,N_17995,N_19202);
or U23657 (N_23657,N_15521,N_15821);
nor U23658 (N_23658,N_17860,N_15957);
nand U23659 (N_23659,N_18554,N_17649);
and U23660 (N_23660,N_17046,N_18186);
nand U23661 (N_23661,N_17003,N_16297);
nand U23662 (N_23662,N_15675,N_15319);
nor U23663 (N_23663,N_16874,N_18169);
or U23664 (N_23664,N_16633,N_18646);
nand U23665 (N_23665,N_18772,N_16553);
xor U23666 (N_23666,N_15560,N_16609);
nand U23667 (N_23667,N_19123,N_19287);
nor U23668 (N_23668,N_19103,N_17173);
or U23669 (N_23669,N_19706,N_19791);
or U23670 (N_23670,N_17012,N_18059);
nor U23671 (N_23671,N_17963,N_16733);
xor U23672 (N_23672,N_18434,N_17732);
or U23673 (N_23673,N_16095,N_16128);
nor U23674 (N_23674,N_17625,N_18001);
nor U23675 (N_23675,N_19483,N_19563);
and U23676 (N_23676,N_19352,N_17252);
xnor U23677 (N_23677,N_16850,N_18420);
xnor U23678 (N_23678,N_17695,N_15739);
nand U23679 (N_23679,N_15938,N_15554);
nor U23680 (N_23680,N_17152,N_19703);
nor U23681 (N_23681,N_15019,N_15841);
xnor U23682 (N_23682,N_19630,N_18879);
or U23683 (N_23683,N_15694,N_17376);
and U23684 (N_23684,N_15240,N_17896);
xor U23685 (N_23685,N_19209,N_18810);
xor U23686 (N_23686,N_15321,N_17173);
or U23687 (N_23687,N_18123,N_19238);
xnor U23688 (N_23688,N_16201,N_19653);
nor U23689 (N_23689,N_19075,N_16522);
nand U23690 (N_23690,N_15990,N_16209);
xor U23691 (N_23691,N_16853,N_18894);
and U23692 (N_23692,N_19206,N_15185);
and U23693 (N_23693,N_15305,N_15207);
or U23694 (N_23694,N_16324,N_18035);
nor U23695 (N_23695,N_16776,N_18802);
nand U23696 (N_23696,N_16895,N_19944);
and U23697 (N_23697,N_18768,N_19470);
xor U23698 (N_23698,N_17355,N_18867);
or U23699 (N_23699,N_17361,N_15053);
or U23700 (N_23700,N_18026,N_17965);
nand U23701 (N_23701,N_16587,N_18557);
and U23702 (N_23702,N_15410,N_19183);
nor U23703 (N_23703,N_17004,N_19511);
and U23704 (N_23704,N_16111,N_19379);
nand U23705 (N_23705,N_19383,N_16481);
xnor U23706 (N_23706,N_19029,N_17248);
or U23707 (N_23707,N_16620,N_15107);
or U23708 (N_23708,N_19663,N_19105);
and U23709 (N_23709,N_15101,N_17871);
xnor U23710 (N_23710,N_17547,N_17209);
nor U23711 (N_23711,N_18407,N_17616);
nor U23712 (N_23712,N_18825,N_19195);
and U23713 (N_23713,N_16983,N_19416);
or U23714 (N_23714,N_18013,N_17269);
xor U23715 (N_23715,N_15706,N_15313);
xor U23716 (N_23716,N_18616,N_17987);
or U23717 (N_23717,N_18592,N_16958);
or U23718 (N_23718,N_19227,N_17175);
nor U23719 (N_23719,N_17642,N_15055);
or U23720 (N_23720,N_19663,N_19362);
or U23721 (N_23721,N_19188,N_18191);
nand U23722 (N_23722,N_19035,N_15411);
nor U23723 (N_23723,N_15330,N_15912);
or U23724 (N_23724,N_18802,N_16839);
xor U23725 (N_23725,N_18258,N_16915);
nor U23726 (N_23726,N_17517,N_19842);
nor U23727 (N_23727,N_19025,N_15133);
or U23728 (N_23728,N_17581,N_17125);
nor U23729 (N_23729,N_15069,N_16643);
xnor U23730 (N_23730,N_15023,N_17375);
and U23731 (N_23731,N_19698,N_15594);
nand U23732 (N_23732,N_18638,N_18392);
and U23733 (N_23733,N_17722,N_17392);
or U23734 (N_23734,N_15305,N_17210);
or U23735 (N_23735,N_19585,N_16975);
and U23736 (N_23736,N_16526,N_18930);
nor U23737 (N_23737,N_18186,N_19409);
xor U23738 (N_23738,N_19000,N_17705);
and U23739 (N_23739,N_17808,N_17606);
or U23740 (N_23740,N_18864,N_16613);
xnor U23741 (N_23741,N_19247,N_18880);
xor U23742 (N_23742,N_15836,N_15976);
nor U23743 (N_23743,N_18529,N_15582);
or U23744 (N_23744,N_18982,N_18682);
xnor U23745 (N_23745,N_16361,N_17007);
nand U23746 (N_23746,N_16689,N_16390);
nand U23747 (N_23747,N_15066,N_16927);
or U23748 (N_23748,N_17515,N_17357);
and U23749 (N_23749,N_15312,N_18202);
nor U23750 (N_23750,N_17797,N_15115);
and U23751 (N_23751,N_18321,N_17126);
nor U23752 (N_23752,N_15854,N_19727);
or U23753 (N_23753,N_17517,N_15493);
and U23754 (N_23754,N_18002,N_17004);
nor U23755 (N_23755,N_17961,N_17549);
nor U23756 (N_23756,N_18178,N_18142);
nand U23757 (N_23757,N_15341,N_19679);
or U23758 (N_23758,N_15667,N_19639);
nand U23759 (N_23759,N_15592,N_18402);
and U23760 (N_23760,N_16825,N_17723);
and U23761 (N_23761,N_18033,N_16772);
or U23762 (N_23762,N_19613,N_16759);
xor U23763 (N_23763,N_19402,N_15208);
nor U23764 (N_23764,N_17735,N_17272);
nor U23765 (N_23765,N_19908,N_15001);
xnor U23766 (N_23766,N_15735,N_15856);
xor U23767 (N_23767,N_19838,N_17004);
nor U23768 (N_23768,N_19006,N_18430);
xnor U23769 (N_23769,N_19539,N_17953);
or U23770 (N_23770,N_19059,N_15407);
nor U23771 (N_23771,N_15685,N_19499);
or U23772 (N_23772,N_17514,N_18892);
nand U23773 (N_23773,N_18623,N_17750);
nand U23774 (N_23774,N_16351,N_15962);
and U23775 (N_23775,N_18957,N_19666);
and U23776 (N_23776,N_19784,N_16901);
and U23777 (N_23777,N_18654,N_17445);
nand U23778 (N_23778,N_16221,N_15397);
xor U23779 (N_23779,N_19883,N_18003);
or U23780 (N_23780,N_17111,N_18037);
nand U23781 (N_23781,N_17437,N_16370);
nand U23782 (N_23782,N_17860,N_18363);
nor U23783 (N_23783,N_16141,N_19358);
and U23784 (N_23784,N_15526,N_18678);
and U23785 (N_23785,N_19140,N_16223);
nor U23786 (N_23786,N_17541,N_19820);
nor U23787 (N_23787,N_19232,N_18479);
nand U23788 (N_23788,N_17958,N_18807);
nand U23789 (N_23789,N_18354,N_19898);
nor U23790 (N_23790,N_16496,N_17999);
nor U23791 (N_23791,N_19994,N_18808);
or U23792 (N_23792,N_15399,N_16996);
xor U23793 (N_23793,N_15663,N_19878);
xor U23794 (N_23794,N_19302,N_17172);
nor U23795 (N_23795,N_17792,N_18989);
or U23796 (N_23796,N_19098,N_17425);
nand U23797 (N_23797,N_19274,N_17919);
xnor U23798 (N_23798,N_19496,N_18986);
nor U23799 (N_23799,N_18043,N_19721);
nand U23800 (N_23800,N_15931,N_17711);
nand U23801 (N_23801,N_15842,N_16017);
or U23802 (N_23802,N_16285,N_18474);
and U23803 (N_23803,N_15510,N_15113);
or U23804 (N_23804,N_16072,N_16530);
nor U23805 (N_23805,N_19839,N_16724);
xnor U23806 (N_23806,N_18719,N_18346);
or U23807 (N_23807,N_17047,N_19804);
or U23808 (N_23808,N_16363,N_17794);
nor U23809 (N_23809,N_18061,N_16836);
and U23810 (N_23810,N_18572,N_19842);
nand U23811 (N_23811,N_19568,N_16374);
nor U23812 (N_23812,N_19395,N_18538);
nand U23813 (N_23813,N_19696,N_19379);
nor U23814 (N_23814,N_16725,N_17293);
nand U23815 (N_23815,N_16314,N_15104);
xnor U23816 (N_23816,N_15720,N_16859);
and U23817 (N_23817,N_18331,N_18541);
nor U23818 (N_23818,N_15119,N_18062);
and U23819 (N_23819,N_16865,N_16992);
nor U23820 (N_23820,N_16970,N_19262);
nor U23821 (N_23821,N_16287,N_15505);
nand U23822 (N_23822,N_15259,N_19765);
nor U23823 (N_23823,N_19982,N_19093);
xnor U23824 (N_23824,N_19937,N_17199);
xor U23825 (N_23825,N_16142,N_19489);
or U23826 (N_23826,N_17234,N_19909);
xnor U23827 (N_23827,N_17940,N_17005);
or U23828 (N_23828,N_19453,N_17977);
xor U23829 (N_23829,N_19809,N_16091);
and U23830 (N_23830,N_18134,N_16222);
or U23831 (N_23831,N_16162,N_19628);
nand U23832 (N_23832,N_16497,N_18946);
nand U23833 (N_23833,N_17443,N_18320);
xor U23834 (N_23834,N_17307,N_18256);
xnor U23835 (N_23835,N_16121,N_19815);
or U23836 (N_23836,N_16335,N_16462);
and U23837 (N_23837,N_18501,N_17417);
nor U23838 (N_23838,N_15848,N_17282);
or U23839 (N_23839,N_15322,N_19117);
xnor U23840 (N_23840,N_18847,N_16047);
or U23841 (N_23841,N_18983,N_18926);
nor U23842 (N_23842,N_17458,N_17418);
nand U23843 (N_23843,N_16308,N_15699);
xnor U23844 (N_23844,N_18121,N_19571);
and U23845 (N_23845,N_19681,N_18317);
nor U23846 (N_23846,N_16891,N_15511);
nor U23847 (N_23847,N_15948,N_19137);
xor U23848 (N_23848,N_16994,N_18923);
and U23849 (N_23849,N_17054,N_17748);
xor U23850 (N_23850,N_15968,N_19938);
nand U23851 (N_23851,N_16244,N_18963);
and U23852 (N_23852,N_17350,N_16869);
and U23853 (N_23853,N_18266,N_16997);
nand U23854 (N_23854,N_19191,N_19001);
nand U23855 (N_23855,N_17173,N_19873);
xor U23856 (N_23856,N_17873,N_15818);
xor U23857 (N_23857,N_17769,N_15039);
nand U23858 (N_23858,N_18844,N_15661);
or U23859 (N_23859,N_15818,N_17225);
nand U23860 (N_23860,N_19484,N_19322);
and U23861 (N_23861,N_17852,N_16912);
and U23862 (N_23862,N_18639,N_19386);
nor U23863 (N_23863,N_19819,N_18645);
nand U23864 (N_23864,N_17340,N_19229);
and U23865 (N_23865,N_19749,N_16655);
xnor U23866 (N_23866,N_17168,N_18869);
or U23867 (N_23867,N_19589,N_16980);
nor U23868 (N_23868,N_15643,N_17973);
nor U23869 (N_23869,N_16040,N_17213);
xnor U23870 (N_23870,N_18090,N_15886);
nor U23871 (N_23871,N_16932,N_16809);
or U23872 (N_23872,N_16974,N_15871);
nand U23873 (N_23873,N_18329,N_17222);
or U23874 (N_23874,N_15596,N_17356);
and U23875 (N_23875,N_18987,N_19147);
or U23876 (N_23876,N_18281,N_19131);
or U23877 (N_23877,N_17322,N_19134);
xnor U23878 (N_23878,N_19962,N_15263);
nand U23879 (N_23879,N_18569,N_19091);
nor U23880 (N_23880,N_18632,N_17214);
nand U23881 (N_23881,N_19976,N_16641);
xnor U23882 (N_23882,N_19183,N_19999);
xnor U23883 (N_23883,N_19146,N_19039);
xor U23884 (N_23884,N_15400,N_15375);
nor U23885 (N_23885,N_19776,N_15383);
or U23886 (N_23886,N_19966,N_19382);
nor U23887 (N_23887,N_16239,N_19837);
and U23888 (N_23888,N_16613,N_17864);
or U23889 (N_23889,N_19661,N_17339);
and U23890 (N_23890,N_16944,N_19911);
and U23891 (N_23891,N_17927,N_17805);
nor U23892 (N_23892,N_17444,N_17982);
nand U23893 (N_23893,N_15695,N_16938);
and U23894 (N_23894,N_16865,N_18602);
or U23895 (N_23895,N_15609,N_16316);
and U23896 (N_23896,N_18838,N_18698);
xor U23897 (N_23897,N_17597,N_17334);
xnor U23898 (N_23898,N_19296,N_15956);
xnor U23899 (N_23899,N_18004,N_15043);
nand U23900 (N_23900,N_15153,N_19874);
and U23901 (N_23901,N_18654,N_17199);
nor U23902 (N_23902,N_16775,N_16149);
nand U23903 (N_23903,N_18896,N_15599);
and U23904 (N_23904,N_18546,N_18459);
and U23905 (N_23905,N_15038,N_19350);
or U23906 (N_23906,N_15687,N_15030);
and U23907 (N_23907,N_15634,N_19081);
xnor U23908 (N_23908,N_16545,N_16342);
nand U23909 (N_23909,N_18026,N_15590);
or U23910 (N_23910,N_17351,N_19468);
xor U23911 (N_23911,N_19954,N_19581);
or U23912 (N_23912,N_19864,N_17430);
xnor U23913 (N_23913,N_17665,N_16845);
nand U23914 (N_23914,N_15720,N_18651);
and U23915 (N_23915,N_15151,N_19278);
and U23916 (N_23916,N_18215,N_19926);
xor U23917 (N_23917,N_19671,N_16771);
nand U23918 (N_23918,N_16645,N_18146);
nor U23919 (N_23919,N_17972,N_17105);
nor U23920 (N_23920,N_17041,N_16170);
or U23921 (N_23921,N_19000,N_15631);
nand U23922 (N_23922,N_17674,N_18114);
nor U23923 (N_23923,N_17370,N_18752);
and U23924 (N_23924,N_18258,N_19949);
and U23925 (N_23925,N_17410,N_19312);
xnor U23926 (N_23926,N_19847,N_16601);
and U23927 (N_23927,N_15221,N_15635);
xor U23928 (N_23928,N_17748,N_15106);
nor U23929 (N_23929,N_17744,N_18769);
and U23930 (N_23930,N_17126,N_17983);
or U23931 (N_23931,N_18447,N_16546);
xor U23932 (N_23932,N_17270,N_18743);
and U23933 (N_23933,N_15057,N_17102);
nor U23934 (N_23934,N_18101,N_17313);
and U23935 (N_23935,N_16853,N_15287);
nand U23936 (N_23936,N_17090,N_16562);
nand U23937 (N_23937,N_18819,N_19046);
or U23938 (N_23938,N_17483,N_19132);
and U23939 (N_23939,N_18483,N_18213);
nor U23940 (N_23940,N_19396,N_17387);
xor U23941 (N_23941,N_15926,N_18827);
xnor U23942 (N_23942,N_19289,N_19752);
xnor U23943 (N_23943,N_15973,N_16514);
nand U23944 (N_23944,N_17166,N_19966);
and U23945 (N_23945,N_17378,N_18032);
xor U23946 (N_23946,N_17841,N_18837);
or U23947 (N_23947,N_17541,N_15789);
or U23948 (N_23948,N_17293,N_19815);
nand U23949 (N_23949,N_17222,N_18126);
nor U23950 (N_23950,N_17662,N_19651);
and U23951 (N_23951,N_15193,N_17594);
and U23952 (N_23952,N_19132,N_19360);
nand U23953 (N_23953,N_18008,N_18798);
nor U23954 (N_23954,N_17891,N_18127);
xnor U23955 (N_23955,N_17465,N_19658);
nand U23956 (N_23956,N_18037,N_15867);
and U23957 (N_23957,N_16872,N_16205);
or U23958 (N_23958,N_17959,N_18188);
nand U23959 (N_23959,N_15442,N_15844);
nor U23960 (N_23960,N_18678,N_19909);
nand U23961 (N_23961,N_17482,N_16147);
and U23962 (N_23962,N_17196,N_16846);
or U23963 (N_23963,N_19706,N_15213);
xor U23964 (N_23964,N_19134,N_17770);
or U23965 (N_23965,N_18277,N_15437);
nor U23966 (N_23966,N_17767,N_19878);
and U23967 (N_23967,N_16551,N_19704);
nor U23968 (N_23968,N_19777,N_18660);
nand U23969 (N_23969,N_17215,N_15212);
xor U23970 (N_23970,N_18157,N_15068);
nand U23971 (N_23971,N_19339,N_16713);
nor U23972 (N_23972,N_15073,N_19999);
xor U23973 (N_23973,N_15578,N_18440);
xor U23974 (N_23974,N_18563,N_15222);
nand U23975 (N_23975,N_16097,N_17089);
and U23976 (N_23976,N_19526,N_16660);
xnor U23977 (N_23977,N_18020,N_17292);
xor U23978 (N_23978,N_16481,N_16284);
nor U23979 (N_23979,N_18248,N_17393);
xnor U23980 (N_23980,N_17372,N_18316);
nor U23981 (N_23981,N_16888,N_18883);
nand U23982 (N_23982,N_17732,N_18305);
xor U23983 (N_23983,N_19085,N_18651);
or U23984 (N_23984,N_17871,N_16507);
nand U23985 (N_23985,N_17670,N_17112);
and U23986 (N_23986,N_16997,N_18464);
and U23987 (N_23987,N_18153,N_15796);
or U23988 (N_23988,N_15767,N_17919);
nor U23989 (N_23989,N_16190,N_17381);
and U23990 (N_23990,N_19759,N_16903);
xnor U23991 (N_23991,N_18548,N_18287);
or U23992 (N_23992,N_18605,N_17396);
nand U23993 (N_23993,N_15330,N_17713);
nor U23994 (N_23994,N_16083,N_18400);
or U23995 (N_23995,N_17388,N_15503);
nor U23996 (N_23996,N_16103,N_17945);
nor U23997 (N_23997,N_17160,N_16432);
nor U23998 (N_23998,N_18843,N_18792);
xor U23999 (N_23999,N_18154,N_17174);
nor U24000 (N_24000,N_15891,N_15355);
xor U24001 (N_24001,N_16370,N_18526);
nand U24002 (N_24002,N_15715,N_19877);
nor U24003 (N_24003,N_16525,N_16554);
nand U24004 (N_24004,N_17837,N_17858);
nand U24005 (N_24005,N_17896,N_18699);
nand U24006 (N_24006,N_17474,N_15705);
nand U24007 (N_24007,N_19853,N_15602);
nor U24008 (N_24008,N_16678,N_16236);
nand U24009 (N_24009,N_18500,N_18008);
xor U24010 (N_24010,N_16948,N_15061);
nand U24011 (N_24011,N_18388,N_17413);
xor U24012 (N_24012,N_16264,N_16871);
and U24013 (N_24013,N_19847,N_17608);
or U24014 (N_24014,N_19070,N_18047);
xor U24015 (N_24015,N_15883,N_16028);
or U24016 (N_24016,N_17165,N_18681);
and U24017 (N_24017,N_16195,N_19339);
nor U24018 (N_24018,N_17136,N_18068);
or U24019 (N_24019,N_15115,N_17144);
nor U24020 (N_24020,N_18076,N_18270);
and U24021 (N_24021,N_17550,N_15794);
xnor U24022 (N_24022,N_17933,N_19576);
and U24023 (N_24023,N_15480,N_16780);
xnor U24024 (N_24024,N_15674,N_16027);
xnor U24025 (N_24025,N_17357,N_19671);
or U24026 (N_24026,N_19058,N_16256);
nand U24027 (N_24027,N_15876,N_18628);
nand U24028 (N_24028,N_17532,N_19599);
or U24029 (N_24029,N_19572,N_15672);
xor U24030 (N_24030,N_15927,N_19210);
xor U24031 (N_24031,N_17640,N_17749);
xor U24032 (N_24032,N_19194,N_19936);
xnor U24033 (N_24033,N_15509,N_19241);
nor U24034 (N_24034,N_17298,N_19743);
xnor U24035 (N_24035,N_15709,N_19134);
or U24036 (N_24036,N_16732,N_17210);
nand U24037 (N_24037,N_19784,N_18206);
and U24038 (N_24038,N_18353,N_19956);
nand U24039 (N_24039,N_15809,N_17406);
and U24040 (N_24040,N_19851,N_15170);
nand U24041 (N_24041,N_18066,N_16580);
nand U24042 (N_24042,N_15047,N_19514);
and U24043 (N_24043,N_16873,N_19487);
nand U24044 (N_24044,N_18937,N_18427);
nand U24045 (N_24045,N_16173,N_15032);
nand U24046 (N_24046,N_19819,N_19920);
and U24047 (N_24047,N_15393,N_16780);
and U24048 (N_24048,N_17508,N_16282);
nand U24049 (N_24049,N_17572,N_15739);
nand U24050 (N_24050,N_19497,N_16032);
xor U24051 (N_24051,N_18781,N_18873);
or U24052 (N_24052,N_16108,N_16158);
nor U24053 (N_24053,N_19490,N_19652);
or U24054 (N_24054,N_15224,N_19323);
nor U24055 (N_24055,N_16414,N_16876);
and U24056 (N_24056,N_16418,N_15099);
xor U24057 (N_24057,N_16137,N_17953);
or U24058 (N_24058,N_17151,N_18871);
xnor U24059 (N_24059,N_16372,N_15729);
or U24060 (N_24060,N_18850,N_17041);
xor U24061 (N_24061,N_19216,N_15102);
and U24062 (N_24062,N_19545,N_16004);
and U24063 (N_24063,N_15846,N_17650);
nor U24064 (N_24064,N_18127,N_18439);
and U24065 (N_24065,N_19245,N_15041);
or U24066 (N_24066,N_17386,N_15566);
xor U24067 (N_24067,N_17114,N_15956);
xnor U24068 (N_24068,N_16641,N_17738);
or U24069 (N_24069,N_18143,N_17805);
nor U24070 (N_24070,N_19835,N_15251);
nor U24071 (N_24071,N_15141,N_18484);
nand U24072 (N_24072,N_19918,N_18740);
or U24073 (N_24073,N_17374,N_15680);
or U24074 (N_24074,N_19451,N_19074);
and U24075 (N_24075,N_18027,N_15872);
nand U24076 (N_24076,N_18983,N_17775);
xor U24077 (N_24077,N_16055,N_15557);
xor U24078 (N_24078,N_17727,N_19348);
and U24079 (N_24079,N_16307,N_18042);
xor U24080 (N_24080,N_17479,N_19644);
and U24081 (N_24081,N_17863,N_19975);
nand U24082 (N_24082,N_15680,N_17066);
nor U24083 (N_24083,N_19505,N_17646);
nor U24084 (N_24084,N_19192,N_15259);
or U24085 (N_24085,N_15137,N_17539);
nor U24086 (N_24086,N_17508,N_15088);
nor U24087 (N_24087,N_18490,N_16434);
and U24088 (N_24088,N_15849,N_18914);
xor U24089 (N_24089,N_15709,N_19531);
xnor U24090 (N_24090,N_16260,N_17350);
nand U24091 (N_24091,N_15581,N_17563);
and U24092 (N_24092,N_16359,N_15648);
nor U24093 (N_24093,N_16896,N_17647);
and U24094 (N_24094,N_16306,N_16597);
and U24095 (N_24095,N_19112,N_15316);
nand U24096 (N_24096,N_18331,N_16494);
and U24097 (N_24097,N_18442,N_17711);
and U24098 (N_24098,N_16955,N_18410);
xor U24099 (N_24099,N_17851,N_15076);
or U24100 (N_24100,N_15205,N_18133);
xnor U24101 (N_24101,N_15848,N_18516);
and U24102 (N_24102,N_18733,N_18291);
and U24103 (N_24103,N_17178,N_16970);
and U24104 (N_24104,N_16767,N_18151);
xnor U24105 (N_24105,N_17004,N_17382);
nand U24106 (N_24106,N_16590,N_15194);
and U24107 (N_24107,N_17177,N_15525);
and U24108 (N_24108,N_17272,N_16258);
nor U24109 (N_24109,N_18554,N_16433);
nand U24110 (N_24110,N_17197,N_19724);
or U24111 (N_24111,N_16826,N_18362);
nor U24112 (N_24112,N_19753,N_15034);
nor U24113 (N_24113,N_17346,N_15716);
nand U24114 (N_24114,N_16853,N_15263);
xnor U24115 (N_24115,N_16737,N_16072);
or U24116 (N_24116,N_15642,N_16443);
xnor U24117 (N_24117,N_17140,N_19658);
or U24118 (N_24118,N_15425,N_17987);
xnor U24119 (N_24119,N_18257,N_17222);
or U24120 (N_24120,N_16592,N_16944);
or U24121 (N_24121,N_17440,N_17813);
nor U24122 (N_24122,N_17526,N_16025);
xnor U24123 (N_24123,N_19053,N_17979);
nor U24124 (N_24124,N_15540,N_19292);
xor U24125 (N_24125,N_17488,N_19058);
xor U24126 (N_24126,N_19272,N_16695);
nor U24127 (N_24127,N_16088,N_15283);
and U24128 (N_24128,N_17701,N_18114);
xor U24129 (N_24129,N_18646,N_15177);
nor U24130 (N_24130,N_19863,N_16427);
or U24131 (N_24131,N_15531,N_16981);
or U24132 (N_24132,N_16456,N_15160);
or U24133 (N_24133,N_19633,N_15566);
and U24134 (N_24134,N_15451,N_16520);
xor U24135 (N_24135,N_19866,N_16509);
nor U24136 (N_24136,N_16267,N_19226);
nand U24137 (N_24137,N_18998,N_19924);
and U24138 (N_24138,N_15386,N_19990);
xor U24139 (N_24139,N_16678,N_16673);
nand U24140 (N_24140,N_18911,N_15964);
nand U24141 (N_24141,N_16447,N_16860);
nor U24142 (N_24142,N_16154,N_17131);
nor U24143 (N_24143,N_18888,N_15093);
nor U24144 (N_24144,N_16170,N_19934);
and U24145 (N_24145,N_18841,N_15795);
and U24146 (N_24146,N_18939,N_16620);
nand U24147 (N_24147,N_19649,N_16910);
and U24148 (N_24148,N_16605,N_18708);
nand U24149 (N_24149,N_16305,N_17134);
or U24150 (N_24150,N_15636,N_17511);
or U24151 (N_24151,N_17430,N_16727);
nand U24152 (N_24152,N_16924,N_15891);
nand U24153 (N_24153,N_18144,N_15083);
and U24154 (N_24154,N_17392,N_18988);
or U24155 (N_24155,N_16608,N_19892);
nand U24156 (N_24156,N_17894,N_17368);
xor U24157 (N_24157,N_17111,N_15781);
xor U24158 (N_24158,N_19868,N_19823);
nor U24159 (N_24159,N_15639,N_18192);
or U24160 (N_24160,N_19580,N_15943);
xor U24161 (N_24161,N_18798,N_16020);
or U24162 (N_24162,N_18095,N_18419);
or U24163 (N_24163,N_16644,N_19975);
xnor U24164 (N_24164,N_19872,N_19765);
nand U24165 (N_24165,N_19202,N_17287);
or U24166 (N_24166,N_17882,N_15598);
or U24167 (N_24167,N_15800,N_15898);
xor U24168 (N_24168,N_18374,N_17144);
and U24169 (N_24169,N_16037,N_18917);
xor U24170 (N_24170,N_15630,N_16528);
or U24171 (N_24171,N_15987,N_16082);
or U24172 (N_24172,N_15513,N_17280);
xor U24173 (N_24173,N_16589,N_15566);
xor U24174 (N_24174,N_18749,N_15353);
nand U24175 (N_24175,N_16650,N_17164);
nand U24176 (N_24176,N_16083,N_17095);
or U24177 (N_24177,N_17773,N_19725);
or U24178 (N_24178,N_17206,N_19965);
xnor U24179 (N_24179,N_16148,N_18856);
and U24180 (N_24180,N_19398,N_17886);
and U24181 (N_24181,N_18307,N_16016);
or U24182 (N_24182,N_19462,N_16321);
nor U24183 (N_24183,N_19897,N_16486);
or U24184 (N_24184,N_18062,N_15902);
xor U24185 (N_24185,N_17580,N_17962);
or U24186 (N_24186,N_19081,N_15885);
or U24187 (N_24187,N_19510,N_19534);
nor U24188 (N_24188,N_15897,N_18710);
and U24189 (N_24189,N_15559,N_19806);
nor U24190 (N_24190,N_19807,N_15627);
xnor U24191 (N_24191,N_15060,N_16163);
and U24192 (N_24192,N_19401,N_15197);
nand U24193 (N_24193,N_16353,N_19471);
nor U24194 (N_24194,N_15180,N_17883);
xor U24195 (N_24195,N_15163,N_15496);
nand U24196 (N_24196,N_17164,N_18810);
xnor U24197 (N_24197,N_16602,N_19656);
and U24198 (N_24198,N_19124,N_15978);
or U24199 (N_24199,N_15438,N_16955);
nand U24200 (N_24200,N_15153,N_15709);
and U24201 (N_24201,N_16388,N_16453);
xnor U24202 (N_24202,N_15107,N_17631);
nor U24203 (N_24203,N_16261,N_19881);
xnor U24204 (N_24204,N_19481,N_17170);
nor U24205 (N_24205,N_19354,N_19800);
nand U24206 (N_24206,N_15629,N_16258);
or U24207 (N_24207,N_15475,N_17227);
or U24208 (N_24208,N_15601,N_17943);
xnor U24209 (N_24209,N_19138,N_15379);
xnor U24210 (N_24210,N_19192,N_18425);
or U24211 (N_24211,N_17346,N_17585);
nor U24212 (N_24212,N_17288,N_18030);
xor U24213 (N_24213,N_17622,N_16233);
nand U24214 (N_24214,N_18037,N_16619);
xor U24215 (N_24215,N_16047,N_19640);
nor U24216 (N_24216,N_16562,N_18880);
xnor U24217 (N_24217,N_16877,N_15506);
and U24218 (N_24218,N_17957,N_18926);
xnor U24219 (N_24219,N_15454,N_16642);
xnor U24220 (N_24220,N_17372,N_15350);
and U24221 (N_24221,N_18857,N_15400);
nand U24222 (N_24222,N_17719,N_19405);
and U24223 (N_24223,N_18519,N_15051);
or U24224 (N_24224,N_19046,N_19580);
nor U24225 (N_24225,N_17746,N_17523);
nor U24226 (N_24226,N_15892,N_18020);
nand U24227 (N_24227,N_19570,N_15369);
or U24228 (N_24228,N_16731,N_19058);
and U24229 (N_24229,N_18695,N_19334);
xnor U24230 (N_24230,N_15981,N_16975);
nand U24231 (N_24231,N_17494,N_16213);
and U24232 (N_24232,N_18012,N_19945);
nand U24233 (N_24233,N_19946,N_15604);
nor U24234 (N_24234,N_17479,N_17906);
nor U24235 (N_24235,N_18550,N_19427);
nand U24236 (N_24236,N_15820,N_18592);
and U24237 (N_24237,N_17025,N_19667);
xor U24238 (N_24238,N_16724,N_19098);
or U24239 (N_24239,N_15063,N_18425);
or U24240 (N_24240,N_17319,N_18527);
nor U24241 (N_24241,N_19515,N_15829);
and U24242 (N_24242,N_17655,N_19766);
nor U24243 (N_24243,N_16442,N_18948);
nor U24244 (N_24244,N_18766,N_18942);
nand U24245 (N_24245,N_15300,N_16753);
nor U24246 (N_24246,N_19619,N_18500);
nor U24247 (N_24247,N_15302,N_17788);
xnor U24248 (N_24248,N_18600,N_18718);
nor U24249 (N_24249,N_17301,N_18926);
xor U24250 (N_24250,N_16850,N_16396);
and U24251 (N_24251,N_18663,N_17633);
nor U24252 (N_24252,N_16930,N_17007);
nor U24253 (N_24253,N_19232,N_17294);
nand U24254 (N_24254,N_15289,N_16738);
and U24255 (N_24255,N_15082,N_17567);
nand U24256 (N_24256,N_18685,N_15779);
and U24257 (N_24257,N_15682,N_19255);
nor U24258 (N_24258,N_15396,N_16217);
or U24259 (N_24259,N_18754,N_16175);
nor U24260 (N_24260,N_17719,N_19278);
nand U24261 (N_24261,N_18755,N_17638);
nand U24262 (N_24262,N_17798,N_15985);
nand U24263 (N_24263,N_15537,N_18485);
or U24264 (N_24264,N_17011,N_16076);
or U24265 (N_24265,N_17457,N_19490);
xnor U24266 (N_24266,N_19785,N_16020);
xor U24267 (N_24267,N_15286,N_15663);
and U24268 (N_24268,N_16317,N_19118);
xnor U24269 (N_24269,N_17233,N_17431);
nor U24270 (N_24270,N_17380,N_17556);
and U24271 (N_24271,N_16633,N_17554);
xnor U24272 (N_24272,N_18596,N_19949);
nand U24273 (N_24273,N_18737,N_19022);
nand U24274 (N_24274,N_19321,N_15753);
xor U24275 (N_24275,N_18885,N_18583);
or U24276 (N_24276,N_18808,N_17980);
nand U24277 (N_24277,N_16096,N_17040);
or U24278 (N_24278,N_17751,N_15335);
and U24279 (N_24279,N_17774,N_17295);
nor U24280 (N_24280,N_17876,N_19390);
and U24281 (N_24281,N_19422,N_17273);
and U24282 (N_24282,N_18273,N_15608);
xor U24283 (N_24283,N_15354,N_17546);
xnor U24284 (N_24284,N_17067,N_17441);
nand U24285 (N_24285,N_19239,N_19092);
nor U24286 (N_24286,N_19898,N_17442);
or U24287 (N_24287,N_17380,N_19686);
and U24288 (N_24288,N_16578,N_18740);
nand U24289 (N_24289,N_18541,N_18376);
nor U24290 (N_24290,N_15517,N_16065);
xnor U24291 (N_24291,N_16557,N_15325);
or U24292 (N_24292,N_17306,N_16676);
and U24293 (N_24293,N_17831,N_15300);
and U24294 (N_24294,N_17801,N_19867);
nand U24295 (N_24295,N_15338,N_17173);
and U24296 (N_24296,N_19515,N_18709);
nand U24297 (N_24297,N_17347,N_18661);
and U24298 (N_24298,N_19706,N_17433);
nor U24299 (N_24299,N_16301,N_19237);
or U24300 (N_24300,N_19766,N_15008);
nand U24301 (N_24301,N_15163,N_19421);
xnor U24302 (N_24302,N_19791,N_16953);
nand U24303 (N_24303,N_15100,N_16681);
xor U24304 (N_24304,N_18673,N_19346);
nand U24305 (N_24305,N_17203,N_16003);
or U24306 (N_24306,N_18556,N_15475);
nor U24307 (N_24307,N_18317,N_15001);
xor U24308 (N_24308,N_17048,N_16057);
or U24309 (N_24309,N_17226,N_17907);
or U24310 (N_24310,N_19838,N_18476);
nand U24311 (N_24311,N_17684,N_19098);
nor U24312 (N_24312,N_15311,N_17807);
or U24313 (N_24313,N_19510,N_18708);
xnor U24314 (N_24314,N_16073,N_15213);
and U24315 (N_24315,N_19167,N_15261);
xor U24316 (N_24316,N_19892,N_19096);
nand U24317 (N_24317,N_19984,N_15389);
and U24318 (N_24318,N_18435,N_17456);
xor U24319 (N_24319,N_19257,N_17485);
nor U24320 (N_24320,N_15863,N_18171);
nor U24321 (N_24321,N_17515,N_17269);
nand U24322 (N_24322,N_16975,N_15788);
and U24323 (N_24323,N_18068,N_17352);
xnor U24324 (N_24324,N_15579,N_18278);
and U24325 (N_24325,N_16616,N_17744);
xor U24326 (N_24326,N_18473,N_16152);
xor U24327 (N_24327,N_15012,N_19443);
nand U24328 (N_24328,N_17471,N_19218);
xor U24329 (N_24329,N_19096,N_19809);
nor U24330 (N_24330,N_17537,N_18933);
nor U24331 (N_24331,N_18553,N_18997);
xor U24332 (N_24332,N_16798,N_19783);
nand U24333 (N_24333,N_19616,N_17657);
or U24334 (N_24334,N_19409,N_17659);
xor U24335 (N_24335,N_19605,N_15714);
nand U24336 (N_24336,N_15143,N_16596);
nor U24337 (N_24337,N_15134,N_15503);
nand U24338 (N_24338,N_17666,N_17569);
xor U24339 (N_24339,N_19543,N_15657);
nand U24340 (N_24340,N_17047,N_16105);
nand U24341 (N_24341,N_17327,N_19296);
nor U24342 (N_24342,N_15271,N_19783);
or U24343 (N_24343,N_15672,N_19113);
and U24344 (N_24344,N_18657,N_18758);
and U24345 (N_24345,N_15954,N_18792);
nand U24346 (N_24346,N_19265,N_19214);
nor U24347 (N_24347,N_18545,N_15884);
xor U24348 (N_24348,N_17619,N_19097);
and U24349 (N_24349,N_15153,N_15323);
xnor U24350 (N_24350,N_15424,N_16740);
xnor U24351 (N_24351,N_15946,N_16578);
xor U24352 (N_24352,N_18094,N_18254);
xnor U24353 (N_24353,N_18335,N_18587);
nand U24354 (N_24354,N_16527,N_18704);
and U24355 (N_24355,N_15116,N_15951);
nor U24356 (N_24356,N_18110,N_18596);
xnor U24357 (N_24357,N_17686,N_15339);
nand U24358 (N_24358,N_18328,N_18466);
nand U24359 (N_24359,N_15918,N_17650);
nand U24360 (N_24360,N_18980,N_18778);
nor U24361 (N_24361,N_15027,N_19304);
nand U24362 (N_24362,N_16827,N_15155);
or U24363 (N_24363,N_17206,N_18981);
nor U24364 (N_24364,N_19072,N_15305);
and U24365 (N_24365,N_19162,N_19093);
nor U24366 (N_24366,N_16127,N_15265);
xnor U24367 (N_24367,N_16889,N_19429);
or U24368 (N_24368,N_17693,N_16301);
and U24369 (N_24369,N_15133,N_16344);
or U24370 (N_24370,N_17675,N_15767);
xnor U24371 (N_24371,N_15735,N_19828);
xor U24372 (N_24372,N_19128,N_15164);
nor U24373 (N_24373,N_16643,N_18398);
xnor U24374 (N_24374,N_16796,N_16261);
and U24375 (N_24375,N_19157,N_16725);
xnor U24376 (N_24376,N_17923,N_16633);
and U24377 (N_24377,N_17291,N_18724);
or U24378 (N_24378,N_16889,N_18863);
nand U24379 (N_24379,N_16215,N_17242);
nor U24380 (N_24380,N_17879,N_15400);
or U24381 (N_24381,N_15891,N_17546);
and U24382 (N_24382,N_19530,N_15758);
or U24383 (N_24383,N_15533,N_19863);
nand U24384 (N_24384,N_17788,N_18131);
nand U24385 (N_24385,N_18233,N_18389);
and U24386 (N_24386,N_16641,N_17482);
nor U24387 (N_24387,N_17005,N_15073);
and U24388 (N_24388,N_15139,N_17597);
nand U24389 (N_24389,N_15854,N_17833);
nand U24390 (N_24390,N_17266,N_18849);
xor U24391 (N_24391,N_16856,N_15955);
nand U24392 (N_24392,N_15520,N_17074);
and U24393 (N_24393,N_18673,N_15823);
and U24394 (N_24394,N_15655,N_18959);
or U24395 (N_24395,N_16687,N_18992);
nor U24396 (N_24396,N_18035,N_15652);
or U24397 (N_24397,N_16922,N_17455);
nand U24398 (N_24398,N_15779,N_16010);
nor U24399 (N_24399,N_19228,N_18935);
nor U24400 (N_24400,N_17855,N_18318);
and U24401 (N_24401,N_19390,N_16320);
or U24402 (N_24402,N_15737,N_15832);
nand U24403 (N_24403,N_18970,N_16053);
xnor U24404 (N_24404,N_16384,N_17395);
xnor U24405 (N_24405,N_17822,N_18691);
xnor U24406 (N_24406,N_15673,N_15788);
nand U24407 (N_24407,N_18242,N_16587);
nand U24408 (N_24408,N_19565,N_16299);
or U24409 (N_24409,N_17374,N_16718);
xor U24410 (N_24410,N_19959,N_16207);
xnor U24411 (N_24411,N_16582,N_16450);
and U24412 (N_24412,N_17013,N_15729);
nand U24413 (N_24413,N_16099,N_18618);
or U24414 (N_24414,N_18580,N_19455);
nor U24415 (N_24415,N_15229,N_16475);
and U24416 (N_24416,N_16383,N_18925);
and U24417 (N_24417,N_17266,N_18227);
nand U24418 (N_24418,N_19079,N_17218);
nand U24419 (N_24419,N_18975,N_17576);
xor U24420 (N_24420,N_18361,N_16676);
nand U24421 (N_24421,N_16031,N_17242);
nand U24422 (N_24422,N_15102,N_19723);
nor U24423 (N_24423,N_18366,N_16418);
xor U24424 (N_24424,N_16019,N_19103);
or U24425 (N_24425,N_19569,N_18234);
nor U24426 (N_24426,N_19381,N_15856);
and U24427 (N_24427,N_18624,N_16139);
nand U24428 (N_24428,N_18101,N_17365);
nor U24429 (N_24429,N_16498,N_18427);
or U24430 (N_24430,N_16762,N_17597);
nor U24431 (N_24431,N_19286,N_17289);
xnor U24432 (N_24432,N_16655,N_17668);
nand U24433 (N_24433,N_18574,N_15112);
nor U24434 (N_24434,N_18429,N_19655);
or U24435 (N_24435,N_18264,N_18256);
or U24436 (N_24436,N_16642,N_17662);
nor U24437 (N_24437,N_19298,N_19663);
nand U24438 (N_24438,N_16192,N_15756);
nand U24439 (N_24439,N_17810,N_15682);
xor U24440 (N_24440,N_19210,N_17503);
and U24441 (N_24441,N_18230,N_18880);
nand U24442 (N_24442,N_16581,N_19671);
or U24443 (N_24443,N_17110,N_17921);
and U24444 (N_24444,N_18032,N_15781);
or U24445 (N_24445,N_19902,N_16380);
nand U24446 (N_24446,N_19301,N_16473);
nand U24447 (N_24447,N_15012,N_15575);
or U24448 (N_24448,N_15926,N_17074);
xnor U24449 (N_24449,N_16089,N_19794);
or U24450 (N_24450,N_17787,N_16702);
nor U24451 (N_24451,N_19127,N_17904);
or U24452 (N_24452,N_16674,N_18164);
or U24453 (N_24453,N_18831,N_15468);
nor U24454 (N_24454,N_16005,N_17509);
nor U24455 (N_24455,N_19412,N_18097);
nor U24456 (N_24456,N_19510,N_19209);
and U24457 (N_24457,N_18898,N_18977);
xnor U24458 (N_24458,N_19084,N_15984);
and U24459 (N_24459,N_18313,N_19538);
and U24460 (N_24460,N_17176,N_15859);
nor U24461 (N_24461,N_18868,N_16113);
nor U24462 (N_24462,N_18901,N_17573);
nor U24463 (N_24463,N_17433,N_18846);
xnor U24464 (N_24464,N_15540,N_17884);
and U24465 (N_24465,N_18041,N_18774);
or U24466 (N_24466,N_19507,N_15276);
or U24467 (N_24467,N_16323,N_19839);
nand U24468 (N_24468,N_15782,N_15975);
or U24469 (N_24469,N_18835,N_16134);
or U24470 (N_24470,N_16680,N_16616);
or U24471 (N_24471,N_16086,N_18178);
and U24472 (N_24472,N_18555,N_15414);
or U24473 (N_24473,N_15464,N_16750);
or U24474 (N_24474,N_19274,N_18712);
xnor U24475 (N_24475,N_19594,N_17906);
xor U24476 (N_24476,N_16771,N_16595);
or U24477 (N_24477,N_16290,N_17508);
nand U24478 (N_24478,N_18827,N_17933);
nor U24479 (N_24479,N_19492,N_17204);
and U24480 (N_24480,N_16610,N_16571);
nand U24481 (N_24481,N_17944,N_15282);
xor U24482 (N_24482,N_16500,N_18884);
xor U24483 (N_24483,N_16549,N_18260);
and U24484 (N_24484,N_19566,N_17667);
or U24485 (N_24485,N_18261,N_16229);
or U24486 (N_24486,N_18549,N_18957);
and U24487 (N_24487,N_18698,N_15303);
xor U24488 (N_24488,N_18990,N_16417);
xnor U24489 (N_24489,N_18421,N_17000);
or U24490 (N_24490,N_16077,N_18759);
xnor U24491 (N_24491,N_15255,N_19914);
xor U24492 (N_24492,N_19580,N_16626);
xnor U24493 (N_24493,N_17513,N_16949);
and U24494 (N_24494,N_16367,N_16673);
and U24495 (N_24495,N_18993,N_18570);
and U24496 (N_24496,N_15134,N_15720);
and U24497 (N_24497,N_15992,N_19338);
and U24498 (N_24498,N_19200,N_16814);
and U24499 (N_24499,N_17148,N_15422);
nand U24500 (N_24500,N_15891,N_16655);
and U24501 (N_24501,N_15473,N_16236);
nand U24502 (N_24502,N_19204,N_19098);
and U24503 (N_24503,N_18042,N_16702);
nand U24504 (N_24504,N_15417,N_15914);
nand U24505 (N_24505,N_19816,N_19622);
nand U24506 (N_24506,N_18358,N_19360);
or U24507 (N_24507,N_18325,N_15944);
or U24508 (N_24508,N_18114,N_17126);
and U24509 (N_24509,N_16861,N_18985);
xnor U24510 (N_24510,N_19622,N_19032);
or U24511 (N_24511,N_19088,N_19676);
xnor U24512 (N_24512,N_16558,N_18806);
xor U24513 (N_24513,N_16199,N_16258);
xor U24514 (N_24514,N_15089,N_16520);
nand U24515 (N_24515,N_19323,N_19741);
or U24516 (N_24516,N_16536,N_17006);
nand U24517 (N_24517,N_19987,N_16825);
or U24518 (N_24518,N_16499,N_15757);
xor U24519 (N_24519,N_18412,N_17616);
xnor U24520 (N_24520,N_18628,N_15377);
nand U24521 (N_24521,N_19967,N_18264);
xor U24522 (N_24522,N_16500,N_17024);
xnor U24523 (N_24523,N_16172,N_16627);
xnor U24524 (N_24524,N_19896,N_15710);
or U24525 (N_24525,N_19475,N_19326);
or U24526 (N_24526,N_15823,N_16767);
and U24527 (N_24527,N_18835,N_16886);
or U24528 (N_24528,N_19088,N_19121);
and U24529 (N_24529,N_18127,N_19696);
xor U24530 (N_24530,N_19137,N_17820);
nand U24531 (N_24531,N_17194,N_16652);
and U24532 (N_24532,N_18454,N_18353);
and U24533 (N_24533,N_16852,N_19636);
nor U24534 (N_24534,N_19847,N_17503);
or U24535 (N_24535,N_16580,N_18510);
or U24536 (N_24536,N_19089,N_17787);
xor U24537 (N_24537,N_18452,N_17012);
and U24538 (N_24538,N_15595,N_17488);
or U24539 (N_24539,N_16868,N_18502);
or U24540 (N_24540,N_16038,N_18244);
xnor U24541 (N_24541,N_19594,N_15579);
xnor U24542 (N_24542,N_19430,N_19144);
xor U24543 (N_24543,N_16336,N_17718);
nor U24544 (N_24544,N_15563,N_16208);
nor U24545 (N_24545,N_18691,N_19233);
and U24546 (N_24546,N_15882,N_19832);
nor U24547 (N_24547,N_17028,N_15432);
nand U24548 (N_24548,N_16228,N_19196);
xor U24549 (N_24549,N_18862,N_18893);
or U24550 (N_24550,N_18069,N_17884);
and U24551 (N_24551,N_17738,N_17172);
or U24552 (N_24552,N_16946,N_18121);
nand U24553 (N_24553,N_18299,N_17004);
nand U24554 (N_24554,N_16242,N_15279);
or U24555 (N_24555,N_17520,N_16854);
and U24556 (N_24556,N_17547,N_18577);
nor U24557 (N_24557,N_16235,N_15567);
and U24558 (N_24558,N_15630,N_19193);
and U24559 (N_24559,N_16917,N_15402);
nand U24560 (N_24560,N_15305,N_16172);
or U24561 (N_24561,N_15480,N_19711);
nand U24562 (N_24562,N_17873,N_19263);
xnor U24563 (N_24563,N_19176,N_15621);
or U24564 (N_24564,N_17333,N_16346);
xor U24565 (N_24565,N_19512,N_16858);
nor U24566 (N_24566,N_16079,N_15989);
nor U24567 (N_24567,N_18396,N_17719);
xnor U24568 (N_24568,N_17773,N_19306);
nor U24569 (N_24569,N_16885,N_17098);
or U24570 (N_24570,N_18028,N_18564);
and U24571 (N_24571,N_15936,N_19758);
and U24572 (N_24572,N_17573,N_18258);
xor U24573 (N_24573,N_17829,N_17183);
and U24574 (N_24574,N_19680,N_18334);
nor U24575 (N_24575,N_17254,N_19310);
or U24576 (N_24576,N_16236,N_17698);
xor U24577 (N_24577,N_16494,N_19672);
and U24578 (N_24578,N_18951,N_19611);
nand U24579 (N_24579,N_15121,N_17096);
or U24580 (N_24580,N_19154,N_18215);
or U24581 (N_24581,N_16497,N_15523);
and U24582 (N_24582,N_17987,N_17603);
and U24583 (N_24583,N_16109,N_16453);
xor U24584 (N_24584,N_16994,N_15485);
nor U24585 (N_24585,N_18533,N_15880);
or U24586 (N_24586,N_18605,N_17087);
or U24587 (N_24587,N_19640,N_19143);
nor U24588 (N_24588,N_19542,N_18873);
nand U24589 (N_24589,N_18491,N_19930);
or U24590 (N_24590,N_15353,N_15922);
and U24591 (N_24591,N_19186,N_17897);
nor U24592 (N_24592,N_18060,N_16903);
nand U24593 (N_24593,N_16951,N_16232);
xor U24594 (N_24594,N_15426,N_16001);
or U24595 (N_24595,N_18475,N_19692);
nand U24596 (N_24596,N_17763,N_16208);
or U24597 (N_24597,N_18380,N_16867);
xor U24598 (N_24598,N_19188,N_15347);
or U24599 (N_24599,N_19360,N_19939);
nand U24600 (N_24600,N_17995,N_16509);
nor U24601 (N_24601,N_17418,N_18656);
nor U24602 (N_24602,N_16091,N_19406);
nor U24603 (N_24603,N_15274,N_15985);
or U24604 (N_24604,N_16112,N_16308);
nor U24605 (N_24605,N_17077,N_19389);
or U24606 (N_24606,N_16256,N_19878);
and U24607 (N_24607,N_16356,N_18783);
nand U24608 (N_24608,N_17083,N_15781);
nor U24609 (N_24609,N_18595,N_18758);
xnor U24610 (N_24610,N_19205,N_17791);
and U24611 (N_24611,N_15848,N_16780);
and U24612 (N_24612,N_15234,N_15839);
xnor U24613 (N_24613,N_17819,N_15461);
nand U24614 (N_24614,N_16859,N_19790);
nor U24615 (N_24615,N_15298,N_18304);
and U24616 (N_24616,N_18564,N_16636);
nor U24617 (N_24617,N_17605,N_17312);
nor U24618 (N_24618,N_19422,N_17096);
or U24619 (N_24619,N_16630,N_16381);
nor U24620 (N_24620,N_18067,N_18385);
or U24621 (N_24621,N_16987,N_17643);
xor U24622 (N_24622,N_19386,N_15907);
nand U24623 (N_24623,N_18532,N_19525);
nor U24624 (N_24624,N_16351,N_17494);
and U24625 (N_24625,N_17543,N_16788);
or U24626 (N_24626,N_17780,N_16489);
nand U24627 (N_24627,N_16727,N_19025);
nor U24628 (N_24628,N_16953,N_17890);
and U24629 (N_24629,N_18792,N_18816);
and U24630 (N_24630,N_16622,N_15214);
xor U24631 (N_24631,N_18451,N_18710);
nand U24632 (N_24632,N_15488,N_17290);
xnor U24633 (N_24633,N_19596,N_15574);
or U24634 (N_24634,N_18272,N_15854);
and U24635 (N_24635,N_17395,N_15013);
nor U24636 (N_24636,N_15688,N_16218);
or U24637 (N_24637,N_15958,N_18914);
nand U24638 (N_24638,N_15143,N_15873);
nor U24639 (N_24639,N_16744,N_15900);
xor U24640 (N_24640,N_16134,N_15127);
nor U24641 (N_24641,N_15396,N_18348);
nand U24642 (N_24642,N_17014,N_19662);
xnor U24643 (N_24643,N_19018,N_18515);
xor U24644 (N_24644,N_16686,N_19539);
and U24645 (N_24645,N_19751,N_17086);
xnor U24646 (N_24646,N_18888,N_17341);
nor U24647 (N_24647,N_19208,N_18850);
nor U24648 (N_24648,N_15526,N_19252);
nand U24649 (N_24649,N_16080,N_19190);
xnor U24650 (N_24650,N_18297,N_19909);
nand U24651 (N_24651,N_15849,N_19596);
and U24652 (N_24652,N_19994,N_17551);
xor U24653 (N_24653,N_18687,N_18870);
xor U24654 (N_24654,N_18983,N_15016);
nor U24655 (N_24655,N_17040,N_18942);
xor U24656 (N_24656,N_17958,N_17006);
or U24657 (N_24657,N_19549,N_15464);
nor U24658 (N_24658,N_17756,N_19320);
and U24659 (N_24659,N_16757,N_16753);
and U24660 (N_24660,N_16752,N_15646);
nor U24661 (N_24661,N_15293,N_19523);
nand U24662 (N_24662,N_19631,N_17845);
nor U24663 (N_24663,N_19689,N_15333);
nand U24664 (N_24664,N_16361,N_17303);
nand U24665 (N_24665,N_16364,N_15251);
xnor U24666 (N_24666,N_19556,N_15472);
xnor U24667 (N_24667,N_16125,N_16671);
and U24668 (N_24668,N_15030,N_15304);
xor U24669 (N_24669,N_17483,N_18687);
or U24670 (N_24670,N_18858,N_18310);
nor U24671 (N_24671,N_17401,N_19705);
or U24672 (N_24672,N_15756,N_15866);
nor U24673 (N_24673,N_18337,N_18489);
nand U24674 (N_24674,N_16256,N_19069);
nand U24675 (N_24675,N_17884,N_17547);
and U24676 (N_24676,N_18451,N_15405);
and U24677 (N_24677,N_17584,N_17138);
xor U24678 (N_24678,N_17163,N_17434);
or U24679 (N_24679,N_17782,N_16057);
xnor U24680 (N_24680,N_16510,N_15256);
or U24681 (N_24681,N_18932,N_15819);
nor U24682 (N_24682,N_19802,N_17932);
nand U24683 (N_24683,N_17426,N_19399);
nor U24684 (N_24684,N_19154,N_19839);
nand U24685 (N_24685,N_16088,N_16420);
or U24686 (N_24686,N_16590,N_18139);
or U24687 (N_24687,N_18866,N_19113);
and U24688 (N_24688,N_16476,N_17022);
and U24689 (N_24689,N_17996,N_17871);
nor U24690 (N_24690,N_15360,N_18336);
or U24691 (N_24691,N_16231,N_19813);
or U24692 (N_24692,N_19415,N_17055);
nor U24693 (N_24693,N_19613,N_16222);
and U24694 (N_24694,N_17878,N_16526);
nor U24695 (N_24695,N_19982,N_18119);
xor U24696 (N_24696,N_17757,N_15859);
xnor U24697 (N_24697,N_15686,N_16886);
xor U24698 (N_24698,N_16529,N_18283);
and U24699 (N_24699,N_17050,N_18843);
or U24700 (N_24700,N_18019,N_16947);
nand U24701 (N_24701,N_15979,N_16317);
nor U24702 (N_24702,N_19117,N_15902);
nor U24703 (N_24703,N_15660,N_17616);
or U24704 (N_24704,N_16529,N_15422);
or U24705 (N_24705,N_16897,N_15271);
or U24706 (N_24706,N_17053,N_18162);
xor U24707 (N_24707,N_17913,N_19450);
nand U24708 (N_24708,N_15084,N_19378);
nor U24709 (N_24709,N_16714,N_18201);
or U24710 (N_24710,N_17998,N_16156);
nor U24711 (N_24711,N_15924,N_15067);
nand U24712 (N_24712,N_17381,N_18000);
nand U24713 (N_24713,N_16792,N_16805);
and U24714 (N_24714,N_16387,N_15184);
xor U24715 (N_24715,N_18138,N_19887);
or U24716 (N_24716,N_17327,N_19229);
nor U24717 (N_24717,N_17341,N_16223);
nor U24718 (N_24718,N_17032,N_16238);
and U24719 (N_24719,N_18332,N_16473);
or U24720 (N_24720,N_19515,N_17083);
nor U24721 (N_24721,N_16317,N_15748);
nand U24722 (N_24722,N_19477,N_19885);
or U24723 (N_24723,N_17725,N_19715);
or U24724 (N_24724,N_15204,N_16190);
nor U24725 (N_24725,N_19383,N_19997);
or U24726 (N_24726,N_15562,N_15539);
nand U24727 (N_24727,N_17731,N_15710);
nand U24728 (N_24728,N_16622,N_18133);
and U24729 (N_24729,N_15248,N_15200);
and U24730 (N_24730,N_17774,N_17928);
or U24731 (N_24731,N_18910,N_15783);
nand U24732 (N_24732,N_17962,N_15212);
and U24733 (N_24733,N_15352,N_16987);
nand U24734 (N_24734,N_15072,N_17547);
xor U24735 (N_24735,N_17466,N_18142);
nor U24736 (N_24736,N_15737,N_19364);
nor U24737 (N_24737,N_16873,N_17525);
xor U24738 (N_24738,N_16431,N_19005);
nor U24739 (N_24739,N_18161,N_18275);
or U24740 (N_24740,N_16024,N_17712);
and U24741 (N_24741,N_17070,N_19537);
xnor U24742 (N_24742,N_18805,N_19927);
and U24743 (N_24743,N_18452,N_19797);
nand U24744 (N_24744,N_15502,N_15926);
nor U24745 (N_24745,N_16549,N_18400);
nand U24746 (N_24746,N_17509,N_16792);
or U24747 (N_24747,N_19226,N_16919);
nand U24748 (N_24748,N_17207,N_17776);
nand U24749 (N_24749,N_18405,N_18203);
nor U24750 (N_24750,N_19564,N_16799);
and U24751 (N_24751,N_15625,N_19372);
or U24752 (N_24752,N_17982,N_18748);
nor U24753 (N_24753,N_15076,N_18557);
nand U24754 (N_24754,N_15388,N_16799);
and U24755 (N_24755,N_16762,N_15993);
nor U24756 (N_24756,N_19568,N_16069);
nand U24757 (N_24757,N_18606,N_16198);
xnor U24758 (N_24758,N_15205,N_18872);
or U24759 (N_24759,N_15912,N_15492);
nor U24760 (N_24760,N_19793,N_19461);
nand U24761 (N_24761,N_17119,N_19550);
nand U24762 (N_24762,N_19037,N_16783);
nand U24763 (N_24763,N_17441,N_15054);
or U24764 (N_24764,N_19712,N_19321);
or U24765 (N_24765,N_17365,N_15276);
xnor U24766 (N_24766,N_19281,N_17477);
or U24767 (N_24767,N_17096,N_19653);
nor U24768 (N_24768,N_19217,N_18625);
and U24769 (N_24769,N_17708,N_15734);
nand U24770 (N_24770,N_19371,N_16880);
and U24771 (N_24771,N_15968,N_19638);
xor U24772 (N_24772,N_19246,N_16236);
nand U24773 (N_24773,N_15005,N_19925);
xor U24774 (N_24774,N_19089,N_15872);
and U24775 (N_24775,N_18623,N_16007);
and U24776 (N_24776,N_15264,N_16615);
xor U24777 (N_24777,N_16860,N_15320);
and U24778 (N_24778,N_15724,N_18444);
xor U24779 (N_24779,N_17441,N_16880);
xnor U24780 (N_24780,N_15007,N_15967);
nand U24781 (N_24781,N_15486,N_19433);
xnor U24782 (N_24782,N_18732,N_17091);
nand U24783 (N_24783,N_18899,N_17622);
xor U24784 (N_24784,N_16742,N_18111);
nand U24785 (N_24785,N_15541,N_17663);
nand U24786 (N_24786,N_18844,N_17011);
and U24787 (N_24787,N_16358,N_19678);
or U24788 (N_24788,N_16726,N_16827);
and U24789 (N_24789,N_15858,N_15035);
xor U24790 (N_24790,N_17313,N_15974);
and U24791 (N_24791,N_19481,N_19604);
and U24792 (N_24792,N_19403,N_17286);
nor U24793 (N_24793,N_16670,N_17500);
nor U24794 (N_24794,N_18992,N_17832);
nand U24795 (N_24795,N_18021,N_18090);
or U24796 (N_24796,N_18037,N_15697);
or U24797 (N_24797,N_17530,N_15631);
nand U24798 (N_24798,N_15655,N_19550);
and U24799 (N_24799,N_17898,N_17344);
or U24800 (N_24800,N_19740,N_15853);
xor U24801 (N_24801,N_17498,N_17850);
or U24802 (N_24802,N_16240,N_15751);
nor U24803 (N_24803,N_18689,N_16621);
nand U24804 (N_24804,N_15246,N_18148);
xnor U24805 (N_24805,N_15245,N_16232);
or U24806 (N_24806,N_17118,N_15994);
nor U24807 (N_24807,N_16576,N_15687);
xor U24808 (N_24808,N_15861,N_19925);
or U24809 (N_24809,N_18332,N_16713);
nand U24810 (N_24810,N_17289,N_18741);
xor U24811 (N_24811,N_15700,N_17716);
xnor U24812 (N_24812,N_17277,N_15594);
and U24813 (N_24813,N_15103,N_15931);
xor U24814 (N_24814,N_17429,N_17251);
and U24815 (N_24815,N_15184,N_18883);
nor U24816 (N_24816,N_15230,N_16727);
or U24817 (N_24817,N_15015,N_16632);
xnor U24818 (N_24818,N_15132,N_15751);
xnor U24819 (N_24819,N_15029,N_19853);
nor U24820 (N_24820,N_19040,N_18537);
nand U24821 (N_24821,N_18943,N_15007);
or U24822 (N_24822,N_18606,N_15311);
and U24823 (N_24823,N_16160,N_16116);
xor U24824 (N_24824,N_18184,N_18062);
nor U24825 (N_24825,N_17030,N_16927);
xnor U24826 (N_24826,N_19281,N_18261);
nand U24827 (N_24827,N_16143,N_16337);
nor U24828 (N_24828,N_19353,N_19111);
nor U24829 (N_24829,N_16173,N_19951);
or U24830 (N_24830,N_16301,N_15587);
or U24831 (N_24831,N_16654,N_15880);
nor U24832 (N_24832,N_15387,N_19850);
nor U24833 (N_24833,N_16886,N_17323);
nor U24834 (N_24834,N_17867,N_17360);
or U24835 (N_24835,N_19249,N_15462);
or U24836 (N_24836,N_19745,N_18949);
and U24837 (N_24837,N_19664,N_15087);
nand U24838 (N_24838,N_18161,N_17470);
or U24839 (N_24839,N_19587,N_18725);
nor U24840 (N_24840,N_19021,N_18667);
or U24841 (N_24841,N_15667,N_18109);
or U24842 (N_24842,N_15974,N_17589);
or U24843 (N_24843,N_18212,N_17205);
or U24844 (N_24844,N_15778,N_17285);
xnor U24845 (N_24845,N_19330,N_16595);
xor U24846 (N_24846,N_15117,N_17625);
xnor U24847 (N_24847,N_19300,N_19648);
nor U24848 (N_24848,N_17872,N_19410);
nor U24849 (N_24849,N_16043,N_15890);
or U24850 (N_24850,N_15004,N_17109);
xnor U24851 (N_24851,N_18004,N_16151);
xor U24852 (N_24852,N_15699,N_19407);
nand U24853 (N_24853,N_15621,N_17495);
or U24854 (N_24854,N_17321,N_18871);
nor U24855 (N_24855,N_17239,N_17958);
and U24856 (N_24856,N_19458,N_19020);
nand U24857 (N_24857,N_19587,N_15075);
or U24858 (N_24858,N_19917,N_19944);
nand U24859 (N_24859,N_17837,N_15607);
and U24860 (N_24860,N_19255,N_18146);
nand U24861 (N_24861,N_19611,N_17697);
or U24862 (N_24862,N_19035,N_18152);
nor U24863 (N_24863,N_17601,N_19358);
nor U24864 (N_24864,N_19169,N_16101);
and U24865 (N_24865,N_19308,N_18197);
nor U24866 (N_24866,N_16265,N_17583);
nand U24867 (N_24867,N_16559,N_17054);
nor U24868 (N_24868,N_18373,N_17217);
and U24869 (N_24869,N_15466,N_17912);
xor U24870 (N_24870,N_19655,N_19783);
nor U24871 (N_24871,N_19135,N_18093);
and U24872 (N_24872,N_15916,N_19404);
nor U24873 (N_24873,N_19304,N_17219);
and U24874 (N_24874,N_17828,N_16268);
xnor U24875 (N_24875,N_15788,N_19171);
nand U24876 (N_24876,N_16620,N_16495);
xor U24877 (N_24877,N_16449,N_17790);
nor U24878 (N_24878,N_18567,N_17346);
or U24879 (N_24879,N_18049,N_17404);
nor U24880 (N_24880,N_16795,N_16566);
nand U24881 (N_24881,N_18276,N_16093);
or U24882 (N_24882,N_17897,N_18745);
and U24883 (N_24883,N_19438,N_19233);
nor U24884 (N_24884,N_18906,N_19984);
or U24885 (N_24885,N_15845,N_19422);
or U24886 (N_24886,N_16772,N_17088);
and U24887 (N_24887,N_18215,N_15432);
nand U24888 (N_24888,N_17795,N_16391);
and U24889 (N_24889,N_18808,N_16345);
nor U24890 (N_24890,N_17150,N_16661);
nor U24891 (N_24891,N_19389,N_17383);
and U24892 (N_24892,N_15606,N_18406);
or U24893 (N_24893,N_16151,N_16286);
and U24894 (N_24894,N_19515,N_16103);
or U24895 (N_24895,N_18563,N_19297);
and U24896 (N_24896,N_16069,N_15956);
nand U24897 (N_24897,N_16336,N_18943);
xor U24898 (N_24898,N_17427,N_18873);
nor U24899 (N_24899,N_16861,N_19872);
xnor U24900 (N_24900,N_19666,N_19818);
and U24901 (N_24901,N_19825,N_18881);
or U24902 (N_24902,N_18501,N_16136);
xor U24903 (N_24903,N_19660,N_19090);
xnor U24904 (N_24904,N_15960,N_16320);
nand U24905 (N_24905,N_16711,N_19903);
nor U24906 (N_24906,N_19809,N_19861);
nor U24907 (N_24907,N_17502,N_16710);
and U24908 (N_24908,N_16126,N_17092);
and U24909 (N_24909,N_19343,N_18839);
nand U24910 (N_24910,N_16511,N_15996);
and U24911 (N_24911,N_19948,N_16158);
nand U24912 (N_24912,N_18981,N_15573);
and U24913 (N_24913,N_17100,N_17121);
nand U24914 (N_24914,N_19625,N_18424);
nor U24915 (N_24915,N_18170,N_18028);
or U24916 (N_24916,N_18406,N_18540);
and U24917 (N_24917,N_19753,N_16636);
nand U24918 (N_24918,N_16456,N_17903);
and U24919 (N_24919,N_17435,N_15799);
nor U24920 (N_24920,N_15933,N_15187);
xor U24921 (N_24921,N_16797,N_18162);
and U24922 (N_24922,N_19391,N_18320);
or U24923 (N_24923,N_15508,N_19181);
xnor U24924 (N_24924,N_15682,N_17089);
or U24925 (N_24925,N_15093,N_15596);
or U24926 (N_24926,N_18654,N_19343);
nor U24927 (N_24927,N_19457,N_18562);
and U24928 (N_24928,N_15163,N_18003);
or U24929 (N_24929,N_18879,N_15766);
xor U24930 (N_24930,N_18839,N_17314);
xnor U24931 (N_24931,N_16189,N_16407);
and U24932 (N_24932,N_18300,N_17196);
xnor U24933 (N_24933,N_19750,N_15499);
or U24934 (N_24934,N_19685,N_15650);
nand U24935 (N_24935,N_18684,N_19553);
nor U24936 (N_24936,N_15252,N_19253);
and U24937 (N_24937,N_16900,N_16402);
and U24938 (N_24938,N_19438,N_16543);
nand U24939 (N_24939,N_19588,N_18504);
nand U24940 (N_24940,N_17255,N_19172);
or U24941 (N_24941,N_17704,N_16879);
or U24942 (N_24942,N_19708,N_18370);
nor U24943 (N_24943,N_16686,N_18993);
or U24944 (N_24944,N_16810,N_16287);
or U24945 (N_24945,N_16674,N_16215);
nand U24946 (N_24946,N_17933,N_16951);
xnor U24947 (N_24947,N_18001,N_17503);
and U24948 (N_24948,N_16109,N_17349);
or U24949 (N_24949,N_19185,N_18582);
nand U24950 (N_24950,N_15810,N_17682);
nand U24951 (N_24951,N_15081,N_18173);
nor U24952 (N_24952,N_16483,N_16681);
or U24953 (N_24953,N_17070,N_18127);
and U24954 (N_24954,N_16451,N_19258);
nor U24955 (N_24955,N_17642,N_16286);
or U24956 (N_24956,N_15459,N_17804);
nand U24957 (N_24957,N_17473,N_17618);
xnor U24958 (N_24958,N_17430,N_18198);
or U24959 (N_24959,N_17078,N_18417);
or U24960 (N_24960,N_15954,N_17893);
or U24961 (N_24961,N_15065,N_17889);
xnor U24962 (N_24962,N_15200,N_15856);
xnor U24963 (N_24963,N_16624,N_15761);
or U24964 (N_24964,N_16363,N_15429);
or U24965 (N_24965,N_19374,N_17490);
and U24966 (N_24966,N_15529,N_16734);
and U24967 (N_24967,N_18945,N_18468);
and U24968 (N_24968,N_15957,N_16979);
nand U24969 (N_24969,N_17452,N_17445);
nor U24970 (N_24970,N_15770,N_15557);
nand U24971 (N_24971,N_17983,N_15123);
nor U24972 (N_24972,N_17547,N_17049);
and U24973 (N_24973,N_19327,N_16749);
xnor U24974 (N_24974,N_18251,N_17614);
or U24975 (N_24975,N_17677,N_19915);
or U24976 (N_24976,N_15038,N_19319);
or U24977 (N_24977,N_15908,N_17610);
and U24978 (N_24978,N_17354,N_16248);
nor U24979 (N_24979,N_19181,N_17700);
nand U24980 (N_24980,N_19800,N_18234);
nand U24981 (N_24981,N_16578,N_18734);
xor U24982 (N_24982,N_16850,N_19706);
or U24983 (N_24983,N_18037,N_19612);
nor U24984 (N_24984,N_16698,N_19133);
nand U24985 (N_24985,N_19150,N_17408);
xor U24986 (N_24986,N_17922,N_19873);
nand U24987 (N_24987,N_16968,N_16439);
xnor U24988 (N_24988,N_19966,N_18002);
xnor U24989 (N_24989,N_16852,N_18364);
nor U24990 (N_24990,N_19964,N_19177);
xor U24991 (N_24991,N_16188,N_19788);
xor U24992 (N_24992,N_18896,N_16393);
or U24993 (N_24993,N_16240,N_16431);
nand U24994 (N_24994,N_15665,N_15788);
nor U24995 (N_24995,N_15122,N_15279);
nand U24996 (N_24996,N_17727,N_18378);
nor U24997 (N_24997,N_15628,N_17358);
nor U24998 (N_24998,N_19808,N_15152);
nor U24999 (N_24999,N_15098,N_19892);
xor U25000 (N_25000,N_21814,N_22714);
xor U25001 (N_25001,N_23917,N_20457);
nor U25002 (N_25002,N_22706,N_22869);
and U25003 (N_25003,N_21025,N_20239);
xor U25004 (N_25004,N_24759,N_21277);
nand U25005 (N_25005,N_24272,N_24020);
or U25006 (N_25006,N_22722,N_22106);
and U25007 (N_25007,N_22801,N_21927);
xnor U25008 (N_25008,N_22710,N_21709);
xnor U25009 (N_25009,N_23550,N_21650);
nand U25010 (N_25010,N_20308,N_22316);
and U25011 (N_25011,N_20458,N_24063);
nor U25012 (N_25012,N_21447,N_21380);
or U25013 (N_25013,N_22118,N_24531);
and U25014 (N_25014,N_22837,N_24089);
or U25015 (N_25015,N_22280,N_21680);
nor U25016 (N_25016,N_22324,N_22450);
and U25017 (N_25017,N_23473,N_23920);
or U25018 (N_25018,N_21142,N_21971);
nand U25019 (N_25019,N_24659,N_21410);
or U25020 (N_25020,N_22603,N_22043);
nand U25021 (N_25021,N_22920,N_22124);
or U25022 (N_25022,N_23266,N_24849);
and U25023 (N_25023,N_21768,N_21887);
nor U25024 (N_25024,N_22519,N_20611);
xnor U25025 (N_25025,N_20718,N_20861);
or U25026 (N_25026,N_21018,N_22277);
and U25027 (N_25027,N_21071,N_21822);
xor U25028 (N_25028,N_23400,N_23648);
xnor U25029 (N_25029,N_22535,N_24707);
xor U25030 (N_25030,N_23376,N_22857);
nor U25031 (N_25031,N_23560,N_22653);
nor U25032 (N_25032,N_20035,N_21537);
nand U25033 (N_25033,N_24958,N_21304);
xnor U25034 (N_25034,N_21500,N_20778);
and U25035 (N_25035,N_21905,N_22629);
or U25036 (N_25036,N_22851,N_22625);
nand U25037 (N_25037,N_23398,N_24794);
nand U25038 (N_25038,N_21098,N_22744);
nor U25039 (N_25039,N_23537,N_23849);
nand U25040 (N_25040,N_24597,N_20670);
xnor U25041 (N_25041,N_23261,N_23252);
nor U25042 (N_25042,N_21384,N_20031);
and U25043 (N_25043,N_20836,N_21212);
nor U25044 (N_25044,N_20801,N_21674);
xnor U25045 (N_25045,N_21843,N_22012);
and U25046 (N_25046,N_24986,N_24665);
nand U25047 (N_25047,N_22850,N_21378);
and U25048 (N_25048,N_24835,N_22594);
and U25049 (N_25049,N_20533,N_24596);
or U25050 (N_25050,N_21206,N_24140);
and U25051 (N_25051,N_23782,N_20513);
xnor U25052 (N_25052,N_23324,N_20311);
and U25053 (N_25053,N_24099,N_21051);
xnor U25054 (N_25054,N_21610,N_23511);
nand U25055 (N_25055,N_22331,N_20994);
xnor U25056 (N_25056,N_24719,N_23612);
xnor U25057 (N_25057,N_21309,N_20580);
nand U25058 (N_25058,N_22478,N_22941);
or U25059 (N_25059,N_24054,N_24810);
nor U25060 (N_25060,N_24534,N_20640);
xnor U25061 (N_25061,N_24834,N_21186);
nor U25062 (N_25062,N_24677,N_20905);
nor U25063 (N_25063,N_22160,N_23978);
nand U25064 (N_25064,N_22269,N_23658);
nor U25065 (N_25065,N_21232,N_24329);
and U25066 (N_25066,N_20741,N_21816);
nand U25067 (N_25067,N_22254,N_22188);
nor U25068 (N_25068,N_21871,N_24942);
and U25069 (N_25069,N_22723,N_23864);
and U25070 (N_25070,N_23565,N_22825);
nand U25071 (N_25071,N_21376,N_24287);
or U25072 (N_25072,N_24268,N_24177);
nor U25073 (N_25073,N_22439,N_24578);
nor U25074 (N_25074,N_23726,N_20983);
nand U25075 (N_25075,N_21823,N_20333);
nor U25076 (N_25076,N_20250,N_21247);
nor U25077 (N_25077,N_21434,N_22695);
xor U25078 (N_25078,N_23985,N_22991);
and U25079 (N_25079,N_21169,N_23772);
nor U25080 (N_25080,N_21008,N_21925);
nor U25081 (N_25081,N_24302,N_20438);
xor U25082 (N_25082,N_24495,N_20134);
and U25083 (N_25083,N_24483,N_20405);
nor U25084 (N_25084,N_20667,N_22334);
or U25085 (N_25085,N_20970,N_24060);
nor U25086 (N_25086,N_22746,N_24565);
nor U25087 (N_25087,N_21585,N_23556);
or U25088 (N_25088,N_20751,N_24740);
or U25089 (N_25089,N_20930,N_23620);
or U25090 (N_25090,N_20017,N_21466);
or U25091 (N_25091,N_21526,N_20747);
nor U25092 (N_25092,N_21554,N_20233);
nand U25093 (N_25093,N_22033,N_22698);
and U25094 (N_25094,N_24783,N_24172);
nor U25095 (N_25095,N_24622,N_24925);
xor U25096 (N_25096,N_21416,N_21483);
and U25097 (N_25097,N_24240,N_24066);
or U25098 (N_25098,N_22347,N_20633);
or U25099 (N_25099,N_22376,N_24123);
or U25100 (N_25100,N_22965,N_21584);
xor U25101 (N_25101,N_23490,N_20610);
nand U25102 (N_25102,N_21108,N_24160);
and U25103 (N_25103,N_24785,N_21937);
nor U25104 (N_25104,N_23545,N_21441);
nand U25105 (N_25105,N_20025,N_23755);
and U25106 (N_25106,N_21245,N_21326);
or U25107 (N_25107,N_22025,N_22247);
and U25108 (N_25108,N_20617,N_23967);
nor U25109 (N_25109,N_23571,N_23223);
nor U25110 (N_25110,N_24638,N_20829);
nand U25111 (N_25111,N_23224,N_23016);
or U25112 (N_25112,N_22844,N_23646);
nor U25113 (N_25113,N_21781,N_22226);
xor U25114 (N_25114,N_24460,N_20126);
xor U25115 (N_25115,N_24344,N_20051);
nand U25116 (N_25116,N_22552,N_20286);
and U25117 (N_25117,N_24148,N_20204);
or U25118 (N_25118,N_23168,N_21015);
nand U25119 (N_25119,N_20365,N_22630);
xor U25120 (N_25120,N_24498,N_22285);
or U25121 (N_25121,N_20603,N_20103);
or U25122 (N_25122,N_23035,N_24038);
or U25123 (N_25123,N_20814,N_24936);
nand U25124 (N_25124,N_20061,N_20429);
nand U25125 (N_25125,N_22125,N_24350);
nor U25126 (N_25126,N_21553,N_20024);
or U25127 (N_25127,N_23981,N_23825);
nor U25128 (N_25128,N_21168,N_23554);
or U25129 (N_25129,N_23691,N_23315);
nand U25130 (N_25130,N_22266,N_24386);
nor U25131 (N_25131,N_22211,N_20472);
and U25132 (N_25132,N_24396,N_23057);
nand U25133 (N_25133,N_24918,N_24203);
or U25134 (N_25134,N_22335,N_21749);
nor U25135 (N_25135,N_24647,N_22894);
xor U25136 (N_25136,N_23583,N_20595);
and U25137 (N_25137,N_22243,N_20825);
nor U25138 (N_25138,N_24171,N_21643);
nand U25139 (N_25139,N_22515,N_24481);
nor U25140 (N_25140,N_23444,N_23258);
nand U25141 (N_25141,N_23445,N_22527);
and U25142 (N_25142,N_24086,N_21608);
or U25143 (N_25143,N_20892,N_20172);
and U25144 (N_25144,N_22927,N_20109);
nand U25145 (N_25145,N_22231,N_23197);
nand U25146 (N_25146,N_24455,N_24157);
nor U25147 (N_25147,N_22040,N_21191);
nor U25148 (N_25148,N_22422,N_23474);
or U25149 (N_25149,N_21923,N_24778);
nor U25150 (N_25150,N_24652,N_22871);
nor U25151 (N_25151,N_23683,N_24011);
and U25152 (N_25152,N_20244,N_20809);
or U25153 (N_25153,N_23878,N_21954);
xor U25154 (N_25154,N_22901,N_22789);
nor U25155 (N_25155,N_21300,N_20171);
and U25156 (N_25156,N_22907,N_20090);
xor U25157 (N_25157,N_20374,N_20556);
and U25158 (N_25158,N_20482,N_24017);
and U25159 (N_25159,N_20433,N_20887);
xor U25160 (N_25160,N_22974,N_22141);
or U25161 (N_25161,N_24681,N_22464);
nand U25162 (N_25162,N_23955,N_23428);
nand U25163 (N_25163,N_24933,N_23267);
xnor U25164 (N_25164,N_22893,N_24446);
nand U25165 (N_25165,N_21528,N_24018);
xor U25166 (N_25166,N_23800,N_22109);
and U25167 (N_25167,N_23734,N_24121);
xnor U25168 (N_25168,N_23065,N_21227);
xor U25169 (N_25169,N_20010,N_20692);
nor U25170 (N_25170,N_22967,N_21053);
or U25171 (N_25171,N_24322,N_23017);
xor U25172 (N_25172,N_21510,N_24723);
or U25173 (N_25173,N_21269,N_20310);
and U25174 (N_25174,N_20476,N_23356);
xnor U25175 (N_25175,N_23650,N_24658);
xor U25176 (N_25176,N_24855,N_22639);
or U25177 (N_25177,N_22836,N_20424);
and U25178 (N_25178,N_22501,N_23941);
and U25179 (N_25179,N_23729,N_20454);
xor U25180 (N_25180,N_24953,N_20373);
nor U25181 (N_25181,N_21884,N_20349);
nand U25182 (N_25182,N_24644,N_22312);
or U25183 (N_25183,N_20984,N_24155);
and U25184 (N_25184,N_22808,N_21173);
nor U25185 (N_25185,N_22624,N_23368);
nand U25186 (N_25186,N_24758,N_23636);
and U25187 (N_25187,N_24765,N_22129);
nor U25188 (N_25188,N_21022,N_23340);
xor U25189 (N_25189,N_22088,N_21363);
nand U25190 (N_25190,N_24726,N_21448);
nor U25191 (N_25191,N_21215,N_21599);
nor U25192 (N_25192,N_21963,N_21698);
xor U25193 (N_25193,N_22453,N_22687);
or U25194 (N_25194,N_20128,N_24634);
nand U25195 (N_25195,N_24375,N_22516);
nand U25196 (N_25196,N_23738,N_22561);
nor U25197 (N_25197,N_20862,N_22089);
xor U25198 (N_25198,N_23670,N_21061);
xor U25199 (N_25199,N_22015,N_22896);
xnor U25200 (N_25200,N_21980,N_22949);
and U25201 (N_25201,N_23641,N_24290);
xnor U25202 (N_25202,N_23750,N_20135);
nor U25203 (N_25203,N_23855,N_22742);
nor U25204 (N_25204,N_20679,N_22934);
and U25205 (N_25205,N_22326,N_23821);
xor U25206 (N_25206,N_23847,N_21714);
nand U25207 (N_25207,N_21032,N_23325);
nand U25208 (N_25208,N_24892,N_23260);
nand U25209 (N_25209,N_21427,N_20860);
and U25210 (N_25210,N_21214,N_24540);
xnor U25211 (N_25211,N_23411,N_22018);
xor U25212 (N_25212,N_24997,N_23723);
or U25213 (N_25213,N_23532,N_22470);
and U25214 (N_25214,N_24888,N_21989);
xnor U25215 (N_25215,N_21868,N_22532);
nor U25216 (N_25216,N_22599,N_21837);
xnor U25217 (N_25217,N_24052,N_22740);
nand U25218 (N_25218,N_23719,N_20947);
nor U25219 (N_25219,N_21414,N_22657);
and U25220 (N_25220,N_21952,N_23054);
nand U25221 (N_25221,N_23921,N_20148);
and U25222 (N_25222,N_22251,N_23627);
and U25223 (N_25223,N_23533,N_20832);
nand U25224 (N_25224,N_23517,N_22217);
xnor U25225 (N_25225,N_22774,N_22474);
or U25226 (N_25226,N_22842,N_21290);
nor U25227 (N_25227,N_24722,N_21660);
nor U25228 (N_25228,N_20332,N_22578);
xor U25229 (N_25229,N_20839,N_20895);
nor U25230 (N_25230,N_23024,N_22606);
nand U25231 (N_25231,N_21405,N_20125);
xor U25232 (N_25232,N_20587,N_23333);
and U25233 (N_25233,N_24238,N_20541);
nor U25234 (N_25234,N_23006,N_24489);
xor U25235 (N_25235,N_21847,N_24232);
nand U25236 (N_25236,N_22708,N_20315);
xor U25237 (N_25237,N_23581,N_20655);
nand U25238 (N_25238,N_22405,N_21628);
or U25239 (N_25239,N_20978,N_21502);
nand U25240 (N_25240,N_23746,N_23048);
nand U25241 (N_25241,N_23283,N_23875);
nor U25242 (N_25242,N_20437,N_24575);
and U25243 (N_25243,N_21170,N_21237);
nand U25244 (N_25244,N_20156,N_21175);
xor U25245 (N_25245,N_20394,N_23924);
nor U25246 (N_25246,N_20601,N_21785);
nor U25247 (N_25247,N_24382,N_20030);
xnor U25248 (N_25248,N_24249,N_23322);
and U25249 (N_25249,N_22411,N_23709);
xor U25250 (N_25250,N_20948,N_20276);
xor U25251 (N_25251,N_21524,N_23991);
and U25252 (N_25252,N_22446,N_24390);
and U25253 (N_25253,N_23044,N_21469);
or U25254 (N_25254,N_21347,N_22737);
or U25255 (N_25255,N_22323,N_23704);
nor U25256 (N_25256,N_24971,N_20515);
xor U25257 (N_25257,N_23766,N_24105);
nand U25258 (N_25258,N_23874,N_23822);
and U25259 (N_25259,N_22973,N_21161);
nand U25260 (N_25260,N_23562,N_21476);
or U25261 (N_25261,N_24860,N_21338);
or U25262 (N_25262,N_20530,N_21836);
and U25263 (N_25263,N_23568,N_23736);
xor U25264 (N_25264,N_21240,N_23717);
nor U25265 (N_25265,N_20672,N_23809);
or U25266 (N_25266,N_24893,N_23475);
or U25267 (N_25267,N_20511,N_20431);
nor U25268 (N_25268,N_21747,N_24970);
xnor U25269 (N_25269,N_24560,N_24229);
nor U25270 (N_25270,N_20184,N_24278);
nor U25271 (N_25271,N_22843,N_23856);
or U25272 (N_25272,N_24899,N_22272);
xnor U25273 (N_25273,N_22403,N_22418);
nand U25274 (N_25274,N_21332,N_23367);
nand U25275 (N_25275,N_24323,N_22220);
and U25276 (N_25276,N_23536,N_24225);
xor U25277 (N_25277,N_21374,N_22267);
or U25278 (N_25278,N_24605,N_24433);
and U25279 (N_25279,N_22371,N_20053);
nor U25280 (N_25280,N_23391,N_23314);
nand U25281 (N_25281,N_22457,N_20188);
nor U25282 (N_25282,N_22385,N_24732);
nor U25283 (N_25283,N_21083,N_23910);
xnor U25284 (N_25284,N_20988,N_23229);
and U25285 (N_25285,N_23876,N_23817);
and U25286 (N_25286,N_24512,N_21146);
or U25287 (N_25287,N_23507,N_20823);
nor U25288 (N_25288,N_22972,N_23089);
xnor U25289 (N_25289,N_23799,N_21305);
xor U25290 (N_25290,N_24820,N_24844);
xor U25291 (N_25291,N_21393,N_22486);
xnor U25292 (N_25292,N_21220,N_23169);
or U25293 (N_25293,N_23491,N_21885);
nand U25294 (N_25294,N_24984,N_24371);
xnor U25295 (N_25295,N_23622,N_20935);
and U25296 (N_25296,N_22374,N_24516);
nand U25297 (N_25297,N_20414,N_23965);
xnor U25298 (N_25298,N_22423,N_24248);
nand U25299 (N_25299,N_24084,N_21404);
xor U25300 (N_25300,N_23128,N_23175);
or U25301 (N_25301,N_22039,N_21111);
and U25302 (N_25302,N_21830,N_22438);
or U25303 (N_25303,N_23439,N_22554);
nand U25304 (N_25304,N_20651,N_22623);
nor U25305 (N_25305,N_22948,N_24866);
and U25306 (N_25306,N_24198,N_21174);
xor U25307 (N_25307,N_22985,N_20499);
nand U25308 (N_25308,N_20281,N_20616);
xor U25309 (N_25309,N_22028,N_21713);
or U25310 (N_25310,N_24989,N_21199);
and U25311 (N_25311,N_20168,N_20083);
nor U25312 (N_25312,N_20466,N_22381);
nand U25313 (N_25313,N_21738,N_24030);
xor U25314 (N_25314,N_24028,N_21361);
nor U25315 (N_25315,N_24760,N_20115);
nand U25316 (N_25316,N_22301,N_20052);
and U25317 (N_25317,N_20650,N_20579);
and U25318 (N_25318,N_22484,N_20399);
nand U25319 (N_25319,N_21895,N_20789);
xor U25320 (N_25320,N_24280,N_21387);
nor U25321 (N_25321,N_24208,N_24064);
nor U25322 (N_25322,N_22051,N_23587);
xnor U25323 (N_25323,N_20737,N_23841);
xor U25324 (N_25324,N_20625,N_21773);
and U25325 (N_25325,N_23030,N_22036);
xnor U25326 (N_25326,N_22279,N_23180);
nand U25327 (N_25327,N_20242,N_24782);
xor U25328 (N_25328,N_20910,N_24956);
or U25329 (N_25329,N_20527,N_23541);
nand U25330 (N_25330,N_22747,N_22739);
nand U25331 (N_25331,N_24475,N_24050);
xor U25332 (N_25332,N_23603,N_22310);
nand U25333 (N_25333,N_24318,N_22077);
nand U25334 (N_25334,N_21348,N_20422);
nand U25335 (N_25335,N_24439,N_22490);
xor U25336 (N_25336,N_22196,N_23238);
nor U25337 (N_25337,N_23932,N_21866);
nand U25338 (N_25338,N_24803,N_21634);
nor U25339 (N_25339,N_22754,N_22890);
or U25340 (N_25340,N_20879,N_24391);
xor U25341 (N_25341,N_24643,N_24562);
and U25342 (N_25342,N_20340,N_21438);
nand U25343 (N_25343,N_22148,N_21828);
and U25344 (N_25344,N_21499,N_20954);
nand U25345 (N_25345,N_24167,N_24563);
and U25346 (N_25346,N_23707,N_23940);
nor U25347 (N_25347,N_22178,N_24828);
xnor U25348 (N_25348,N_21110,N_20305);
xor U25349 (N_25349,N_20914,N_22105);
nand U25350 (N_25350,N_24853,N_23538);
or U25351 (N_25351,N_21433,N_23903);
nor U25352 (N_25352,N_20802,N_21021);
nor U25353 (N_25353,N_23547,N_20881);
xor U25354 (N_25354,N_20137,N_21360);
nand U25355 (N_25355,N_21944,N_21473);
nand U25356 (N_25356,N_23961,N_21330);
nor U25357 (N_25357,N_24742,N_24372);
nor U25358 (N_25358,N_23988,N_21957);
nor U25359 (N_25359,N_23975,N_20059);
nor U25360 (N_25360,N_20312,N_24246);
xor U25361 (N_25361,N_20254,N_21693);
and U25362 (N_25362,N_23983,N_22047);
or U25363 (N_25363,N_20612,N_20868);
xor U25364 (N_25364,N_24134,N_22509);
nand U25365 (N_25365,N_21057,N_24113);
nor U25366 (N_25366,N_24291,N_23412);
xor U25367 (N_25367,N_20641,N_22875);
nand U25368 (N_25368,N_22539,N_23773);
and U25369 (N_25369,N_20195,N_23243);
nand U25370 (N_25370,N_24370,N_23335);
xor U25371 (N_25371,N_20409,N_23640);
and U25372 (N_25372,N_23501,N_22265);
nor U25373 (N_25373,N_21106,N_21182);
or U25374 (N_25374,N_20506,N_24403);
nand U25375 (N_25375,N_22669,N_21266);
and U25376 (N_25376,N_23743,N_20807);
and U25377 (N_25377,N_22407,N_21196);
and U25378 (N_25378,N_23497,N_22868);
or U25379 (N_25379,N_22465,N_22780);
nand U25380 (N_25380,N_21088,N_23804);
nor U25381 (N_25381,N_23403,N_22919);
nand U25382 (N_25382,N_24425,N_23850);
or U25383 (N_25383,N_22170,N_21664);
nor U25384 (N_25384,N_20341,N_23278);
and U25385 (N_25385,N_24027,N_22971);
nor U25386 (N_25386,N_21800,N_20943);
nor U25387 (N_25387,N_23344,N_22664);
xnor U25388 (N_25388,N_21243,N_22066);
or U25389 (N_25389,N_23796,N_23482);
or U25390 (N_25390,N_22117,N_21334);
and U25391 (N_25391,N_20371,N_22344);
and U25392 (N_25392,N_23279,N_21398);
nand U25393 (N_25393,N_24960,N_23112);
nor U25394 (N_25394,N_24006,N_24222);
xor U25395 (N_25395,N_20992,N_22946);
and U25396 (N_25396,N_21964,N_22019);
or U25397 (N_25397,N_24195,N_21236);
nor U25398 (N_25398,N_22963,N_21246);
and U25399 (N_25399,N_21419,N_24144);
or U25400 (N_25400,N_24436,N_21718);
or U25401 (N_25401,N_23381,N_20039);
and U25402 (N_25402,N_22727,N_24388);
or U25403 (N_25403,N_20143,N_20926);
and U25404 (N_25404,N_21350,N_23594);
and U25405 (N_25405,N_20937,N_24270);
or U25406 (N_25406,N_21565,N_21546);
nand U25407 (N_25407,N_21997,N_22879);
xnor U25408 (N_25408,N_20800,N_23184);
nor U25409 (N_25409,N_24260,N_24093);
and U25410 (N_25410,N_23639,N_22618);
nor U25411 (N_25411,N_24932,N_21582);
and U25412 (N_25412,N_24341,N_24947);
xor U25413 (N_25413,N_21415,N_23787);
or U25414 (N_25414,N_24902,N_24786);
nor U25415 (N_25415,N_21623,N_21904);
nand U25416 (N_25416,N_24231,N_20586);
nand U25417 (N_25417,N_21225,N_24915);
and U25418 (N_25418,N_20798,N_23710);
or U25419 (N_25419,N_23461,N_23610);
xor U25420 (N_25420,N_22565,N_24669);
and U25421 (N_25421,N_20222,N_21624);
and U25422 (N_25422,N_21813,N_23564);
xnor U25423 (N_25423,N_20484,N_20263);
and U25424 (N_25424,N_22736,N_22139);
xor U25425 (N_25425,N_23759,N_21055);
nor U25426 (N_25426,N_22577,N_22512);
nand U25427 (N_25427,N_24750,N_23775);
and U25428 (N_25428,N_21936,N_22122);
nor U25429 (N_25429,N_22998,N_24474);
or U25430 (N_25430,N_21996,N_20289);
xnor U25431 (N_25431,N_22293,N_23867);
nand U25432 (N_25432,N_21189,N_20744);
nand U25433 (N_25433,N_20664,N_21226);
nand U25434 (N_25434,N_23761,N_23840);
nand U25435 (N_25435,N_21038,N_22800);
and U25436 (N_25436,N_22839,N_23202);
xor U25437 (N_25437,N_23588,N_22962);
xor U25438 (N_25438,N_21986,N_20119);
xor U25439 (N_25439,N_22969,N_23740);
xnor U25440 (N_25440,N_20569,N_22360);
xor U25441 (N_25441,N_22341,N_21221);
xor U25442 (N_25442,N_20848,N_21981);
or U25443 (N_25443,N_23392,N_24022);
or U25444 (N_25444,N_21757,N_22818);
xor U25445 (N_25445,N_20081,N_21133);
nand U25446 (N_25446,N_22976,N_23050);
and U25447 (N_25447,N_20346,N_23606);
or U25448 (N_25448,N_21732,N_23320);
and U25449 (N_25449,N_23259,N_23575);
nand U25450 (N_25450,N_21876,N_20058);
or U25451 (N_25451,N_23797,N_21459);
nor U25452 (N_25452,N_23093,N_23369);
xnor U25453 (N_25453,N_21481,N_24126);
and U25454 (N_25454,N_24791,N_21708);
xnor U25455 (N_25455,N_20336,N_20658);
nand U25456 (N_25456,N_22716,N_23601);
nand U25457 (N_25457,N_22302,N_22154);
or U25458 (N_25458,N_20563,N_20562);
nor U25459 (N_25459,N_24746,N_22074);
nand U25460 (N_25460,N_21091,N_24935);
xnor U25461 (N_25461,N_22044,N_23366);
nand U25462 (N_25462,N_23156,N_22617);
and U25463 (N_25463,N_21203,N_22147);
or U25464 (N_25464,N_20451,N_23115);
or U25465 (N_25465,N_22573,N_23069);
and U25466 (N_25466,N_20334,N_22298);
nand U25467 (N_25467,N_21178,N_22169);
nand U25468 (N_25468,N_22270,N_23330);
xor U25469 (N_25469,N_20283,N_20260);
and U25470 (N_25470,N_20094,N_21292);
and U25471 (N_25471,N_23861,N_20567);
xor U25472 (N_25472,N_21854,N_22460);
nand U25473 (N_25473,N_23768,N_24704);
or U25474 (N_25474,N_24200,N_21820);
and U25475 (N_25475,N_21257,N_24158);
and U25476 (N_25476,N_23883,N_23264);
nand U25477 (N_25477,N_24470,N_23929);
nor U25478 (N_25478,N_23793,N_23968);
nand U25479 (N_25479,N_22305,N_23012);
or U25480 (N_25480,N_22820,N_23508);
or U25481 (N_25481,N_22441,N_22770);
nor U25482 (N_25482,N_23590,N_23306);
nor U25483 (N_25483,N_23938,N_20478);
nand U25484 (N_25484,N_23879,N_21297);
xnor U25485 (N_25485,N_20342,N_20459);
and U25486 (N_25486,N_23725,N_20318);
xor U25487 (N_25487,N_20036,N_22050);
xor U25488 (N_25488,N_22583,N_20764);
nand U25489 (N_25489,N_20291,N_21670);
and U25490 (N_25490,N_21355,N_22321);
xor U25491 (N_25491,N_21548,N_21857);
or U25492 (N_25492,N_22416,N_22459);
and U25493 (N_25493,N_22127,N_23698);
and U25494 (N_25494,N_23614,N_20114);
or U25495 (N_25495,N_24021,N_21922);
nor U25496 (N_25496,N_20867,N_23798);
nand U25497 (N_25497,N_22549,N_22612);
nand U25498 (N_25498,N_22317,N_20497);
xnor U25499 (N_25499,N_22114,N_21990);
and U25500 (N_25500,N_24003,N_23268);
or U25501 (N_25501,N_22156,N_22913);
xnor U25502 (N_25502,N_24812,N_22646);
or U25503 (N_25503,N_20956,N_21569);
xor U25504 (N_25504,N_21171,N_21901);
nor U25505 (N_25505,N_22887,N_22725);
nor U25506 (N_25506,N_24295,N_24747);
and U25507 (N_25507,N_23770,N_23074);
nor U25508 (N_25508,N_22576,N_21354);
nor U25509 (N_25509,N_20535,N_24537);
nand U25510 (N_25510,N_24908,N_20712);
and U25511 (N_25511,N_22795,N_23728);
and U25512 (N_25512,N_22046,N_22707);
or U25513 (N_25513,N_24987,N_21275);
and U25514 (N_25514,N_21331,N_21933);
or U25515 (N_25515,N_20526,N_21557);
nor U25516 (N_25516,N_23312,N_22308);
nand U25517 (N_25517,N_23808,N_20547);
nand U25518 (N_25518,N_20982,N_23617);
and U25519 (N_25519,N_22174,N_20415);
and U25520 (N_25520,N_20357,N_20834);
nand U25521 (N_25521,N_20996,N_24642);
nand U25522 (N_25522,N_23346,N_23352);
xnor U25523 (N_25523,N_23302,N_24090);
nand U25524 (N_25524,N_23853,N_24657);
and U25525 (N_25525,N_20685,N_20668);
and U25526 (N_25526,N_20054,N_23980);
nand U25527 (N_25527,N_22982,N_22332);
and U25528 (N_25528,N_24503,N_20411);
nor U25529 (N_25529,N_22604,N_24939);
nand U25530 (N_25530,N_21293,N_22437);
and U25531 (N_25531,N_21181,N_22236);
nand U25532 (N_25532,N_21163,N_22327);
xor U25533 (N_25533,N_23466,N_24887);
nand U25534 (N_25534,N_24805,N_20001);
and U25535 (N_25535,N_20656,N_24550);
xnor U25536 (N_25536,N_21042,N_23173);
xor U25537 (N_25537,N_21728,N_20042);
or U25538 (N_25538,N_21609,N_21003);
or U25539 (N_25539,N_23845,N_21946);
xnor U25540 (N_25540,N_24694,N_20161);
xnor U25541 (N_25541,N_23724,N_24507);
and U25542 (N_25542,N_23890,N_24755);
or U25543 (N_25543,N_23582,N_22677);
and U25544 (N_25544,N_24088,N_21470);
xnor U25545 (N_25545,N_22208,N_24827);
and U25546 (N_25546,N_21529,N_24409);
nand U25547 (N_25547,N_23711,N_21615);
xor U25548 (N_25548,N_24176,N_21219);
nand U25549 (N_25549,N_20124,N_21908);
nor U25550 (N_25550,N_21043,N_21748);
nor U25551 (N_25551,N_22675,N_24532);
nor U25552 (N_25552,N_24948,N_20091);
xnor U25553 (N_25553,N_20756,N_20863);
and U25554 (N_25554,N_21894,N_21652);
and U25555 (N_25555,N_23913,N_24153);
or U25556 (N_25556,N_24502,N_23986);
or U25557 (N_25557,N_23481,N_21037);
xor U25558 (N_25558,N_21035,N_20331);
xnor U25559 (N_25559,N_21085,N_21468);
nor U25560 (N_25560,N_24648,N_21112);
or U25561 (N_25561,N_20991,N_20470);
nor U25562 (N_25562,N_21618,N_20966);
and U25563 (N_25563,N_22702,N_22398);
or U25564 (N_25564,N_21806,N_22020);
or U25565 (N_25565,N_21251,N_24656);
and U25566 (N_25566,N_21479,N_20316);
or U25567 (N_25567,N_24944,N_22100);
nand U25568 (N_25568,N_23483,N_20518);
xor U25569 (N_25569,N_23029,N_21155);
or U25570 (N_25570,N_22116,N_20037);
nor U25571 (N_25571,N_23801,N_23962);
and U25572 (N_25572,N_21048,N_24991);
nor U25573 (N_25573,N_23688,N_22921);
nor U25574 (N_25574,N_20849,N_23101);
or U25575 (N_25575,N_22362,N_22348);
and U25576 (N_25576,N_24300,N_20776);
and U25577 (N_25577,N_24445,N_24818);
or U25578 (N_25578,N_23751,N_22026);
or U25579 (N_25579,N_24243,N_23553);
nor U25580 (N_25580,N_24301,N_21033);
nand U25581 (N_25581,N_23270,N_24766);
or U25582 (N_25582,N_21289,N_20927);
nand U25583 (N_25583,N_20576,N_20696);
xnor U25584 (N_25584,N_22922,N_23457);
and U25585 (N_25585,N_24870,N_22977);
or U25586 (N_25586,N_24611,N_20642);
and U25587 (N_25587,N_22216,N_22654);
and U25588 (N_25588,N_23647,N_23731);
or U25589 (N_25589,N_20919,N_24588);
or U25590 (N_25590,N_21924,N_20245);
xor U25591 (N_25591,N_21764,N_24600);
nand U25592 (N_25592,N_22369,N_23129);
and U25593 (N_25593,N_21123,N_23385);
and U25594 (N_25594,N_23928,N_22882);
and U25595 (N_25595,N_22522,N_23332);
or U25596 (N_25596,N_20716,N_20898);
and U25597 (N_25597,N_20503,N_22511);
and U25598 (N_25598,N_24245,N_23659);
or U25599 (N_25599,N_21795,N_22417);
nor U25600 (N_25600,N_21741,N_22158);
nand U25601 (N_25601,N_24864,N_24762);
nor U25602 (N_25602,N_21667,N_20510);
or U25603 (N_25603,N_22180,N_20504);
nor U25604 (N_25604,N_23014,N_23769);
or U25605 (N_25605,N_24809,N_24352);
and U25606 (N_25606,N_22093,N_23702);
and U25607 (N_25607,N_22759,N_20682);
xor U25608 (N_25608,N_21322,N_24062);
nor U25609 (N_25609,N_23301,N_22872);
or U25610 (N_25610,N_23685,N_24883);
nand U25611 (N_25611,N_20969,N_20133);
nand U25612 (N_25612,N_24954,N_20469);
and U25613 (N_25613,N_24161,N_24992);
nor U25614 (N_25614,N_21004,N_24836);
or U25615 (N_25615,N_20181,N_21783);
nand U25616 (N_25616,N_24488,N_22286);
and U25617 (N_25617,N_20072,N_21518);
nor U25618 (N_25618,N_22908,N_21377);
and U25619 (N_25619,N_21559,N_24367);
nor U25620 (N_25620,N_24660,N_20977);
or U25621 (N_25621,N_24538,N_24718);
and U25622 (N_25622,N_22526,N_24389);
nor U25623 (N_25623,N_22479,N_20099);
and U25624 (N_25624,N_23739,N_22111);
and U25625 (N_25625,N_22847,N_22250);
nand U25626 (N_25626,N_22673,N_21394);
nor U25627 (N_25627,N_20906,N_23071);
nand U25628 (N_25628,N_20453,N_21756);
or U25629 (N_25629,N_24102,N_24206);
and U25630 (N_25630,N_20840,N_21262);
nor U25631 (N_25631,N_24598,N_22809);
or U25632 (N_25632,N_22543,N_21023);
xor U25633 (N_25633,N_23790,N_23831);
or U25634 (N_25634,N_20217,N_23189);
nand U25635 (N_25635,N_21725,N_20649);
and U25636 (N_25636,N_22199,N_22935);
or U25637 (N_25637,N_22113,N_22057);
xor U25638 (N_25638,N_23471,N_20273);
nor U25639 (N_25639,N_20767,N_24316);
nand U25640 (N_25640,N_21802,N_22658);
and U25641 (N_25641,N_24056,N_21019);
nand U25642 (N_25642,N_23441,N_20908);
nor U25643 (N_25643,N_24339,N_21832);
and U25644 (N_25644,N_20951,N_20752);
nor U25645 (N_25645,N_22002,N_22396);
nor U25646 (N_25646,N_21077,N_22469);
nor U25647 (N_25647,N_20043,N_22359);
xnor U25648 (N_25648,N_20669,N_24579);
nor U25649 (N_25649,N_20599,N_20304);
xnor U25650 (N_25650,N_21686,N_21515);
xor U25651 (N_25651,N_20174,N_21364);
nand U25652 (N_25652,N_23757,N_21397);
or U25653 (N_25653,N_24357,N_23188);
nand U25654 (N_25654,N_22567,N_24312);
and U25655 (N_25655,N_21060,N_22553);
or U25656 (N_25656,N_22413,N_21353);
nand U25657 (N_25657,N_24592,N_22585);
nor U25658 (N_25658,N_21150,N_23514);
nor U25659 (N_25659,N_20093,N_22004);
or U25660 (N_25660,N_21819,N_21829);
xnor U25661 (N_25661,N_20038,N_23254);
or U25662 (N_25662,N_24205,N_20266);
or U25663 (N_25663,N_22814,N_22504);
nor U25664 (N_25664,N_24504,N_20295);
and U25665 (N_25665,N_22692,N_22917);
xnor U25666 (N_25666,N_22775,N_21442);
nand U25667 (N_25667,N_21654,N_22961);
and U25668 (N_25668,N_22060,N_23105);
or U25669 (N_25669,N_23215,N_21918);
nand U25670 (N_25670,N_21786,N_21669);
xnor U25671 (N_25671,N_21159,N_24019);
xor U25672 (N_25672,N_23172,N_24146);
nand U25673 (N_25673,N_21792,N_23486);
nand U25674 (N_25674,N_24359,N_21064);
xor U25675 (N_25675,N_20366,N_22330);
nor U25676 (N_25676,N_20062,N_20225);
or U25677 (N_25677,N_22686,N_20153);
nand U25678 (N_25678,N_23205,N_23700);
nand U25679 (N_25679,N_24995,N_22500);
xor U25680 (N_25680,N_24983,N_24725);
nor U25681 (N_25681,N_20615,N_21835);
nand U25682 (N_25682,N_20465,N_21320);
nor U25683 (N_25683,N_21346,N_23321);
or U25684 (N_25684,N_23525,N_20452);
and U25685 (N_25685,N_21411,N_20362);
or U25686 (N_25686,N_20178,N_20824);
or U25687 (N_25687,N_23055,N_20939);
or U25688 (N_25688,N_23784,N_20775);
nor U25689 (N_25689,N_20613,N_21026);
or U25690 (N_25690,N_23811,N_22128);
xnor U25691 (N_25691,N_22001,N_23146);
and U25692 (N_25692,N_24497,N_24815);
and U25693 (N_25693,N_21633,N_24196);
xor U25694 (N_25694,N_20445,N_22239);
nor U25695 (N_25695,N_21097,N_22518);
or U25696 (N_25696,N_24826,N_22926);
nand U25697 (N_25697,N_24034,N_20901);
or U25698 (N_25698,N_23308,N_21272);
xnor U25699 (N_25699,N_23506,N_22131);
or U25700 (N_25700,N_23994,N_24002);
xnor U25701 (N_25701,N_20695,N_21535);
xor U25702 (N_25702,N_20117,N_22287);
and U25703 (N_25703,N_23298,N_20026);
nor U25704 (N_25704,N_23404,N_23025);
or U25705 (N_25705,N_22173,N_22670);
nor U25706 (N_25706,N_20076,N_21794);
and U25707 (N_25707,N_23122,N_22593);
or U25708 (N_25708,N_20750,N_22694);
nand U25709 (N_25709,N_22102,N_23294);
or U25710 (N_25710,N_24307,N_24686);
nor U25711 (N_25711,N_24116,N_21995);
and U25712 (N_25712,N_20661,N_24410);
xnor U25713 (N_25713,N_20997,N_21859);
or U25714 (N_25714,N_21817,N_20018);
nor U25715 (N_25715,N_21611,N_20732);
and U25716 (N_25716,N_22471,N_23679);
and U25717 (N_25717,N_20960,N_21367);
and U25718 (N_25718,N_21362,N_21551);
nor U25719 (N_25719,N_22990,N_24789);
xnor U25720 (N_25720,N_22943,N_21642);
nand U25721 (N_25721,N_21440,N_24679);
and U25722 (N_25722,N_22197,N_24649);
xnor U25723 (N_25723,N_21154,N_23531);
xnor U25724 (N_25724,N_20757,N_20151);
xnor U25725 (N_25725,N_23289,N_20296);
xor U25726 (N_25726,N_22333,N_21572);
nor U25727 (N_25727,N_22819,N_23791);
xor U25728 (N_25728,N_24071,N_24143);
xnor U25729 (N_25729,N_23274,N_21024);
nand U25730 (N_25730,N_24711,N_23785);
nor U25731 (N_25731,N_21271,N_24373);
nand U25732 (N_25732,N_21391,N_24639);
and U25733 (N_25733,N_20875,N_20121);
and U25734 (N_25734,N_23914,N_23415);
and U25735 (N_25735,N_21877,N_24548);
or U25736 (N_25736,N_24424,N_23815);
or U25737 (N_25737,N_20475,N_20558);
xnor U25738 (N_25738,N_20843,N_23781);
xnor U25739 (N_25739,N_22401,N_21103);
and U25740 (N_25740,N_21012,N_23378);
xor U25741 (N_25741,N_20327,N_24486);
and U25742 (N_25742,N_21640,N_24363);
and U25743 (N_25743,N_22276,N_21072);
xnor U25744 (N_25744,N_21530,N_23138);
or U25745 (N_25745,N_21325,N_23269);
or U25746 (N_25746,N_24241,N_24724);
or U25747 (N_25747,N_22906,N_24552);
or U25748 (N_25748,N_23083,N_21961);
or U25749 (N_25749,N_21465,N_22258);
or U25750 (N_25750,N_22099,N_24365);
xor U25751 (N_25751,N_23211,N_21166);
and U25752 (N_25752,N_22273,N_23094);
or U25753 (N_25753,N_21193,N_21917);
nor U25754 (N_25754,N_20955,N_20631);
nand U25755 (N_25755,N_21396,N_23563);
and U25756 (N_25756,N_22322,N_24910);
nor U25757 (N_25757,N_23179,N_24780);
xor U25758 (N_25758,N_21696,N_24476);
nand U25759 (N_25759,N_22354,N_20734);
or U25760 (N_25760,N_24361,N_20388);
nor U25761 (N_25761,N_20498,N_24982);
or U25762 (N_25762,N_23446,N_23618);
nor U25763 (N_25763,N_23680,N_24926);
xor U25764 (N_25764,N_21090,N_20360);
nor U25765 (N_25765,N_22107,N_20545);
xnor U25766 (N_25766,N_21216,N_24520);
nand U25767 (N_25767,N_24955,N_22261);
xnor U25768 (N_25768,N_22730,N_22430);
nor U25769 (N_25769,N_23696,N_22499);
nor U25770 (N_25770,N_20688,N_22406);
nor U25771 (N_25771,N_24182,N_24456);
nand U25772 (N_25772,N_20264,N_24727);
nor U25773 (N_25773,N_20395,N_21413);
or U25774 (N_25774,N_24931,N_22380);
and U25775 (N_25775,N_22172,N_24349);
and U25776 (N_25776,N_20777,N_23349);
or U25777 (N_25777,N_20364,N_23735);
and U25778 (N_25778,N_22939,N_20447);
nor U25779 (N_25779,N_23602,N_22320);
or U25780 (N_25780,N_24135,N_20607);
or U25781 (N_25781,N_20635,N_21128);
nor U25782 (N_25782,N_20448,N_23480);
xnor U25783 (N_25783,N_24862,N_20317);
or U25784 (N_25784,N_21009,N_22424);
xnor U25785 (N_25785,N_22619,N_22076);
nand U25786 (N_25786,N_21844,N_23529);
nor U25787 (N_25787,N_23272,N_22764);
or U25788 (N_25788,N_20762,N_24934);
nor U25789 (N_25789,N_24427,N_21993);
xor U25790 (N_25790,N_21780,N_20353);
or U25791 (N_25791,N_23893,N_24304);
or U25792 (N_25792,N_24186,N_20857);
nand U25793 (N_25793,N_23748,N_21648);
nand U25794 (N_25794,N_24044,N_22984);
nor U25795 (N_25795,N_23084,N_22823);
nand U25796 (N_25796,N_21590,N_24087);
nor U25797 (N_25797,N_20045,N_22633);
xnor U25798 (N_25798,N_21278,N_23100);
nor U25799 (N_25799,N_20319,N_23887);
xnor U25800 (N_25800,N_21942,N_21943);
xnor U25801 (N_25801,N_21436,N_20069);
xor U25802 (N_25802,N_23063,N_23578);
nor U25803 (N_25803,N_21344,N_24539);
xnor U25804 (N_25804,N_24774,N_24744);
nand U25805 (N_25805,N_22885,N_20820);
and U25806 (N_25806,N_22763,N_20993);
xnor U25807 (N_25807,N_24583,N_23317);
nand U25808 (N_25808,N_20516,N_24577);
nor U25809 (N_25809,N_20637,N_23135);
nand U25810 (N_25810,N_21379,N_24553);
nand U25811 (N_25811,N_22605,N_21370);
or U25812 (N_25812,N_22591,N_21520);
or U25813 (N_25813,N_23214,N_21544);
or U25814 (N_25814,N_22191,N_22634);
nand U25815 (N_25815,N_23121,N_21242);
or U25816 (N_25816,N_24745,N_23389);
nand U25817 (N_25817,N_23871,N_24612);
and U25818 (N_25818,N_20468,N_24430);
and U25819 (N_25819,N_20379,N_20702);
nand U25820 (N_25820,N_22514,N_20435);
nand U25821 (N_25821,N_20423,N_22589);
or U25822 (N_25822,N_24506,N_20517);
and U25823 (N_25823,N_21920,N_20522);
and U25824 (N_25824,N_21228,N_23795);
nor U25825 (N_25825,N_23145,N_21497);
and U25826 (N_25826,N_20831,N_20290);
and U25827 (N_25827,N_23966,N_24264);
nand U25828 (N_25828,N_20890,N_24204);
nor U25829 (N_25829,N_24894,N_22587);
nor U25830 (N_25830,N_22665,N_20816);
xor U25831 (N_25831,N_24024,N_23216);
and U25832 (N_25832,N_22925,N_22753);
or U25833 (N_25833,N_21074,N_22548);
nand U25834 (N_25834,N_22898,N_22062);
xnor U25835 (N_25835,N_22614,N_22195);
nor U25836 (N_25836,N_20110,N_23245);
nand U25837 (N_25837,N_20323,N_20755);
xnor U25838 (N_25838,N_22035,N_21627);
or U25839 (N_25839,N_22475,N_22791);
xor U25840 (N_25840,N_20220,N_23470);
xnor U25841 (N_25841,N_21486,N_22149);
and U25842 (N_25842,N_21059,N_23526);
nand U25843 (N_25843,N_24417,N_23881);
nand U25844 (N_25844,N_20203,N_23051);
or U25845 (N_25845,N_21812,N_24277);
and U25846 (N_25846,N_20008,N_22363);
nor U25847 (N_25847,N_20307,N_24690);
xnor U25848 (N_25848,N_21291,N_23608);
xnor U25849 (N_25849,N_21604,N_21039);
xnor U25850 (N_25850,N_24900,N_21512);
nor U25851 (N_25851,N_22075,N_24392);
nand U25852 (N_25852,N_24945,N_23540);
nand U25853 (N_25853,N_23859,N_22824);
xor U25854 (N_25854,N_23854,N_22802);
or U25855 (N_25855,N_23524,N_23160);
nor U25856 (N_25856,N_21295,N_21602);
and U25857 (N_25857,N_23431,N_23221);
nand U25858 (N_25858,N_21694,N_24735);
nor U25859 (N_25859,N_22292,N_21007);
and U25860 (N_25860,N_24581,N_20597);
and U25861 (N_25861,N_21914,N_23807);
and U25862 (N_25862,N_20550,N_22688);
xor U25863 (N_25863,N_24584,N_23280);
xor U25864 (N_25864,N_22482,N_23584);
nor U25865 (N_25865,N_20758,N_21672);
nor U25866 (N_25866,N_20686,N_22408);
xor U25867 (N_25867,N_22318,N_20907);
nand U25868 (N_25868,N_21095,N_22205);
nor U25869 (N_25869,N_21568,N_22337);
and U25870 (N_25870,N_22186,N_20743);
nor U25871 (N_25871,N_22115,N_22349);
or U25872 (N_25872,N_21595,N_21027);
xor U25873 (N_25873,N_20713,N_20419);
and U25874 (N_25874,N_21503,N_20086);
and U25875 (N_25875,N_24252,N_24441);
nor U25876 (N_25876,N_23977,N_23465);
or U25877 (N_25877,N_21153,N_21753);
nor U25878 (N_25878,N_22676,N_22831);
or U25879 (N_25879,N_21881,N_20107);
nand U25880 (N_25880,N_22126,N_22145);
or U25881 (N_25881,N_23712,N_22083);
or U25882 (N_25882,N_24334,N_24288);
or U25883 (N_25883,N_24994,N_22024);
xnor U25884 (N_25884,N_23326,N_23159);
nand U25885 (N_25885,N_22559,N_20218);
xnor U25886 (N_25886,N_20087,N_23246);
nand U25887 (N_25887,N_21666,N_21607);
or U25888 (N_25888,N_24342,N_24174);
nor U25889 (N_25889,N_24437,N_24731);
xnor U25890 (N_25890,N_24331,N_23779);
or U25891 (N_25891,N_24697,N_24737);
xor U25892 (N_25892,N_23747,N_21767);
or U25893 (N_25893,N_24282,N_21789);
nor U25894 (N_25894,N_24976,N_20790);
or U25895 (N_25895,N_22339,N_24524);
or U25896 (N_25896,N_22840,N_21720);
or U25897 (N_25897,N_20645,N_21424);
and U25898 (N_25898,N_24109,N_24626);
nand U25899 (N_25899,N_23090,N_21047);
xnor U25900 (N_25900,N_20496,N_22480);
nor U25901 (N_25901,N_22534,N_20320);
or U25902 (N_25902,N_20033,N_22489);
xor U25903 (N_25903,N_21555,N_20427);
nand U25904 (N_25904,N_24244,N_21704);
xnor U25905 (N_25905,N_20620,N_24114);
or U25906 (N_25906,N_23416,N_22914);
or U25907 (N_25907,N_20406,N_23462);
nand U25908 (N_25908,N_20963,N_23458);
xor U25909 (N_25909,N_23637,N_20396);
xor U25910 (N_25910,N_23181,N_21864);
nand U25911 (N_25911,N_21149,N_21371);
and U25912 (N_25912,N_22414,N_24543);
nor U25913 (N_25913,N_23756,N_22378);
or U25914 (N_25914,N_21094,N_23982);
xor U25915 (N_25915,N_24979,N_23886);
and U25916 (N_25916,N_21485,N_23504);
and U25917 (N_25917,N_23765,N_21538);
nand U25918 (N_25918,N_24434,N_23305);
and U25919 (N_25919,N_24029,N_21673);
or U25920 (N_25920,N_22013,N_20236);
nand U25921 (N_25921,N_21636,N_20158);
and U25922 (N_25922,N_21856,N_23889);
xor U25923 (N_25923,N_22352,N_20169);
or U25924 (N_25924,N_24589,N_24173);
xor U25925 (N_25925,N_20894,N_23672);
xnor U25926 (N_25926,N_24682,N_22884);
or U25927 (N_25927,N_20287,N_21390);
nand U25928 (N_25928,N_20474,N_23362);
nand U25929 (N_25929,N_23714,N_22880);
nand U25930 (N_25930,N_22905,N_24641);
xor U25931 (N_25931,N_24336,N_22130);
or U25932 (N_25932,N_22058,N_24793);
or U25933 (N_25933,N_21700,N_20255);
nand U25934 (N_25934,N_21945,N_20401);
nand U25935 (N_25935,N_21701,N_22953);
or U25936 (N_25936,N_20888,N_22709);
nand U25937 (N_25937,N_23833,N_23034);
or U25938 (N_25938,N_22627,N_24345);
xnor U25939 (N_25939,N_22910,N_20917);
and U25940 (N_25940,N_21452,N_21953);
or U25941 (N_25941,N_22206,N_23299);
xnor U25942 (N_25942,N_20720,N_24508);
xnor U25943 (N_25943,N_23353,N_20889);
nand U25944 (N_25944,N_20208,N_21498);
xor U25945 (N_25945,N_21603,N_20175);
and U25946 (N_25946,N_22175,N_24041);
and U25947 (N_25947,N_20856,N_20918);
or U25948 (N_25948,N_24397,N_23435);
or U25949 (N_25949,N_20020,N_22388);
xnor U25950 (N_25950,N_24777,N_20215);
or U25951 (N_25951,N_22048,N_24414);
xnor U25952 (N_25952,N_20973,N_23771);
or U25953 (N_25953,N_22784,N_20976);
nor U25954 (N_25954,N_23767,N_23905);
nand U25955 (N_25955,N_22562,N_21282);
xnor U25956 (N_25956,N_22886,N_20193);
and U25957 (N_25957,N_23476,N_23149);
or U25958 (N_25958,N_24154,N_22968);
xnor U25959 (N_25959,N_22628,N_22300);
xor U25960 (N_25960,N_24840,N_24804);
xnor U25961 (N_25961,N_20878,N_24333);
xor U25962 (N_25962,N_20596,N_21965);
nor U25963 (N_25963,N_22244,N_21761);
or U25964 (N_25964,N_21494,N_20194);
or U25965 (N_25965,N_24787,N_24699);
or U25966 (N_25966,N_24362,N_23190);
nor U25967 (N_25967,N_22582,N_23318);
nand U25968 (N_25968,N_20339,N_23092);
nand U25969 (N_25969,N_23402,N_20560);
or U25970 (N_25970,N_22805,N_23290);
nor U25971 (N_25971,N_20460,N_23693);
nand U25972 (N_25972,N_22640,N_24254);
nor U25973 (N_25973,N_21147,N_20376);
or U25974 (N_25974,N_21210,N_20534);
nand U25975 (N_25975,N_21533,N_20272);
or U25976 (N_25976,N_21941,N_20157);
nand U25977 (N_25977,N_21211,N_22242);
or U25978 (N_25978,N_20231,N_23950);
and U25979 (N_25979,N_22190,N_23593);
xor U25980 (N_25980,N_22930,N_21724);
xnor U25981 (N_25981,N_24717,N_24676);
nand U25982 (N_25982,N_22626,N_21430);
and U25983 (N_25983,N_24193,N_21522);
nand U25984 (N_25984,N_24555,N_21729);
nor U25985 (N_25985,N_24980,N_24824);
or U25986 (N_25986,N_21934,N_21862);
or U25987 (N_25987,N_20865,N_24449);
or U25988 (N_25988,N_24214,N_21689);
nor U25989 (N_25989,N_21067,N_20794);
and U25990 (N_25990,N_23193,N_20196);
or U25991 (N_25991,N_24513,N_20989);
or U25992 (N_25992,N_22315,N_20931);
nand U25993 (N_25993,N_23806,N_24128);
or U25994 (N_25994,N_22528,N_24518);
xnor U25995 (N_25995,N_20847,N_21827);
nand U25996 (N_25996,N_23579,N_20561);
xor U25997 (N_25997,N_22521,N_20754);
xnor U25998 (N_25998,N_24779,N_21543);
and U25999 (N_25999,N_22445,N_24092);
xor U26000 (N_26000,N_23559,N_21591);
or U26001 (N_26001,N_21902,N_24920);
and U26002 (N_26002,N_22392,N_24379);
and U26003 (N_26003,N_23558,N_24591);
or U26004 (N_26004,N_22159,N_24668);
nand U26005 (N_26005,N_23028,N_23952);
and U26006 (N_26006,N_23139,N_24773);
and U26007 (N_26007,N_21324,N_22741);
nor U26008 (N_26008,N_20896,N_24216);
xor U26009 (N_26009,N_22859,N_21695);
or U26010 (N_26010,N_22144,N_21579);
nand U26011 (N_26011,N_22544,N_23170);
nor U26012 (N_26012,N_22493,N_20965);
nand U26013 (N_26013,N_20830,N_22361);
xor U26014 (N_26014,N_23203,N_22022);
or U26015 (N_26015,N_24880,N_20129);
nor U26016 (N_26016,N_23329,N_23039);
or U26017 (N_26017,N_23361,N_21176);
or U26018 (N_26018,N_23085,N_20826);
and U26019 (N_26019,N_20932,N_22987);
xnor U26020 (N_26020,N_22164,N_20082);
nand U26021 (N_26021,N_20293,N_24816);
nand U26022 (N_26022,N_21592,N_21549);
and U26023 (N_26023,N_20570,N_21766);
nand U26024 (N_26024,N_23426,N_22719);
and U26025 (N_26025,N_24872,N_20127);
or U26026 (N_26026,N_23448,N_20278);
nand U26027 (N_26027,N_24005,N_23192);
and U26028 (N_26028,N_23363,N_22485);
or U26029 (N_26029,N_24556,N_23857);
nor U26030 (N_26030,N_21992,N_24909);
nor U26031 (N_26031,N_23959,N_21016);
nor U26032 (N_26032,N_23058,N_22602);
nor U26033 (N_26033,N_21475,N_23043);
or U26034 (N_26034,N_23042,N_21148);
nand U26035 (N_26035,N_22072,N_21461);
xnor U26036 (N_26036,N_21845,N_21341);
nand U26037 (N_26037,N_23674,N_22765);
and U26038 (N_26038,N_22379,N_21867);
nand U26039 (N_26039,N_21279,N_21070);
xor U26040 (N_26040,N_24377,N_21213);
and U26041 (N_26041,N_22529,N_22431);
or U26042 (N_26042,N_24014,N_23056);
xor U26043 (N_26043,N_24885,N_24817);
or U26044 (N_26044,N_21737,N_23943);
nand U26045 (N_26045,N_20041,N_20113);
and U26046 (N_26046,N_22409,N_21467);
nand U26047 (N_26047,N_21403,N_21754);
nand U26048 (N_26048,N_23577,N_20815);
or U26049 (N_26049,N_24007,N_23222);
or U26050 (N_26050,N_21907,N_20538);
nor U26051 (N_26051,N_22933,N_24073);
and U26052 (N_26052,N_20780,N_21775);
xnor U26053 (N_26053,N_23377,N_24541);
nand U26054 (N_26054,N_22712,N_23918);
and U26055 (N_26055,N_23535,N_23176);
or U26056 (N_26056,N_20397,N_23240);
nand U26057 (N_26057,N_24743,N_22762);
nor U26058 (N_26058,N_24530,N_20671);
xor U26059 (N_26059,N_22497,N_24236);
and U26060 (N_26060,N_23990,N_24529);
or U26061 (N_26061,N_22790,N_23653);
or U26062 (N_26062,N_24975,N_21471);
and U26063 (N_26063,N_24447,N_23331);
or U26064 (N_26064,N_22635,N_21312);
xor U26065 (N_26065,N_24471,N_20950);
nand U26066 (N_26066,N_20391,N_22865);
nand U26067 (N_26067,N_24645,N_23624);
nor U26068 (N_26068,N_22011,N_22053);
or U26069 (N_26069,N_22517,N_24458);
or U26070 (N_26070,N_23082,N_20608);
or U26071 (N_26071,N_22684,N_23384);
xnor U26072 (N_26072,N_20050,N_20098);
and U26073 (N_26073,N_21798,N_22950);
xnor U26074 (N_26074,N_22596,N_24219);
xnor U26075 (N_26075,N_23574,N_22568);
xnor U26076 (N_26076,N_23127,N_23040);
or U26077 (N_26077,N_20066,N_20152);
or U26078 (N_26078,N_23638,N_24884);
nor U26079 (N_26079,N_20490,N_20710);
nor U26080 (N_26080,N_24004,N_23923);
nand U26081 (N_26081,N_20726,N_20488);
nor U26082 (N_26082,N_20130,N_22645);
xnor U26083 (N_26083,N_22536,N_22997);
xnor U26084 (N_26084,N_21935,N_22045);
and U26085 (N_26085,N_24962,N_21201);
nand U26086 (N_26086,N_24950,N_23027);
nor U26087 (N_26087,N_21909,N_23960);
xor U26088 (N_26088,N_24118,N_24383);
nand U26089 (N_26089,N_24298,N_23778);
xnor U26090 (N_26090,N_24526,N_20639);
or U26091 (N_26091,N_22542,N_22936);
nor U26092 (N_26092,N_22537,N_23999);
and U26093 (N_26093,N_21622,N_23678);
or U26094 (N_26094,N_24608,N_23148);
and U26095 (N_26095,N_23374,N_24919);
nand U26096 (N_26096,N_23561,N_22032);
xor U26097 (N_26097,N_20428,N_20235);
and U26098 (N_26098,N_24124,N_24142);
nand U26099 (N_26099,N_20268,N_21573);
and U26100 (N_26100,N_20882,N_20883);
or U26101 (N_26101,N_23123,N_23307);
nand U26102 (N_26102,N_21287,N_21903);
or U26103 (N_26103,N_22207,N_20788);
or U26104 (N_26104,N_23472,N_22983);
or U26105 (N_26105,N_22054,N_24265);
nor U26106 (N_26106,N_22123,N_24250);
or U26107 (N_26107,N_24967,N_20559);
or U26108 (N_26108,N_24795,N_23478);
or U26109 (N_26109,N_22915,N_21677);
xor U26110 (N_26110,N_21132,N_20795);
and U26111 (N_26111,N_23877,N_23891);
and U26112 (N_26112,N_20064,N_24227);
or U26113 (N_26113,N_24763,N_21840);
nand U26114 (N_26114,N_24185,N_24618);
nand U26115 (N_26115,N_22494,N_23705);
xor U26116 (N_26116,N_22538,N_22679);
nor U26117 (N_26117,N_21703,N_24175);
or U26118 (N_26118,N_24472,N_21671);
nand U26119 (N_26119,N_21152,N_23523);
and U26120 (N_26120,N_21897,N_20705);
nor U26121 (N_26121,N_22637,N_21185);
xor U26122 (N_26122,N_20210,N_21900);
xnor U26123 (N_26123,N_24103,N_24218);
xor U26124 (N_26124,N_24798,N_21099);
xor U26125 (N_26125,N_22049,N_24136);
and U26126 (N_26126,N_23141,N_21567);
and U26127 (N_26127,N_24442,N_24825);
and U26128 (N_26128,N_22729,N_21321);
xor U26129 (N_26129,N_23495,N_21597);
xor U26130 (N_26130,N_22389,N_22787);
and U26131 (N_26131,N_21574,N_23147);
or U26132 (N_26132,N_22931,N_20230);
nand U26133 (N_26133,N_22999,N_21841);
and U26134 (N_26134,N_23073,N_24091);
or U26135 (N_26135,N_22705,N_22717);
and U26136 (N_26136,N_24813,N_21373);
and U26137 (N_26137,N_21423,N_21065);
nor U26138 (N_26138,N_20262,N_23662);
nor U26139 (N_26139,N_24881,N_23835);
nand U26140 (N_26140,N_20136,N_24429);
and U26141 (N_26141,N_22476,N_20933);
nand U26142 (N_26142,N_23763,N_21204);
xor U26143 (N_26143,N_20845,N_23516);
nand U26144 (N_26144,N_22918,N_20706);
and U26145 (N_26145,N_21253,N_20494);
or U26146 (N_26146,N_20199,N_21769);
nor U26147 (N_26147,N_22525,N_22451);
or U26148 (N_26148,N_23816,N_24607);
nor U26149 (N_26149,N_22454,N_22755);
nand U26150 (N_26150,N_24197,N_22680);
nor U26151 (N_26151,N_21265,N_20551);
xor U26152 (N_26152,N_20582,N_22297);
or U26153 (N_26153,N_21223,N_20185);
and U26154 (N_26154,N_22855,N_20913);
nor U26155 (N_26155,N_23038,N_24621);
xor U26156 (N_26156,N_24454,N_24974);
nand U26157 (N_26157,N_22607,N_24457);
nor U26158 (N_26158,N_20588,N_21209);
xor U26159 (N_26159,N_20543,N_22311);
nor U26160 (N_26160,N_22652,N_21406);
nand U26161 (N_26161,N_21639,N_20828);
or U26162 (N_26162,N_23919,N_22621);
nor U26163 (N_26163,N_21839,N_23241);
nor U26164 (N_26164,N_24355,N_24720);
and U26165 (N_26165,N_22253,N_22237);
nand U26166 (N_26166,N_21028,N_23296);
or U26167 (N_26167,N_21357,N_23519);
and U26168 (N_26168,N_24179,N_20606);
nand U26169 (N_26169,N_23212,N_20390);
or U26170 (N_26170,N_23623,N_23695);
nand U26171 (N_26171,N_20502,N_21796);
nand U26172 (N_26172,N_23489,N_21519);
nor U26173 (N_26173,N_22443,N_20028);
nand U26174 (N_26174,N_24698,N_21612);
nand U26175 (N_26175,N_21270,N_23357);
or U26176 (N_26176,N_21217,N_22353);
nand U26177 (N_26177,N_21855,N_22592);
or U26178 (N_26178,N_24432,N_21252);
xor U26179 (N_26179,N_24426,N_22071);
xnor U26180 (N_26180,N_20249,N_23132);
xnor U26181 (N_26181,N_21959,N_20392);
or U26182 (N_26182,N_21891,N_21092);
or U26183 (N_26183,N_20232,N_23520);
and U26184 (N_26184,N_22966,N_24451);
and U26185 (N_26185,N_24462,N_21644);
xnor U26186 (N_26186,N_20864,N_23760);
or U26187 (N_26187,N_20105,N_21873);
nand U26188 (N_26188,N_23605,N_24515);
xnor U26189 (N_26189,N_22550,N_20284);
or U26190 (N_26190,N_24784,N_21958);
and U26191 (N_26191,N_23649,N_23061);
nor U26192 (N_26192,N_23484,N_24374);
and U26193 (N_26193,N_20084,N_22541);
or U26194 (N_26194,N_24043,N_23971);
and U26195 (N_26195,N_23689,N_24633);
and U26196 (N_26196,N_24385,N_24049);
nor U26197 (N_26197,N_23492,N_21385);
and U26198 (N_26198,N_21575,N_20501);
nor U26199 (N_26199,N_20048,N_20352);
or U26200 (N_26200,N_24393,N_22201);
nor U26201 (N_26201,N_21504,N_23780);
nand U26202 (N_26202,N_20111,N_23477);
nand U26203 (N_26203,N_21259,N_21735);
or U26204 (N_26204,N_20441,N_23713);
xnor U26205 (N_26205,N_20426,N_20646);
or U26206 (N_26206,N_22030,N_22651);
nand U26207 (N_26207,N_23964,N_21771);
xor U26208 (N_26208,N_24101,N_20080);
nand U26209 (N_26209,N_23001,N_20243);
nand U26210 (N_26210,N_20787,N_23200);
or U26211 (N_26211,N_21561,N_24710);
or U26212 (N_26212,N_20205,N_21029);
nand U26213 (N_26213,N_20626,N_20553);
and U26214 (N_26214,N_23078,N_24069);
and U26215 (N_26215,N_20730,N_20444);
nor U26216 (N_26216,N_20149,N_22835);
xnor U26217 (N_26217,N_20118,N_24258);
or U26218 (N_26218,N_23842,N_22750);
or U26219 (N_26219,N_22162,N_22693);
nand U26220 (N_26220,N_20812,N_23271);
nand U26221 (N_26221,N_23663,N_24402);
nand U26222 (N_26222,N_23820,N_22346);
and U26223 (N_26223,N_24494,N_20480);
and U26224 (N_26224,N_23114,N_24187);
or U26225 (N_26225,N_22862,N_20393);
xor U26226 (N_26226,N_23863,N_21195);
or U26227 (N_26227,N_23888,N_20012);
xnor U26228 (N_26228,N_20581,N_21093);
or U26229 (N_26229,N_22377,N_22449);
nor U26230 (N_26230,N_24112,N_22861);
nand U26231 (N_26231,N_21143,N_24963);
xor U26232 (N_26232,N_23210,N_21102);
nand U26233 (N_26233,N_24604,N_20300);
nand U26234 (N_26234,N_24680,N_21540);
nor U26235 (N_26235,N_21948,N_22432);
or U26236 (N_26236,N_24147,N_22834);
nand U26237 (N_26237,N_21138,N_24640);
or U26238 (N_26238,N_23467,N_22284);
nor U26239 (N_26239,N_20765,N_21619);
and U26240 (N_26240,N_23247,N_24761);
nor U26241 (N_26241,N_20141,N_20725);
and U26242 (N_26242,N_22873,N_23237);
or U26243 (N_26243,N_21630,N_20068);
nor U26244 (N_26244,N_24428,N_21013);
nand U26245 (N_26245,N_23297,N_20886);
xor U26246 (N_26246,N_23303,N_21613);
and U26247 (N_26247,N_20922,N_24480);
and U26248 (N_26248,N_22182,N_22531);
nand U26249 (N_26249,N_22166,N_21172);
nand U26250 (N_26250,N_21342,N_20032);
nor U26251 (N_26251,N_24190,N_22296);
xor U26252 (N_26252,N_23036,N_22897);
or U26253 (N_26253,N_20542,N_20015);
nor U26254 (N_26254,N_23479,N_24180);
nand U26255 (N_26255,N_21114,N_21740);
and U26256 (N_26256,N_21307,N_24993);
xor U26257 (N_26257,N_24443,N_24366);
nand U26258 (N_26258,N_22735,N_21617);
and U26259 (N_26259,N_21455,N_24201);
nor U26260 (N_26260,N_20122,N_21888);
and U26261 (N_26261,N_20408,N_24199);
xor U26262 (N_26262,N_23902,N_22733);
nor U26263 (N_26263,N_21928,N_23291);
nor U26264 (N_26264,N_22821,N_22822);
nand U26265 (N_26265,N_22841,N_24941);
nor U26266 (N_26266,N_24192,N_23372);
and U26267 (N_26267,N_22481,N_21653);
nand U26268 (N_26268,N_23880,N_22683);
nand U26269 (N_26269,N_21726,N_23118);
xnor U26270 (N_26270,N_24416,N_22372);
nand U26271 (N_26271,N_24233,N_23829);
and U26272 (N_26272,N_24896,N_22364);
and U26273 (N_26273,N_24702,N_22027);
nand U26274 (N_26274,N_23493,N_23998);
nor U26275 (N_26275,N_24940,N_24830);
and U26276 (N_26276,N_23953,N_21495);
or U26277 (N_26277,N_22487,N_22082);
xor U26278 (N_26278,N_24617,N_20277);
nand U26279 (N_26279,N_24125,N_23716);
nand U26280 (N_26280,N_21303,N_21001);
and U26281 (N_26281,N_20240,N_23824);
nand U26282 (N_26282,N_20736,N_22546);
and U26283 (N_26283,N_22980,N_24822);
xnor U26284 (N_26284,N_22798,N_24865);
nor U26285 (N_26285,N_22771,N_23885);
nand U26286 (N_26286,N_22757,N_21359);
nand U26287 (N_26287,N_22691,N_20531);
or U26288 (N_26288,N_20131,N_20338);
xnor U26289 (N_26289,N_22436,N_24875);
or U26290 (N_26290,N_22610,N_21256);
xor U26291 (N_26291,N_21382,N_22502);
or U26292 (N_26292,N_22350,N_24294);
and U26293 (N_26293,N_23898,N_22580);
nor U26294 (N_26294,N_21889,N_22367);
nand U26295 (N_26295,N_20495,N_21435);
xor U26296 (N_26296,N_22203,N_21752);
nand U26297 (N_26297,N_21306,N_22461);
nor U26298 (N_26298,N_21443,N_21082);
and U26299 (N_26299,N_24012,N_21493);
xnor U26300 (N_26300,N_20971,N_21861);
xnor U26301 (N_26301,N_20690,N_20487);
and U26302 (N_26302,N_20536,N_23509);
nor U26303 (N_26303,N_21705,N_24464);
nand U26304 (N_26304,N_22387,N_20309);
nor U26305 (N_26305,N_22342,N_24220);
and U26306 (N_26306,N_23708,N_22383);
or U26307 (N_26307,N_20280,N_23020);
or U26308 (N_26308,N_20912,N_21809);
nor U26309 (N_26309,N_20238,N_20680);
and U26310 (N_26310,N_23207,N_23157);
and U26311 (N_26311,N_22307,N_23884);
xor U26312 (N_26312,N_24164,N_22151);
nor U26313 (N_26313,N_20841,N_21685);
nor U26314 (N_26314,N_23546,N_21587);
nor U26315 (N_26315,N_21050,N_22812);
nor U26316 (N_26316,N_23862,N_24687);
and U26317 (N_26317,N_20473,N_21807);
nand U26318 (N_26318,N_23064,N_20256);
or U26319 (N_26319,N_21014,N_20489);
nand U26320 (N_26320,N_21337,N_24683);
nand U26321 (N_26321,N_24890,N_21898);
and U26322 (N_26322,N_21545,N_23436);
nand U26323 (N_26323,N_23595,N_20198);
xnor U26324 (N_26324,N_24713,N_21444);
xnor U26325 (N_26325,N_21784,N_22137);
nand U26326 (N_26326,N_24856,N_24978);
and U26327 (N_26327,N_22507,N_23487);
or U26328 (N_26328,N_22557,N_20972);
nor U26329 (N_26329,N_21790,N_20389);
nor U26330 (N_26330,N_23164,N_24303);
xor U26331 (N_26331,N_23916,N_22155);
nor U26332 (N_26332,N_20410,N_23163);
xnor U26333 (N_26333,N_23130,N_20368);
nor U26334 (N_26334,N_21600,N_20164);
nor U26335 (N_26335,N_23976,N_20962);
or U26336 (N_26336,N_22238,N_22923);
xor U26337 (N_26337,N_23178,N_21951);
nor U26338 (N_26338,N_22473,N_20492);
or U26339 (N_26339,N_24595,N_20014);
nand U26340 (N_26340,N_23832,N_22400);
nor U26341 (N_26341,N_24921,N_22830);
or U26342 (N_26342,N_21489,N_23665);
xnor U26343 (N_26343,N_21774,N_24895);
xor U26344 (N_26344,N_22584,N_21151);
nor U26345 (N_26345,N_20486,N_24730);
nor U26346 (N_26346,N_20979,N_22826);
xnor U26347 (N_26347,N_22179,N_21165);
xor U26348 (N_26348,N_23185,N_23126);
and U26349 (N_26349,N_20463,N_21389);
nor U26350 (N_26350,N_24448,N_21874);
and U26351 (N_26351,N_20628,N_22171);
nand U26352 (N_26352,N_24308,N_24675);
nor U26353 (N_26353,N_20717,N_22883);
xnor U26354 (N_26354,N_23915,N_23655);
nand U26355 (N_26355,N_23080,N_23619);
xnor U26356 (N_26356,N_20749,N_24083);
xnor U26357 (N_26357,N_24097,N_23414);
or U26358 (N_26358,N_22005,N_24381);
nor U26359 (N_26359,N_22245,N_23409);
or U26360 (N_26360,N_23354,N_24914);
or U26361 (N_26361,N_21160,N_24191);
or U26362 (N_26362,N_22397,N_20259);
or U26363 (N_26363,N_20177,N_24104);
nand U26364 (N_26364,N_21388,N_21872);
and U26365 (N_26365,N_23345,N_22271);
or U26366 (N_26366,N_23718,N_23022);
and U26367 (N_26367,N_24081,N_21852);
xor U26368 (N_26368,N_21002,N_23199);
nor U26369 (N_26369,N_24854,N_20768);
and U26370 (N_26370,N_23031,N_20946);
xnor U26371 (N_26371,N_24587,N_21803);
or U26372 (N_26372,N_21665,N_21488);
and U26373 (N_26373,N_21477,N_22615);
nand U26374 (N_26374,N_24977,N_23171);
or U26375 (N_26375,N_22468,N_23161);
and U26376 (N_26376,N_20554,N_23687);
xnor U26377 (N_26377,N_24821,N_23334);
nor U26378 (N_26378,N_20442,N_24211);
xnor U26379 (N_26379,N_23262,N_22530);
xor U26380 (N_26380,N_24557,N_24867);
nor U26381 (N_26381,N_22268,N_20968);
nand U26382 (N_26382,N_23969,N_20804);
xnor U26383 (N_26383,N_23232,N_21973);
nor U26384 (N_26384,N_21853,N_22846);
or U26385 (N_26385,N_20727,N_21578);
xnor U26386 (N_26386,N_21190,N_23350);
nand U26387 (N_26387,N_20652,N_21267);
nand U26388 (N_26388,N_24008,N_24566);
nand U26389 (N_26389,N_22034,N_22421);
or U26390 (N_26390,N_24801,N_22230);
or U26391 (N_26391,N_23313,N_23037);
xnor U26392 (N_26392,N_21456,N_23644);
and U26393 (N_26393,N_24059,N_21096);
or U26394 (N_26394,N_22087,N_22932);
or U26395 (N_26395,N_23927,N_23812);
or U26396 (N_26396,N_23979,N_20221);
or U26397 (N_26397,N_23866,N_22410);
and U26398 (N_26398,N_24478,N_24631);
nand U26399 (N_26399,N_22492,N_23459);
nor U26400 (N_26400,N_21539,N_22817);
or U26401 (N_26401,N_23219,N_23873);
xor U26402 (N_26402,N_23008,N_20874);
xnor U26403 (N_26403,N_22212,N_20753);
and U26404 (N_26404,N_23295,N_22697);
or U26405 (N_26405,N_21676,N_24137);
nand U26406 (N_26406,N_23430,N_21734);
or U26407 (N_26407,N_21972,N_22064);
nand U26408 (N_26408,N_22138,N_20575);
nand U26409 (N_26409,N_23463,N_20227);
or U26410 (N_26410,N_22696,N_22952);
and U26411 (N_26411,N_20095,N_24917);
or U26412 (N_26412,N_23000,N_21999);
nand U26413 (N_26413,N_24882,N_23087);
nand U26414 (N_26414,N_20998,N_24353);
or U26415 (N_26415,N_22204,N_22343);
nor U26416 (N_26416,N_21950,N_23865);
nor U26417 (N_26417,N_21621,N_20745);
nand U26418 (N_26418,N_20806,N_24263);
nor U26419 (N_26419,N_22994,N_24876);
nand U26420 (N_26420,N_23722,N_22864);
nor U26421 (N_26421,N_21657,N_24602);
nand U26422 (N_26422,N_20034,N_22488);
xnor U26423 (N_26423,N_23450,N_20044);
nand U26424 (N_26424,N_22533,N_23794);
and U26425 (N_26425,N_24637,N_22957);
nand U26426 (N_26426,N_22037,N_23802);
or U26427 (N_26427,N_22382,N_23136);
or U26428 (N_26428,N_24712,N_23277);
xnor U26429 (N_26429,N_20002,N_23894);
nor U26430 (N_26430,N_20782,N_22853);
xor U26431 (N_26431,N_23762,N_20214);
and U26432 (N_26432,N_23452,N_22912);
nor U26433 (N_26433,N_20760,N_23285);
and U26434 (N_26434,N_22827,N_22425);
and U26435 (N_26435,N_21261,N_22662);
nor U26436 (N_26436,N_20481,N_21614);
xnor U26437 (N_26437,N_20248,N_23764);
nor U26438 (N_26438,N_21906,N_24404);
xnor U26439 (N_26439,N_21298,N_24184);
nand U26440 (N_26440,N_21581,N_20146);
xor U26441 (N_26441,N_21349,N_23706);
nand U26442 (N_26442,N_20773,N_20891);
xnor U26443 (N_26443,N_20723,N_21200);
nand U26444 (N_26444,N_23451,N_21222);
xnor U26445 (N_26445,N_21006,N_21340);
nand U26446 (N_26446,N_21005,N_20241);
xor U26447 (N_26447,N_24422,N_20715);
or U26448 (N_26448,N_22246,N_23552);
xnor U26449 (N_26449,N_21248,N_24023);
or U26450 (N_26450,N_21976,N_24296);
and U26451 (N_26451,N_24110,N_24606);
and U26452 (N_26452,N_20691,N_20821);
nor U26453 (N_26453,N_21870,N_22570);
nand U26454 (N_26454,N_21460,N_20271);
nand U26455 (N_26455,N_24151,N_22052);
and U26456 (N_26456,N_24688,N_20381);
xor U26457 (N_26457,N_20384,N_22904);
or U26458 (N_26458,N_20916,N_21682);
nor U26459 (N_26459,N_22329,N_21658);
nand U26460 (N_26460,N_24297,N_23837);
nor U26461 (N_26461,N_21462,N_24998);
nand U26462 (N_26462,N_24223,N_20402);
nand U26463 (N_26463,N_21962,N_23993);
or U26464 (N_26464,N_20733,N_20742);
nand U26465 (N_26465,N_20301,N_20206);
nor U26466 (N_26466,N_21721,N_21301);
nand U26467 (N_26467,N_22023,N_22294);
nor U26468 (N_26468,N_23549,N_22447);
nand U26469 (N_26469,N_24938,N_22336);
and U26470 (N_26470,N_21967,N_24324);
or U26471 (N_26471,N_23062,N_20719);
nor U26472 (N_26472,N_22993,N_24347);
xnor U26473 (N_26473,N_21496,N_22574);
or U26474 (N_26474,N_22815,N_20155);
nand U26475 (N_26475,N_21333,N_22415);
xnor U26476 (N_26476,N_20434,N_24705);
xnor U26477 (N_26477,N_24492,N_23548);
nor U26478 (N_26478,N_23814,N_23442);
nand U26479 (N_26479,N_20144,N_22900);
xor U26480 (N_26480,N_24033,N_22638);
nand U26481 (N_26481,N_24585,N_24547);
nand U26482 (N_26482,N_21407,N_20614);
or U26483 (N_26483,N_22351,N_24306);
and U26484 (N_26484,N_21345,N_22319);
nor U26485 (N_26485,N_20618,N_23379);
nor U26486 (N_26486,N_24913,N_24916);
and U26487 (N_26487,N_21550,N_20833);
nor U26488 (N_26488,N_23947,N_22523);
nor U26489 (N_26489,N_21730,N_24261);
or U26490 (N_26490,N_21365,N_21472);
or U26491 (N_26491,N_21120,N_21281);
and U26492 (N_26492,N_20949,N_20370);
nor U26493 (N_26493,N_23774,N_24459);
or U26494 (N_26494,N_24015,N_24072);
nand U26495 (N_26495,N_21280,N_24067);
and U26496 (N_26496,N_21167,N_22142);
xnor U26497 (N_26497,N_20928,N_20029);
or U26498 (N_26498,N_20004,N_21541);
and U26499 (N_26499,N_20007,N_21702);
xor U26500 (N_26500,N_24453,N_24337);
xnor U26501 (N_26501,N_23813,N_23925);
nor U26502 (N_26502,N_23293,N_21750);
and U26503 (N_26503,N_24736,N_21890);
or U26504 (N_26504,N_22498,N_24903);
and U26505 (N_26505,N_23684,N_21319);
nand U26506 (N_26506,N_20555,N_24729);
and U26507 (N_26507,N_21690,N_22202);
nand U26508 (N_26508,N_21929,N_21536);
and U26509 (N_26509,N_21745,N_23182);
and U26510 (N_26510,N_20400,N_22314);
nand U26511 (N_26511,N_20023,N_21787);
xor U26512 (N_26512,N_24491,N_20818);
nand U26513 (N_26513,N_21117,N_23502);
nand U26514 (N_26514,N_23408,N_23067);
nand U26515 (N_26515,N_24806,N_20251);
or U26516 (N_26516,N_22442,N_22274);
xor U26517 (N_26517,N_23720,N_21202);
nor U26518 (N_26518,N_22393,N_20343);
and U26519 (N_26519,N_20257,N_21688);
xor U26520 (N_26520,N_20957,N_22084);
nor U26521 (N_26521,N_21431,N_24599);
or U26522 (N_26522,N_23937,N_24217);
and U26523 (N_26523,N_23425,N_21234);
nand U26524 (N_26524,N_21121,N_20074);
nor U26525 (N_26525,N_21358,N_24259);
nor U26526 (N_26526,N_20781,N_22080);
nor U26527 (N_26527,N_23542,N_23503);
xnor U26528 (N_26528,N_20246,N_20684);
and U26529 (N_26529,N_23830,N_20102);
or U26530 (N_26530,N_24546,N_20528);
nand U26531 (N_26531,N_21328,N_20552);
xnor U26532 (N_26532,N_22682,N_22215);
or U26533 (N_26533,N_21136,N_23908);
or U26534 (N_26534,N_21046,N_20746);
nand U26535 (N_26535,N_24852,N_21449);
xor U26536 (N_26536,N_21484,N_20627);
and U26537 (N_26537,N_24380,N_20088);
and U26538 (N_26538,N_20842,N_22803);
or U26539 (N_26539,N_20643,N_24079);
xnor U26540 (N_26540,N_20980,N_21421);
xnor U26541 (N_26541,N_24150,N_24042);
xor U26542 (N_26542,N_20663,N_24685);
and U26543 (N_26543,N_23963,N_23496);
nand U26544 (N_26544,N_21659,N_24609);
and U26545 (N_26545,N_22793,N_24695);
and U26546 (N_26546,N_20285,N_24273);
nor U26547 (N_26547,N_21087,N_24650);
nand U26548 (N_26548,N_22328,N_22213);
xnor U26549 (N_26549,N_21645,N_24897);
nand U26550 (N_26550,N_21145,N_20483);
xnor U26551 (N_26551,N_24159,N_20288);
and U26552 (N_26552,N_23041,N_24420);
or U26553 (N_26553,N_21969,N_20549);
nand U26554 (N_26554,N_23852,N_24461);
or U26555 (N_26555,N_24692,N_23086);
xor U26556 (N_26556,N_21231,N_21880);
nor U26557 (N_26557,N_24907,N_22055);
or U26558 (N_26558,N_22219,N_20412);
nor U26559 (N_26559,N_24283,N_20785);
or U26560 (N_26560,N_23075,N_23848);
or U26561 (N_26561,N_22229,N_24706);
nand U26562 (N_26562,N_22429,N_20279);
xnor U26563 (N_26563,N_24586,N_21930);
nand U26564 (N_26564,N_22209,N_22290);
nor U26565 (N_26565,N_22143,N_23137);
xor U26566 (N_26566,N_20844,N_21719);
and U26567 (N_26567,N_23576,N_24868);
xor U26568 (N_26568,N_21860,N_23858);
nor U26569 (N_26569,N_21966,N_22929);
nand U26570 (N_26570,N_21525,N_20508);
xnor U26571 (N_26571,N_24415,N_22161);
xor U26572 (N_26572,N_22483,N_21731);
nand U26573 (N_26573,N_24636,N_20852);
nand U26574 (N_26574,N_22849,N_24814);
nand U26575 (N_26575,N_22452,N_22068);
and U26576 (N_26576,N_21583,N_20591);
nor U26577 (N_26577,N_22644,N_20759);
xor U26578 (N_26578,N_20523,N_24395);
nand U26579 (N_26579,N_20589,N_20761);
nor U26580 (N_26580,N_21439,N_24832);
and U26581 (N_26581,N_23046,N_21949);
nor U26582 (N_26582,N_20055,N_22600);
xor U26583 (N_26583,N_21192,N_21896);
and U26584 (N_26584,N_23634,N_20116);
xnor U26585 (N_26585,N_22641,N_22876);
or U26586 (N_26586,N_22833,N_23669);
xor U26587 (N_26587,N_23359,N_22427);
and U26588 (N_26588,N_24721,N_21534);
nand U26589 (N_26589,N_20944,N_20724);
nand U26590 (N_26590,N_20253,N_20681);
nand U26591 (N_26591,N_21144,N_23505);
nor U26592 (N_26592,N_22563,N_20953);
nor U26593 (N_26593,N_22609,N_23945);
nor U26594 (N_26594,N_24625,N_20940);
nand U26595 (N_26595,N_22572,N_20282);
nand U26596 (N_26596,N_22721,N_20525);
nand U26597 (N_26597,N_23018,N_22909);
and U26598 (N_26598,N_22373,N_22781);
xnor U26599 (N_26599,N_24398,N_21742);
and U26600 (N_26600,N_24235,N_24162);
and U26601 (N_26601,N_21194,N_23422);
xor U26602 (N_26602,N_20348,N_21825);
xnor U26603 (N_26603,N_23752,N_21960);
nand U26604 (N_26604,N_20799,N_20902);
nand U26605 (N_26605,N_22891,N_22112);
or U26606 (N_26606,N_23107,N_22685);
xnor U26607 (N_26607,N_23341,N_24614);
nand U26608 (N_26608,N_23421,N_24181);
or U26609 (N_26609,N_22419,N_22081);
and U26610 (N_26610,N_22506,N_23868);
xor U26611 (N_26611,N_21283,N_24922);
or U26612 (N_26612,N_24886,N_20329);
nand U26613 (N_26613,N_24039,N_20774);
nand U26614 (N_26614,N_22505,N_22234);
xor U26615 (N_26615,N_21589,N_24544);
nand U26616 (N_26616,N_24078,N_21104);
or U26617 (N_26617,N_23066,N_23244);
nor U26618 (N_26618,N_23906,N_20140);
xor U26619 (N_26619,N_23635,N_22959);
nand U26620 (N_26620,N_21733,N_23958);
xnor U26621 (N_26621,N_22608,N_23839);
nand U26622 (N_26622,N_20089,N_20166);
nand U26623 (N_26623,N_23498,N_23936);
nor U26624 (N_26624,N_24663,N_20566);
xnor U26625 (N_26625,N_23900,N_20302);
or U26626 (N_26626,N_24364,N_21985);
nor U26627 (N_26627,N_21777,N_22150);
nand U26628 (N_26628,N_24781,N_22807);
nand U26629 (N_26629,N_21368,N_24624);
nand U26630 (N_26630,N_24418,N_21501);
or U26631 (N_26631,N_21119,N_23106);
nand U26632 (N_26632,N_24117,N_21372);
and U26633 (N_26633,N_20491,N_23239);
nand U26634 (N_26634,N_21107,N_24037);
nor U26635 (N_26635,N_20077,N_21566);
and U26636 (N_26636,N_22558,N_21031);
and U26637 (N_26637,N_23803,N_20987);
and U26638 (N_26638,N_23406,N_20636);
nand U26639 (N_26639,N_23004,N_23860);
or U26640 (N_26640,N_24239,N_20383);
xor U26641 (N_26641,N_24423,N_20446);
or U26642 (N_26642,N_21056,N_23399);
nand U26643 (N_26643,N_22288,N_20985);
xnor U26644 (N_26644,N_23383,N_20160);
nand U26645 (N_26645,N_24952,N_22786);
xnor U26646 (N_26646,N_24255,N_24904);
or U26647 (N_26647,N_20000,N_21834);
and U26648 (N_26648,N_20694,N_20139);
nor U26649 (N_26649,N_22096,N_21044);
or U26650 (N_26650,N_20722,N_24661);
or U26651 (N_26651,N_21302,N_22065);
nand U26652 (N_26652,N_24152,N_21034);
nor U26653 (N_26653,N_21308,N_21987);
nand U26654 (N_26654,N_23899,N_23521);
nand U26655 (N_26655,N_24620,N_21453);
and U26656 (N_26656,N_23673,N_22992);
xnor U26657 (N_26657,N_24843,N_20529);
nor U26658 (N_26658,N_20003,N_21765);
nor U26659 (N_26659,N_20577,N_21818);
and U26660 (N_26660,N_22176,N_21118);
nand U26661 (N_26661,N_24368,N_22132);
nand U26662 (N_26662,N_22745,N_24313);
and U26663 (N_26663,N_24823,N_24076);
and U26664 (N_26664,N_20876,N_24194);
and U26665 (N_26665,N_24085,N_21113);
nor U26666 (N_26666,N_21316,N_22611);
and U26667 (N_26667,N_22241,N_20321);
or U26668 (N_26668,N_20096,N_24799);
xor U26669 (N_26669,N_22021,N_22185);
xnor U26670 (N_26670,N_21183,N_22672);
or U26671 (N_26671,N_22223,N_22975);
nor U26672 (N_26672,N_20739,N_21218);
xnor U26673 (N_26673,N_21299,N_22845);
xnor U26674 (N_26674,N_21706,N_23047);
nor U26675 (N_26675,N_24399,N_20326);
xnor U26676 (N_26676,N_24582,N_22513);
or U26677 (N_26677,N_22899,N_22340);
nor U26678 (N_26678,N_23187,N_23596);
nand U26679 (N_26679,N_22659,N_24930);
or U26680 (N_26680,N_22874,N_20584);
and U26681 (N_26681,N_22656,N_23438);
xor U26682 (N_26682,N_24074,N_22877);
and U26683 (N_26683,N_22358,N_20200);
nor U26684 (N_26684,N_23604,N_22104);
and U26685 (N_26685,N_23300,N_23134);
or U26686 (N_26686,N_22181,N_21716);
xnor U26687 (N_26687,N_21386,N_21523);
xnor U26688 (N_26688,N_20398,N_24048);
nand U26689 (N_26689,N_20859,N_20269);
nand U26690 (N_26690,N_23727,N_20880);
or U26691 (N_26691,N_21804,N_23256);
and U26692 (N_26692,N_24224,N_20698);
and U26693 (N_26693,N_21879,N_21580);
nand U26694 (N_26694,N_22856,N_22588);
or U26695 (N_26695,N_22282,N_21139);
nor U26696 (N_26696,N_20049,N_21375);
and U26697 (N_26697,N_20981,N_20104);
or U26698 (N_26698,N_21049,N_23681);
or U26699 (N_26699,N_22942,N_22704);
xor U26700 (N_26700,N_23420,N_21356);
or U26701 (N_26701,N_22412,N_24068);
xor U26702 (N_26702,N_20274,N_21632);
and U26703 (N_26703,N_20413,N_24851);
or U26704 (N_26704,N_20011,N_20165);
xor U26705 (N_26705,N_24802,N_23697);
or U26706 (N_26706,N_22232,N_20609);
or U26707 (N_26707,N_21631,N_23737);
or U26708 (N_26708,N_21516,N_22010);
xor U26709 (N_26709,N_23609,N_24466);
nand U26710 (N_26710,N_24733,N_20073);
xor U26711 (N_26711,N_24335,N_24769);
and U26712 (N_26712,N_23033,N_22101);
xor U26713 (N_26713,N_21606,N_24946);
nor U26714 (N_26714,N_22520,N_22951);
and U26715 (N_26715,N_22564,N_23539);
nor U26716 (N_26716,N_24514,N_20945);
nor U26717 (N_26717,N_22860,N_23423);
or U26718 (N_26718,N_24748,N_24988);
xor U26719 (N_26719,N_21233,N_22395);
xnor U26720 (N_26720,N_20509,N_22503);
xor U26721 (N_26721,N_20766,N_22233);
nand U26722 (N_26722,N_24309,N_23124);
nor U26723 (N_26723,N_23997,N_20853);
and U26724 (N_26724,N_21919,N_23652);
nor U26725 (N_26725,N_20092,N_23288);
nand U26726 (N_26726,N_24163,N_22870);
and U26727 (N_26727,N_24501,N_24670);
xor U26728 (N_26728,N_24891,N_24846);
xor U26729 (N_26729,N_21883,N_22370);
nor U26730 (N_26730,N_22404,N_21336);
xor U26731 (N_26731,N_22540,N_24406);
and U26732 (N_26732,N_23375,N_24138);
or U26733 (N_26733,N_20432,N_22938);
xnor U26734 (N_26734,N_23049,N_20418);
nand U26735 (N_26735,N_21412,N_23598);
nor U26736 (N_26736,N_24139,N_20071);
or U26737 (N_26737,N_23208,N_21760);
nor U26738 (N_26738,N_23201,N_24061);
or U26739 (N_26739,N_24905,N_20594);
and U26740 (N_26740,N_23177,N_22547);
xnor U26741 (N_26741,N_24156,N_20546);
nand U26742 (N_26742,N_22986,N_24407);
xnor U26743 (N_26743,N_24741,N_20936);
xnor U26744 (N_26744,N_22586,N_24284);
or U26745 (N_26745,N_21521,N_24286);
nor U26746 (N_26746,N_24561,N_23826);
nor U26747 (N_26747,N_22508,N_23671);
nor U26748 (N_26748,N_23844,N_21036);
nor U26749 (N_26749,N_24911,N_22257);
nor U26750 (N_26750,N_23777,N_20085);
nor U26751 (N_26751,N_22249,N_20120);
xor U26752 (N_26752,N_22325,N_23944);
nand U26753 (N_26753,N_20938,N_20247);
or U26754 (N_26754,N_23607,N_21947);
nor U26755 (N_26755,N_22070,N_21668);
xor U26756 (N_26756,N_22008,N_21779);
nor U26757 (N_26757,N_23615,N_22955);
nor U26758 (N_26758,N_20224,N_23235);
nand U26759 (N_26759,N_20328,N_21833);
and U26760 (N_26760,N_23733,N_21131);
xor U26761 (N_26761,N_20659,N_24149);
or U26762 (N_26762,N_24527,N_22788);
nor U26763 (N_26763,N_23131,N_20183);
xnor U26764 (N_26764,N_23895,N_24990);
nand U26765 (N_26765,N_23443,N_20952);
or U26766 (N_26766,N_24593,N_23869);
and U26767 (N_26767,N_24098,N_21849);
or U26768 (N_26768,N_24861,N_21882);
xor U26769 (N_26769,N_24001,N_23656);
nand U26770 (N_26770,N_22007,N_22668);
or U26771 (N_26771,N_20911,N_23570);
nor U26772 (N_26772,N_24848,N_24275);
xor U26773 (N_26773,N_24369,N_23633);
nand U26774 (N_26774,N_24354,N_24053);
or U26775 (N_26775,N_22792,N_22810);
and U26776 (N_26776,N_21125,N_24521);
nor U26777 (N_26777,N_22278,N_23432);
nand U26778 (N_26778,N_22177,N_23077);
and U26779 (N_26779,N_22263,N_22368);
xor U26780 (N_26780,N_23419,N_20229);
xnor U26781 (N_26781,N_20006,N_24010);
nand U26782 (N_26782,N_24340,N_24189);
or U26783 (N_26783,N_20187,N_21507);
nor U26784 (N_26784,N_24912,N_24570);
xor U26785 (N_26785,N_20056,N_20493);
or U26786 (N_26786,N_22041,N_20299);
xnor U26787 (N_26787,N_21068,N_22748);
nand U26788 (N_26788,N_23120,N_22813);
nand U26789 (N_26789,N_23059,N_21101);
nand U26790 (N_26790,N_23591,N_22366);
xnor U26791 (N_26791,N_22309,N_23870);
and U26792 (N_26792,N_20132,N_20697);
xor U26793 (N_26793,N_20995,N_23522);
nor U26794 (N_26794,N_20173,N_20351);
or U26795 (N_26795,N_22655,N_24655);
nand U26796 (N_26796,N_23417,N_23433);
and U26797 (N_26797,N_20769,N_20337);
nor U26798 (N_26798,N_20226,N_22390);
nor U26799 (N_26799,N_21970,N_23754);
nor U26800 (N_26800,N_21678,N_21417);
xnor U26801 (N_26801,N_22768,N_21323);
nor U26802 (N_26802,N_22718,N_24025);
nor U26803 (N_26803,N_22092,N_24107);
xor U26804 (N_26804,N_20180,N_21249);
and U26805 (N_26805,N_21712,N_22590);
and U26806 (N_26806,N_22495,N_22189);
nand U26807 (N_26807,N_20735,N_22235);
xnor U26808 (N_26808,N_22140,N_22136);
xor U26809 (N_26809,N_20430,N_22399);
xnor U26810 (N_26810,N_24221,N_22743);
nand U26811 (N_26811,N_23327,N_20267);
and U26812 (N_26812,N_24266,N_21129);
nand U26813 (N_26813,N_23677,N_21268);
or U26814 (N_26814,N_20835,N_22598);
nor U26815 (N_26815,N_21052,N_20201);
nor U26816 (N_26816,N_20770,N_23846);
or U26817 (N_26817,N_23103,N_22794);
xnor U26818 (N_26818,N_21230,N_24985);
and U26819 (N_26819,N_23010,N_23110);
or U26820 (N_26820,N_23666,N_24635);
xor U26821 (N_26821,N_24708,N_23676);
or U26822 (N_26822,N_24847,N_23081);
or U26823 (N_26823,N_22643,N_21717);
xnor U26824 (N_26824,N_24026,N_23226);
xor U26825 (N_26825,N_21727,N_24487);
nand U26826 (N_26826,N_24927,N_23512);
nand U26827 (N_26827,N_21284,N_24808);
and U26828 (N_26828,N_23500,N_24673);
nand U26829 (N_26829,N_21858,N_20520);
and U26830 (N_26830,N_24096,N_23792);
or U26831 (N_26831,N_21983,N_24226);
and U26832 (N_26832,N_23323,N_22715);
or U26833 (N_26833,N_23153,N_20223);
and U26834 (N_26834,N_20578,N_22783);
and U26835 (N_26835,N_24525,N_21863);
nor U26836 (N_26836,N_21810,N_21638);
or U26837 (N_26837,N_21255,N_21744);
and U26838 (N_26838,N_20920,N_22167);
xor U26839 (N_26839,N_21010,N_21100);
xor U26840 (N_26840,N_21428,N_24551);
nand U26841 (N_26841,N_21366,N_21691);
nand U26842 (N_26842,N_24999,N_20532);
nand U26843 (N_26843,N_21080,N_21445);
or U26844 (N_26844,N_21776,N_21978);
xor U26845 (N_26845,N_23805,N_22103);
nor U26846 (N_26846,N_20150,N_20191);
or U26847 (N_26847,N_22597,N_23052);
and U26848 (N_26848,N_21751,N_23166);
or U26849 (N_26849,N_22785,N_21315);
nand U26850 (N_26850,N_20046,N_21327);
xnor U26851 (N_26851,N_21994,N_24653);
nand U26852 (N_26852,N_22073,N_23469);
and U26853 (N_26853,N_21134,N_23621);
and U26854 (N_26854,N_23394,N_20022);
xnor U26855 (N_26855,N_20803,N_22981);
or U26856 (N_26856,N_22491,N_23464);
xor U26857 (N_26857,N_21979,N_23907);
xor U26858 (N_26858,N_24082,N_23045);
and U26859 (N_26859,N_20461,N_22119);
nand U26860 (N_26860,N_24509,N_22690);
and U26861 (N_26861,N_24615,N_23003);
nor U26862 (N_26862,N_21458,N_22749);
and U26863 (N_26863,N_22524,N_23113);
and U26864 (N_26864,N_21939,N_22444);
and U26865 (N_26865,N_20693,N_24776);
xnor U26866 (N_26866,N_22440,N_24253);
and U26867 (N_26867,N_24924,N_21229);
and U26868 (N_26868,N_21020,N_22681);
and U26869 (N_26869,N_24819,N_20638);
or U26870 (N_26870,N_21655,N_22848);
or U26871 (N_26871,N_22782,N_21317);
nor U26872 (N_26872,N_21899,N_24376);
or U26873 (N_26873,N_21552,N_20449);
or U26874 (N_26874,N_23786,N_23513);
nand U26875 (N_26875,N_24400,N_20101);
nand U26876 (N_26876,N_22711,N_21739);
xor U26877 (N_26877,N_20709,N_23904);
nand U26878 (N_26878,N_21084,N_23566);
or U26879 (N_26879,N_20990,N_23152);
xnor U26880 (N_26880,N_22477,N_24672);
xor U26881 (N_26881,N_20884,N_23996);
nand U26882 (N_26882,N_22356,N_20934);
nand U26883 (N_26883,N_21838,N_22703);
or U26884 (N_26884,N_24237,N_21089);
or U26885 (N_26885,N_20186,N_24343);
nand U26886 (N_26886,N_21073,N_22152);
and U26887 (N_26887,N_23721,N_20467);
and U26888 (N_26888,N_24077,N_22110);
nor U26889 (N_26889,N_22881,N_23339);
or U26890 (N_26890,N_23690,N_20324);
xnor U26891 (N_26891,N_22313,N_20294);
xor U26892 (N_26892,N_20792,N_23198);
and U26893 (N_26893,N_22797,N_20728);
or U26894 (N_26894,N_20443,N_21383);
and U26895 (N_26895,N_21463,N_23388);
and U26896 (N_26896,N_20345,N_24351);
xnor U26897 (N_26897,N_23095,N_20537);
or U26898 (N_26898,N_22303,N_20154);
nor U26899 (N_26899,N_20704,N_21490);
or U26900 (N_26900,N_23236,N_24145);
xor U26901 (N_26901,N_21140,N_20593);
and U26902 (N_26902,N_21062,N_23373);
or U26903 (N_26903,N_22184,N_24906);
nand U26904 (N_26904,N_22391,N_21570);
or U26905 (N_26905,N_24394,N_24716);
and U26906 (N_26906,N_22194,N_23109);
or U26907 (N_26907,N_20335,N_23155);
nand U26908 (N_26908,N_22218,N_22752);
nor U26909 (N_26909,N_21432,N_24119);
xor U26910 (N_26910,N_20805,N_21274);
nand U26911 (N_26911,N_24115,N_23741);
nand U26912 (N_26912,N_24438,N_23454);
and U26913 (N_26913,N_20786,N_24646);
xor U26914 (N_26914,N_20779,N_21422);
and U26915 (N_26915,N_24207,N_23253);
and U26916 (N_26916,N_20660,N_20524);
nand U26917 (N_26917,N_20662,N_22545);
and U26918 (N_26918,N_24796,N_20585);
nand U26919 (N_26919,N_24289,N_24473);
xnor U26920 (N_26920,N_20479,N_20189);
or U26921 (N_26921,N_22225,N_22979);
nor U26922 (N_26922,N_22275,N_23818);
nor U26923 (N_26923,N_22394,N_21017);
and U26924 (N_26924,N_24564,N_20275);
nor U26925 (N_26925,N_21598,N_20893);
xnor U26926 (N_26926,N_20462,N_24757);
xnor U26927 (N_26927,N_23098,N_21177);
nor U26928 (N_26928,N_24477,N_21505);
nor U26929 (N_26929,N_23453,N_22255);
nor U26930 (N_26930,N_23407,N_23287);
and U26931 (N_26931,N_20900,N_23401);
nand U26932 (N_26932,N_24632,N_21310);
or U26933 (N_26933,N_23580,N_23935);
nor U26934 (N_26934,N_23447,N_21576);
nand U26935 (N_26935,N_20622,N_20897);
nand U26936 (N_26936,N_20234,N_21596);
nand U26937 (N_26937,N_23460,N_22031);
nand U26938 (N_26938,N_24031,N_23682);
nor U26939 (N_26939,N_20871,N_21723);
nor U26940 (N_26940,N_23275,N_23167);
nor U26941 (N_26941,N_21926,N_21915);
xnor U26942 (N_26942,N_22838,N_22163);
and U26943 (N_26943,N_21791,N_21369);
nor U26944 (N_26944,N_23140,N_21799);
and U26945 (N_26945,N_24678,N_22566);
xor U26946 (N_26946,N_24408,N_24465);
and U26947 (N_26947,N_22467,N_22384);
xor U26948 (N_26948,N_21758,N_22056);
nand U26949 (N_26949,N_24845,N_22779);
xor U26950 (N_26950,N_21241,N_20519);
xnor U26951 (N_26951,N_22769,N_24257);
xor U26952 (N_26952,N_24000,N_22551);
xor U26953 (N_26953,N_24055,N_21649);
nor U26954 (N_26954,N_22067,N_20163);
nor U26955 (N_26955,N_23645,N_24629);
nand U26956 (N_26956,N_20145,N_24269);
nand U26957 (N_26957,N_23342,N_20674);
and U26958 (N_26958,N_24511,N_22726);
nand U26959 (N_26959,N_23616,N_21646);
and U26960 (N_26960,N_24674,N_24325);
nand U26961 (N_26961,N_24311,N_23657);
or U26962 (N_26962,N_23013,N_21276);
nand U26963 (N_26963,N_21314,N_22281);
or U26964 (N_26964,N_24837,N_24571);
nor U26965 (N_26965,N_24479,N_22365);
or U26966 (N_26966,N_24996,N_21801);
nor U26967 (N_26967,N_22811,N_23872);
or U26968 (N_26968,N_20624,N_23072);
nor U26969 (N_26969,N_23309,N_20382);
nand U26970 (N_26970,N_20729,N_24493);
and U26971 (N_26971,N_21395,N_21661);
or U26972 (N_26972,N_21207,N_23437);
nand U26973 (N_26973,N_20605,N_23664);
or U26974 (N_26974,N_23418,N_24739);
xnor U26975 (N_26975,N_23882,N_22091);
nor U26976 (N_26976,N_21474,N_22017);
xor U26977 (N_26977,N_24170,N_24080);
or U26978 (N_26978,N_24328,N_23009);
and U26979 (N_26979,N_20590,N_23079);
or U26980 (N_26980,N_23405,N_20106);
xor U26981 (N_26981,N_23926,N_22198);
nor U26982 (N_26982,N_20817,N_23032);
nor U26983 (N_26983,N_20797,N_21105);
nor U26984 (N_26984,N_21755,N_21821);
nor U26985 (N_26985,N_20923,N_24966);
xnor U26986 (N_26986,N_23144,N_23183);
or U26987 (N_26987,N_22902,N_21115);
nor U26988 (N_26988,N_24256,N_23206);
and U26989 (N_26989,N_20211,N_23364);
xor U26990 (N_26990,N_20485,N_21288);
nor U26991 (N_26991,N_20810,N_21778);
and U26992 (N_26992,N_24070,N_24106);
and U26993 (N_26993,N_20306,N_22227);
nand U26994 (N_26994,N_24166,N_21910);
or U26995 (N_26995,N_20147,N_22616);
nor U26996 (N_26996,N_20252,N_21940);
nor U26997 (N_26997,N_21418,N_22079);
nand U26998 (N_26998,N_21662,N_23233);
nand U26999 (N_26999,N_23892,N_21869);
nand U27000 (N_27000,N_24450,N_24601);
nand U27001 (N_27001,N_20540,N_23273);
xor U27002 (N_27002,N_21179,N_24267);
nor U27003 (N_27003,N_23628,N_22357);
nand U27004 (N_27004,N_23776,N_22183);
and U27005 (N_27005,N_24700,N_23068);
and U27006 (N_27006,N_24411,N_24360);
nand U27007 (N_27007,N_21656,N_21982);
nand U27008 (N_27008,N_21244,N_21605);
or U27009 (N_27009,N_24928,N_23186);
nand U27010 (N_27010,N_24691,N_20846);
nand U27011 (N_27011,N_24949,N_24169);
and U27012 (N_27012,N_24533,N_21511);
nand U27013 (N_27013,N_24499,N_23753);
nor U27014 (N_27014,N_20456,N_20521);
nor U27015 (N_27015,N_24714,N_24141);
or U27016 (N_27016,N_22134,N_22571);
nor U27017 (N_27017,N_21399,N_20377);
nand U27018 (N_27018,N_20138,N_24542);
or U27019 (N_27019,N_24569,N_23987);
or U27020 (N_27020,N_21069,N_24387);
xor U27021 (N_27021,N_23371,N_21352);
xor U27022 (N_27022,N_21571,N_22581);
xnor U27023 (N_27023,N_21651,N_24574);
nand U27024 (N_27024,N_20855,N_21426);
xnor U27025 (N_27025,N_21141,N_23613);
or U27026 (N_27026,N_20903,N_22778);
nor U27027 (N_27027,N_20416,N_21054);
or U27028 (N_27028,N_24703,N_24558);
and U27029 (N_27029,N_22435,N_23265);
nand U27030 (N_27030,N_23592,N_21826);
nor U27031 (N_27031,N_20027,N_21188);
nand U27032 (N_27032,N_23142,N_20796);
or U27033 (N_27033,N_23543,N_20167);
or U27034 (N_27034,N_22299,N_20367);
nor U27035 (N_27035,N_22661,N_20386);
nor U27036 (N_27036,N_24035,N_21402);
xor U27037 (N_27037,N_22042,N_20784);
nor U27038 (N_27038,N_20772,N_22029);
nor U27039 (N_27039,N_20665,N_23828);
or U27040 (N_27040,N_24567,N_21264);
nand U27041 (N_27041,N_21492,N_24800);
xnor U27042 (N_27042,N_24517,N_23510);
nand U27043 (N_27043,N_20378,N_21513);
or U27044 (N_27044,N_24929,N_20237);
or U27045 (N_27045,N_21974,N_22496);
nand U27046 (N_27046,N_24709,N_23116);
or U27047 (N_27047,N_22210,N_23225);
xor U27048 (N_27048,N_22888,N_22636);
or U27049 (N_27049,N_20942,N_21066);
and U27050 (N_27050,N_24850,N_23586);
nor U27051 (N_27051,N_20877,N_21451);
and U27052 (N_27052,N_23133,N_22165);
xor U27053 (N_27053,N_24871,N_24957);
nand U27054 (N_27054,N_21078,N_23227);
nand U27055 (N_27055,N_20325,N_24613);
or U27056 (N_27056,N_23626,N_21446);
xnor U27057 (N_27057,N_24317,N_21180);
nor U27058 (N_27058,N_22355,N_23455);
xor U27059 (N_27059,N_20683,N_23002);
nor U27060 (N_27060,N_23019,N_23946);
or U27061 (N_27061,N_22228,N_24877);
or U27062 (N_27062,N_21075,N_24923);
or U27063 (N_27063,N_23694,N_21620);
nor U27064 (N_27064,N_22063,N_20067);
or U27065 (N_27065,N_22940,N_23974);
and U27066 (N_27066,N_24734,N_24274);
and U27067 (N_27067,N_24320,N_20322);
and U27068 (N_27068,N_22345,N_20512);
nand U27069 (N_27069,N_22995,N_21681);
nor U27070 (N_27070,N_21392,N_23263);
or U27071 (N_27071,N_24901,N_24684);
or U27072 (N_27072,N_21558,N_21875);
and U27073 (N_27073,N_22699,N_22192);
nor U27074 (N_27074,N_24095,N_23703);
xor U27075 (N_27075,N_24401,N_24505);
nor U27076 (N_27076,N_23099,N_21586);
or U27077 (N_27077,N_21335,N_22632);
nand U27078 (N_27078,N_24122,N_21921);
or U27079 (N_27079,N_24545,N_23111);
or U27080 (N_27080,N_20941,N_24230);
xor U27081 (N_27081,N_24829,N_23930);
xor U27082 (N_27082,N_21772,N_22766);
xnor U27083 (N_27083,N_20123,N_24961);
xor U27084 (N_27084,N_21736,N_22678);
and U27085 (N_27085,N_20359,N_20678);
and U27086 (N_27086,N_23661,N_20298);
nor U27087 (N_27087,N_24338,N_24559);
or U27088 (N_27088,N_22701,N_21137);
or U27089 (N_27089,N_24667,N_22700);
nand U27090 (N_27090,N_22014,N_21770);
xnor U27091 (N_27091,N_23530,N_20159);
nand U27092 (N_27092,N_21684,N_21824);
nand U27093 (N_27093,N_23686,N_23026);
nand U27094 (N_27094,N_23911,N_24715);
and U27095 (N_27095,N_20356,N_21556);
nand U27096 (N_27096,N_23154,N_22958);
and U27097 (N_27097,N_20619,N_20564);
nand U27098 (N_27098,N_21850,N_22863);
nor U27099 (N_27099,N_23625,N_22650);
xor U27100 (N_27100,N_24751,N_21715);
and U27101 (N_27101,N_22937,N_22756);
and U27102 (N_27102,N_21450,N_24315);
xor U27103 (N_27103,N_21697,N_21224);
xor U27104 (N_27104,N_21205,N_20539);
nand U27105 (N_27105,N_23758,N_20703);
nand U27106 (N_27106,N_23151,N_23527);
nor U27107 (N_27107,N_23281,N_23316);
nand U27108 (N_27108,N_21687,N_23162);
nor U27109 (N_27109,N_24628,N_24045);
or U27110 (N_27110,N_22720,N_22016);
nand U27111 (N_27111,N_21931,N_24234);
xor U27112 (N_27112,N_20909,N_21124);
xor U27113 (N_27113,N_21968,N_20647);
xor U27114 (N_27114,N_23897,N_22575);
xnor U27115 (N_27115,N_22689,N_22944);
and U27116 (N_27116,N_20657,N_21208);
or U27117 (N_27117,N_24120,N_24753);
and U27118 (N_27118,N_22135,N_22259);
nand U27119 (N_27119,N_24630,N_20964);
nand U27120 (N_27120,N_24775,N_20079);
xnor U27121 (N_27121,N_20925,N_23642);
nand U27122 (N_27122,N_20013,N_22772);
nor U27123 (N_27123,N_20421,N_20568);
nor U27124 (N_27124,N_23360,N_24627);
nor U27125 (N_27125,N_23573,N_22078);
nand U27126 (N_27126,N_20986,N_21482);
nor U27127 (N_27127,N_23749,N_21184);
and U27128 (N_27128,N_21329,N_22295);
and U27129 (N_27129,N_23942,N_21480);
nand U27130 (N_27130,N_23745,N_21401);
nor U27131 (N_27131,N_22854,N_20929);
or U27132 (N_27132,N_22009,N_23732);
or U27133 (N_27133,N_20477,N_20009);
xor U27134 (N_27134,N_23585,N_22631);
nor U27135 (N_27135,N_20075,N_24666);
nand U27136 (N_27136,N_21235,N_23951);
or U27137 (N_27137,N_23076,N_20999);
and U27138 (N_27138,N_22773,N_20213);
or U27139 (N_27139,N_20838,N_21629);
nor U27140 (N_27140,N_24535,N_21679);
and U27141 (N_27141,N_21977,N_24279);
xnor U27142 (N_27142,N_23195,N_20975);
xor U27143 (N_27143,N_24768,N_22555);
nor U27144 (N_27144,N_22858,N_24771);
xnor U27145 (N_27145,N_22649,N_24378);
nor U27146 (N_27146,N_24788,N_22734);
nor U27147 (N_27147,N_24285,N_20544);
and U27148 (N_27148,N_22666,N_21707);
or U27149 (N_27149,N_21563,N_21998);
or U27150 (N_27150,N_24132,N_20548);
and U27151 (N_27151,N_24075,N_21878);
or U27152 (N_27152,N_22945,N_22256);
and U27153 (N_27153,N_22867,N_21239);
or U27154 (N_27154,N_20314,N_24482);
nor U27155 (N_27155,N_22291,N_23007);
xnor U27156 (N_27156,N_24468,N_24058);
nor U27157 (N_27157,N_22947,N_23989);
and U27158 (N_27158,N_24590,N_23434);
nor U27159 (N_27159,N_21408,N_21041);
xnor U27160 (N_27160,N_20924,N_22472);
nand U27161 (N_27161,N_21491,N_22108);
or U27162 (N_27162,N_21187,N_20313);
or U27163 (N_27163,N_23248,N_22094);
or U27164 (N_27164,N_20666,N_20176);
xor U27165 (N_27165,N_24032,N_23311);
xnor U27166 (N_27166,N_20060,N_22069);
nor U27167 (N_27167,N_23348,N_22816);
and U27168 (N_27168,N_20827,N_21746);
nand U27169 (N_27169,N_23257,N_24276);
and U27170 (N_27170,N_23355,N_23096);
nor U27171 (N_27171,N_20644,N_23611);
and U27172 (N_27172,N_21975,N_24412);
nor U27173 (N_27173,N_23286,N_21675);
nor U27174 (N_27174,N_22420,N_21116);
or U27175 (N_27175,N_20634,N_21846);
nand U27176 (N_27176,N_22642,N_21625);
nor U27177 (N_27177,N_24046,N_23242);
and U27178 (N_27178,N_23395,N_24767);
nor U27179 (N_27179,N_22911,N_21063);
nor U27180 (N_27180,N_20598,N_24210);
and U27181 (N_27181,N_22988,N_22097);
xnor U27182 (N_27182,N_24972,N_24764);
nand U27183 (N_27183,N_22448,N_23660);
or U27184 (N_27184,N_24959,N_24327);
or U27185 (N_27185,N_21250,N_22455);
nor U27186 (N_27186,N_24405,N_22090);
and U27187 (N_27187,N_21162,N_22260);
xnor U27188 (N_27188,N_20197,N_21506);
or U27189 (N_27189,N_20700,N_24754);
and U27190 (N_27190,N_23528,N_23220);
or U27191 (N_27191,N_23319,N_22402);
nor U27192 (N_27192,N_20707,N_20870);
xnor U27193 (N_27193,N_21641,N_21637);
xor U27194 (N_27194,N_21011,N_20557);
xor U27195 (N_27195,N_23150,N_22731);
and U27196 (N_27196,N_22804,N_22248);
and U27197 (N_27197,N_20959,N_21420);
and U27198 (N_27198,N_22595,N_23922);
nor U27199 (N_27199,N_24016,N_23119);
and U27200 (N_27200,N_23933,N_22767);
nand U27201 (N_27201,N_23413,N_22832);
xor U27202 (N_27202,N_23097,N_20961);
or U27203 (N_27203,N_21429,N_20330);
nand U27204 (N_27204,N_21916,N_21197);
or U27205 (N_27205,N_20070,N_22283);
and U27206 (N_27206,N_20573,N_21722);
nor U27207 (N_27207,N_24431,N_23213);
xor U27208 (N_27208,N_20699,N_23518);
or U27209 (N_27209,N_20500,N_23393);
nor U27210 (N_27210,N_24133,N_23021);
xor U27211 (N_27211,N_23382,N_21842);
xnor U27212 (N_27212,N_20212,N_22222);
or U27213 (N_27213,N_24973,N_21130);
or U27214 (N_27214,N_23427,N_22289);
and U27215 (N_27215,N_24797,N_22466);
or U27216 (N_27216,N_21260,N_24326);
xor U27217 (N_27217,N_20771,N_23204);
nand U27218 (N_27218,N_20574,N_23931);
and U27219 (N_27219,N_20358,N_24965);
or U27220 (N_27220,N_21286,N_24898);
xnor U27221 (N_27221,N_20632,N_21699);
or U27222 (N_27222,N_24209,N_20439);
and U27223 (N_27223,N_22989,N_20347);
and U27224 (N_27224,N_22895,N_24616);
xor U27225 (N_27225,N_22852,N_22157);
or U27226 (N_27226,N_20958,N_21127);
xor U27227 (N_27227,N_21663,N_24964);
xor U27228 (N_27228,N_23397,N_24943);
nor U27229 (N_27229,N_23255,N_24651);
xnor U27230 (N_27230,N_20292,N_23948);
and U27231 (N_27231,N_23984,N_20097);
xor U27232 (N_27232,N_20572,N_20450);
and U27233 (N_27233,N_21743,N_23730);
and U27234 (N_27234,N_23125,N_24467);
or U27235 (N_27235,N_22059,N_23336);
and U27236 (N_27236,N_22674,N_23934);
or U27237 (N_27237,N_20505,N_20380);
and U27238 (N_27238,N_21710,N_22306);
nand U27239 (N_27239,N_20621,N_21793);
or U27240 (N_27240,N_23534,N_24969);
nor U27241 (N_27241,N_21913,N_22338);
nand U27242 (N_27242,N_20270,N_20207);
xor U27243 (N_27243,N_20455,N_24968);
xor U27244 (N_27244,N_21601,N_22434);
nor U27245 (N_27245,N_23304,N_21683);
and U27246 (N_27246,N_24857,N_21564);
nor U27247 (N_27247,N_23834,N_22964);
nand U27248 (N_27248,N_24108,N_21647);
nor U27249 (N_27249,N_23231,N_24807);
nand U27250 (N_27250,N_21487,N_22829);
nor U27251 (N_27251,N_21532,N_21157);
nor U27252 (N_27252,N_22751,N_23410);
xor U27253 (N_27253,N_21343,N_21635);
or U27254 (N_27254,N_21339,N_23485);
and U27255 (N_27255,N_22828,N_22954);
nand U27256 (N_27256,N_23909,N_21938);
nor U27257 (N_27257,N_21711,N_23249);
nor U27258 (N_27258,N_23643,N_22796);
and U27259 (N_27259,N_21531,N_20142);
xnor U27260 (N_27260,N_24728,N_20192);
or U27261 (N_27261,N_21984,N_23569);
or U27262 (N_27262,N_21122,N_22510);
nand U27263 (N_27263,N_21156,N_23599);
or U27264 (N_27264,N_22153,N_24790);
nor U27265 (N_27265,N_24490,N_20811);
nor U27266 (N_27266,N_20654,N_23091);
and U27267 (N_27267,N_20714,N_20021);
and U27268 (N_27268,N_22667,N_23390);
and U27269 (N_27269,N_22663,N_24215);
and U27270 (N_27270,N_20793,N_22620);
nand U27271 (N_27271,N_23667,N_24833);
nor U27272 (N_27272,N_22433,N_24811);
and U27273 (N_27273,N_24603,N_20974);
xor U27274 (N_27274,N_20571,N_21542);
or U27275 (N_27275,N_24662,N_21258);
nor U27276 (N_27276,N_23701,N_20100);
or U27277 (N_27277,N_23365,N_23972);
xnor U27278 (N_27278,N_22221,N_20675);
xor U27279 (N_27279,N_23851,N_21865);
nand U27280 (N_27280,N_21081,N_24858);
xor U27281 (N_27281,N_24051,N_24752);
nor U27282 (N_27282,N_24863,N_21759);
nor U27283 (N_27283,N_22426,N_23358);
and U27284 (N_27284,N_22622,N_20005);
nor U27285 (N_27285,N_23191,N_24131);
or U27286 (N_27286,N_21000,N_21273);
and U27287 (N_27287,N_23250,N_23174);
nor U27288 (N_27288,N_21988,N_23819);
xor U27289 (N_27289,N_23810,N_24572);
nand U27290 (N_27290,N_20065,N_22120);
xor U27291 (N_27291,N_23836,N_24869);
nand U27292 (N_27292,N_21616,N_20216);
nand U27293 (N_27293,N_24183,N_20202);
nor U27294 (N_27294,N_21805,N_22003);
nor U27295 (N_27295,N_23551,N_22193);
xnor U27296 (N_27296,N_23011,N_24654);
nor U27297 (N_27297,N_23675,N_24485);
nor U27298 (N_27298,N_24469,N_22262);
xnor U27299 (N_27299,N_24484,N_20604);
or U27300 (N_27300,N_21254,N_22187);
and U27301 (N_27301,N_23515,N_24281);
nor U27302 (N_27302,N_20209,N_21912);
and U27303 (N_27303,N_22866,N_21030);
or U27304 (N_27304,N_21588,N_23158);
and U27305 (N_27305,N_20676,N_24756);
and U27306 (N_27306,N_23370,N_21514);
and U27307 (N_27307,N_24213,N_20354);
nor U27308 (N_27308,N_20763,N_21381);
nor U27309 (N_27309,N_24013,N_20063);
nand U27310 (N_27310,N_23060,N_20689);
or U27311 (N_27311,N_24165,N_20019);
xor U27312 (N_27312,N_20740,N_21517);
nor U27313 (N_27313,N_23957,N_23347);
or U27314 (N_27314,N_21311,N_23449);
nor U27315 (N_27315,N_21086,N_21425);
nand U27316 (N_27316,N_22240,N_22647);
and U27317 (N_27317,N_23788,N_24358);
nand U27318 (N_27318,N_23544,N_20179);
nor U27319 (N_27319,N_21238,N_24792);
or U27320 (N_27320,N_20854,N_24111);
nand U27321 (N_27321,N_20355,N_20219);
or U27322 (N_27322,N_22264,N_24738);
xor U27323 (N_27323,N_20813,N_21263);
or U27324 (N_27324,N_23555,N_21076);
nand U27325 (N_27325,N_21892,N_23654);
and U27326 (N_27326,N_23973,N_20677);
and U27327 (N_27327,N_24549,N_22660);
nand U27328 (N_27328,N_24937,N_20904);
or U27329 (N_27329,N_22095,N_22928);
nor U27330 (N_27330,N_24594,N_21886);
nand U27331 (N_27331,N_20350,N_22761);
nor U27332 (N_27332,N_20303,N_21815);
nor U27333 (N_27333,N_24188,N_24981);
and U27334 (N_27334,N_23440,N_24356);
and U27335 (N_27335,N_23783,N_20648);
nor U27336 (N_27336,N_20403,N_22462);
or U27337 (N_27337,N_20592,N_24671);
or U27338 (N_27338,N_22121,N_22560);
xnor U27339 (N_27339,N_24522,N_23949);
nand U27340 (N_27340,N_21109,N_24435);
xnor U27341 (N_27341,N_22006,N_21762);
or U27342 (N_27342,N_23015,N_24305);
nand U27343 (N_27343,N_20040,N_24510);
or U27344 (N_27344,N_23992,N_21893);
nand U27345 (N_27345,N_23328,N_21285);
nor U27346 (N_27346,N_21560,N_22648);
xor U27347 (N_27347,N_23896,N_22613);
and U27348 (N_27348,N_23630,N_20297);
nand U27349 (N_27349,N_20899,N_24523);
or U27350 (N_27350,N_24842,N_23251);
or U27351 (N_27351,N_20866,N_24168);
xnor U27352 (N_27352,N_20873,N_23557);
nand U27353 (N_27353,N_24444,N_22878);
or U27354 (N_27354,N_22061,N_23912);
xor U27355 (N_27355,N_23023,N_23600);
and U27356 (N_27356,N_23789,N_23456);
nand U27357 (N_27357,N_23494,N_24292);
nand U27358 (N_27358,N_22168,N_22758);
and U27359 (N_27359,N_21351,N_21045);
and U27360 (N_27360,N_20858,N_21126);
xor U27361 (N_27361,N_23629,N_24440);
nand U27362 (N_27362,N_21454,N_22924);
and U27363 (N_27363,N_23499,N_24580);
or U27364 (N_27364,N_23218,N_20885);
and U27365 (N_27365,N_20387,N_20057);
and U27366 (N_27366,N_22200,N_20808);
nand U27367 (N_27367,N_20721,N_24664);
or U27368 (N_27368,N_23597,N_21991);
or U27369 (N_27369,N_21911,N_20514);
nor U27370 (N_27370,N_23429,N_23104);
and U27371 (N_27371,N_22000,N_20673);
xnor U27372 (N_27372,N_20375,N_20108);
xnor U27373 (N_27373,N_20404,N_23143);
and U27374 (N_27374,N_21409,N_23234);
or U27375 (N_27375,N_23165,N_20921);
or U27376 (N_27376,N_24696,N_20748);
nor U27377 (N_27377,N_20182,N_20869);
nand U27378 (N_27378,N_22732,N_24330);
nand U27379 (N_27379,N_23970,N_22146);
and U27380 (N_27380,N_24094,N_23088);
nor U27381 (N_27381,N_24242,N_24040);
or U27382 (N_27382,N_20623,N_24879);
xor U27383 (N_27383,N_24212,N_24749);
and U27384 (N_27384,N_20731,N_23194);
nor U27385 (N_27385,N_22456,N_24693);
or U27386 (N_27386,N_21782,N_24951);
xor U27387 (N_27387,N_20016,N_22970);
nand U27388 (N_27388,N_20440,N_23424);
nor U27389 (N_27389,N_24576,N_21956);
nand U27390 (N_27390,N_20162,N_24841);
nand U27391 (N_27391,N_20361,N_24619);
xnor U27392 (N_27392,N_21478,N_20425);
or U27393 (N_27393,N_20363,N_20738);
and U27394 (N_27394,N_24500,N_23337);
nor U27395 (N_27395,N_22304,N_24889);
nor U27396 (N_27396,N_20851,N_23954);
or U27397 (N_27397,N_24319,N_22889);
nand U27398 (N_27398,N_24859,N_22760);
or U27399 (N_27399,N_21527,N_24036);
nor U27400 (N_27400,N_24346,N_21692);
nor U27401 (N_27401,N_23715,N_22671);
nor U27402 (N_27402,N_24129,N_20258);
and U27403 (N_27403,N_21135,N_21808);
and U27404 (N_27404,N_20600,N_24419);
nand U27405 (N_27405,N_23744,N_24568);
and U27406 (N_27406,N_24047,N_21562);
nor U27407 (N_27407,N_24831,N_21831);
nor U27408 (N_27408,N_22713,N_23230);
or U27409 (N_27409,N_23117,N_22806);
xor U27410 (N_27410,N_22776,N_24247);
nand U27411 (N_27411,N_21811,N_23589);
xnor U27412 (N_27412,N_21788,N_23939);
nor U27413 (N_27413,N_20407,N_24332);
xnor U27414 (N_27414,N_23396,N_24873);
nand U27415 (N_27415,N_23292,N_20629);
nor U27416 (N_27416,N_22601,N_20344);
xor U27417 (N_27417,N_24348,N_20464);
or U27418 (N_27418,N_23387,N_24413);
or U27419 (N_27419,N_21079,N_20420);
nor U27420 (N_27420,N_21763,N_23631);
xnor U27421 (N_27421,N_20819,N_22038);
and U27422 (N_27422,N_24251,N_23995);
nor U27423 (N_27423,N_23956,N_24452);
or U27424 (N_27424,N_23338,N_21040);
xor U27425 (N_27425,N_23196,N_23217);
xnor U27426 (N_27426,N_22892,N_20047);
xor U27427 (N_27427,N_24178,N_22133);
or U27428 (N_27428,N_21457,N_24839);
and U27429 (N_27429,N_20837,N_20872);
and U27430 (N_27430,N_24536,N_23108);
nor U27431 (N_27431,N_24057,N_22428);
and U27432 (N_27432,N_20653,N_23053);
nand U27433 (N_27433,N_20471,N_24874);
nor U27434 (N_27434,N_20630,N_22252);
nand U27435 (N_27435,N_23310,N_24130);
nand U27436 (N_27436,N_21547,N_22903);
and U27437 (N_27437,N_21851,N_20190);
nor U27438 (N_27438,N_23102,N_24689);
and U27439 (N_27439,N_22569,N_23668);
xnor U27440 (N_27440,N_20967,N_20687);
nand U27441 (N_27441,N_22086,N_24100);
xnor U27442 (N_27442,N_21955,N_24384);
and U27443 (N_27443,N_22724,N_22960);
nor U27444 (N_27444,N_22463,N_24838);
nand U27445 (N_27445,N_24271,N_20436);
or U27446 (N_27446,N_23209,N_20369);
or U27447 (N_27447,N_20372,N_24421);
nand U27448 (N_27448,N_20783,N_20711);
nor U27449 (N_27449,N_24528,N_22738);
xor U27450 (N_27450,N_24293,N_21577);
xor U27451 (N_27451,N_20915,N_23843);
xor U27452 (N_27452,N_21593,N_24009);
nand U27453 (N_27453,N_23386,N_23228);
nor U27454 (N_27454,N_20112,N_20507);
and U27455 (N_27455,N_20417,N_23284);
nor U27456 (N_27456,N_22098,N_24321);
xor U27457 (N_27457,N_20228,N_23699);
or U27458 (N_27458,N_20791,N_23488);
and U27459 (N_27459,N_24701,N_24770);
nand U27460 (N_27460,N_20822,N_23343);
or U27461 (N_27461,N_21848,N_24310);
xor U27462 (N_27462,N_22556,N_22214);
or U27463 (N_27463,N_20170,N_21508);
xor U27464 (N_27464,N_20385,N_20708);
and U27465 (N_27465,N_23282,N_23823);
and U27466 (N_27466,N_21464,N_24463);
and U27467 (N_27467,N_20261,N_24314);
or U27468 (N_27468,N_21313,N_24262);
xnor U27469 (N_27469,N_24623,N_23838);
and U27470 (N_27470,N_21509,N_20701);
nand U27471 (N_27471,N_22978,N_24772);
and U27472 (N_27472,N_23070,N_23901);
nor U27473 (N_27473,N_22799,N_24519);
or U27474 (N_27474,N_24573,N_21198);
and U27475 (N_27475,N_22579,N_21400);
or U27476 (N_27476,N_23276,N_24299);
and U27477 (N_27477,N_23567,N_22777);
nor U27478 (N_27478,N_23742,N_23651);
xor U27479 (N_27479,N_24202,N_21626);
nor U27480 (N_27480,N_21158,N_23827);
or U27481 (N_27481,N_24610,N_23692);
and U27482 (N_27482,N_22996,N_22375);
nand U27483 (N_27483,N_21318,N_24554);
and U27484 (N_27484,N_21058,N_23572);
or U27485 (N_27485,N_21294,N_21797);
or U27486 (N_27486,N_20078,N_21437);
xnor U27487 (N_27487,N_24127,N_24496);
and U27488 (N_27488,N_21296,N_23632);
nand U27489 (N_27489,N_22458,N_23005);
and U27490 (N_27490,N_20583,N_23468);
nor U27491 (N_27491,N_24228,N_22386);
and U27492 (N_27492,N_20265,N_22956);
xor U27493 (N_27493,N_22728,N_22085);
nor U27494 (N_27494,N_23380,N_24065);
xnor U27495 (N_27495,N_21164,N_22224);
xnor U27496 (N_27496,N_21932,N_23351);
nand U27497 (N_27497,N_20602,N_22916);
nand U27498 (N_27498,N_24878,N_20565);
xor U27499 (N_27499,N_21594,N_20850);
and U27500 (N_27500,N_23706,N_23099);
xnor U27501 (N_27501,N_21347,N_20487);
nor U27502 (N_27502,N_20891,N_22194);
xor U27503 (N_27503,N_22264,N_22192);
xnor U27504 (N_27504,N_24118,N_22858);
xor U27505 (N_27505,N_22689,N_24747);
xnor U27506 (N_27506,N_21693,N_24977);
or U27507 (N_27507,N_20049,N_24247);
xnor U27508 (N_27508,N_20033,N_24538);
nand U27509 (N_27509,N_22385,N_20738);
xor U27510 (N_27510,N_22019,N_21861);
or U27511 (N_27511,N_23389,N_20285);
and U27512 (N_27512,N_21611,N_21682);
nand U27513 (N_27513,N_24148,N_20224);
nor U27514 (N_27514,N_24418,N_20953);
and U27515 (N_27515,N_21618,N_20339);
nor U27516 (N_27516,N_21150,N_24088);
and U27517 (N_27517,N_23520,N_23988);
and U27518 (N_27518,N_24595,N_22825);
or U27519 (N_27519,N_20707,N_22420);
nor U27520 (N_27520,N_22525,N_22181);
nand U27521 (N_27521,N_24283,N_20653);
nor U27522 (N_27522,N_21594,N_21901);
nor U27523 (N_27523,N_24293,N_22186);
or U27524 (N_27524,N_22832,N_24267);
and U27525 (N_27525,N_24837,N_24595);
and U27526 (N_27526,N_22686,N_20174);
xnor U27527 (N_27527,N_22489,N_24339);
nor U27528 (N_27528,N_20951,N_23757);
or U27529 (N_27529,N_24815,N_24867);
nand U27530 (N_27530,N_21759,N_22036);
and U27531 (N_27531,N_21670,N_24953);
xor U27532 (N_27532,N_24748,N_21397);
nand U27533 (N_27533,N_24796,N_22253);
and U27534 (N_27534,N_24533,N_22612);
nand U27535 (N_27535,N_23566,N_22144);
and U27536 (N_27536,N_22337,N_24202);
xor U27537 (N_27537,N_21520,N_22224);
nand U27538 (N_27538,N_24757,N_24453);
nand U27539 (N_27539,N_20783,N_23948);
and U27540 (N_27540,N_23120,N_20840);
nand U27541 (N_27541,N_20049,N_22844);
or U27542 (N_27542,N_22775,N_20710);
and U27543 (N_27543,N_20142,N_21468);
xnor U27544 (N_27544,N_20338,N_23348);
or U27545 (N_27545,N_21936,N_23370);
xnor U27546 (N_27546,N_24841,N_24009);
and U27547 (N_27547,N_23074,N_22788);
and U27548 (N_27548,N_22601,N_22570);
xor U27549 (N_27549,N_23291,N_23908);
nand U27550 (N_27550,N_21604,N_21972);
nand U27551 (N_27551,N_23574,N_21211);
and U27552 (N_27552,N_21663,N_20506);
nand U27553 (N_27553,N_24326,N_23248);
xor U27554 (N_27554,N_21414,N_22431);
or U27555 (N_27555,N_23098,N_22752);
or U27556 (N_27556,N_20694,N_22674);
or U27557 (N_27557,N_24847,N_23049);
and U27558 (N_27558,N_23633,N_24947);
nor U27559 (N_27559,N_23678,N_20357);
nor U27560 (N_27560,N_20753,N_23384);
nand U27561 (N_27561,N_23587,N_20973);
and U27562 (N_27562,N_20380,N_22415);
nand U27563 (N_27563,N_24851,N_24507);
and U27564 (N_27564,N_22399,N_24195);
and U27565 (N_27565,N_22447,N_24527);
xnor U27566 (N_27566,N_23604,N_22183);
nor U27567 (N_27567,N_22087,N_21446);
nor U27568 (N_27568,N_24679,N_22532);
nor U27569 (N_27569,N_20184,N_24794);
or U27570 (N_27570,N_22348,N_20565);
or U27571 (N_27571,N_23148,N_22474);
or U27572 (N_27572,N_20718,N_20362);
or U27573 (N_27573,N_24448,N_22488);
nand U27574 (N_27574,N_24352,N_22118);
xor U27575 (N_27575,N_22135,N_23909);
and U27576 (N_27576,N_21023,N_24001);
xnor U27577 (N_27577,N_22610,N_22304);
and U27578 (N_27578,N_24173,N_23302);
and U27579 (N_27579,N_23587,N_24408);
and U27580 (N_27580,N_20960,N_23747);
xnor U27581 (N_27581,N_23406,N_21990);
and U27582 (N_27582,N_22185,N_20398);
xnor U27583 (N_27583,N_24863,N_23272);
or U27584 (N_27584,N_23416,N_20965);
and U27585 (N_27585,N_24681,N_21661);
or U27586 (N_27586,N_22544,N_20449);
or U27587 (N_27587,N_24565,N_20856);
nand U27588 (N_27588,N_24519,N_23859);
and U27589 (N_27589,N_20224,N_21475);
and U27590 (N_27590,N_20290,N_20508);
nand U27591 (N_27591,N_24748,N_24279);
and U27592 (N_27592,N_22644,N_24951);
nor U27593 (N_27593,N_20554,N_23544);
and U27594 (N_27594,N_22474,N_23945);
xor U27595 (N_27595,N_24406,N_22102);
and U27596 (N_27596,N_22224,N_20098);
or U27597 (N_27597,N_22471,N_21390);
or U27598 (N_27598,N_23707,N_20969);
xor U27599 (N_27599,N_21439,N_21758);
nor U27600 (N_27600,N_23585,N_20790);
nor U27601 (N_27601,N_21636,N_24351);
nor U27602 (N_27602,N_23797,N_20340);
and U27603 (N_27603,N_22933,N_21668);
xor U27604 (N_27604,N_24575,N_22439);
and U27605 (N_27605,N_20939,N_20995);
and U27606 (N_27606,N_22411,N_24498);
xor U27607 (N_27607,N_21749,N_22609);
nand U27608 (N_27608,N_20424,N_21194);
and U27609 (N_27609,N_20518,N_20618);
or U27610 (N_27610,N_20571,N_23575);
and U27611 (N_27611,N_22774,N_20329);
and U27612 (N_27612,N_21902,N_24601);
xor U27613 (N_27613,N_24193,N_21301);
xor U27614 (N_27614,N_20793,N_24512);
or U27615 (N_27615,N_21998,N_21843);
nor U27616 (N_27616,N_22351,N_23797);
or U27617 (N_27617,N_20039,N_21390);
nand U27618 (N_27618,N_21520,N_21380);
xor U27619 (N_27619,N_21700,N_20892);
nand U27620 (N_27620,N_22306,N_21125);
and U27621 (N_27621,N_23016,N_22249);
or U27622 (N_27622,N_20173,N_21546);
nor U27623 (N_27623,N_22891,N_24590);
xor U27624 (N_27624,N_20697,N_23319);
xnor U27625 (N_27625,N_21419,N_22323);
and U27626 (N_27626,N_22763,N_22628);
xor U27627 (N_27627,N_21698,N_24733);
and U27628 (N_27628,N_24609,N_22159);
or U27629 (N_27629,N_20027,N_23110);
xnor U27630 (N_27630,N_23744,N_24010);
or U27631 (N_27631,N_20029,N_22942);
and U27632 (N_27632,N_23508,N_22427);
nor U27633 (N_27633,N_22299,N_20598);
xor U27634 (N_27634,N_20436,N_24146);
and U27635 (N_27635,N_20419,N_21531);
nor U27636 (N_27636,N_21535,N_22160);
nand U27637 (N_27637,N_22335,N_21770);
xor U27638 (N_27638,N_23852,N_20851);
nor U27639 (N_27639,N_22969,N_21177);
or U27640 (N_27640,N_24838,N_20299);
nand U27641 (N_27641,N_20365,N_23938);
and U27642 (N_27642,N_21308,N_24513);
nor U27643 (N_27643,N_21379,N_20649);
and U27644 (N_27644,N_23614,N_22309);
nor U27645 (N_27645,N_21747,N_22039);
nand U27646 (N_27646,N_24199,N_23956);
and U27647 (N_27647,N_22777,N_23761);
or U27648 (N_27648,N_24333,N_22617);
and U27649 (N_27649,N_20943,N_23309);
nand U27650 (N_27650,N_22076,N_22614);
nor U27651 (N_27651,N_23609,N_24882);
nor U27652 (N_27652,N_22007,N_24777);
nand U27653 (N_27653,N_23710,N_21060);
or U27654 (N_27654,N_22315,N_24833);
xnor U27655 (N_27655,N_20381,N_21878);
xor U27656 (N_27656,N_21850,N_22258);
or U27657 (N_27657,N_23115,N_22358);
and U27658 (N_27658,N_20001,N_20428);
nor U27659 (N_27659,N_21514,N_20150);
or U27660 (N_27660,N_24318,N_24370);
or U27661 (N_27661,N_20488,N_22478);
xor U27662 (N_27662,N_20855,N_21288);
or U27663 (N_27663,N_23059,N_22841);
nor U27664 (N_27664,N_21378,N_22305);
or U27665 (N_27665,N_24572,N_24502);
nand U27666 (N_27666,N_22750,N_21156);
nor U27667 (N_27667,N_23143,N_22353);
nor U27668 (N_27668,N_24455,N_24720);
nor U27669 (N_27669,N_22775,N_24451);
and U27670 (N_27670,N_23351,N_20370);
nor U27671 (N_27671,N_20703,N_21779);
nor U27672 (N_27672,N_23541,N_20354);
xnor U27673 (N_27673,N_21281,N_20776);
xnor U27674 (N_27674,N_24156,N_21069);
nor U27675 (N_27675,N_22727,N_23430);
nor U27676 (N_27676,N_21533,N_23752);
nor U27677 (N_27677,N_20366,N_22994);
and U27678 (N_27678,N_24770,N_23620);
or U27679 (N_27679,N_21309,N_21344);
and U27680 (N_27680,N_20424,N_20544);
or U27681 (N_27681,N_23326,N_22151);
and U27682 (N_27682,N_24456,N_21163);
xor U27683 (N_27683,N_23552,N_22341);
nand U27684 (N_27684,N_20733,N_23864);
nor U27685 (N_27685,N_23831,N_24913);
nor U27686 (N_27686,N_21482,N_24522);
and U27687 (N_27687,N_22993,N_20700);
nand U27688 (N_27688,N_24735,N_23027);
and U27689 (N_27689,N_20429,N_23583);
nand U27690 (N_27690,N_21024,N_24388);
xnor U27691 (N_27691,N_21315,N_24455);
or U27692 (N_27692,N_24105,N_23636);
and U27693 (N_27693,N_20505,N_20775);
and U27694 (N_27694,N_22963,N_24538);
xor U27695 (N_27695,N_21835,N_22298);
nor U27696 (N_27696,N_20124,N_24604);
nor U27697 (N_27697,N_22279,N_22057);
or U27698 (N_27698,N_20376,N_23060);
or U27699 (N_27699,N_23442,N_24370);
and U27700 (N_27700,N_20248,N_23823);
nand U27701 (N_27701,N_22332,N_23493);
nand U27702 (N_27702,N_20853,N_24497);
or U27703 (N_27703,N_20518,N_22606);
nand U27704 (N_27704,N_24029,N_21279);
and U27705 (N_27705,N_20289,N_21395);
xor U27706 (N_27706,N_20813,N_20635);
nor U27707 (N_27707,N_21646,N_24723);
nand U27708 (N_27708,N_22428,N_24428);
nor U27709 (N_27709,N_21484,N_21287);
and U27710 (N_27710,N_23993,N_22801);
xnor U27711 (N_27711,N_22448,N_24161);
or U27712 (N_27712,N_23157,N_21452);
or U27713 (N_27713,N_23111,N_23369);
nor U27714 (N_27714,N_21753,N_21012);
nand U27715 (N_27715,N_20277,N_21609);
xor U27716 (N_27716,N_24901,N_23040);
xnor U27717 (N_27717,N_20669,N_22682);
or U27718 (N_27718,N_21696,N_20878);
nand U27719 (N_27719,N_22693,N_23106);
and U27720 (N_27720,N_23850,N_23581);
nor U27721 (N_27721,N_24754,N_23057);
nor U27722 (N_27722,N_22360,N_21243);
nor U27723 (N_27723,N_21538,N_20127);
nor U27724 (N_27724,N_23663,N_22787);
xnor U27725 (N_27725,N_24943,N_21813);
or U27726 (N_27726,N_22670,N_21106);
and U27727 (N_27727,N_23952,N_21862);
nor U27728 (N_27728,N_22547,N_21993);
nor U27729 (N_27729,N_24296,N_22752);
nand U27730 (N_27730,N_24175,N_24362);
xor U27731 (N_27731,N_20746,N_24219);
nor U27732 (N_27732,N_22066,N_20211);
or U27733 (N_27733,N_22531,N_22330);
or U27734 (N_27734,N_21051,N_24306);
and U27735 (N_27735,N_21446,N_21473);
and U27736 (N_27736,N_22437,N_24615);
xnor U27737 (N_27737,N_21260,N_20037);
nand U27738 (N_27738,N_22125,N_24842);
nand U27739 (N_27739,N_20182,N_22950);
nand U27740 (N_27740,N_22856,N_24866);
and U27741 (N_27741,N_22903,N_24456);
nor U27742 (N_27742,N_21410,N_22641);
nor U27743 (N_27743,N_24270,N_23955);
or U27744 (N_27744,N_20037,N_23513);
nor U27745 (N_27745,N_22350,N_20210);
nand U27746 (N_27746,N_22151,N_22995);
nand U27747 (N_27747,N_21442,N_24015);
xnor U27748 (N_27748,N_20946,N_20325);
xor U27749 (N_27749,N_20265,N_22278);
or U27750 (N_27750,N_20089,N_23813);
xor U27751 (N_27751,N_21219,N_20900);
and U27752 (N_27752,N_23805,N_23813);
nor U27753 (N_27753,N_20269,N_21441);
or U27754 (N_27754,N_24762,N_24823);
nor U27755 (N_27755,N_22450,N_21334);
and U27756 (N_27756,N_24087,N_21680);
and U27757 (N_27757,N_23336,N_24046);
and U27758 (N_27758,N_20663,N_24100);
xor U27759 (N_27759,N_21086,N_23500);
and U27760 (N_27760,N_20538,N_23854);
or U27761 (N_27761,N_21205,N_20326);
xnor U27762 (N_27762,N_24583,N_22918);
nand U27763 (N_27763,N_21481,N_22426);
nand U27764 (N_27764,N_24499,N_20400);
and U27765 (N_27765,N_22239,N_22905);
or U27766 (N_27766,N_22626,N_20813);
xor U27767 (N_27767,N_23364,N_22197);
nor U27768 (N_27768,N_20672,N_20537);
nor U27769 (N_27769,N_23420,N_20696);
nor U27770 (N_27770,N_24082,N_24474);
or U27771 (N_27771,N_20292,N_21842);
nor U27772 (N_27772,N_24434,N_21669);
or U27773 (N_27773,N_23641,N_21798);
xor U27774 (N_27774,N_24706,N_21817);
or U27775 (N_27775,N_21237,N_20899);
or U27776 (N_27776,N_21152,N_20290);
nand U27777 (N_27777,N_20309,N_24845);
nor U27778 (N_27778,N_22829,N_21581);
nand U27779 (N_27779,N_20187,N_24288);
xnor U27780 (N_27780,N_20704,N_21143);
xnor U27781 (N_27781,N_22427,N_20391);
and U27782 (N_27782,N_22331,N_20400);
or U27783 (N_27783,N_22105,N_22233);
nor U27784 (N_27784,N_22736,N_20612);
and U27785 (N_27785,N_23166,N_22728);
nand U27786 (N_27786,N_23026,N_21159);
nor U27787 (N_27787,N_21380,N_24691);
nand U27788 (N_27788,N_22934,N_23287);
xor U27789 (N_27789,N_20710,N_21070);
nand U27790 (N_27790,N_24635,N_22462);
nand U27791 (N_27791,N_24178,N_24409);
and U27792 (N_27792,N_20431,N_21622);
xnor U27793 (N_27793,N_24307,N_21244);
nor U27794 (N_27794,N_23837,N_20382);
or U27795 (N_27795,N_20210,N_24575);
xor U27796 (N_27796,N_24379,N_23984);
or U27797 (N_27797,N_21766,N_22143);
and U27798 (N_27798,N_22857,N_21207);
nor U27799 (N_27799,N_22131,N_22469);
and U27800 (N_27800,N_21042,N_23014);
and U27801 (N_27801,N_23303,N_21270);
or U27802 (N_27802,N_20847,N_20819);
and U27803 (N_27803,N_24331,N_20871);
xnor U27804 (N_27804,N_23493,N_20864);
and U27805 (N_27805,N_20845,N_23078);
xnor U27806 (N_27806,N_23985,N_23023);
nor U27807 (N_27807,N_21164,N_23877);
or U27808 (N_27808,N_24087,N_21794);
nand U27809 (N_27809,N_24495,N_23059);
and U27810 (N_27810,N_21872,N_22750);
xnor U27811 (N_27811,N_23789,N_24341);
and U27812 (N_27812,N_20325,N_22331);
or U27813 (N_27813,N_21694,N_22971);
or U27814 (N_27814,N_23058,N_24099);
xor U27815 (N_27815,N_22831,N_20687);
xnor U27816 (N_27816,N_20905,N_23645);
nand U27817 (N_27817,N_22472,N_20465);
nor U27818 (N_27818,N_22067,N_21461);
xnor U27819 (N_27819,N_21859,N_21073);
and U27820 (N_27820,N_23345,N_20037);
nand U27821 (N_27821,N_20623,N_24838);
nand U27822 (N_27822,N_23340,N_22582);
nand U27823 (N_27823,N_23759,N_21801);
or U27824 (N_27824,N_24773,N_20024);
xnor U27825 (N_27825,N_21819,N_23149);
xor U27826 (N_27826,N_23062,N_22598);
or U27827 (N_27827,N_21788,N_21490);
or U27828 (N_27828,N_22257,N_20412);
xnor U27829 (N_27829,N_21469,N_21966);
xor U27830 (N_27830,N_21278,N_21879);
nand U27831 (N_27831,N_23604,N_20181);
nand U27832 (N_27832,N_20278,N_24386);
and U27833 (N_27833,N_23572,N_20388);
nand U27834 (N_27834,N_23606,N_22396);
xor U27835 (N_27835,N_21314,N_24283);
nand U27836 (N_27836,N_20463,N_20112);
nand U27837 (N_27837,N_22737,N_21798);
nor U27838 (N_27838,N_22799,N_21031);
nand U27839 (N_27839,N_23769,N_21761);
xnor U27840 (N_27840,N_21785,N_24563);
xnor U27841 (N_27841,N_24791,N_20012);
nor U27842 (N_27842,N_21113,N_24778);
xor U27843 (N_27843,N_21265,N_21235);
nor U27844 (N_27844,N_22140,N_24434);
and U27845 (N_27845,N_21670,N_20712);
nor U27846 (N_27846,N_23058,N_24773);
and U27847 (N_27847,N_24882,N_21020);
or U27848 (N_27848,N_21183,N_20547);
and U27849 (N_27849,N_23903,N_20514);
and U27850 (N_27850,N_24158,N_22816);
nand U27851 (N_27851,N_21711,N_22505);
or U27852 (N_27852,N_21451,N_20282);
xnor U27853 (N_27853,N_24242,N_20011);
and U27854 (N_27854,N_23086,N_22750);
xor U27855 (N_27855,N_24078,N_20304);
and U27856 (N_27856,N_22346,N_23501);
xor U27857 (N_27857,N_24891,N_20860);
nor U27858 (N_27858,N_24002,N_24940);
xor U27859 (N_27859,N_24438,N_22961);
xor U27860 (N_27860,N_21983,N_23476);
nor U27861 (N_27861,N_23395,N_22329);
nor U27862 (N_27862,N_23347,N_21118);
xor U27863 (N_27863,N_21186,N_21602);
and U27864 (N_27864,N_21802,N_21614);
and U27865 (N_27865,N_20804,N_20193);
nand U27866 (N_27866,N_21272,N_24927);
and U27867 (N_27867,N_22131,N_20272);
xor U27868 (N_27868,N_22483,N_23524);
or U27869 (N_27869,N_21640,N_24213);
and U27870 (N_27870,N_23328,N_22645);
nor U27871 (N_27871,N_22547,N_20477);
or U27872 (N_27872,N_21782,N_20696);
and U27873 (N_27873,N_23295,N_23296);
and U27874 (N_27874,N_24192,N_21903);
nand U27875 (N_27875,N_21077,N_24933);
xor U27876 (N_27876,N_22990,N_23261);
nor U27877 (N_27877,N_22084,N_22247);
nand U27878 (N_27878,N_21959,N_22061);
nor U27879 (N_27879,N_22484,N_24707);
xor U27880 (N_27880,N_20891,N_23966);
nand U27881 (N_27881,N_21480,N_24258);
or U27882 (N_27882,N_24699,N_22204);
or U27883 (N_27883,N_21785,N_24599);
or U27884 (N_27884,N_20483,N_22853);
xnor U27885 (N_27885,N_21579,N_20661);
or U27886 (N_27886,N_20378,N_24580);
xnor U27887 (N_27887,N_21067,N_21503);
nand U27888 (N_27888,N_24830,N_23602);
xnor U27889 (N_27889,N_23685,N_20020);
nand U27890 (N_27890,N_24855,N_20156);
and U27891 (N_27891,N_24132,N_21279);
and U27892 (N_27892,N_20776,N_20421);
nand U27893 (N_27893,N_20508,N_22980);
xor U27894 (N_27894,N_22651,N_20302);
and U27895 (N_27895,N_20205,N_20426);
and U27896 (N_27896,N_24183,N_22930);
xor U27897 (N_27897,N_21130,N_21572);
nand U27898 (N_27898,N_23948,N_24157);
xnor U27899 (N_27899,N_20181,N_22742);
nand U27900 (N_27900,N_24415,N_20383);
nand U27901 (N_27901,N_24267,N_20989);
nor U27902 (N_27902,N_24154,N_20537);
or U27903 (N_27903,N_22510,N_20696);
xor U27904 (N_27904,N_24870,N_23290);
nand U27905 (N_27905,N_24891,N_22237);
nor U27906 (N_27906,N_22441,N_20639);
and U27907 (N_27907,N_21960,N_21239);
nor U27908 (N_27908,N_23992,N_23559);
nor U27909 (N_27909,N_24543,N_20035);
and U27910 (N_27910,N_20107,N_24564);
nor U27911 (N_27911,N_20410,N_23401);
or U27912 (N_27912,N_20403,N_20446);
nand U27913 (N_27913,N_22251,N_24160);
and U27914 (N_27914,N_20115,N_22441);
xor U27915 (N_27915,N_22405,N_23798);
nor U27916 (N_27916,N_22205,N_22614);
and U27917 (N_27917,N_24640,N_21524);
nand U27918 (N_27918,N_20588,N_23822);
nand U27919 (N_27919,N_23910,N_21938);
nor U27920 (N_27920,N_23081,N_24228);
nor U27921 (N_27921,N_20199,N_20160);
nand U27922 (N_27922,N_21605,N_21647);
and U27923 (N_27923,N_24287,N_20277);
or U27924 (N_27924,N_20576,N_22662);
nand U27925 (N_27925,N_21473,N_24142);
or U27926 (N_27926,N_22055,N_20560);
and U27927 (N_27927,N_20333,N_22390);
nor U27928 (N_27928,N_24906,N_24314);
nor U27929 (N_27929,N_20260,N_22975);
and U27930 (N_27930,N_21172,N_20666);
nand U27931 (N_27931,N_22772,N_24578);
xor U27932 (N_27932,N_24452,N_24640);
and U27933 (N_27933,N_24289,N_20346);
or U27934 (N_27934,N_22776,N_24504);
or U27935 (N_27935,N_21207,N_23067);
xor U27936 (N_27936,N_23371,N_21707);
nand U27937 (N_27937,N_23961,N_24190);
or U27938 (N_27938,N_21013,N_21514);
and U27939 (N_27939,N_22423,N_20912);
or U27940 (N_27940,N_22337,N_22751);
nand U27941 (N_27941,N_20749,N_22842);
xnor U27942 (N_27942,N_21927,N_21141);
nand U27943 (N_27943,N_23536,N_24458);
or U27944 (N_27944,N_23765,N_21338);
and U27945 (N_27945,N_24147,N_20963);
and U27946 (N_27946,N_22508,N_22494);
nand U27947 (N_27947,N_23004,N_20854);
or U27948 (N_27948,N_22012,N_24188);
nand U27949 (N_27949,N_21584,N_21891);
nand U27950 (N_27950,N_21365,N_21092);
or U27951 (N_27951,N_22370,N_22054);
and U27952 (N_27952,N_24626,N_22477);
and U27953 (N_27953,N_21844,N_20084);
nand U27954 (N_27954,N_21997,N_20903);
nor U27955 (N_27955,N_23771,N_20040);
or U27956 (N_27956,N_21543,N_20152);
or U27957 (N_27957,N_22009,N_23602);
xor U27958 (N_27958,N_20120,N_24874);
nand U27959 (N_27959,N_22596,N_23998);
xnor U27960 (N_27960,N_23795,N_21548);
or U27961 (N_27961,N_23613,N_24372);
and U27962 (N_27962,N_22196,N_22283);
or U27963 (N_27963,N_21748,N_24495);
xnor U27964 (N_27964,N_23855,N_23599);
nand U27965 (N_27965,N_22816,N_24083);
nor U27966 (N_27966,N_21436,N_21968);
nor U27967 (N_27967,N_21340,N_24637);
and U27968 (N_27968,N_23428,N_24827);
and U27969 (N_27969,N_22744,N_23634);
nor U27970 (N_27970,N_24065,N_24192);
and U27971 (N_27971,N_24602,N_22207);
and U27972 (N_27972,N_22765,N_22386);
and U27973 (N_27973,N_20275,N_21228);
nor U27974 (N_27974,N_20517,N_20575);
or U27975 (N_27975,N_24119,N_20319);
xnor U27976 (N_27976,N_21404,N_22987);
nand U27977 (N_27977,N_21010,N_23260);
nor U27978 (N_27978,N_20368,N_23070);
nand U27979 (N_27979,N_20487,N_22548);
or U27980 (N_27980,N_23084,N_21496);
xnor U27981 (N_27981,N_22156,N_21491);
xor U27982 (N_27982,N_21275,N_21614);
or U27983 (N_27983,N_22478,N_21333);
nand U27984 (N_27984,N_21822,N_23116);
nor U27985 (N_27985,N_20915,N_24277);
xor U27986 (N_27986,N_21947,N_23722);
and U27987 (N_27987,N_23247,N_23550);
nand U27988 (N_27988,N_24833,N_20328);
nand U27989 (N_27989,N_22675,N_21639);
nand U27990 (N_27990,N_23521,N_20950);
or U27991 (N_27991,N_20520,N_20749);
nor U27992 (N_27992,N_24166,N_24079);
nand U27993 (N_27993,N_22856,N_21547);
and U27994 (N_27994,N_21355,N_20167);
or U27995 (N_27995,N_23310,N_23629);
nor U27996 (N_27996,N_22820,N_22213);
and U27997 (N_27997,N_21864,N_23629);
and U27998 (N_27998,N_20599,N_20946);
and U27999 (N_27999,N_21834,N_20252);
xor U28000 (N_28000,N_24285,N_22647);
nor U28001 (N_28001,N_21455,N_21597);
xor U28002 (N_28002,N_20193,N_21284);
or U28003 (N_28003,N_22192,N_22740);
xnor U28004 (N_28004,N_24515,N_24745);
or U28005 (N_28005,N_22236,N_20803);
nor U28006 (N_28006,N_21844,N_21448);
and U28007 (N_28007,N_20695,N_23023);
and U28008 (N_28008,N_22927,N_21380);
xor U28009 (N_28009,N_23329,N_22787);
nand U28010 (N_28010,N_23407,N_23011);
xnor U28011 (N_28011,N_20034,N_24520);
or U28012 (N_28012,N_21680,N_23504);
xor U28013 (N_28013,N_20689,N_23087);
or U28014 (N_28014,N_23883,N_20838);
nand U28015 (N_28015,N_23894,N_20311);
and U28016 (N_28016,N_24900,N_21229);
nand U28017 (N_28017,N_23045,N_22750);
nor U28018 (N_28018,N_20289,N_24796);
and U28019 (N_28019,N_23259,N_24874);
or U28020 (N_28020,N_21959,N_21660);
nand U28021 (N_28021,N_22052,N_20498);
nand U28022 (N_28022,N_24788,N_24442);
nor U28023 (N_28023,N_24144,N_23646);
nor U28024 (N_28024,N_22589,N_23378);
xnor U28025 (N_28025,N_24075,N_20144);
xnor U28026 (N_28026,N_20572,N_21213);
nor U28027 (N_28027,N_24070,N_21918);
nand U28028 (N_28028,N_20443,N_20841);
and U28029 (N_28029,N_24944,N_24041);
xnor U28030 (N_28030,N_22907,N_22312);
and U28031 (N_28031,N_22772,N_22020);
nand U28032 (N_28032,N_24753,N_21429);
nand U28033 (N_28033,N_24578,N_21747);
nand U28034 (N_28034,N_24651,N_20115);
and U28035 (N_28035,N_23310,N_24892);
nand U28036 (N_28036,N_23883,N_24269);
nand U28037 (N_28037,N_20649,N_20217);
nand U28038 (N_28038,N_23829,N_20692);
xor U28039 (N_28039,N_22338,N_21405);
or U28040 (N_28040,N_24199,N_23883);
nand U28041 (N_28041,N_24651,N_24335);
nor U28042 (N_28042,N_21012,N_21405);
nand U28043 (N_28043,N_23831,N_23083);
xor U28044 (N_28044,N_22551,N_21184);
or U28045 (N_28045,N_21360,N_22739);
nand U28046 (N_28046,N_24357,N_20248);
xor U28047 (N_28047,N_24139,N_22270);
xnor U28048 (N_28048,N_23254,N_22150);
nand U28049 (N_28049,N_24036,N_20286);
xnor U28050 (N_28050,N_23045,N_20796);
and U28051 (N_28051,N_24414,N_21786);
nor U28052 (N_28052,N_24207,N_22804);
or U28053 (N_28053,N_21314,N_23670);
nor U28054 (N_28054,N_24507,N_21089);
nand U28055 (N_28055,N_22209,N_23214);
or U28056 (N_28056,N_21041,N_23234);
nand U28057 (N_28057,N_23285,N_20052);
nand U28058 (N_28058,N_21100,N_23876);
nand U28059 (N_28059,N_21657,N_23144);
xnor U28060 (N_28060,N_24754,N_23879);
xnor U28061 (N_28061,N_22133,N_23553);
nor U28062 (N_28062,N_21209,N_21804);
and U28063 (N_28063,N_24057,N_23159);
nor U28064 (N_28064,N_23165,N_23497);
and U28065 (N_28065,N_24979,N_22419);
or U28066 (N_28066,N_20136,N_22787);
and U28067 (N_28067,N_23250,N_21360);
or U28068 (N_28068,N_22375,N_23902);
nand U28069 (N_28069,N_24964,N_21634);
and U28070 (N_28070,N_20325,N_21345);
or U28071 (N_28071,N_21353,N_24521);
or U28072 (N_28072,N_22465,N_24989);
nor U28073 (N_28073,N_21966,N_22063);
nor U28074 (N_28074,N_20830,N_21085);
or U28075 (N_28075,N_23855,N_23409);
and U28076 (N_28076,N_24291,N_22972);
nand U28077 (N_28077,N_21458,N_21151);
nand U28078 (N_28078,N_21665,N_20779);
nor U28079 (N_28079,N_23147,N_20085);
or U28080 (N_28080,N_20363,N_21096);
or U28081 (N_28081,N_24626,N_23463);
nor U28082 (N_28082,N_20090,N_21719);
or U28083 (N_28083,N_20833,N_22880);
nor U28084 (N_28084,N_22607,N_22938);
nor U28085 (N_28085,N_23371,N_22364);
and U28086 (N_28086,N_21428,N_24135);
and U28087 (N_28087,N_24586,N_22898);
nor U28088 (N_28088,N_24576,N_22690);
nor U28089 (N_28089,N_23755,N_24502);
nand U28090 (N_28090,N_20909,N_24140);
xor U28091 (N_28091,N_21856,N_24062);
xnor U28092 (N_28092,N_23180,N_20589);
and U28093 (N_28093,N_21973,N_22481);
nor U28094 (N_28094,N_20605,N_23331);
nand U28095 (N_28095,N_23488,N_22511);
and U28096 (N_28096,N_22136,N_21067);
nor U28097 (N_28097,N_24834,N_21620);
nor U28098 (N_28098,N_22883,N_23733);
nand U28099 (N_28099,N_20630,N_22668);
xor U28100 (N_28100,N_20283,N_22941);
xnor U28101 (N_28101,N_21175,N_20224);
and U28102 (N_28102,N_22370,N_21704);
xnor U28103 (N_28103,N_20667,N_23653);
and U28104 (N_28104,N_21505,N_23000);
nor U28105 (N_28105,N_23440,N_21216);
nand U28106 (N_28106,N_20375,N_24625);
xor U28107 (N_28107,N_23672,N_24319);
nor U28108 (N_28108,N_21520,N_20000);
and U28109 (N_28109,N_22235,N_23600);
nand U28110 (N_28110,N_22409,N_20859);
and U28111 (N_28111,N_24519,N_22924);
nand U28112 (N_28112,N_23160,N_22294);
and U28113 (N_28113,N_24373,N_21212);
xnor U28114 (N_28114,N_22673,N_24425);
and U28115 (N_28115,N_22661,N_20549);
nor U28116 (N_28116,N_24619,N_23449);
or U28117 (N_28117,N_21432,N_22916);
or U28118 (N_28118,N_20082,N_20559);
xnor U28119 (N_28119,N_23680,N_23242);
xnor U28120 (N_28120,N_23848,N_24926);
xor U28121 (N_28121,N_24420,N_23071);
nand U28122 (N_28122,N_20497,N_21424);
xor U28123 (N_28123,N_23457,N_24611);
nand U28124 (N_28124,N_22855,N_20449);
and U28125 (N_28125,N_23646,N_20880);
nand U28126 (N_28126,N_21633,N_21241);
or U28127 (N_28127,N_24260,N_24911);
nand U28128 (N_28128,N_24657,N_24890);
xnor U28129 (N_28129,N_24245,N_23605);
or U28130 (N_28130,N_22813,N_20888);
nor U28131 (N_28131,N_23990,N_20602);
xnor U28132 (N_28132,N_24268,N_22493);
xnor U28133 (N_28133,N_24045,N_23317);
or U28134 (N_28134,N_21143,N_21985);
and U28135 (N_28135,N_20944,N_21301);
or U28136 (N_28136,N_23923,N_22243);
or U28137 (N_28137,N_22248,N_21835);
and U28138 (N_28138,N_23317,N_24914);
nand U28139 (N_28139,N_22259,N_22868);
or U28140 (N_28140,N_20464,N_21573);
nand U28141 (N_28141,N_22408,N_23769);
and U28142 (N_28142,N_24331,N_20000);
nor U28143 (N_28143,N_23201,N_20008);
nor U28144 (N_28144,N_20741,N_21190);
nand U28145 (N_28145,N_20056,N_24903);
nand U28146 (N_28146,N_20650,N_21708);
nor U28147 (N_28147,N_20088,N_21064);
or U28148 (N_28148,N_23419,N_23845);
nand U28149 (N_28149,N_24599,N_20011);
and U28150 (N_28150,N_20535,N_20576);
xor U28151 (N_28151,N_20087,N_21521);
nand U28152 (N_28152,N_20728,N_23605);
xnor U28153 (N_28153,N_20444,N_24770);
xnor U28154 (N_28154,N_21495,N_21157);
xor U28155 (N_28155,N_20389,N_21306);
xnor U28156 (N_28156,N_21389,N_20912);
or U28157 (N_28157,N_24701,N_21454);
or U28158 (N_28158,N_20652,N_22068);
nand U28159 (N_28159,N_24476,N_22776);
nor U28160 (N_28160,N_20167,N_20813);
and U28161 (N_28161,N_23083,N_22579);
nor U28162 (N_28162,N_21525,N_21565);
xor U28163 (N_28163,N_23788,N_23288);
and U28164 (N_28164,N_20946,N_23944);
nand U28165 (N_28165,N_24877,N_20230);
or U28166 (N_28166,N_23095,N_23222);
and U28167 (N_28167,N_23733,N_21138);
nand U28168 (N_28168,N_22890,N_22143);
nor U28169 (N_28169,N_22705,N_22134);
and U28170 (N_28170,N_20131,N_23908);
xnor U28171 (N_28171,N_23001,N_24132);
nor U28172 (N_28172,N_20175,N_22970);
or U28173 (N_28173,N_24840,N_21065);
xor U28174 (N_28174,N_22577,N_22587);
nor U28175 (N_28175,N_20805,N_22073);
and U28176 (N_28176,N_23736,N_21029);
xnor U28177 (N_28177,N_24108,N_20953);
nand U28178 (N_28178,N_23233,N_24226);
or U28179 (N_28179,N_20999,N_24101);
or U28180 (N_28180,N_24052,N_21484);
and U28181 (N_28181,N_24854,N_21067);
and U28182 (N_28182,N_24819,N_20957);
nand U28183 (N_28183,N_23748,N_24560);
and U28184 (N_28184,N_24295,N_23240);
nor U28185 (N_28185,N_21229,N_24204);
nand U28186 (N_28186,N_24592,N_24319);
or U28187 (N_28187,N_23770,N_23968);
xor U28188 (N_28188,N_20984,N_21746);
or U28189 (N_28189,N_20458,N_22700);
xnor U28190 (N_28190,N_22831,N_24814);
nand U28191 (N_28191,N_23497,N_24164);
nor U28192 (N_28192,N_20777,N_21948);
and U28193 (N_28193,N_20304,N_21298);
nor U28194 (N_28194,N_20461,N_24692);
xnor U28195 (N_28195,N_23424,N_21748);
nand U28196 (N_28196,N_20702,N_23940);
xnor U28197 (N_28197,N_24605,N_21694);
nor U28198 (N_28198,N_24467,N_24169);
or U28199 (N_28199,N_23418,N_22496);
or U28200 (N_28200,N_24780,N_22483);
or U28201 (N_28201,N_20270,N_23553);
xnor U28202 (N_28202,N_24817,N_20480);
xor U28203 (N_28203,N_21570,N_24174);
or U28204 (N_28204,N_21340,N_22255);
nor U28205 (N_28205,N_20337,N_24556);
xor U28206 (N_28206,N_20389,N_24196);
xnor U28207 (N_28207,N_22220,N_24014);
nor U28208 (N_28208,N_22964,N_24992);
xnor U28209 (N_28209,N_24572,N_20344);
nor U28210 (N_28210,N_20492,N_23107);
nor U28211 (N_28211,N_21612,N_21100);
nor U28212 (N_28212,N_24270,N_21345);
xnor U28213 (N_28213,N_21011,N_20830);
nand U28214 (N_28214,N_23200,N_23652);
xnor U28215 (N_28215,N_22434,N_23636);
nor U28216 (N_28216,N_24454,N_22011);
nand U28217 (N_28217,N_20394,N_20987);
nand U28218 (N_28218,N_21825,N_20847);
nor U28219 (N_28219,N_21224,N_21856);
or U28220 (N_28220,N_20225,N_23366);
nand U28221 (N_28221,N_23646,N_22549);
or U28222 (N_28222,N_20951,N_24304);
nor U28223 (N_28223,N_24467,N_23373);
and U28224 (N_28224,N_22471,N_24425);
xor U28225 (N_28225,N_23275,N_23005);
or U28226 (N_28226,N_22115,N_23474);
or U28227 (N_28227,N_20071,N_23904);
xor U28228 (N_28228,N_22335,N_24419);
and U28229 (N_28229,N_22607,N_21475);
nor U28230 (N_28230,N_21840,N_23216);
or U28231 (N_28231,N_22400,N_21133);
or U28232 (N_28232,N_21560,N_24419);
nor U28233 (N_28233,N_23942,N_20792);
xor U28234 (N_28234,N_23354,N_23664);
nor U28235 (N_28235,N_20793,N_22243);
nand U28236 (N_28236,N_20602,N_22588);
nand U28237 (N_28237,N_21549,N_20718);
or U28238 (N_28238,N_20235,N_21669);
or U28239 (N_28239,N_21196,N_24526);
or U28240 (N_28240,N_23164,N_23561);
nand U28241 (N_28241,N_24785,N_21630);
nor U28242 (N_28242,N_23209,N_24652);
nor U28243 (N_28243,N_22127,N_21075);
nand U28244 (N_28244,N_24137,N_20701);
nor U28245 (N_28245,N_21609,N_20077);
xnor U28246 (N_28246,N_22007,N_21944);
xor U28247 (N_28247,N_22581,N_20496);
or U28248 (N_28248,N_22170,N_24563);
nor U28249 (N_28249,N_23667,N_20755);
nor U28250 (N_28250,N_22376,N_24242);
and U28251 (N_28251,N_21502,N_23438);
nand U28252 (N_28252,N_20146,N_24219);
nor U28253 (N_28253,N_21396,N_20394);
and U28254 (N_28254,N_24767,N_21583);
xor U28255 (N_28255,N_23643,N_24459);
nor U28256 (N_28256,N_22017,N_23426);
or U28257 (N_28257,N_23882,N_23704);
and U28258 (N_28258,N_22262,N_23813);
or U28259 (N_28259,N_24105,N_20361);
xnor U28260 (N_28260,N_23657,N_22480);
and U28261 (N_28261,N_22339,N_21498);
nor U28262 (N_28262,N_23507,N_21152);
xnor U28263 (N_28263,N_22654,N_24325);
nand U28264 (N_28264,N_21312,N_23478);
xnor U28265 (N_28265,N_20113,N_22739);
or U28266 (N_28266,N_21712,N_20676);
nor U28267 (N_28267,N_21341,N_22372);
or U28268 (N_28268,N_22761,N_24955);
nand U28269 (N_28269,N_23520,N_24550);
nor U28270 (N_28270,N_20942,N_24450);
xnor U28271 (N_28271,N_24382,N_24264);
nor U28272 (N_28272,N_24536,N_23756);
xnor U28273 (N_28273,N_24425,N_23837);
or U28274 (N_28274,N_22037,N_23439);
nor U28275 (N_28275,N_23683,N_22869);
and U28276 (N_28276,N_23507,N_21261);
nor U28277 (N_28277,N_24470,N_21693);
and U28278 (N_28278,N_24856,N_20981);
or U28279 (N_28279,N_23793,N_24745);
nand U28280 (N_28280,N_23993,N_23713);
and U28281 (N_28281,N_21491,N_22483);
and U28282 (N_28282,N_20164,N_23359);
nor U28283 (N_28283,N_23610,N_22429);
nor U28284 (N_28284,N_20197,N_24322);
xor U28285 (N_28285,N_21905,N_22857);
nand U28286 (N_28286,N_20284,N_22344);
or U28287 (N_28287,N_22710,N_23387);
xor U28288 (N_28288,N_23773,N_22442);
and U28289 (N_28289,N_20654,N_20680);
and U28290 (N_28290,N_22793,N_23839);
nor U28291 (N_28291,N_20481,N_22253);
nor U28292 (N_28292,N_23000,N_20407);
xnor U28293 (N_28293,N_22121,N_21136);
and U28294 (N_28294,N_20966,N_22309);
and U28295 (N_28295,N_22287,N_21900);
nor U28296 (N_28296,N_23230,N_23938);
xor U28297 (N_28297,N_20645,N_24127);
nor U28298 (N_28298,N_22173,N_24778);
and U28299 (N_28299,N_23037,N_24390);
xor U28300 (N_28300,N_23784,N_20976);
nand U28301 (N_28301,N_23853,N_20763);
nor U28302 (N_28302,N_24460,N_23793);
and U28303 (N_28303,N_20376,N_22791);
xor U28304 (N_28304,N_20707,N_23689);
nand U28305 (N_28305,N_21722,N_22504);
or U28306 (N_28306,N_22212,N_22456);
and U28307 (N_28307,N_23777,N_21468);
nand U28308 (N_28308,N_20274,N_20703);
or U28309 (N_28309,N_20476,N_24754);
xor U28310 (N_28310,N_22036,N_23405);
or U28311 (N_28311,N_21217,N_21015);
nand U28312 (N_28312,N_21475,N_23721);
nand U28313 (N_28313,N_24130,N_21067);
nor U28314 (N_28314,N_24106,N_24275);
nand U28315 (N_28315,N_21762,N_23712);
and U28316 (N_28316,N_24395,N_24619);
xnor U28317 (N_28317,N_23768,N_20633);
and U28318 (N_28318,N_24760,N_24381);
and U28319 (N_28319,N_23728,N_20060);
nand U28320 (N_28320,N_20838,N_24416);
nor U28321 (N_28321,N_21358,N_20401);
or U28322 (N_28322,N_20434,N_22606);
xnor U28323 (N_28323,N_24229,N_20824);
or U28324 (N_28324,N_21366,N_20454);
and U28325 (N_28325,N_22122,N_21739);
and U28326 (N_28326,N_22823,N_23259);
nand U28327 (N_28327,N_20631,N_22096);
nor U28328 (N_28328,N_20312,N_23071);
nor U28329 (N_28329,N_23947,N_20343);
nor U28330 (N_28330,N_20880,N_20567);
and U28331 (N_28331,N_23966,N_24543);
xor U28332 (N_28332,N_20789,N_22021);
and U28333 (N_28333,N_24489,N_21633);
nand U28334 (N_28334,N_21698,N_20326);
nor U28335 (N_28335,N_22548,N_23694);
nor U28336 (N_28336,N_21168,N_20700);
xor U28337 (N_28337,N_23646,N_23418);
nand U28338 (N_28338,N_24919,N_24809);
or U28339 (N_28339,N_20713,N_22026);
nor U28340 (N_28340,N_24324,N_24660);
or U28341 (N_28341,N_24170,N_21705);
nand U28342 (N_28342,N_20953,N_21479);
and U28343 (N_28343,N_24862,N_20040);
nand U28344 (N_28344,N_23693,N_23316);
nand U28345 (N_28345,N_23621,N_21001);
and U28346 (N_28346,N_24807,N_23645);
or U28347 (N_28347,N_23915,N_22360);
and U28348 (N_28348,N_21015,N_21322);
nand U28349 (N_28349,N_23102,N_21882);
nand U28350 (N_28350,N_21806,N_24035);
nor U28351 (N_28351,N_22807,N_24877);
nand U28352 (N_28352,N_22449,N_22015);
or U28353 (N_28353,N_22226,N_21930);
and U28354 (N_28354,N_20416,N_20556);
or U28355 (N_28355,N_22868,N_20534);
xor U28356 (N_28356,N_20744,N_23047);
and U28357 (N_28357,N_23309,N_23790);
and U28358 (N_28358,N_22596,N_20614);
nor U28359 (N_28359,N_21565,N_21090);
nand U28360 (N_28360,N_21101,N_20282);
nor U28361 (N_28361,N_23383,N_21248);
or U28362 (N_28362,N_22933,N_21008);
nand U28363 (N_28363,N_24688,N_22609);
xor U28364 (N_28364,N_24977,N_21711);
nor U28365 (N_28365,N_22492,N_24897);
nand U28366 (N_28366,N_21539,N_20565);
or U28367 (N_28367,N_22977,N_23029);
nor U28368 (N_28368,N_24935,N_20804);
and U28369 (N_28369,N_21787,N_21086);
xor U28370 (N_28370,N_22995,N_21175);
and U28371 (N_28371,N_21817,N_21662);
nor U28372 (N_28372,N_22012,N_22565);
and U28373 (N_28373,N_20563,N_23895);
nand U28374 (N_28374,N_20480,N_21257);
nor U28375 (N_28375,N_24388,N_20327);
nor U28376 (N_28376,N_23199,N_21666);
nor U28377 (N_28377,N_21598,N_20891);
xor U28378 (N_28378,N_22892,N_24257);
and U28379 (N_28379,N_21276,N_24118);
or U28380 (N_28380,N_23753,N_22830);
and U28381 (N_28381,N_24896,N_21119);
xnor U28382 (N_28382,N_21389,N_21450);
xnor U28383 (N_28383,N_21708,N_20875);
xor U28384 (N_28384,N_20926,N_23416);
or U28385 (N_28385,N_21032,N_24032);
or U28386 (N_28386,N_24405,N_21824);
or U28387 (N_28387,N_22234,N_22660);
or U28388 (N_28388,N_21028,N_23445);
xnor U28389 (N_28389,N_23384,N_20109);
nand U28390 (N_28390,N_24921,N_23993);
nor U28391 (N_28391,N_20636,N_20012);
nor U28392 (N_28392,N_24317,N_22891);
or U28393 (N_28393,N_23135,N_21518);
or U28394 (N_28394,N_24212,N_24413);
xor U28395 (N_28395,N_22892,N_24403);
nor U28396 (N_28396,N_23330,N_21551);
nand U28397 (N_28397,N_20105,N_20179);
or U28398 (N_28398,N_20314,N_22412);
nor U28399 (N_28399,N_24933,N_22241);
nor U28400 (N_28400,N_23359,N_24098);
xor U28401 (N_28401,N_20312,N_20833);
xor U28402 (N_28402,N_23037,N_22987);
and U28403 (N_28403,N_24297,N_20517);
or U28404 (N_28404,N_21467,N_21885);
nand U28405 (N_28405,N_24995,N_22187);
nor U28406 (N_28406,N_24879,N_22707);
nand U28407 (N_28407,N_22006,N_21212);
and U28408 (N_28408,N_23152,N_21785);
nand U28409 (N_28409,N_22796,N_22583);
xor U28410 (N_28410,N_24596,N_21884);
or U28411 (N_28411,N_21497,N_24304);
xor U28412 (N_28412,N_24133,N_22706);
or U28413 (N_28413,N_21032,N_20950);
or U28414 (N_28414,N_20399,N_20858);
xor U28415 (N_28415,N_21895,N_21823);
or U28416 (N_28416,N_23204,N_20811);
nor U28417 (N_28417,N_21648,N_20628);
or U28418 (N_28418,N_21149,N_22886);
and U28419 (N_28419,N_24960,N_22707);
nand U28420 (N_28420,N_22814,N_24968);
and U28421 (N_28421,N_21787,N_20377);
nand U28422 (N_28422,N_21858,N_21105);
nor U28423 (N_28423,N_23387,N_22794);
and U28424 (N_28424,N_22601,N_23114);
xor U28425 (N_28425,N_21275,N_24420);
nand U28426 (N_28426,N_24620,N_22164);
and U28427 (N_28427,N_22845,N_24981);
and U28428 (N_28428,N_22758,N_20240);
xor U28429 (N_28429,N_20933,N_23608);
and U28430 (N_28430,N_22260,N_20077);
nor U28431 (N_28431,N_21235,N_24801);
nor U28432 (N_28432,N_24533,N_20167);
nor U28433 (N_28433,N_24508,N_24764);
or U28434 (N_28434,N_22708,N_24456);
or U28435 (N_28435,N_20044,N_22995);
or U28436 (N_28436,N_24646,N_20633);
or U28437 (N_28437,N_24854,N_20178);
or U28438 (N_28438,N_20155,N_23409);
nand U28439 (N_28439,N_23450,N_21535);
nor U28440 (N_28440,N_22826,N_22078);
or U28441 (N_28441,N_22993,N_23531);
and U28442 (N_28442,N_24396,N_21705);
and U28443 (N_28443,N_22495,N_22297);
xnor U28444 (N_28444,N_22415,N_24289);
nor U28445 (N_28445,N_23990,N_24025);
xor U28446 (N_28446,N_21679,N_24978);
and U28447 (N_28447,N_24068,N_23251);
or U28448 (N_28448,N_20502,N_23579);
or U28449 (N_28449,N_23197,N_23646);
xnor U28450 (N_28450,N_20922,N_21768);
nand U28451 (N_28451,N_23795,N_20883);
or U28452 (N_28452,N_20581,N_23849);
nor U28453 (N_28453,N_24443,N_23478);
nor U28454 (N_28454,N_21543,N_22173);
xnor U28455 (N_28455,N_21905,N_23351);
nor U28456 (N_28456,N_23519,N_21975);
and U28457 (N_28457,N_21161,N_20225);
nor U28458 (N_28458,N_24422,N_20770);
nor U28459 (N_28459,N_24504,N_24302);
nand U28460 (N_28460,N_22666,N_24311);
xor U28461 (N_28461,N_20800,N_22189);
nand U28462 (N_28462,N_22756,N_23661);
xnor U28463 (N_28463,N_23521,N_24732);
nor U28464 (N_28464,N_23620,N_23475);
nor U28465 (N_28465,N_23853,N_21566);
xor U28466 (N_28466,N_24449,N_24283);
xor U28467 (N_28467,N_22798,N_20039);
and U28468 (N_28468,N_23478,N_22802);
nand U28469 (N_28469,N_21839,N_23620);
and U28470 (N_28470,N_23572,N_22341);
nand U28471 (N_28471,N_24716,N_22855);
or U28472 (N_28472,N_21598,N_20472);
xnor U28473 (N_28473,N_21699,N_23746);
nor U28474 (N_28474,N_22822,N_24686);
nor U28475 (N_28475,N_20135,N_23059);
nand U28476 (N_28476,N_24190,N_24321);
nand U28477 (N_28477,N_21954,N_21999);
nand U28478 (N_28478,N_22849,N_22003);
xnor U28479 (N_28479,N_24040,N_24545);
nor U28480 (N_28480,N_23903,N_23101);
nand U28481 (N_28481,N_22844,N_21874);
or U28482 (N_28482,N_21272,N_22700);
and U28483 (N_28483,N_22296,N_23870);
nand U28484 (N_28484,N_23014,N_24089);
and U28485 (N_28485,N_23278,N_22983);
and U28486 (N_28486,N_22464,N_22104);
nor U28487 (N_28487,N_24833,N_24304);
and U28488 (N_28488,N_24266,N_24799);
nand U28489 (N_28489,N_21821,N_20587);
or U28490 (N_28490,N_22934,N_23405);
xor U28491 (N_28491,N_22235,N_22003);
or U28492 (N_28492,N_20130,N_20693);
or U28493 (N_28493,N_20552,N_20683);
and U28494 (N_28494,N_20029,N_21078);
nand U28495 (N_28495,N_21202,N_21164);
nand U28496 (N_28496,N_23636,N_23974);
and U28497 (N_28497,N_22387,N_23719);
xor U28498 (N_28498,N_22887,N_20715);
and U28499 (N_28499,N_23198,N_23090);
xor U28500 (N_28500,N_21375,N_21737);
xor U28501 (N_28501,N_20894,N_20934);
or U28502 (N_28502,N_20016,N_20400);
nor U28503 (N_28503,N_23404,N_22909);
nand U28504 (N_28504,N_22968,N_23071);
nor U28505 (N_28505,N_23459,N_23524);
or U28506 (N_28506,N_23960,N_23399);
or U28507 (N_28507,N_24259,N_21382);
nor U28508 (N_28508,N_24874,N_22822);
and U28509 (N_28509,N_22134,N_21675);
nor U28510 (N_28510,N_20805,N_21350);
or U28511 (N_28511,N_21695,N_22472);
nand U28512 (N_28512,N_20487,N_24996);
nand U28513 (N_28513,N_24913,N_23043);
xnor U28514 (N_28514,N_22592,N_22654);
and U28515 (N_28515,N_23331,N_24593);
or U28516 (N_28516,N_23629,N_22533);
and U28517 (N_28517,N_23313,N_20513);
xor U28518 (N_28518,N_20945,N_20917);
and U28519 (N_28519,N_20464,N_24882);
nand U28520 (N_28520,N_22738,N_22290);
and U28521 (N_28521,N_22091,N_23363);
nand U28522 (N_28522,N_20804,N_21520);
xnor U28523 (N_28523,N_20537,N_23760);
and U28524 (N_28524,N_24176,N_22460);
and U28525 (N_28525,N_20036,N_20244);
nand U28526 (N_28526,N_23561,N_21519);
or U28527 (N_28527,N_24196,N_23655);
nand U28528 (N_28528,N_23091,N_20829);
or U28529 (N_28529,N_22655,N_21519);
nor U28530 (N_28530,N_23741,N_22469);
xnor U28531 (N_28531,N_24080,N_21143);
or U28532 (N_28532,N_24816,N_21574);
xnor U28533 (N_28533,N_21341,N_22580);
nor U28534 (N_28534,N_21962,N_20640);
or U28535 (N_28535,N_23764,N_20214);
xnor U28536 (N_28536,N_24541,N_22019);
xnor U28537 (N_28537,N_24725,N_22358);
xnor U28538 (N_28538,N_20540,N_22489);
and U28539 (N_28539,N_24050,N_20569);
xor U28540 (N_28540,N_24013,N_22037);
nor U28541 (N_28541,N_22512,N_21115);
xnor U28542 (N_28542,N_23570,N_20158);
xnor U28543 (N_28543,N_23098,N_23120);
or U28544 (N_28544,N_24395,N_21627);
xnor U28545 (N_28545,N_20095,N_23025);
and U28546 (N_28546,N_20766,N_24596);
nor U28547 (N_28547,N_24726,N_23186);
and U28548 (N_28548,N_24464,N_24783);
nor U28549 (N_28549,N_22585,N_23207);
and U28550 (N_28550,N_24653,N_23045);
nand U28551 (N_28551,N_24065,N_24579);
nor U28552 (N_28552,N_22085,N_23030);
xor U28553 (N_28553,N_21685,N_22734);
xnor U28554 (N_28554,N_22721,N_22576);
nand U28555 (N_28555,N_23808,N_23172);
or U28556 (N_28556,N_20422,N_20259);
nor U28557 (N_28557,N_23426,N_24870);
nor U28558 (N_28558,N_20389,N_21197);
xor U28559 (N_28559,N_20333,N_22741);
nand U28560 (N_28560,N_22826,N_22772);
nor U28561 (N_28561,N_21358,N_22408);
nor U28562 (N_28562,N_23110,N_20436);
nand U28563 (N_28563,N_20294,N_22009);
or U28564 (N_28564,N_20806,N_23532);
and U28565 (N_28565,N_23112,N_23024);
nor U28566 (N_28566,N_24329,N_20116);
and U28567 (N_28567,N_20294,N_24707);
nand U28568 (N_28568,N_21609,N_22393);
or U28569 (N_28569,N_20164,N_20393);
and U28570 (N_28570,N_22197,N_24726);
or U28571 (N_28571,N_21778,N_24260);
nor U28572 (N_28572,N_21565,N_22214);
xor U28573 (N_28573,N_23078,N_20575);
nor U28574 (N_28574,N_24679,N_21229);
nand U28575 (N_28575,N_24503,N_23742);
nand U28576 (N_28576,N_23376,N_21989);
nand U28577 (N_28577,N_24787,N_22591);
xnor U28578 (N_28578,N_21044,N_23190);
nand U28579 (N_28579,N_24274,N_21201);
nand U28580 (N_28580,N_21756,N_21353);
nor U28581 (N_28581,N_23279,N_20883);
xor U28582 (N_28582,N_24636,N_22946);
and U28583 (N_28583,N_23317,N_24813);
or U28584 (N_28584,N_24180,N_23812);
nor U28585 (N_28585,N_22531,N_20149);
and U28586 (N_28586,N_22117,N_21872);
and U28587 (N_28587,N_24377,N_20280);
nand U28588 (N_28588,N_23292,N_21413);
and U28589 (N_28589,N_23615,N_21412);
nand U28590 (N_28590,N_24804,N_20832);
nor U28591 (N_28591,N_21314,N_24603);
nor U28592 (N_28592,N_20669,N_21154);
xnor U28593 (N_28593,N_24516,N_22272);
and U28594 (N_28594,N_20503,N_21006);
nor U28595 (N_28595,N_22359,N_21595);
nor U28596 (N_28596,N_21266,N_24475);
nand U28597 (N_28597,N_20740,N_23475);
xor U28598 (N_28598,N_21658,N_20781);
nand U28599 (N_28599,N_21923,N_24575);
or U28600 (N_28600,N_23857,N_22595);
xor U28601 (N_28601,N_22649,N_23563);
or U28602 (N_28602,N_24137,N_24394);
and U28603 (N_28603,N_20509,N_22137);
nor U28604 (N_28604,N_24502,N_22342);
nor U28605 (N_28605,N_23976,N_21753);
and U28606 (N_28606,N_24809,N_22782);
nor U28607 (N_28607,N_21974,N_23796);
nor U28608 (N_28608,N_21950,N_23743);
or U28609 (N_28609,N_23341,N_21904);
nor U28610 (N_28610,N_24479,N_23251);
and U28611 (N_28611,N_24178,N_22419);
nand U28612 (N_28612,N_23361,N_20175);
nand U28613 (N_28613,N_20009,N_23460);
xnor U28614 (N_28614,N_24486,N_20838);
nand U28615 (N_28615,N_21118,N_22660);
or U28616 (N_28616,N_20530,N_24115);
nand U28617 (N_28617,N_24447,N_20312);
nand U28618 (N_28618,N_24197,N_24261);
or U28619 (N_28619,N_21029,N_20007);
nand U28620 (N_28620,N_22675,N_21559);
and U28621 (N_28621,N_20760,N_20415);
or U28622 (N_28622,N_20029,N_23487);
or U28623 (N_28623,N_22213,N_23950);
and U28624 (N_28624,N_20398,N_21024);
nor U28625 (N_28625,N_23091,N_20544);
xor U28626 (N_28626,N_23210,N_24763);
xor U28627 (N_28627,N_23650,N_23708);
nor U28628 (N_28628,N_24427,N_23920);
or U28629 (N_28629,N_20012,N_22505);
nor U28630 (N_28630,N_21508,N_20345);
nand U28631 (N_28631,N_24327,N_23084);
or U28632 (N_28632,N_24012,N_21447);
and U28633 (N_28633,N_24824,N_20900);
nand U28634 (N_28634,N_24262,N_24567);
nor U28635 (N_28635,N_20596,N_20188);
nor U28636 (N_28636,N_22561,N_23809);
or U28637 (N_28637,N_22283,N_22981);
or U28638 (N_28638,N_20948,N_21969);
nor U28639 (N_28639,N_20846,N_22252);
nand U28640 (N_28640,N_20852,N_20538);
nand U28641 (N_28641,N_22754,N_20579);
nor U28642 (N_28642,N_21850,N_23738);
xor U28643 (N_28643,N_21287,N_23449);
and U28644 (N_28644,N_22598,N_23036);
and U28645 (N_28645,N_21680,N_24637);
nor U28646 (N_28646,N_20029,N_23009);
and U28647 (N_28647,N_22542,N_20545);
xor U28648 (N_28648,N_24450,N_23343);
nand U28649 (N_28649,N_24605,N_23257);
nand U28650 (N_28650,N_21405,N_22196);
xnor U28651 (N_28651,N_22821,N_21125);
nand U28652 (N_28652,N_24144,N_24648);
nand U28653 (N_28653,N_21206,N_20723);
xor U28654 (N_28654,N_22639,N_22643);
nand U28655 (N_28655,N_20334,N_22284);
or U28656 (N_28656,N_22595,N_24718);
nor U28657 (N_28657,N_23295,N_22090);
nor U28658 (N_28658,N_23004,N_21016);
nor U28659 (N_28659,N_21717,N_22038);
nand U28660 (N_28660,N_20261,N_24277);
nand U28661 (N_28661,N_21241,N_23383);
or U28662 (N_28662,N_21292,N_24713);
and U28663 (N_28663,N_24453,N_22675);
nor U28664 (N_28664,N_20518,N_24774);
and U28665 (N_28665,N_24151,N_24118);
or U28666 (N_28666,N_20555,N_22530);
xor U28667 (N_28667,N_22552,N_22805);
and U28668 (N_28668,N_20342,N_24118);
xor U28669 (N_28669,N_24466,N_20412);
nand U28670 (N_28670,N_22053,N_24765);
nand U28671 (N_28671,N_21097,N_20285);
xor U28672 (N_28672,N_24242,N_23251);
nand U28673 (N_28673,N_20769,N_23825);
nand U28674 (N_28674,N_21413,N_20664);
or U28675 (N_28675,N_21906,N_22463);
nand U28676 (N_28676,N_22294,N_24539);
xor U28677 (N_28677,N_21119,N_22545);
xor U28678 (N_28678,N_22865,N_22569);
and U28679 (N_28679,N_22086,N_22215);
nor U28680 (N_28680,N_23157,N_22007);
and U28681 (N_28681,N_23537,N_20464);
or U28682 (N_28682,N_22876,N_20823);
or U28683 (N_28683,N_21752,N_24759);
nor U28684 (N_28684,N_24684,N_20190);
xnor U28685 (N_28685,N_20116,N_23121);
or U28686 (N_28686,N_23540,N_23712);
and U28687 (N_28687,N_23998,N_21991);
nor U28688 (N_28688,N_23683,N_21261);
nor U28689 (N_28689,N_20579,N_24348);
or U28690 (N_28690,N_20289,N_22460);
nand U28691 (N_28691,N_22687,N_21834);
xor U28692 (N_28692,N_20259,N_20443);
nor U28693 (N_28693,N_23304,N_20886);
nand U28694 (N_28694,N_20007,N_22305);
xor U28695 (N_28695,N_21009,N_23796);
nor U28696 (N_28696,N_23718,N_24282);
xnor U28697 (N_28697,N_24683,N_20169);
nand U28698 (N_28698,N_24766,N_21185);
nor U28699 (N_28699,N_23122,N_20376);
nor U28700 (N_28700,N_21375,N_22597);
nor U28701 (N_28701,N_21153,N_20336);
or U28702 (N_28702,N_22679,N_23021);
nand U28703 (N_28703,N_23896,N_23459);
or U28704 (N_28704,N_21024,N_21062);
nand U28705 (N_28705,N_21137,N_22977);
xor U28706 (N_28706,N_23864,N_23505);
and U28707 (N_28707,N_20580,N_22985);
nor U28708 (N_28708,N_21680,N_23253);
nor U28709 (N_28709,N_20012,N_24980);
or U28710 (N_28710,N_21349,N_20346);
nand U28711 (N_28711,N_22582,N_23824);
nand U28712 (N_28712,N_22081,N_20661);
xor U28713 (N_28713,N_22105,N_24419);
nand U28714 (N_28714,N_21225,N_20217);
or U28715 (N_28715,N_24873,N_23633);
or U28716 (N_28716,N_22091,N_21024);
or U28717 (N_28717,N_20474,N_24672);
nand U28718 (N_28718,N_23196,N_23064);
and U28719 (N_28719,N_24228,N_21776);
nand U28720 (N_28720,N_22967,N_21278);
nand U28721 (N_28721,N_23109,N_21368);
and U28722 (N_28722,N_23383,N_22640);
and U28723 (N_28723,N_20310,N_24483);
or U28724 (N_28724,N_23750,N_21855);
or U28725 (N_28725,N_23487,N_21754);
and U28726 (N_28726,N_22565,N_22539);
xor U28727 (N_28727,N_20894,N_20591);
nor U28728 (N_28728,N_23631,N_24148);
nor U28729 (N_28729,N_23559,N_22640);
and U28730 (N_28730,N_23381,N_21885);
xor U28731 (N_28731,N_21580,N_21348);
nor U28732 (N_28732,N_23351,N_20421);
or U28733 (N_28733,N_21765,N_23327);
or U28734 (N_28734,N_20905,N_21477);
nand U28735 (N_28735,N_21018,N_23895);
nand U28736 (N_28736,N_23213,N_22646);
xnor U28737 (N_28737,N_23981,N_23286);
or U28738 (N_28738,N_23826,N_22501);
or U28739 (N_28739,N_24711,N_20477);
or U28740 (N_28740,N_23004,N_23378);
xor U28741 (N_28741,N_23256,N_23961);
and U28742 (N_28742,N_22270,N_22746);
xor U28743 (N_28743,N_20788,N_20781);
or U28744 (N_28744,N_24996,N_23589);
xnor U28745 (N_28745,N_22994,N_23703);
nand U28746 (N_28746,N_24415,N_21899);
nor U28747 (N_28747,N_24177,N_22194);
xnor U28748 (N_28748,N_21856,N_22256);
and U28749 (N_28749,N_24066,N_23218);
or U28750 (N_28750,N_20870,N_23468);
nor U28751 (N_28751,N_20269,N_20097);
and U28752 (N_28752,N_22607,N_23383);
xor U28753 (N_28753,N_22739,N_20534);
xor U28754 (N_28754,N_24064,N_22819);
xor U28755 (N_28755,N_22977,N_21049);
nor U28756 (N_28756,N_21632,N_21963);
and U28757 (N_28757,N_20663,N_23307);
or U28758 (N_28758,N_20994,N_23499);
nor U28759 (N_28759,N_24682,N_23122);
xor U28760 (N_28760,N_22504,N_20984);
and U28761 (N_28761,N_23081,N_21502);
nand U28762 (N_28762,N_20371,N_23236);
nand U28763 (N_28763,N_20955,N_20862);
xnor U28764 (N_28764,N_24299,N_23290);
nand U28765 (N_28765,N_20717,N_20382);
or U28766 (N_28766,N_24708,N_24552);
or U28767 (N_28767,N_24893,N_24479);
nand U28768 (N_28768,N_22189,N_22112);
nand U28769 (N_28769,N_22213,N_21919);
and U28770 (N_28770,N_20633,N_24914);
nand U28771 (N_28771,N_21777,N_22804);
xor U28772 (N_28772,N_22082,N_20835);
or U28773 (N_28773,N_20225,N_20007);
nand U28774 (N_28774,N_20045,N_22761);
nor U28775 (N_28775,N_21118,N_21511);
or U28776 (N_28776,N_20032,N_23607);
nor U28777 (N_28777,N_20990,N_24420);
and U28778 (N_28778,N_22885,N_22286);
nand U28779 (N_28779,N_24634,N_20007);
and U28780 (N_28780,N_21422,N_22857);
nor U28781 (N_28781,N_22035,N_21935);
xnor U28782 (N_28782,N_20409,N_20372);
or U28783 (N_28783,N_21637,N_24531);
nor U28784 (N_28784,N_22192,N_21536);
nand U28785 (N_28785,N_23192,N_24691);
and U28786 (N_28786,N_21936,N_22908);
and U28787 (N_28787,N_20847,N_21054);
or U28788 (N_28788,N_20540,N_20199);
or U28789 (N_28789,N_23878,N_24530);
nor U28790 (N_28790,N_22492,N_22643);
and U28791 (N_28791,N_22148,N_23598);
and U28792 (N_28792,N_22069,N_20425);
or U28793 (N_28793,N_20367,N_22849);
and U28794 (N_28794,N_24332,N_24765);
xor U28795 (N_28795,N_21720,N_22957);
nor U28796 (N_28796,N_24952,N_23263);
or U28797 (N_28797,N_20673,N_20074);
or U28798 (N_28798,N_24472,N_21660);
and U28799 (N_28799,N_23487,N_22445);
and U28800 (N_28800,N_21878,N_21476);
or U28801 (N_28801,N_23318,N_23455);
xnor U28802 (N_28802,N_21636,N_24613);
and U28803 (N_28803,N_24325,N_22809);
nand U28804 (N_28804,N_20117,N_23649);
nor U28805 (N_28805,N_24168,N_20455);
nor U28806 (N_28806,N_23545,N_22485);
xnor U28807 (N_28807,N_21034,N_21881);
and U28808 (N_28808,N_24742,N_21525);
nand U28809 (N_28809,N_22289,N_24749);
xor U28810 (N_28810,N_22428,N_21124);
and U28811 (N_28811,N_24755,N_21077);
and U28812 (N_28812,N_22985,N_20833);
and U28813 (N_28813,N_20244,N_24605);
or U28814 (N_28814,N_20216,N_20883);
and U28815 (N_28815,N_24078,N_24465);
or U28816 (N_28816,N_20881,N_20769);
xor U28817 (N_28817,N_21325,N_22370);
nand U28818 (N_28818,N_22259,N_21139);
nand U28819 (N_28819,N_20657,N_22835);
nor U28820 (N_28820,N_20535,N_21563);
nand U28821 (N_28821,N_20689,N_23844);
xnor U28822 (N_28822,N_24784,N_21447);
nand U28823 (N_28823,N_20844,N_24373);
nand U28824 (N_28824,N_22123,N_21587);
xor U28825 (N_28825,N_23697,N_21756);
nand U28826 (N_28826,N_21004,N_24324);
nand U28827 (N_28827,N_22402,N_24021);
nor U28828 (N_28828,N_20061,N_23019);
or U28829 (N_28829,N_23079,N_21448);
nor U28830 (N_28830,N_21527,N_24144);
or U28831 (N_28831,N_24572,N_24373);
nand U28832 (N_28832,N_20037,N_22530);
and U28833 (N_28833,N_24743,N_23657);
and U28834 (N_28834,N_21450,N_21889);
and U28835 (N_28835,N_22009,N_21614);
or U28836 (N_28836,N_23712,N_21671);
and U28837 (N_28837,N_23800,N_24939);
xor U28838 (N_28838,N_24314,N_23855);
and U28839 (N_28839,N_21948,N_22795);
nor U28840 (N_28840,N_20922,N_22830);
and U28841 (N_28841,N_21041,N_22347);
or U28842 (N_28842,N_23677,N_23888);
or U28843 (N_28843,N_21276,N_20616);
and U28844 (N_28844,N_21776,N_21117);
and U28845 (N_28845,N_23607,N_22751);
or U28846 (N_28846,N_23189,N_20550);
xor U28847 (N_28847,N_22850,N_23242);
and U28848 (N_28848,N_24469,N_22838);
nand U28849 (N_28849,N_20056,N_22625);
or U28850 (N_28850,N_21973,N_21328);
and U28851 (N_28851,N_20566,N_23553);
nor U28852 (N_28852,N_24090,N_21834);
xor U28853 (N_28853,N_23403,N_21659);
and U28854 (N_28854,N_23952,N_24447);
or U28855 (N_28855,N_24158,N_23194);
nand U28856 (N_28856,N_24310,N_24787);
and U28857 (N_28857,N_24912,N_23645);
nand U28858 (N_28858,N_23435,N_20939);
or U28859 (N_28859,N_20447,N_23070);
or U28860 (N_28860,N_24563,N_24067);
or U28861 (N_28861,N_22408,N_24650);
nand U28862 (N_28862,N_24114,N_20833);
nand U28863 (N_28863,N_24191,N_22632);
and U28864 (N_28864,N_22991,N_20813);
and U28865 (N_28865,N_21689,N_20934);
nor U28866 (N_28866,N_22283,N_20248);
xor U28867 (N_28867,N_23697,N_23471);
xnor U28868 (N_28868,N_23649,N_23240);
xnor U28869 (N_28869,N_22026,N_22602);
xnor U28870 (N_28870,N_24698,N_22006);
xor U28871 (N_28871,N_21413,N_22203);
or U28872 (N_28872,N_21931,N_21941);
and U28873 (N_28873,N_20568,N_20855);
or U28874 (N_28874,N_21656,N_23960);
xor U28875 (N_28875,N_21906,N_21034);
xnor U28876 (N_28876,N_23602,N_22923);
and U28877 (N_28877,N_24050,N_20897);
nand U28878 (N_28878,N_20655,N_24820);
xnor U28879 (N_28879,N_23060,N_22957);
xnor U28880 (N_28880,N_24111,N_23143);
xor U28881 (N_28881,N_21836,N_24678);
nand U28882 (N_28882,N_21170,N_24969);
nand U28883 (N_28883,N_21772,N_24771);
and U28884 (N_28884,N_23249,N_21138);
nor U28885 (N_28885,N_21087,N_24858);
nand U28886 (N_28886,N_21404,N_23099);
and U28887 (N_28887,N_21753,N_22632);
or U28888 (N_28888,N_21290,N_21897);
and U28889 (N_28889,N_20559,N_23820);
nor U28890 (N_28890,N_20736,N_20758);
nand U28891 (N_28891,N_20938,N_22263);
xnor U28892 (N_28892,N_24029,N_22561);
or U28893 (N_28893,N_21669,N_24578);
and U28894 (N_28894,N_20687,N_22693);
and U28895 (N_28895,N_22964,N_22887);
nor U28896 (N_28896,N_20214,N_22795);
xnor U28897 (N_28897,N_24745,N_21800);
nand U28898 (N_28898,N_20584,N_24538);
xor U28899 (N_28899,N_23971,N_20554);
xnor U28900 (N_28900,N_22294,N_24235);
nor U28901 (N_28901,N_22028,N_22933);
or U28902 (N_28902,N_20201,N_24458);
and U28903 (N_28903,N_22045,N_23745);
xnor U28904 (N_28904,N_23520,N_23234);
xnor U28905 (N_28905,N_23132,N_24940);
or U28906 (N_28906,N_20719,N_24162);
xor U28907 (N_28907,N_24143,N_24862);
nand U28908 (N_28908,N_22565,N_23551);
nand U28909 (N_28909,N_24341,N_22443);
nor U28910 (N_28910,N_21670,N_23476);
xor U28911 (N_28911,N_23179,N_21750);
nor U28912 (N_28912,N_21951,N_20980);
xor U28913 (N_28913,N_23835,N_20109);
nor U28914 (N_28914,N_20465,N_22476);
or U28915 (N_28915,N_22333,N_24944);
or U28916 (N_28916,N_24680,N_24710);
nand U28917 (N_28917,N_23506,N_22847);
xor U28918 (N_28918,N_23211,N_20970);
or U28919 (N_28919,N_22562,N_20880);
and U28920 (N_28920,N_21242,N_21324);
and U28921 (N_28921,N_20142,N_21656);
nor U28922 (N_28922,N_21758,N_24046);
and U28923 (N_28923,N_20181,N_23352);
or U28924 (N_28924,N_21023,N_21733);
xor U28925 (N_28925,N_23921,N_22939);
or U28926 (N_28926,N_23053,N_22019);
nand U28927 (N_28927,N_22771,N_22105);
and U28928 (N_28928,N_23935,N_24698);
or U28929 (N_28929,N_20602,N_20056);
nor U28930 (N_28930,N_20541,N_22578);
or U28931 (N_28931,N_22508,N_23261);
or U28932 (N_28932,N_21105,N_24056);
nor U28933 (N_28933,N_24860,N_22821);
xnor U28934 (N_28934,N_23709,N_22737);
xor U28935 (N_28935,N_20702,N_20809);
or U28936 (N_28936,N_23898,N_20312);
nand U28937 (N_28937,N_22524,N_22395);
nand U28938 (N_28938,N_20448,N_20819);
nor U28939 (N_28939,N_21422,N_22305);
nor U28940 (N_28940,N_20954,N_21022);
xnor U28941 (N_28941,N_22894,N_21781);
nor U28942 (N_28942,N_22264,N_22342);
xnor U28943 (N_28943,N_22872,N_21774);
nor U28944 (N_28944,N_24185,N_23508);
or U28945 (N_28945,N_23456,N_20776);
nor U28946 (N_28946,N_24984,N_22805);
or U28947 (N_28947,N_20370,N_22991);
nor U28948 (N_28948,N_20951,N_22314);
nor U28949 (N_28949,N_21387,N_20309);
and U28950 (N_28950,N_20936,N_20614);
nand U28951 (N_28951,N_22049,N_24557);
nand U28952 (N_28952,N_20915,N_20422);
nor U28953 (N_28953,N_22969,N_24816);
nor U28954 (N_28954,N_20923,N_20598);
and U28955 (N_28955,N_23529,N_23641);
and U28956 (N_28956,N_22831,N_21054);
xnor U28957 (N_28957,N_20634,N_24707);
or U28958 (N_28958,N_24151,N_24495);
nand U28959 (N_28959,N_24388,N_22039);
nor U28960 (N_28960,N_20047,N_23790);
nor U28961 (N_28961,N_23332,N_21197);
nor U28962 (N_28962,N_22114,N_22719);
nand U28963 (N_28963,N_20063,N_22398);
or U28964 (N_28964,N_22635,N_21498);
nor U28965 (N_28965,N_24723,N_21900);
and U28966 (N_28966,N_24929,N_22136);
and U28967 (N_28967,N_23610,N_21850);
or U28968 (N_28968,N_22990,N_24260);
nand U28969 (N_28969,N_20445,N_21911);
or U28970 (N_28970,N_20281,N_24796);
nand U28971 (N_28971,N_20362,N_23675);
and U28972 (N_28972,N_23878,N_21278);
nand U28973 (N_28973,N_21082,N_21325);
nor U28974 (N_28974,N_21400,N_24792);
nand U28975 (N_28975,N_24392,N_23138);
xor U28976 (N_28976,N_22436,N_20486);
and U28977 (N_28977,N_24954,N_21443);
xor U28978 (N_28978,N_22633,N_23263);
or U28979 (N_28979,N_22654,N_24533);
nand U28980 (N_28980,N_21589,N_22895);
xor U28981 (N_28981,N_21297,N_20803);
and U28982 (N_28982,N_21109,N_21809);
or U28983 (N_28983,N_23786,N_23069);
nor U28984 (N_28984,N_20350,N_22700);
xor U28985 (N_28985,N_23065,N_22815);
nand U28986 (N_28986,N_20820,N_23433);
xnor U28987 (N_28987,N_21250,N_21393);
or U28988 (N_28988,N_21861,N_20518);
nand U28989 (N_28989,N_24053,N_22209);
xor U28990 (N_28990,N_21305,N_22645);
xor U28991 (N_28991,N_21226,N_20746);
nand U28992 (N_28992,N_22519,N_24675);
and U28993 (N_28993,N_24744,N_21916);
or U28994 (N_28994,N_22451,N_24299);
nor U28995 (N_28995,N_20213,N_23020);
xor U28996 (N_28996,N_24661,N_20308);
nand U28997 (N_28997,N_23171,N_24260);
nand U28998 (N_28998,N_21016,N_22668);
and U28999 (N_28999,N_20931,N_24513);
and U29000 (N_29000,N_22721,N_22562);
xnor U29001 (N_29001,N_22115,N_24071);
nand U29002 (N_29002,N_21905,N_22831);
nor U29003 (N_29003,N_24389,N_24588);
or U29004 (N_29004,N_23273,N_23944);
xor U29005 (N_29005,N_23592,N_21000);
and U29006 (N_29006,N_21908,N_20113);
or U29007 (N_29007,N_21661,N_24440);
nor U29008 (N_29008,N_24162,N_21087);
and U29009 (N_29009,N_24769,N_22864);
xor U29010 (N_29010,N_24101,N_20712);
nor U29011 (N_29011,N_21029,N_20511);
nand U29012 (N_29012,N_20000,N_23369);
and U29013 (N_29013,N_20899,N_23385);
nor U29014 (N_29014,N_21217,N_23948);
nor U29015 (N_29015,N_23069,N_24682);
nand U29016 (N_29016,N_20107,N_24646);
and U29017 (N_29017,N_22076,N_21975);
and U29018 (N_29018,N_21616,N_22426);
and U29019 (N_29019,N_23814,N_20050);
or U29020 (N_29020,N_21384,N_20412);
or U29021 (N_29021,N_21468,N_20791);
nor U29022 (N_29022,N_20148,N_24666);
or U29023 (N_29023,N_22368,N_20448);
and U29024 (N_29024,N_22437,N_23065);
xor U29025 (N_29025,N_22769,N_23268);
and U29026 (N_29026,N_22971,N_24163);
or U29027 (N_29027,N_20084,N_24908);
nor U29028 (N_29028,N_20297,N_23791);
and U29029 (N_29029,N_21461,N_22303);
nand U29030 (N_29030,N_20749,N_21127);
nor U29031 (N_29031,N_21072,N_20560);
xor U29032 (N_29032,N_21948,N_21539);
and U29033 (N_29033,N_21204,N_24172);
nand U29034 (N_29034,N_24473,N_21655);
or U29035 (N_29035,N_23307,N_21596);
nand U29036 (N_29036,N_20188,N_22508);
and U29037 (N_29037,N_20096,N_20157);
nor U29038 (N_29038,N_20618,N_20017);
nand U29039 (N_29039,N_22766,N_20348);
or U29040 (N_29040,N_20107,N_24035);
and U29041 (N_29041,N_22281,N_23086);
nand U29042 (N_29042,N_21061,N_22004);
or U29043 (N_29043,N_20435,N_22361);
nor U29044 (N_29044,N_24276,N_21753);
xnor U29045 (N_29045,N_23087,N_20407);
nand U29046 (N_29046,N_24876,N_23396);
xnor U29047 (N_29047,N_24132,N_24083);
nand U29048 (N_29048,N_24600,N_23709);
or U29049 (N_29049,N_21323,N_22518);
nor U29050 (N_29050,N_20738,N_21055);
xor U29051 (N_29051,N_20409,N_23049);
xnor U29052 (N_29052,N_20183,N_23874);
or U29053 (N_29053,N_22280,N_21866);
and U29054 (N_29054,N_20533,N_20903);
or U29055 (N_29055,N_22376,N_23630);
or U29056 (N_29056,N_20708,N_21197);
nor U29057 (N_29057,N_23541,N_23733);
and U29058 (N_29058,N_23629,N_22926);
or U29059 (N_29059,N_21243,N_22376);
nand U29060 (N_29060,N_22184,N_24745);
and U29061 (N_29061,N_20425,N_20115);
and U29062 (N_29062,N_20073,N_23125);
and U29063 (N_29063,N_20027,N_21985);
and U29064 (N_29064,N_21878,N_20989);
nand U29065 (N_29065,N_23228,N_21887);
xor U29066 (N_29066,N_22331,N_24987);
nand U29067 (N_29067,N_21074,N_23696);
nor U29068 (N_29068,N_21672,N_21762);
or U29069 (N_29069,N_23838,N_22087);
xnor U29070 (N_29070,N_22617,N_23066);
xor U29071 (N_29071,N_20292,N_22409);
nor U29072 (N_29072,N_22940,N_22063);
and U29073 (N_29073,N_24071,N_21232);
and U29074 (N_29074,N_20490,N_22517);
nor U29075 (N_29075,N_20066,N_22707);
or U29076 (N_29076,N_21625,N_22135);
nor U29077 (N_29077,N_20351,N_23925);
nor U29078 (N_29078,N_24537,N_21316);
or U29079 (N_29079,N_23952,N_22745);
or U29080 (N_29080,N_24271,N_22909);
and U29081 (N_29081,N_23360,N_23394);
nand U29082 (N_29082,N_22098,N_24041);
xor U29083 (N_29083,N_20861,N_21974);
nor U29084 (N_29084,N_21769,N_23402);
nor U29085 (N_29085,N_20373,N_20255);
nor U29086 (N_29086,N_20045,N_22339);
and U29087 (N_29087,N_23382,N_24976);
nand U29088 (N_29088,N_22566,N_23972);
nand U29089 (N_29089,N_23893,N_21449);
nand U29090 (N_29090,N_20800,N_24518);
or U29091 (N_29091,N_23488,N_24383);
or U29092 (N_29092,N_20643,N_20700);
nand U29093 (N_29093,N_21405,N_21757);
or U29094 (N_29094,N_20887,N_23428);
and U29095 (N_29095,N_22373,N_22081);
and U29096 (N_29096,N_20618,N_21415);
nand U29097 (N_29097,N_23403,N_23236);
nor U29098 (N_29098,N_21000,N_22496);
nor U29099 (N_29099,N_21694,N_24590);
nor U29100 (N_29100,N_24452,N_23942);
or U29101 (N_29101,N_23082,N_22296);
nor U29102 (N_29102,N_20000,N_23755);
and U29103 (N_29103,N_21235,N_20152);
or U29104 (N_29104,N_21837,N_21929);
or U29105 (N_29105,N_21868,N_21431);
nor U29106 (N_29106,N_22381,N_23946);
nand U29107 (N_29107,N_24875,N_21954);
and U29108 (N_29108,N_23040,N_23980);
nand U29109 (N_29109,N_24312,N_24293);
nor U29110 (N_29110,N_21729,N_20831);
nor U29111 (N_29111,N_23823,N_23396);
or U29112 (N_29112,N_20938,N_20142);
nand U29113 (N_29113,N_21525,N_24357);
or U29114 (N_29114,N_22499,N_21926);
xnor U29115 (N_29115,N_22298,N_22597);
nand U29116 (N_29116,N_20633,N_20699);
or U29117 (N_29117,N_21390,N_21833);
nor U29118 (N_29118,N_20948,N_20980);
nand U29119 (N_29119,N_22317,N_21806);
and U29120 (N_29120,N_23739,N_24928);
or U29121 (N_29121,N_21331,N_24087);
nand U29122 (N_29122,N_20475,N_22207);
xnor U29123 (N_29123,N_21391,N_23753);
xnor U29124 (N_29124,N_22552,N_22407);
nor U29125 (N_29125,N_21554,N_24793);
and U29126 (N_29126,N_23484,N_21633);
or U29127 (N_29127,N_23677,N_24597);
and U29128 (N_29128,N_20907,N_23283);
nand U29129 (N_29129,N_20164,N_21939);
nand U29130 (N_29130,N_21382,N_20408);
nor U29131 (N_29131,N_20374,N_22049);
and U29132 (N_29132,N_21040,N_23108);
nor U29133 (N_29133,N_23328,N_24520);
xnor U29134 (N_29134,N_20662,N_22770);
nor U29135 (N_29135,N_20748,N_23988);
and U29136 (N_29136,N_24513,N_22849);
and U29137 (N_29137,N_24103,N_20189);
nor U29138 (N_29138,N_21297,N_22583);
or U29139 (N_29139,N_21887,N_21046);
xnor U29140 (N_29140,N_20902,N_22691);
nor U29141 (N_29141,N_21648,N_20051);
xnor U29142 (N_29142,N_24251,N_22136);
nor U29143 (N_29143,N_23189,N_21345);
or U29144 (N_29144,N_20157,N_23466);
or U29145 (N_29145,N_23276,N_23953);
and U29146 (N_29146,N_20545,N_24720);
xnor U29147 (N_29147,N_23754,N_20002);
and U29148 (N_29148,N_24720,N_23592);
nand U29149 (N_29149,N_23739,N_23842);
or U29150 (N_29150,N_21589,N_20475);
and U29151 (N_29151,N_22433,N_22745);
nand U29152 (N_29152,N_24637,N_22637);
and U29153 (N_29153,N_24676,N_21140);
xor U29154 (N_29154,N_24448,N_22110);
and U29155 (N_29155,N_23052,N_23873);
nor U29156 (N_29156,N_21083,N_21991);
or U29157 (N_29157,N_22282,N_22624);
or U29158 (N_29158,N_21744,N_22780);
nand U29159 (N_29159,N_23894,N_24715);
nor U29160 (N_29160,N_23960,N_24089);
nor U29161 (N_29161,N_24280,N_24744);
xnor U29162 (N_29162,N_21603,N_21195);
and U29163 (N_29163,N_20294,N_21565);
and U29164 (N_29164,N_22849,N_21362);
xor U29165 (N_29165,N_23647,N_21703);
nand U29166 (N_29166,N_22091,N_20282);
and U29167 (N_29167,N_22146,N_24316);
nand U29168 (N_29168,N_22296,N_23376);
and U29169 (N_29169,N_23907,N_23073);
and U29170 (N_29170,N_21575,N_20626);
nand U29171 (N_29171,N_23635,N_23612);
nor U29172 (N_29172,N_22080,N_23807);
nor U29173 (N_29173,N_21957,N_21425);
nor U29174 (N_29174,N_20007,N_22707);
or U29175 (N_29175,N_22707,N_21444);
and U29176 (N_29176,N_24639,N_22391);
xnor U29177 (N_29177,N_24664,N_24714);
nand U29178 (N_29178,N_24109,N_22626);
xnor U29179 (N_29179,N_20501,N_21525);
and U29180 (N_29180,N_22649,N_22127);
and U29181 (N_29181,N_21440,N_24198);
nor U29182 (N_29182,N_24681,N_22563);
nor U29183 (N_29183,N_24566,N_23149);
nor U29184 (N_29184,N_21703,N_20959);
nand U29185 (N_29185,N_23625,N_20722);
nor U29186 (N_29186,N_22639,N_21159);
nor U29187 (N_29187,N_20116,N_24544);
and U29188 (N_29188,N_23403,N_24722);
or U29189 (N_29189,N_23847,N_22468);
xnor U29190 (N_29190,N_24673,N_20122);
nand U29191 (N_29191,N_23287,N_24491);
or U29192 (N_29192,N_22557,N_22900);
nor U29193 (N_29193,N_22945,N_21416);
nand U29194 (N_29194,N_24637,N_20799);
and U29195 (N_29195,N_20834,N_24398);
nand U29196 (N_29196,N_24765,N_24192);
xnor U29197 (N_29197,N_22213,N_23242);
or U29198 (N_29198,N_21690,N_23163);
or U29199 (N_29199,N_21116,N_22257);
xnor U29200 (N_29200,N_23631,N_21424);
xor U29201 (N_29201,N_24781,N_20205);
or U29202 (N_29202,N_22110,N_21828);
xor U29203 (N_29203,N_23571,N_22920);
nand U29204 (N_29204,N_23869,N_21148);
or U29205 (N_29205,N_24286,N_24082);
or U29206 (N_29206,N_22011,N_21278);
nand U29207 (N_29207,N_22713,N_22687);
nand U29208 (N_29208,N_21380,N_23660);
nor U29209 (N_29209,N_20149,N_23266);
or U29210 (N_29210,N_24674,N_24087);
or U29211 (N_29211,N_21330,N_23563);
nor U29212 (N_29212,N_24462,N_22408);
or U29213 (N_29213,N_22895,N_24118);
nand U29214 (N_29214,N_24826,N_23403);
and U29215 (N_29215,N_20828,N_22628);
nand U29216 (N_29216,N_21506,N_20477);
and U29217 (N_29217,N_24333,N_20207);
or U29218 (N_29218,N_23860,N_24386);
nand U29219 (N_29219,N_21709,N_23877);
xor U29220 (N_29220,N_22974,N_20894);
or U29221 (N_29221,N_21057,N_22876);
and U29222 (N_29222,N_23617,N_24007);
nand U29223 (N_29223,N_21124,N_24154);
xnor U29224 (N_29224,N_24357,N_23975);
xor U29225 (N_29225,N_23357,N_20728);
nand U29226 (N_29226,N_23830,N_21596);
and U29227 (N_29227,N_21693,N_22431);
xor U29228 (N_29228,N_21327,N_22340);
and U29229 (N_29229,N_20542,N_22502);
and U29230 (N_29230,N_22322,N_24917);
nand U29231 (N_29231,N_23079,N_21152);
and U29232 (N_29232,N_22263,N_20720);
nor U29233 (N_29233,N_24197,N_20915);
xnor U29234 (N_29234,N_20504,N_22389);
xor U29235 (N_29235,N_23039,N_24721);
nand U29236 (N_29236,N_20752,N_23161);
and U29237 (N_29237,N_24168,N_24416);
or U29238 (N_29238,N_22995,N_24112);
nor U29239 (N_29239,N_22219,N_20533);
nor U29240 (N_29240,N_20184,N_21109);
nand U29241 (N_29241,N_24111,N_23455);
and U29242 (N_29242,N_21247,N_23049);
or U29243 (N_29243,N_22473,N_22448);
nor U29244 (N_29244,N_22561,N_23931);
xor U29245 (N_29245,N_21318,N_24784);
or U29246 (N_29246,N_23977,N_23777);
nor U29247 (N_29247,N_22042,N_23215);
or U29248 (N_29248,N_23300,N_24448);
nor U29249 (N_29249,N_23177,N_22628);
nand U29250 (N_29250,N_20508,N_22338);
nand U29251 (N_29251,N_22599,N_22443);
xnor U29252 (N_29252,N_21564,N_23754);
nand U29253 (N_29253,N_23855,N_24048);
and U29254 (N_29254,N_22764,N_23947);
nor U29255 (N_29255,N_23743,N_22315);
nand U29256 (N_29256,N_20753,N_24250);
nand U29257 (N_29257,N_20537,N_24622);
and U29258 (N_29258,N_22020,N_23884);
and U29259 (N_29259,N_20008,N_20181);
and U29260 (N_29260,N_23182,N_21180);
or U29261 (N_29261,N_21322,N_23822);
xnor U29262 (N_29262,N_23486,N_23849);
xor U29263 (N_29263,N_23789,N_20465);
nor U29264 (N_29264,N_23342,N_22283);
nor U29265 (N_29265,N_21896,N_22796);
nor U29266 (N_29266,N_20588,N_21860);
and U29267 (N_29267,N_20859,N_21551);
xnor U29268 (N_29268,N_24025,N_22374);
or U29269 (N_29269,N_20199,N_20001);
nand U29270 (N_29270,N_23477,N_21432);
xnor U29271 (N_29271,N_21837,N_21632);
nand U29272 (N_29272,N_22828,N_21762);
or U29273 (N_29273,N_22383,N_22682);
nor U29274 (N_29274,N_23912,N_21901);
and U29275 (N_29275,N_23587,N_21455);
xnor U29276 (N_29276,N_21244,N_21526);
xnor U29277 (N_29277,N_21405,N_24334);
or U29278 (N_29278,N_20193,N_24756);
xnor U29279 (N_29279,N_24626,N_22505);
or U29280 (N_29280,N_24657,N_20283);
or U29281 (N_29281,N_22096,N_21141);
and U29282 (N_29282,N_20063,N_20224);
and U29283 (N_29283,N_21692,N_22772);
nand U29284 (N_29284,N_23820,N_20548);
and U29285 (N_29285,N_22641,N_21259);
nor U29286 (N_29286,N_21310,N_22202);
or U29287 (N_29287,N_23881,N_20421);
and U29288 (N_29288,N_24151,N_20913);
and U29289 (N_29289,N_20017,N_24944);
nand U29290 (N_29290,N_24297,N_24304);
and U29291 (N_29291,N_24428,N_20261);
nand U29292 (N_29292,N_22432,N_22272);
nor U29293 (N_29293,N_24575,N_20770);
or U29294 (N_29294,N_24466,N_23909);
and U29295 (N_29295,N_20927,N_24440);
or U29296 (N_29296,N_24989,N_24198);
xnor U29297 (N_29297,N_21564,N_23036);
or U29298 (N_29298,N_24484,N_22856);
or U29299 (N_29299,N_22502,N_24184);
xnor U29300 (N_29300,N_22558,N_20156);
nor U29301 (N_29301,N_23465,N_23102);
nor U29302 (N_29302,N_21262,N_22522);
or U29303 (N_29303,N_22740,N_23628);
xor U29304 (N_29304,N_20387,N_21898);
and U29305 (N_29305,N_22157,N_24104);
and U29306 (N_29306,N_23378,N_24685);
or U29307 (N_29307,N_22311,N_22107);
and U29308 (N_29308,N_20317,N_22801);
nor U29309 (N_29309,N_21656,N_22079);
nand U29310 (N_29310,N_23510,N_22550);
and U29311 (N_29311,N_24856,N_24776);
or U29312 (N_29312,N_22214,N_23787);
xnor U29313 (N_29313,N_22490,N_21869);
nand U29314 (N_29314,N_22902,N_22719);
xnor U29315 (N_29315,N_23058,N_22693);
nor U29316 (N_29316,N_23332,N_20812);
nor U29317 (N_29317,N_24835,N_24337);
or U29318 (N_29318,N_22756,N_23407);
and U29319 (N_29319,N_20893,N_23596);
and U29320 (N_29320,N_23966,N_23291);
nand U29321 (N_29321,N_23767,N_23138);
xnor U29322 (N_29322,N_20850,N_24297);
nor U29323 (N_29323,N_23578,N_22521);
nand U29324 (N_29324,N_22810,N_22522);
xnor U29325 (N_29325,N_20877,N_22640);
and U29326 (N_29326,N_24199,N_20559);
xor U29327 (N_29327,N_23004,N_24174);
nand U29328 (N_29328,N_21255,N_20727);
and U29329 (N_29329,N_24178,N_21782);
or U29330 (N_29330,N_23771,N_20794);
or U29331 (N_29331,N_22685,N_23450);
or U29332 (N_29332,N_22829,N_22347);
nor U29333 (N_29333,N_24962,N_22080);
nand U29334 (N_29334,N_23378,N_23594);
nand U29335 (N_29335,N_20878,N_20319);
xor U29336 (N_29336,N_24304,N_23912);
and U29337 (N_29337,N_24825,N_22231);
nand U29338 (N_29338,N_24463,N_23418);
and U29339 (N_29339,N_22188,N_22765);
and U29340 (N_29340,N_23759,N_23226);
nand U29341 (N_29341,N_21363,N_22082);
nand U29342 (N_29342,N_24661,N_21839);
nand U29343 (N_29343,N_23435,N_22678);
xor U29344 (N_29344,N_24801,N_20691);
and U29345 (N_29345,N_24645,N_21450);
and U29346 (N_29346,N_24315,N_20796);
nor U29347 (N_29347,N_20330,N_23493);
nor U29348 (N_29348,N_24575,N_24152);
nor U29349 (N_29349,N_21969,N_24553);
xor U29350 (N_29350,N_20443,N_22622);
nand U29351 (N_29351,N_23591,N_20970);
and U29352 (N_29352,N_24872,N_20241);
xnor U29353 (N_29353,N_23722,N_21666);
and U29354 (N_29354,N_22160,N_22783);
nand U29355 (N_29355,N_21169,N_20855);
nand U29356 (N_29356,N_21413,N_21691);
xor U29357 (N_29357,N_24047,N_20511);
nor U29358 (N_29358,N_23198,N_23877);
and U29359 (N_29359,N_22855,N_22492);
xnor U29360 (N_29360,N_22286,N_24010);
nand U29361 (N_29361,N_20364,N_23022);
nor U29362 (N_29362,N_23364,N_24343);
xnor U29363 (N_29363,N_21625,N_21688);
or U29364 (N_29364,N_23573,N_23259);
nand U29365 (N_29365,N_23445,N_22017);
and U29366 (N_29366,N_24222,N_20266);
nand U29367 (N_29367,N_20318,N_24999);
or U29368 (N_29368,N_24922,N_20745);
or U29369 (N_29369,N_20919,N_21536);
nor U29370 (N_29370,N_24934,N_21660);
xnor U29371 (N_29371,N_20839,N_21430);
nand U29372 (N_29372,N_20463,N_20323);
and U29373 (N_29373,N_21947,N_22620);
nand U29374 (N_29374,N_21815,N_20881);
or U29375 (N_29375,N_20344,N_22497);
xor U29376 (N_29376,N_22229,N_24774);
nor U29377 (N_29377,N_21626,N_24636);
or U29378 (N_29378,N_21043,N_23215);
nand U29379 (N_29379,N_21801,N_24909);
nor U29380 (N_29380,N_22036,N_21722);
and U29381 (N_29381,N_24796,N_22344);
or U29382 (N_29382,N_24817,N_21165);
nand U29383 (N_29383,N_20996,N_20656);
and U29384 (N_29384,N_20801,N_21277);
or U29385 (N_29385,N_21013,N_23097);
xnor U29386 (N_29386,N_21947,N_22941);
xor U29387 (N_29387,N_24805,N_21342);
nor U29388 (N_29388,N_22767,N_24322);
xor U29389 (N_29389,N_22526,N_24125);
nand U29390 (N_29390,N_23585,N_20486);
nand U29391 (N_29391,N_23081,N_20374);
xor U29392 (N_29392,N_21958,N_23297);
and U29393 (N_29393,N_20242,N_24420);
nand U29394 (N_29394,N_22336,N_21251);
nand U29395 (N_29395,N_20090,N_22168);
xnor U29396 (N_29396,N_20534,N_22742);
xor U29397 (N_29397,N_21294,N_21480);
nor U29398 (N_29398,N_24794,N_23377);
nand U29399 (N_29399,N_21696,N_21538);
or U29400 (N_29400,N_21798,N_22873);
xnor U29401 (N_29401,N_21053,N_24038);
xor U29402 (N_29402,N_24660,N_22338);
or U29403 (N_29403,N_24996,N_24333);
xor U29404 (N_29404,N_22908,N_23357);
or U29405 (N_29405,N_23276,N_23678);
nor U29406 (N_29406,N_20473,N_20039);
or U29407 (N_29407,N_22928,N_24344);
nand U29408 (N_29408,N_23428,N_23772);
nor U29409 (N_29409,N_21431,N_24266);
nor U29410 (N_29410,N_22837,N_21467);
and U29411 (N_29411,N_23272,N_24303);
nor U29412 (N_29412,N_21974,N_24605);
and U29413 (N_29413,N_21139,N_20909);
nor U29414 (N_29414,N_24132,N_23936);
or U29415 (N_29415,N_20609,N_20494);
or U29416 (N_29416,N_22204,N_24903);
nand U29417 (N_29417,N_24379,N_24640);
nand U29418 (N_29418,N_23963,N_20235);
nor U29419 (N_29419,N_21778,N_24270);
and U29420 (N_29420,N_22429,N_21635);
or U29421 (N_29421,N_23903,N_23955);
nand U29422 (N_29422,N_21478,N_24022);
nand U29423 (N_29423,N_21976,N_21463);
nor U29424 (N_29424,N_20118,N_20156);
nor U29425 (N_29425,N_21847,N_21800);
or U29426 (N_29426,N_20761,N_20049);
xnor U29427 (N_29427,N_23924,N_22381);
nor U29428 (N_29428,N_23529,N_23944);
nor U29429 (N_29429,N_22523,N_23268);
and U29430 (N_29430,N_22332,N_20265);
or U29431 (N_29431,N_20902,N_20480);
or U29432 (N_29432,N_22655,N_21083);
nor U29433 (N_29433,N_20348,N_22140);
nor U29434 (N_29434,N_20297,N_22022);
and U29435 (N_29435,N_24689,N_23848);
xnor U29436 (N_29436,N_23552,N_23263);
or U29437 (N_29437,N_20489,N_22739);
xor U29438 (N_29438,N_21535,N_24497);
nor U29439 (N_29439,N_23036,N_20181);
and U29440 (N_29440,N_24342,N_20784);
nand U29441 (N_29441,N_22804,N_23431);
xor U29442 (N_29442,N_22800,N_21275);
or U29443 (N_29443,N_23045,N_23174);
nand U29444 (N_29444,N_21691,N_22761);
nand U29445 (N_29445,N_22756,N_24311);
xor U29446 (N_29446,N_21520,N_20533);
nand U29447 (N_29447,N_23779,N_23526);
nand U29448 (N_29448,N_23853,N_23399);
or U29449 (N_29449,N_23763,N_24774);
nand U29450 (N_29450,N_23235,N_24368);
nor U29451 (N_29451,N_21719,N_22232);
xor U29452 (N_29452,N_20259,N_20500);
and U29453 (N_29453,N_22874,N_23866);
nor U29454 (N_29454,N_20058,N_22662);
nand U29455 (N_29455,N_24220,N_22448);
and U29456 (N_29456,N_20402,N_24766);
xnor U29457 (N_29457,N_24629,N_21002);
nand U29458 (N_29458,N_21716,N_23393);
xor U29459 (N_29459,N_23565,N_24125);
xnor U29460 (N_29460,N_24482,N_22938);
and U29461 (N_29461,N_21567,N_24032);
xnor U29462 (N_29462,N_21177,N_21491);
nand U29463 (N_29463,N_22310,N_24051);
nor U29464 (N_29464,N_21321,N_23447);
nor U29465 (N_29465,N_20832,N_21996);
and U29466 (N_29466,N_20642,N_22135);
nand U29467 (N_29467,N_24603,N_24021);
and U29468 (N_29468,N_23850,N_24035);
or U29469 (N_29469,N_23096,N_23244);
xnor U29470 (N_29470,N_20515,N_22506);
and U29471 (N_29471,N_24919,N_21890);
or U29472 (N_29472,N_22066,N_24791);
or U29473 (N_29473,N_24923,N_21174);
or U29474 (N_29474,N_23773,N_23917);
xor U29475 (N_29475,N_24083,N_21710);
nor U29476 (N_29476,N_23783,N_23449);
nand U29477 (N_29477,N_23706,N_20565);
nor U29478 (N_29478,N_23179,N_23377);
xor U29479 (N_29479,N_23620,N_22880);
nand U29480 (N_29480,N_21335,N_23124);
nor U29481 (N_29481,N_20242,N_21580);
or U29482 (N_29482,N_24412,N_22723);
or U29483 (N_29483,N_22425,N_23839);
nor U29484 (N_29484,N_22864,N_22589);
or U29485 (N_29485,N_24279,N_22325);
or U29486 (N_29486,N_20181,N_22284);
nor U29487 (N_29487,N_23576,N_24039);
nand U29488 (N_29488,N_20023,N_20794);
nor U29489 (N_29489,N_21722,N_21944);
xnor U29490 (N_29490,N_23943,N_24569);
xor U29491 (N_29491,N_20329,N_23778);
and U29492 (N_29492,N_21777,N_21565);
nor U29493 (N_29493,N_23275,N_22564);
xnor U29494 (N_29494,N_22111,N_21184);
nor U29495 (N_29495,N_22205,N_23307);
nand U29496 (N_29496,N_21337,N_23805);
and U29497 (N_29497,N_22001,N_20915);
xnor U29498 (N_29498,N_24437,N_24250);
nand U29499 (N_29499,N_20778,N_24741);
and U29500 (N_29500,N_20623,N_24712);
nand U29501 (N_29501,N_21129,N_23795);
nor U29502 (N_29502,N_21862,N_23300);
or U29503 (N_29503,N_24756,N_23042);
nor U29504 (N_29504,N_20702,N_20329);
xnor U29505 (N_29505,N_20857,N_20013);
nor U29506 (N_29506,N_22730,N_23765);
or U29507 (N_29507,N_24729,N_21107);
or U29508 (N_29508,N_24224,N_23456);
nand U29509 (N_29509,N_21866,N_23677);
nor U29510 (N_29510,N_22376,N_21472);
nor U29511 (N_29511,N_23610,N_22040);
nand U29512 (N_29512,N_21117,N_20129);
xor U29513 (N_29513,N_24107,N_22580);
and U29514 (N_29514,N_23452,N_22834);
and U29515 (N_29515,N_22996,N_20761);
or U29516 (N_29516,N_24005,N_21498);
nand U29517 (N_29517,N_21737,N_22356);
or U29518 (N_29518,N_23475,N_24013);
nand U29519 (N_29519,N_21791,N_24327);
or U29520 (N_29520,N_24336,N_24130);
nor U29521 (N_29521,N_20994,N_21662);
xnor U29522 (N_29522,N_24140,N_23988);
nor U29523 (N_29523,N_22142,N_22823);
nor U29524 (N_29524,N_20014,N_20872);
xor U29525 (N_29525,N_24175,N_20105);
xnor U29526 (N_29526,N_20664,N_23495);
nor U29527 (N_29527,N_20495,N_23231);
or U29528 (N_29528,N_21660,N_24180);
nor U29529 (N_29529,N_24975,N_22316);
nor U29530 (N_29530,N_21009,N_21007);
and U29531 (N_29531,N_24969,N_20498);
xnor U29532 (N_29532,N_21028,N_20686);
or U29533 (N_29533,N_23101,N_20795);
xnor U29534 (N_29534,N_21460,N_22620);
and U29535 (N_29535,N_23571,N_21652);
nor U29536 (N_29536,N_20229,N_22086);
nand U29537 (N_29537,N_24862,N_20845);
or U29538 (N_29538,N_23544,N_21323);
or U29539 (N_29539,N_22887,N_20075);
or U29540 (N_29540,N_21602,N_24573);
nor U29541 (N_29541,N_23109,N_24448);
nand U29542 (N_29542,N_23647,N_20205);
xor U29543 (N_29543,N_24999,N_20064);
and U29544 (N_29544,N_21292,N_24859);
nor U29545 (N_29545,N_23170,N_22666);
nand U29546 (N_29546,N_24019,N_21430);
xnor U29547 (N_29547,N_21942,N_21748);
or U29548 (N_29548,N_21666,N_21524);
or U29549 (N_29549,N_22723,N_21149);
and U29550 (N_29550,N_20639,N_21838);
and U29551 (N_29551,N_23143,N_20144);
nor U29552 (N_29552,N_20751,N_23777);
or U29553 (N_29553,N_23850,N_21162);
xor U29554 (N_29554,N_20812,N_21341);
and U29555 (N_29555,N_24998,N_23783);
nor U29556 (N_29556,N_23009,N_22823);
nor U29557 (N_29557,N_22475,N_22017);
and U29558 (N_29558,N_22685,N_22093);
and U29559 (N_29559,N_23641,N_21003);
nand U29560 (N_29560,N_24915,N_22770);
xor U29561 (N_29561,N_20653,N_24826);
and U29562 (N_29562,N_24907,N_22855);
or U29563 (N_29563,N_21757,N_23576);
nand U29564 (N_29564,N_20106,N_23973);
and U29565 (N_29565,N_20771,N_20809);
nor U29566 (N_29566,N_21767,N_21014);
and U29567 (N_29567,N_21045,N_21154);
nand U29568 (N_29568,N_21160,N_24291);
xor U29569 (N_29569,N_21154,N_20987);
nor U29570 (N_29570,N_21614,N_21738);
nor U29571 (N_29571,N_21258,N_22052);
nor U29572 (N_29572,N_22535,N_20885);
nor U29573 (N_29573,N_23536,N_23439);
and U29574 (N_29574,N_24285,N_22682);
and U29575 (N_29575,N_21864,N_20501);
and U29576 (N_29576,N_23931,N_22599);
nor U29577 (N_29577,N_22553,N_21234);
xnor U29578 (N_29578,N_21787,N_20609);
xor U29579 (N_29579,N_23466,N_23576);
or U29580 (N_29580,N_24136,N_21400);
xor U29581 (N_29581,N_21286,N_21969);
or U29582 (N_29582,N_24079,N_22619);
and U29583 (N_29583,N_20716,N_24738);
or U29584 (N_29584,N_24936,N_23357);
or U29585 (N_29585,N_24978,N_20994);
xor U29586 (N_29586,N_23266,N_24756);
nor U29587 (N_29587,N_20031,N_24502);
xnor U29588 (N_29588,N_21112,N_22277);
and U29589 (N_29589,N_21047,N_20939);
and U29590 (N_29590,N_22872,N_22530);
or U29591 (N_29591,N_21539,N_24344);
nand U29592 (N_29592,N_21371,N_24006);
xor U29593 (N_29593,N_24703,N_22967);
nand U29594 (N_29594,N_20945,N_21229);
or U29595 (N_29595,N_24408,N_20794);
nor U29596 (N_29596,N_23281,N_24419);
xnor U29597 (N_29597,N_20652,N_21488);
nand U29598 (N_29598,N_23956,N_21006);
xnor U29599 (N_29599,N_20645,N_21113);
nor U29600 (N_29600,N_24447,N_22543);
and U29601 (N_29601,N_24155,N_23245);
xnor U29602 (N_29602,N_24048,N_23211);
nor U29603 (N_29603,N_20028,N_21577);
nor U29604 (N_29604,N_20965,N_22595);
xnor U29605 (N_29605,N_20604,N_23029);
and U29606 (N_29606,N_20449,N_20731);
nand U29607 (N_29607,N_20617,N_20803);
nand U29608 (N_29608,N_20570,N_22428);
or U29609 (N_29609,N_21125,N_21285);
and U29610 (N_29610,N_21553,N_22166);
nand U29611 (N_29611,N_21863,N_24429);
and U29612 (N_29612,N_24984,N_24818);
nor U29613 (N_29613,N_23612,N_23203);
nand U29614 (N_29614,N_22595,N_22714);
or U29615 (N_29615,N_22283,N_23384);
nor U29616 (N_29616,N_21739,N_22238);
nand U29617 (N_29617,N_24406,N_23176);
or U29618 (N_29618,N_21451,N_21042);
nor U29619 (N_29619,N_24222,N_23539);
or U29620 (N_29620,N_20723,N_24586);
or U29621 (N_29621,N_21853,N_23021);
or U29622 (N_29622,N_24130,N_23977);
nor U29623 (N_29623,N_20962,N_23620);
and U29624 (N_29624,N_23544,N_21106);
or U29625 (N_29625,N_24647,N_20097);
and U29626 (N_29626,N_24231,N_21164);
nand U29627 (N_29627,N_20148,N_20609);
nand U29628 (N_29628,N_20293,N_22731);
nor U29629 (N_29629,N_20708,N_21064);
nand U29630 (N_29630,N_20542,N_24379);
or U29631 (N_29631,N_22767,N_23878);
nand U29632 (N_29632,N_24078,N_20721);
nand U29633 (N_29633,N_20820,N_20268);
or U29634 (N_29634,N_23802,N_23599);
nor U29635 (N_29635,N_20233,N_20910);
nor U29636 (N_29636,N_22268,N_21271);
xor U29637 (N_29637,N_21598,N_24700);
nand U29638 (N_29638,N_20493,N_24175);
or U29639 (N_29639,N_22775,N_20546);
nor U29640 (N_29640,N_24950,N_24145);
xor U29641 (N_29641,N_20898,N_24941);
or U29642 (N_29642,N_23885,N_21188);
xor U29643 (N_29643,N_20425,N_22802);
and U29644 (N_29644,N_24449,N_24864);
or U29645 (N_29645,N_22748,N_24365);
nor U29646 (N_29646,N_23696,N_21110);
xnor U29647 (N_29647,N_21097,N_21433);
nand U29648 (N_29648,N_20054,N_22571);
and U29649 (N_29649,N_20488,N_23513);
nand U29650 (N_29650,N_24725,N_24336);
xor U29651 (N_29651,N_21839,N_21910);
xnor U29652 (N_29652,N_24499,N_24978);
and U29653 (N_29653,N_23913,N_24463);
and U29654 (N_29654,N_23779,N_21012);
nand U29655 (N_29655,N_24308,N_20711);
nor U29656 (N_29656,N_24106,N_22785);
nor U29657 (N_29657,N_20499,N_22892);
and U29658 (N_29658,N_20317,N_24755);
or U29659 (N_29659,N_24717,N_24238);
nand U29660 (N_29660,N_21686,N_24083);
or U29661 (N_29661,N_23223,N_20094);
nor U29662 (N_29662,N_24137,N_24690);
or U29663 (N_29663,N_23265,N_23746);
xnor U29664 (N_29664,N_24088,N_24452);
nor U29665 (N_29665,N_24202,N_23203);
xor U29666 (N_29666,N_23971,N_20884);
and U29667 (N_29667,N_21272,N_21951);
nor U29668 (N_29668,N_22005,N_22892);
or U29669 (N_29669,N_20155,N_20933);
nand U29670 (N_29670,N_23307,N_23635);
or U29671 (N_29671,N_23459,N_22114);
or U29672 (N_29672,N_23002,N_21068);
nand U29673 (N_29673,N_20294,N_21855);
and U29674 (N_29674,N_23457,N_24348);
nor U29675 (N_29675,N_24473,N_21185);
nand U29676 (N_29676,N_23845,N_23985);
or U29677 (N_29677,N_21455,N_22785);
nor U29678 (N_29678,N_24356,N_22577);
xnor U29679 (N_29679,N_20330,N_24628);
nor U29680 (N_29680,N_20359,N_23947);
nor U29681 (N_29681,N_20213,N_23806);
and U29682 (N_29682,N_23671,N_24526);
nor U29683 (N_29683,N_20556,N_20849);
nor U29684 (N_29684,N_20872,N_24061);
nand U29685 (N_29685,N_20890,N_22904);
nor U29686 (N_29686,N_23088,N_20741);
or U29687 (N_29687,N_22314,N_21005);
nor U29688 (N_29688,N_23535,N_21799);
and U29689 (N_29689,N_20728,N_23709);
or U29690 (N_29690,N_24039,N_23598);
nor U29691 (N_29691,N_22956,N_21275);
or U29692 (N_29692,N_24309,N_22653);
nor U29693 (N_29693,N_24116,N_22866);
nor U29694 (N_29694,N_24143,N_24254);
nand U29695 (N_29695,N_21776,N_22218);
or U29696 (N_29696,N_21442,N_20219);
xnor U29697 (N_29697,N_20739,N_22295);
nor U29698 (N_29698,N_24365,N_21059);
nor U29699 (N_29699,N_23380,N_23012);
nor U29700 (N_29700,N_22748,N_20985);
xor U29701 (N_29701,N_24502,N_21898);
nand U29702 (N_29702,N_23917,N_24603);
nand U29703 (N_29703,N_23128,N_22005);
and U29704 (N_29704,N_23424,N_23528);
xnor U29705 (N_29705,N_21384,N_22243);
or U29706 (N_29706,N_22612,N_22251);
xor U29707 (N_29707,N_21251,N_23041);
xnor U29708 (N_29708,N_21764,N_20375);
nand U29709 (N_29709,N_22234,N_22573);
xor U29710 (N_29710,N_21898,N_23102);
nor U29711 (N_29711,N_21595,N_20969);
or U29712 (N_29712,N_21098,N_21666);
xnor U29713 (N_29713,N_24966,N_22793);
nand U29714 (N_29714,N_24415,N_24781);
nand U29715 (N_29715,N_21045,N_22003);
nor U29716 (N_29716,N_22818,N_20362);
nor U29717 (N_29717,N_24871,N_21676);
nand U29718 (N_29718,N_24025,N_22302);
nor U29719 (N_29719,N_22566,N_20988);
xnor U29720 (N_29720,N_22553,N_24513);
or U29721 (N_29721,N_24703,N_23521);
nand U29722 (N_29722,N_20339,N_23655);
nand U29723 (N_29723,N_20509,N_23440);
xnor U29724 (N_29724,N_22382,N_24015);
and U29725 (N_29725,N_23385,N_21766);
or U29726 (N_29726,N_24516,N_24434);
and U29727 (N_29727,N_20604,N_22690);
or U29728 (N_29728,N_22846,N_20791);
and U29729 (N_29729,N_24921,N_21080);
and U29730 (N_29730,N_20770,N_22652);
and U29731 (N_29731,N_21594,N_21341);
nor U29732 (N_29732,N_24780,N_23295);
or U29733 (N_29733,N_21683,N_24194);
xnor U29734 (N_29734,N_21075,N_23635);
and U29735 (N_29735,N_22199,N_22271);
xnor U29736 (N_29736,N_20805,N_24652);
xnor U29737 (N_29737,N_24626,N_23390);
nor U29738 (N_29738,N_23853,N_23109);
and U29739 (N_29739,N_23754,N_21882);
nor U29740 (N_29740,N_24198,N_20728);
nor U29741 (N_29741,N_23558,N_23137);
xor U29742 (N_29742,N_23226,N_22086);
nand U29743 (N_29743,N_21547,N_22926);
and U29744 (N_29744,N_21110,N_22721);
or U29745 (N_29745,N_20752,N_21726);
nor U29746 (N_29746,N_22491,N_20851);
or U29747 (N_29747,N_21888,N_23185);
nand U29748 (N_29748,N_20257,N_21170);
and U29749 (N_29749,N_24487,N_20735);
nand U29750 (N_29750,N_22153,N_21809);
nor U29751 (N_29751,N_23294,N_22248);
and U29752 (N_29752,N_23397,N_21374);
nand U29753 (N_29753,N_20099,N_20888);
nor U29754 (N_29754,N_21473,N_24099);
nand U29755 (N_29755,N_23622,N_23108);
or U29756 (N_29756,N_20482,N_20386);
or U29757 (N_29757,N_24698,N_24362);
nor U29758 (N_29758,N_22171,N_24901);
or U29759 (N_29759,N_20030,N_24534);
nor U29760 (N_29760,N_22567,N_21200);
and U29761 (N_29761,N_23388,N_21035);
or U29762 (N_29762,N_20998,N_21002);
xor U29763 (N_29763,N_24224,N_22653);
nor U29764 (N_29764,N_21111,N_23374);
nor U29765 (N_29765,N_22194,N_22938);
and U29766 (N_29766,N_22684,N_23061);
nor U29767 (N_29767,N_21960,N_23845);
nor U29768 (N_29768,N_21709,N_22478);
nand U29769 (N_29769,N_22945,N_24317);
and U29770 (N_29770,N_21105,N_20905);
nor U29771 (N_29771,N_20353,N_21946);
xor U29772 (N_29772,N_23527,N_22310);
or U29773 (N_29773,N_21642,N_21575);
nor U29774 (N_29774,N_24591,N_22192);
and U29775 (N_29775,N_21005,N_20080);
xnor U29776 (N_29776,N_23921,N_21658);
xor U29777 (N_29777,N_21055,N_21222);
nand U29778 (N_29778,N_23806,N_20584);
nor U29779 (N_29779,N_24431,N_20142);
or U29780 (N_29780,N_24241,N_22254);
nand U29781 (N_29781,N_24476,N_20296);
or U29782 (N_29782,N_24368,N_23697);
and U29783 (N_29783,N_21820,N_22645);
or U29784 (N_29784,N_24950,N_20092);
or U29785 (N_29785,N_21953,N_20005);
nand U29786 (N_29786,N_20680,N_24998);
or U29787 (N_29787,N_24620,N_20019);
xor U29788 (N_29788,N_20013,N_23815);
and U29789 (N_29789,N_24495,N_20933);
and U29790 (N_29790,N_20362,N_24674);
xor U29791 (N_29791,N_24868,N_20254);
xor U29792 (N_29792,N_20472,N_24184);
or U29793 (N_29793,N_21999,N_22425);
xnor U29794 (N_29794,N_23597,N_20253);
or U29795 (N_29795,N_24586,N_20694);
nor U29796 (N_29796,N_23116,N_22994);
and U29797 (N_29797,N_22391,N_22381);
nor U29798 (N_29798,N_21236,N_21090);
or U29799 (N_29799,N_24836,N_21034);
xor U29800 (N_29800,N_21024,N_20184);
xnor U29801 (N_29801,N_22303,N_24096);
and U29802 (N_29802,N_23495,N_23517);
nand U29803 (N_29803,N_24517,N_24436);
xor U29804 (N_29804,N_23569,N_21205);
nor U29805 (N_29805,N_23688,N_23552);
and U29806 (N_29806,N_23318,N_21703);
or U29807 (N_29807,N_20249,N_24614);
xnor U29808 (N_29808,N_21119,N_22810);
and U29809 (N_29809,N_23656,N_24251);
and U29810 (N_29810,N_24032,N_23915);
nor U29811 (N_29811,N_21627,N_23866);
nand U29812 (N_29812,N_21084,N_20262);
and U29813 (N_29813,N_24686,N_23033);
or U29814 (N_29814,N_24240,N_21351);
nor U29815 (N_29815,N_20884,N_22845);
nor U29816 (N_29816,N_22186,N_21459);
nand U29817 (N_29817,N_23309,N_23849);
or U29818 (N_29818,N_22851,N_24565);
or U29819 (N_29819,N_24763,N_23272);
or U29820 (N_29820,N_20618,N_22255);
and U29821 (N_29821,N_23955,N_20616);
nor U29822 (N_29822,N_23475,N_24765);
or U29823 (N_29823,N_21373,N_24963);
or U29824 (N_29824,N_20000,N_20290);
or U29825 (N_29825,N_20323,N_24280);
or U29826 (N_29826,N_21423,N_22565);
nor U29827 (N_29827,N_20312,N_21619);
or U29828 (N_29828,N_23150,N_22212);
nor U29829 (N_29829,N_24436,N_24129);
nand U29830 (N_29830,N_21475,N_21681);
xnor U29831 (N_29831,N_23410,N_21518);
xor U29832 (N_29832,N_22219,N_20973);
nor U29833 (N_29833,N_20736,N_21795);
and U29834 (N_29834,N_20665,N_22406);
nor U29835 (N_29835,N_21993,N_21609);
nand U29836 (N_29836,N_21992,N_22479);
xnor U29837 (N_29837,N_24965,N_24688);
nand U29838 (N_29838,N_21184,N_23732);
or U29839 (N_29839,N_23391,N_20339);
nor U29840 (N_29840,N_21624,N_20161);
nand U29841 (N_29841,N_21885,N_20194);
xnor U29842 (N_29842,N_20838,N_20904);
nor U29843 (N_29843,N_22671,N_21436);
and U29844 (N_29844,N_20066,N_23932);
nand U29845 (N_29845,N_24924,N_24126);
and U29846 (N_29846,N_21933,N_23976);
or U29847 (N_29847,N_20805,N_22726);
xor U29848 (N_29848,N_24365,N_24840);
nor U29849 (N_29849,N_23729,N_20634);
xor U29850 (N_29850,N_22007,N_22859);
xor U29851 (N_29851,N_21384,N_22013);
nor U29852 (N_29852,N_22762,N_21681);
nand U29853 (N_29853,N_20571,N_22644);
nand U29854 (N_29854,N_20252,N_20561);
nand U29855 (N_29855,N_22857,N_21909);
nor U29856 (N_29856,N_24690,N_24435);
nor U29857 (N_29857,N_20909,N_21636);
or U29858 (N_29858,N_22339,N_21357);
xnor U29859 (N_29859,N_23810,N_20069);
nand U29860 (N_29860,N_23210,N_23375);
and U29861 (N_29861,N_23021,N_20692);
nand U29862 (N_29862,N_21774,N_21042);
xnor U29863 (N_29863,N_22347,N_24425);
nor U29864 (N_29864,N_24316,N_24628);
nor U29865 (N_29865,N_22993,N_20517);
nor U29866 (N_29866,N_20614,N_24372);
or U29867 (N_29867,N_22317,N_22052);
xnor U29868 (N_29868,N_22403,N_20276);
xor U29869 (N_29869,N_20103,N_22489);
nor U29870 (N_29870,N_21211,N_21955);
nor U29871 (N_29871,N_21300,N_23506);
nand U29872 (N_29872,N_21554,N_23514);
or U29873 (N_29873,N_23959,N_23101);
and U29874 (N_29874,N_23932,N_20787);
and U29875 (N_29875,N_21444,N_22089);
xnor U29876 (N_29876,N_20493,N_24334);
xnor U29877 (N_29877,N_24458,N_21729);
or U29878 (N_29878,N_24267,N_20078);
nor U29879 (N_29879,N_24234,N_22891);
and U29880 (N_29880,N_20284,N_21970);
nor U29881 (N_29881,N_21096,N_20940);
nor U29882 (N_29882,N_23975,N_24685);
nor U29883 (N_29883,N_24218,N_22014);
or U29884 (N_29884,N_21709,N_22738);
nand U29885 (N_29885,N_23786,N_22183);
and U29886 (N_29886,N_23707,N_20506);
and U29887 (N_29887,N_24627,N_23555);
nand U29888 (N_29888,N_21838,N_20422);
or U29889 (N_29889,N_22297,N_23566);
nand U29890 (N_29890,N_23314,N_20253);
xor U29891 (N_29891,N_20072,N_22420);
or U29892 (N_29892,N_23537,N_20262);
or U29893 (N_29893,N_20465,N_23032);
xor U29894 (N_29894,N_22475,N_24118);
xor U29895 (N_29895,N_20597,N_23842);
or U29896 (N_29896,N_22638,N_22963);
or U29897 (N_29897,N_20772,N_22810);
or U29898 (N_29898,N_20588,N_21484);
xor U29899 (N_29899,N_24907,N_23724);
or U29900 (N_29900,N_22423,N_23519);
and U29901 (N_29901,N_21920,N_21328);
xor U29902 (N_29902,N_21274,N_20546);
and U29903 (N_29903,N_23974,N_24466);
or U29904 (N_29904,N_20652,N_20810);
nand U29905 (N_29905,N_21061,N_24062);
or U29906 (N_29906,N_22839,N_23214);
nor U29907 (N_29907,N_20856,N_23538);
or U29908 (N_29908,N_20065,N_21802);
or U29909 (N_29909,N_24996,N_24787);
xor U29910 (N_29910,N_23261,N_20934);
nand U29911 (N_29911,N_21584,N_20991);
nand U29912 (N_29912,N_22883,N_24915);
and U29913 (N_29913,N_20240,N_22143);
or U29914 (N_29914,N_21538,N_23783);
nor U29915 (N_29915,N_23881,N_24369);
xor U29916 (N_29916,N_24728,N_20976);
nand U29917 (N_29917,N_20378,N_21491);
or U29918 (N_29918,N_22277,N_24206);
xor U29919 (N_29919,N_20354,N_24071);
xor U29920 (N_29920,N_21697,N_20782);
nand U29921 (N_29921,N_20568,N_21648);
or U29922 (N_29922,N_22345,N_21449);
nand U29923 (N_29923,N_21008,N_22648);
or U29924 (N_29924,N_22274,N_22184);
nand U29925 (N_29925,N_21648,N_23348);
and U29926 (N_29926,N_20637,N_21394);
nor U29927 (N_29927,N_21070,N_22529);
nor U29928 (N_29928,N_23058,N_24532);
nor U29929 (N_29929,N_23887,N_21250);
nand U29930 (N_29930,N_23332,N_22834);
nor U29931 (N_29931,N_20154,N_24253);
nor U29932 (N_29932,N_20531,N_23548);
or U29933 (N_29933,N_24032,N_21974);
nand U29934 (N_29934,N_20146,N_21982);
nand U29935 (N_29935,N_20871,N_21047);
nor U29936 (N_29936,N_22721,N_24771);
nor U29937 (N_29937,N_24476,N_22751);
xor U29938 (N_29938,N_20111,N_24383);
nor U29939 (N_29939,N_22976,N_21029);
or U29940 (N_29940,N_22387,N_23052);
or U29941 (N_29941,N_23012,N_20892);
or U29942 (N_29942,N_22163,N_24704);
nand U29943 (N_29943,N_21516,N_22629);
and U29944 (N_29944,N_20187,N_22489);
nor U29945 (N_29945,N_21815,N_24173);
and U29946 (N_29946,N_20347,N_21485);
or U29947 (N_29947,N_23993,N_23700);
or U29948 (N_29948,N_20376,N_23718);
nor U29949 (N_29949,N_20278,N_24091);
or U29950 (N_29950,N_20059,N_20374);
nand U29951 (N_29951,N_22419,N_20868);
or U29952 (N_29952,N_22128,N_22847);
and U29953 (N_29953,N_20021,N_21646);
or U29954 (N_29954,N_24604,N_21997);
xor U29955 (N_29955,N_24478,N_23156);
and U29956 (N_29956,N_23437,N_24799);
or U29957 (N_29957,N_22598,N_24843);
xnor U29958 (N_29958,N_22301,N_20896);
nand U29959 (N_29959,N_21009,N_23666);
nor U29960 (N_29960,N_21890,N_24247);
nor U29961 (N_29961,N_24145,N_24344);
or U29962 (N_29962,N_22332,N_24343);
nand U29963 (N_29963,N_24218,N_24045);
nand U29964 (N_29964,N_22073,N_24075);
nand U29965 (N_29965,N_21419,N_20988);
nor U29966 (N_29966,N_22382,N_22931);
and U29967 (N_29967,N_20933,N_22354);
nand U29968 (N_29968,N_24907,N_22842);
nand U29969 (N_29969,N_20960,N_24643);
nor U29970 (N_29970,N_24741,N_21328);
nor U29971 (N_29971,N_23097,N_23476);
and U29972 (N_29972,N_21610,N_24448);
and U29973 (N_29973,N_24856,N_21043);
nand U29974 (N_29974,N_20141,N_24467);
or U29975 (N_29975,N_21125,N_21752);
and U29976 (N_29976,N_23772,N_23329);
or U29977 (N_29977,N_22315,N_22668);
and U29978 (N_29978,N_24191,N_20300);
nand U29979 (N_29979,N_23376,N_21935);
and U29980 (N_29980,N_20074,N_24997);
xnor U29981 (N_29981,N_21120,N_20662);
xor U29982 (N_29982,N_20991,N_20909);
nand U29983 (N_29983,N_23685,N_24791);
and U29984 (N_29984,N_20090,N_22245);
or U29985 (N_29985,N_20236,N_23007);
or U29986 (N_29986,N_23250,N_20193);
or U29987 (N_29987,N_23575,N_24298);
xor U29988 (N_29988,N_21265,N_24751);
and U29989 (N_29989,N_23604,N_20823);
or U29990 (N_29990,N_21997,N_21437);
nor U29991 (N_29991,N_21897,N_20391);
nand U29992 (N_29992,N_22234,N_23245);
nand U29993 (N_29993,N_20643,N_20126);
nor U29994 (N_29994,N_20406,N_24615);
and U29995 (N_29995,N_21556,N_22580);
nor U29996 (N_29996,N_21194,N_21738);
xnor U29997 (N_29997,N_24887,N_23666);
nand U29998 (N_29998,N_20404,N_23087);
and U29999 (N_29999,N_24712,N_22943);
xnor U30000 (N_30000,N_29332,N_28476);
and U30001 (N_30001,N_28194,N_25732);
and U30002 (N_30002,N_29531,N_29011);
or U30003 (N_30003,N_26483,N_26355);
nor U30004 (N_30004,N_26017,N_27066);
or U30005 (N_30005,N_29914,N_28157);
or U30006 (N_30006,N_25139,N_29862);
nor U30007 (N_30007,N_28585,N_25045);
or U30008 (N_30008,N_28793,N_26030);
xnor U30009 (N_30009,N_26124,N_28572);
nor U30010 (N_30010,N_28415,N_29805);
and U30011 (N_30011,N_27745,N_27634);
nor U30012 (N_30012,N_27923,N_27186);
xor U30013 (N_30013,N_25105,N_28436);
or U30014 (N_30014,N_29334,N_27029);
nor U30015 (N_30015,N_25231,N_26477);
nor U30016 (N_30016,N_26648,N_28899);
and U30017 (N_30017,N_27289,N_27319);
xnor U30018 (N_30018,N_28959,N_25903);
and U30019 (N_30019,N_29442,N_27939);
xnor U30020 (N_30020,N_29021,N_28792);
xnor U30021 (N_30021,N_29809,N_27181);
nor U30022 (N_30022,N_26877,N_26734);
nand U30023 (N_30023,N_27638,N_25845);
or U30024 (N_30024,N_28734,N_29698);
and U30025 (N_30025,N_29704,N_26994);
nor U30026 (N_30026,N_28231,N_25500);
and U30027 (N_30027,N_29070,N_28576);
and U30028 (N_30028,N_25747,N_27099);
xnor U30029 (N_30029,N_25919,N_28529);
and U30030 (N_30030,N_26963,N_26398);
nor U30031 (N_30031,N_29228,N_28803);
nor U30032 (N_30032,N_29926,N_27534);
xnor U30033 (N_30033,N_27320,N_28552);
and U30034 (N_30034,N_26338,N_25068);
nand U30035 (N_30035,N_28731,N_27052);
nand U30036 (N_30036,N_29633,N_29202);
and U30037 (N_30037,N_29373,N_29192);
xnor U30038 (N_30038,N_28080,N_29830);
xor U30039 (N_30039,N_26950,N_29231);
or U30040 (N_30040,N_25456,N_29340);
nand U30041 (N_30041,N_25171,N_29595);
and U30042 (N_30042,N_26039,N_29753);
nor U30043 (N_30043,N_28049,N_26695);
nor U30044 (N_30044,N_26104,N_26050);
nand U30045 (N_30045,N_25294,N_25061);
or U30046 (N_30046,N_26746,N_27844);
or U30047 (N_30047,N_29445,N_27587);
nand U30048 (N_30048,N_26100,N_26558);
or U30049 (N_30049,N_25965,N_25963);
and U30050 (N_30050,N_28314,N_29745);
or U30051 (N_30051,N_28862,N_29291);
or U30052 (N_30052,N_29648,N_29839);
or U30053 (N_30053,N_27911,N_25311);
and U30054 (N_30054,N_29514,N_26468);
xnor U30055 (N_30055,N_26774,N_28113);
or U30056 (N_30056,N_25084,N_26072);
or U30057 (N_30057,N_25388,N_26917);
and U30058 (N_30058,N_27197,N_26741);
nand U30059 (N_30059,N_29191,N_28325);
xnor U30060 (N_30060,N_28238,N_25148);
nand U30061 (N_30061,N_26564,N_26560);
and U30062 (N_30062,N_25938,N_28167);
or U30063 (N_30063,N_25077,N_25270);
nor U30064 (N_30064,N_25382,N_28624);
and U30065 (N_30065,N_28747,N_27619);
and U30066 (N_30066,N_29296,N_26952);
or U30067 (N_30067,N_27965,N_27170);
or U30068 (N_30068,N_27218,N_25094);
nand U30069 (N_30069,N_26207,N_29924);
nand U30070 (N_30070,N_28254,N_25447);
nand U30071 (N_30071,N_26766,N_28025);
xor U30072 (N_30072,N_28941,N_28383);
and U30073 (N_30073,N_25931,N_28685);
nor U30074 (N_30074,N_29016,N_25907);
nand U30075 (N_30075,N_25727,N_27018);
nor U30076 (N_30076,N_26377,N_29242);
and U30077 (N_30077,N_25947,N_27140);
nor U30078 (N_30078,N_27904,N_29229);
nor U30079 (N_30079,N_27726,N_29186);
and U30080 (N_30080,N_27035,N_25174);
xnor U30081 (N_30081,N_29087,N_27653);
nor U30082 (N_30082,N_28953,N_25768);
xnor U30083 (N_30083,N_29972,N_29183);
or U30084 (N_30084,N_26969,N_25295);
nor U30085 (N_30085,N_25650,N_29437);
xnor U30086 (N_30086,N_26902,N_28335);
nor U30087 (N_30087,N_29164,N_25746);
nor U30088 (N_30088,N_26624,N_26983);
or U30089 (N_30089,N_29925,N_25133);
nand U30090 (N_30090,N_29454,N_28195);
or U30091 (N_30091,N_26269,N_27135);
xnor U30092 (N_30092,N_27825,N_26496);
nor U30093 (N_30093,N_28183,N_27157);
and U30094 (N_30094,N_25262,N_29563);
nand U30095 (N_30095,N_25708,N_25423);
nand U30096 (N_30096,N_26553,N_27705);
xnor U30097 (N_30097,N_28896,N_27956);
or U30098 (N_30098,N_28962,N_25868);
nand U30099 (N_30099,N_26528,N_28506);
nor U30100 (N_30100,N_25553,N_27881);
nor U30101 (N_30101,N_29705,N_27327);
nand U30102 (N_30102,N_26710,N_28557);
nand U30103 (N_30103,N_28055,N_28575);
and U30104 (N_30104,N_28939,N_27623);
and U30105 (N_30105,N_26008,N_29835);
nand U30106 (N_30106,N_28091,N_26432);
nand U30107 (N_30107,N_28640,N_25943);
or U30108 (N_30108,N_29497,N_26006);
nor U30109 (N_30109,N_29324,N_29582);
nand U30110 (N_30110,N_29721,N_26526);
xnor U30111 (N_30111,N_28121,N_29451);
xnor U30112 (N_30112,N_29396,N_25352);
xor U30113 (N_30113,N_27301,N_29273);
xnor U30114 (N_30114,N_26972,N_27516);
nor U30115 (N_30115,N_25597,N_25327);
and U30116 (N_30116,N_26886,N_25433);
xnor U30117 (N_30117,N_25592,N_27611);
xnor U30118 (N_30118,N_26587,N_27642);
nand U30119 (N_30119,N_28701,N_25435);
or U30120 (N_30120,N_28785,N_27973);
and U30121 (N_30121,N_29712,N_27440);
xnor U30122 (N_30122,N_29979,N_28706);
nand U30123 (N_30123,N_26677,N_28606);
xor U30124 (N_30124,N_25624,N_26479);
xnor U30125 (N_30125,N_26307,N_29931);
or U30126 (N_30126,N_28587,N_26586);
and U30127 (N_30127,N_29892,N_27968);
nand U30128 (N_30128,N_25001,N_27699);
xor U30129 (N_30129,N_26942,N_27577);
or U30130 (N_30130,N_28482,N_28742);
nand U30131 (N_30131,N_27941,N_28942);
and U30132 (N_30132,N_29247,N_28020);
xnor U30133 (N_30133,N_27127,N_28367);
xnor U30134 (N_30134,N_28802,N_25242);
or U30135 (N_30135,N_28257,N_27455);
xor U30136 (N_30136,N_29064,N_25857);
nor U30137 (N_30137,N_28381,N_28819);
and U30138 (N_30138,N_28535,N_29529);
nand U30139 (N_30139,N_27171,N_26260);
and U30140 (N_30140,N_28635,N_25682);
nand U30141 (N_30141,N_26051,N_25793);
and U30142 (N_30142,N_29299,N_28344);
xnor U30143 (N_30143,N_26295,N_29626);
nand U30144 (N_30144,N_28727,N_29592);
and U30145 (N_30145,N_29995,N_27158);
nor U30146 (N_30146,N_28339,N_25124);
or U30147 (N_30147,N_25810,N_29300);
nor U30148 (N_30148,N_26612,N_28102);
nor U30149 (N_30149,N_26843,N_25924);
or U30150 (N_30150,N_26700,N_28908);
and U30151 (N_30151,N_26054,N_25802);
and U30152 (N_30152,N_28846,N_25059);
nor U30153 (N_30153,N_26473,N_26805);
xnor U30154 (N_30154,N_26725,N_28361);
and U30155 (N_30155,N_27692,N_26313);
and U30156 (N_30156,N_28117,N_26406);
and U30157 (N_30157,N_25686,N_28935);
or U30158 (N_30158,N_25959,N_29473);
and U30159 (N_30159,N_25414,N_28142);
or U30160 (N_30160,N_29967,N_26788);
nand U30161 (N_30161,N_28350,N_28919);
nor U30162 (N_30162,N_26064,N_25999);
nor U30163 (N_30163,N_28300,N_29621);
or U30164 (N_30164,N_28418,N_29657);
and U30165 (N_30165,N_25897,N_25318);
and U30166 (N_30166,N_28712,N_29692);
xnor U30167 (N_30167,N_25257,N_28777);
xnor U30168 (N_30168,N_28695,N_26012);
or U30169 (N_30169,N_25787,N_25770);
xnor U30170 (N_30170,N_25641,N_25291);
or U30171 (N_30171,N_27354,N_27445);
xor U30172 (N_30172,N_26209,N_29703);
nor U30173 (N_30173,N_27629,N_28402);
and U30174 (N_30174,N_26530,N_26484);
or U30175 (N_30175,N_26565,N_25154);
xnor U30176 (N_30176,N_25333,N_28312);
nor U30177 (N_30177,N_25712,N_25507);
xor U30178 (N_30178,N_28869,N_25426);
or U30179 (N_30179,N_28505,N_27925);
nor U30180 (N_30180,N_27994,N_27296);
and U30181 (N_30181,N_28541,N_29928);
nor U30182 (N_30182,N_29121,N_27818);
and U30183 (N_30183,N_27156,N_27584);
xnor U30184 (N_30184,N_27433,N_25410);
nor U30185 (N_30185,N_27441,N_26164);
nor U30186 (N_30186,N_29927,N_26614);
nor U30187 (N_30187,N_25019,N_28251);
and U30188 (N_30188,N_29655,N_25347);
and U30189 (N_30189,N_26491,N_25156);
xnor U30190 (N_30190,N_28276,N_26354);
or U30191 (N_30191,N_26544,N_29173);
nand U30192 (N_30192,N_27614,N_27085);
nand U30193 (N_30193,N_26711,N_27697);
nor U30194 (N_30194,N_26489,N_25620);
nor U30195 (N_30195,N_25518,N_26556);
nand U30196 (N_30196,N_28663,N_27276);
and U30197 (N_30197,N_25520,N_26997);
nor U30198 (N_30198,N_27672,N_26729);
and U30199 (N_30199,N_29863,N_29135);
xor U30200 (N_30200,N_26593,N_29249);
xnor U30201 (N_30201,N_25536,N_26380);
and U30202 (N_30202,N_29586,N_29735);
nand U30203 (N_30203,N_25767,N_26144);
nor U30204 (N_30204,N_29158,N_26539);
xnor U30205 (N_30205,N_25669,N_27793);
nand U30206 (N_30206,N_26792,N_27179);
xnor U30207 (N_30207,N_28061,N_28244);
nor U30208 (N_30208,N_28648,N_26719);
or U30209 (N_30209,N_25182,N_28448);
nor U30210 (N_30210,N_29329,N_29864);
or U30211 (N_30211,N_26933,N_27328);
nand U30212 (N_30212,N_26824,N_27631);
and U30213 (N_30213,N_29777,N_25250);
and U30214 (N_30214,N_28378,N_29195);
and U30215 (N_30215,N_25769,N_28444);
or U30216 (N_30216,N_26737,N_29620);
nand U30217 (N_30217,N_27252,N_26438);
nor U30218 (N_30218,N_28915,N_27717);
xor U30219 (N_30219,N_29938,N_26524);
nor U30220 (N_30220,N_29985,N_28387);
nand U30221 (N_30221,N_25086,N_25815);
and U30222 (N_30222,N_28767,N_27620);
xnor U30223 (N_30223,N_28211,N_29447);
nand U30224 (N_30224,N_28216,N_26718);
xnor U30225 (N_30225,N_29106,N_26186);
xnor U30226 (N_30226,N_29569,N_26178);
nor U30227 (N_30227,N_26841,N_26829);
nor U30228 (N_30228,N_28385,N_25934);
or U30229 (N_30229,N_28997,N_28374);
or U30230 (N_30230,N_27131,N_29312);
xor U30231 (N_30231,N_25535,N_26557);
xnor U30232 (N_30232,N_28769,N_28514);
nor U30233 (N_30233,N_25187,N_28096);
nand U30234 (N_30234,N_27972,N_27800);
and U30235 (N_30235,N_27601,N_27564);
nand U30236 (N_30236,N_28945,N_29916);
nor U30237 (N_30237,N_29872,N_27500);
or U30238 (N_30238,N_29096,N_28138);
xor U30239 (N_30239,N_25269,N_28203);
nor U30240 (N_30240,N_26617,N_27869);
nand U30241 (N_30241,N_25474,N_28399);
and U30242 (N_30242,N_26421,N_26762);
xnor U30243 (N_30243,N_26757,N_29791);
nor U30244 (N_30244,N_27287,N_25396);
xnor U30245 (N_30245,N_29711,N_25673);
or U30246 (N_30246,N_29891,N_25194);
nand U30247 (N_30247,N_28499,N_26937);
nor U30248 (N_30248,N_27801,N_26311);
xor U30249 (N_30249,N_28283,N_29257);
nor U30250 (N_30250,N_28468,N_26023);
and U30251 (N_30251,N_29554,N_29899);
nand U30252 (N_30252,N_26516,N_26031);
xor U30253 (N_30253,N_27123,N_27547);
or U30254 (N_30254,N_25288,N_28007);
and U30255 (N_30255,N_25973,N_27325);
nand U30256 (N_30256,N_28323,N_25853);
or U30257 (N_30257,N_25180,N_26964);
and U30258 (N_30258,N_27698,N_26328);
nand U30259 (N_30259,N_25796,N_28594);
xnor U30260 (N_30260,N_27443,N_26517);
or U30261 (N_30261,N_29510,N_25825);
and U30262 (N_30262,N_26267,N_25894);
nor U30263 (N_30263,N_25705,N_26702);
nor U30264 (N_30264,N_26263,N_28322);
nor U30265 (N_30265,N_26436,N_27989);
and U30266 (N_30266,N_29720,N_28353);
nand U30267 (N_30267,N_28311,N_26724);
nand U30268 (N_30268,N_29093,N_27714);
and U30269 (N_30269,N_26029,N_29198);
nand U30270 (N_30270,N_29271,N_27466);
xnor U30271 (N_30271,N_29025,N_26845);
or U30272 (N_30272,N_29117,N_26900);
nor U30273 (N_30273,N_28441,N_29264);
xor U30274 (N_30274,N_27036,N_27074);
or U30275 (N_30275,N_28437,N_28355);
or U30276 (N_30276,N_28303,N_29362);
nor U30277 (N_30277,N_26274,N_25877);
xnor U30278 (N_30278,N_25567,N_25995);
and U30279 (N_30279,N_27935,N_29277);
and U30280 (N_30280,N_27647,N_25029);
nor U30281 (N_30281,N_27876,N_25008);
or U30282 (N_30282,N_28934,N_25750);
nor U30283 (N_30283,N_25736,N_27020);
nand U30284 (N_30284,N_25632,N_25207);
nor U30285 (N_30285,N_29804,N_26992);
xnor U30286 (N_30286,N_27464,N_26063);
and U30287 (N_30287,N_29218,N_25030);
nand U30288 (N_30288,N_29983,N_27811);
nor U30289 (N_30289,N_27779,N_26576);
or U30290 (N_30290,N_29150,N_26674);
nand U30291 (N_30291,N_29499,N_26767);
xor U30292 (N_30292,N_26455,N_29343);
or U30293 (N_30293,N_27244,N_29841);
or U30294 (N_30294,N_29347,N_27583);
or U30295 (N_30295,N_27435,N_27612);
or U30296 (N_30296,N_26424,N_25366);
and U30297 (N_30297,N_28460,N_29583);
or U30298 (N_30298,N_26084,N_25885);
nor U30299 (N_30299,N_25883,N_26508);
nand U30300 (N_30300,N_27145,N_26894);
nor U30301 (N_30301,N_26794,N_26219);
nor U30302 (N_30302,N_25255,N_28109);
nand U30303 (N_30303,N_28659,N_27960);
or U30304 (N_30304,N_26704,N_27648);
nor U30305 (N_30305,N_25576,N_28574);
xor U30306 (N_30306,N_29762,N_29868);
nand U30307 (N_30307,N_26233,N_26132);
and U30308 (N_30308,N_28044,N_28008);
nor U30309 (N_30309,N_25007,N_28545);
nand U30310 (N_30310,N_25861,N_25609);
nor U30311 (N_30311,N_27804,N_25646);
xor U30312 (N_30312,N_29207,N_26641);
or U30313 (N_30313,N_28459,N_29115);
and U30314 (N_30314,N_29842,N_26388);
nand U30315 (N_30315,N_29047,N_27058);
nor U30316 (N_30316,N_28440,N_26381);
xor U30317 (N_30317,N_26128,N_25132);
and U30318 (N_30318,N_25819,N_29923);
or U30319 (N_30319,N_26465,N_29513);
nor U30320 (N_30320,N_25354,N_28174);
nand U30321 (N_30321,N_27755,N_25342);
xor U30322 (N_30322,N_26828,N_29425);
nand U30323 (N_30323,N_27909,N_27368);
nand U30324 (N_30324,N_27971,N_27662);
nor U30325 (N_30325,N_27429,N_27679);
xnor U30326 (N_30326,N_29538,N_25711);
nand U30327 (N_30327,N_26428,N_29256);
nand U30328 (N_30328,N_26172,N_27861);
nand U30329 (N_30329,N_27199,N_27856);
xor U30330 (N_30330,N_27588,N_27412);
xnor U30331 (N_30331,N_27567,N_25450);
or U30332 (N_30332,N_25582,N_25748);
xor U30333 (N_30333,N_27835,N_28450);
nand U30334 (N_30334,N_26303,N_29001);
xor U30335 (N_30335,N_25742,N_26601);
xor U30336 (N_30336,N_28295,N_29520);
or U30337 (N_30337,N_25698,N_28957);
nand U30338 (N_30338,N_29659,N_29145);
nand U30339 (N_30339,N_29859,N_25540);
nor U30340 (N_30340,N_28334,N_28029);
and U30341 (N_30341,N_26271,N_25461);
or U30342 (N_30342,N_27509,N_26745);
or U30343 (N_30343,N_26330,N_29706);
nor U30344 (N_30344,N_26515,N_29978);
xnor U30345 (N_30345,N_25689,N_29729);
and U30346 (N_30346,N_28419,N_25782);
and U30347 (N_30347,N_26159,N_29541);
nor U30348 (N_30348,N_28732,N_25982);
or U30349 (N_30349,N_26345,N_27084);
or U30350 (N_30350,N_25038,N_27905);
nor U30351 (N_30351,N_29843,N_25904);
and U30352 (N_30352,N_25674,N_28841);
xnor U30353 (N_30353,N_29873,N_26510);
or U30354 (N_30354,N_25716,N_26290);
and U30355 (N_30355,N_27845,N_28829);
and U30356 (N_30356,N_25521,N_26554);
xnor U30357 (N_30357,N_29128,N_28360);
or U30358 (N_30358,N_27855,N_25545);
xor U30359 (N_30359,N_27729,N_29302);
nor U30360 (N_30360,N_27091,N_27075);
and U30361 (N_30361,N_27312,N_28446);
xnor U30362 (N_30362,N_28682,N_26108);
and U30363 (N_30363,N_28876,N_29727);
xnor U30364 (N_30364,N_27759,N_27109);
xor U30365 (N_30365,N_26343,N_28817);
or U30366 (N_30366,N_25983,N_25072);
xnor U30367 (N_30367,N_29204,N_27880);
nand U30368 (N_30368,N_29308,N_25618);
nor U30369 (N_30369,N_28347,N_29602);
xnor U30370 (N_30370,N_27532,N_29895);
nor U30371 (N_30371,N_26226,N_27947);
nand U30372 (N_30372,N_29475,N_29686);
and U30373 (N_30373,N_28464,N_29053);
nand U30374 (N_30374,N_29966,N_29758);
and U30375 (N_30375,N_29774,N_28779);
nand U30376 (N_30376,N_25566,N_26385);
and U30377 (N_30377,N_29459,N_29635);
and U30378 (N_30378,N_27786,N_28521);
and U30379 (N_30379,N_26301,N_28001);
or U30380 (N_30380,N_28813,N_27465);
or U30381 (N_30381,N_29682,N_29759);
nand U30382 (N_30382,N_27832,N_27342);
xnor U30383 (N_30383,N_29787,N_26273);
nor U30384 (N_30384,N_29007,N_27038);
nor U30385 (N_30385,N_27051,N_28062);
nor U30386 (N_30386,N_25756,N_25699);
or U30387 (N_30387,N_26906,N_28252);
nor U30388 (N_30388,N_26005,N_29004);
xnor U30389 (N_30389,N_26364,N_29200);
or U30390 (N_30390,N_25169,N_26333);
nand U30391 (N_30391,N_26187,N_29063);
and U30392 (N_30392,N_26120,N_27754);
nand U30393 (N_30393,N_25277,N_26370);
and U30394 (N_30394,N_25106,N_27830);
and U30395 (N_30395,N_28234,N_29609);
nand U30396 (N_30396,N_26125,N_25981);
and U30397 (N_30397,N_26044,N_25593);
nand U30398 (N_30398,N_26324,N_25543);
nand U30399 (N_30399,N_29709,N_26189);
xnor U30400 (N_30400,N_25078,N_27859);
nor U30401 (N_30401,N_29060,N_25702);
and U30402 (N_30402,N_26412,N_29912);
or U30403 (N_30403,N_26856,N_28844);
or U30404 (N_30404,N_27434,N_27682);
xor U30405 (N_30405,N_29248,N_27457);
and U30406 (N_30406,N_29515,N_25490);
nand U30407 (N_30407,N_26019,N_27841);
nand U30408 (N_30408,N_28463,N_26591);
xnor U30409 (N_30409,N_26103,N_26811);
nor U30410 (N_30410,N_25737,N_29996);
nand U30411 (N_30411,N_27528,N_29412);
and U30412 (N_30412,N_25523,N_27995);
xnor U30413 (N_30413,N_28198,N_26860);
nand U30414 (N_30414,N_28038,N_29401);
nand U30415 (N_30415,N_28782,N_27579);
and U30416 (N_30416,N_27271,N_29293);
xor U30417 (N_30417,N_29405,N_27883);
or U30418 (N_30418,N_28160,N_26686);
nand U30419 (N_30419,N_26904,N_27599);
and U30420 (N_30420,N_26237,N_29687);
nor U30421 (N_30421,N_26649,N_29439);
nor U30422 (N_30422,N_27888,N_28032);
xnor U30423 (N_30423,N_27016,N_27826);
or U30424 (N_30424,N_26775,N_29095);
xor U30425 (N_30425,N_25577,N_29147);
and U30426 (N_30426,N_26141,N_28797);
nor U30427 (N_30427,N_28187,N_27749);
and U30428 (N_30428,N_26352,N_28166);
nor U30429 (N_30429,N_26098,N_27162);
xor U30430 (N_30430,N_25123,N_29527);
nor U30431 (N_30431,N_27982,N_28758);
nand U30432 (N_30432,N_27565,N_25684);
nor U30433 (N_30433,N_28559,N_27913);
or U30434 (N_30434,N_25253,N_25126);
and U30435 (N_30435,N_29304,N_25345);
nand U30436 (N_30436,N_29153,N_27760);
nor U30437 (N_30437,N_27794,N_29986);
and U30438 (N_30438,N_25188,N_26129);
xnor U30439 (N_30439,N_27828,N_25147);
nand U30440 (N_30440,N_27149,N_29301);
nor U30441 (N_30441,N_27380,N_25228);
and U30442 (N_30442,N_26447,N_28425);
and U30443 (N_30443,N_25704,N_27226);
or U30444 (N_30444,N_25120,N_27558);
or U30445 (N_30445,N_25402,N_27894);
and U30446 (N_30446,N_29723,N_26683);
nor U30447 (N_30447,N_28391,N_29642);
xnor U30448 (N_30448,N_25913,N_29309);
nor U30449 (N_30449,N_29888,N_28920);
and U30450 (N_30450,N_28968,N_27411);
or U30451 (N_30451,N_25879,N_27508);
nand U30452 (N_30452,N_25890,N_29988);
and U30453 (N_30453,N_28705,N_29666);
or U30454 (N_30454,N_26196,N_25751);
nand U30455 (N_30455,N_26135,N_25488);
xnor U30456 (N_30456,N_29270,N_27616);
nor U30457 (N_30457,N_27424,N_26032);
and U30458 (N_30458,N_29816,N_25780);
xor U30459 (N_30459,N_28787,N_25557);
nand U30460 (N_30460,N_27964,N_26344);
nand U30461 (N_30461,N_27555,N_25267);
nand U30462 (N_30462,N_25788,N_27180);
nand U30463 (N_30463,N_25168,N_26152);
nand U30464 (N_30464,N_25099,N_28313);
or U30465 (N_30465,N_28814,N_27257);
xnor U30466 (N_30466,N_29357,N_29665);
xnor U30467 (N_30467,N_27039,N_28465);
and U30468 (N_30468,N_28087,N_29356);
nor U30469 (N_30469,N_26948,N_27292);
or U30470 (N_30470,N_27379,N_29002);
or U30471 (N_30471,N_27061,N_27782);
xor U30472 (N_30472,N_27177,N_27645);
xor U30473 (N_30473,N_26208,N_26374);
nor U30474 (N_30474,N_26855,N_28615);
nor U30475 (N_30475,N_29321,N_27879);
and U30476 (N_30476,N_25263,N_25478);
xor U30477 (N_30477,N_27849,N_28280);
or U30478 (N_30478,N_29137,N_26882);
nor U30479 (N_30479,N_27491,N_27329);
and U30480 (N_30480,N_28726,N_26033);
or U30481 (N_30481,N_28201,N_29382);
and U30482 (N_30482,N_29913,N_29812);
xor U30483 (N_30483,N_25854,N_26583);
xor U30484 (N_30484,N_29619,N_26346);
and U30485 (N_30485,N_27143,N_28530);
xor U30486 (N_30486,N_29831,N_28879);
and U30487 (N_30487,N_29189,N_27545);
xnor U30488 (N_30488,N_25212,N_29311);
nor U30489 (N_30489,N_29870,N_28578);
nor U30490 (N_30490,N_28642,N_29084);
xnor U30491 (N_30491,N_28916,N_27453);
or U30492 (N_30492,N_28242,N_28644);
or U30493 (N_30493,N_25741,N_25541);
xor U30494 (N_30494,N_25390,N_25367);
or U30495 (N_30495,N_25547,N_25365);
and U30496 (N_30496,N_29467,N_26940);
or U30497 (N_30497,N_25492,N_25626);
nor U30498 (N_30498,N_25469,N_25297);
and U30499 (N_30499,N_27476,N_29607);
nor U30500 (N_30500,N_29533,N_27418);
or U30501 (N_30501,N_25595,N_28728);
nand U30502 (N_30502,N_28389,N_26859);
and U30503 (N_30503,N_29427,N_25745);
xnor U30504 (N_30504,N_26760,N_28564);
nand U30505 (N_30505,N_29756,N_27695);
and U30506 (N_30506,N_27696,N_28317);
nor U30507 (N_30507,N_28703,N_25240);
nor U30508 (N_30508,N_26234,N_28759);
xnor U30509 (N_30509,N_28825,N_29702);
nand U30510 (N_30510,N_26444,N_26761);
nor U30511 (N_30511,N_25697,N_28762);
or U30512 (N_30512,N_26314,N_28306);
xor U30513 (N_30513,N_25637,N_26679);
nor U30514 (N_30514,N_29157,N_28843);
nand U30515 (N_30515,N_25803,N_25146);
nor U30516 (N_30516,N_28004,N_27802);
xor U30517 (N_30517,N_26655,N_27920);
nand U30518 (N_30518,N_29904,N_28443);
or U30519 (N_30519,N_27966,N_25688);
and U30520 (N_30520,N_25118,N_28660);
and U30521 (N_30521,N_27395,N_28963);
xor U30522 (N_30522,N_27150,N_25628);
nand U30523 (N_30523,N_29165,N_28076);
and U30524 (N_30524,N_29568,N_25052);
xor U30525 (N_30525,N_26742,N_26357);
nand U30526 (N_30526,N_29601,N_28979);
or U30527 (N_30527,N_26013,N_28509);
and U30528 (N_30528,N_27919,N_26606);
nand U30529 (N_30529,N_27944,N_25792);
and U30530 (N_30530,N_29325,N_27137);
nand U30531 (N_30531,N_27813,N_25895);
nor U30532 (N_30532,N_26903,N_27420);
nand U30533 (N_30533,N_25383,N_25067);
nor U30534 (N_30534,N_25644,N_25887);
and U30535 (N_30535,N_27656,N_27912);
or U30536 (N_30536,N_26632,N_27931);
nor U30537 (N_30537,N_29650,N_28193);
nor U30538 (N_30538,N_25163,N_26699);
and U30539 (N_30539,N_29502,N_28667);
or U30540 (N_30540,N_27549,N_29422);
nor U30541 (N_30541,N_29457,N_28451);
and U30542 (N_30542,N_27111,N_28580);
and U30543 (N_30543,N_28152,N_28179);
nor U30544 (N_30544,N_27796,N_26779);
nor U30545 (N_30545,N_29654,N_27200);
nor U30546 (N_30546,N_29960,N_27267);
nand U30547 (N_30547,N_29822,N_29530);
or U30548 (N_30548,N_28743,N_25041);
nand U30549 (N_30549,N_29470,N_28154);
nor U30550 (N_30550,N_29180,N_27820);
nand U30551 (N_30551,N_25549,N_27928);
xnor U30552 (N_30552,N_28591,N_25872);
and U30553 (N_30553,N_29251,N_27142);
or U30554 (N_30554,N_26685,N_29739);
nor U30555 (N_30555,N_26002,N_28855);
xnor U30556 (N_30556,N_27169,N_28998);
and U30557 (N_30557,N_26839,N_28593);
nor U30558 (N_30558,N_25216,N_25477);
xnor U30559 (N_30559,N_27005,N_26383);
xor U30560 (N_30560,N_27812,N_25571);
nand U30561 (N_30561,N_29844,N_26361);
and U30562 (N_30562,N_28761,N_28128);
xnor U30563 (N_30563,N_28538,N_26981);
or U30564 (N_30564,N_29585,N_28611);
nand U30565 (N_30565,N_25213,N_28866);
or U30566 (N_30566,N_29974,N_27165);
or U30567 (N_30567,N_25744,N_27734);
nand U30568 (N_30568,N_26153,N_27363);
nor U30569 (N_30569,N_26472,N_27750);
xor U30570 (N_30570,N_27416,N_25016);
nand U30571 (N_30571,N_26763,N_29946);
or U30572 (N_30572,N_29213,N_26238);
or U30573 (N_30573,N_27961,N_28699);
and U30574 (N_30574,N_29867,N_28255);
or U30575 (N_30575,N_27206,N_27073);
nand U30576 (N_30576,N_29446,N_29837);
nor U30577 (N_30577,N_29464,N_25326);
or U30578 (N_30578,N_25125,N_29882);
nor U30579 (N_30579,N_25419,N_29989);
or U30580 (N_30580,N_26397,N_26636);
nor U30581 (N_30581,N_26927,N_26971);
xor U30582 (N_30582,N_26188,N_29539);
nand U30583 (N_30583,N_29193,N_29840);
xor U30584 (N_30584,N_25131,N_29005);
and U30585 (N_30585,N_29393,N_29107);
xnor U30586 (N_30586,N_26095,N_25457);
and U30587 (N_30587,N_29155,N_25489);
and U30588 (N_30588,N_29184,N_27377);
nor U30589 (N_30589,N_25584,N_26982);
or U30590 (N_30590,N_27580,N_25773);
and U30591 (N_30591,N_27447,N_27980);
nor U30592 (N_30592,N_25665,N_26861);
nand U30593 (N_30593,N_26025,N_29825);
and U30594 (N_30594,N_29632,N_29122);
and U30595 (N_30595,N_29677,N_29922);
and U30596 (N_30596,N_29900,N_28428);
nor U30597 (N_30597,N_28411,N_26411);
xnor U30598 (N_30598,N_29348,N_29715);
and U30599 (N_30599,N_29941,N_25760);
nor U30600 (N_30600,N_28895,N_27489);
xor U30601 (N_30601,N_25860,N_29801);
nand U30602 (N_30602,N_27034,N_28995);
or U30603 (N_30603,N_28345,N_25411);
or U30604 (N_30604,N_28133,N_27799);
and U30605 (N_30605,N_28485,N_28240);
xnor U30606 (N_30606,N_26671,N_25247);
nor U30607 (N_30607,N_27553,N_28687);
or U30608 (N_30608,N_28577,N_25925);
nand U30609 (N_30609,N_27637,N_28694);
and U30610 (N_30610,N_27151,N_26907);
xnor U30611 (N_30611,N_29546,N_29489);
nand U30612 (N_30612,N_27371,N_25300);
nand U30613 (N_30613,N_25918,N_29987);
xnor U30614 (N_30614,N_29567,N_26901);
and U30615 (N_30615,N_29736,N_29460);
xnor U30616 (N_30616,N_28292,N_26998);
nand U30617 (N_30617,N_29500,N_26895);
or U30618 (N_30618,N_29163,N_26905);
or U30619 (N_30619,N_27846,N_27272);
and U30620 (N_30620,N_25344,N_29280);
nor U30621 (N_30621,N_29639,N_25173);
nand U30622 (N_30622,N_26668,N_29557);
or U30623 (N_30623,N_26118,N_27358);
or U30624 (N_30624,N_28735,N_27521);
or U30625 (N_30625,N_28504,N_27356);
xor U30626 (N_30626,N_26797,N_28698);
nor U30627 (N_30627,N_25800,N_28217);
xor U30628 (N_30628,N_29765,N_28277);
and U30629 (N_30629,N_27011,N_28341);
xnor U30630 (N_30630,N_25685,N_28110);
or U30631 (N_30631,N_28164,N_26224);
or U30632 (N_30632,N_28188,N_27988);
nand U30633 (N_30633,N_27333,N_29779);
or U30634 (N_30634,N_28966,N_25946);
or U30635 (N_30635,N_28548,N_27929);
or U30636 (N_30636,N_29092,N_27615);
and U30637 (N_30637,N_25006,N_27556);
nor U30638 (N_30638,N_27068,N_28275);
nand U30639 (N_30639,N_26240,N_28205);
and U30640 (N_30640,N_27108,N_28471);
xnor U30641 (N_30641,N_29094,N_25606);
and U30642 (N_30642,N_26535,N_25984);
nor U30643 (N_30643,N_27872,N_29430);
xnor U30644 (N_30644,N_29059,N_26831);
nor U30645 (N_30645,N_25839,N_25088);
or U30646 (N_30646,N_26419,N_26470);
and U30647 (N_30647,N_25614,N_25048);
or U30648 (N_30648,N_25002,N_29934);
xnor U30649 (N_30649,N_26332,N_25372);
nand U30650 (N_30650,N_29043,N_29336);
or U30651 (N_30651,N_26995,N_27816);
nand U30652 (N_30652,N_28708,N_29866);
nor U30653 (N_30653,N_26551,N_29030);
or U30654 (N_30654,N_27847,N_27985);
nand U30655 (N_30655,N_29641,N_28219);
nor U30656 (N_30656,N_27317,N_25337);
nand U30657 (N_30657,N_28299,N_29486);
xnor U30658 (N_30658,N_28666,N_25151);
and U30659 (N_30659,N_25331,N_26572);
or U30660 (N_30660,N_29245,N_27336);
and U30661 (N_30661,N_29294,N_29333);
nand U30662 (N_30662,N_25590,N_28511);
or U30663 (N_30663,N_28668,N_27386);
or U30664 (N_30664,N_27625,N_25781);
nor U30665 (N_30665,N_25962,N_25233);
or U30666 (N_30666,N_28409,N_28643);
nor U30667 (N_30667,N_25987,N_25720);
nand U30668 (N_30668,N_25799,N_29181);
and U30669 (N_30669,N_29684,N_25676);
nor U30670 (N_30670,N_27047,N_29253);
and U30671 (N_30671,N_27590,N_26834);
and U30672 (N_30672,N_25412,N_26358);
xor U30673 (N_30673,N_29250,N_27212);
nor U30674 (N_30674,N_25511,N_25656);
nor U30675 (N_30675,N_26949,N_26951);
xnor U30676 (N_30676,N_25466,N_26190);
nand U30677 (N_30677,N_27807,N_29283);
and U30678 (N_30678,N_25908,N_25930);
and U30679 (N_30679,N_29477,N_28260);
nand U30680 (N_30680,N_26283,N_25399);
or U30681 (N_30681,N_27764,N_25141);
nand U30682 (N_30682,N_25643,N_28620);
and U30683 (N_30683,N_25954,N_27536);
nand U30684 (N_30684,N_28097,N_28253);
or U30685 (N_30685,N_25696,N_28487);
or U30686 (N_30686,N_28191,N_28297);
and U30687 (N_30687,N_29696,N_28554);
nand U30688 (N_30688,N_27027,N_28073);
or U30689 (N_30689,N_25243,N_26106);
or U30690 (N_30690,N_27144,N_26276);
or U30691 (N_30691,N_28078,N_29783);
or U30692 (N_30692,N_28500,N_26248);
xor U30693 (N_30693,N_27251,N_28362);
and U30694 (N_30694,N_27087,N_27242);
and U30695 (N_30695,N_29468,N_27249);
nor U30696 (N_30696,N_26778,N_28043);
nand U30697 (N_30697,N_26140,N_28247);
or U30698 (N_30698,N_28799,N_27851);
nor U30699 (N_30699,N_26401,N_26650);
or U30700 (N_30700,N_26921,N_28495);
xnor U30701 (N_30701,N_28661,N_28880);
nand U30702 (N_30702,N_28931,N_25276);
and U30703 (N_30703,N_29858,N_28290);
nand U30704 (N_30704,N_25301,N_27196);
xor U30705 (N_30705,N_29646,N_26168);
or U30706 (N_30706,N_26529,N_28664);
xor U30707 (N_30707,N_28481,N_29879);
nand U30708 (N_30708,N_28720,N_27562);
nor U30709 (N_30709,N_26936,N_26243);
nand U30710 (N_30710,N_25310,N_29824);
and U30711 (N_30711,N_25935,N_28881);
nand U30712 (N_30712,N_29320,N_25451);
nor U30713 (N_30713,N_26071,N_26356);
nor U30714 (N_30714,N_27809,N_25512);
and U30715 (N_30715,N_26522,N_29846);
xor U30716 (N_30716,N_29488,N_27046);
nand U30717 (N_30717,N_29918,N_26058);
xnor U30718 (N_30718,N_27787,N_29424);
nor U30719 (N_30719,N_28520,N_27795);
nor U30720 (N_30720,N_29950,N_29576);
or U30721 (N_30721,N_28823,N_28954);
and U30722 (N_30722,N_27167,N_25635);
nor U30723 (N_30723,N_27821,N_25942);
xnor U30724 (N_30724,N_28852,N_28691);
nor U30725 (N_30725,N_25258,N_26755);
xor U30726 (N_30726,N_27375,N_26403);
or U30727 (N_30727,N_27785,N_26490);
xnor U30728 (N_30728,N_28207,N_26869);
and U30729 (N_30729,N_28236,N_28479);
xor U30730 (N_30730,N_27054,N_27733);
xor U30731 (N_30731,N_25957,N_25612);
nor U30732 (N_30732,N_26111,N_25091);
nor U30733 (N_30733,N_27862,N_25526);
xor U30734 (N_30734,N_29932,N_29435);
nor U30735 (N_30735,N_25766,N_26386);
nor U30736 (N_30736,N_28909,N_27889);
nor U30737 (N_30737,N_28269,N_28438);
xor U30738 (N_30738,N_29061,N_28723);
or U30739 (N_30739,N_29484,N_28832);
and U30740 (N_30740,N_28549,N_29662);
xnor U30741 (N_30741,N_26059,N_27538);
and U30742 (N_30742,N_29605,N_25241);
nor U30743 (N_30743,N_29290,N_25065);
nor U30744 (N_30744,N_29588,N_27089);
nand U30745 (N_30745,N_26566,N_27550);
xnor U30746 (N_30746,N_26373,N_26418);
nor U30747 (N_30747,N_27768,N_26993);
xor U30748 (N_30748,N_28396,N_25401);
xnor U30749 (N_30749,N_27506,N_27891);
nand U30750 (N_30750,N_25558,N_29429);
or U30751 (N_30751,N_25098,N_28386);
nand U30752 (N_30752,N_29151,N_29883);
nand U30753 (N_30753,N_27792,N_26562);
and U30754 (N_30754,N_25814,N_28516);
nor U30755 (N_30755,N_28922,N_26919);
or U30756 (N_30756,N_26770,N_28861);
nand U30757 (N_30757,N_25322,N_25538);
xor U30758 (N_30758,N_27783,N_29337);
or U30759 (N_30759,N_27227,N_28757);
nor U30760 (N_30760,N_27680,N_25143);
nand U30761 (N_30761,N_28358,N_25274);
xnor U30762 (N_30762,N_26789,N_27594);
nand U30763 (N_30763,N_27351,N_25611);
or U30764 (N_30764,N_26815,N_28239);
nand U30765 (N_30765,N_25725,N_29136);
and U30766 (N_30766,N_25057,N_29113);
and U30767 (N_30767,N_29058,N_28359);
or U30768 (N_30768,N_28632,N_27667);
xor U30769 (N_30769,N_26842,N_26609);
xor U30770 (N_30770,N_29139,N_27348);
xnor U30771 (N_30771,N_28984,N_27529);
nand U30772 (N_30772,N_25260,N_26218);
xor U30773 (N_30773,N_26469,N_26220);
xnor U30774 (N_30774,N_25308,N_28744);
or U30775 (N_30775,N_29074,N_29593);
or U30776 (N_30776,N_27063,N_28938);
and U30777 (N_30777,N_29784,N_25285);
or U30778 (N_30778,N_25391,N_28037);
nand U30779 (N_30779,N_27322,N_29544);
nor U30780 (N_30780,N_28289,N_26507);
nand U30781 (N_30781,N_25970,N_26471);
nor U30782 (N_30782,N_27537,N_29610);
and U30783 (N_30783,N_28647,N_28563);
or U30784 (N_30784,N_27663,N_25647);
nand U30785 (N_30785,N_25384,N_28461);
and U30786 (N_30786,N_28204,N_29330);
or U30787 (N_30787,N_27539,N_27752);
nand U30788 (N_30788,N_26015,N_26256);
or U30789 (N_30789,N_29227,N_25040);
and U30790 (N_30790,N_25082,N_25755);
nor U30791 (N_30791,N_29980,N_25821);
nor U30792 (N_30792,N_27589,N_28738);
nand U30793 (N_30793,N_26962,N_28952);
xnor U30794 (N_30794,N_25884,N_25049);
or U30795 (N_30795,N_25893,N_28783);
and U30796 (N_30796,N_29476,N_26057);
xor U30797 (N_30797,N_27277,N_29263);
nand U30798 (N_30798,N_29323,N_26266);
or U30799 (N_30799,N_28512,N_29675);
and U30800 (N_30800,N_29645,N_28330);
and U30801 (N_30801,N_28950,N_29262);
nand U30802 (N_30802,N_25873,N_28400);
xnor U30803 (N_30803,N_27209,N_26546);
or U30804 (N_30804,N_29827,N_27670);
or U30805 (N_30805,N_28867,N_26004);
nor U30806 (N_30806,N_29553,N_29077);
and U30807 (N_30807,N_29776,N_27969);
or U30808 (N_30808,N_26083,N_28863);
and U30809 (N_30809,N_28151,N_26367);
or U30810 (N_30810,N_26221,N_26682);
or U30811 (N_30811,N_29808,N_29881);
xnor U30812 (N_30812,N_25976,N_29948);
nor U30813 (N_30813,N_26826,N_26193);
and U30814 (N_30814,N_25190,N_29085);
nor U30815 (N_30815,N_28775,N_27059);
nand U30816 (N_30816,N_28616,N_26748);
nor U30817 (N_30817,N_28937,N_28657);
nor U30818 (N_30818,N_28949,N_29496);
nand U30819 (N_30819,N_26000,N_29773);
nand U30820 (N_30820,N_26020,N_29999);
and U30821 (N_30821,N_27878,N_29608);
nor U30822 (N_30822,N_27299,N_28617);
nor U30823 (N_30823,N_26954,N_26646);
nor U30824 (N_30824,N_29860,N_29224);
nor U30825 (N_30825,N_27918,N_26434);
nand U30826 (N_30826,N_27139,N_25820);
nor U30827 (N_30827,N_27582,N_25204);
nand U30828 (N_30828,N_27668,N_26337);
and U30829 (N_30829,N_26410,N_29313);
nand U30830 (N_30830,N_29078,N_27469);
or U30831 (N_30831,N_26116,N_26200);
nand U30832 (N_30832,N_25949,N_27535);
or U30833 (N_30833,N_26532,N_29012);
nor U30834 (N_30834,N_27789,N_26804);
or U30835 (N_30835,N_29955,N_26450);
nand U30836 (N_30836,N_29511,N_25726);
or U30837 (N_30837,N_28424,N_29722);
nand U30838 (N_30838,N_27953,N_25044);
nor U30839 (N_30839,N_28902,N_26261);
or U30840 (N_30840,N_26924,N_29977);
and U30841 (N_30841,N_28357,N_25275);
nor U30842 (N_30842,N_29453,N_29419);
or U30843 (N_30843,N_29307,N_27391);
nand U30844 (N_30844,N_28181,N_29611);
and U30845 (N_30845,N_26932,N_25460);
and U30846 (N_30846,N_29219,N_26250);
and U30847 (N_30847,N_25636,N_28870);
and U30848 (N_30848,N_29614,N_25223);
nand U30849 (N_30849,N_28473,N_26010);
nand U30850 (N_30850,N_29921,N_25459);
xnor U30851 (N_30851,N_27732,N_26844);
and U30852 (N_30852,N_28014,N_26651);
nand U30853 (N_30853,N_27940,N_28103);
or U30854 (N_30854,N_26965,N_27124);
nor U30855 (N_30855,N_26980,N_26744);
and U30856 (N_30856,N_27661,N_26105);
or U30857 (N_30857,N_28679,N_26547);
nand U30858 (N_30858,N_28537,N_28082);
or U30859 (N_30859,N_29143,N_25373);
or U30860 (N_30860,N_29818,N_26185);
or U30861 (N_30861,N_26049,N_26520);
nand U30862 (N_30862,N_29742,N_28948);
xnor U30863 (N_30863,N_29149,N_27148);
xnor U30864 (N_30864,N_29288,N_28887);
xor U30865 (N_30865,N_29010,N_27414);
nand U30866 (N_30866,N_28918,N_28637);
nand U30867 (N_30867,N_26396,N_29823);
or U30868 (N_30868,N_29699,N_29524);
xor U30869 (N_30869,N_25565,N_26372);
xor U30870 (N_30870,N_26756,N_28136);
nor U30871 (N_30871,N_28980,N_27952);
or U30872 (N_30872,N_29017,N_26353);
nand U30873 (N_30873,N_28327,N_27086);
or U30874 (N_30874,N_25239,N_29190);
nand U30875 (N_30875,N_29057,N_26619);
nor U30876 (N_30876,N_29737,N_28089);
or U30877 (N_30877,N_25096,N_25428);
and U30878 (N_30878,N_29161,N_27417);
nand U30879 (N_30879,N_28993,N_29154);
and U30880 (N_30880,N_27510,N_25136);
nor U30881 (N_30881,N_29743,N_26166);
xnor U30882 (N_30882,N_27452,N_26109);
xnor U30883 (N_30883,N_29098,N_28375);
nand U30884 (N_30884,N_28689,N_29472);
and U30885 (N_30885,N_27613,N_28268);
nand U30886 (N_30886,N_28053,N_25855);
nand U30887 (N_30887,N_25293,N_26289);
nor U30888 (N_30888,N_29973,N_28992);
xnor U30889 (N_30889,N_25880,N_29141);
or U30890 (N_30890,N_26304,N_26423);
xor U30891 (N_30891,N_27644,N_27460);
and U30892 (N_30892,N_26934,N_26214);
nand U30893 (N_30893,N_26326,N_29024);
nor U30894 (N_30894,N_26688,N_28772);
or U30895 (N_30895,N_29266,N_26731);
nor U30896 (N_30896,N_28454,N_29055);
nor U30897 (N_30897,N_26620,N_25134);
nand U30898 (N_30898,N_29479,N_27188);
nor U30899 (N_30899,N_29730,N_28218);
or U30900 (N_30900,N_25679,N_29998);
nor U30901 (N_30901,N_25053,N_27404);
and U30902 (N_30902,N_25916,N_25831);
nor U30903 (N_30903,N_29306,N_25856);
nor U30904 (N_30904,N_25498,N_27850);
nand U30905 (N_30905,N_27049,N_29695);
or U30906 (N_30906,N_29885,N_25248);
nor U30907 (N_30907,N_28982,N_28965);
xnor U30908 (N_30908,N_25977,N_25119);
xnor U30909 (N_30909,N_27958,N_28688);
xor U30910 (N_30910,N_28083,N_29658);
nand U30911 (N_30911,N_27643,N_26038);
and U30912 (N_30912,N_26772,N_29088);
or U30913 (N_30913,N_26836,N_26603);
or U30914 (N_30914,N_26173,N_28108);
nor U30915 (N_30915,N_29731,N_25138);
and U30916 (N_30916,N_25031,N_25974);
xor U30917 (N_30917,N_26288,N_27933);
nor U30918 (N_30918,N_27178,N_25515);
nor U30919 (N_30919,N_27021,N_29381);
and U30920 (N_30920,N_26046,N_27007);
nand U30921 (N_30921,N_25302,N_26776);
nor U30922 (N_30922,N_25070,N_25579);
nand U30923 (N_30923,N_27974,N_29952);
xor U30924 (N_30924,N_25762,N_28702);
nor U30925 (N_30925,N_25771,N_26588);
or U30926 (N_30926,N_26268,N_28222);
nor U30927 (N_30927,N_25493,N_28501);
nor U30928 (N_30928,N_28776,N_27766);
and U30929 (N_30929,N_29399,N_29169);
or U30930 (N_30930,N_29945,N_27246);
xnor U30931 (N_30931,N_26060,N_27294);
or U30932 (N_30932,N_25012,N_27834);
or U30933 (N_30933,N_29140,N_25369);
or U30934 (N_30934,N_25621,N_27104);
or U30935 (N_30935,N_26360,N_27201);
nand U30936 (N_30936,N_25761,N_28649);
and U30937 (N_30937,N_29965,N_28366);
and U30938 (N_30938,N_28771,N_29214);
nor U30939 (N_30939,N_26968,N_25838);
or U30940 (N_30940,N_28175,N_27559);
nor U30941 (N_30941,N_28898,N_28302);
nand U30942 (N_30942,N_26308,N_28414);
xnor U30943 (N_30943,N_29901,N_27313);
xor U30944 (N_30944,N_26457,N_27773);
nand U30945 (N_30945,N_29778,N_27805);
nand U30946 (N_30946,N_28822,N_28447);
nor U30947 (N_30947,N_29993,N_27585);
or U30948 (N_30948,N_27718,N_26073);
nor U30949 (N_30949,N_28533,N_26707);
xnor U30950 (N_30950,N_28176,N_27959);
xor U30951 (N_30951,N_27874,N_25440);
or U30952 (N_30952,N_25629,N_28213);
nand U30953 (N_30953,N_26464,N_25491);
nor U30954 (N_30954,N_25953,N_28161);
and U30955 (N_30955,N_26052,N_26339);
or U30956 (N_30956,N_25881,N_29364);
xnor U30957 (N_30957,N_25738,N_27239);
nor U30958 (N_30958,N_29944,N_29376);
xnor U30959 (N_30959,N_29339,N_26525);
nand U30960 (N_30960,N_26325,N_26899);
and U30961 (N_30961,N_27134,N_26584);
and U30962 (N_30962,N_29767,N_26379);
nor U30963 (N_30963,N_28910,N_25554);
or U30964 (N_30964,N_26158,N_26085);
and U30965 (N_30965,N_26596,N_28077);
and U30966 (N_30966,N_29172,N_26228);
xnor U30967 (N_30967,N_27596,N_28741);
xnor U30968 (N_30968,N_25282,N_27230);
xor U30969 (N_30969,N_28655,N_29491);
nand U30970 (N_30970,N_28749,N_26368);
nand U30971 (N_30971,N_29465,N_26918);
and U30972 (N_30972,N_28069,N_27997);
xnor U30973 (N_30973,N_26175,N_28258);
nor U30974 (N_30974,N_29083,N_25950);
nand U30975 (N_30975,N_26908,N_25871);
or U30976 (N_30976,N_28592,N_26759);
nor U30977 (N_30977,N_25710,N_26456);
nand U30978 (N_30978,N_27210,N_29146);
nor U30979 (N_30979,N_29751,N_27349);
or U30980 (N_30980,N_26293,N_26148);
or U30981 (N_30981,N_26034,N_26732);
xnor U30982 (N_30982,N_26493,N_29953);
nor U30983 (N_30983,N_26941,N_27873);
nand U30984 (N_30984,N_27784,N_27771);
or U30985 (N_30985,N_29880,N_27942);
nor U30986 (N_30986,N_29690,N_28877);
nand U30987 (N_30987,N_28304,N_26872);
or U30988 (N_30988,N_26849,N_25851);
and U30989 (N_30989,N_28433,N_28673);
xor U30990 (N_30990,N_25922,N_29754);
xor U30991 (N_30991,N_27566,N_29469);
and U30992 (N_30992,N_27479,N_28671);
nand U30993 (N_30993,N_27530,N_29596);
or U30994 (N_30994,N_27254,N_29389);
nor U30995 (N_30995,N_28805,N_27525);
or U30996 (N_30996,N_28491,N_29409);
or U30997 (N_30997,N_28693,N_27427);
nor U30998 (N_30998,N_29981,N_26837);
xnor U30999 (N_30999,N_28141,N_26286);
and U31000 (N_31000,N_28232,N_29548);
nand U31001 (N_31001,N_29046,N_25218);
nand U31002 (N_31002,N_29579,N_26149);
nor U31003 (N_31003,N_25662,N_29281);
xor U31004 (N_31004,N_28890,N_25809);
nand U31005 (N_31005,N_25740,N_27999);
nand U31006 (N_31006,N_27266,N_25927);
nor U31007 (N_31007,N_28927,N_25778);
and U31008 (N_31008,N_26506,N_27161);
nor U31009 (N_31009,N_26703,N_29810);
nor U31010 (N_31010,N_28406,N_26117);
or U31011 (N_31011,N_27331,N_25037);
xnor U31012 (N_31012,N_27078,N_27945);
nand U31013 (N_31013,N_28973,N_26798);
and U31014 (N_31014,N_28790,N_27632);
nand U31015 (N_31015,N_25329,N_26595);
nand U31016 (N_31016,N_29028,N_25920);
and U31017 (N_31017,N_26440,N_28212);
nor U31018 (N_31018,N_25797,N_27362);
nand U31019 (N_31019,N_29800,N_28010);
xor U31020 (N_31020,N_27211,N_26121);
or U31021 (N_31021,N_28609,N_29571);
nand U31022 (N_31022,N_25442,N_29062);
xnor U31023 (N_31023,N_27172,N_26387);
or U31024 (N_31024,N_29649,N_25936);
and U31025 (N_31025,N_25055,N_29898);
xnor U31026 (N_31026,N_25150,N_25385);
nand U31027 (N_31027,N_26167,N_26573);
nor U31028 (N_31028,N_25281,N_29045);
nor U31029 (N_31029,N_27189,N_28305);
xnor U31030 (N_31030,N_25539,N_27270);
nand U31031 (N_31031,N_28893,N_27822);
nand U31032 (N_31032,N_28773,N_27410);
and U31033 (N_31033,N_26577,N_27655);
or U31034 (N_31034,N_29636,N_27438);
nor U31035 (N_31035,N_27248,N_26296);
or U31036 (N_31036,N_26027,N_25166);
or U31037 (N_31037,N_27635,N_26399);
nor U31038 (N_31038,N_27790,N_27693);
nand U31039 (N_31039,N_26446,N_25734);
or U31040 (N_31040,N_26504,N_25501);
nand U31041 (N_31041,N_26204,N_26197);
or U31042 (N_31042,N_26176,N_28839);
nand U31043 (N_31043,N_28928,N_27191);
xor U31044 (N_31044,N_25574,N_27374);
nor U31045 (N_31045,N_29782,N_28859);
or U31046 (N_31046,N_26830,N_29305);
and U31047 (N_31047,N_25555,N_28434);
or U31048 (N_31048,N_25642,N_25866);
or U31049 (N_31049,N_28555,N_29772);
nand U31050 (N_31050,N_28143,N_25779);
nand U31051 (N_31051,N_28107,N_28721);
or U31052 (N_31052,N_26203,N_28542);
nand U31053 (N_31053,N_29363,N_25694);
nor U31054 (N_31054,N_27370,N_27990);
or U31055 (N_31055,N_27743,N_27934);
nor U31056 (N_31056,N_25160,N_28894);
and U31057 (N_31057,N_27776,N_26923);
nand U31058 (N_31058,N_25062,N_25162);
xnor U31059 (N_31059,N_27198,N_26885);
xor U31060 (N_31060,N_27761,N_29174);
nor U31061 (N_31061,N_27430,N_25208);
xnor U31062 (N_31062,N_27263,N_28271);
nor U31063 (N_31063,N_28189,N_28050);
or U31064 (N_31064,N_28508,N_25840);
nand U31065 (N_31065,N_29877,N_25852);
xnor U31066 (N_31066,N_28907,N_25254);
or U31067 (N_31067,N_25531,N_28281);
xor U31068 (N_31068,N_29957,N_28192);
nor U31069 (N_31069,N_25550,N_26542);
or U31070 (N_31070,N_25355,N_25013);
xnor U31071 (N_31071,N_25027,N_25655);
nand U31072 (N_31072,N_26626,N_29215);
nand U31073 (N_31073,N_26653,N_28565);
xor U31074 (N_31074,N_25184,N_25978);
or U31075 (N_31075,N_29785,N_28225);
nand U31076 (N_31076,N_29316,N_27012);
xor U31077 (N_31077,N_28639,N_29246);
and U31078 (N_31078,N_25397,N_26171);
or U31079 (N_31079,N_28809,N_27937);
or U31080 (N_31080,N_25060,N_26819);
and U31081 (N_31081,N_25937,N_26880);
and U31082 (N_31082,N_26018,N_27660);
or U31083 (N_31083,N_25170,N_27033);
xor U31084 (N_31084,N_29237,N_26024);
and U31085 (N_31085,N_25272,N_27593);
nand U31086 (N_31086,N_29072,N_26393);
and U31087 (N_31087,N_28602,N_26402);
and U31088 (N_31088,N_27076,N_26467);
nor U31089 (N_31089,N_29615,N_25654);
xnor U31090 (N_31090,N_27606,N_25505);
nor U31091 (N_31091,N_29235,N_27369);
xnor U31092 (N_31092,N_29075,N_29521);
nor U31093 (N_31093,N_25036,N_25446);
and U31094 (N_31094,N_26101,N_29188);
nand U31095 (N_31095,N_27657,N_27025);
xor U31096 (N_31096,N_28684,N_26292);
nor U31097 (N_31097,N_28531,N_26462);
nor U31098 (N_31098,N_25537,N_28475);
and U31099 (N_31099,N_27738,N_26747);
nor U31100 (N_31100,N_28221,N_29624);
nor U31101 (N_31101,N_25524,N_25387);
xnor U31102 (N_31102,N_27017,N_25142);
nor U31103 (N_31103,N_27205,N_27977);
xnor U31104 (N_31104,N_27646,N_28622);
nand U31105 (N_31105,N_25018,N_26056);
nor U31106 (N_31106,N_25966,N_25955);
nand U31107 (N_31107,N_27602,N_29480);
nand U31108 (N_31108,N_27915,N_25824);
nor U31109 (N_31109,N_28099,N_27691);
and U31110 (N_31110,N_28124,N_26946);
or U31111 (N_31111,N_27808,N_26987);
xnor U31112 (N_31112,N_29507,N_25530);
nor U31113 (N_31113,N_28364,N_26521);
and U31114 (N_31114,N_27105,N_29573);
xnor U31115 (N_31115,N_28127,N_29958);
nand U31116 (N_31116,N_29503,N_27507);
xor U31117 (N_31117,N_27719,N_27604);
and U31118 (N_31118,N_25339,N_29871);
nor U31119 (N_31119,N_28618,N_28036);
and U31120 (N_31120,N_28285,N_28336);
nor U31121 (N_31121,N_27957,N_25014);
and U31122 (N_31122,N_25680,N_26977);
nor U31123 (N_31123,N_26984,N_29564);
or U31124 (N_31124,N_29565,N_28298);
xnor U31125 (N_31125,N_26713,N_28518);
or U31126 (N_31126,N_27857,N_28282);
xnor U31127 (N_31127,N_28256,N_25801);
xnor U31128 (N_31128,N_26863,N_26916);
nand U31129 (N_31129,N_28370,N_28393);
and U31130 (N_31130,N_26911,N_25201);
nor U31131 (N_31131,N_26850,N_25217);
xor U31132 (N_31132,N_25836,N_28135);
nand U31133 (N_31133,N_25508,N_27684);
or U31134 (N_31134,N_25968,N_25357);
and U31135 (N_31135,N_26832,N_28229);
nand U31136 (N_31136,N_27392,N_29814);
xor U31137 (N_31137,N_27232,N_27877);
and U31138 (N_31138,N_26068,N_25534);
xnor U31139 (N_31139,N_25487,N_26953);
and U31140 (N_31140,N_27595,N_27385);
and U31141 (N_31141,N_29355,N_26316);
or U31142 (N_31142,N_25497,N_25404);
xnor U31143 (N_31143,N_26482,N_25717);
and U31144 (N_31144,N_27444,N_28864);
nor U31145 (N_31145,N_25774,N_25325);
nand U31146 (N_31146,N_28057,N_27473);
and U31147 (N_31147,N_25227,N_29598);
nor U31148 (N_31148,N_29732,N_26442);
and U31149 (N_31149,N_27238,N_28155);
and U31150 (N_31150,N_27557,N_27708);
or U31151 (N_31151,N_27182,N_27658);
nor U31152 (N_31152,N_27128,N_28380);
xnor U31153 (N_31153,N_28196,N_28621);
and U31154 (N_31154,N_27069,N_26569);
and U31155 (N_31155,N_28426,N_27450);
nand U31156 (N_31156,N_26279,N_26555);
nand U31157 (N_31157,N_27518,N_25519);
and U31158 (N_31158,N_25653,N_27748);
nor U31159 (N_31159,N_26138,N_27902);
nand U31160 (N_31160,N_25896,N_29710);
nor U31161 (N_31161,N_29217,N_26644);
xor U31162 (N_31162,N_27863,N_29081);
xnor U31163 (N_31163,N_27159,N_29388);
xor U31164 (N_31164,N_27384,N_26509);
nor U31165 (N_31165,N_26165,N_26822);
and U31166 (N_31166,N_29428,N_26957);
or U31167 (N_31167,N_25721,N_28106);
xor U31168 (N_31168,N_28153,N_29509);
nor U31169 (N_31169,N_26405,N_28882);
or U31170 (N_31170,N_28146,N_28745);
xnor U31171 (N_31171,N_27618,N_25116);
or U31172 (N_31172,N_29082,N_29752);
nand U31173 (N_31173,N_26910,N_28470);
or U31174 (N_31174,N_27381,N_25651);
or U31175 (N_31175,N_29505,N_28833);
and U31176 (N_31176,N_29850,N_27753);
and U31177 (N_31177,N_29051,N_25586);
xnor U31178 (N_31178,N_26673,N_29688);
nor U31179 (N_31179,N_28478,N_25476);
xnor U31180 (N_31180,N_25998,N_26790);
or U31181 (N_31181,N_25613,N_29105);
and U31182 (N_31182,N_27302,N_26808);
nor U31183 (N_31183,N_26865,N_28856);
and U31184 (N_31184,N_27399,N_25775);
nor U31185 (N_31185,N_26112,N_25284);
or U31186 (N_31186,N_29915,N_26272);
or U31187 (N_31187,N_25080,N_27352);
or U31188 (N_31188,N_26803,N_25657);
xnor U31189 (N_31189,N_29048,N_26284);
xor U31190 (N_31190,N_25429,N_27810);
nand U31191 (N_31191,N_28697,N_27081);
or U31192 (N_31192,N_26966,N_29540);
or U31193 (N_31193,N_27298,N_25706);
or U31194 (N_31194,N_29550,N_29994);
nor U31195 (N_31195,N_27814,N_26821);
nor U31196 (N_31196,N_28369,N_25332);
or U31197 (N_31197,N_28801,N_28318);
nor U31198 (N_31198,N_26570,N_29240);
nor U31199 (N_31199,N_26676,N_27998);
xor U31200 (N_31200,N_26048,N_26007);
and U31201 (N_31201,N_29448,N_25728);
or U31202 (N_31202,N_26478,N_25479);
or U31203 (N_31203,N_27906,N_25035);
nor U31204 (N_31204,N_28670,N_27119);
nand U31205 (N_31205,N_26503,N_26961);
and U31206 (N_31206,N_26958,N_26257);
nand U31207 (N_31207,N_28392,N_25448);
or U31208 (N_31208,N_29561,N_29350);
nand U31209 (N_31209,N_29594,N_29845);
or U31210 (N_31210,N_27630,N_28770);
or U31211 (N_31211,N_27831,N_26868);
nand U31212 (N_31212,N_26502,N_26730);
nand U31213 (N_31213,N_28519,N_25348);
xnor U31214 (N_31214,N_26009,N_27442);
and U31215 (N_31215,N_25324,N_25486);
nand U31216 (N_31216,N_29331,N_29878);
and U31217 (N_31217,N_25874,N_27916);
xnor U31218 (N_31218,N_27848,N_27951);
and U31219 (N_31219,N_25729,N_26669);
nor U31220 (N_31220,N_28394,N_29449);
nor U31221 (N_31221,N_25630,N_29265);
and U31222 (N_31222,N_27865,N_27118);
nand U31223 (N_31223,N_25359,N_28571);
nand U31224 (N_31224,N_27229,N_26752);
xnor U31225 (N_31225,N_29390,N_26139);
xor U31226 (N_31226,N_28892,N_25765);
or U31227 (N_31227,N_29861,N_25572);
nand U31228 (N_31228,N_27777,N_25485);
or U31229 (N_31229,N_26801,N_29090);
nand U31230 (N_31230,N_28607,N_29407);
nor U31231 (N_31231,N_29345,N_26974);
or U31232 (N_31232,N_28794,N_25028);
or U31233 (N_31233,N_25958,N_29875);
xnor U31234 (N_31234,N_26391,N_26154);
and U31235 (N_31235,N_27284,N_25832);
nor U31236 (N_31236,N_28768,N_26162);
and U31237 (N_31237,N_29628,N_26945);
xnor U31238 (N_31238,N_29420,N_26067);
and U31239 (N_31239,N_29797,N_27640);
nor U31240 (N_31240,N_28676,N_26433);
or U31241 (N_31241,N_29326,N_28717);
and U31242 (N_31242,N_26817,N_26881);
and U31243 (N_31243,N_25432,N_27092);
nor U31244 (N_31244,N_29728,N_27346);
or U31245 (N_31245,N_28139,N_29014);
nand U31246 (N_31246,N_27295,N_27575);
and U31247 (N_31247,N_28940,N_29315);
nor U31248 (N_31248,N_25152,N_29936);
and U31249 (N_31249,N_28791,N_25266);
and U31250 (N_31250,N_27949,N_25316);
or U31251 (N_31251,N_28975,N_28714);
nor U31252 (N_31252,N_26114,N_29209);
xnor U31253 (N_31253,N_29485,N_28854);
and U31254 (N_31254,N_29604,N_25183);
nand U31255 (N_31255,N_27285,N_26523);
nor U31256 (N_31256,N_25677,N_25914);
and U31257 (N_31257,N_27671,N_27048);
and U31258 (N_31258,N_25875,N_28051);
nor U31259 (N_31259,N_28796,N_27110);
xor U31260 (N_31260,N_28543,N_27026);
nand U31261 (N_31261,N_28926,N_26764);
nor U31262 (N_31262,N_28376,N_29258);
nor U31263 (N_31263,N_26889,N_29990);
xnor U31264 (N_31264,N_28308,N_28065);
nor U31265 (N_31265,N_29226,N_29853);
nand U31266 (N_31266,N_28005,N_25026);
xor U31267 (N_31267,N_26897,N_28006);
nand U31268 (N_31268,N_25784,N_29275);
or U31269 (N_31269,N_25023,N_26785);
and U31270 (N_31270,N_25252,N_28112);
xor U31271 (N_31271,N_28798,N_25602);
and U31272 (N_31272,N_28079,N_27674);
nand U31273 (N_31273,N_26113,N_26864);
nand U31274 (N_31274,N_29225,N_29371);
and U31275 (N_31275,N_25473,N_26970);
or U31276 (N_31276,N_28093,N_29618);
nand U31277 (N_31277,N_27459,N_26610);
nand U31278 (N_31278,N_25425,N_28999);
or U31279 (N_31279,N_26749,N_25594);
nand U31280 (N_31280,N_25847,N_25064);
and U31281 (N_31281,N_29959,N_27300);
or U31282 (N_31282,N_26110,N_29627);
nor U31283 (N_31283,N_27910,N_25236);
nand U31284 (N_31284,N_26390,N_29118);
or U31285 (N_31285,N_29232,N_29656);
nor U31286 (N_31286,N_27742,N_29456);
xnor U31287 (N_31287,N_27372,N_29156);
nor U31288 (N_31288,N_27394,N_28484);
and U31289 (N_31289,N_27053,N_26896);
xor U31290 (N_31290,N_29634,N_26458);
nand U31291 (N_31291,N_25376,N_25374);
nor U31292 (N_31292,N_27315,N_26690);
and U31293 (N_31293,N_26739,N_28122);
xnor U31294 (N_31294,N_25996,N_26568);
and U31295 (N_31295,N_28748,N_28646);
or U31296 (N_31296,N_29124,N_25575);
nor U31297 (N_31297,N_29631,N_26378);
xnor U31298 (N_31298,N_29268,N_28737);
xnor U31299 (N_31299,N_25865,N_29441);
and U31300 (N_31300,N_28031,N_27273);
and U31301 (N_31301,N_29116,N_25424);
nand U31302 (N_31302,N_27155,N_28596);
nor U31303 (N_31303,N_27681,N_25910);
or U31304 (N_31304,N_26893,N_25438);
or U31305 (N_31305,N_25341,N_29889);
nand U31306 (N_31306,N_29668,N_29194);
nand U31307 (N_31307,N_28058,N_25022);
nand U31308 (N_31308,N_29876,N_25573);
or U31309 (N_31309,N_29386,N_29671);
or U31310 (N_31310,N_29259,N_26835);
nor U31311 (N_31311,N_26407,N_26198);
xnor U31312 (N_31312,N_28835,N_29466);
and U31313 (N_31313,N_28913,N_25463);
nor U31314 (N_31314,N_28766,N_25668);
and U31315 (N_31315,N_26210,N_26206);
nor U31316 (N_31316,N_26161,N_27291);
nand U31317 (N_31317,N_27817,N_25480);
xor U31318 (N_31318,N_29854,N_26930);
or U31319 (N_31319,N_27574,N_27183);
nor U31320 (N_31320,N_28725,N_29295);
or U31321 (N_31321,N_28826,N_26363);
or U31322 (N_31322,N_25063,N_29747);
and U31323 (N_31323,N_25159,N_26852);
or U31324 (N_31324,N_29884,N_25172);
nor U31325 (N_31325,N_27339,N_29111);
nand U31326 (N_31326,N_26635,N_29205);
or U31327 (N_31327,N_28597,N_28830);
or U31328 (N_31328,N_29580,N_25164);
nand U31329 (N_31329,N_25533,N_25826);
nor U31330 (N_31330,N_27501,N_25024);
nor U31331 (N_31331,N_29284,N_28733);
and U31332 (N_31332,N_28352,N_25828);
nand U31333 (N_31333,N_25046,N_26922);
or U31334 (N_31334,N_26229,N_27064);
and U31335 (N_31335,N_26365,N_27274);
nor U31336 (N_31336,N_28818,N_29292);
nand U31337 (N_31337,N_26631,N_28439);
nor U31338 (N_31338,N_26656,N_25113);
or U31339 (N_31339,N_27827,N_29397);
xor U31340 (N_31340,N_29897,N_26235);
nor U31341 (N_31341,N_27767,N_25244);
xor U31342 (N_31342,N_29673,N_25011);
nor U31343 (N_31343,N_26715,N_26873);
and U31344 (N_31344,N_25230,N_28811);
nor U31345 (N_31345,N_29968,N_25952);
nand U31346 (N_31346,N_28115,N_26016);
and U31347 (N_31347,N_26317,N_29643);
or U31348 (N_31348,N_27515,N_28296);
and U31349 (N_31349,N_26319,N_28180);
or U31350 (N_31350,N_26781,N_29803);
xor U31351 (N_31351,N_28522,N_26488);
and U31352 (N_31352,N_28009,N_25198);
nand U31353 (N_31353,N_28781,N_26422);
nand U31354 (N_31354,N_29385,N_25988);
nand U31355 (N_31355,N_28126,N_27364);
nor U31356 (N_31356,N_27603,N_26675);
xor U31357 (N_31357,N_27174,N_27723);
and U31358 (N_31358,N_28163,N_29310);
xor U31359 (N_31359,N_29338,N_27687);
nor U31360 (N_31360,N_28850,N_28332);
nor U31361 (N_31361,N_29734,N_26306);
nor U31362 (N_31362,N_25189,N_28990);
or U31363 (N_31363,N_28806,N_26131);
nand U31364 (N_31364,N_28429,N_27927);
xor U31365 (N_31365,N_28363,N_25221);
nand U31366 (N_31366,N_27715,N_27000);
nand U31367 (N_31367,N_28947,N_26145);
or U31368 (N_31368,N_27495,N_26126);
nand U31369 (N_31369,N_26409,N_26578);
nand U31370 (N_31370,N_25054,N_28384);
nor U31371 (N_31371,N_25251,N_28410);
and U31372 (N_31372,N_28235,N_25956);
nand U31373 (N_31373,N_26533,N_29052);
nor U31374 (N_31374,N_28488,N_26545);
or U31375 (N_31375,N_25975,N_29110);
or U31376 (N_31376,N_26169,N_28489);
nand U31377 (N_31377,N_27838,N_25017);
xor U31378 (N_31378,N_28458,N_29741);
nor U31379 (N_31379,N_28286,N_27639);
and U31380 (N_31380,N_28605,N_27884);
xnor U31381 (N_31381,N_26765,N_27788);
nor U31382 (N_31382,N_29663,N_29152);
and U31383 (N_31383,N_28696,N_25972);
and U31384 (N_31384,N_28490,N_28209);
xor U31385 (N_31385,N_29170,N_29781);
and U31386 (N_31386,N_26331,N_29365);
nand U31387 (N_31387,N_28333,N_29719);
nand U31388 (N_31388,N_29120,N_27703);
xor U31389 (N_31389,N_27350,N_27781);
or U31390 (N_31390,N_27001,N_27527);
or U31391 (N_31391,N_27402,N_25743);
xor U31392 (N_31392,N_25232,N_27586);
or U31393 (N_31393,N_28838,N_28739);
or U31394 (N_31394,N_25103,N_25661);
and U31395 (N_31395,N_29910,N_25034);
and U31396 (N_31396,N_29584,N_25405);
nor U31397 (N_31397,N_29276,N_28272);
or U31398 (N_31398,N_25351,N_27673);
nand U31399 (N_31399,N_26672,N_28033);
or U31400 (N_31400,N_25101,N_28397);
and U31401 (N_31401,N_29764,N_27095);
nor U31402 (N_31402,N_26461,N_27730);
xnor U31403 (N_31403,N_27936,N_26142);
or U31404 (N_31404,N_28837,N_29707);
xor U31405 (N_31405,N_25776,N_28413);
nand U31406 (N_31406,N_27478,N_29947);
or U31407 (N_31407,N_26041,N_28650);
nor U31408 (N_31408,N_28951,N_25718);
or U31409 (N_31409,N_27735,N_26633);
xnor U31410 (N_31410,N_27367,N_28547);
nand U31411 (N_31411,N_25502,N_27383);
nor U31412 (N_31412,N_25583,N_29050);
nor U31413 (N_31413,N_29893,N_27269);
xor U31414 (N_31414,N_26687,N_27725);
xor U31415 (N_31415,N_28828,N_25564);
nand U31416 (N_31416,N_25882,N_27898);
nand U31417 (N_31417,N_26252,N_27423);
or U31418 (N_31418,N_28170,N_25757);
and U31419 (N_31419,N_25596,N_27240);
xor U31420 (N_31420,N_25074,N_29022);
nor U31421 (N_31421,N_27930,N_28638);
or U31422 (N_31422,N_29572,N_25361);
nand U31423 (N_31423,N_25196,N_25004);
xnor U31424 (N_31424,N_28331,N_29894);
and U31425 (N_31425,N_28348,N_29112);
nor U31426 (N_31426,N_25178,N_25349);
nand U31427 (N_31427,N_25033,N_28502);
or U31428 (N_31428,N_26985,N_28634);
xnor U31429 (N_31429,N_26035,N_27720);
or U31430 (N_31430,N_27676,N_29244);
nand U31431 (N_31431,N_28569,N_28435);
or U31432 (N_31432,N_27899,N_29716);
xnor U31433 (N_31433,N_25199,N_25109);
and U31434 (N_31434,N_28068,N_27224);
nand U31435 (N_31435,N_28858,N_25986);
nor U31436 (N_31436,N_26155,N_25193);
nand U31437 (N_31437,N_28765,N_28996);
xor U31438 (N_31438,N_26717,N_25229);
nand U31439 (N_31439,N_29606,N_27288);
and U31440 (N_31440,N_26914,N_25806);
or U31441 (N_31441,N_27102,N_25867);
xor U31442 (N_31442,N_28150,N_29917);
nand U31443 (N_31443,N_27065,N_28656);
nor U31444 (N_31444,N_29462,N_26181);
and U31445 (N_31445,N_26943,N_27842);
nor U31446 (N_31446,N_28064,N_29423);
xnor U31447 (N_31447,N_27694,N_29613);
xnor U31448 (N_31448,N_26001,N_25130);
nor U31449 (N_31449,N_28472,N_27505);
or U31450 (N_31450,N_29820,N_26174);
xnor U31451 (N_31451,N_26627,N_29108);
nor U31452 (N_31452,N_26847,N_26512);
and U31453 (N_31453,N_25627,N_25107);
nand U31454 (N_31454,N_26750,N_26630);
xnor U31455 (N_31455,N_25923,N_26429);
or U31456 (N_31456,N_26691,N_26920);
and U31457 (N_31457,N_26939,N_29971);
and U31458 (N_31458,N_28831,N_27114);
nand U31459 (N_31459,N_25483,N_29746);
and U31460 (N_31460,N_27649,N_28763);
nand U31461 (N_31461,N_28755,N_28753);
nor U31462 (N_31462,N_28224,N_28483);
nand U31463 (N_31463,N_25844,N_28729);
xor U31464 (N_31464,N_28989,N_26334);
and U31465 (N_31465,N_29103,N_27758);
or U31466 (N_31466,N_28377,N_25849);
xnor U31467 (N_31467,N_27303,N_26179);
or U31468 (N_31468,N_25153,N_29768);
nand U31469 (N_31469,N_27023,N_27932);
and U31470 (N_31470,N_25563,N_28746);
nand U31471 (N_31471,N_29319,N_26680);
nor U31472 (N_31472,N_28371,N_26780);
xnor U31473 (N_31473,N_27598,N_26809);
xnor U31474 (N_31474,N_28680,N_28503);
nand U31475 (N_31475,N_28230,N_29179);
nor U31476 (N_31476,N_29689,N_26258);
xnor U31477 (N_31477,N_26931,N_25634);
nor U31478 (N_31478,N_28462,N_29370);
xnor U31479 (N_31479,N_25177,N_26959);
or U31480 (N_31480,N_26813,N_25888);
nand U31481 (N_31481,N_28614,N_27496);
or U31482 (N_31482,N_29487,N_29848);
xnor U31483 (N_31483,N_26598,N_29964);
and U31484 (N_31484,N_29026,N_25993);
nand U31485 (N_31485,N_28148,N_25307);
xnor U31486 (N_31486,N_26299,N_26615);
xor U31487 (N_31487,N_25155,N_29896);
and U31488 (N_31488,N_28288,N_26816);
and U31489 (N_31489,N_28625,N_26087);
or U31490 (N_31490,N_25368,N_28629);
xnor U31491 (N_31491,N_27332,N_25559);
nand U31492 (N_31492,N_26851,N_27727);
nand U31493 (N_31493,N_29286,N_27431);
nor U31494 (N_31494,N_28071,N_28786);
nand U31495 (N_31495,N_29387,N_28056);
and U31496 (N_31496,N_28084,N_25985);
and U31497 (N_31497,N_27765,N_29252);
nor U31498 (N_31498,N_25371,N_28408);
xnor U31499 (N_31499,N_26011,N_26321);
nor U31500 (N_31500,N_26362,N_28287);
nand U31501 (N_31501,N_25683,N_28967);
xnor U31502 (N_31502,N_25527,N_25278);
and U31503 (N_31503,N_27617,N_27477);
nand U31504 (N_31504,N_26913,N_26047);
or U31505 (N_31505,N_29852,N_29236);
nor U31506 (N_31506,N_28293,N_28713);
and U31507 (N_31507,N_28265,N_25715);
and U31508 (N_31508,N_29353,N_25317);
nor U31509 (N_31509,N_28675,N_28452);
or U31510 (N_31510,N_28199,N_28423);
and U31511 (N_31511,N_27741,N_27216);
xnor U31512 (N_31512,N_29826,N_26297);
and U31513 (N_31513,N_29560,N_27425);
and U31514 (N_31514,N_29667,N_28604);
or U31515 (N_31515,N_28513,N_27243);
nand U31516 (N_31516,N_29354,N_25899);
xor U31517 (N_31517,N_26647,N_28090);
and U31518 (N_31518,N_26194,N_28704);
nor U31519 (N_31519,N_29352,N_25238);
nand U31520 (N_31520,N_27770,N_28626);
nand U31521 (N_31521,N_28540,N_26278);
and U31522 (N_31522,N_25010,N_25335);
xor U31523 (N_31523,N_27345,N_26500);
or U31524 (N_31524,N_27560,N_29033);
xnor U31525 (N_31525,N_29463,N_26599);
or U31526 (N_31526,N_25176,N_26213);
nand U31527 (N_31527,N_29443,N_25092);
nor U31528 (N_31528,N_25431,N_27101);
nand U31529 (N_31529,N_29069,N_27493);
nor U31530 (N_31530,N_25025,N_26497);
or U31531 (N_31531,N_28816,N_26320);
nor U31532 (N_31532,N_27664,N_28030);
or U31533 (N_31533,N_26827,N_28619);
nand U31534 (N_31534,N_27406,N_29119);
or U31535 (N_31535,N_28903,N_29402);
xnor U31536 (N_31536,N_28202,N_28567);
or U31537 (N_31537,N_26548,N_26329);
or U31538 (N_31538,N_25562,N_28897);
nor U31539 (N_31539,N_25605,N_26091);
or U31540 (N_31540,N_27071,N_28365);
nor U31541 (N_31541,N_28821,N_28226);
xnor U31542 (N_31542,N_26884,N_27056);
and U31543 (N_31543,N_25690,N_25939);
nand U31544 (N_31544,N_27042,N_26078);
nand U31545 (N_31545,N_25735,N_29436);
nor U31546 (N_31546,N_25752,N_25561);
and U31547 (N_31547,N_28711,N_26452);
xnor U31548 (N_31548,N_26143,N_29440);
and U31549 (N_31549,N_27987,N_29458);
nor U31550 (N_31550,N_26796,N_25090);
nor U31551 (N_31551,N_25330,N_27975);
or U31552 (N_31552,N_26925,N_28279);
or U31553 (N_31553,N_29278,N_28338);
nor U31554 (N_31554,N_26192,N_26666);
and U31555 (N_31555,N_25900,N_26090);
nor U31556 (N_31556,N_28474,N_29815);
nor U31557 (N_31557,N_27867,N_27542);
and U31558 (N_31558,N_29920,N_26769);
and U31559 (N_31559,N_28784,N_27419);
xnor U31560 (N_31560,N_29481,N_28891);
nor U31561 (N_31561,N_29780,N_29589);
and U31562 (N_31562,N_25246,N_26417);
xor U31563 (N_31563,N_25789,N_29375);
nor U31564 (N_31564,N_25544,N_26123);
and U31565 (N_31565,N_26459,N_28368);
xor U31566 (N_31566,N_27890,N_26281);
nor U31567 (N_31567,N_28197,N_27512);
xnor U31568 (N_31568,N_29114,N_25971);
and U31569 (N_31569,N_29346,N_25816);
xnor U31570 (N_31570,N_28719,N_28795);
or U31571 (N_31571,N_25709,N_27487);
or U31572 (N_31572,N_25320,N_27716);
nor U31573 (N_31573,N_29185,N_27214);
and U31574 (N_31574,N_27736,N_28827);
nand U31575 (N_31575,N_29426,N_27837);
nand U31576 (N_31576,N_25991,N_28808);
and U31577 (N_31577,N_29199,N_27474);
and U31578 (N_31578,N_25649,N_25315);
or U31579 (N_31579,N_25135,N_28162);
or U31580 (N_31580,N_27279,N_25817);
nor U31581 (N_31581,N_29474,N_26823);
or U31582 (N_31582,N_27686,N_29478);
and U31583 (N_31583,N_29241,N_29492);
xor U31584 (N_31584,N_28301,N_27893);
xnor U31585 (N_31585,N_28034,N_29997);
nand U31586 (N_31586,N_27208,N_29452);
xnor U31587 (N_31587,N_27389,N_29597);
xor U31588 (N_31588,N_28558,N_26086);
or U31589 (N_31589,N_27040,N_29498);
or U31590 (N_31590,N_29694,N_29769);
nor U31591 (N_31591,N_25546,N_27887);
or U31592 (N_31592,N_27712,N_26818);
nor U31593 (N_31593,N_27261,N_25083);
nand U31594 (N_31594,N_26026,N_26786);
and U31595 (N_31595,N_25909,N_27548);
nand U31596 (N_31596,N_25211,N_28165);
xnor U31597 (N_31597,N_25271,N_27463);
and U31598 (N_31598,N_28812,N_26956);
xnor U31599 (N_31599,N_29125,N_29079);
nor U31600 (N_31600,N_25081,N_25249);
xor U31601 (N_31601,N_28981,N_26242);
nor U31602 (N_31602,N_26451,N_27907);
or U31603 (N_31603,N_28101,N_27685);
nor U31604 (N_31604,N_27636,N_25529);
nor U31605 (N_31605,N_25102,N_29911);
and U31606 (N_31606,N_26879,N_26431);
nand U31607 (N_31607,N_29798,N_27062);
and U31608 (N_31608,N_28692,N_29206);
xor U31609 (N_31609,N_25032,N_29625);
and U31610 (N_31610,N_27946,N_28878);
nand U31611 (N_31611,N_25321,N_25551);
xor U31612 (N_31612,N_29444,N_28936);
nor U31613 (N_31613,N_25499,N_26579);
nand U31614 (N_31614,N_28182,N_27387);
or U31615 (N_31615,N_26079,N_25085);
xnor U31616 (N_31616,N_29222,N_28430);
xnor U31617 (N_31617,N_25110,N_27451);
or U31618 (N_31618,N_28883,N_29679);
nand U31619 (N_31619,N_25129,N_25692);
xnor U31620 (N_31620,N_28294,N_27112);
xnor U31621 (N_31621,N_29811,N_28824);
xnor U31622 (N_31622,N_28523,N_28551);
or U31623 (N_31623,N_27706,N_27517);
nor U31624 (N_31624,N_27260,N_25009);
xnor U31625 (N_31625,N_28857,N_29067);
nor U31626 (N_31626,N_27338,N_28526);
or U31627 (N_31627,N_28873,N_25304);
and U31628 (N_31628,N_27581,N_25992);
and U31629 (N_31629,N_27798,N_27572);
nand U31630 (N_31630,N_29956,N_29374);
xor U31631 (N_31631,N_29159,N_29080);
nor U31632 (N_31632,N_29638,N_28486);
and U31633 (N_31633,N_26701,N_27523);
or U31634 (N_31634,N_27791,N_26427);
xor U31635 (N_31635,N_25305,N_28917);
and U31636 (N_31636,N_26231,N_28847);
nor U31637 (N_31637,N_25772,N_29285);
xor U31638 (N_31638,N_28145,N_27504);
nand U31639 (N_31639,N_28888,N_26753);
nand U31640 (N_31640,N_28774,N_28432);
xnor U31641 (N_31641,N_28654,N_29786);
xor U31642 (N_31642,N_29123,N_25724);
nor U31643 (N_31643,N_25370,N_29790);
and U31644 (N_31644,N_27004,N_25670);
xnor U31645 (N_31645,N_28601,N_29097);
and U31646 (N_31646,N_26714,N_25600);
xnor U31647 (N_31647,N_27763,N_27486);
and U31648 (N_31648,N_25504,N_29652);
nand U31649 (N_31649,N_28233,N_28023);
and U31650 (N_31650,N_26793,N_27481);
nand U31651 (N_31651,N_29203,N_26582);
nand U31652 (N_31652,N_26561,N_29303);
nand U31653 (N_31653,N_27983,N_29577);
nor U31654 (N_31654,N_29187,N_27100);
and U31655 (N_31655,N_26898,N_28035);
nand U31656 (N_31656,N_25671,N_26180);
xor U31657 (N_31657,N_27152,N_26351);
nor U31658 (N_31658,N_26955,N_26045);
and U31659 (N_31659,N_25444,N_25794);
and U31660 (N_31660,N_26062,N_27954);
and U31661 (N_31661,N_29269,N_28961);
or U31662 (N_31662,N_27722,N_25818);
nor U31663 (N_31663,N_28228,N_26102);
nor U31664 (N_31664,N_27938,N_29282);
xnor U31665 (N_31665,N_26608,N_27432);
xor U31666 (N_31666,N_25158,N_25813);
and U31667 (N_31667,N_26247,N_28098);
xnor U31668 (N_31668,N_28964,N_25777);
or U31669 (N_31669,N_27449,N_26754);
nand U31670 (N_31670,N_27485,N_28974);
xnor U31671 (N_31671,N_28422,N_26222);
nand U31672 (N_31672,N_29434,N_27702);
xor U31673 (N_31673,N_28983,N_29056);
or U31674 (N_31674,N_29937,N_25210);
or U31675 (N_31675,N_29578,N_25245);
and U31676 (N_31676,N_26727,N_29431);
xnor U31677 (N_31677,N_26563,N_29651);
or U31678 (N_31678,N_26758,N_25785);
nand U31679 (N_31679,N_25658,N_26654);
xor U31680 (N_31680,N_28492,N_27498);
nor U31681 (N_31681,N_28807,N_26988);
nand U31682 (N_31682,N_28544,N_27353);
or U31683 (N_31683,N_29006,N_29943);
xnor U31684 (N_31684,N_29238,N_29653);
nand U31685 (N_31685,N_26975,N_26294);
nand U31686 (N_31686,N_26783,N_25623);
nor U31687 (N_31687,N_27278,N_29543);
nor U31688 (N_31688,N_28405,N_25990);
and U31689 (N_31689,N_28130,N_28715);
xnor U31690 (N_31690,N_26658,N_26327);
nand U31691 (N_31691,N_25764,N_28469);
nand U31692 (N_31692,N_26474,N_27022);
nand U31693 (N_31693,N_26212,N_26857);
xor U31694 (N_31694,N_27324,N_27195);
nor U31695 (N_31695,N_26973,N_25578);
and U31696 (N_31696,N_25842,N_25645);
and U31697 (N_31697,N_28662,N_27357);
and U31698 (N_31698,N_28273,N_25506);
nor U31699 (N_31699,N_27471,N_28100);
and U31700 (N_31700,N_25560,N_26382);
nor U31701 (N_31701,N_28724,N_28379);
and U31702 (N_31702,N_28590,N_25687);
nand U31703 (N_31703,N_29566,N_27569);
and U31704 (N_31704,N_29482,N_28003);
or U31705 (N_31705,N_25200,N_28820);
or U31706 (N_31706,N_27187,N_28550);
nand U31707 (N_31707,N_27462,N_28382);
xor U31708 (N_31708,N_25334,N_26514);
or U31709 (N_31709,N_28027,N_25675);
nor U31710 (N_31710,N_26014,N_27737);
nor U31711 (N_31711,N_27901,N_26205);
nand U31712 (N_31712,N_27650,N_29733);
nor U31713 (N_31713,N_25823,N_26454);
nand U31714 (N_31714,N_27689,N_29789);
or U31715 (N_31715,N_29216,N_27917);
or U31716 (N_31716,N_27225,N_29761);
xor U31717 (N_31717,N_25869,N_26136);
nor U31718 (N_31718,N_28610,N_29556);
nand U31719 (N_31719,N_25876,N_26494);
nor U31720 (N_31720,N_26659,N_25587);
and U31721 (N_31721,N_28274,N_26400);
and U31722 (N_31722,N_27125,N_27057);
or U31723 (N_31723,N_29379,N_26870);
or U31724 (N_31724,N_28700,N_27868);
xor U31725 (N_31725,N_27624,N_27570);
and U31726 (N_31726,N_29744,N_26628);
xor U31727 (N_31727,N_29066,N_28583);
nand U31728 (N_31728,N_28052,N_27217);
nand U31729 (N_31729,N_27096,N_28120);
nor U31730 (N_31730,N_26130,N_29160);
xor U31731 (N_31731,N_26876,N_27175);
nand U31732 (N_31732,N_25841,N_26425);
nor U31733 (N_31733,N_26437,N_26137);
xor U31734 (N_31734,N_28494,N_28536);
xor U31735 (N_31735,N_26552,N_25161);
nand U31736 (N_31736,N_27222,N_28208);
nor U31737 (N_31737,N_26538,N_27236);
xnor U31738 (N_31738,N_28716,N_25406);
nand U31739 (N_31739,N_29162,N_28215);
or U31740 (N_31740,N_25862,N_27136);
nand U31741 (N_31741,N_29130,N_26915);
or U31742 (N_31742,N_25691,N_27323);
nor U31743 (N_31743,N_26782,N_29455);
nor U31744 (N_31744,N_26151,N_25837);
nor U31745 (N_31745,N_29669,N_26099);
and U31746 (N_31746,N_25000,N_27234);
xor U31747 (N_31747,N_28466,N_25622);
or U31748 (N_31748,N_27094,N_26840);
xor U31749 (N_31749,N_26795,N_27710);
xnor U31750 (N_31750,N_28132,N_28683);
xor U31751 (N_31751,N_27436,N_26938);
and U31752 (N_31752,N_27067,N_25834);
and U31753 (N_31753,N_29962,N_29433);
xnor U31754 (N_31754,N_29148,N_27554);
nor U31755 (N_31755,N_27468,N_26122);
xor U31756 (N_31756,N_25759,N_27045);
xor U31757 (N_31757,N_25056,N_25465);
nand U31758 (N_31758,N_27194,N_27138);
nand U31759 (N_31759,N_26426,N_28756);
xnor U31760 (N_31760,N_26287,N_28528);
and U31761 (N_31761,N_26812,N_29421);
nor U31762 (N_31762,N_26430,N_29757);
and U31763 (N_31763,N_26230,N_25312);
or U31764 (N_31764,N_26708,N_25585);
or U31765 (N_31765,N_26740,N_27122);
xor U31766 (N_31766,N_28328,N_29261);
or U31767 (N_31767,N_28094,N_26395);
or U31768 (N_31768,N_27097,N_25754);
xor U31769 (N_31769,N_25798,N_26236);
nand U31770 (N_31770,N_29591,N_29167);
nand U31771 (N_31771,N_29874,N_25470);
nand U31772 (N_31772,N_28911,N_29416);
nor U31773 (N_31773,N_25237,N_25749);
nand U31774 (N_31774,N_29272,N_29905);
nor U31775 (N_31775,N_25167,N_27355);
nand U31776 (N_31776,N_27502,N_27690);
and U31777 (N_31777,N_27044,N_28836);
nand U31778 (N_31778,N_27948,N_25648);
or U31779 (N_31779,N_27050,N_25969);
and U31780 (N_31780,N_25042,N_26960);
nand U31781 (N_31781,N_27597,N_27337);
xnor U31782 (N_31782,N_27153,N_27032);
nand U31783 (N_31783,N_29054,N_26495);
and U31784 (N_31784,N_25580,N_27120);
nand U31785 (N_31785,N_25400,N_28568);
or U31786 (N_31786,N_29857,N_29289);
and U31787 (N_31787,N_25701,N_26678);
or U31788 (N_31788,N_27220,N_26537);
and U31789 (N_31789,N_25289,N_28497);
nor U31790 (N_31790,N_29223,N_27461);
nor U31791 (N_31791,N_27775,N_28810);
nor U31792 (N_31792,N_27400,N_29000);
nor U31793 (N_31793,N_27376,N_27490);
and U31794 (N_31794,N_29177,N_27665);
nor U31795 (N_31795,N_28403,N_26298);
nand U31796 (N_31796,N_28584,N_26575);
nand U31797 (N_31797,N_25261,N_27290);
and U31798 (N_31798,N_27163,N_28971);
xor U31799 (N_31799,N_29037,N_26420);
and U31800 (N_31800,N_25235,N_28496);
or U31801 (N_31801,N_28081,N_25467);
and U31802 (N_31802,N_27133,N_27797);
nand U31803 (N_31803,N_29640,N_28329);
nand U31804 (N_31804,N_26947,N_28985);
nand U31805 (N_31805,N_28912,N_28075);
nor U31806 (N_31806,N_26076,N_26498);
nor U31807 (N_31807,N_25693,N_27472);
nand U31808 (N_31808,N_26486,N_27806);
xnor U31809 (N_31809,N_26585,N_29178);
or U31810 (N_31810,N_25427,N_27409);
or U31811 (N_31811,N_27093,N_27321);
nor U31812 (N_31812,N_29438,N_27037);
xor U31813 (N_31813,N_27544,N_27552);
nor U31814 (N_31814,N_27008,N_29939);
and U31815 (N_31815,N_27082,N_29432);
and U31816 (N_31816,N_25051,N_25020);
or U31817 (N_31817,N_26662,N_29523);
xor U31818 (N_31818,N_28929,N_28987);
nor U31819 (N_31819,N_26481,N_28986);
and U31820 (N_31820,N_25517,N_26622);
and U31821 (N_31821,N_25878,N_26559);
nor U31822 (N_31822,N_27439,N_26639);
xor U31823 (N_31823,N_26597,N_26280);
or U31824 (N_31824,N_27605,N_25157);
nor U31825 (N_31825,N_27030,N_25481);
nor U31826 (N_31826,N_27019,N_26246);
nor U31827 (N_31827,N_25514,N_26156);
xor U31828 (N_31828,N_27591,N_28586);
nand U31829 (N_31829,N_29220,N_26133);
and U31830 (N_31830,N_26348,N_25093);
or U31831 (N_31831,N_28159,N_29681);
and U31832 (N_31832,N_28177,N_29359);
nor U31833 (N_31833,N_29674,N_26574);
nor U31834 (N_31834,N_26802,N_25015);
nor U31835 (N_31835,N_29562,N_27514);
xnor U31836 (N_31836,N_29713,N_25513);
or U31837 (N_31837,N_25902,N_28147);
xor U31838 (N_31838,N_28900,N_27541);
nor U31839 (N_31839,N_28848,N_25989);
nand U31840 (N_31840,N_26074,N_27926);
and U31841 (N_31841,N_26638,N_28011);
xor U31842 (N_31842,N_28914,N_28562);
and U31843 (N_31843,N_26312,N_28800);
nand U31844 (N_31844,N_27146,N_28190);
and U31845 (N_31845,N_26875,N_29700);
nor U31846 (N_31846,N_29929,N_29044);
nand U31847 (N_31847,N_29738,N_28868);
nor U31848 (N_31848,N_29535,N_26613);
nand U31849 (N_31849,N_25280,N_25422);
nor U31850 (N_31850,N_29991,N_25418);
xnor U31851 (N_31851,N_29817,N_26976);
or U31852 (N_31852,N_27258,N_26107);
nand U31853 (N_31853,N_28672,N_27724);
nor U31854 (N_31854,N_27398,N_29600);
and U31855 (N_31855,N_25117,N_26689);
or U31856 (N_31856,N_26061,N_25525);
xor U31857 (N_31857,N_25287,N_29701);
nor U31858 (N_31858,N_27546,N_25980);
xnor U31859 (N_31859,N_29664,N_29335);
nor U31860 (N_31860,N_26735,N_26389);
nor U31861 (N_31861,N_28018,N_25306);
or U31862 (N_31862,N_29073,N_26825);
nand U31863 (N_31863,N_27335,N_27340);
or U31864 (N_31864,N_27055,N_27707);
and U31865 (N_31865,N_27202,N_29142);
or U31866 (N_31866,N_25100,N_26618);
nor U31867 (N_31867,N_28340,N_27126);
nand U31868 (N_31868,N_25127,N_29490);
and U31869 (N_31869,N_25864,N_25290);
and U31870 (N_31870,N_28123,N_29697);
nand U31871 (N_31871,N_28579,N_27458);
xor U31872 (N_31872,N_25667,N_25203);
nand U31873 (N_31873,N_26501,N_25733);
xnor U31874 (N_31874,N_28088,N_25323);
nand U31875 (N_31875,N_26733,N_27213);
and U31876 (N_31876,N_25268,N_28114);
xor U31877 (N_31877,N_26492,N_27824);
or U31878 (N_31878,N_25791,N_25863);
and U31879 (N_31879,N_25468,N_25197);
xor U31880 (N_31880,N_25069,N_26990);
nor U31881 (N_31881,N_25360,N_25891);
xor U31882 (N_31882,N_27176,N_29519);
xor U31883 (N_31883,N_27041,N_25607);
nor U31884 (N_31884,N_27259,N_28570);
nor U31885 (N_31885,N_26245,N_27524);
nor U31886 (N_31886,N_26075,N_26340);
and U31887 (N_31887,N_25569,N_28553);
xnor U31888 (N_31888,N_28416,N_29975);
and U31889 (N_31889,N_26743,N_26605);
and U31890 (N_31890,N_29144,N_27829);
xnor U31891 (N_31891,N_25205,N_26611);
or U31892 (N_31892,N_27885,N_26404);
or U31893 (N_31893,N_26534,N_29175);
and U31894 (N_31894,N_25445,N_26592);
xnor U31895 (N_31895,N_27255,N_28874);
nand U31896 (N_31896,N_27223,N_25265);
or U31897 (N_31897,N_29003,N_26392);
nand U31898 (N_31898,N_29493,N_27576);
xor U31899 (N_31899,N_29408,N_29599);
and U31900 (N_31900,N_29534,N_28309);
nand U31901 (N_31901,N_25542,N_29683);
xnor U31902 (N_31902,N_25353,N_25666);
and U31903 (N_31903,N_28588,N_26435);
nor U31904 (N_31904,N_26642,N_29201);
nand U31905 (N_31905,N_28395,N_26692);
nor U31906 (N_31906,N_27297,N_29545);
xor U31907 (N_31907,N_25377,N_27709);
and U31908 (N_31908,N_26858,N_29788);
or U31909 (N_31909,N_26519,N_26453);
xor U31910 (N_31910,N_28002,N_28046);
nor U31911 (N_31911,N_26527,N_27446);
and U31912 (N_31912,N_25039,N_28972);
or U31913 (N_31913,N_29833,N_25416);
xor U31914 (N_31914,N_28337,N_26021);
nand U31915 (N_31915,N_28645,N_29380);
and U31916 (N_31916,N_28600,N_29821);
or U31917 (N_31917,N_25224,N_28431);
nor U31918 (N_31918,N_29127,N_27875);
nor U31919 (N_31919,N_28156,N_27475);
and U31920 (N_31920,N_28390,N_28924);
or U31921 (N_31921,N_25905,N_29298);
xor U31922 (N_31922,N_27823,N_27129);
xor U31923 (N_31923,N_27116,N_25601);
nand U31924 (N_31924,N_25804,N_29168);
nand U31925 (N_31925,N_25700,N_29027);
nor U31926 (N_31926,N_26999,N_28651);
and U31927 (N_31927,N_27943,N_26810);
nand U31928 (N_31928,N_29522,N_28040);
nor U31929 (N_31929,N_28373,N_28186);
or U31930 (N_31930,N_29504,N_28140);
xor U31931 (N_31931,N_27967,N_27467);
nor U31932 (N_31932,N_27903,N_28398);
nor U31933 (N_31933,N_28988,N_28184);
and U31934 (N_31934,N_26147,N_27308);
nor U31935 (N_31935,N_25095,N_26414);
or U31936 (N_31936,N_25808,N_26227);
or U31937 (N_31937,N_25420,N_26874);
nand U31938 (N_31938,N_25413,N_26241);
and U31939 (N_31939,N_29171,N_27130);
nor U31940 (N_31940,N_29672,N_27166);
or U31941 (N_31941,N_27366,N_26182);
or U31942 (N_31942,N_29239,N_26846);
nand U31943 (N_31943,N_27207,N_25951);
or U31944 (N_31944,N_29395,N_29341);
nand U31945 (N_31945,N_25617,N_26150);
or U31946 (N_31946,N_25403,N_26590);
nor U31947 (N_31947,N_26066,N_28261);
and U31948 (N_31948,N_26696,N_27769);
and U31949 (N_31949,N_25496,N_29930);
nor U31950 (N_31950,N_29132,N_27621);
xnor U31951 (N_31951,N_27231,N_27950);
or U31952 (N_31952,N_29349,N_28354);
nand U31953 (N_31953,N_28220,N_28589);
nand U31954 (N_31954,N_27772,N_28477);
nor U31955 (N_31955,N_29954,N_28930);
nand U31956 (N_31956,N_25296,N_27359);
nand U31957 (N_31957,N_25588,N_27896);
and U31958 (N_31958,N_25314,N_28131);
and U31959 (N_31959,N_29940,N_29869);
xor U31960 (N_31960,N_29849,N_28278);
and U31961 (N_31961,N_29517,N_29691);
and U31962 (N_31962,N_26342,N_28342);
or U31963 (N_31963,N_27892,N_25462);
and U31964 (N_31964,N_29961,N_26667);
nand U31965 (N_31965,N_27293,N_28595);
or U31966 (N_31966,N_25633,N_28752);
nor U31967 (N_31967,N_28227,N_25209);
or U31968 (N_31968,N_25848,N_25128);
xnor U31969 (N_31969,N_25681,N_25115);
nand U31970 (N_31970,N_29775,N_26336);
or U31971 (N_31971,N_25191,N_25625);
and U31972 (N_31972,N_25664,N_29342);
nand U31973 (N_31973,N_29392,N_28245);
and U31974 (N_31974,N_25638,N_29071);
or U31975 (N_31975,N_28105,N_27010);
nand U31976 (N_31976,N_26979,N_26996);
nor U31977 (N_31977,N_26661,N_28627);
nor U31978 (N_31978,N_29714,N_26259);
or U31979 (N_31979,N_28118,N_25395);
nor U31980 (N_31980,N_29254,N_29102);
nor U31981 (N_31981,N_28507,N_26706);
xor U31982 (N_31982,N_28168,N_25659);
or U31983 (N_31983,N_25730,N_25219);
nor U31984 (N_31984,N_25206,N_25441);
xnor U31985 (N_31985,N_28851,N_29036);
or U31986 (N_31986,N_29660,N_27963);
xor U31987 (N_31987,N_27984,N_25933);
and U31988 (N_31988,N_26216,N_26487);
xnor U31989 (N_31989,N_25917,N_26705);
and U31990 (N_31990,N_28709,N_25570);
or U31991 (N_31991,N_27522,N_25510);
nand U31992 (N_31992,N_27347,N_28525);
nor U31993 (N_31993,N_25434,N_27334);
nor U31994 (N_31994,N_25455,N_27306);
xor U31995 (N_31995,N_27922,N_28237);
or U31996 (N_31996,N_25443,N_29603);
and U31997 (N_31997,N_25075,N_29902);
nor U31998 (N_31998,N_29676,N_25581);
xor U31999 (N_31999,N_25912,N_27280);
or U32000 (N_32000,N_26784,N_27921);
nand U32001 (N_32001,N_26089,N_25640);
nand U32002 (N_32002,N_26134,N_27215);
nand U32003 (N_32003,N_26375,N_29366);
xnor U32004 (N_32004,N_29933,N_25494);
xnor U32005 (N_32005,N_27072,N_25398);
nor U32006 (N_32006,N_25340,N_25475);
nor U32007 (N_32007,N_29411,N_26712);
and U32008 (N_32008,N_28946,N_25889);
nand U32009 (N_32009,N_27853,N_29629);
nor U32010 (N_32010,N_26384,N_28445);
and U32011 (N_32011,N_29483,N_25758);
nor U32012 (N_32012,N_26270,N_28678);
nand U32013 (N_32013,N_26867,N_25356);
xnor U32014 (N_32014,N_26645,N_29795);
nor U32015 (N_32015,N_25926,N_28977);
and U32016 (N_32016,N_28493,N_26549);
nor U32017 (N_32017,N_28019,N_28674);
and U32018 (N_32018,N_28532,N_27962);
and U32019 (N_32019,N_26616,N_27190);
or U32020 (N_32020,N_29410,N_28246);
or U32021 (N_32021,N_25713,N_26736);
xnor U32022 (N_32022,N_29260,N_29836);
xor U32023 (N_32023,N_26239,N_29984);
and U32024 (N_32024,N_25948,N_29019);
nor U32025 (N_32025,N_26511,N_25058);
xor U32026 (N_32026,N_27184,N_26097);
nand U32027 (N_32027,N_28884,N_25108);
or U32028 (N_32028,N_27316,N_27083);
nor U32029 (N_32029,N_28041,N_26621);
nand U32030 (N_32030,N_27895,N_28412);
xnor U32031 (N_32031,N_28351,N_27318);
nor U32032 (N_32032,N_26787,N_29693);
xnor U32033 (N_32033,N_28172,N_26862);
nand U32034 (N_32034,N_27897,N_29089);
nor U32035 (N_32035,N_27415,N_29182);
nor U32036 (N_32036,N_29516,N_26800);
nand U32037 (N_32037,N_25795,N_26791);
nor U32038 (N_32038,N_29976,N_26305);
or U32039 (N_32039,N_29549,N_29109);
nand U32040 (N_32040,N_29637,N_26531);
xnor U32041 (N_32041,N_26967,N_28976);
or U32042 (N_32042,N_27578,N_29708);
nand U32043 (N_32043,N_28111,N_27854);
nor U32044 (N_32044,N_29855,N_26201);
and U32045 (N_32045,N_29267,N_25079);
and U32046 (N_32046,N_28923,N_27739);
nor U32047 (N_32047,N_28241,N_27815);
nand U32048 (N_32048,N_28407,N_27286);
and U32049 (N_32049,N_25279,N_25495);
nand U32050 (N_32050,N_25631,N_29210);
xnor U32051 (N_32051,N_26721,N_29018);
nor U32052 (N_32052,N_28024,N_26848);
xor U32053 (N_32053,N_26441,N_28420);
or U32054 (N_32054,N_26323,N_25089);
or U32055 (N_32055,N_26663,N_27511);
nand U32056 (N_32056,N_25234,N_26589);
nand U32057 (N_32057,N_28958,N_29008);
nand U32058 (N_32058,N_26543,N_27711);
or U32059 (N_32059,N_29234,N_29126);
xor U32060 (N_32060,N_27600,N_26082);
and U32061 (N_32061,N_29274,N_29547);
nor U32062 (N_32062,N_27307,N_26202);
and U32063 (N_32063,N_28066,N_28599);
and U32064 (N_32064,N_28886,N_26069);
or U32065 (N_32065,N_28129,N_28690);
nand U32066 (N_32066,N_26629,N_29647);
nor U32067 (N_32067,N_28206,N_25858);
and U32068 (N_32068,N_25112,N_29100);
xor U32069 (N_32069,N_26146,N_26127);
nor U32070 (N_32070,N_26660,N_25859);
xnor U32071 (N_32071,N_26466,N_27173);
nor U32072 (N_32072,N_29755,N_26890);
or U32073 (N_32073,N_27484,N_29406);
nor U32074 (N_32074,N_25226,N_25313);
nand U32075 (N_32075,N_27627,N_29314);
or U32076 (N_32076,N_27390,N_28789);
nand U32077 (N_32077,N_26887,N_25003);
or U32078 (N_32078,N_27740,N_27268);
or U32079 (N_32079,N_27488,N_28556);
and U32080 (N_32080,N_29361,N_28457);
xnor U32081 (N_32081,N_26698,N_25087);
or U32082 (N_32082,N_27652,N_29322);
and U32083 (N_32083,N_27981,N_25449);
or U32084 (N_32084,N_27103,N_27043);
nor U32085 (N_32085,N_29176,N_28116);
or U32086 (N_32086,N_28677,N_28249);
nand U32087 (N_32087,N_26077,N_26376);
nor U32088 (N_32088,N_25214,N_25822);
xor U32089 (N_32089,N_28266,N_29404);
xnor U32090 (N_32090,N_25695,N_27677);
nand U32091 (N_32091,N_29020,N_25140);
or U32092 (N_32092,N_29351,N_26625);
or U32093 (N_32093,N_27088,N_26318);
nand U32094 (N_32094,N_27626,N_29542);
or U32095 (N_32095,N_26475,N_26070);
or U32096 (N_32096,N_28085,N_26541);
and U32097 (N_32097,N_27311,N_28815);
and U32098 (N_32098,N_29403,N_25921);
xor U32099 (N_32099,N_27756,N_25484);
or U32100 (N_32100,N_27421,N_26416);
nor U32101 (N_32101,N_29518,N_27275);
nor U32102 (N_32102,N_25378,N_27456);
xnor U32103 (N_32103,N_27666,N_27310);
or U32104 (N_32104,N_25122,N_29590);
or U32105 (N_32105,N_29763,N_26571);
nand U32106 (N_32106,N_26643,N_27908);
xor U32107 (N_32107,N_26600,N_28045);
xnor U32108 (N_32108,N_28534,N_28070);
nor U32109 (N_32109,N_28904,N_29581);
nand U32110 (N_32110,N_27361,N_26989);
and U32111 (N_32111,N_26991,N_28778);
or U32112 (N_32112,N_25532,N_26369);
or U32113 (N_32113,N_27836,N_25835);
xor U32114 (N_32114,N_28310,N_28016);
and U32115 (N_32115,N_27373,N_26694);
and U32116 (N_32116,N_26771,N_28901);
nand U32117 (N_32117,N_26251,N_27422);
nor U32118 (N_32118,N_28442,N_28686);
and U32119 (N_32119,N_25901,N_25608);
or U32120 (N_32120,N_28652,N_26665);
and U32121 (N_32121,N_27265,N_26215);
or U32122 (N_32122,N_27006,N_26195);
or U32123 (N_32123,N_27344,N_28561);
and U32124 (N_32124,N_28875,N_25591);
xnor U32125 (N_32125,N_25928,N_25940);
or U32126 (N_32126,N_29906,N_28214);
nor U32127 (N_32127,N_29865,N_25556);
xnor U32128 (N_32128,N_29068,N_29887);
nor U32129 (N_32129,N_25071,N_26728);
nor U32130 (N_32130,N_29748,N_25186);
xor U32131 (N_32131,N_27609,N_29750);
xor U32132 (N_32132,N_25458,N_26518);
nor U32133 (N_32133,N_29015,N_27744);
or U32134 (N_32134,N_27731,N_25598);
or U32135 (N_32135,N_27407,N_29233);
and U32136 (N_32136,N_26773,N_28267);
nand U32137 (N_32137,N_29034,N_28054);
nand U32138 (N_32138,N_29023,N_27675);
nor U32139 (N_32139,N_29398,N_28262);
or U32140 (N_32140,N_29031,N_28264);
or U32141 (N_32141,N_28012,N_26634);
or U32142 (N_32142,N_28710,N_26347);
nand U32143 (N_32143,N_27024,N_29766);
or U32144 (N_32144,N_27571,N_27678);
and U32145 (N_32145,N_27700,N_25829);
nor U32146 (N_32146,N_27513,N_26986);
nand U32147 (N_32147,N_29587,N_27002);
and U32148 (N_32148,N_28582,N_26716);
or U32149 (N_32149,N_25421,N_25753);
nor U32150 (N_32150,N_28834,N_26037);
xor U32151 (N_32151,N_28925,N_26394);
and U32152 (N_32152,N_28248,N_25870);
or U32153 (N_32153,N_26225,N_25394);
and U32154 (N_32154,N_29908,N_27121);
and U32155 (N_32155,N_26550,N_27864);
nor U32156 (N_32156,N_27628,N_26217);
and U32157 (N_32157,N_27991,N_29138);
xnor U32158 (N_32158,N_28015,N_25783);
and U32159 (N_32159,N_25997,N_28169);
or U32160 (N_32160,N_29536,N_28780);
nor U32161 (N_32161,N_26944,N_25941);
nand U32162 (N_32162,N_28853,N_26244);
and U32163 (N_32163,N_25050,N_29035);
nand U32164 (N_32164,N_25509,N_29726);
nand U32165 (N_32165,N_27882,N_27774);
nand U32166 (N_32166,N_27778,N_27914);
nand U32167 (N_32167,N_26255,N_25892);
xnor U32168 (N_32168,N_27314,N_25283);
nand U32169 (N_32169,N_29951,N_25528);
nor U32170 (N_32170,N_28480,N_27610);
and U32171 (N_32171,N_26359,N_27401);
nor U32172 (N_32172,N_28427,N_28612);
xor U32173 (N_32173,N_29506,N_29838);
and U32174 (N_32174,N_25722,N_28943);
and U32175 (N_32175,N_26157,N_28608);
nor U32176 (N_32176,N_28707,N_26854);
xnor U32177 (N_32177,N_27237,N_28158);
xnor U32178 (N_32178,N_26726,N_25195);
nand U32179 (N_32179,N_28842,N_25114);
and U32180 (N_32180,N_27704,N_28250);
or U32181 (N_32181,N_27540,N_29328);
or U32182 (N_32182,N_25453,N_27573);
nor U32183 (N_32183,N_26065,N_25731);
and U32184 (N_32184,N_29344,N_25336);
nor U32185 (N_32185,N_28417,N_25979);
nand U32186 (N_32186,N_26183,N_25408);
nand U32187 (N_32187,N_27437,N_28060);
or U32188 (N_32188,N_25363,N_26768);
nor U32189 (N_32189,N_25407,N_28517);
nor U32190 (N_32190,N_27757,N_29949);
nor U32191 (N_32191,N_27426,N_29383);
and U32192 (N_32192,N_29013,N_27264);
xor U32193 (N_32193,N_29413,N_27701);
and U32194 (N_32194,N_27221,N_28560);
or U32195 (N_32195,N_26448,N_28613);
xor U32196 (N_32196,N_29091,N_28291);
nor U32197 (N_32197,N_25616,N_27492);
nor U32198 (N_32198,N_26853,N_29378);
or U32199 (N_32199,N_25482,N_27448);
or U32200 (N_32200,N_29570,N_25471);
xor U32201 (N_32201,N_26670,N_29134);
or U32202 (N_32202,N_28119,N_27683);
nor U32203 (N_32203,N_29129,N_28028);
nor U32204 (N_32204,N_28063,N_26322);
nor U32205 (N_32205,N_27454,N_26043);
or U32206 (N_32206,N_25472,N_25192);
or U32207 (N_32207,N_27955,N_28933);
and U32208 (N_32208,N_28885,N_27326);
nand U32209 (N_32209,N_29368,N_26567);
nor U32210 (N_32210,N_26580,N_27608);
nand U32211 (N_32211,N_25906,N_26366);
xnor U32212 (N_32212,N_29612,N_28730);
nand U32213 (N_32213,N_26349,N_26335);
xor U32214 (N_32214,N_29039,N_27746);
and U32215 (N_32215,N_28449,N_28658);
or U32216 (N_32216,N_28104,N_27147);
nor U32217 (N_32217,N_28356,N_29725);
nand U32218 (N_32218,N_25338,N_28000);
xor U32219 (N_32219,N_26463,N_29196);
nand U32220 (N_32220,N_28804,N_26300);
nor U32221 (N_32221,N_27858,N_25222);
xnor U32222 (N_32222,N_27090,N_25392);
or U32223 (N_32223,N_29367,N_27079);
and U32224 (N_32224,N_26036,N_25362);
or U32225 (N_32225,N_29802,N_28546);
nand U32226 (N_32226,N_27563,N_25043);
nand U32227 (N_32227,N_27996,N_29616);
or U32228 (N_32228,N_27986,N_26723);
xnor U32229 (N_32229,N_29099,N_28598);
and U32230 (N_32230,N_26871,N_27413);
xnor U32231 (N_32231,N_29806,N_25104);
nand U32232 (N_32232,N_25807,N_25672);
and U32233 (N_32233,N_29526,N_26191);
and U32234 (N_32234,N_26777,N_28072);
or U32235 (N_32235,N_28263,N_29558);
xor U32236 (N_32236,N_28524,N_26265);
and U32237 (N_32237,N_27009,N_25319);
nand U32238 (N_32238,N_29369,N_28059);
nand U32239 (N_32239,N_26681,N_26684);
nor U32240 (N_32240,N_26253,N_29847);
nor U32241 (N_32241,N_27343,N_29770);
xnor U32242 (N_32242,N_27470,N_25723);
nor U32243 (N_32243,N_25915,N_29555);
or U32244 (N_32244,N_27117,N_25452);
or U32245 (N_32245,N_27651,N_27378);
nand U32246 (N_32246,N_28346,N_28994);
nor U32247 (N_32247,N_27728,N_28581);
nand U32248 (N_32248,N_25073,N_27497);
and U32249 (N_32249,N_28404,N_26177);
nor U32250 (N_32250,N_29208,N_25111);
or U32251 (N_32251,N_28173,N_27843);
xor U32252 (N_32252,N_25185,N_25663);
nor U32253 (N_32253,N_29828,N_27721);
nor U32254 (N_32254,N_28047,N_26480);
nor U32255 (N_32255,N_28498,N_27641);
xnor U32256 (N_32256,N_26476,N_26664);
nand U32257 (N_32257,N_25145,N_28944);
xor U32258 (N_32258,N_29501,N_29029);
nand U32259 (N_32259,N_29935,N_25439);
or U32260 (N_32260,N_25652,N_29969);
xnor U32261 (N_32261,N_27341,N_28307);
nand U32262 (N_32262,N_28316,N_25328);
and U32263 (N_32263,N_26878,N_25960);
or U32264 (N_32264,N_28641,N_29532);
and U32265 (N_32265,N_26053,N_25144);
or U32266 (N_32266,N_28991,N_28125);
nand U32267 (N_32267,N_29508,N_25389);
nor U32268 (N_32268,N_28750,N_27482);
nor U32269 (N_32269,N_28623,N_26093);
or U32270 (N_32270,N_28067,N_27228);
nor U32271 (N_32271,N_28017,N_26536);
and U32272 (N_32272,N_26751,N_26623);
xnor U32273 (N_32273,N_26088,N_25827);
and U32274 (N_32274,N_26640,N_29279);
xor U32275 (N_32275,N_29793,N_25165);
xor U32276 (N_32276,N_27203,N_29559);
xnor U32277 (N_32277,N_26262,N_28840);
nor U32278 (N_32278,N_25805,N_25097);
nor U32279 (N_32279,N_27403,N_27533);
or U32280 (N_32280,N_26040,N_28324);
or U32281 (N_32281,N_25516,N_29909);
or U32282 (N_32282,N_25552,N_29221);
nand U32283 (N_32283,N_29551,N_29630);
nor U32284 (N_32284,N_28200,N_29661);
or U32285 (N_32285,N_27262,N_28421);
nor U32286 (N_32286,N_26978,N_27393);
nand U32287 (N_32287,N_25292,N_25417);
nand U32288 (N_32288,N_25380,N_25615);
or U32289 (N_32289,N_25503,N_26232);
or U32290 (N_32290,N_29537,N_27713);
and U32291 (N_32291,N_28270,N_27028);
or U32292 (N_32292,N_25604,N_28969);
and U32293 (N_32293,N_27520,N_29718);
and U32294 (N_32294,N_28144,N_26833);
xor U32295 (N_32295,N_29794,N_26291);
xnor U32296 (N_32296,N_26928,N_26408);
and U32297 (N_32297,N_25215,N_26807);
and U32298 (N_32298,N_25994,N_28760);
or U32299 (N_32299,N_28906,N_28566);
xnor U32300 (N_32300,N_29372,N_28527);
xnor U32301 (N_32301,N_28388,N_27483);
and U32302 (N_32302,N_27031,N_28074);
and U32303 (N_32303,N_27164,N_28149);
nor U32304 (N_32304,N_26838,N_27543);
or U32305 (N_32305,N_29287,N_29919);
and U32306 (N_32306,N_28960,N_27305);
xor U32307 (N_32307,N_26277,N_28653);
nand U32308 (N_32308,N_27592,N_26607);
xnor U32309 (N_32309,N_29851,N_28455);
xor U32310 (N_32310,N_28905,N_26310);
or U32311 (N_32311,N_26170,N_28669);
xor U32312 (N_32312,N_27250,N_27304);
or U32313 (N_32313,N_25181,N_28401);
nand U32314 (N_32314,N_29494,N_28178);
nand U32315 (N_32315,N_29450,N_27388);
or U32316 (N_32316,N_26022,N_27098);
and U32317 (N_32317,N_28740,N_27245);
or U32318 (N_32318,N_27866,N_26720);
nand U32319 (N_32319,N_25137,N_27160);
xnor U32320 (N_32320,N_28259,N_29813);
or U32321 (N_32321,N_28718,N_29685);
nor U32322 (N_32322,N_28860,N_29358);
and U32323 (N_32323,N_27561,N_29678);
nor U32324 (N_32324,N_27659,N_28349);
nor U32325 (N_32325,N_25454,N_26604);
nor U32326 (N_32326,N_27803,N_25149);
and U32327 (N_32327,N_25393,N_25066);
nor U32328 (N_32328,N_27106,N_26926);
or U32329 (N_32329,N_26282,N_25961);
nor U32330 (N_32330,N_29856,N_25522);
xor U32331 (N_32331,N_25786,N_27499);
nand U32332 (N_32332,N_26912,N_29211);
nand U32333 (N_32333,N_26499,N_28048);
nand U32334 (N_32334,N_27060,N_26657);
nand U32335 (N_32335,N_29907,N_28013);
xor U32336 (N_32336,N_26891,N_28872);
xnor U32337 (N_32337,N_25610,N_27780);
or U32338 (N_32338,N_28319,N_29819);
nor U32339 (N_32339,N_26028,N_26315);
and U32340 (N_32340,N_29680,N_26371);
nand U32341 (N_32341,N_25790,N_27852);
nor U32342 (N_32342,N_29890,N_26929);
nand U32343 (N_32343,N_26866,N_29982);
or U32344 (N_32344,N_28137,N_25299);
nand U32345 (N_32345,N_29724,N_26042);
xnor U32346 (N_32346,N_27330,N_29243);
or U32347 (N_32347,N_27247,N_29942);
or U32348 (N_32348,N_28510,N_26199);
nor U32349 (N_32349,N_27365,N_27978);
and U32350 (N_32350,N_29525,N_29740);
nand U32351 (N_32351,N_27077,N_27405);
nand U32352 (N_32352,N_27382,N_26709);
nor U32353 (N_32353,N_25256,N_27839);
xor U32354 (N_32354,N_28022,N_25619);
nand U32355 (N_32355,N_27503,N_28665);
nand U32356 (N_32356,N_27070,N_26722);
nand U32357 (N_32357,N_25707,N_25599);
or U32358 (N_32358,N_28134,N_28754);
xor U32359 (N_32359,N_27014,N_25259);
or U32360 (N_32360,N_27860,N_28539);
nor U32361 (N_32361,N_29076,N_26302);
xor U32362 (N_32362,N_27762,N_29963);
and U32363 (N_32363,N_25179,N_25932);
xor U32364 (N_32364,N_25346,N_25409);
nor U32365 (N_32365,N_28849,N_27253);
and U32366 (N_32366,N_28628,N_27871);
xor U32367 (N_32367,N_25719,N_27976);
and U32368 (N_32368,N_29461,N_27900);
or U32369 (N_32369,N_26814,N_26439);
xnor U32370 (N_32370,N_27397,N_26415);
or U32371 (N_32371,N_26935,N_25850);
nor U32372 (N_32372,N_25964,N_28185);
nand U32373 (N_32373,N_25714,N_27154);
nand U32374 (N_32374,N_27633,N_25309);
xor U32375 (N_32375,N_26081,N_25603);
nor U32376 (N_32376,N_26211,N_29512);
or U32377 (N_32377,N_29886,N_29327);
or U32378 (N_32378,N_27622,N_27204);
and U32379 (N_32379,N_27833,N_29829);
or U32380 (N_32380,N_26909,N_25076);
nand U32381 (N_32381,N_27494,N_29417);
and U32382 (N_32382,N_25929,N_28764);
or U32383 (N_32383,N_27281,N_27747);
xnor U32384 (N_32384,N_27979,N_26413);
nor U32385 (N_32385,N_27519,N_25548);
nor U32386 (N_32386,N_27283,N_29670);
or U32387 (N_32387,N_27568,N_25886);
nor U32388 (N_32388,N_28243,N_29086);
or U32389 (N_32389,N_25298,N_25833);
nand U32390 (N_32390,N_29166,N_25639);
nand U32391 (N_32391,N_26163,N_29384);
nor U32392 (N_32392,N_27282,N_27115);
and U32393 (N_32393,N_25589,N_25121);
nand U32394 (N_32394,N_25464,N_29418);
nor U32395 (N_32395,N_29414,N_26652);
nor U32396 (N_32396,N_28372,N_25703);
or U32397 (N_32397,N_27480,N_29796);
or U32398 (N_32398,N_29009,N_26092);
xnor U32399 (N_32399,N_29101,N_26888);
nor U32400 (N_32400,N_28633,N_28321);
nor U32401 (N_32401,N_25375,N_25830);
and U32402 (N_32402,N_25047,N_29317);
or U32403 (N_32403,N_29771,N_27924);
nor U32404 (N_32404,N_27309,N_25005);
nor U32405 (N_32405,N_28284,N_28095);
or U32406 (N_32406,N_28736,N_27870);
and U32407 (N_32407,N_25225,N_25437);
and U32408 (N_32408,N_25415,N_26350);
and U32409 (N_32409,N_27669,N_28042);
or U32410 (N_32410,N_26223,N_29574);
and U32411 (N_32411,N_28021,N_29970);
nand U32412 (N_32412,N_25358,N_29360);
nand U32413 (N_32413,N_29038,N_25846);
or U32414 (N_32414,N_26055,N_26341);
nor U32415 (N_32415,N_27185,N_26249);
and U32416 (N_32416,N_26080,N_29230);
nand U32417 (N_32417,N_25898,N_27751);
xnor U32418 (N_32418,N_25763,N_29903);
nor U32419 (N_32419,N_26309,N_27654);
nand U32420 (N_32420,N_27531,N_27886);
nand U32421 (N_32421,N_27428,N_28751);
nand U32422 (N_32422,N_28343,N_26581);
nor U32423 (N_32423,N_29644,N_28845);
and U32424 (N_32424,N_29717,N_28932);
or U32425 (N_32425,N_27233,N_26637);
nor U32426 (N_32426,N_26485,N_27241);
and U32427 (N_32427,N_26119,N_25381);
or U32428 (N_32428,N_28092,N_27256);
and U32429 (N_32429,N_27013,N_27607);
xor U32430 (N_32430,N_29040,N_29394);
nand U32431 (N_32431,N_29792,N_28788);
or U32432 (N_32432,N_25568,N_27819);
and U32433 (N_32433,N_29471,N_28086);
nor U32434 (N_32434,N_29749,N_29552);
or U32435 (N_32435,N_27992,N_27396);
xnor U32436 (N_32436,N_26820,N_28681);
nor U32437 (N_32437,N_28210,N_28467);
or U32438 (N_32438,N_27132,N_29807);
nor U32439 (N_32439,N_28315,N_25021);
or U32440 (N_32440,N_25303,N_26892);
nor U32441 (N_32441,N_26264,N_25343);
nand U32442 (N_32442,N_29318,N_26693);
and U32443 (N_32443,N_29212,N_26697);
xnor U32444 (N_32444,N_26513,N_29255);
nand U32445 (N_32445,N_26160,N_26443);
xor U32446 (N_32446,N_25678,N_25811);
nand U32447 (N_32447,N_29495,N_27219);
nand U32448 (N_32448,N_29528,N_27192);
xnor U32449 (N_32449,N_25967,N_27408);
and U32450 (N_32450,N_26540,N_29133);
nor U32451 (N_32451,N_26445,N_28889);
or U32452 (N_32452,N_27688,N_26505);
and U32453 (N_32453,N_29297,N_26738);
or U32454 (N_32454,N_25350,N_28955);
xor U32455 (N_32455,N_29197,N_29065);
and U32456 (N_32456,N_25430,N_29377);
or U32457 (N_32457,N_25379,N_26602);
nor U32458 (N_32458,N_25739,N_27970);
and U32459 (N_32459,N_29760,N_25202);
nand U32460 (N_32460,N_25175,N_27168);
or U32461 (N_32461,N_27107,N_29400);
and U32462 (N_32462,N_26883,N_28978);
xnor U32463 (N_32463,N_28326,N_29617);
or U32464 (N_32464,N_27141,N_27551);
xor U32465 (N_32465,N_28453,N_29391);
or U32466 (N_32466,N_27840,N_28630);
and U32467 (N_32467,N_29575,N_29623);
nand U32468 (N_32468,N_28865,N_28603);
nand U32469 (N_32469,N_28631,N_29799);
nand U32470 (N_32470,N_26115,N_26096);
nor U32471 (N_32471,N_25386,N_28026);
and U32472 (N_32472,N_25660,N_28970);
and U32473 (N_32473,N_28456,N_29032);
or U32474 (N_32474,N_29622,N_26799);
nor U32475 (N_32475,N_28956,N_29834);
nor U32476 (N_32476,N_25273,N_26003);
and U32477 (N_32477,N_26275,N_28515);
xnor U32478 (N_32478,N_28636,N_29832);
and U32479 (N_32479,N_27526,N_27193);
or U32480 (N_32480,N_29131,N_27113);
nor U32481 (N_32481,N_25812,N_26285);
or U32482 (N_32482,N_25945,N_28171);
xnor U32483 (N_32483,N_26460,N_27993);
nand U32484 (N_32484,N_28871,N_26184);
nor U32485 (N_32485,N_29042,N_26449);
and U32486 (N_32486,N_26594,N_25220);
nand U32487 (N_32487,N_28223,N_26094);
or U32488 (N_32488,N_29049,N_29992);
or U32489 (N_32489,N_27080,N_26806);
or U32490 (N_32490,N_25944,N_25843);
nor U32491 (N_32491,N_28921,N_28039);
nand U32492 (N_32492,N_25264,N_26254);
nor U32493 (N_32493,N_27015,N_28573);
and U32494 (N_32494,N_27003,N_27235);
or U32495 (N_32495,N_29415,N_25911);
xor U32496 (N_32496,N_27360,N_28722);
xnor U32497 (N_32497,N_25286,N_25364);
and U32498 (N_32498,N_25436,N_29104);
or U32499 (N_32499,N_28320,N_29041);
xor U32500 (N_32500,N_26114,N_27554);
or U32501 (N_32501,N_26644,N_28883);
xor U32502 (N_32502,N_25709,N_28320);
xor U32503 (N_32503,N_27721,N_26573);
and U32504 (N_32504,N_29690,N_29917);
nor U32505 (N_32505,N_26509,N_27242);
xnor U32506 (N_32506,N_26837,N_27404);
xor U32507 (N_32507,N_28613,N_27131);
nand U32508 (N_32508,N_27201,N_25990);
nand U32509 (N_32509,N_25621,N_27113);
nand U32510 (N_32510,N_26151,N_29832);
and U32511 (N_32511,N_28959,N_29446);
or U32512 (N_32512,N_25319,N_26088);
nand U32513 (N_32513,N_25929,N_25264);
nor U32514 (N_32514,N_28894,N_28398);
nand U32515 (N_32515,N_26838,N_29230);
nor U32516 (N_32516,N_28530,N_27220);
or U32517 (N_32517,N_29060,N_25064);
nor U32518 (N_32518,N_25901,N_28265);
and U32519 (N_32519,N_28771,N_29173);
nand U32520 (N_32520,N_28753,N_26808);
or U32521 (N_32521,N_29539,N_26668);
xor U32522 (N_32522,N_25495,N_29348);
nor U32523 (N_32523,N_28764,N_27904);
nand U32524 (N_32524,N_27950,N_29002);
and U32525 (N_32525,N_25284,N_28166);
or U32526 (N_32526,N_26152,N_29107);
and U32527 (N_32527,N_28476,N_29063);
xnor U32528 (N_32528,N_27481,N_27761);
nor U32529 (N_32529,N_26471,N_26407);
and U32530 (N_32530,N_27414,N_28261);
xnor U32531 (N_32531,N_28594,N_27384);
nor U32532 (N_32532,N_28372,N_27000);
or U32533 (N_32533,N_28354,N_27060);
xor U32534 (N_32534,N_27660,N_27493);
nand U32535 (N_32535,N_25083,N_27760);
or U32536 (N_32536,N_29679,N_27757);
nand U32537 (N_32537,N_26686,N_28699);
and U32538 (N_32538,N_25210,N_26241);
nor U32539 (N_32539,N_29075,N_29052);
nor U32540 (N_32540,N_27331,N_25678);
or U32541 (N_32541,N_28826,N_28306);
and U32542 (N_32542,N_27471,N_29376);
nor U32543 (N_32543,N_27636,N_25596);
nand U32544 (N_32544,N_25110,N_26397);
nor U32545 (N_32545,N_29108,N_28531);
and U32546 (N_32546,N_25170,N_29435);
nor U32547 (N_32547,N_29402,N_26037);
nand U32548 (N_32548,N_26411,N_28069);
xnor U32549 (N_32549,N_25334,N_28727);
and U32550 (N_32550,N_27962,N_26049);
nor U32551 (N_32551,N_28515,N_27424);
and U32552 (N_32552,N_27651,N_28297);
nor U32553 (N_32553,N_28125,N_26419);
or U32554 (N_32554,N_28753,N_25881);
nor U32555 (N_32555,N_25986,N_26744);
and U32556 (N_32556,N_27458,N_27755);
or U32557 (N_32557,N_25230,N_29247);
and U32558 (N_32558,N_26215,N_25734);
xor U32559 (N_32559,N_29243,N_26661);
nand U32560 (N_32560,N_29375,N_26433);
nand U32561 (N_32561,N_27102,N_26046);
nand U32562 (N_32562,N_26417,N_26097);
xor U32563 (N_32563,N_28787,N_29699);
and U32564 (N_32564,N_27494,N_28850);
xnor U32565 (N_32565,N_25052,N_26240);
nand U32566 (N_32566,N_25512,N_28265);
and U32567 (N_32567,N_26485,N_29145);
nor U32568 (N_32568,N_25672,N_28867);
xnor U32569 (N_32569,N_25850,N_27267);
nand U32570 (N_32570,N_29882,N_28748);
and U32571 (N_32571,N_25220,N_28395);
nor U32572 (N_32572,N_28140,N_28169);
nand U32573 (N_32573,N_29012,N_26371);
nor U32574 (N_32574,N_26795,N_28811);
nor U32575 (N_32575,N_26295,N_28732);
xor U32576 (N_32576,N_27958,N_28769);
nand U32577 (N_32577,N_27294,N_27895);
nor U32578 (N_32578,N_28530,N_28235);
xor U32579 (N_32579,N_27173,N_28065);
xnor U32580 (N_32580,N_29236,N_26807);
nand U32581 (N_32581,N_26448,N_26847);
or U32582 (N_32582,N_25227,N_26997);
xnor U32583 (N_32583,N_25316,N_27371);
nand U32584 (N_32584,N_26720,N_26047);
or U32585 (N_32585,N_26191,N_27288);
nand U32586 (N_32586,N_25398,N_29004);
nand U32587 (N_32587,N_28721,N_25191);
nor U32588 (N_32588,N_27436,N_28088);
nand U32589 (N_32589,N_28706,N_27062);
nand U32590 (N_32590,N_29993,N_25428);
and U32591 (N_32591,N_29606,N_27781);
and U32592 (N_32592,N_26688,N_25430);
or U32593 (N_32593,N_26814,N_26808);
nor U32594 (N_32594,N_25385,N_26755);
or U32595 (N_32595,N_27890,N_25982);
nand U32596 (N_32596,N_25554,N_29030);
and U32597 (N_32597,N_28142,N_25814);
nand U32598 (N_32598,N_28055,N_27661);
xnor U32599 (N_32599,N_25641,N_27908);
and U32600 (N_32600,N_25606,N_28070);
xnor U32601 (N_32601,N_28232,N_26730);
or U32602 (N_32602,N_25090,N_25374);
nand U32603 (N_32603,N_28131,N_29672);
nor U32604 (N_32604,N_25764,N_29692);
and U32605 (N_32605,N_28788,N_28985);
and U32606 (N_32606,N_25837,N_28729);
xor U32607 (N_32607,N_26816,N_29855);
nand U32608 (N_32608,N_25265,N_29158);
or U32609 (N_32609,N_29554,N_28848);
nand U32610 (N_32610,N_28248,N_27387);
xor U32611 (N_32611,N_28753,N_29911);
nand U32612 (N_32612,N_25029,N_26069);
nand U32613 (N_32613,N_26238,N_26684);
xor U32614 (N_32614,N_26780,N_25619);
xor U32615 (N_32615,N_29489,N_27799);
nor U32616 (N_32616,N_25737,N_27242);
and U32617 (N_32617,N_29155,N_26042);
xnor U32618 (N_32618,N_28939,N_26161);
and U32619 (N_32619,N_28960,N_27441);
nand U32620 (N_32620,N_29800,N_25722);
and U32621 (N_32621,N_28011,N_29951);
xnor U32622 (N_32622,N_26664,N_27342);
xor U32623 (N_32623,N_25575,N_27556);
and U32624 (N_32624,N_28759,N_25767);
nand U32625 (N_32625,N_28216,N_27178);
nor U32626 (N_32626,N_29716,N_28370);
nor U32627 (N_32627,N_28181,N_28717);
nand U32628 (N_32628,N_28177,N_27450);
and U32629 (N_32629,N_28383,N_28748);
nor U32630 (N_32630,N_29817,N_26462);
or U32631 (N_32631,N_25273,N_27557);
and U32632 (N_32632,N_28796,N_25307);
or U32633 (N_32633,N_29271,N_29578);
and U32634 (N_32634,N_27118,N_27300);
xor U32635 (N_32635,N_25560,N_29588);
or U32636 (N_32636,N_29266,N_27795);
nand U32637 (N_32637,N_29248,N_28556);
xor U32638 (N_32638,N_25526,N_28175);
nor U32639 (N_32639,N_29023,N_29649);
nand U32640 (N_32640,N_28213,N_26297);
xnor U32641 (N_32641,N_27458,N_25746);
nand U32642 (N_32642,N_29996,N_29895);
nor U32643 (N_32643,N_29907,N_28475);
or U32644 (N_32644,N_28456,N_28201);
nand U32645 (N_32645,N_25409,N_26370);
xnor U32646 (N_32646,N_25843,N_26777);
and U32647 (N_32647,N_27757,N_28452);
and U32648 (N_32648,N_29842,N_25312);
nand U32649 (N_32649,N_25047,N_26636);
nand U32650 (N_32650,N_29361,N_27221);
nand U32651 (N_32651,N_28111,N_28324);
nor U32652 (N_32652,N_28533,N_26818);
and U32653 (N_32653,N_25104,N_25995);
nor U32654 (N_32654,N_26285,N_29460);
and U32655 (N_32655,N_29699,N_28904);
and U32656 (N_32656,N_28308,N_29565);
and U32657 (N_32657,N_27748,N_27362);
xor U32658 (N_32658,N_28687,N_26376);
or U32659 (N_32659,N_26129,N_29994);
or U32660 (N_32660,N_26844,N_28937);
and U32661 (N_32661,N_28762,N_25663);
nand U32662 (N_32662,N_27334,N_29143);
xor U32663 (N_32663,N_26323,N_25125);
and U32664 (N_32664,N_26852,N_28181);
nor U32665 (N_32665,N_27035,N_27760);
nor U32666 (N_32666,N_28489,N_28356);
nand U32667 (N_32667,N_27971,N_27515);
or U32668 (N_32668,N_26840,N_26671);
nor U32669 (N_32669,N_28992,N_29192);
xor U32670 (N_32670,N_25918,N_25606);
or U32671 (N_32671,N_25014,N_26927);
nor U32672 (N_32672,N_25632,N_27512);
nand U32673 (N_32673,N_27794,N_26727);
xor U32674 (N_32674,N_28474,N_27800);
nor U32675 (N_32675,N_29725,N_28933);
xnor U32676 (N_32676,N_25411,N_25426);
and U32677 (N_32677,N_28623,N_25901);
xor U32678 (N_32678,N_29984,N_28166);
xnor U32679 (N_32679,N_26943,N_28524);
xnor U32680 (N_32680,N_28528,N_28946);
xor U32681 (N_32681,N_26525,N_28130);
nor U32682 (N_32682,N_26479,N_27017);
and U32683 (N_32683,N_27462,N_25620);
nor U32684 (N_32684,N_25150,N_25657);
nor U32685 (N_32685,N_27081,N_27456);
or U32686 (N_32686,N_28475,N_26931);
xnor U32687 (N_32687,N_25613,N_28974);
nand U32688 (N_32688,N_29347,N_27081);
nand U32689 (N_32689,N_25778,N_27989);
and U32690 (N_32690,N_27897,N_28787);
nand U32691 (N_32691,N_27574,N_27477);
nor U32692 (N_32692,N_26743,N_28701);
nor U32693 (N_32693,N_25889,N_25335);
and U32694 (N_32694,N_28861,N_25197);
and U32695 (N_32695,N_27564,N_28019);
nor U32696 (N_32696,N_27186,N_25105);
and U32697 (N_32697,N_29873,N_28750);
xor U32698 (N_32698,N_28168,N_25044);
xnor U32699 (N_32699,N_28807,N_29223);
xor U32700 (N_32700,N_29285,N_25716);
xor U32701 (N_32701,N_29921,N_29107);
and U32702 (N_32702,N_27200,N_27259);
xnor U32703 (N_32703,N_25820,N_25965);
and U32704 (N_32704,N_26028,N_25264);
or U32705 (N_32705,N_25886,N_28102);
xnor U32706 (N_32706,N_26194,N_27030);
or U32707 (N_32707,N_29388,N_29863);
or U32708 (N_32708,N_25341,N_25560);
nor U32709 (N_32709,N_25367,N_27164);
nand U32710 (N_32710,N_25394,N_28956);
nand U32711 (N_32711,N_25837,N_27942);
or U32712 (N_32712,N_25299,N_25533);
xnor U32713 (N_32713,N_25900,N_26422);
nand U32714 (N_32714,N_28611,N_26087);
and U32715 (N_32715,N_29051,N_28610);
nor U32716 (N_32716,N_25684,N_28895);
xor U32717 (N_32717,N_25900,N_26309);
or U32718 (N_32718,N_28554,N_25074);
nor U32719 (N_32719,N_29942,N_25260);
nor U32720 (N_32720,N_29730,N_29412);
nand U32721 (N_32721,N_26132,N_28728);
or U32722 (N_32722,N_25154,N_29394);
xnor U32723 (N_32723,N_27458,N_26868);
xor U32724 (N_32724,N_29833,N_29278);
and U32725 (N_32725,N_29057,N_25077);
nor U32726 (N_32726,N_29746,N_27256);
nor U32727 (N_32727,N_29268,N_29537);
nor U32728 (N_32728,N_25734,N_29136);
xor U32729 (N_32729,N_28021,N_27237);
nor U32730 (N_32730,N_28146,N_26404);
xnor U32731 (N_32731,N_25403,N_27934);
nand U32732 (N_32732,N_29473,N_26935);
nor U32733 (N_32733,N_28180,N_26700);
nor U32734 (N_32734,N_27659,N_26006);
xor U32735 (N_32735,N_27877,N_26312);
and U32736 (N_32736,N_25615,N_29144);
xnor U32737 (N_32737,N_25182,N_29992);
nor U32738 (N_32738,N_28445,N_28069);
xor U32739 (N_32739,N_27279,N_29215);
nor U32740 (N_32740,N_25866,N_25994);
and U32741 (N_32741,N_28091,N_27223);
nand U32742 (N_32742,N_27995,N_25339);
nand U32743 (N_32743,N_29195,N_27205);
nor U32744 (N_32744,N_27183,N_25025);
or U32745 (N_32745,N_28942,N_26808);
or U32746 (N_32746,N_26736,N_25216);
or U32747 (N_32747,N_29474,N_29884);
nor U32748 (N_32748,N_27126,N_28543);
nand U32749 (N_32749,N_26832,N_25390);
nor U32750 (N_32750,N_29632,N_29031);
and U32751 (N_32751,N_27808,N_27962);
xor U32752 (N_32752,N_27223,N_28918);
and U32753 (N_32753,N_26030,N_27503);
or U32754 (N_32754,N_25873,N_29702);
nand U32755 (N_32755,N_26989,N_29881);
nor U32756 (N_32756,N_25109,N_27637);
nor U32757 (N_32757,N_29351,N_27621);
nand U32758 (N_32758,N_26174,N_26682);
nor U32759 (N_32759,N_25819,N_26173);
and U32760 (N_32760,N_27307,N_25597);
and U32761 (N_32761,N_28432,N_28161);
xnor U32762 (N_32762,N_28404,N_26284);
nand U32763 (N_32763,N_26213,N_29737);
or U32764 (N_32764,N_28807,N_27101);
xnor U32765 (N_32765,N_27565,N_29612);
or U32766 (N_32766,N_27510,N_27164);
xor U32767 (N_32767,N_25176,N_28289);
and U32768 (N_32768,N_25438,N_29536);
and U32769 (N_32769,N_25745,N_28086);
nand U32770 (N_32770,N_28252,N_28528);
nor U32771 (N_32771,N_27402,N_29026);
and U32772 (N_32772,N_26915,N_28954);
or U32773 (N_32773,N_28292,N_25100);
xnor U32774 (N_32774,N_27617,N_28944);
nor U32775 (N_32775,N_29920,N_26292);
xnor U32776 (N_32776,N_27035,N_29080);
nor U32777 (N_32777,N_25944,N_25091);
xor U32778 (N_32778,N_28829,N_29953);
and U32779 (N_32779,N_26818,N_28028);
xnor U32780 (N_32780,N_25720,N_29882);
nand U32781 (N_32781,N_25035,N_25629);
nand U32782 (N_32782,N_27280,N_28048);
or U32783 (N_32783,N_29793,N_28174);
xor U32784 (N_32784,N_28557,N_28834);
nand U32785 (N_32785,N_25884,N_28599);
or U32786 (N_32786,N_25868,N_28586);
nor U32787 (N_32787,N_26526,N_26605);
or U32788 (N_32788,N_28923,N_29988);
xor U32789 (N_32789,N_28927,N_27803);
xor U32790 (N_32790,N_28099,N_28015);
nand U32791 (N_32791,N_29566,N_25640);
and U32792 (N_32792,N_29049,N_28807);
or U32793 (N_32793,N_29308,N_29559);
nor U32794 (N_32794,N_27981,N_26730);
xnor U32795 (N_32795,N_28387,N_28267);
or U32796 (N_32796,N_29391,N_28900);
xnor U32797 (N_32797,N_28008,N_27838);
or U32798 (N_32798,N_27499,N_26440);
and U32799 (N_32799,N_29275,N_27180);
xnor U32800 (N_32800,N_29052,N_27595);
nand U32801 (N_32801,N_27195,N_29082);
xor U32802 (N_32802,N_25460,N_25089);
or U32803 (N_32803,N_26618,N_26202);
or U32804 (N_32804,N_26663,N_25344);
or U32805 (N_32805,N_25706,N_25447);
nand U32806 (N_32806,N_26051,N_28710);
xor U32807 (N_32807,N_29930,N_26725);
nor U32808 (N_32808,N_25956,N_25090);
and U32809 (N_32809,N_26604,N_27744);
nor U32810 (N_32810,N_25268,N_28670);
nand U32811 (N_32811,N_29157,N_29631);
and U32812 (N_32812,N_26745,N_29634);
and U32813 (N_32813,N_27029,N_29068);
or U32814 (N_32814,N_26443,N_29320);
and U32815 (N_32815,N_28882,N_27713);
and U32816 (N_32816,N_25857,N_26759);
nor U32817 (N_32817,N_27623,N_25814);
nand U32818 (N_32818,N_27190,N_25083);
nor U32819 (N_32819,N_29525,N_28470);
nand U32820 (N_32820,N_27302,N_28092);
or U32821 (N_32821,N_25138,N_28397);
or U32822 (N_32822,N_29388,N_29132);
and U32823 (N_32823,N_28417,N_26722);
and U32824 (N_32824,N_25375,N_27867);
or U32825 (N_32825,N_27450,N_26436);
nand U32826 (N_32826,N_29972,N_25953);
nand U32827 (N_32827,N_29035,N_28693);
or U32828 (N_32828,N_27967,N_26782);
nor U32829 (N_32829,N_26978,N_26182);
or U32830 (N_32830,N_26488,N_29250);
nor U32831 (N_32831,N_26874,N_29293);
and U32832 (N_32832,N_26763,N_25356);
xnor U32833 (N_32833,N_28051,N_25734);
nor U32834 (N_32834,N_25514,N_27773);
nand U32835 (N_32835,N_25842,N_28630);
nor U32836 (N_32836,N_25993,N_29980);
xnor U32837 (N_32837,N_28182,N_26186);
or U32838 (N_32838,N_26161,N_27084);
and U32839 (N_32839,N_26433,N_25409);
and U32840 (N_32840,N_29882,N_28977);
or U32841 (N_32841,N_27591,N_26792);
nand U32842 (N_32842,N_29653,N_27013);
nand U32843 (N_32843,N_29404,N_29965);
and U32844 (N_32844,N_26854,N_25675);
xnor U32845 (N_32845,N_25548,N_25877);
and U32846 (N_32846,N_28198,N_25639);
xor U32847 (N_32847,N_26967,N_29493);
nand U32848 (N_32848,N_27217,N_25780);
and U32849 (N_32849,N_26791,N_28792);
and U32850 (N_32850,N_25612,N_28309);
nand U32851 (N_32851,N_29068,N_25101);
xnor U32852 (N_32852,N_27242,N_25028);
or U32853 (N_32853,N_29490,N_27960);
nor U32854 (N_32854,N_25362,N_27958);
nand U32855 (N_32855,N_26192,N_26602);
nor U32856 (N_32856,N_28622,N_29521);
xnor U32857 (N_32857,N_27569,N_28640);
or U32858 (N_32858,N_27839,N_26905);
and U32859 (N_32859,N_28748,N_28764);
and U32860 (N_32860,N_25568,N_29255);
and U32861 (N_32861,N_29663,N_25537);
xor U32862 (N_32862,N_27653,N_27359);
and U32863 (N_32863,N_28357,N_27161);
xor U32864 (N_32864,N_28282,N_28717);
nand U32865 (N_32865,N_28181,N_29316);
nand U32866 (N_32866,N_29312,N_28868);
nand U32867 (N_32867,N_29937,N_26126);
and U32868 (N_32868,N_27645,N_28008);
or U32869 (N_32869,N_28578,N_29163);
xnor U32870 (N_32870,N_26419,N_27479);
xor U32871 (N_32871,N_26504,N_28162);
nor U32872 (N_32872,N_25544,N_27538);
xor U32873 (N_32873,N_26288,N_27487);
nand U32874 (N_32874,N_28249,N_25466);
and U32875 (N_32875,N_29373,N_28449);
xnor U32876 (N_32876,N_29140,N_25612);
xor U32877 (N_32877,N_25399,N_29588);
nand U32878 (N_32878,N_25317,N_25467);
and U32879 (N_32879,N_27800,N_26085);
or U32880 (N_32880,N_28213,N_26584);
and U32881 (N_32881,N_29897,N_28129);
xor U32882 (N_32882,N_26306,N_26552);
or U32883 (N_32883,N_28491,N_28485);
xor U32884 (N_32884,N_26642,N_26308);
nor U32885 (N_32885,N_28736,N_25508);
and U32886 (N_32886,N_25757,N_26638);
and U32887 (N_32887,N_28355,N_28102);
nor U32888 (N_32888,N_25280,N_28744);
nand U32889 (N_32889,N_28910,N_25404);
or U32890 (N_32890,N_26148,N_27962);
xnor U32891 (N_32891,N_28060,N_25348);
nor U32892 (N_32892,N_29307,N_26112);
nor U32893 (N_32893,N_28619,N_25764);
and U32894 (N_32894,N_27257,N_27410);
nand U32895 (N_32895,N_28295,N_28893);
and U32896 (N_32896,N_29479,N_26187);
xor U32897 (N_32897,N_27392,N_28490);
nand U32898 (N_32898,N_26736,N_28642);
nand U32899 (N_32899,N_27373,N_25246);
nand U32900 (N_32900,N_28076,N_26556);
xnor U32901 (N_32901,N_26014,N_28257);
nand U32902 (N_32902,N_26323,N_29988);
nor U32903 (N_32903,N_27199,N_25070);
nor U32904 (N_32904,N_26158,N_29659);
nor U32905 (N_32905,N_26491,N_29985);
xor U32906 (N_32906,N_27790,N_29643);
xor U32907 (N_32907,N_29335,N_25763);
xor U32908 (N_32908,N_27248,N_25099);
and U32909 (N_32909,N_29181,N_25537);
or U32910 (N_32910,N_29804,N_29834);
nor U32911 (N_32911,N_28439,N_27187);
and U32912 (N_32912,N_25312,N_26222);
or U32913 (N_32913,N_27267,N_29324);
nor U32914 (N_32914,N_28394,N_28096);
xor U32915 (N_32915,N_28151,N_27034);
or U32916 (N_32916,N_25551,N_26846);
nor U32917 (N_32917,N_25574,N_28776);
xor U32918 (N_32918,N_29015,N_25914);
and U32919 (N_32919,N_25671,N_27653);
and U32920 (N_32920,N_26415,N_28950);
nor U32921 (N_32921,N_25280,N_27514);
nor U32922 (N_32922,N_26425,N_28153);
or U32923 (N_32923,N_25846,N_26783);
and U32924 (N_32924,N_29906,N_26114);
nand U32925 (N_32925,N_29160,N_27043);
nand U32926 (N_32926,N_27175,N_29639);
nand U32927 (N_32927,N_25727,N_27549);
nor U32928 (N_32928,N_25826,N_27807);
nand U32929 (N_32929,N_27311,N_25190);
nor U32930 (N_32930,N_25248,N_25782);
nor U32931 (N_32931,N_29935,N_26966);
nor U32932 (N_32932,N_29824,N_29548);
and U32933 (N_32933,N_28071,N_25950);
or U32934 (N_32934,N_25813,N_26743);
and U32935 (N_32935,N_27415,N_26598);
nand U32936 (N_32936,N_28295,N_25928);
or U32937 (N_32937,N_26062,N_28438);
nand U32938 (N_32938,N_25880,N_28297);
or U32939 (N_32939,N_27380,N_27878);
nor U32940 (N_32940,N_27730,N_27128);
nand U32941 (N_32941,N_25529,N_27541);
and U32942 (N_32942,N_27628,N_25430);
or U32943 (N_32943,N_28420,N_28796);
xnor U32944 (N_32944,N_28325,N_27084);
nor U32945 (N_32945,N_25169,N_25669);
and U32946 (N_32946,N_26086,N_25092);
xnor U32947 (N_32947,N_26433,N_25416);
or U32948 (N_32948,N_25539,N_28293);
nand U32949 (N_32949,N_25294,N_26219);
nor U32950 (N_32950,N_28224,N_25661);
xor U32951 (N_32951,N_26462,N_28477);
nand U32952 (N_32952,N_29250,N_29195);
and U32953 (N_32953,N_26352,N_29346);
nand U32954 (N_32954,N_27617,N_27428);
and U32955 (N_32955,N_27709,N_28286);
nor U32956 (N_32956,N_29871,N_29276);
and U32957 (N_32957,N_25942,N_27984);
xnor U32958 (N_32958,N_29723,N_27051);
nor U32959 (N_32959,N_28035,N_28729);
nand U32960 (N_32960,N_28327,N_25127);
or U32961 (N_32961,N_26520,N_29919);
nand U32962 (N_32962,N_28419,N_28481);
nor U32963 (N_32963,N_28634,N_26929);
nand U32964 (N_32964,N_26857,N_29533);
nand U32965 (N_32965,N_28119,N_26988);
nand U32966 (N_32966,N_27238,N_29720);
or U32967 (N_32967,N_25376,N_28199);
or U32968 (N_32968,N_26246,N_28694);
nand U32969 (N_32969,N_26855,N_28652);
or U32970 (N_32970,N_27354,N_25630);
nand U32971 (N_32971,N_29784,N_28425);
nand U32972 (N_32972,N_27331,N_28803);
or U32973 (N_32973,N_27336,N_25951);
nor U32974 (N_32974,N_26000,N_27365);
xnor U32975 (N_32975,N_25151,N_25206);
nand U32976 (N_32976,N_28781,N_29048);
and U32977 (N_32977,N_29585,N_27307);
nor U32978 (N_32978,N_27717,N_27076);
xnor U32979 (N_32979,N_29915,N_26410);
and U32980 (N_32980,N_25959,N_25649);
nor U32981 (N_32981,N_26169,N_28982);
nand U32982 (N_32982,N_28406,N_28162);
and U32983 (N_32983,N_29562,N_28490);
xor U32984 (N_32984,N_26817,N_26110);
xor U32985 (N_32985,N_25227,N_29916);
nor U32986 (N_32986,N_26064,N_26315);
and U32987 (N_32987,N_29067,N_29816);
or U32988 (N_32988,N_25231,N_27946);
nor U32989 (N_32989,N_26036,N_25110);
nor U32990 (N_32990,N_26421,N_26575);
xnor U32991 (N_32991,N_28730,N_27503);
or U32992 (N_32992,N_28522,N_26646);
or U32993 (N_32993,N_28825,N_27836);
or U32994 (N_32994,N_28537,N_26028);
nor U32995 (N_32995,N_27675,N_29737);
or U32996 (N_32996,N_28102,N_27927);
and U32997 (N_32997,N_28255,N_25781);
xnor U32998 (N_32998,N_29090,N_26651);
or U32999 (N_32999,N_26145,N_29318);
or U33000 (N_33000,N_26745,N_28012);
and U33001 (N_33001,N_27520,N_28184);
and U33002 (N_33002,N_29814,N_29678);
or U33003 (N_33003,N_29313,N_27785);
or U33004 (N_33004,N_29730,N_29561);
or U33005 (N_33005,N_27520,N_26998);
nor U33006 (N_33006,N_29497,N_25509);
or U33007 (N_33007,N_26746,N_27204);
nor U33008 (N_33008,N_27323,N_28861);
xnor U33009 (N_33009,N_27175,N_25766);
nor U33010 (N_33010,N_26296,N_29518);
nand U33011 (N_33011,N_27008,N_28245);
or U33012 (N_33012,N_27860,N_26234);
nand U33013 (N_33013,N_27156,N_26290);
nor U33014 (N_33014,N_26388,N_28974);
or U33015 (N_33015,N_26017,N_28464);
nand U33016 (N_33016,N_25583,N_25399);
nor U33017 (N_33017,N_26875,N_25746);
or U33018 (N_33018,N_27998,N_26094);
or U33019 (N_33019,N_28427,N_27499);
and U33020 (N_33020,N_26569,N_29547);
xnor U33021 (N_33021,N_25862,N_26442);
or U33022 (N_33022,N_27831,N_28350);
xor U33023 (N_33023,N_26404,N_28041);
xor U33024 (N_33024,N_25730,N_27656);
or U33025 (N_33025,N_26651,N_29040);
or U33026 (N_33026,N_25509,N_29934);
and U33027 (N_33027,N_29599,N_27730);
or U33028 (N_33028,N_27334,N_27046);
xnor U33029 (N_33029,N_29997,N_28425);
nor U33030 (N_33030,N_29806,N_26405);
nor U33031 (N_33031,N_27601,N_27242);
nand U33032 (N_33032,N_29996,N_25917);
nand U33033 (N_33033,N_26689,N_25843);
nor U33034 (N_33034,N_28577,N_27302);
nand U33035 (N_33035,N_29342,N_29189);
xor U33036 (N_33036,N_26726,N_27953);
nor U33037 (N_33037,N_28643,N_26525);
and U33038 (N_33038,N_26654,N_26447);
and U33039 (N_33039,N_26891,N_27822);
xor U33040 (N_33040,N_25835,N_27835);
xor U33041 (N_33041,N_25698,N_25615);
and U33042 (N_33042,N_29244,N_25254);
nand U33043 (N_33043,N_28485,N_27935);
or U33044 (N_33044,N_26615,N_27347);
nor U33045 (N_33045,N_25895,N_29358);
nand U33046 (N_33046,N_29549,N_25491);
and U33047 (N_33047,N_26099,N_27098);
and U33048 (N_33048,N_28097,N_25765);
xnor U33049 (N_33049,N_28682,N_27771);
xor U33050 (N_33050,N_25371,N_25992);
nand U33051 (N_33051,N_25784,N_28328);
xnor U33052 (N_33052,N_27290,N_27575);
or U33053 (N_33053,N_26418,N_26900);
xor U33054 (N_33054,N_26939,N_28498);
nor U33055 (N_33055,N_27297,N_26046);
nand U33056 (N_33056,N_28671,N_28601);
or U33057 (N_33057,N_25040,N_28848);
nand U33058 (N_33058,N_28209,N_29032);
or U33059 (N_33059,N_29907,N_26774);
xor U33060 (N_33060,N_28619,N_29138);
nand U33061 (N_33061,N_26693,N_27661);
xor U33062 (N_33062,N_25877,N_27220);
or U33063 (N_33063,N_27167,N_27132);
nor U33064 (N_33064,N_27309,N_27788);
xor U33065 (N_33065,N_25511,N_26729);
xor U33066 (N_33066,N_27928,N_29547);
nor U33067 (N_33067,N_26568,N_29274);
and U33068 (N_33068,N_28116,N_29125);
nor U33069 (N_33069,N_28909,N_29231);
and U33070 (N_33070,N_26278,N_26284);
or U33071 (N_33071,N_28191,N_29412);
xnor U33072 (N_33072,N_25355,N_28109);
nand U33073 (N_33073,N_28786,N_27994);
xor U33074 (N_33074,N_27766,N_27950);
nor U33075 (N_33075,N_28702,N_26823);
nand U33076 (N_33076,N_28565,N_25081);
or U33077 (N_33077,N_26684,N_28931);
nor U33078 (N_33078,N_29641,N_25402);
and U33079 (N_33079,N_29028,N_29738);
nor U33080 (N_33080,N_25037,N_26351);
and U33081 (N_33081,N_27939,N_28259);
nand U33082 (N_33082,N_26971,N_28501);
nand U33083 (N_33083,N_25323,N_25798);
nand U33084 (N_33084,N_27922,N_29814);
xnor U33085 (N_33085,N_26352,N_27803);
nor U33086 (N_33086,N_28365,N_29617);
xnor U33087 (N_33087,N_27473,N_25504);
nand U33088 (N_33088,N_27703,N_25568);
and U33089 (N_33089,N_28318,N_28456);
nor U33090 (N_33090,N_25727,N_28796);
and U33091 (N_33091,N_27761,N_29056);
nand U33092 (N_33092,N_28269,N_29805);
nand U33093 (N_33093,N_28545,N_29857);
or U33094 (N_33094,N_29785,N_26313);
xnor U33095 (N_33095,N_26644,N_25332);
and U33096 (N_33096,N_29733,N_25052);
nor U33097 (N_33097,N_26230,N_25280);
or U33098 (N_33098,N_27130,N_29391);
nand U33099 (N_33099,N_26966,N_25267);
or U33100 (N_33100,N_26943,N_25464);
or U33101 (N_33101,N_26856,N_26596);
nor U33102 (N_33102,N_27479,N_28243);
xor U33103 (N_33103,N_26709,N_27663);
nor U33104 (N_33104,N_25791,N_25687);
and U33105 (N_33105,N_28771,N_25328);
nand U33106 (N_33106,N_26628,N_26570);
or U33107 (N_33107,N_25930,N_28482);
nand U33108 (N_33108,N_29576,N_27779);
nor U33109 (N_33109,N_25151,N_29482);
or U33110 (N_33110,N_28670,N_25419);
nor U33111 (N_33111,N_27979,N_25624);
nand U33112 (N_33112,N_26823,N_25328);
nand U33113 (N_33113,N_29399,N_28742);
or U33114 (N_33114,N_26181,N_29094);
and U33115 (N_33115,N_29886,N_25707);
nor U33116 (N_33116,N_28559,N_29332);
and U33117 (N_33117,N_28430,N_26827);
nor U33118 (N_33118,N_28258,N_27635);
nand U33119 (N_33119,N_27675,N_25732);
nand U33120 (N_33120,N_26671,N_26715);
nand U33121 (N_33121,N_29613,N_27328);
or U33122 (N_33122,N_25321,N_29961);
or U33123 (N_33123,N_29182,N_27723);
nand U33124 (N_33124,N_25598,N_25096);
xor U33125 (N_33125,N_29449,N_25062);
or U33126 (N_33126,N_29371,N_29863);
nor U33127 (N_33127,N_29722,N_25590);
nor U33128 (N_33128,N_29097,N_27680);
or U33129 (N_33129,N_25359,N_26942);
nor U33130 (N_33130,N_25407,N_27936);
and U33131 (N_33131,N_26395,N_25491);
nor U33132 (N_33132,N_26766,N_28253);
xor U33133 (N_33133,N_29960,N_29961);
xnor U33134 (N_33134,N_26001,N_28123);
nand U33135 (N_33135,N_29615,N_25145);
xnor U33136 (N_33136,N_27981,N_26581);
or U33137 (N_33137,N_29110,N_25020);
nand U33138 (N_33138,N_28288,N_27528);
or U33139 (N_33139,N_28435,N_28985);
nand U33140 (N_33140,N_27489,N_26870);
nor U33141 (N_33141,N_27362,N_27753);
and U33142 (N_33142,N_28991,N_25706);
or U33143 (N_33143,N_28560,N_28995);
or U33144 (N_33144,N_29582,N_29978);
and U33145 (N_33145,N_27205,N_26247);
xor U33146 (N_33146,N_27960,N_29376);
nand U33147 (N_33147,N_26132,N_25755);
or U33148 (N_33148,N_26891,N_26434);
xnor U33149 (N_33149,N_27077,N_26760);
and U33150 (N_33150,N_25918,N_26803);
nor U33151 (N_33151,N_26304,N_26574);
and U33152 (N_33152,N_29753,N_26445);
and U33153 (N_33153,N_27829,N_27397);
and U33154 (N_33154,N_28500,N_28334);
or U33155 (N_33155,N_25965,N_26983);
nand U33156 (N_33156,N_26401,N_25897);
or U33157 (N_33157,N_26446,N_25977);
nor U33158 (N_33158,N_29123,N_25184);
or U33159 (N_33159,N_28683,N_29378);
nand U33160 (N_33160,N_29983,N_27020);
xnor U33161 (N_33161,N_29988,N_25103);
xor U33162 (N_33162,N_27919,N_27871);
nand U33163 (N_33163,N_27181,N_29868);
and U33164 (N_33164,N_27374,N_27045);
xnor U33165 (N_33165,N_26279,N_25038);
or U33166 (N_33166,N_26661,N_29045);
or U33167 (N_33167,N_28391,N_25033);
or U33168 (N_33168,N_27149,N_26488);
and U33169 (N_33169,N_28031,N_25321);
and U33170 (N_33170,N_27717,N_26417);
xnor U33171 (N_33171,N_28351,N_28589);
or U33172 (N_33172,N_29153,N_28541);
nand U33173 (N_33173,N_26324,N_25168);
and U33174 (N_33174,N_27444,N_26844);
nand U33175 (N_33175,N_26098,N_28317);
or U33176 (N_33176,N_29211,N_28550);
xnor U33177 (N_33177,N_25910,N_25105);
nand U33178 (N_33178,N_28188,N_29246);
or U33179 (N_33179,N_25715,N_29903);
nand U33180 (N_33180,N_26704,N_25416);
nor U33181 (N_33181,N_29856,N_25413);
xor U33182 (N_33182,N_26837,N_29127);
or U33183 (N_33183,N_29350,N_26017);
and U33184 (N_33184,N_25479,N_27363);
or U33185 (N_33185,N_26174,N_27707);
nand U33186 (N_33186,N_28049,N_25376);
or U33187 (N_33187,N_27165,N_28392);
or U33188 (N_33188,N_25889,N_27739);
xnor U33189 (N_33189,N_26799,N_28640);
nand U33190 (N_33190,N_29086,N_28649);
xnor U33191 (N_33191,N_26422,N_27534);
nor U33192 (N_33192,N_29343,N_29613);
or U33193 (N_33193,N_26688,N_25052);
xnor U33194 (N_33194,N_26820,N_29923);
and U33195 (N_33195,N_27790,N_29451);
and U33196 (N_33196,N_29199,N_26237);
nand U33197 (N_33197,N_26555,N_29415);
xnor U33198 (N_33198,N_25710,N_27902);
and U33199 (N_33199,N_26914,N_26945);
and U33200 (N_33200,N_28966,N_26922);
nor U33201 (N_33201,N_29342,N_29164);
and U33202 (N_33202,N_25805,N_29350);
nor U33203 (N_33203,N_29647,N_25850);
and U33204 (N_33204,N_25727,N_28131);
xnor U33205 (N_33205,N_29955,N_28322);
xnor U33206 (N_33206,N_28155,N_27013);
xor U33207 (N_33207,N_28834,N_28674);
or U33208 (N_33208,N_29541,N_26539);
xnor U33209 (N_33209,N_28618,N_28320);
nand U33210 (N_33210,N_26091,N_29526);
or U33211 (N_33211,N_26212,N_27255);
nand U33212 (N_33212,N_25275,N_29976);
nand U33213 (N_33213,N_27407,N_29827);
or U33214 (N_33214,N_25226,N_28297);
or U33215 (N_33215,N_29509,N_26348);
and U33216 (N_33216,N_25530,N_29339);
or U33217 (N_33217,N_27937,N_29951);
or U33218 (N_33218,N_29470,N_29303);
nor U33219 (N_33219,N_29594,N_27085);
or U33220 (N_33220,N_25020,N_27697);
xor U33221 (N_33221,N_25900,N_28022);
nor U33222 (N_33222,N_28129,N_28491);
and U33223 (N_33223,N_28243,N_29798);
or U33224 (N_33224,N_28446,N_28558);
and U33225 (N_33225,N_29018,N_28463);
nor U33226 (N_33226,N_25745,N_29950);
xor U33227 (N_33227,N_26394,N_27417);
nor U33228 (N_33228,N_29084,N_25418);
and U33229 (N_33229,N_25553,N_28337);
nand U33230 (N_33230,N_26962,N_26310);
xor U33231 (N_33231,N_27443,N_26639);
nand U33232 (N_33232,N_28082,N_28415);
and U33233 (N_33233,N_26560,N_27279);
nand U33234 (N_33234,N_27182,N_26073);
nand U33235 (N_33235,N_27701,N_25048);
or U33236 (N_33236,N_26565,N_27836);
nor U33237 (N_33237,N_28059,N_28292);
nand U33238 (N_33238,N_28635,N_27342);
and U33239 (N_33239,N_29142,N_28568);
nor U33240 (N_33240,N_25962,N_25585);
nand U33241 (N_33241,N_26604,N_29566);
or U33242 (N_33242,N_25646,N_29907);
nor U33243 (N_33243,N_25503,N_29922);
nor U33244 (N_33244,N_27687,N_29092);
and U33245 (N_33245,N_29578,N_29135);
and U33246 (N_33246,N_28716,N_25766);
nor U33247 (N_33247,N_26660,N_26724);
xnor U33248 (N_33248,N_28927,N_27409);
nand U33249 (N_33249,N_26316,N_28341);
nor U33250 (N_33250,N_28619,N_29538);
xor U33251 (N_33251,N_27675,N_25798);
nor U33252 (N_33252,N_28358,N_26706);
or U33253 (N_33253,N_28259,N_26592);
or U33254 (N_33254,N_26892,N_26942);
xnor U33255 (N_33255,N_26180,N_29690);
or U33256 (N_33256,N_26166,N_28116);
and U33257 (N_33257,N_26342,N_28891);
or U33258 (N_33258,N_26332,N_26471);
or U33259 (N_33259,N_28291,N_25414);
xnor U33260 (N_33260,N_26584,N_26981);
xor U33261 (N_33261,N_27630,N_28732);
and U33262 (N_33262,N_29412,N_28730);
nor U33263 (N_33263,N_28265,N_25545);
or U33264 (N_33264,N_25667,N_25578);
and U33265 (N_33265,N_28018,N_26149);
nor U33266 (N_33266,N_25550,N_27111);
xnor U33267 (N_33267,N_26576,N_25124);
nor U33268 (N_33268,N_27660,N_27218);
and U33269 (N_33269,N_27730,N_26269);
nand U33270 (N_33270,N_29454,N_29311);
nor U33271 (N_33271,N_26669,N_25909);
nand U33272 (N_33272,N_28633,N_29020);
or U33273 (N_33273,N_28520,N_27263);
nand U33274 (N_33274,N_27234,N_27726);
or U33275 (N_33275,N_26038,N_25034);
xor U33276 (N_33276,N_25267,N_29312);
nor U33277 (N_33277,N_29679,N_29394);
or U33278 (N_33278,N_29971,N_26712);
and U33279 (N_33279,N_27436,N_28383);
nand U33280 (N_33280,N_28662,N_26023);
nand U33281 (N_33281,N_25018,N_25934);
nand U33282 (N_33282,N_25004,N_29863);
nand U33283 (N_33283,N_29267,N_27435);
nor U33284 (N_33284,N_29138,N_29036);
or U33285 (N_33285,N_26181,N_29694);
xnor U33286 (N_33286,N_28717,N_26086);
xnor U33287 (N_33287,N_27080,N_28628);
and U33288 (N_33288,N_27517,N_25980);
xnor U33289 (N_33289,N_28701,N_28028);
xor U33290 (N_33290,N_25227,N_28238);
xor U33291 (N_33291,N_27457,N_28042);
nor U33292 (N_33292,N_29446,N_27569);
nand U33293 (N_33293,N_25781,N_27034);
xor U33294 (N_33294,N_29991,N_28690);
xor U33295 (N_33295,N_27419,N_27934);
or U33296 (N_33296,N_25451,N_26800);
and U33297 (N_33297,N_29321,N_28351);
and U33298 (N_33298,N_28170,N_29200);
nand U33299 (N_33299,N_27151,N_29358);
xnor U33300 (N_33300,N_27374,N_27169);
and U33301 (N_33301,N_27211,N_26352);
or U33302 (N_33302,N_25266,N_28697);
nor U33303 (N_33303,N_27096,N_29478);
and U33304 (N_33304,N_27558,N_26137);
nand U33305 (N_33305,N_26067,N_28211);
and U33306 (N_33306,N_25176,N_25312);
or U33307 (N_33307,N_28198,N_27903);
or U33308 (N_33308,N_27152,N_29508);
and U33309 (N_33309,N_25422,N_29622);
xnor U33310 (N_33310,N_25644,N_28821);
nor U33311 (N_33311,N_25028,N_27528);
or U33312 (N_33312,N_29673,N_26391);
xnor U33313 (N_33313,N_25536,N_28842);
or U33314 (N_33314,N_28441,N_25413);
and U33315 (N_33315,N_26911,N_25595);
nand U33316 (N_33316,N_27823,N_29313);
nor U33317 (N_33317,N_26620,N_28015);
nand U33318 (N_33318,N_26007,N_28874);
nor U33319 (N_33319,N_28486,N_29069);
or U33320 (N_33320,N_27914,N_25369);
or U33321 (N_33321,N_27118,N_27454);
nand U33322 (N_33322,N_26003,N_26362);
or U33323 (N_33323,N_29154,N_27717);
nor U33324 (N_33324,N_27643,N_28127);
nor U33325 (N_33325,N_27498,N_28619);
xnor U33326 (N_33326,N_26497,N_25886);
xor U33327 (N_33327,N_29334,N_29715);
and U33328 (N_33328,N_29665,N_27232);
xor U33329 (N_33329,N_28952,N_26739);
xnor U33330 (N_33330,N_25179,N_26145);
nand U33331 (N_33331,N_26562,N_29131);
nand U33332 (N_33332,N_26426,N_28971);
or U33333 (N_33333,N_26708,N_29660);
or U33334 (N_33334,N_25687,N_29185);
or U33335 (N_33335,N_27752,N_26534);
nand U33336 (N_33336,N_29516,N_28319);
and U33337 (N_33337,N_28746,N_29630);
xor U33338 (N_33338,N_26581,N_25770);
nand U33339 (N_33339,N_26700,N_27637);
xnor U33340 (N_33340,N_29937,N_25522);
or U33341 (N_33341,N_29022,N_27498);
and U33342 (N_33342,N_27920,N_28966);
or U33343 (N_33343,N_26391,N_26929);
and U33344 (N_33344,N_27177,N_27261);
or U33345 (N_33345,N_26050,N_29167);
nand U33346 (N_33346,N_27212,N_29747);
nor U33347 (N_33347,N_28841,N_25736);
or U33348 (N_33348,N_27584,N_27836);
or U33349 (N_33349,N_27752,N_27876);
and U33350 (N_33350,N_29813,N_26479);
nor U33351 (N_33351,N_28996,N_29000);
nand U33352 (N_33352,N_26192,N_26990);
xor U33353 (N_33353,N_26086,N_29468);
xnor U33354 (N_33354,N_28387,N_25871);
nand U33355 (N_33355,N_29760,N_25764);
and U33356 (N_33356,N_26922,N_29680);
nand U33357 (N_33357,N_25587,N_29719);
nand U33358 (N_33358,N_25902,N_29384);
or U33359 (N_33359,N_28683,N_28057);
or U33360 (N_33360,N_29183,N_26459);
or U33361 (N_33361,N_27236,N_29011);
or U33362 (N_33362,N_29573,N_26376);
xnor U33363 (N_33363,N_26132,N_28402);
xor U33364 (N_33364,N_29683,N_25062);
and U33365 (N_33365,N_28808,N_25812);
and U33366 (N_33366,N_25981,N_25645);
and U33367 (N_33367,N_27912,N_25403);
nor U33368 (N_33368,N_26183,N_26374);
xor U33369 (N_33369,N_27198,N_25871);
and U33370 (N_33370,N_27298,N_26237);
nor U33371 (N_33371,N_26709,N_29373);
and U33372 (N_33372,N_25695,N_29750);
or U33373 (N_33373,N_26564,N_27611);
nand U33374 (N_33374,N_26270,N_25251);
nand U33375 (N_33375,N_27410,N_27902);
nand U33376 (N_33376,N_26066,N_28154);
xnor U33377 (N_33377,N_29937,N_27320);
and U33378 (N_33378,N_29134,N_25623);
nor U33379 (N_33379,N_25744,N_26228);
xor U33380 (N_33380,N_29002,N_25698);
nand U33381 (N_33381,N_29384,N_25418);
and U33382 (N_33382,N_27517,N_26693);
and U33383 (N_33383,N_25305,N_26607);
and U33384 (N_33384,N_28199,N_28761);
nor U33385 (N_33385,N_25299,N_26282);
or U33386 (N_33386,N_26616,N_26475);
nand U33387 (N_33387,N_26562,N_25966);
and U33388 (N_33388,N_28175,N_27000);
nor U33389 (N_33389,N_27732,N_26800);
nor U33390 (N_33390,N_25145,N_29391);
xnor U33391 (N_33391,N_29836,N_25311);
nand U33392 (N_33392,N_29017,N_26183);
nand U33393 (N_33393,N_29932,N_26020);
xor U33394 (N_33394,N_28015,N_26519);
and U33395 (N_33395,N_26702,N_25837);
xnor U33396 (N_33396,N_28184,N_25219);
or U33397 (N_33397,N_29420,N_28348);
and U33398 (N_33398,N_25629,N_28174);
nor U33399 (N_33399,N_26805,N_26776);
xor U33400 (N_33400,N_27241,N_28788);
or U33401 (N_33401,N_28246,N_27506);
xor U33402 (N_33402,N_25232,N_26065);
and U33403 (N_33403,N_29693,N_26418);
or U33404 (N_33404,N_25475,N_26879);
nand U33405 (N_33405,N_28833,N_26290);
or U33406 (N_33406,N_27640,N_28304);
nor U33407 (N_33407,N_25352,N_25812);
and U33408 (N_33408,N_25772,N_28734);
nand U33409 (N_33409,N_26077,N_27901);
nor U33410 (N_33410,N_28609,N_25475);
xnor U33411 (N_33411,N_25860,N_29372);
or U33412 (N_33412,N_26362,N_27461);
and U33413 (N_33413,N_29165,N_26049);
nand U33414 (N_33414,N_25564,N_28290);
nand U33415 (N_33415,N_29180,N_25799);
or U33416 (N_33416,N_27663,N_29291);
or U33417 (N_33417,N_29921,N_28495);
nor U33418 (N_33418,N_27361,N_25647);
xnor U33419 (N_33419,N_27017,N_26732);
or U33420 (N_33420,N_26800,N_26216);
nand U33421 (N_33421,N_27247,N_26686);
nor U33422 (N_33422,N_26284,N_26732);
and U33423 (N_33423,N_29473,N_28098);
nor U33424 (N_33424,N_26059,N_26013);
nor U33425 (N_33425,N_26594,N_25864);
xor U33426 (N_33426,N_27280,N_26852);
or U33427 (N_33427,N_29904,N_28154);
nand U33428 (N_33428,N_27700,N_26920);
nand U33429 (N_33429,N_29935,N_28482);
nor U33430 (N_33430,N_29130,N_26813);
and U33431 (N_33431,N_26159,N_26941);
and U33432 (N_33432,N_27735,N_26187);
nor U33433 (N_33433,N_28413,N_27670);
and U33434 (N_33434,N_26453,N_29869);
xor U33435 (N_33435,N_27975,N_27322);
nor U33436 (N_33436,N_27166,N_25486);
nand U33437 (N_33437,N_25989,N_28959);
or U33438 (N_33438,N_29227,N_25031);
or U33439 (N_33439,N_25836,N_29491);
xnor U33440 (N_33440,N_26770,N_26712);
and U33441 (N_33441,N_27446,N_29595);
and U33442 (N_33442,N_29897,N_29041);
and U33443 (N_33443,N_27426,N_27512);
nor U33444 (N_33444,N_25485,N_29400);
nand U33445 (N_33445,N_27812,N_27544);
nand U33446 (N_33446,N_25142,N_28056);
nor U33447 (N_33447,N_26515,N_29172);
and U33448 (N_33448,N_28174,N_29812);
or U33449 (N_33449,N_25317,N_26213);
nor U33450 (N_33450,N_28376,N_29483);
nor U33451 (N_33451,N_29243,N_29020);
and U33452 (N_33452,N_28909,N_25001);
nor U33453 (N_33453,N_29441,N_28333);
xnor U33454 (N_33454,N_29546,N_28394);
nand U33455 (N_33455,N_28938,N_29972);
or U33456 (N_33456,N_27018,N_29121);
xnor U33457 (N_33457,N_25621,N_25564);
or U33458 (N_33458,N_26974,N_26969);
xnor U33459 (N_33459,N_28941,N_25112);
and U33460 (N_33460,N_27518,N_26646);
and U33461 (N_33461,N_29910,N_28681);
nor U33462 (N_33462,N_27000,N_25534);
nand U33463 (N_33463,N_27935,N_28900);
and U33464 (N_33464,N_29900,N_27426);
or U33465 (N_33465,N_28613,N_26515);
and U33466 (N_33466,N_26322,N_25876);
and U33467 (N_33467,N_25179,N_29985);
or U33468 (N_33468,N_29730,N_29245);
nand U33469 (N_33469,N_25621,N_29266);
or U33470 (N_33470,N_29941,N_27070);
xnor U33471 (N_33471,N_28701,N_26977);
nand U33472 (N_33472,N_27032,N_27057);
nor U33473 (N_33473,N_25795,N_28969);
and U33474 (N_33474,N_27585,N_25878);
nand U33475 (N_33475,N_26702,N_28037);
xnor U33476 (N_33476,N_27210,N_29920);
or U33477 (N_33477,N_26267,N_28375);
nor U33478 (N_33478,N_25200,N_28984);
nand U33479 (N_33479,N_29933,N_28439);
or U33480 (N_33480,N_26262,N_29655);
nand U33481 (N_33481,N_28021,N_25951);
or U33482 (N_33482,N_25506,N_28293);
xor U33483 (N_33483,N_25330,N_26434);
xnor U33484 (N_33484,N_25748,N_27474);
nor U33485 (N_33485,N_26104,N_27319);
xnor U33486 (N_33486,N_26200,N_25975);
nor U33487 (N_33487,N_29754,N_25849);
nand U33488 (N_33488,N_25471,N_28969);
and U33489 (N_33489,N_27089,N_27249);
nand U33490 (N_33490,N_28929,N_25143);
and U33491 (N_33491,N_26973,N_27732);
or U33492 (N_33492,N_26080,N_29293);
nor U33493 (N_33493,N_25845,N_28105);
nor U33494 (N_33494,N_25759,N_25854);
nor U33495 (N_33495,N_25773,N_26138);
and U33496 (N_33496,N_29156,N_29471);
nor U33497 (N_33497,N_26630,N_27077);
and U33498 (N_33498,N_28927,N_25252);
or U33499 (N_33499,N_26671,N_25837);
nand U33500 (N_33500,N_28634,N_26205);
and U33501 (N_33501,N_25765,N_28283);
xor U33502 (N_33502,N_25197,N_27998);
and U33503 (N_33503,N_26460,N_28585);
nor U33504 (N_33504,N_28408,N_28486);
nand U33505 (N_33505,N_27567,N_25402);
or U33506 (N_33506,N_27725,N_29887);
nand U33507 (N_33507,N_27270,N_25884);
nor U33508 (N_33508,N_26489,N_28327);
and U33509 (N_33509,N_29151,N_25207);
xnor U33510 (N_33510,N_27885,N_25224);
or U33511 (N_33511,N_29103,N_26386);
and U33512 (N_33512,N_25383,N_25528);
or U33513 (N_33513,N_27280,N_28975);
nand U33514 (N_33514,N_28699,N_27918);
or U33515 (N_33515,N_25833,N_26801);
nor U33516 (N_33516,N_25975,N_25383);
xnor U33517 (N_33517,N_25764,N_27348);
nand U33518 (N_33518,N_25932,N_27112);
nand U33519 (N_33519,N_28751,N_27256);
nand U33520 (N_33520,N_25518,N_28473);
xor U33521 (N_33521,N_25370,N_29661);
xor U33522 (N_33522,N_25246,N_29357);
xor U33523 (N_33523,N_28346,N_28265);
nand U33524 (N_33524,N_26949,N_29400);
and U33525 (N_33525,N_28775,N_28752);
and U33526 (N_33526,N_26774,N_29326);
and U33527 (N_33527,N_29500,N_25186);
and U33528 (N_33528,N_29704,N_28299);
and U33529 (N_33529,N_27337,N_29796);
or U33530 (N_33530,N_25394,N_29366);
nand U33531 (N_33531,N_29265,N_27551);
xnor U33532 (N_33532,N_28702,N_28557);
nor U33533 (N_33533,N_25050,N_27859);
nor U33534 (N_33534,N_26372,N_28934);
xnor U33535 (N_33535,N_27809,N_29380);
nand U33536 (N_33536,N_29856,N_28982);
or U33537 (N_33537,N_25888,N_29865);
xor U33538 (N_33538,N_26224,N_26867);
or U33539 (N_33539,N_26208,N_26554);
nor U33540 (N_33540,N_26889,N_25629);
or U33541 (N_33541,N_26563,N_25847);
and U33542 (N_33542,N_29658,N_25534);
and U33543 (N_33543,N_27091,N_25896);
and U33544 (N_33544,N_28296,N_26240);
or U33545 (N_33545,N_26298,N_29687);
and U33546 (N_33546,N_29450,N_25983);
nand U33547 (N_33547,N_27567,N_28563);
nand U33548 (N_33548,N_29914,N_28896);
or U33549 (N_33549,N_28160,N_25052);
xor U33550 (N_33550,N_28555,N_25402);
nand U33551 (N_33551,N_27973,N_25945);
or U33552 (N_33552,N_29404,N_28880);
or U33553 (N_33553,N_28597,N_28366);
nor U33554 (N_33554,N_27383,N_26994);
or U33555 (N_33555,N_25507,N_29412);
and U33556 (N_33556,N_27872,N_27137);
and U33557 (N_33557,N_28786,N_28231);
and U33558 (N_33558,N_25797,N_27448);
nand U33559 (N_33559,N_27811,N_28530);
or U33560 (N_33560,N_26466,N_26339);
nor U33561 (N_33561,N_25309,N_26781);
nand U33562 (N_33562,N_28527,N_26459);
xnor U33563 (N_33563,N_29203,N_27888);
or U33564 (N_33564,N_29184,N_29310);
nand U33565 (N_33565,N_26701,N_25771);
nand U33566 (N_33566,N_27783,N_27538);
xor U33567 (N_33567,N_26293,N_26506);
or U33568 (N_33568,N_26819,N_28896);
xnor U33569 (N_33569,N_27396,N_26249);
nand U33570 (N_33570,N_27954,N_25838);
or U33571 (N_33571,N_25560,N_27655);
xor U33572 (N_33572,N_28864,N_26467);
nand U33573 (N_33573,N_25493,N_26234);
and U33574 (N_33574,N_27322,N_28184);
nand U33575 (N_33575,N_25402,N_25144);
and U33576 (N_33576,N_28820,N_25306);
and U33577 (N_33577,N_27695,N_27558);
nor U33578 (N_33578,N_26237,N_26226);
xnor U33579 (N_33579,N_26417,N_26750);
nand U33580 (N_33580,N_28128,N_26976);
nor U33581 (N_33581,N_29321,N_26452);
xor U33582 (N_33582,N_25484,N_26303);
and U33583 (N_33583,N_28875,N_26307);
xor U33584 (N_33584,N_29959,N_26562);
nor U33585 (N_33585,N_26458,N_28760);
nand U33586 (N_33586,N_29693,N_25087);
xor U33587 (N_33587,N_25201,N_27507);
nand U33588 (N_33588,N_25232,N_27885);
nor U33589 (N_33589,N_27612,N_29301);
nand U33590 (N_33590,N_27814,N_25835);
and U33591 (N_33591,N_28188,N_26543);
nor U33592 (N_33592,N_25949,N_25728);
xnor U33593 (N_33593,N_27035,N_29067);
or U33594 (N_33594,N_26693,N_26244);
xor U33595 (N_33595,N_25755,N_29071);
nand U33596 (N_33596,N_25599,N_27351);
xor U33597 (N_33597,N_29586,N_29218);
nand U33598 (N_33598,N_29400,N_28110);
nor U33599 (N_33599,N_29358,N_28210);
or U33600 (N_33600,N_29423,N_25206);
or U33601 (N_33601,N_28664,N_29423);
xnor U33602 (N_33602,N_26847,N_27968);
or U33603 (N_33603,N_25046,N_26001);
or U33604 (N_33604,N_25182,N_28392);
nor U33605 (N_33605,N_27765,N_29505);
xnor U33606 (N_33606,N_25525,N_29612);
or U33607 (N_33607,N_26694,N_29401);
nand U33608 (N_33608,N_29230,N_27966);
nor U33609 (N_33609,N_29639,N_29121);
or U33610 (N_33610,N_28827,N_26016);
or U33611 (N_33611,N_27751,N_27630);
nor U33612 (N_33612,N_29910,N_25994);
or U33613 (N_33613,N_29842,N_28846);
xor U33614 (N_33614,N_25389,N_25139);
or U33615 (N_33615,N_29281,N_26836);
xnor U33616 (N_33616,N_29472,N_26829);
or U33617 (N_33617,N_29698,N_29429);
and U33618 (N_33618,N_28289,N_25529);
xor U33619 (N_33619,N_25785,N_29074);
or U33620 (N_33620,N_26160,N_26346);
nand U33621 (N_33621,N_26292,N_27699);
and U33622 (N_33622,N_29527,N_27536);
or U33623 (N_33623,N_28832,N_27812);
nor U33624 (N_33624,N_25917,N_28248);
xor U33625 (N_33625,N_29617,N_29116);
and U33626 (N_33626,N_27115,N_25885);
nor U33627 (N_33627,N_27030,N_25679);
nor U33628 (N_33628,N_25856,N_27263);
nor U33629 (N_33629,N_26389,N_25952);
or U33630 (N_33630,N_28900,N_26665);
nor U33631 (N_33631,N_26268,N_27798);
nor U33632 (N_33632,N_29272,N_26008);
and U33633 (N_33633,N_29660,N_29514);
nand U33634 (N_33634,N_29110,N_28224);
nand U33635 (N_33635,N_29907,N_29878);
nand U33636 (N_33636,N_25777,N_26384);
nand U33637 (N_33637,N_27753,N_27929);
nor U33638 (N_33638,N_27558,N_25215);
nor U33639 (N_33639,N_25756,N_29451);
or U33640 (N_33640,N_29386,N_27675);
nand U33641 (N_33641,N_29906,N_25505);
or U33642 (N_33642,N_25223,N_29369);
and U33643 (N_33643,N_29337,N_28583);
and U33644 (N_33644,N_27449,N_26791);
xnor U33645 (N_33645,N_27116,N_27760);
nand U33646 (N_33646,N_25928,N_25733);
or U33647 (N_33647,N_27120,N_26811);
nand U33648 (N_33648,N_27941,N_26033);
and U33649 (N_33649,N_28514,N_28052);
or U33650 (N_33650,N_26068,N_26931);
and U33651 (N_33651,N_28717,N_25491);
and U33652 (N_33652,N_27528,N_29491);
or U33653 (N_33653,N_27578,N_25453);
and U33654 (N_33654,N_28882,N_27931);
nor U33655 (N_33655,N_26086,N_26404);
or U33656 (N_33656,N_29350,N_28194);
or U33657 (N_33657,N_26547,N_27163);
nor U33658 (N_33658,N_27320,N_28449);
nand U33659 (N_33659,N_25865,N_27262);
or U33660 (N_33660,N_29354,N_28054);
nand U33661 (N_33661,N_25307,N_28849);
and U33662 (N_33662,N_28212,N_29039);
nor U33663 (N_33663,N_28464,N_27366);
nor U33664 (N_33664,N_26752,N_29484);
nor U33665 (N_33665,N_27960,N_29634);
or U33666 (N_33666,N_27453,N_25561);
xor U33667 (N_33667,N_26127,N_26205);
or U33668 (N_33668,N_28416,N_29069);
xnor U33669 (N_33669,N_28074,N_29173);
or U33670 (N_33670,N_28195,N_29782);
nor U33671 (N_33671,N_28348,N_25652);
nand U33672 (N_33672,N_25601,N_29283);
nand U33673 (N_33673,N_29042,N_29909);
or U33674 (N_33674,N_28808,N_28846);
or U33675 (N_33675,N_28362,N_27806);
xor U33676 (N_33676,N_27086,N_29846);
and U33677 (N_33677,N_27248,N_25375);
nor U33678 (N_33678,N_28293,N_27976);
nor U33679 (N_33679,N_25529,N_29046);
nand U33680 (N_33680,N_29452,N_26716);
xor U33681 (N_33681,N_26840,N_25378);
xor U33682 (N_33682,N_26764,N_28307);
and U33683 (N_33683,N_27268,N_25421);
and U33684 (N_33684,N_28577,N_29316);
nand U33685 (N_33685,N_28957,N_29832);
nor U33686 (N_33686,N_28526,N_28380);
and U33687 (N_33687,N_29062,N_29697);
nor U33688 (N_33688,N_29741,N_25829);
or U33689 (N_33689,N_25535,N_26620);
and U33690 (N_33690,N_26973,N_28569);
nor U33691 (N_33691,N_25083,N_29490);
xnor U33692 (N_33692,N_28402,N_26270);
xnor U33693 (N_33693,N_25235,N_29465);
xor U33694 (N_33694,N_28871,N_28741);
xor U33695 (N_33695,N_29860,N_28322);
nor U33696 (N_33696,N_29806,N_27804);
xor U33697 (N_33697,N_27538,N_27773);
nand U33698 (N_33698,N_29514,N_27461);
xor U33699 (N_33699,N_27623,N_28381);
nand U33700 (N_33700,N_26895,N_26343);
or U33701 (N_33701,N_26956,N_28268);
nand U33702 (N_33702,N_26904,N_28089);
nor U33703 (N_33703,N_27575,N_26713);
and U33704 (N_33704,N_25519,N_26067);
nor U33705 (N_33705,N_25925,N_27859);
nor U33706 (N_33706,N_29517,N_29466);
nor U33707 (N_33707,N_28536,N_28046);
xor U33708 (N_33708,N_26769,N_27377);
xor U33709 (N_33709,N_27159,N_28358);
nor U33710 (N_33710,N_26907,N_26772);
xnor U33711 (N_33711,N_25052,N_26905);
nand U33712 (N_33712,N_27375,N_25345);
or U33713 (N_33713,N_29360,N_27538);
xnor U33714 (N_33714,N_29600,N_29952);
nor U33715 (N_33715,N_26589,N_29650);
xnor U33716 (N_33716,N_27273,N_26680);
or U33717 (N_33717,N_26970,N_27064);
xnor U33718 (N_33718,N_27332,N_25602);
and U33719 (N_33719,N_27245,N_28619);
nand U33720 (N_33720,N_28653,N_27697);
or U33721 (N_33721,N_25923,N_29296);
xor U33722 (N_33722,N_29141,N_26478);
and U33723 (N_33723,N_26658,N_29007);
and U33724 (N_33724,N_29678,N_29321);
nor U33725 (N_33725,N_25926,N_27846);
xnor U33726 (N_33726,N_29629,N_25254);
or U33727 (N_33727,N_28511,N_26245);
and U33728 (N_33728,N_27482,N_25112);
nor U33729 (N_33729,N_26556,N_27834);
nor U33730 (N_33730,N_28142,N_27116);
and U33731 (N_33731,N_28071,N_28028);
and U33732 (N_33732,N_29203,N_26885);
and U33733 (N_33733,N_25310,N_26511);
nand U33734 (N_33734,N_27561,N_28368);
nand U33735 (N_33735,N_28747,N_25500);
or U33736 (N_33736,N_26596,N_28938);
and U33737 (N_33737,N_28740,N_25896);
and U33738 (N_33738,N_27514,N_25507);
or U33739 (N_33739,N_28169,N_26473);
nor U33740 (N_33740,N_29474,N_27236);
or U33741 (N_33741,N_29415,N_28233);
xor U33742 (N_33742,N_26421,N_28030);
and U33743 (N_33743,N_27902,N_27690);
xor U33744 (N_33744,N_28801,N_26256);
nor U33745 (N_33745,N_28536,N_25294);
nor U33746 (N_33746,N_29001,N_26912);
or U33747 (N_33747,N_25591,N_27753);
nand U33748 (N_33748,N_25523,N_27189);
or U33749 (N_33749,N_29531,N_26273);
xor U33750 (N_33750,N_25239,N_29130);
nor U33751 (N_33751,N_29124,N_26078);
or U33752 (N_33752,N_29006,N_27460);
and U33753 (N_33753,N_28651,N_28579);
xnor U33754 (N_33754,N_28961,N_25837);
or U33755 (N_33755,N_25079,N_29937);
xnor U33756 (N_33756,N_28430,N_29784);
nand U33757 (N_33757,N_27924,N_26623);
nand U33758 (N_33758,N_25771,N_26707);
nand U33759 (N_33759,N_29167,N_26461);
nor U33760 (N_33760,N_29430,N_25274);
and U33761 (N_33761,N_25775,N_26151);
nor U33762 (N_33762,N_28716,N_26171);
xnor U33763 (N_33763,N_26524,N_26858);
xnor U33764 (N_33764,N_28713,N_29452);
or U33765 (N_33765,N_29924,N_29121);
and U33766 (N_33766,N_28181,N_29392);
or U33767 (N_33767,N_29606,N_28977);
nor U33768 (N_33768,N_29379,N_25744);
xnor U33769 (N_33769,N_29962,N_29631);
xnor U33770 (N_33770,N_27744,N_25938);
nand U33771 (N_33771,N_26470,N_27531);
or U33772 (N_33772,N_28305,N_27877);
and U33773 (N_33773,N_25455,N_26212);
nor U33774 (N_33774,N_28342,N_26322);
or U33775 (N_33775,N_29051,N_29303);
nand U33776 (N_33776,N_29178,N_26896);
xnor U33777 (N_33777,N_27626,N_26976);
nand U33778 (N_33778,N_25632,N_29098);
nor U33779 (N_33779,N_25422,N_25902);
xnor U33780 (N_33780,N_25564,N_28664);
or U33781 (N_33781,N_25329,N_28108);
xnor U33782 (N_33782,N_29366,N_27670);
or U33783 (N_33783,N_25705,N_29944);
or U33784 (N_33784,N_25184,N_29468);
nor U33785 (N_33785,N_27264,N_29168);
and U33786 (N_33786,N_27803,N_29104);
nor U33787 (N_33787,N_27504,N_26838);
xor U33788 (N_33788,N_29848,N_25867);
or U33789 (N_33789,N_26179,N_25797);
nand U33790 (N_33790,N_25617,N_25180);
xnor U33791 (N_33791,N_28661,N_26075);
nor U33792 (N_33792,N_29161,N_29014);
nor U33793 (N_33793,N_29361,N_29038);
and U33794 (N_33794,N_25571,N_26734);
nor U33795 (N_33795,N_25767,N_26364);
and U33796 (N_33796,N_28430,N_28192);
nand U33797 (N_33797,N_27551,N_28030);
and U33798 (N_33798,N_27270,N_29962);
xnor U33799 (N_33799,N_26371,N_26636);
nand U33800 (N_33800,N_29968,N_25183);
or U33801 (N_33801,N_25745,N_29255);
and U33802 (N_33802,N_27772,N_28216);
nand U33803 (N_33803,N_27927,N_29058);
nand U33804 (N_33804,N_27282,N_29418);
nor U33805 (N_33805,N_28580,N_26994);
nor U33806 (N_33806,N_29988,N_29586);
nor U33807 (N_33807,N_29074,N_25043);
or U33808 (N_33808,N_26816,N_26198);
xor U33809 (N_33809,N_28212,N_26236);
or U33810 (N_33810,N_28075,N_26668);
nand U33811 (N_33811,N_25081,N_29321);
and U33812 (N_33812,N_26786,N_25151);
and U33813 (N_33813,N_25981,N_26323);
or U33814 (N_33814,N_29517,N_27354);
and U33815 (N_33815,N_28184,N_29799);
xor U33816 (N_33816,N_25571,N_26347);
xnor U33817 (N_33817,N_25815,N_26704);
nor U33818 (N_33818,N_25963,N_28229);
or U33819 (N_33819,N_27055,N_29606);
nand U33820 (N_33820,N_25688,N_26950);
and U33821 (N_33821,N_27494,N_25151);
nor U33822 (N_33822,N_27005,N_28051);
xor U33823 (N_33823,N_26879,N_26444);
nand U33824 (N_33824,N_28222,N_29143);
nand U33825 (N_33825,N_25804,N_28720);
and U33826 (N_33826,N_29242,N_26655);
xnor U33827 (N_33827,N_28011,N_28481);
nor U33828 (N_33828,N_29783,N_28669);
and U33829 (N_33829,N_26810,N_26051);
and U33830 (N_33830,N_25471,N_27295);
nor U33831 (N_33831,N_28893,N_25604);
nand U33832 (N_33832,N_29021,N_25700);
or U33833 (N_33833,N_26465,N_29831);
nand U33834 (N_33834,N_26381,N_26971);
nand U33835 (N_33835,N_28816,N_26044);
nor U33836 (N_33836,N_28769,N_25614);
xor U33837 (N_33837,N_29714,N_26332);
and U33838 (N_33838,N_28754,N_29876);
and U33839 (N_33839,N_28433,N_25575);
nand U33840 (N_33840,N_29839,N_28296);
and U33841 (N_33841,N_28896,N_27806);
nand U33842 (N_33842,N_26116,N_27982);
nor U33843 (N_33843,N_28900,N_27043);
or U33844 (N_33844,N_28773,N_25834);
nor U33845 (N_33845,N_26679,N_29100);
nand U33846 (N_33846,N_29856,N_27003);
and U33847 (N_33847,N_26898,N_25294);
and U33848 (N_33848,N_29102,N_27594);
nand U33849 (N_33849,N_27456,N_25234);
xnor U33850 (N_33850,N_29506,N_28722);
xnor U33851 (N_33851,N_29064,N_28618);
nor U33852 (N_33852,N_27806,N_29964);
nand U33853 (N_33853,N_28951,N_27947);
nand U33854 (N_33854,N_26944,N_27411);
or U33855 (N_33855,N_28938,N_27702);
nand U33856 (N_33856,N_29402,N_28391);
or U33857 (N_33857,N_25771,N_26909);
nand U33858 (N_33858,N_27743,N_26691);
nand U33859 (N_33859,N_26780,N_28240);
and U33860 (N_33860,N_27891,N_27479);
nand U33861 (N_33861,N_25979,N_28162);
xnor U33862 (N_33862,N_29738,N_26567);
nand U33863 (N_33863,N_27017,N_27889);
and U33864 (N_33864,N_28042,N_28089);
nand U33865 (N_33865,N_27915,N_27726);
nand U33866 (N_33866,N_27761,N_28228);
and U33867 (N_33867,N_25168,N_25271);
or U33868 (N_33868,N_25108,N_25300);
or U33869 (N_33869,N_26103,N_28100);
xor U33870 (N_33870,N_27314,N_25343);
and U33871 (N_33871,N_29393,N_26904);
xor U33872 (N_33872,N_28887,N_29908);
nand U33873 (N_33873,N_25340,N_25807);
and U33874 (N_33874,N_26034,N_29385);
xnor U33875 (N_33875,N_28463,N_25796);
or U33876 (N_33876,N_29905,N_26504);
or U33877 (N_33877,N_27886,N_28639);
xor U33878 (N_33878,N_27425,N_29141);
and U33879 (N_33879,N_25199,N_28482);
or U33880 (N_33880,N_29124,N_25670);
xnor U33881 (N_33881,N_28971,N_27498);
nor U33882 (N_33882,N_29320,N_26011);
and U33883 (N_33883,N_27845,N_27491);
nor U33884 (N_33884,N_26301,N_27061);
and U33885 (N_33885,N_26729,N_25381);
nor U33886 (N_33886,N_26683,N_26776);
or U33887 (N_33887,N_26995,N_27712);
and U33888 (N_33888,N_26644,N_27943);
xnor U33889 (N_33889,N_29926,N_29542);
nand U33890 (N_33890,N_27556,N_25528);
nor U33891 (N_33891,N_25482,N_27240);
and U33892 (N_33892,N_27641,N_28276);
nor U33893 (N_33893,N_26897,N_26223);
or U33894 (N_33894,N_25182,N_26788);
and U33895 (N_33895,N_28847,N_25089);
nor U33896 (N_33896,N_26488,N_29767);
nor U33897 (N_33897,N_27643,N_28426);
nor U33898 (N_33898,N_26992,N_27660);
or U33899 (N_33899,N_25334,N_25508);
or U33900 (N_33900,N_28252,N_27146);
xor U33901 (N_33901,N_26081,N_28833);
nand U33902 (N_33902,N_25521,N_29075);
or U33903 (N_33903,N_29791,N_27007);
xor U33904 (N_33904,N_25894,N_29176);
xnor U33905 (N_33905,N_26083,N_28867);
or U33906 (N_33906,N_25663,N_28849);
or U33907 (N_33907,N_29120,N_25828);
or U33908 (N_33908,N_28798,N_28318);
and U33909 (N_33909,N_26157,N_26742);
nor U33910 (N_33910,N_27900,N_29079);
nor U33911 (N_33911,N_25571,N_29252);
nand U33912 (N_33912,N_27726,N_28676);
nand U33913 (N_33913,N_27077,N_27500);
and U33914 (N_33914,N_28592,N_26651);
or U33915 (N_33915,N_27939,N_25900);
nand U33916 (N_33916,N_29500,N_27319);
or U33917 (N_33917,N_25752,N_27855);
or U33918 (N_33918,N_25206,N_28985);
nand U33919 (N_33919,N_28195,N_29469);
xnor U33920 (N_33920,N_29172,N_29030);
nor U33921 (N_33921,N_29137,N_29425);
or U33922 (N_33922,N_28325,N_26836);
and U33923 (N_33923,N_29537,N_28653);
and U33924 (N_33924,N_29354,N_26495);
nand U33925 (N_33925,N_29890,N_28939);
or U33926 (N_33926,N_25910,N_25654);
xor U33927 (N_33927,N_29964,N_26143);
nand U33928 (N_33928,N_27701,N_25736);
xor U33929 (N_33929,N_25972,N_29512);
nand U33930 (N_33930,N_28324,N_27962);
xnor U33931 (N_33931,N_28034,N_25989);
or U33932 (N_33932,N_26254,N_29437);
and U33933 (N_33933,N_28770,N_27355);
xor U33934 (N_33934,N_28596,N_26239);
or U33935 (N_33935,N_27822,N_28463);
or U33936 (N_33936,N_28459,N_29033);
nor U33937 (N_33937,N_28191,N_28939);
nor U33938 (N_33938,N_27621,N_29330);
or U33939 (N_33939,N_28139,N_25326);
nor U33940 (N_33940,N_27965,N_27041);
or U33941 (N_33941,N_27623,N_27962);
nand U33942 (N_33942,N_26524,N_25300);
nor U33943 (N_33943,N_26748,N_26843);
or U33944 (N_33944,N_29053,N_26667);
and U33945 (N_33945,N_28225,N_29088);
xor U33946 (N_33946,N_29972,N_29266);
nor U33947 (N_33947,N_27701,N_26117);
or U33948 (N_33948,N_25088,N_25316);
xnor U33949 (N_33949,N_25839,N_29418);
or U33950 (N_33950,N_28964,N_27460);
xnor U33951 (N_33951,N_28598,N_29146);
nor U33952 (N_33952,N_25976,N_27174);
and U33953 (N_33953,N_27360,N_28725);
nor U33954 (N_33954,N_25365,N_25546);
nor U33955 (N_33955,N_28049,N_25480);
xor U33956 (N_33956,N_26141,N_26016);
nor U33957 (N_33957,N_26785,N_29582);
and U33958 (N_33958,N_27950,N_29547);
nor U33959 (N_33959,N_28800,N_26349);
and U33960 (N_33960,N_26848,N_28302);
or U33961 (N_33961,N_25247,N_25654);
or U33962 (N_33962,N_28899,N_25585);
nor U33963 (N_33963,N_26930,N_29417);
nor U33964 (N_33964,N_25156,N_27110);
nor U33965 (N_33965,N_25537,N_28893);
nand U33966 (N_33966,N_27007,N_29312);
or U33967 (N_33967,N_28434,N_26599);
or U33968 (N_33968,N_29014,N_27756);
or U33969 (N_33969,N_25298,N_25794);
xnor U33970 (N_33970,N_27842,N_25111);
nand U33971 (N_33971,N_26792,N_26650);
or U33972 (N_33972,N_28367,N_28449);
xnor U33973 (N_33973,N_27792,N_27986);
or U33974 (N_33974,N_29507,N_28590);
or U33975 (N_33975,N_27998,N_26400);
and U33976 (N_33976,N_28712,N_27535);
nand U33977 (N_33977,N_25328,N_26390);
xor U33978 (N_33978,N_27785,N_25914);
nor U33979 (N_33979,N_25729,N_25972);
nor U33980 (N_33980,N_26072,N_26728);
nor U33981 (N_33981,N_29602,N_26094);
xor U33982 (N_33982,N_27677,N_25627);
and U33983 (N_33983,N_28350,N_28735);
and U33984 (N_33984,N_29696,N_27234);
xnor U33985 (N_33985,N_29302,N_27806);
nor U33986 (N_33986,N_25962,N_25193);
and U33987 (N_33987,N_26013,N_25047);
nor U33988 (N_33988,N_26386,N_27572);
xor U33989 (N_33989,N_26273,N_28671);
or U33990 (N_33990,N_28068,N_25546);
nor U33991 (N_33991,N_25270,N_28579);
nand U33992 (N_33992,N_27147,N_28746);
nor U33993 (N_33993,N_27796,N_27545);
nor U33994 (N_33994,N_25500,N_26748);
xnor U33995 (N_33995,N_26214,N_29100);
xor U33996 (N_33996,N_27515,N_27750);
xor U33997 (N_33997,N_28839,N_25508);
nor U33998 (N_33998,N_29982,N_29324);
or U33999 (N_33999,N_29976,N_28280);
or U34000 (N_34000,N_28197,N_29189);
or U34001 (N_34001,N_25606,N_26451);
or U34002 (N_34002,N_25284,N_25910);
nor U34003 (N_34003,N_27363,N_26182);
or U34004 (N_34004,N_29376,N_28344);
and U34005 (N_34005,N_27489,N_25297);
nor U34006 (N_34006,N_28837,N_29391);
xnor U34007 (N_34007,N_26432,N_27323);
xor U34008 (N_34008,N_27578,N_26923);
or U34009 (N_34009,N_29469,N_26096);
xor U34010 (N_34010,N_25573,N_26799);
and U34011 (N_34011,N_25664,N_27528);
nand U34012 (N_34012,N_27322,N_28748);
nand U34013 (N_34013,N_27108,N_26887);
nor U34014 (N_34014,N_28212,N_28319);
nor U34015 (N_34015,N_26068,N_28598);
nor U34016 (N_34016,N_27745,N_29610);
or U34017 (N_34017,N_26447,N_25366);
and U34018 (N_34018,N_29719,N_25224);
nor U34019 (N_34019,N_26939,N_28175);
nor U34020 (N_34020,N_28004,N_28942);
or U34021 (N_34021,N_25411,N_25776);
or U34022 (N_34022,N_25544,N_26760);
nor U34023 (N_34023,N_28047,N_29025);
nand U34024 (N_34024,N_25924,N_25945);
or U34025 (N_34025,N_28186,N_26063);
nand U34026 (N_34026,N_27221,N_26644);
nand U34027 (N_34027,N_25478,N_29874);
nor U34028 (N_34028,N_26845,N_25535);
or U34029 (N_34029,N_29316,N_25696);
nor U34030 (N_34030,N_25275,N_26068);
nor U34031 (N_34031,N_27471,N_25808);
and U34032 (N_34032,N_27809,N_29093);
nand U34033 (N_34033,N_28249,N_25135);
xnor U34034 (N_34034,N_29606,N_29781);
xnor U34035 (N_34035,N_28953,N_27850);
and U34036 (N_34036,N_27994,N_29282);
nor U34037 (N_34037,N_28558,N_25456);
nor U34038 (N_34038,N_26590,N_28188);
xnor U34039 (N_34039,N_28580,N_26868);
or U34040 (N_34040,N_29860,N_29385);
and U34041 (N_34041,N_26586,N_29919);
nor U34042 (N_34042,N_27230,N_29422);
xor U34043 (N_34043,N_29458,N_28966);
and U34044 (N_34044,N_26332,N_25462);
nand U34045 (N_34045,N_26294,N_29900);
and U34046 (N_34046,N_27116,N_29302);
nand U34047 (N_34047,N_28703,N_25340);
and U34048 (N_34048,N_26015,N_28718);
xnor U34049 (N_34049,N_29797,N_25378);
and U34050 (N_34050,N_28478,N_25065);
xor U34051 (N_34051,N_29155,N_28276);
nor U34052 (N_34052,N_27340,N_28143);
xor U34053 (N_34053,N_29801,N_28495);
xnor U34054 (N_34054,N_29614,N_28077);
and U34055 (N_34055,N_26746,N_26638);
or U34056 (N_34056,N_29880,N_27883);
and U34057 (N_34057,N_29425,N_27375);
nand U34058 (N_34058,N_29892,N_25600);
and U34059 (N_34059,N_28416,N_25359);
or U34060 (N_34060,N_29715,N_26050);
or U34061 (N_34061,N_25676,N_29783);
and U34062 (N_34062,N_27115,N_29915);
nor U34063 (N_34063,N_29089,N_27177);
nand U34064 (N_34064,N_28382,N_27759);
and U34065 (N_34065,N_28724,N_27789);
nor U34066 (N_34066,N_26997,N_26268);
or U34067 (N_34067,N_25121,N_29618);
and U34068 (N_34068,N_28451,N_27260);
nand U34069 (N_34069,N_26401,N_25535);
or U34070 (N_34070,N_27773,N_29806);
or U34071 (N_34071,N_29490,N_27701);
or U34072 (N_34072,N_26646,N_28792);
and U34073 (N_34073,N_27297,N_28175);
or U34074 (N_34074,N_28583,N_26344);
nor U34075 (N_34075,N_25399,N_27327);
nor U34076 (N_34076,N_28016,N_26513);
nand U34077 (N_34077,N_27016,N_29195);
nor U34078 (N_34078,N_28102,N_27889);
and U34079 (N_34079,N_28074,N_27006);
nor U34080 (N_34080,N_25433,N_27688);
xor U34081 (N_34081,N_27320,N_28734);
or U34082 (N_34082,N_26253,N_25063);
and U34083 (N_34083,N_26098,N_25285);
nor U34084 (N_34084,N_26724,N_25544);
xnor U34085 (N_34085,N_26603,N_28740);
and U34086 (N_34086,N_26487,N_26808);
and U34087 (N_34087,N_25348,N_26407);
or U34088 (N_34088,N_28407,N_29969);
or U34089 (N_34089,N_26700,N_27537);
nand U34090 (N_34090,N_25025,N_25633);
and U34091 (N_34091,N_29952,N_26118);
nand U34092 (N_34092,N_26508,N_27336);
xnor U34093 (N_34093,N_27980,N_26956);
or U34094 (N_34094,N_25720,N_28997);
nand U34095 (N_34095,N_26151,N_26808);
and U34096 (N_34096,N_28068,N_25103);
and U34097 (N_34097,N_25842,N_27013);
nand U34098 (N_34098,N_25829,N_27751);
and U34099 (N_34099,N_26212,N_26612);
nand U34100 (N_34100,N_29101,N_29703);
nor U34101 (N_34101,N_29533,N_28032);
xor U34102 (N_34102,N_28628,N_25182);
xor U34103 (N_34103,N_28357,N_29418);
nand U34104 (N_34104,N_26862,N_27554);
nor U34105 (N_34105,N_28641,N_28732);
xnor U34106 (N_34106,N_26020,N_25108);
nand U34107 (N_34107,N_29134,N_25596);
and U34108 (N_34108,N_29894,N_25884);
nand U34109 (N_34109,N_26388,N_29801);
and U34110 (N_34110,N_25725,N_28013);
nand U34111 (N_34111,N_27223,N_28950);
nand U34112 (N_34112,N_26686,N_29817);
or U34113 (N_34113,N_28451,N_27624);
and U34114 (N_34114,N_27178,N_29219);
nor U34115 (N_34115,N_29419,N_26706);
nand U34116 (N_34116,N_26955,N_29214);
nor U34117 (N_34117,N_26552,N_29886);
nand U34118 (N_34118,N_29548,N_28773);
nand U34119 (N_34119,N_27918,N_28391);
xnor U34120 (N_34120,N_25669,N_28992);
or U34121 (N_34121,N_29753,N_26480);
and U34122 (N_34122,N_25138,N_26943);
xnor U34123 (N_34123,N_27577,N_29012);
nor U34124 (N_34124,N_28226,N_29619);
and U34125 (N_34125,N_26499,N_28565);
nand U34126 (N_34126,N_26507,N_28176);
or U34127 (N_34127,N_26808,N_28490);
and U34128 (N_34128,N_28501,N_26603);
and U34129 (N_34129,N_26351,N_26156);
and U34130 (N_34130,N_26331,N_29497);
xnor U34131 (N_34131,N_29699,N_26266);
nor U34132 (N_34132,N_29482,N_29979);
xor U34133 (N_34133,N_25791,N_28086);
nand U34134 (N_34134,N_27484,N_29757);
nor U34135 (N_34135,N_25563,N_26377);
nor U34136 (N_34136,N_26846,N_28422);
xor U34137 (N_34137,N_28909,N_27780);
or U34138 (N_34138,N_28901,N_27374);
nand U34139 (N_34139,N_29783,N_28095);
xnor U34140 (N_34140,N_27035,N_29051);
nand U34141 (N_34141,N_25375,N_25297);
nand U34142 (N_34142,N_27568,N_26695);
or U34143 (N_34143,N_25665,N_26099);
xor U34144 (N_34144,N_25568,N_28288);
nand U34145 (N_34145,N_28853,N_25962);
xor U34146 (N_34146,N_29520,N_27799);
nor U34147 (N_34147,N_28136,N_26943);
and U34148 (N_34148,N_25085,N_28825);
and U34149 (N_34149,N_25546,N_27156);
or U34150 (N_34150,N_26056,N_27156);
nor U34151 (N_34151,N_27661,N_28822);
xnor U34152 (N_34152,N_29887,N_29408);
or U34153 (N_34153,N_29009,N_26696);
xnor U34154 (N_34154,N_26401,N_25731);
nor U34155 (N_34155,N_25329,N_25144);
nand U34156 (N_34156,N_29125,N_26265);
nor U34157 (N_34157,N_27002,N_29725);
and U34158 (N_34158,N_29211,N_28792);
xor U34159 (N_34159,N_28758,N_28071);
nand U34160 (N_34160,N_29658,N_25864);
nand U34161 (N_34161,N_28783,N_27554);
nand U34162 (N_34162,N_27091,N_26818);
xor U34163 (N_34163,N_25085,N_25700);
or U34164 (N_34164,N_29493,N_27601);
or U34165 (N_34165,N_29421,N_27355);
or U34166 (N_34166,N_26004,N_27357);
and U34167 (N_34167,N_27292,N_27534);
and U34168 (N_34168,N_27922,N_28635);
xnor U34169 (N_34169,N_26442,N_29764);
and U34170 (N_34170,N_26320,N_29910);
nor U34171 (N_34171,N_29610,N_28815);
or U34172 (N_34172,N_27386,N_25800);
nor U34173 (N_34173,N_29672,N_28283);
xnor U34174 (N_34174,N_25223,N_29870);
or U34175 (N_34175,N_26062,N_25083);
and U34176 (N_34176,N_28999,N_28683);
or U34177 (N_34177,N_28647,N_25288);
nor U34178 (N_34178,N_25625,N_27582);
or U34179 (N_34179,N_26596,N_27418);
xnor U34180 (N_34180,N_28407,N_25749);
nor U34181 (N_34181,N_25048,N_28297);
or U34182 (N_34182,N_29294,N_25162);
nand U34183 (N_34183,N_27103,N_26946);
xnor U34184 (N_34184,N_26883,N_29485);
xor U34185 (N_34185,N_28522,N_27795);
and U34186 (N_34186,N_29370,N_28129);
xnor U34187 (N_34187,N_25647,N_28178);
and U34188 (N_34188,N_25210,N_28082);
nand U34189 (N_34189,N_29698,N_29837);
nand U34190 (N_34190,N_29650,N_26477);
and U34191 (N_34191,N_28611,N_29982);
nand U34192 (N_34192,N_28444,N_26054);
nand U34193 (N_34193,N_26582,N_29445);
or U34194 (N_34194,N_27819,N_29029);
nand U34195 (N_34195,N_29417,N_29654);
xor U34196 (N_34196,N_28879,N_29607);
nor U34197 (N_34197,N_26683,N_29055);
and U34198 (N_34198,N_26037,N_27685);
and U34199 (N_34199,N_26105,N_28586);
and U34200 (N_34200,N_28329,N_27856);
nand U34201 (N_34201,N_29510,N_25292);
or U34202 (N_34202,N_25155,N_29061);
and U34203 (N_34203,N_28242,N_25974);
nor U34204 (N_34204,N_28372,N_25320);
nand U34205 (N_34205,N_28470,N_27347);
nor U34206 (N_34206,N_25067,N_29394);
xnor U34207 (N_34207,N_26965,N_25585);
or U34208 (N_34208,N_29450,N_29097);
and U34209 (N_34209,N_25865,N_28348);
xor U34210 (N_34210,N_28935,N_25459);
xor U34211 (N_34211,N_28876,N_25571);
or U34212 (N_34212,N_25425,N_28613);
or U34213 (N_34213,N_28864,N_26572);
nand U34214 (N_34214,N_29767,N_25703);
and U34215 (N_34215,N_27878,N_28725);
nor U34216 (N_34216,N_26028,N_25895);
nor U34217 (N_34217,N_25540,N_25765);
nor U34218 (N_34218,N_28880,N_29669);
nor U34219 (N_34219,N_26133,N_26563);
xnor U34220 (N_34220,N_27578,N_29482);
nand U34221 (N_34221,N_25082,N_29274);
xor U34222 (N_34222,N_25641,N_26514);
and U34223 (N_34223,N_28609,N_29271);
xnor U34224 (N_34224,N_28309,N_25180);
nor U34225 (N_34225,N_27381,N_27036);
and U34226 (N_34226,N_29061,N_25930);
nor U34227 (N_34227,N_29138,N_28327);
and U34228 (N_34228,N_28370,N_25372);
xor U34229 (N_34229,N_26928,N_25114);
nand U34230 (N_34230,N_27094,N_26713);
nor U34231 (N_34231,N_29275,N_27015);
xnor U34232 (N_34232,N_28302,N_27002);
nor U34233 (N_34233,N_26500,N_25991);
and U34234 (N_34234,N_25064,N_28103);
xor U34235 (N_34235,N_25491,N_29523);
or U34236 (N_34236,N_29344,N_28985);
nor U34237 (N_34237,N_25134,N_28304);
xor U34238 (N_34238,N_26391,N_25216);
nand U34239 (N_34239,N_27029,N_28377);
or U34240 (N_34240,N_27536,N_26243);
and U34241 (N_34241,N_26837,N_26883);
nand U34242 (N_34242,N_26421,N_27443);
or U34243 (N_34243,N_27936,N_28550);
or U34244 (N_34244,N_26001,N_29278);
nand U34245 (N_34245,N_27239,N_28125);
nand U34246 (N_34246,N_29527,N_25622);
and U34247 (N_34247,N_27777,N_29890);
nor U34248 (N_34248,N_25710,N_29770);
nand U34249 (N_34249,N_29095,N_25326);
or U34250 (N_34250,N_28910,N_29543);
or U34251 (N_34251,N_26181,N_29229);
nand U34252 (N_34252,N_29908,N_26564);
or U34253 (N_34253,N_29194,N_27949);
nor U34254 (N_34254,N_26383,N_29720);
nand U34255 (N_34255,N_28422,N_29062);
nor U34256 (N_34256,N_29181,N_28032);
nand U34257 (N_34257,N_26645,N_25608);
and U34258 (N_34258,N_28945,N_27237);
nor U34259 (N_34259,N_25808,N_29909);
nand U34260 (N_34260,N_26096,N_26011);
nand U34261 (N_34261,N_27163,N_26846);
and U34262 (N_34262,N_29671,N_25353);
nor U34263 (N_34263,N_27488,N_27084);
nand U34264 (N_34264,N_27117,N_25051);
nor U34265 (N_34265,N_28903,N_28679);
nor U34266 (N_34266,N_27533,N_25089);
and U34267 (N_34267,N_28047,N_29418);
xor U34268 (N_34268,N_27644,N_25531);
or U34269 (N_34269,N_25116,N_29038);
nand U34270 (N_34270,N_26576,N_28779);
or U34271 (N_34271,N_26538,N_26724);
and U34272 (N_34272,N_25592,N_28247);
xor U34273 (N_34273,N_26834,N_28248);
and U34274 (N_34274,N_26213,N_25612);
xnor U34275 (N_34275,N_25723,N_27601);
xor U34276 (N_34276,N_27715,N_26495);
and U34277 (N_34277,N_25227,N_29368);
or U34278 (N_34278,N_29504,N_29437);
nor U34279 (N_34279,N_25047,N_25050);
and U34280 (N_34280,N_26640,N_29937);
or U34281 (N_34281,N_28776,N_29438);
or U34282 (N_34282,N_25719,N_28462);
nor U34283 (N_34283,N_27077,N_28696);
xnor U34284 (N_34284,N_28547,N_28114);
or U34285 (N_34285,N_27538,N_27507);
xor U34286 (N_34286,N_27740,N_28120);
nor U34287 (N_34287,N_28605,N_29743);
or U34288 (N_34288,N_28611,N_29962);
nand U34289 (N_34289,N_27027,N_27216);
xnor U34290 (N_34290,N_26113,N_25947);
nand U34291 (N_34291,N_27591,N_25217);
xor U34292 (N_34292,N_29258,N_26798);
nand U34293 (N_34293,N_26722,N_26684);
nand U34294 (N_34294,N_27786,N_29473);
xnor U34295 (N_34295,N_25935,N_28041);
or U34296 (N_34296,N_29815,N_29013);
nand U34297 (N_34297,N_27510,N_27245);
nand U34298 (N_34298,N_27593,N_27094);
xnor U34299 (N_34299,N_28411,N_28052);
nand U34300 (N_34300,N_25942,N_29008);
xor U34301 (N_34301,N_26708,N_25840);
and U34302 (N_34302,N_29363,N_27792);
nand U34303 (N_34303,N_27036,N_28604);
nand U34304 (N_34304,N_27215,N_29166);
nor U34305 (N_34305,N_26382,N_29144);
and U34306 (N_34306,N_28795,N_26656);
and U34307 (N_34307,N_29181,N_29763);
or U34308 (N_34308,N_25601,N_29217);
xnor U34309 (N_34309,N_29223,N_29193);
nor U34310 (N_34310,N_26312,N_29887);
and U34311 (N_34311,N_25007,N_26976);
or U34312 (N_34312,N_25046,N_28233);
or U34313 (N_34313,N_29831,N_25186);
nor U34314 (N_34314,N_29658,N_28951);
and U34315 (N_34315,N_27978,N_29172);
or U34316 (N_34316,N_25123,N_28105);
and U34317 (N_34317,N_27699,N_27550);
or U34318 (N_34318,N_26150,N_28617);
and U34319 (N_34319,N_26804,N_27196);
nand U34320 (N_34320,N_29420,N_25951);
or U34321 (N_34321,N_28055,N_27550);
nor U34322 (N_34322,N_29589,N_26301);
or U34323 (N_34323,N_27196,N_28148);
nand U34324 (N_34324,N_27060,N_28959);
nand U34325 (N_34325,N_25260,N_28687);
or U34326 (N_34326,N_25423,N_29100);
and U34327 (N_34327,N_29304,N_25244);
xnor U34328 (N_34328,N_28010,N_26953);
xor U34329 (N_34329,N_25688,N_25611);
and U34330 (N_34330,N_28447,N_28601);
xor U34331 (N_34331,N_26801,N_26837);
nand U34332 (N_34332,N_26196,N_28039);
or U34333 (N_34333,N_27781,N_28981);
nand U34334 (N_34334,N_28662,N_28783);
xor U34335 (N_34335,N_25952,N_26658);
nor U34336 (N_34336,N_28413,N_27254);
nand U34337 (N_34337,N_29836,N_28421);
or U34338 (N_34338,N_25841,N_28868);
nor U34339 (N_34339,N_25914,N_27613);
xnor U34340 (N_34340,N_26889,N_26425);
xnor U34341 (N_34341,N_27606,N_27020);
or U34342 (N_34342,N_26237,N_28462);
or U34343 (N_34343,N_27951,N_28018);
nand U34344 (N_34344,N_29319,N_29340);
nor U34345 (N_34345,N_26152,N_29019);
xnor U34346 (N_34346,N_25916,N_26803);
and U34347 (N_34347,N_25799,N_27130);
nor U34348 (N_34348,N_29263,N_27566);
or U34349 (N_34349,N_26128,N_28923);
nor U34350 (N_34350,N_28640,N_29685);
and U34351 (N_34351,N_26436,N_25817);
nor U34352 (N_34352,N_29036,N_27619);
xnor U34353 (N_34353,N_25484,N_29166);
nand U34354 (N_34354,N_25770,N_29258);
nor U34355 (N_34355,N_27356,N_26014);
and U34356 (N_34356,N_29214,N_29948);
nor U34357 (N_34357,N_27299,N_26523);
nand U34358 (N_34358,N_26807,N_26501);
xor U34359 (N_34359,N_27077,N_25208);
xor U34360 (N_34360,N_25553,N_29091);
and U34361 (N_34361,N_28313,N_27455);
nand U34362 (N_34362,N_27065,N_26316);
nor U34363 (N_34363,N_26045,N_27889);
nor U34364 (N_34364,N_25847,N_28304);
and U34365 (N_34365,N_29681,N_25081);
or U34366 (N_34366,N_27820,N_25202);
or U34367 (N_34367,N_26394,N_26902);
and U34368 (N_34368,N_25968,N_29481);
xor U34369 (N_34369,N_26896,N_29756);
nor U34370 (N_34370,N_27897,N_26845);
nand U34371 (N_34371,N_29329,N_28095);
or U34372 (N_34372,N_27652,N_27632);
xnor U34373 (N_34373,N_28505,N_26422);
and U34374 (N_34374,N_28658,N_28064);
or U34375 (N_34375,N_26415,N_25195);
and U34376 (N_34376,N_29147,N_28307);
xnor U34377 (N_34377,N_25529,N_27043);
nand U34378 (N_34378,N_25688,N_28031);
and U34379 (N_34379,N_25250,N_28233);
nand U34380 (N_34380,N_26392,N_25801);
nand U34381 (N_34381,N_25588,N_25880);
or U34382 (N_34382,N_27277,N_28644);
and U34383 (N_34383,N_26724,N_27953);
or U34384 (N_34384,N_26067,N_26303);
or U34385 (N_34385,N_25497,N_27991);
nor U34386 (N_34386,N_29590,N_25365);
nor U34387 (N_34387,N_28584,N_26196);
nor U34388 (N_34388,N_28718,N_25545);
nand U34389 (N_34389,N_27777,N_25493);
or U34390 (N_34390,N_26210,N_29169);
xnor U34391 (N_34391,N_25289,N_26486);
and U34392 (N_34392,N_26851,N_28931);
nand U34393 (N_34393,N_27091,N_28053);
nand U34394 (N_34394,N_29927,N_28494);
nand U34395 (N_34395,N_26702,N_25693);
nor U34396 (N_34396,N_27292,N_26285);
nand U34397 (N_34397,N_25800,N_28169);
or U34398 (N_34398,N_25282,N_25520);
nor U34399 (N_34399,N_26309,N_26183);
or U34400 (N_34400,N_29914,N_27787);
xor U34401 (N_34401,N_25839,N_25262);
nor U34402 (N_34402,N_28272,N_25535);
xor U34403 (N_34403,N_27760,N_28532);
nor U34404 (N_34404,N_28848,N_28904);
or U34405 (N_34405,N_28867,N_29991);
and U34406 (N_34406,N_25969,N_29534);
nor U34407 (N_34407,N_29797,N_29208);
nor U34408 (N_34408,N_25367,N_28927);
nand U34409 (N_34409,N_27548,N_28655);
xnor U34410 (N_34410,N_28435,N_25987);
and U34411 (N_34411,N_25303,N_29635);
nor U34412 (N_34412,N_28785,N_29143);
or U34413 (N_34413,N_28950,N_29812);
nor U34414 (N_34414,N_25221,N_29080);
or U34415 (N_34415,N_28848,N_26920);
or U34416 (N_34416,N_27452,N_25373);
nor U34417 (N_34417,N_29040,N_27834);
nor U34418 (N_34418,N_29064,N_27500);
nand U34419 (N_34419,N_26600,N_27684);
nor U34420 (N_34420,N_27002,N_27015);
or U34421 (N_34421,N_29612,N_29438);
xor U34422 (N_34422,N_27106,N_29607);
and U34423 (N_34423,N_27900,N_29038);
nand U34424 (N_34424,N_26763,N_26748);
or U34425 (N_34425,N_29015,N_29307);
or U34426 (N_34426,N_29674,N_26468);
xnor U34427 (N_34427,N_27903,N_28836);
and U34428 (N_34428,N_29343,N_25188);
nand U34429 (N_34429,N_28101,N_25602);
nor U34430 (N_34430,N_29046,N_28230);
nor U34431 (N_34431,N_27634,N_25919);
nor U34432 (N_34432,N_25604,N_29572);
nor U34433 (N_34433,N_27043,N_26863);
nor U34434 (N_34434,N_28718,N_28247);
or U34435 (N_34435,N_29253,N_25167);
nand U34436 (N_34436,N_29937,N_25949);
nand U34437 (N_34437,N_29347,N_27178);
nor U34438 (N_34438,N_29454,N_26585);
and U34439 (N_34439,N_27184,N_25085);
or U34440 (N_34440,N_25696,N_26463);
or U34441 (N_34441,N_28465,N_29098);
nor U34442 (N_34442,N_27526,N_29133);
nand U34443 (N_34443,N_28690,N_27169);
and U34444 (N_34444,N_28256,N_28704);
nor U34445 (N_34445,N_28819,N_25692);
and U34446 (N_34446,N_26816,N_27461);
nor U34447 (N_34447,N_28483,N_27370);
nand U34448 (N_34448,N_26820,N_29598);
nand U34449 (N_34449,N_28438,N_25137);
or U34450 (N_34450,N_28655,N_26805);
nand U34451 (N_34451,N_29476,N_28439);
xnor U34452 (N_34452,N_28824,N_25434);
xnor U34453 (N_34453,N_26730,N_27277);
nand U34454 (N_34454,N_25601,N_28319);
and U34455 (N_34455,N_26556,N_28873);
xor U34456 (N_34456,N_25254,N_27900);
nor U34457 (N_34457,N_25983,N_27177);
nor U34458 (N_34458,N_28351,N_25185);
and U34459 (N_34459,N_27520,N_27408);
xor U34460 (N_34460,N_28584,N_29598);
nor U34461 (N_34461,N_25499,N_28840);
xnor U34462 (N_34462,N_27041,N_26017);
nor U34463 (N_34463,N_26175,N_25585);
and U34464 (N_34464,N_29377,N_26495);
xnor U34465 (N_34465,N_27806,N_29718);
nand U34466 (N_34466,N_29658,N_25195);
and U34467 (N_34467,N_25333,N_26914);
xnor U34468 (N_34468,N_28406,N_25112);
nor U34469 (N_34469,N_28895,N_26602);
nor U34470 (N_34470,N_26779,N_26541);
xnor U34471 (N_34471,N_25438,N_26330);
nand U34472 (N_34472,N_25108,N_29303);
xnor U34473 (N_34473,N_27464,N_26441);
nand U34474 (N_34474,N_28769,N_27744);
nor U34475 (N_34475,N_25257,N_26653);
and U34476 (N_34476,N_29835,N_26339);
or U34477 (N_34477,N_26420,N_29987);
nor U34478 (N_34478,N_29899,N_28173);
or U34479 (N_34479,N_25660,N_26638);
or U34480 (N_34480,N_26755,N_26651);
xnor U34481 (N_34481,N_25731,N_29151);
xnor U34482 (N_34482,N_25671,N_26311);
and U34483 (N_34483,N_27433,N_27637);
and U34484 (N_34484,N_28069,N_29436);
and U34485 (N_34485,N_27754,N_29324);
or U34486 (N_34486,N_27481,N_26567);
nand U34487 (N_34487,N_25012,N_27664);
xor U34488 (N_34488,N_25782,N_28761);
or U34489 (N_34489,N_28749,N_25587);
nor U34490 (N_34490,N_26003,N_26084);
nand U34491 (N_34491,N_29660,N_28461);
nand U34492 (N_34492,N_25009,N_26065);
or U34493 (N_34493,N_26728,N_25473);
or U34494 (N_34494,N_27412,N_27847);
nor U34495 (N_34495,N_26233,N_25185);
xor U34496 (N_34496,N_25184,N_26345);
and U34497 (N_34497,N_27555,N_29252);
or U34498 (N_34498,N_27391,N_25373);
and U34499 (N_34499,N_26648,N_25746);
xnor U34500 (N_34500,N_29844,N_29349);
nand U34501 (N_34501,N_25074,N_28924);
nor U34502 (N_34502,N_27022,N_29028);
or U34503 (N_34503,N_26790,N_26873);
nand U34504 (N_34504,N_29158,N_28117);
and U34505 (N_34505,N_29397,N_27516);
and U34506 (N_34506,N_25186,N_25991);
nor U34507 (N_34507,N_27305,N_27441);
and U34508 (N_34508,N_25268,N_29109);
xor U34509 (N_34509,N_28672,N_26182);
nand U34510 (N_34510,N_25654,N_25695);
or U34511 (N_34511,N_27619,N_25215);
or U34512 (N_34512,N_25661,N_27238);
nand U34513 (N_34513,N_27000,N_27404);
nand U34514 (N_34514,N_27321,N_25511);
or U34515 (N_34515,N_27165,N_29800);
nor U34516 (N_34516,N_28275,N_25639);
nor U34517 (N_34517,N_25921,N_29323);
or U34518 (N_34518,N_25748,N_29570);
or U34519 (N_34519,N_25177,N_27148);
nand U34520 (N_34520,N_27311,N_29287);
xor U34521 (N_34521,N_27947,N_27498);
or U34522 (N_34522,N_27319,N_29117);
nor U34523 (N_34523,N_29403,N_29599);
xnor U34524 (N_34524,N_25871,N_27112);
and U34525 (N_34525,N_29852,N_28431);
or U34526 (N_34526,N_26654,N_26093);
and U34527 (N_34527,N_28884,N_27635);
nand U34528 (N_34528,N_26755,N_29987);
and U34529 (N_34529,N_27982,N_25295);
nand U34530 (N_34530,N_29898,N_28131);
nand U34531 (N_34531,N_29110,N_26551);
xnor U34532 (N_34532,N_25818,N_28711);
and U34533 (N_34533,N_26907,N_29913);
nor U34534 (N_34534,N_27570,N_25845);
nand U34535 (N_34535,N_29399,N_29464);
xor U34536 (N_34536,N_26190,N_28572);
nand U34537 (N_34537,N_29092,N_27971);
or U34538 (N_34538,N_27930,N_27385);
nand U34539 (N_34539,N_27421,N_29995);
nor U34540 (N_34540,N_29911,N_27951);
and U34541 (N_34541,N_29567,N_28325);
and U34542 (N_34542,N_29947,N_27836);
nand U34543 (N_34543,N_27824,N_28503);
nand U34544 (N_34544,N_28795,N_29826);
and U34545 (N_34545,N_26972,N_25008);
xnor U34546 (N_34546,N_26510,N_29171);
xor U34547 (N_34547,N_25720,N_28632);
xor U34548 (N_34548,N_29419,N_29715);
or U34549 (N_34549,N_25572,N_27666);
and U34550 (N_34550,N_26851,N_27916);
and U34551 (N_34551,N_27970,N_26126);
and U34552 (N_34552,N_28441,N_25516);
nand U34553 (N_34553,N_29786,N_27854);
and U34554 (N_34554,N_29484,N_29925);
or U34555 (N_34555,N_28038,N_25027);
and U34556 (N_34556,N_27328,N_27197);
nor U34557 (N_34557,N_27692,N_26608);
nor U34558 (N_34558,N_25094,N_25495);
and U34559 (N_34559,N_29400,N_25552);
nand U34560 (N_34560,N_27355,N_25637);
nor U34561 (N_34561,N_29998,N_25100);
and U34562 (N_34562,N_29066,N_29654);
and U34563 (N_34563,N_28557,N_25001);
nor U34564 (N_34564,N_29926,N_29073);
nand U34565 (N_34565,N_28866,N_28431);
nand U34566 (N_34566,N_29572,N_28241);
xor U34567 (N_34567,N_26666,N_27510);
nor U34568 (N_34568,N_27530,N_27759);
nand U34569 (N_34569,N_26374,N_27531);
nor U34570 (N_34570,N_29799,N_25881);
or U34571 (N_34571,N_29786,N_25234);
and U34572 (N_34572,N_29208,N_27343);
or U34573 (N_34573,N_28591,N_27802);
and U34574 (N_34574,N_25259,N_25476);
nor U34575 (N_34575,N_28025,N_27057);
xnor U34576 (N_34576,N_27752,N_27112);
or U34577 (N_34577,N_26504,N_27282);
or U34578 (N_34578,N_26157,N_26780);
or U34579 (N_34579,N_27372,N_25400);
xor U34580 (N_34580,N_29056,N_28133);
and U34581 (N_34581,N_26927,N_28475);
nand U34582 (N_34582,N_27334,N_25212);
and U34583 (N_34583,N_27155,N_29876);
xor U34584 (N_34584,N_27605,N_27039);
xnor U34585 (N_34585,N_29973,N_29983);
nor U34586 (N_34586,N_29478,N_28993);
nor U34587 (N_34587,N_25211,N_29282);
nor U34588 (N_34588,N_29561,N_26070);
and U34589 (N_34589,N_29654,N_25286);
and U34590 (N_34590,N_26454,N_26624);
nand U34591 (N_34591,N_26014,N_25522);
nand U34592 (N_34592,N_26430,N_28063);
nor U34593 (N_34593,N_29735,N_28587);
or U34594 (N_34594,N_27755,N_29887);
nand U34595 (N_34595,N_26869,N_25488);
nand U34596 (N_34596,N_27811,N_29102);
nand U34597 (N_34597,N_27663,N_26485);
xnor U34598 (N_34598,N_25362,N_25868);
nand U34599 (N_34599,N_29068,N_29434);
or U34600 (N_34600,N_26827,N_29696);
nor U34601 (N_34601,N_29557,N_29386);
xnor U34602 (N_34602,N_25251,N_29862);
nand U34603 (N_34603,N_27462,N_27682);
nand U34604 (N_34604,N_28746,N_27004);
xnor U34605 (N_34605,N_29927,N_25714);
and U34606 (N_34606,N_27641,N_25766);
or U34607 (N_34607,N_26745,N_25053);
xor U34608 (N_34608,N_26631,N_25239);
nand U34609 (N_34609,N_25726,N_25973);
and U34610 (N_34610,N_29958,N_25401);
xnor U34611 (N_34611,N_29822,N_26652);
or U34612 (N_34612,N_29304,N_29793);
or U34613 (N_34613,N_27738,N_27361);
and U34614 (N_34614,N_28248,N_26373);
nor U34615 (N_34615,N_28497,N_25996);
or U34616 (N_34616,N_26361,N_27123);
and U34617 (N_34617,N_25247,N_27077);
and U34618 (N_34618,N_28130,N_27072);
xnor U34619 (N_34619,N_29688,N_29986);
or U34620 (N_34620,N_27555,N_26357);
nor U34621 (N_34621,N_27245,N_29544);
nand U34622 (N_34622,N_25616,N_26633);
nand U34623 (N_34623,N_26717,N_28596);
or U34624 (N_34624,N_27615,N_28112);
or U34625 (N_34625,N_28815,N_25890);
nor U34626 (N_34626,N_29151,N_25391);
or U34627 (N_34627,N_25669,N_28626);
and U34628 (N_34628,N_29438,N_28833);
nand U34629 (N_34629,N_27066,N_26648);
xor U34630 (N_34630,N_26725,N_29184);
nand U34631 (N_34631,N_25545,N_28331);
or U34632 (N_34632,N_26237,N_28455);
and U34633 (N_34633,N_28561,N_29124);
xnor U34634 (N_34634,N_25530,N_25498);
xor U34635 (N_34635,N_28806,N_29024);
or U34636 (N_34636,N_27754,N_28918);
xnor U34637 (N_34637,N_25050,N_28560);
xor U34638 (N_34638,N_29806,N_27023);
and U34639 (N_34639,N_26468,N_27160);
or U34640 (N_34640,N_27714,N_26019);
and U34641 (N_34641,N_26715,N_29848);
nand U34642 (N_34642,N_25981,N_25666);
xor U34643 (N_34643,N_29567,N_28378);
xnor U34644 (N_34644,N_28741,N_28129);
xnor U34645 (N_34645,N_29452,N_25866);
nor U34646 (N_34646,N_29166,N_25300);
or U34647 (N_34647,N_27046,N_28260);
nand U34648 (N_34648,N_28278,N_29005);
and U34649 (N_34649,N_29599,N_28225);
nor U34650 (N_34650,N_26951,N_27178);
nor U34651 (N_34651,N_25910,N_29251);
nor U34652 (N_34652,N_28272,N_29560);
nor U34653 (N_34653,N_26205,N_29833);
xnor U34654 (N_34654,N_25007,N_25168);
or U34655 (N_34655,N_27158,N_26789);
xor U34656 (N_34656,N_26226,N_26662);
nand U34657 (N_34657,N_29710,N_25367);
nand U34658 (N_34658,N_25607,N_28850);
or U34659 (N_34659,N_25628,N_25107);
nand U34660 (N_34660,N_27662,N_29973);
and U34661 (N_34661,N_25723,N_27700);
and U34662 (N_34662,N_25125,N_29999);
xor U34663 (N_34663,N_26043,N_28846);
or U34664 (N_34664,N_28260,N_25401);
or U34665 (N_34665,N_27299,N_26100);
or U34666 (N_34666,N_29972,N_29578);
xor U34667 (N_34667,N_27766,N_25046);
nand U34668 (N_34668,N_26296,N_25944);
and U34669 (N_34669,N_27399,N_29137);
or U34670 (N_34670,N_26340,N_27371);
nand U34671 (N_34671,N_27662,N_25135);
nand U34672 (N_34672,N_29283,N_26716);
xor U34673 (N_34673,N_28440,N_25138);
xor U34674 (N_34674,N_25462,N_27662);
nor U34675 (N_34675,N_27229,N_25238);
xnor U34676 (N_34676,N_29916,N_28994);
and U34677 (N_34677,N_29355,N_29761);
and U34678 (N_34678,N_26337,N_29191);
or U34679 (N_34679,N_27738,N_25421);
xnor U34680 (N_34680,N_29364,N_28398);
and U34681 (N_34681,N_26504,N_26486);
or U34682 (N_34682,N_25225,N_26179);
and U34683 (N_34683,N_29590,N_26743);
nor U34684 (N_34684,N_25191,N_26132);
nand U34685 (N_34685,N_25047,N_26565);
nand U34686 (N_34686,N_26608,N_28323);
or U34687 (N_34687,N_25908,N_28876);
xor U34688 (N_34688,N_28930,N_26608);
nor U34689 (N_34689,N_29452,N_25282);
nand U34690 (N_34690,N_28453,N_28817);
or U34691 (N_34691,N_28129,N_29209);
or U34692 (N_34692,N_27145,N_29301);
or U34693 (N_34693,N_29727,N_29261);
nor U34694 (N_34694,N_25425,N_29690);
xor U34695 (N_34695,N_28273,N_25350);
xnor U34696 (N_34696,N_28004,N_28457);
nor U34697 (N_34697,N_29809,N_29900);
nor U34698 (N_34698,N_27000,N_27835);
nor U34699 (N_34699,N_27702,N_27347);
nand U34700 (N_34700,N_25957,N_26245);
and U34701 (N_34701,N_25251,N_28666);
or U34702 (N_34702,N_29653,N_26511);
nand U34703 (N_34703,N_26767,N_26580);
and U34704 (N_34704,N_28899,N_27479);
or U34705 (N_34705,N_29776,N_29493);
and U34706 (N_34706,N_28745,N_27161);
or U34707 (N_34707,N_25378,N_27265);
nor U34708 (N_34708,N_28119,N_29851);
and U34709 (N_34709,N_26569,N_26838);
nor U34710 (N_34710,N_25280,N_29463);
or U34711 (N_34711,N_27573,N_28740);
and U34712 (N_34712,N_28521,N_26323);
xnor U34713 (N_34713,N_26580,N_26147);
or U34714 (N_34714,N_29041,N_27946);
and U34715 (N_34715,N_25853,N_25357);
xor U34716 (N_34716,N_27775,N_26122);
xor U34717 (N_34717,N_25508,N_28909);
nand U34718 (N_34718,N_28696,N_27600);
nand U34719 (N_34719,N_28924,N_29536);
nor U34720 (N_34720,N_28173,N_26410);
xor U34721 (N_34721,N_25539,N_25345);
nor U34722 (N_34722,N_25253,N_28226);
nand U34723 (N_34723,N_27035,N_26463);
and U34724 (N_34724,N_26878,N_25755);
or U34725 (N_34725,N_25640,N_25143);
nand U34726 (N_34726,N_28191,N_26587);
nand U34727 (N_34727,N_26331,N_29245);
xnor U34728 (N_34728,N_29343,N_27465);
xor U34729 (N_34729,N_27487,N_25906);
nor U34730 (N_34730,N_28262,N_25156);
nand U34731 (N_34731,N_26554,N_25784);
nor U34732 (N_34732,N_25667,N_28836);
or U34733 (N_34733,N_29384,N_25604);
xor U34734 (N_34734,N_27828,N_26303);
nand U34735 (N_34735,N_28396,N_28561);
xnor U34736 (N_34736,N_29476,N_29078);
and U34737 (N_34737,N_29061,N_25948);
or U34738 (N_34738,N_26604,N_27039);
nor U34739 (N_34739,N_27404,N_28231);
and U34740 (N_34740,N_26309,N_27812);
or U34741 (N_34741,N_28487,N_26692);
nor U34742 (N_34742,N_28593,N_26234);
or U34743 (N_34743,N_28354,N_27871);
or U34744 (N_34744,N_26647,N_29660);
and U34745 (N_34745,N_26565,N_29658);
or U34746 (N_34746,N_25033,N_26043);
and U34747 (N_34747,N_29935,N_29352);
nor U34748 (N_34748,N_25299,N_25767);
xor U34749 (N_34749,N_27731,N_28995);
nor U34750 (N_34750,N_27680,N_28704);
xnor U34751 (N_34751,N_26585,N_26035);
nand U34752 (N_34752,N_25671,N_26797);
xnor U34753 (N_34753,N_27872,N_29473);
xor U34754 (N_34754,N_29654,N_29305);
xor U34755 (N_34755,N_27917,N_26474);
nor U34756 (N_34756,N_29406,N_27927);
nor U34757 (N_34757,N_27504,N_25768);
nand U34758 (N_34758,N_26316,N_26311);
and U34759 (N_34759,N_26591,N_28357);
nor U34760 (N_34760,N_27065,N_29543);
or U34761 (N_34761,N_26834,N_25511);
and U34762 (N_34762,N_25443,N_27279);
xor U34763 (N_34763,N_27961,N_26909);
and U34764 (N_34764,N_27110,N_26075);
nand U34765 (N_34765,N_29616,N_26490);
nand U34766 (N_34766,N_26954,N_25323);
and U34767 (N_34767,N_27506,N_26328);
or U34768 (N_34768,N_29088,N_29390);
xnor U34769 (N_34769,N_29848,N_26561);
or U34770 (N_34770,N_27501,N_29860);
and U34771 (N_34771,N_25031,N_26564);
and U34772 (N_34772,N_25658,N_29297);
nand U34773 (N_34773,N_27110,N_26592);
nand U34774 (N_34774,N_27723,N_26223);
or U34775 (N_34775,N_29890,N_26088);
and U34776 (N_34776,N_27320,N_28124);
and U34777 (N_34777,N_27342,N_28196);
nand U34778 (N_34778,N_26575,N_29494);
xor U34779 (N_34779,N_27070,N_25412);
and U34780 (N_34780,N_25786,N_25877);
nor U34781 (N_34781,N_25368,N_28640);
or U34782 (N_34782,N_26655,N_29054);
and U34783 (N_34783,N_29678,N_27689);
xnor U34784 (N_34784,N_25271,N_29804);
or U34785 (N_34785,N_25329,N_26212);
or U34786 (N_34786,N_29201,N_25017);
nand U34787 (N_34787,N_26761,N_28163);
or U34788 (N_34788,N_28446,N_29739);
and U34789 (N_34789,N_26744,N_28530);
xnor U34790 (N_34790,N_28247,N_27528);
nor U34791 (N_34791,N_28739,N_25168);
xnor U34792 (N_34792,N_27119,N_28156);
and U34793 (N_34793,N_28781,N_25087);
nand U34794 (N_34794,N_28354,N_28661);
and U34795 (N_34795,N_29485,N_28158);
and U34796 (N_34796,N_25886,N_26005);
xnor U34797 (N_34797,N_29607,N_26301);
nor U34798 (N_34798,N_26023,N_27609);
nand U34799 (N_34799,N_26387,N_27246);
xnor U34800 (N_34800,N_25303,N_29540);
xnor U34801 (N_34801,N_25854,N_27645);
nor U34802 (N_34802,N_27093,N_28513);
and U34803 (N_34803,N_29421,N_27026);
nor U34804 (N_34804,N_29695,N_27376);
nand U34805 (N_34805,N_26567,N_29228);
nand U34806 (N_34806,N_25504,N_26696);
or U34807 (N_34807,N_27197,N_28892);
and U34808 (N_34808,N_25971,N_25638);
xor U34809 (N_34809,N_28151,N_25161);
or U34810 (N_34810,N_27649,N_26207);
nand U34811 (N_34811,N_25644,N_27310);
nor U34812 (N_34812,N_29514,N_28757);
or U34813 (N_34813,N_25899,N_27976);
or U34814 (N_34814,N_26550,N_27080);
and U34815 (N_34815,N_25154,N_26768);
xnor U34816 (N_34816,N_26158,N_25814);
and U34817 (N_34817,N_25442,N_29906);
and U34818 (N_34818,N_28949,N_27016);
nor U34819 (N_34819,N_27030,N_27735);
nand U34820 (N_34820,N_27102,N_25725);
or U34821 (N_34821,N_26070,N_29417);
and U34822 (N_34822,N_25657,N_27331);
nand U34823 (N_34823,N_25485,N_25537);
and U34824 (N_34824,N_27219,N_28177);
or U34825 (N_34825,N_25782,N_26484);
nand U34826 (N_34826,N_25451,N_26988);
or U34827 (N_34827,N_29644,N_29304);
nand U34828 (N_34828,N_26908,N_25891);
nor U34829 (N_34829,N_27487,N_26940);
nand U34830 (N_34830,N_29234,N_25939);
or U34831 (N_34831,N_25822,N_25252);
nor U34832 (N_34832,N_25519,N_27271);
nand U34833 (N_34833,N_25774,N_29420);
or U34834 (N_34834,N_26890,N_29433);
or U34835 (N_34835,N_26682,N_28938);
nand U34836 (N_34836,N_25721,N_28006);
and U34837 (N_34837,N_28363,N_29509);
nand U34838 (N_34838,N_26684,N_29090);
nor U34839 (N_34839,N_25026,N_27025);
xnor U34840 (N_34840,N_25077,N_26844);
or U34841 (N_34841,N_27982,N_25729);
nor U34842 (N_34842,N_25751,N_25219);
nor U34843 (N_34843,N_28931,N_28050);
and U34844 (N_34844,N_25934,N_27543);
xor U34845 (N_34845,N_25807,N_26617);
or U34846 (N_34846,N_27377,N_28554);
nor U34847 (N_34847,N_26819,N_29576);
or U34848 (N_34848,N_25334,N_29421);
nand U34849 (N_34849,N_28449,N_25604);
and U34850 (N_34850,N_26553,N_28708);
or U34851 (N_34851,N_28196,N_26159);
nand U34852 (N_34852,N_26524,N_25486);
nor U34853 (N_34853,N_26115,N_29735);
xor U34854 (N_34854,N_29320,N_29664);
or U34855 (N_34855,N_25906,N_26298);
nor U34856 (N_34856,N_26106,N_25502);
or U34857 (N_34857,N_25373,N_27797);
xnor U34858 (N_34858,N_25883,N_29997);
or U34859 (N_34859,N_27172,N_26158);
and U34860 (N_34860,N_25563,N_26798);
xor U34861 (N_34861,N_28894,N_29952);
nand U34862 (N_34862,N_26638,N_26751);
xor U34863 (N_34863,N_28399,N_25637);
or U34864 (N_34864,N_25061,N_27618);
nor U34865 (N_34865,N_25619,N_27335);
nor U34866 (N_34866,N_29070,N_25605);
and U34867 (N_34867,N_28309,N_27616);
nor U34868 (N_34868,N_29699,N_29063);
nand U34869 (N_34869,N_25206,N_26152);
and U34870 (N_34870,N_28457,N_25604);
and U34871 (N_34871,N_29954,N_29277);
xor U34872 (N_34872,N_28195,N_29593);
xnor U34873 (N_34873,N_26138,N_26449);
or U34874 (N_34874,N_28033,N_26954);
nor U34875 (N_34875,N_29503,N_25529);
nor U34876 (N_34876,N_28957,N_27075);
xor U34877 (N_34877,N_26017,N_28056);
and U34878 (N_34878,N_28014,N_27935);
nand U34879 (N_34879,N_29968,N_28278);
or U34880 (N_34880,N_27711,N_26445);
nor U34881 (N_34881,N_28402,N_27395);
and U34882 (N_34882,N_28062,N_28714);
or U34883 (N_34883,N_28838,N_29776);
or U34884 (N_34884,N_28590,N_26648);
or U34885 (N_34885,N_26884,N_26167);
or U34886 (N_34886,N_27228,N_25605);
or U34887 (N_34887,N_28655,N_29376);
nand U34888 (N_34888,N_28542,N_25413);
nand U34889 (N_34889,N_27835,N_25380);
nor U34890 (N_34890,N_25672,N_26745);
nor U34891 (N_34891,N_28227,N_25925);
nand U34892 (N_34892,N_26234,N_25454);
xor U34893 (N_34893,N_26287,N_25425);
nor U34894 (N_34894,N_27429,N_27541);
xor U34895 (N_34895,N_25100,N_25901);
nand U34896 (N_34896,N_29736,N_29140);
nor U34897 (N_34897,N_29224,N_25440);
xor U34898 (N_34898,N_26551,N_26303);
or U34899 (N_34899,N_28210,N_28302);
and U34900 (N_34900,N_25734,N_25302);
nor U34901 (N_34901,N_25324,N_27094);
xor U34902 (N_34902,N_28184,N_25878);
xor U34903 (N_34903,N_28132,N_27283);
and U34904 (N_34904,N_26073,N_27331);
and U34905 (N_34905,N_28896,N_26676);
nand U34906 (N_34906,N_26412,N_26683);
and U34907 (N_34907,N_27030,N_28692);
nand U34908 (N_34908,N_26966,N_26401);
and U34909 (N_34909,N_26634,N_25205);
and U34910 (N_34910,N_28245,N_27464);
and U34911 (N_34911,N_25607,N_27908);
nand U34912 (N_34912,N_28283,N_28425);
and U34913 (N_34913,N_26226,N_26558);
nand U34914 (N_34914,N_26722,N_28452);
nor U34915 (N_34915,N_28386,N_28912);
nor U34916 (N_34916,N_29275,N_25441);
nor U34917 (N_34917,N_29999,N_29991);
nand U34918 (N_34918,N_28122,N_29841);
or U34919 (N_34919,N_25033,N_25018);
xnor U34920 (N_34920,N_25715,N_26034);
xor U34921 (N_34921,N_26710,N_27146);
nand U34922 (N_34922,N_27343,N_28848);
nand U34923 (N_34923,N_29609,N_27101);
and U34924 (N_34924,N_26191,N_29047);
or U34925 (N_34925,N_25823,N_27577);
nor U34926 (N_34926,N_29183,N_25833);
and U34927 (N_34927,N_29335,N_26701);
xnor U34928 (N_34928,N_25576,N_29063);
xnor U34929 (N_34929,N_26222,N_25431);
and U34930 (N_34930,N_25185,N_29703);
and U34931 (N_34931,N_27521,N_27983);
xnor U34932 (N_34932,N_28703,N_26020);
nand U34933 (N_34933,N_29470,N_26882);
and U34934 (N_34934,N_28591,N_25753);
nand U34935 (N_34935,N_27286,N_29533);
xnor U34936 (N_34936,N_25667,N_25777);
or U34937 (N_34937,N_27571,N_28817);
nand U34938 (N_34938,N_29704,N_26533);
xor U34939 (N_34939,N_26591,N_28564);
xnor U34940 (N_34940,N_29932,N_25533);
and U34941 (N_34941,N_26677,N_27400);
xor U34942 (N_34942,N_29659,N_29255);
xor U34943 (N_34943,N_26469,N_25718);
nor U34944 (N_34944,N_25393,N_29585);
and U34945 (N_34945,N_26138,N_25914);
nand U34946 (N_34946,N_26511,N_28041);
nand U34947 (N_34947,N_25345,N_26377);
xnor U34948 (N_34948,N_26244,N_25912);
or U34949 (N_34949,N_28717,N_25659);
xor U34950 (N_34950,N_29151,N_25235);
and U34951 (N_34951,N_28229,N_25688);
xnor U34952 (N_34952,N_28405,N_25031);
and U34953 (N_34953,N_27897,N_25442);
or U34954 (N_34954,N_26174,N_25458);
or U34955 (N_34955,N_26712,N_28979);
nand U34956 (N_34956,N_28397,N_26154);
or U34957 (N_34957,N_29481,N_28010);
and U34958 (N_34958,N_29205,N_26863);
nand U34959 (N_34959,N_27367,N_26379);
xor U34960 (N_34960,N_26069,N_27630);
or U34961 (N_34961,N_27832,N_28284);
nand U34962 (N_34962,N_25533,N_27547);
xor U34963 (N_34963,N_26817,N_28867);
or U34964 (N_34964,N_25411,N_29828);
xor U34965 (N_34965,N_27469,N_29100);
xor U34966 (N_34966,N_28326,N_27613);
nand U34967 (N_34967,N_29629,N_29844);
and U34968 (N_34968,N_29410,N_25078);
xor U34969 (N_34969,N_25148,N_27772);
or U34970 (N_34970,N_28780,N_28095);
xnor U34971 (N_34971,N_25636,N_29618);
xor U34972 (N_34972,N_26559,N_29201);
xor U34973 (N_34973,N_28966,N_26956);
nor U34974 (N_34974,N_25441,N_26701);
or U34975 (N_34975,N_26018,N_29211);
nor U34976 (N_34976,N_29495,N_25996);
xor U34977 (N_34977,N_28111,N_26395);
or U34978 (N_34978,N_26616,N_25332);
xor U34979 (N_34979,N_28139,N_26690);
or U34980 (N_34980,N_25866,N_27241);
and U34981 (N_34981,N_26930,N_27628);
nand U34982 (N_34982,N_27074,N_26014);
nor U34983 (N_34983,N_25681,N_29472);
nand U34984 (N_34984,N_26321,N_28024);
nor U34985 (N_34985,N_27267,N_29123);
xor U34986 (N_34986,N_28314,N_27899);
nand U34987 (N_34987,N_27556,N_29584);
and U34988 (N_34988,N_27142,N_28010);
xor U34989 (N_34989,N_26831,N_27736);
or U34990 (N_34990,N_25680,N_29178);
or U34991 (N_34991,N_27462,N_29527);
xor U34992 (N_34992,N_26041,N_29621);
and U34993 (N_34993,N_25427,N_25830);
nand U34994 (N_34994,N_28862,N_25302);
nor U34995 (N_34995,N_25666,N_29331);
and U34996 (N_34996,N_28292,N_27187);
or U34997 (N_34997,N_27812,N_27292);
nand U34998 (N_34998,N_25412,N_28194);
and U34999 (N_34999,N_28840,N_25458);
and U35000 (N_35000,N_31109,N_34597);
xor U35001 (N_35001,N_33163,N_34017);
and U35002 (N_35002,N_30170,N_32042);
and U35003 (N_35003,N_33250,N_32775);
and U35004 (N_35004,N_31042,N_31657);
or U35005 (N_35005,N_32223,N_31519);
or U35006 (N_35006,N_31735,N_31580);
xnor U35007 (N_35007,N_30870,N_33754);
or U35008 (N_35008,N_32591,N_34709);
nand U35009 (N_35009,N_30216,N_30364);
nor U35010 (N_35010,N_32045,N_34820);
nor U35011 (N_35011,N_34927,N_32531);
or U35012 (N_35012,N_31771,N_30142);
nor U35013 (N_35013,N_34288,N_34572);
xor U35014 (N_35014,N_33888,N_31597);
or U35015 (N_35015,N_33029,N_34278);
nor U35016 (N_35016,N_32150,N_34953);
or U35017 (N_35017,N_34656,N_32702);
nand U35018 (N_35018,N_34168,N_31670);
nand U35019 (N_35019,N_31856,N_34635);
and U35020 (N_35020,N_34480,N_33130);
nand U35021 (N_35021,N_34557,N_31116);
nor U35022 (N_35022,N_31062,N_34190);
or U35023 (N_35023,N_30827,N_33697);
and U35024 (N_35024,N_33168,N_32035);
nor U35025 (N_35025,N_31774,N_31700);
xor U35026 (N_35026,N_34984,N_32827);
and U35027 (N_35027,N_33789,N_34083);
nand U35028 (N_35028,N_30409,N_33613);
xor U35029 (N_35029,N_34834,N_33334);
nand U35030 (N_35030,N_34523,N_33696);
nor U35031 (N_35031,N_34677,N_30382);
nand U35032 (N_35032,N_31563,N_31325);
nor U35033 (N_35033,N_34718,N_30109);
and U35034 (N_35034,N_31345,N_34366);
nand U35035 (N_35035,N_31592,N_30988);
xnor U35036 (N_35036,N_32247,N_33700);
nand U35037 (N_35037,N_33680,N_33237);
nor U35038 (N_35038,N_31051,N_31830);
nand U35039 (N_35039,N_32790,N_30854);
nand U35040 (N_35040,N_32294,N_30708);
nor U35041 (N_35041,N_34397,N_31476);
and U35042 (N_35042,N_33928,N_33894);
nor U35043 (N_35043,N_31643,N_30631);
or U35044 (N_35044,N_34121,N_30043);
and U35045 (N_35045,N_32895,N_31527);
or U35046 (N_35046,N_31413,N_34883);
nand U35047 (N_35047,N_33953,N_31259);
and U35048 (N_35048,N_32388,N_31258);
xnor U35049 (N_35049,N_33002,N_32421);
nor U35050 (N_35050,N_33837,N_34080);
or U35051 (N_35051,N_31512,N_32009);
or U35052 (N_35052,N_34568,N_31965);
or U35053 (N_35053,N_30837,N_32707);
nor U35054 (N_35054,N_33982,N_33795);
xor U35055 (N_35055,N_30363,N_34165);
or U35056 (N_35056,N_34056,N_32161);
nand U35057 (N_35057,N_33213,N_34669);
or U35058 (N_35058,N_34072,N_32744);
xor U35059 (N_35059,N_31434,N_32530);
xnor U35060 (N_35060,N_33351,N_30129);
nor U35061 (N_35061,N_33620,N_31860);
nand U35062 (N_35062,N_32348,N_33821);
and U35063 (N_35063,N_32039,N_34211);
or U35064 (N_35064,N_30789,N_32711);
and U35065 (N_35065,N_33025,N_34286);
nor U35066 (N_35066,N_30121,N_30374);
nand U35067 (N_35067,N_34571,N_34443);
or U35068 (N_35068,N_33436,N_34719);
xnor U35069 (N_35069,N_34336,N_30327);
nor U35070 (N_35070,N_30989,N_30038);
nand U35071 (N_35071,N_33364,N_33793);
and U35072 (N_35072,N_32489,N_30978);
xnor U35073 (N_35073,N_33882,N_30405);
and U35074 (N_35074,N_34796,N_32867);
and U35075 (N_35075,N_33156,N_33994);
nor U35076 (N_35076,N_34529,N_32111);
or U35077 (N_35077,N_33373,N_32140);
and U35078 (N_35078,N_31869,N_34987);
and U35079 (N_35079,N_30065,N_31544);
and U35080 (N_35080,N_30307,N_32426);
xnor U35081 (N_35081,N_33021,N_32669);
or U35082 (N_35082,N_34029,N_34573);
nor U35083 (N_35083,N_33398,N_32667);
nand U35084 (N_35084,N_32468,N_34531);
or U35085 (N_35085,N_32355,N_32411);
nor U35086 (N_35086,N_30135,N_32728);
xnor U35087 (N_35087,N_32301,N_31163);
or U35088 (N_35088,N_30194,N_32651);
and U35089 (N_35089,N_34684,N_34031);
nand U35090 (N_35090,N_33157,N_30270);
or U35091 (N_35091,N_32948,N_34372);
or U35092 (N_35092,N_31990,N_31154);
xor U35093 (N_35093,N_31407,N_30696);
and U35094 (N_35094,N_31352,N_33312);
nand U35095 (N_35095,N_30034,N_34099);
or U35096 (N_35096,N_32491,N_31740);
nand U35097 (N_35097,N_32692,N_32668);
and U35098 (N_35098,N_30919,N_34246);
xnor U35099 (N_35099,N_31056,N_34837);
nor U35100 (N_35100,N_31862,N_30895);
and U35101 (N_35101,N_34651,N_32276);
and U35102 (N_35102,N_30261,N_33410);
or U35103 (N_35103,N_32783,N_30878);
nand U35104 (N_35104,N_31347,N_34590);
nand U35105 (N_35105,N_30259,N_33149);
xnor U35106 (N_35106,N_32072,N_32563);
and U35107 (N_35107,N_32008,N_34600);
nor U35108 (N_35108,N_33178,N_32753);
or U35109 (N_35109,N_30277,N_34346);
nand U35110 (N_35110,N_30795,N_30190);
xor U35111 (N_35111,N_34063,N_34673);
nand U35112 (N_35112,N_33191,N_30301);
or U35113 (N_35113,N_34822,N_33097);
nand U35114 (N_35114,N_31606,N_33641);
and U35115 (N_35115,N_33689,N_30380);
xor U35116 (N_35116,N_34505,N_30175);
xor U35117 (N_35117,N_32506,N_33577);
or U35118 (N_35118,N_33408,N_30045);
xnor U35119 (N_35119,N_31703,N_31080);
and U35120 (N_35120,N_31686,N_32525);
and U35121 (N_35121,N_33425,N_31736);
nand U35122 (N_35122,N_31414,N_32133);
nor U35123 (N_35123,N_32318,N_31857);
and U35124 (N_35124,N_31999,N_33561);
or U35125 (N_35125,N_31130,N_30164);
nand U35126 (N_35126,N_32834,N_31161);
nor U35127 (N_35127,N_34409,N_34995);
and U35128 (N_35128,N_34581,N_32049);
and U35129 (N_35129,N_34304,N_34858);
and U35130 (N_35130,N_33703,N_32710);
or U35131 (N_35131,N_30544,N_32110);
and U35132 (N_35132,N_31293,N_32210);
or U35133 (N_35133,N_33595,N_33659);
or U35134 (N_35134,N_31859,N_34267);
nand U35135 (N_35135,N_33397,N_30250);
nor U35136 (N_35136,N_31150,N_33511);
and U35137 (N_35137,N_34695,N_30757);
and U35138 (N_35138,N_30794,N_31764);
nor U35139 (N_35139,N_34191,N_31840);
nor U35140 (N_35140,N_31674,N_31377);
and U35141 (N_35141,N_32630,N_33433);
or U35142 (N_35142,N_32296,N_32966);
nand U35143 (N_35143,N_31212,N_31672);
and U35144 (N_35144,N_32921,N_31782);
or U35145 (N_35145,N_32311,N_32559);
or U35146 (N_35146,N_32521,N_34806);
xor U35147 (N_35147,N_32016,N_34956);
and U35148 (N_35148,N_32738,N_34892);
nor U35149 (N_35149,N_34844,N_34354);
and U35150 (N_35150,N_34838,N_34716);
or U35151 (N_35151,N_32583,N_31788);
nand U35152 (N_35152,N_33188,N_31270);
xnor U35153 (N_35153,N_32218,N_31283);
nand U35154 (N_35154,N_30566,N_31517);
nor U35155 (N_35155,N_32891,N_32507);
nor U35156 (N_35156,N_32899,N_32097);
nor U35157 (N_35157,N_32604,N_32396);
nor U35158 (N_35158,N_34789,N_32944);
nor U35159 (N_35159,N_33284,N_33485);
nor U35160 (N_35160,N_30630,N_33540);
xnor U35161 (N_35161,N_34298,N_31732);
xnor U35162 (N_35162,N_30984,N_34075);
nor U35163 (N_35163,N_30830,N_34810);
and U35164 (N_35164,N_33639,N_33495);
and U35165 (N_35165,N_30114,N_33277);
nor U35166 (N_35166,N_33767,N_31392);
or U35167 (N_35167,N_34242,N_32767);
or U35168 (N_35168,N_34608,N_32733);
or U35169 (N_35169,N_30865,N_33228);
nand U35170 (N_35170,N_30267,N_30859);
xor U35171 (N_35171,N_33083,N_31421);
or U35172 (N_35172,N_31077,N_34282);
or U35173 (N_35173,N_34853,N_33472);
nand U35174 (N_35174,N_31743,N_32758);
nor U35175 (N_35175,N_32328,N_33497);
nor U35176 (N_35176,N_32973,N_31280);
and U35177 (N_35177,N_31692,N_31813);
nand U35178 (N_35178,N_33819,N_31490);
nand U35179 (N_35179,N_30366,N_34429);
or U35180 (N_35180,N_30019,N_34813);
xnor U35181 (N_35181,N_31004,N_34802);
xnor U35182 (N_35182,N_34711,N_34322);
nand U35183 (N_35183,N_34509,N_30613);
nor U35184 (N_35184,N_32061,N_31677);
xnor U35185 (N_35185,N_33326,N_33216);
or U35186 (N_35186,N_33275,N_30262);
nand U35187 (N_35187,N_32685,N_32490);
or U35188 (N_35188,N_33897,N_34335);
or U35189 (N_35189,N_34012,N_32969);
nor U35190 (N_35190,N_32504,N_34680);
xnor U35191 (N_35191,N_34983,N_34283);
or U35192 (N_35192,N_34408,N_30758);
or U35193 (N_35193,N_34065,N_33839);
nor U35194 (N_35194,N_33499,N_31711);
nand U35195 (N_35195,N_30947,N_33962);
xor U35196 (N_35196,N_30044,N_30029);
and U35197 (N_35197,N_30873,N_33856);
xor U35198 (N_35198,N_33124,N_33193);
and U35199 (N_35199,N_30841,N_31954);
xnor U35200 (N_35200,N_32107,N_31909);
or U35201 (N_35201,N_31484,N_30941);
nor U35202 (N_35202,N_32300,N_34726);
or U35203 (N_35203,N_31913,N_30428);
nand U35204 (N_35204,N_31494,N_31986);
nand U35205 (N_35205,N_31292,N_31667);
or U35206 (N_35206,N_32467,N_30658);
or U35207 (N_35207,N_34163,N_34952);
and U35208 (N_35208,N_30931,N_34937);
nand U35209 (N_35209,N_32508,N_34139);
nand U35210 (N_35210,N_32401,N_30300);
nand U35211 (N_35211,N_34042,N_34700);
xor U35212 (N_35212,N_31214,N_30271);
nor U35213 (N_35213,N_34876,N_33782);
xor U35214 (N_35214,N_31011,N_33267);
nor U35215 (N_35215,N_31734,N_33208);
xor U35216 (N_35216,N_31048,N_31107);
or U35217 (N_35217,N_32013,N_31317);
or U35218 (N_35218,N_34708,N_30542);
nand U35219 (N_35219,N_33809,N_30539);
nand U35220 (N_35220,N_34639,N_33073);
xnor U35221 (N_35221,N_31149,N_31611);
nand U35222 (N_35222,N_30704,N_31466);
nor U35223 (N_35223,N_32385,N_34423);
nand U35224 (N_35224,N_32060,N_32093);
or U35225 (N_35225,N_33868,N_34237);
nand U35226 (N_35226,N_32309,N_30231);
xnor U35227 (N_35227,N_30625,N_30897);
nand U35228 (N_35228,N_34173,N_30191);
nand U35229 (N_35229,N_31851,N_33644);
and U35230 (N_35230,N_30751,N_30755);
nor U35231 (N_35231,N_31063,N_33921);
and U35232 (N_35232,N_32449,N_32356);
nor U35233 (N_35233,N_33936,N_34281);
or U35234 (N_35234,N_30681,N_31125);
and U35235 (N_35235,N_32122,N_34650);
xor U35236 (N_35236,N_30229,N_33672);
nor U35237 (N_35237,N_30750,N_34317);
or U35238 (N_35238,N_32345,N_31268);
nand U35239 (N_35239,N_30531,N_34384);
xnor U35240 (N_35240,N_31508,N_30399);
nand U35241 (N_35241,N_34392,N_33406);
xor U35242 (N_35242,N_31791,N_34847);
xor U35243 (N_35243,N_30986,N_30078);
or U35244 (N_35244,N_33350,N_30575);
nand U35245 (N_35245,N_32430,N_30239);
xor U35246 (N_35246,N_33448,N_33377);
or U35247 (N_35247,N_30268,N_33652);
or U35248 (N_35248,N_34389,N_32602);
or U35249 (N_35249,N_30381,N_30936);
xnor U35250 (N_35250,N_33777,N_31844);
or U35251 (N_35251,N_32147,N_33480);
and U35252 (N_35252,N_31397,N_32701);
nor U35253 (N_35253,N_34448,N_33610);
and U35254 (N_35254,N_32120,N_31600);
xnor U35255 (N_35255,N_32516,N_32386);
nand U35256 (N_35256,N_31418,N_32237);
xnor U35257 (N_35257,N_30313,N_31309);
or U35258 (N_35258,N_30990,N_32908);
nand U35259 (N_35259,N_32798,N_34138);
nor U35260 (N_35260,N_34763,N_30740);
or U35261 (N_35261,N_34713,N_32561);
nor U35262 (N_35262,N_30959,N_31892);
nor U35263 (N_35263,N_33983,N_33832);
nor U35264 (N_35264,N_33504,N_31942);
xnor U35265 (N_35265,N_30025,N_34969);
nand U35266 (N_35266,N_30545,N_34117);
nor U35267 (N_35267,N_32132,N_30149);
or U35268 (N_35268,N_32863,N_30384);
and U35269 (N_35269,N_33999,N_31819);
nor U35270 (N_35270,N_31654,N_31474);
or U35271 (N_35271,N_33943,N_34044);
nor U35272 (N_35272,N_30773,N_34747);
nor U35273 (N_35273,N_33354,N_30334);
xor U35274 (N_35274,N_34106,N_31562);
and U35275 (N_35275,N_34536,N_33089);
xnor U35276 (N_35276,N_32314,N_31530);
and U35277 (N_35277,N_32519,N_33833);
nand U35278 (N_35278,N_30953,N_34107);
nor U35279 (N_35279,N_33707,N_30768);
or U35280 (N_35280,N_32987,N_33612);
nor U35281 (N_35281,N_32073,N_34947);
and U35282 (N_35282,N_33023,N_30281);
nor U35283 (N_35283,N_32463,N_34825);
and U35284 (N_35284,N_31394,N_33517);
nor U35285 (N_35285,N_34164,N_34229);
and U35286 (N_35286,N_32493,N_34733);
or U35287 (N_35287,N_34334,N_30097);
xnor U35288 (N_35288,N_30588,N_32212);
or U35289 (N_35289,N_30514,N_30030);
nand U35290 (N_35290,N_30533,N_33296);
nand U35291 (N_35291,N_30100,N_31708);
or U35292 (N_35292,N_32533,N_32569);
and U35293 (N_35293,N_31447,N_30922);
xor U35294 (N_35294,N_32466,N_34402);
or U35295 (N_35295,N_31083,N_31425);
and U35296 (N_35296,N_31303,N_30252);
or U35297 (N_35297,N_32780,N_31789);
and U35298 (N_35298,N_34040,N_34606);
or U35299 (N_35299,N_33173,N_31579);
or U35300 (N_35300,N_32004,N_30118);
xnor U35301 (N_35301,N_30450,N_30883);
nor U35302 (N_35302,N_33456,N_31261);
or U35303 (N_35303,N_32104,N_31284);
or U35304 (N_35304,N_31874,N_31045);
xnor U35305 (N_35305,N_31390,N_32960);
nor U35306 (N_35306,N_31324,N_30822);
and U35307 (N_35307,N_30171,N_30429);
nand U35308 (N_35308,N_30565,N_33584);
nor U35309 (N_35309,N_31142,N_34540);
nor U35310 (N_35310,N_30182,N_30629);
xor U35311 (N_35311,N_34902,N_34033);
and U35312 (N_35312,N_31427,N_30911);
xnor U35313 (N_35313,N_30217,N_32677);
or U35314 (N_35314,N_30339,N_31137);
nand U35315 (N_35315,N_33830,N_33581);
xnor U35316 (N_35316,N_33760,N_31491);
nand U35317 (N_35317,N_34330,N_31391);
and U35318 (N_35318,N_33585,N_31968);
nor U35319 (N_35319,N_32295,N_32354);
nor U35320 (N_35320,N_33370,N_32285);
and U35321 (N_35321,N_34574,N_32620);
and U35322 (N_35322,N_32760,N_32026);
nand U35323 (N_35323,N_30155,N_31076);
or U35324 (N_35324,N_34375,N_34218);
and U35325 (N_35325,N_30784,N_33715);
or U35326 (N_35326,N_31523,N_30102);
or U35327 (N_35327,N_34855,N_32607);
and U35328 (N_35328,N_32818,N_33817);
nand U35329 (N_35329,N_34258,N_30511);
nor U35330 (N_35330,N_30688,N_33508);
nand U35331 (N_35331,N_34933,N_32458);
xor U35332 (N_35332,N_32250,N_34666);
xor U35333 (N_35333,N_34048,N_30361);
and U35334 (N_35334,N_31797,N_34074);
and U35335 (N_35335,N_33304,N_32081);
xor U35336 (N_35336,N_32919,N_34565);
and U35337 (N_35337,N_32197,N_32433);
nand U35338 (N_35338,N_33298,N_33392);
nand U35339 (N_35339,N_31961,N_32706);
xnor U35340 (N_35340,N_30985,N_33486);
or U35341 (N_35341,N_34846,N_33941);
nand U35342 (N_35342,N_33388,N_32913);
nand U35343 (N_35343,N_33162,N_31437);
nor U35344 (N_35344,N_34634,N_34496);
or U35345 (N_35345,N_33805,N_31897);
xor U35346 (N_35346,N_31974,N_34771);
xnor U35347 (N_35347,N_30085,N_34626);
nand U35348 (N_35348,N_34110,N_32100);
nor U35349 (N_35349,N_30265,N_31945);
xnor U35350 (N_35350,N_31542,N_34207);
nor U35351 (N_35351,N_31420,N_31572);
xnor U35352 (N_35352,N_33963,N_30520);
or U35353 (N_35353,N_34875,N_33474);
or U35354 (N_35354,N_30521,N_33128);
and U35355 (N_35355,N_30394,N_31911);
nand U35356 (N_35356,N_31973,N_34146);
and U35357 (N_35357,N_32587,N_32886);
xnor U35358 (N_35358,N_34889,N_30360);
xor U35359 (N_35359,N_33196,N_32618);
or U35360 (N_35360,N_31683,N_30786);
nor U35361 (N_35361,N_34897,N_34046);
and U35362 (N_35362,N_32043,N_33104);
nor U35363 (N_35363,N_31768,N_33217);
and U35364 (N_35364,N_32189,N_30202);
nor U35365 (N_35365,N_32741,N_34662);
xnor U35366 (N_35366,N_30156,N_32326);
and U35367 (N_35367,N_34470,N_32954);
nand U35368 (N_35368,N_32130,N_31402);
nor U35369 (N_35369,N_31332,N_30567);
xor U35370 (N_35370,N_34344,N_34051);
nand U35371 (N_35371,N_33428,N_32750);
and U35372 (N_35372,N_32898,N_34501);
and U35373 (N_35373,N_30316,N_33690);
and U35374 (N_35374,N_32379,N_30189);
and U35375 (N_35375,N_33010,N_32912);
and U35376 (N_35376,N_33602,N_34235);
nand U35377 (N_35377,N_32378,N_30151);
nor U35378 (N_35378,N_33297,N_32119);
or U35379 (N_35379,N_30791,N_33692);
or U35380 (N_35380,N_32795,N_30040);
xnor U35381 (N_35381,N_34493,N_30280);
nor U35382 (N_35382,N_30375,N_33653);
or U35383 (N_35383,N_34527,N_30130);
nand U35384 (N_35384,N_32383,N_34754);
nor U35385 (N_35385,N_31240,N_32633);
xor U35386 (N_35386,N_33000,N_33513);
nor U35387 (N_35387,N_33569,N_33253);
nor U35388 (N_35388,N_32070,N_31406);
and U35389 (N_35389,N_33147,N_32310);
and U35390 (N_35390,N_30258,N_33704);
nand U35391 (N_35391,N_31753,N_30403);
and U35392 (N_35392,N_31323,N_32283);
and U35393 (N_35393,N_34602,N_31891);
nand U35394 (N_35394,N_34585,N_33496);
and U35395 (N_35395,N_34691,N_32206);
nand U35396 (N_35396,N_34123,N_30965);
and U35397 (N_35397,N_31610,N_32828);
and U35398 (N_35398,N_33554,N_31087);
and U35399 (N_35399,N_33186,N_30298);
or U35400 (N_35400,N_32321,N_31464);
and U35401 (N_35401,N_30951,N_30310);
or U35402 (N_35402,N_31767,N_31289);
xnor U35403 (N_35403,N_32968,N_30508);
xor U35404 (N_35404,N_30734,N_32796);
and U35405 (N_35405,N_33725,N_31409);
nor U35406 (N_35406,N_30433,N_31801);
nand U35407 (N_35407,N_30410,N_34406);
nor U35408 (N_35408,N_31669,N_30586);
nor U35409 (N_35409,N_31747,N_30718);
and U35410 (N_35410,N_30318,N_31858);
or U35411 (N_35411,N_33950,N_32395);
xnor U35412 (N_35412,N_33289,N_32882);
and U35413 (N_35413,N_32901,N_30338);
or U35414 (N_35414,N_30477,N_32512);
xor U35415 (N_35415,N_33457,N_31059);
and U35416 (N_35416,N_30284,N_33062);
or U35417 (N_35417,N_34688,N_34415);
nor U35418 (N_35418,N_31662,N_31918);
and U35419 (N_35419,N_31445,N_30139);
nand U35420 (N_35420,N_30103,N_31628);
nor U35421 (N_35421,N_30769,N_34021);
xnor U35422 (N_35422,N_30179,N_31805);
and U35423 (N_35423,N_30411,N_34434);
nor U35424 (N_35424,N_31925,N_33067);
xor U35425 (N_35425,N_31110,N_32588);
nor U35426 (N_35426,N_30094,N_33568);
xnor U35427 (N_35427,N_30903,N_34228);
and U35428 (N_35428,N_34016,N_31064);
xor U35429 (N_35429,N_31031,N_32505);
nor U35430 (N_35430,N_34545,N_32922);
nand U35431 (N_35431,N_31988,N_33774);
xor U35432 (N_35432,N_31314,N_34950);
nor U35433 (N_35433,N_34214,N_30016);
and U35434 (N_35434,N_34206,N_34414);
nand U35435 (N_35435,N_32459,N_34013);
xor U35436 (N_35436,N_34714,N_34226);
nor U35437 (N_35437,N_33039,N_32590);
or U35438 (N_35438,N_34913,N_33240);
nor U35439 (N_35439,N_34821,N_31236);
nand U35440 (N_35440,N_31179,N_32251);
nand U35441 (N_35441,N_33077,N_30020);
or U35442 (N_35442,N_34364,N_32353);
or U35443 (N_35443,N_30816,N_31403);
nor U35444 (N_35444,N_34584,N_32156);
nor U35445 (N_35445,N_31356,N_32625);
and U35446 (N_35446,N_30920,N_33658);
nor U35447 (N_35447,N_34332,N_31567);
or U35448 (N_35448,N_30862,N_33638);
xnor U35449 (N_35449,N_34549,N_33553);
nor U35450 (N_35450,N_31569,N_33970);
nor U35451 (N_35451,N_32934,N_33027);
or U35452 (N_35452,N_31224,N_30927);
or U35453 (N_35453,N_33931,N_31924);
and U35454 (N_35454,N_33100,N_32190);
nor U35455 (N_35455,N_33319,N_30236);
nor U35456 (N_35456,N_34184,N_34753);
nor U35457 (N_35457,N_32437,N_31376);
and U35458 (N_35458,N_32033,N_33714);
nor U35459 (N_35459,N_34233,N_33290);
nand U35460 (N_35460,N_33902,N_33650);
nor U35461 (N_35461,N_33682,N_33601);
or U35462 (N_35462,N_31694,N_32144);
xnor U35463 (N_35463,N_32135,N_33929);
nand U35464 (N_35464,N_32752,N_34935);
nand U35465 (N_35465,N_34511,N_30749);
or U35466 (N_35466,N_31652,N_33740);
nor U35467 (N_35467,N_31576,N_30594);
xnor U35468 (N_35468,N_33965,N_30219);
nand U35469 (N_35469,N_30225,N_33635);
xor U35470 (N_35470,N_33563,N_32078);
nor U35471 (N_35471,N_34959,N_32054);
or U35472 (N_35472,N_34617,N_32200);
and U35473 (N_35473,N_32801,N_31176);
nor U35474 (N_35474,N_34614,N_32945);
and U35475 (N_35475,N_34028,N_31796);
xnor U35476 (N_35476,N_32258,N_34605);
nand U35477 (N_35477,N_33735,N_31455);
and U35478 (N_35478,N_34552,N_33851);
nor U35479 (N_35479,N_34234,N_31207);
or U35480 (N_35480,N_33857,N_32647);
and U35481 (N_35481,N_33906,N_31472);
or U35482 (N_35482,N_32170,N_34604);
nand U35483 (N_35483,N_33528,N_33222);
and U35484 (N_35484,N_32793,N_31069);
xnor U35485 (N_35485,N_32833,N_32876);
nor U35486 (N_35486,N_32268,N_31539);
or U35487 (N_35487,N_33048,N_34532);
nand U35488 (N_35488,N_33022,N_33566);
xor U35489 (N_35489,N_32782,N_31758);
nand U35490 (N_35490,N_33242,N_32371);
and U35491 (N_35491,N_30147,N_34393);
nor U35492 (N_35492,N_32609,N_33801);
xnor U35493 (N_35493,N_30036,N_30592);
and U35494 (N_35494,N_34119,N_30548);
or U35495 (N_35495,N_30948,N_34737);
or U35496 (N_35496,N_33309,N_33985);
xnor U35497 (N_35497,N_33243,N_34522);
nor U35498 (N_35498,N_33792,N_34920);
xor U35499 (N_35499,N_32209,N_31671);
nor U35500 (N_35500,N_33961,N_34310);
and U35501 (N_35501,N_33260,N_34469);
nand U35502 (N_35502,N_32671,N_34054);
or U35503 (N_35503,N_32703,N_33478);
nor U35504 (N_35504,N_30185,N_30672);
nand U35505 (N_35505,N_34140,N_34273);
or U35506 (N_35506,N_34538,N_30703);
nor U35507 (N_35507,N_34516,N_33356);
and U35508 (N_35508,N_30073,N_32979);
xnor U35509 (N_35509,N_34851,N_32905);
nand U35510 (N_35510,N_34512,N_30196);
xor U35511 (N_35511,N_30110,N_34868);
and U35512 (N_35512,N_31296,N_34380);
nor U35513 (N_35513,N_30146,N_32304);
xor U35514 (N_35514,N_30160,N_30224);
or U35515 (N_35515,N_31777,N_31290);
nor U35516 (N_35516,N_32362,N_32484);
or U35517 (N_35517,N_34161,N_33286);
nand U35518 (N_35518,N_34670,N_30107);
xor U35519 (N_35519,N_31646,N_30343);
nor U35520 (N_35520,N_31095,N_30591);
nand U35521 (N_35521,N_33731,N_30908);
or U35522 (N_35522,N_33806,N_34045);
or U35523 (N_35523,N_33915,N_30181);
nand U35524 (N_35524,N_31651,N_32090);
nor U35525 (N_35525,N_30494,N_34292);
and U35526 (N_35526,N_30652,N_32694);
and U35527 (N_35527,N_33020,N_30812);
and U35528 (N_35528,N_34504,N_30446);
nor U35529 (N_35529,N_33925,N_33401);
nor U35530 (N_35530,N_30101,N_32866);
nor U35531 (N_35531,N_30639,N_31022);
nand U35532 (N_35532,N_30476,N_33649);
xnor U35533 (N_35533,N_32101,N_34800);
and U35534 (N_35534,N_30711,N_34739);
nand U35535 (N_35535,N_30350,N_31886);
nand U35536 (N_35536,N_33139,N_31326);
nand U35537 (N_35537,N_33539,N_31800);
xnor U35538 (N_35538,N_32679,N_31907);
xor U35539 (N_35539,N_31099,N_32403);
xor U35540 (N_35540,N_33103,N_30120);
nor U35541 (N_35541,N_32288,N_33694);
nor U35542 (N_35542,N_30952,N_32334);
and U35543 (N_35543,N_33307,N_32672);
xnor U35544 (N_35544,N_32704,N_31273);
or U35545 (N_35545,N_31802,N_31308);
xnor U35546 (N_35546,N_34945,N_34559);
xnor U35547 (N_35547,N_34486,N_31552);
or U35548 (N_35548,N_31917,N_30669);
or U35549 (N_35549,N_34848,N_34582);
nor U35550 (N_35550,N_32293,N_30444);
or U35551 (N_35551,N_31175,N_32089);
nor U35552 (N_35552,N_32617,N_34633);
and U35553 (N_35553,N_33623,N_34961);
and U35554 (N_35554,N_31003,N_30500);
or U35555 (N_35555,N_34791,N_34717);
and U35556 (N_35556,N_34951,N_33873);
nand U35557 (N_35557,N_33849,N_33885);
nor U35558 (N_35558,N_30095,N_32769);
nand U35559 (N_35559,N_33316,N_31543);
xor U35560 (N_35560,N_33151,N_32523);
nand U35561 (N_35561,N_32718,N_30379);
and U35562 (N_35562,N_30848,N_32932);
and U35563 (N_35563,N_32528,N_31384);
xor U35564 (N_35564,N_34481,N_31603);
xnor U35565 (N_35565,N_33241,N_34564);
nand U35566 (N_35566,N_31915,N_34580);
or U35567 (N_35567,N_30372,N_32977);
nor U35568 (N_35568,N_33609,N_34641);
xor U35569 (N_35569,N_31310,N_30678);
nand U35570 (N_35570,N_30855,N_30165);
or U35571 (N_35571,N_30408,N_31638);
nor U35572 (N_35572,N_31726,N_32229);
nor U35573 (N_35573,N_32929,N_30434);
or U35574 (N_35574,N_32785,N_34832);
nor U35575 (N_35575,N_30049,N_33150);
nand U35576 (N_35576,N_32845,N_33498);
and U35577 (N_35577,N_33546,N_34862);
xnor U35578 (N_35578,N_33552,N_34035);
xor U35579 (N_35579,N_33069,N_34795);
xor U35580 (N_35580,N_31254,N_33590);
or U35581 (N_35581,N_31922,N_31556);
nor U35582 (N_35582,N_32594,N_33986);
nand U35583 (N_35583,N_32656,N_32946);
xnor U35584 (N_35584,N_32415,N_34784);
or U35585 (N_35585,N_30835,N_31609);
xor U35586 (N_35586,N_32823,N_32691);
or U35587 (N_35587,N_33246,N_30892);
or U35588 (N_35588,N_31693,N_31962);
and U35589 (N_35589,N_30605,N_30723);
nand U35590 (N_35590,N_31301,N_31315);
or U35591 (N_35591,N_34069,N_33604);
xor U35592 (N_35592,N_33949,N_33667);
or U35593 (N_35593,N_33521,N_31463);
nand U35594 (N_35594,N_33861,N_33621);
and U35595 (N_35595,N_32699,N_33850);
nor U35596 (N_35596,N_32359,N_33660);
or U35597 (N_35597,N_31887,N_34009);
or U35598 (N_35598,N_34144,N_30254);
nor U35599 (N_35599,N_31478,N_32400);
nand U35600 (N_35600,N_34197,N_31719);
xnor U35601 (N_35601,N_33034,N_32011);
and U35602 (N_35602,N_30062,N_32440);
nor U35603 (N_35603,N_30643,N_32065);
nor U35604 (N_35604,N_33558,N_31027);
and U35605 (N_35605,N_33688,N_34204);
or U35606 (N_35606,N_32211,N_34859);
and U35607 (N_35607,N_30329,N_31165);
nand U35608 (N_35608,N_32844,N_33108);
and U35609 (N_35609,N_30440,N_30466);
nand U35610 (N_35610,N_32327,N_32053);
xor U35611 (N_35611,N_32207,N_34989);
nor U35612 (N_35612,N_34036,N_32322);
nand U35613 (N_35613,N_31424,N_31111);
nor U35614 (N_35614,N_31364,N_33913);
nor U35615 (N_35615,N_32280,N_31685);
and U35616 (N_35616,N_31504,N_31043);
xor U35617 (N_35617,N_30414,N_33405);
nand U35618 (N_35618,N_32071,N_32010);
xor U35619 (N_35619,N_31944,N_30633);
and U35620 (N_35620,N_34178,N_31633);
nor U35621 (N_35621,N_33838,N_31931);
and U35622 (N_35622,N_31910,N_31313);
xnor U35623 (N_35623,N_34663,N_31465);
nand U35624 (N_35624,N_33329,N_30425);
nand U35625 (N_35625,N_32227,N_31875);
or U35626 (N_35626,N_31241,N_30368);
xnor U35627 (N_35627,N_34452,N_34874);
and U35628 (N_35628,N_33026,N_30154);
and U35629 (N_35629,N_31071,N_31479);
or U35630 (N_35630,N_31873,N_34112);
and U35631 (N_35631,N_31015,N_32778);
xnor U35632 (N_35632,N_31092,N_34979);
and U35633 (N_35633,N_30935,N_34271);
and U35634 (N_35634,N_33693,N_32978);
or U35635 (N_35635,N_34542,N_31269);
and U35636 (N_35636,N_32487,N_34526);
nand U35637 (N_35637,N_33107,N_30760);
nor U35638 (N_35638,N_33989,N_33848);
xnor U35639 (N_35639,N_30589,N_30517);
xnor U35640 (N_35640,N_34973,N_34223);
xor U35641 (N_35641,N_33520,N_31795);
nor U35642 (N_35642,N_31034,N_30707);
or U35643 (N_35643,N_30641,N_33315);
or U35644 (N_35644,N_31591,N_31147);
or U35645 (N_35645,N_34141,N_33185);
nor U35646 (N_35646,N_34769,N_33959);
nand U35647 (N_35647,N_30725,N_34290);
or U35648 (N_35648,N_34108,N_32117);
xnor U35649 (N_35649,N_33327,N_31981);
nor U35650 (N_35650,N_31370,N_30472);
nor U35651 (N_35651,N_32526,N_30233);
or U35652 (N_35652,N_31678,N_33368);
or U35653 (N_35653,N_30255,N_30330);
or U35654 (N_35654,N_31227,N_31180);
xor U35655 (N_35655,N_33352,N_34906);
nand U35656 (N_35656,N_32809,N_31281);
nand U35657 (N_35657,N_32575,N_33645);
nand U35658 (N_35658,N_33677,N_31607);
and U35659 (N_35659,N_30468,N_30485);
xor U35660 (N_35660,N_30851,N_30162);
and U35661 (N_35661,N_33825,N_34872);
xor U35662 (N_35662,N_31721,N_30295);
and U35663 (N_35663,N_33030,N_31598);
and U35664 (N_35664,N_33909,N_34946);
nand U35665 (N_35665,N_32622,N_30798);
or U35666 (N_35666,N_33732,N_32974);
xor U35667 (N_35667,N_34120,N_30793);
nor U35668 (N_35668,N_30805,N_34297);
nand U35669 (N_35669,N_32495,N_31632);
or U35670 (N_35670,N_31160,N_34374);
or U35671 (N_35671,N_33664,N_34823);
xnor U35672 (N_35672,N_33761,N_31191);
xnor U35673 (N_35673,N_32194,N_33955);
or U35674 (N_35674,N_32020,N_34801);
xnor U35675 (N_35675,N_32428,N_30436);
nor U35676 (N_35676,N_33183,N_34284);
or U35677 (N_35677,N_31133,N_31153);
or U35678 (N_35678,N_33591,N_33182);
or U35679 (N_35679,N_31803,N_33699);
xor U35680 (N_35680,N_30312,N_30611);
nor U35681 (N_35681,N_34611,N_32159);
xnor U35682 (N_35682,N_32971,N_32306);
and U35683 (N_35683,N_34478,N_31612);
nand U35684 (N_35684,N_32116,N_30766);
xor U35685 (N_35685,N_31361,N_32086);
nor U35686 (N_35686,N_30212,N_33131);
nand U35687 (N_35687,N_30293,N_33203);
and U35688 (N_35688,N_34213,N_34915);
nor U35689 (N_35689,N_33134,N_32366);
nand U35690 (N_35690,N_31825,N_30337);
xor U35691 (N_35691,N_34285,N_32501);
and U35692 (N_35692,N_30697,N_30137);
and U35693 (N_35693,N_32413,N_34436);
nand U35694 (N_35694,N_30180,N_33333);
xnor U35695 (N_35695,N_34300,N_34064);
xor U35696 (N_35696,N_31631,N_34623);
xnor U35697 (N_35697,N_34232,N_30090);
nor U35698 (N_35698,N_32184,N_34314);
nand U35699 (N_35699,N_31927,N_33453);
or U35700 (N_35700,N_32063,N_31625);
and U35701 (N_35701,N_34530,N_32721);
or U35702 (N_35702,N_33360,N_33946);
nor U35703 (N_35703,N_32900,N_30091);
or U35704 (N_35704,N_33076,N_34787);
xor U35705 (N_35705,N_31751,N_32196);
nor U35706 (N_35706,N_33044,N_30844);
nor U35707 (N_35707,N_34456,N_30995);
xnor U35708 (N_35708,N_31838,N_34175);
xor U35709 (N_35709,N_30754,N_33464);
xnor U35710 (N_35710,N_30071,N_34477);
xor U35711 (N_35711,N_30807,N_31404);
nand U35712 (N_35712,N_32372,N_30082);
xor U35713 (N_35713,N_33078,N_31746);
nand U35714 (N_35714,N_30096,N_30055);
nand U35715 (N_35715,N_30846,N_30615);
and U35716 (N_35716,N_34272,N_31380);
and U35717 (N_35717,N_34845,N_31656);
nor U35718 (N_35718,N_33175,N_33998);
or U35719 (N_35719,N_34347,N_32631);
and U35720 (N_35720,N_34351,N_33087);
xor U35721 (N_35721,N_34311,N_33608);
nor U35722 (N_35722,N_31467,N_34096);
or U35723 (N_35723,N_30820,N_32320);
or U35724 (N_35724,N_31620,N_30398);
nand U35725 (N_35725,N_33626,N_31706);
nand U35726 (N_35726,N_30288,N_33670);
nor U35727 (N_35727,N_34359,N_34554);
or U35728 (N_35728,N_32547,N_31680);
xor U35729 (N_35729,N_30898,N_32582);
and U35730 (N_35730,N_31335,N_32290);
and U35731 (N_35731,N_30218,N_34901);
nor U35732 (N_35732,N_32859,N_32854);
or U35733 (N_35733,N_33647,N_34627);
xnor U35734 (N_35734,N_33958,N_33860);
xnor U35735 (N_35735,N_30651,N_34465);
nor U35736 (N_35736,N_33443,N_31088);
or U35737 (N_35737,N_34212,N_34816);
and U35738 (N_35738,N_33948,N_32198);
or U35739 (N_35739,N_30680,N_31890);
nand U35740 (N_35740,N_31220,N_30413);
nor U35741 (N_35741,N_33811,N_31182);
xnor U35742 (N_35742,N_33133,N_30064);
nand U35743 (N_35743,N_31246,N_34071);
nand U35744 (N_35744,N_33017,N_30731);
or U35745 (N_35745,N_34648,N_33200);
and U35746 (N_35746,N_31636,N_32792);
nor U35747 (N_35747,N_30039,N_30746);
nor U35748 (N_35748,N_30627,N_30685);
or U35749 (N_35749,N_34269,N_33771);
nand U35750 (N_35750,N_31518,N_32805);
and U35751 (N_35751,N_33445,N_30532);
nand U35752 (N_35752,N_34241,N_31824);
xnor U35753 (N_35753,N_31604,N_34262);
nand U35754 (N_35754,N_33935,N_30365);
xnor U35755 (N_35755,N_34391,N_34199);
or U35756 (N_35756,N_33633,N_32514);
nand U35757 (N_35757,N_30868,N_32203);
and U35758 (N_35758,N_33778,N_33180);
nand U35759 (N_35759,N_34924,N_33024);
xor U35760 (N_35760,N_31449,N_33747);
nor U35761 (N_35761,N_31934,N_30014);
nand U35762 (N_35762,N_34475,N_31156);
or U35763 (N_35763,N_34975,N_33828);
or U35764 (N_35764,N_32762,N_34998);
nor U35765 (N_35765,N_32308,N_31028);
and U35766 (N_35766,N_33583,N_32096);
or U35767 (N_35767,N_34439,N_31081);
and U35768 (N_35768,N_33560,N_32853);
xnor U35769 (N_35769,N_31798,N_33923);
and U35770 (N_35770,N_34741,N_31201);
nor U35771 (N_35771,N_34756,N_34537);
or U35772 (N_35772,N_33636,N_30745);
and U35773 (N_35773,N_33422,N_34653);
nor U35774 (N_35774,N_31696,N_31987);
xnor U35775 (N_35775,N_34598,N_32723);
nand U35776 (N_35776,N_30447,N_31930);
nand U35777 (N_35777,N_33964,N_30946);
nor U35778 (N_35778,N_32579,N_31054);
xnor U35779 (N_35779,N_33537,N_32695);
and U35780 (N_35780,N_33995,N_31033);
and U35781 (N_35781,N_34073,N_31018);
xor U35782 (N_35782,N_32548,N_30549);
xor U35783 (N_35783,N_34279,N_34636);
nand U35784 (N_35784,N_34494,N_34729);
and U35785 (N_35785,N_31829,N_33375);
and U35786 (N_35786,N_31237,N_33567);
xnor U35787 (N_35787,N_32872,N_33038);
nand U35788 (N_35788,N_34350,N_32226);
and U35789 (N_35789,N_30084,N_33407);
xnor U35790 (N_35790,N_30742,N_30238);
or U35791 (N_35791,N_31834,N_30840);
nor U35792 (N_35792,N_30068,N_34428);
and U35793 (N_35793,N_32984,N_30776);
nand U35794 (N_35794,N_32244,N_30161);
nor U35795 (N_35795,N_33143,N_33956);
or U35796 (N_35796,N_31655,N_33631);
or U35797 (N_35797,N_33322,N_30081);
nand U35798 (N_35798,N_34333,N_32399);
nand U35799 (N_35799,N_32279,N_31668);
xnor U35800 (N_35800,N_33052,N_30465);
and U35801 (N_35801,N_30510,N_33877);
nand U35802 (N_35802,N_34052,N_30557);
nand U35803 (N_35803,N_32649,N_34383);
and U35804 (N_35804,N_32082,N_34426);
or U35805 (N_35805,N_30602,N_30461);
xor U35806 (N_35806,N_32756,N_34440);
nand U35807 (N_35807,N_30222,N_30975);
nor U35808 (N_35808,N_34134,N_32639);
and U35809 (N_35809,N_32478,N_33043);
nand U35810 (N_35810,N_30223,N_30527);
nand U35811 (N_35811,N_31570,N_32612);
nor U35812 (N_35812,N_33910,N_32850);
nand U35813 (N_35813,N_34459,N_31820);
nand U35814 (N_35814,N_34799,N_31367);
nand U35815 (N_35815,N_32890,N_30918);
or U35816 (N_35816,N_31928,N_34607);
nand U35817 (N_35817,N_32181,N_30905);
or U35818 (N_35818,N_33046,N_31451);
nor U35819 (N_35819,N_32032,N_34301);
nor U35820 (N_35820,N_30079,N_34977);
nor U35821 (N_35821,N_31348,N_34302);
xor U35822 (N_35822,N_33166,N_33068);
xnor U35823 (N_35823,N_34129,N_33974);
or U35824 (N_35824,N_32103,N_31733);
or U35825 (N_35825,N_33502,N_31766);
xnor U35826 (N_35826,N_31577,N_34624);
nor U35827 (N_35827,N_32666,N_33119);
and U35828 (N_35828,N_30845,N_30220);
or U35829 (N_35829,N_32643,N_30714);
nand U35830 (N_35830,N_34949,N_30821);
or U35831 (N_35831,N_30663,N_32145);
or U35832 (N_35832,N_32180,N_31817);
xnor U35833 (N_35833,N_34958,N_32727);
nand U35834 (N_35834,N_31300,N_33090);
and U35835 (N_35835,N_32842,N_33896);
or U35836 (N_35836,N_33763,N_33281);
or U35837 (N_35837,N_30246,N_34553);
and U35838 (N_35838,N_32051,N_31024);
xor U35839 (N_35839,N_31846,N_32915);
or U35840 (N_35840,N_31439,N_32451);
xor U35841 (N_35841,N_31929,N_33501);
and U35842 (N_35842,N_34417,N_31554);
and U35843 (N_35843,N_33272,N_33481);
nand U35844 (N_35844,N_33807,N_33161);
or U35845 (N_35845,N_33120,N_30981);
and U35846 (N_35846,N_31521,N_33091);
xnor U35847 (N_35847,N_32307,N_30509);
nand U35848 (N_35848,N_34775,N_34525);
or U35849 (N_35849,N_34067,N_30353);
nor U35850 (N_35850,N_31762,N_30387);
nor U35851 (N_35851,N_31499,N_31114);
or U35852 (N_35852,N_34011,N_34205);
and U35853 (N_35853,N_30356,N_33355);
nand U35854 (N_35854,N_34167,N_33934);
and U35855 (N_35855,N_33820,N_30172);
nand U35856 (N_35856,N_33990,N_32347);
xor U35857 (N_35857,N_33914,N_30515);
and U35858 (N_35858,N_31101,N_32910);
nand U35859 (N_35859,N_34751,N_30809);
or U35860 (N_35860,N_34321,N_30317);
nand U35861 (N_35861,N_34405,N_33064);
or U35862 (N_35862,N_33573,N_31781);
nor U35863 (N_35863,N_33912,N_32178);
xor U35864 (N_35864,N_34488,N_31811);
nor U35865 (N_35865,N_33571,N_34340);
xor U35866 (N_35866,N_31975,N_34320);
nand U35867 (N_35867,N_31017,N_33579);
nor U35868 (N_35868,N_34299,N_33146);
and U35869 (N_35869,N_31588,N_32410);
or U35870 (N_35870,N_32423,N_31168);
or U35871 (N_35871,N_31216,N_32059);
nor U35872 (N_35872,N_33898,N_30022);
or U35873 (N_35873,N_31266,N_31980);
nand U35874 (N_35874,N_33523,N_30263);
nor U35875 (N_35875,N_31705,N_33476);
nor U35876 (N_35876,N_33122,N_32019);
and U35877 (N_35877,N_32357,N_34378);
and U35878 (N_35878,N_31333,N_31396);
nand U35879 (N_35879,N_30679,N_31511);
and U35880 (N_35880,N_30547,N_31794);
xnor U35881 (N_35881,N_30140,N_32248);
xor U35882 (N_35882,N_32435,N_30958);
nor U35883 (N_35883,N_31381,N_33337);
xor U35884 (N_35884,N_31104,N_31010);
or U35885 (N_35885,N_30026,N_32817);
xnor U35886 (N_35886,N_33978,N_30756);
nand U35887 (N_35887,N_31866,N_34329);
nor U35888 (N_35888,N_30909,N_32036);
and U35889 (N_35889,N_31122,N_32511);
and U35890 (N_35890,N_30783,N_34370);
nand U35891 (N_35891,N_31410,N_30153);
or U35892 (N_35892,N_31908,N_32163);
xnor U35893 (N_35893,N_33063,N_31248);
nand U35894 (N_35894,N_30423,N_31371);
nand U35895 (N_35895,N_31792,N_31438);
nor U35896 (N_35896,N_32460,N_30503);
nor U35897 (N_35897,N_33473,N_32673);
nor U35898 (N_35898,N_31821,N_32924);
and U35899 (N_35899,N_33646,N_32496);
or U35900 (N_35900,N_30665,N_33519);
nor U35901 (N_35901,N_34111,N_31342);
or U35902 (N_35902,N_32001,N_34419);
xnor U35903 (N_35903,N_31100,N_32957);
xnor U35904 (N_35904,N_32281,N_30027);
or U35905 (N_35905,N_32191,N_34689);
xor U35906 (N_35906,N_34808,N_34721);
or U35907 (N_35907,N_33578,N_30421);
nor U35908 (N_35908,N_34388,N_30644);
or U35909 (N_35909,N_31665,N_34331);
nor U35910 (N_35910,N_32139,N_33344);
or U35911 (N_35911,N_30657,N_33109);
nand U35912 (N_35912,N_33981,N_34625);
nor U35913 (N_35913,N_33416,N_32538);
or U35914 (N_35914,N_30569,N_34122);
nor U35915 (N_35915,N_33145,N_33348);
or U35916 (N_35916,N_31085,N_32215);
or U35917 (N_35917,N_31871,N_30686);
xor U35918 (N_35918,N_30737,N_33755);
nand U35919 (N_35919,N_34463,N_34575);
or U35920 (N_35920,N_34755,N_33924);
xor U35921 (N_35921,N_30272,N_31775);
nor U35922 (N_35922,N_34293,N_30213);
and U35923 (N_35923,N_33512,N_33042);
nor U35924 (N_35924,N_32848,N_32906);
and U35925 (N_35925,N_33702,N_32524);
nor U35926 (N_35926,N_34654,N_30117);
or U35927 (N_35927,N_31784,N_30228);
and U35928 (N_35928,N_34577,N_34882);
nand U35929 (N_35929,N_34116,N_33993);
nand U35930 (N_35930,N_32888,N_33975);
nand U35931 (N_35931,N_32402,N_31937);
and U35932 (N_35932,N_33287,N_32062);
and U35933 (N_35933,N_34811,N_33854);
nor U35934 (N_35934,N_32470,N_30648);
nand U35935 (N_35935,N_31780,N_30269);
and U35936 (N_35936,N_30564,N_33016);
xor U35937 (N_35937,N_31888,N_32549);
or U35938 (N_35938,N_34773,N_34484);
nor U35939 (N_35939,N_32041,N_30122);
nand U35940 (N_35940,N_34683,N_34318);
nand U35941 (N_35941,N_30882,N_32603);
and U35942 (N_35942,N_31026,N_31978);
and U35943 (N_35943,N_30186,N_30853);
xnor U35944 (N_35944,N_32800,N_34621);
nand U35945 (N_35945,N_31094,N_30093);
nand U35946 (N_35946,N_34831,N_30866);
and U35947 (N_35947,N_30273,N_31790);
and U35948 (N_35948,N_34244,N_32022);
xnor U35949 (N_35949,N_33285,N_34790);
nor U35950 (N_35950,N_32720,N_31264);
nand U35951 (N_35951,N_32964,N_31757);
nand U35952 (N_35952,N_32131,N_30199);
nand U35953 (N_35953,N_30516,N_30169);
or U35954 (N_35954,N_32064,N_32349);
or U35955 (N_35955,N_33468,N_30471);
nand U35956 (N_35956,N_34991,N_30584);
nand U35957 (N_35957,N_31717,N_32567);
xor U35958 (N_35958,N_30890,N_34661);
or U35959 (N_35959,N_31608,N_33944);
and U35960 (N_35960,N_30763,N_33098);
nand U35961 (N_35961,N_30653,N_33705);
nand U35962 (N_35962,N_32342,N_34715);
xor U35963 (N_35963,N_34502,N_30650);
nand U35964 (N_35964,N_34253,N_33642);
and U35965 (N_35965,N_30046,N_34151);
xnor U35966 (N_35966,N_33205,N_33776);
and U35967 (N_35967,N_31843,N_33001);
nor U35968 (N_35968,N_33332,N_31379);
nor U35969 (N_35969,N_30028,N_31709);
nor U35970 (N_35970,N_30907,N_34555);
nor U35971 (N_35971,N_34765,N_32282);
and U35972 (N_35972,N_34259,N_34997);
nor U35973 (N_35973,N_33588,N_32838);
nand U35974 (N_35974,N_31008,N_30765);
nor U35975 (N_35975,N_30944,N_31500);
xnor U35976 (N_35976,N_30683,N_31525);
or U35977 (N_35977,N_34996,N_32777);
nand U35978 (N_35978,N_33265,N_32874);
nor U35979 (N_35979,N_33442,N_32261);
and U35980 (N_35980,N_31255,N_31561);
xor U35981 (N_35981,N_33813,N_30119);
or U35982 (N_35982,N_31132,N_33187);
nor U35983 (N_35983,N_31731,N_32482);
nand U35984 (N_35984,N_34696,N_34890);
and U35985 (N_35985,N_33283,N_33615);
nand U35986 (N_35986,N_30860,N_33225);
or U35987 (N_35987,N_33229,N_33784);
and U35988 (N_35988,N_32887,N_30242);
or U35989 (N_35989,N_31140,N_34308);
and U35990 (N_35990,N_32255,N_34101);
or U35991 (N_35991,N_31957,N_33335);
xor U35992 (N_35992,N_32748,N_34887);
nor U35993 (N_35993,N_30983,N_31400);
and U35994 (N_35994,N_34910,N_34744);
nand U35995 (N_35995,N_34255,N_33259);
nor U35996 (N_35996,N_31477,N_33920);
nand U35997 (N_35997,N_34422,N_33726);
xor U35998 (N_35998,N_30595,N_33969);
and U35999 (N_35999,N_32317,N_33437);
xnor U36000 (N_36000,N_30056,N_33310);
nand U36001 (N_36001,N_34356,N_34362);
or U36002 (N_36002,N_31256,N_34510);
nor U36003 (N_36003,N_33469,N_32098);
nor U36004 (N_36004,N_33414,N_34148);
or U36005 (N_36005,N_31039,N_31187);
xor U36006 (N_36006,N_31884,N_30701);
nor U36007 (N_36007,N_33890,N_33927);
nand U36008 (N_36008,N_32018,N_34015);
nor U36009 (N_36009,N_33158,N_31905);
nand U36010 (N_36010,N_31557,N_31343);
or U36011 (N_36011,N_34749,N_31661);
or U36012 (N_36012,N_33752,N_31307);
xor U36013 (N_36013,N_30204,N_30735);
and U36014 (N_36014,N_32784,N_32759);
nor U36015 (N_36015,N_31787,N_32439);
and U36016 (N_36016,N_31528,N_33079);
and U36017 (N_36017,N_32537,N_33233);
nor U36018 (N_36018,N_34830,N_30138);
xor U36019 (N_36019,N_31835,N_32187);
xor U36020 (N_36020,N_30210,N_34038);
and U36021 (N_36021,N_34561,N_30912);
nor U36022 (N_36022,N_31555,N_32398);
and U36023 (N_36023,N_31870,N_32412);
and U36024 (N_36024,N_33911,N_33279);
nand U36025 (N_36025,N_33112,N_34194);
nand U36026 (N_36026,N_30698,N_33261);
xor U36027 (N_36027,N_32242,N_30717);
xnor U36028 (N_36028,N_33671,N_34252);
nand U36029 (N_36029,N_31000,N_32158);
or U36030 (N_36030,N_32902,N_31440);
nor U36031 (N_36031,N_32949,N_30035);
xnor U36032 (N_36032,N_31203,N_30144);
and U36033 (N_36033,N_31471,N_33788);
nor U36034 (N_36034,N_32757,N_34081);
nor U36035 (N_36035,N_33594,N_34560);
and U36036 (N_36036,N_31167,N_33979);
nor U36037 (N_36037,N_34418,N_33908);
nor U36038 (N_36038,N_33562,N_31949);
nand U36039 (N_36039,N_30050,N_34757);
nor U36040 (N_36040,N_30741,N_32856);
nor U36041 (N_36041,N_33892,N_33426);
and U36042 (N_36042,N_31131,N_33582);
nand U36043 (N_36043,N_34342,N_31898);
and U36044 (N_36044,N_31642,N_31959);
xnor U36045 (N_36045,N_30489,N_33254);
nor U36046 (N_36046,N_30390,N_33804);
nand U36047 (N_36047,N_33713,N_33459);
or U36048 (N_36048,N_30634,N_30772);
or U36049 (N_36049,N_32265,N_32935);
and U36050 (N_36050,N_34570,N_33891);
and U36051 (N_36051,N_34734,N_34324);
and U36052 (N_36052,N_34487,N_30577);
nand U36053 (N_36053,N_32773,N_31778);
xor U36054 (N_36054,N_34460,N_34738);
or U36055 (N_36055,N_30954,N_34710);
or U36056 (N_36056,N_34748,N_31912);
xor U36057 (N_36057,N_30487,N_34200);
nand U36058 (N_36058,N_30858,N_30456);
and U36059 (N_36059,N_31996,N_34609);
or U36060 (N_36060,N_30554,N_33471);
xnor U36061 (N_36061,N_32659,N_31067);
nand U36062 (N_36062,N_34992,N_30666);
or U36063 (N_36063,N_31329,N_33939);
or U36064 (N_36064,N_33053,N_30808);
nor U36065 (N_36065,N_33880,N_30482);
nand U36066 (N_36066,N_33037,N_31995);
nand U36067 (N_36067,N_33197,N_34618);
nand U36068 (N_36068,N_32230,N_31061);
nor U36069 (N_36069,N_34221,N_34160);
xnor U36070 (N_36070,N_34309,N_32262);
nor U36071 (N_36071,N_31295,N_32953);
nor U36072 (N_36072,N_32755,N_33661);
and U36073 (N_36073,N_34345,N_34569);
and U36074 (N_36074,N_31172,N_33614);
nand U36075 (N_36075,N_31487,N_30702);
xor U36076 (N_36076,N_34482,N_32907);
nand U36077 (N_36077,N_31431,N_31933);
xnor U36078 (N_36078,N_30507,N_34147);
or U36079 (N_36079,N_32697,N_30753);
nand U36080 (N_36080,N_32920,N_31492);
nand U36081 (N_36081,N_32259,N_33419);
or U36082 (N_36082,N_31985,N_33282);
or U36083 (N_36083,N_34742,N_34327);
or U36084 (N_36084,N_30901,N_33901);
or U36085 (N_36085,N_33808,N_31193);
nand U36086 (N_36086,N_33557,N_31650);
nor U36087 (N_36087,N_32127,N_30847);
nor U36088 (N_36088,N_31009,N_31952);
xor U36089 (N_36089,N_31263,N_30722);
or U36090 (N_36090,N_30127,N_31423);
xnor U36091 (N_36091,N_34770,N_30645);
and U36092 (N_36092,N_30352,N_31997);
and U36093 (N_36093,N_31943,N_34466);
nor U36094 (N_36094,N_31113,N_31089);
and U36095 (N_36095,N_33380,N_31035);
nor U36096 (N_36096,N_33654,N_31864);
or U36097 (N_36097,N_30347,N_32000);
xnor U36098 (N_36098,N_32660,N_32726);
nor U36099 (N_36099,N_31038,N_33102);
nor U36100 (N_36100,N_32909,N_34404);
nor U36101 (N_36101,N_33625,N_32562);
xnor U36102 (N_36102,N_31756,N_34198);
or U36103 (N_36103,N_34084,N_33592);
or U36104 (N_36104,N_30622,N_30777);
and U36105 (N_36105,N_31302,N_30274);
and U36106 (N_36106,N_32732,N_32708);
and U36107 (N_36107,N_34192,N_33836);
xor U36108 (N_36108,N_30439,N_32883);
xor U36109 (N_36109,N_33617,N_31613);
nand U36110 (N_36110,N_31641,N_32360);
nand U36111 (N_36111,N_30885,N_34010);
nor U36112 (N_36112,N_33942,N_32841);
or U36113 (N_36113,N_34766,N_33220);
or U36114 (N_36114,N_32648,N_34668);
nor U36115 (N_36115,N_33510,N_30836);
or U36116 (N_36116,N_32791,N_33695);
nor U36117 (N_36117,N_32678,N_32650);
xnor U36118 (N_36118,N_30264,N_33548);
or U36119 (N_36119,N_30719,N_30884);
nor U36120 (N_36120,N_32469,N_32997);
or U36121 (N_36121,N_33114,N_33212);
nand U36122 (N_36122,N_32068,N_34085);
and U36123 (N_36123,N_30292,N_32637);
and U36124 (N_36124,N_31953,N_32169);
nand U36125 (N_36125,N_30206,N_34326);
and U36126 (N_36126,N_32552,N_33050);
xor U36127 (N_36127,N_34592,N_31200);
xnor U36128 (N_36128,N_33988,N_31584);
nor U36129 (N_36129,N_34312,N_32640);
or U36130 (N_36130,N_30070,N_30214);
and U36131 (N_36131,N_34367,N_32652);
nand U36132 (N_36132,N_34895,N_33051);
and U36133 (N_36133,N_34705,N_34006);
nand U36134 (N_36134,N_32970,N_30052);
xnor U36135 (N_36135,N_31346,N_34578);
and U36136 (N_36136,N_33148,N_34251);
xor U36137 (N_36137,N_33842,N_30991);
xor U36138 (N_36138,N_34166,N_34965);
and U36139 (N_36139,N_34917,N_32763);
nand U36140 (N_36140,N_32316,N_30406);
or U36141 (N_36141,N_34245,N_30400);
nand U36142 (N_36142,N_30992,N_31338);
or U36143 (N_36143,N_34352,N_31582);
and U36144 (N_36144,N_32142,N_32675);
xnor U36145 (N_36145,N_33231,N_34407);
and U36146 (N_36146,N_30929,N_31208);
nor U36147 (N_36147,N_33570,N_33556);
and U36148 (N_36148,N_31593,N_31605);
and U36149 (N_36149,N_33787,N_31596);
and U36150 (N_36150,N_34435,N_31982);
nor U36151 (N_36151,N_31906,N_30057);
or U36152 (N_36152,N_33431,N_32808);
or U36153 (N_36153,N_32608,N_30321);
nor U36154 (N_36154,N_31435,N_32734);
or U36155 (N_36155,N_32779,N_34513);
nand U36156 (N_36156,N_33099,N_31084);
or U36157 (N_36157,N_31291,N_30247);
and U36158 (N_36158,N_34225,N_33477);
and U36159 (N_36159,N_30834,N_32928);
nand U36160 (N_36160,N_33031,N_34450);
or U36161 (N_36161,N_33657,N_33746);
nor U36162 (N_36162,N_30015,N_32028);
xnor U36163 (N_36163,N_33541,N_32731);
and U36164 (N_36164,N_32743,N_34681);
xnor U36165 (N_36165,N_31286,N_32923);
nor U36166 (N_36166,N_33358,N_30342);
and U36167 (N_36167,N_30198,N_32121);
nand U36168 (N_36168,N_31178,N_30211);
nor U36169 (N_36169,N_34798,N_32453);
nor U36170 (N_36170,N_34098,N_34622);
nor U36171 (N_36171,N_32555,N_31331);
and U36172 (N_36172,N_34137,N_31230);
and U36173 (N_36173,N_32416,N_31288);
nand U36174 (N_36174,N_31701,N_32389);
and U36175 (N_36175,N_32108,N_33783);
nand U36176 (N_36176,N_33721,N_34421);
or U36177 (N_36177,N_30568,N_30451);
or U36178 (N_36178,N_33843,N_34005);
nand U36179 (N_36179,N_32397,N_33547);
nand U36180 (N_36180,N_34932,N_33729);
and U36181 (N_36181,N_32425,N_34079);
xnor U36182 (N_36182,N_32933,N_32162);
xor U36183 (N_36183,N_33727,N_32619);
nand U36184 (N_36184,N_31070,N_30367);
nor U36185 (N_36185,N_34863,N_32186);
nand U36186 (N_36186,N_30606,N_31702);
and U36187 (N_36187,N_30453,N_33827);
nand U36188 (N_36188,N_32074,N_30843);
nor U36189 (N_36189,N_34907,N_30973);
xnor U36190 (N_36190,N_31234,N_32446);
or U36191 (N_36191,N_30303,N_31106);
and U36192 (N_36192,N_33675,N_34492);
and U36193 (N_36193,N_34195,N_31852);
or U36194 (N_36194,N_33420,N_33291);
xor U36195 (N_36195,N_34341,N_30518);
nand U36196 (N_36196,N_31565,N_30512);
or U36197 (N_36197,N_30003,N_30286);
or U36198 (N_36198,N_32655,N_31454);
and U36199 (N_36199,N_30880,N_34962);
and U36200 (N_36200,N_31358,N_34824);
and U36201 (N_36201,N_31515,N_30257);
nand U36202 (N_36202,N_32628,N_34222);
and U36203 (N_36203,N_31617,N_34185);
nor U36204 (N_36204,N_32869,N_30571);
and U36205 (N_36205,N_33492,N_34153);
xnor U36206 (N_36206,N_32715,N_34257);
or U36207 (N_36207,N_30431,N_30781);
nor U36208 (N_36208,N_34174,N_31093);
nand U36209 (N_36209,N_30673,N_34102);
and U36210 (N_36210,N_30099,N_31976);
and U36211 (N_36211,N_34985,N_31493);
nand U36212 (N_36212,N_33385,N_33153);
nand U36213 (N_36213,N_30047,N_34803);
and U36214 (N_36214,N_32125,N_33734);
or U36215 (N_36215,N_33341,N_30283);
nor U36216 (N_36216,N_31833,N_32424);
and U36217 (N_36217,N_30962,N_32461);
and U36218 (N_36218,N_34368,N_31614);
xnor U36219 (N_36219,N_32188,N_32927);
and U36220 (N_36220,N_33424,N_34550);
and U36221 (N_36221,N_31849,N_31430);
nor U36222 (N_36222,N_34468,N_33303);
or U36223 (N_36223,N_33933,N_32407);
or U36224 (N_36224,N_31573,N_32171);
nand U36225 (N_36225,N_32030,N_32781);
and U36226 (N_36226,N_33271,N_31653);
nand U36227 (N_36227,N_33543,N_33011);
xor U36228 (N_36228,N_32298,N_33766);
and U36229 (N_36229,N_31522,N_34699);
and U36230 (N_36230,N_34877,N_31828);
and U36231 (N_36231,N_31872,N_32153);
nor U36232 (N_36232,N_31855,N_32027);
nand U36233 (N_36233,N_30455,N_31145);
xor U36234 (N_36234,N_34595,N_32788);
or U36235 (N_36235,N_31202,N_31001);
nand U36236 (N_36236,N_34003,N_30867);
or U36237 (N_36237,N_31041,N_30141);
or U36238 (N_36238,N_31387,N_31550);
and U36239 (N_36239,N_30128,N_33930);
and U36240 (N_36240,N_31742,N_31393);
xor U36241 (N_36241,N_31553,N_31164);
xnor U36242 (N_36242,N_32165,N_33033);
and U36243 (N_36243,N_31275,N_34472);
nand U36244 (N_36244,N_32824,N_32940);
nor U36245 (N_36245,N_33085,N_30133);
or U36246 (N_36246,N_34925,N_33359);
or U36247 (N_36247,N_33245,N_34551);
xnor U36248 (N_36248,N_34657,N_31057);
or U36249 (N_36249,N_30693,N_32690);
xnor U36250 (N_36250,N_34760,N_34774);
and U36251 (N_36251,N_32381,N_33248);
nand U36252 (N_36252,N_30955,N_33059);
nor U36253 (N_36253,N_33387,N_31659);
and U36254 (N_36254,N_30445,N_33878);
and U36255 (N_36255,N_30069,N_32208);
nor U36256 (N_36256,N_31426,N_31566);
xnor U36257 (N_36257,N_31882,N_31899);
or U36258 (N_36258,N_31082,N_33141);
xnor U36259 (N_36259,N_33488,N_34566);
or U36260 (N_36260,N_31998,N_30480);
nor U36261 (N_36261,N_32404,N_30415);
xor U36262 (N_36262,N_32626,N_31713);
and U36263 (N_36263,N_30810,N_32535);
or U36264 (N_36264,N_32092,N_30483);
and U36265 (N_36265,N_34781,N_33009);
nand U36266 (N_36266,N_34224,N_30125);
nand U36267 (N_36267,N_33460,N_34603);
nor U36268 (N_36268,N_30801,N_31893);
xor U36269 (N_36269,N_30124,N_33662);
nor U36270 (N_36270,N_30111,N_30354);
xor U36271 (N_36271,N_32596,N_31229);
nand U36272 (N_36272,N_31148,N_31639);
and U36273 (N_36273,N_34216,N_31935);
or U36274 (N_36274,N_33991,N_33907);
nand U36275 (N_36275,N_32712,N_34676);
nor U36276 (N_36276,N_30066,N_33106);
nand U36277 (N_36277,N_32736,N_31861);
nor U36278 (N_36278,N_34287,N_34520);
nand U36279 (N_36279,N_32228,N_30524);
and U36280 (N_36280,N_33201,N_31046);
nor U36281 (N_36281,N_32503,N_32870);
nand U36282 (N_36282,N_33338,N_34697);
or U36283 (N_36283,N_31319,N_33336);
or U36284 (N_36284,N_31068,N_31049);
xnor U36285 (N_36285,N_33138,N_32471);
nor U36286 (N_36286,N_33479,N_32112);
or U36287 (N_36287,N_34861,N_34880);
nand U36288 (N_36288,N_31502,N_33852);
or U36289 (N_36289,N_31244,N_32683);
nand U36290 (N_36290,N_32284,N_34156);
or U36291 (N_36291,N_31272,N_30470);
xor U36292 (N_36292,N_32835,N_31754);
xnor U36293 (N_36293,N_32350,N_32114);
or U36294 (N_36294,N_33278,N_32332);
xor U36295 (N_36295,N_33984,N_34157);
xor U36296 (N_36296,N_30176,N_34105);
nand U36297 (N_36297,N_31250,N_32240);
and U36298 (N_36298,N_30596,N_31885);
nor U36299 (N_36299,N_31253,N_31330);
nand U36300 (N_36300,N_31428,N_33698);
xor U36301 (N_36301,N_31853,N_33270);
nor U36302 (N_36302,N_32136,N_31417);
or U36303 (N_36303,N_32713,N_34857);
or U36304 (N_36304,N_33884,N_33400);
or U36305 (N_36305,N_30276,N_33632);
or U36306 (N_36306,N_31278,N_32722);
or U36307 (N_36307,N_33177,N_32409);
or U36308 (N_36308,N_30598,N_32632);
and U36309 (N_36309,N_31716,N_30243);
xnor U36310 (N_36310,N_31408,N_32646);
or U36311 (N_36311,N_30197,N_30788);
or U36312 (N_36312,N_32217,N_34812);
nand U36313 (N_36313,N_34647,N_30857);
or U36314 (N_36314,N_30829,N_32972);
or U36315 (N_36315,N_31072,N_30618);
nand U36316 (N_36316,N_33113,N_30635);
nor U36317 (N_36317,N_32154,N_34797);
or U36318 (N_36318,N_34115,N_30585);
nor U36319 (N_36319,N_31249,N_31804);
nand U36320 (N_36320,N_30475,N_33932);
and U36321 (N_36321,N_34731,N_34941);
xnor U36322 (N_36322,N_32106,N_34619);
nor U36323 (N_36323,N_32896,N_31305);
nor U36324 (N_36324,N_30610,N_34249);
nand U36325 (N_36325,N_31826,N_34103);
or U36326 (N_36326,N_32951,N_34794);
xor U36327 (N_36327,N_34776,N_32442);
nor U36328 (N_36328,N_34136,N_33004);
nor U36329 (N_36329,N_34971,N_34772);
xor U36330 (N_36330,N_31940,N_32193);
or U36331 (N_36331,N_30656,N_30009);
nor U36332 (N_36332,N_34919,N_30534);
xor U36333 (N_36333,N_31073,N_30979);
or U36334 (N_36334,N_30136,N_34159);
nand U36335 (N_36335,N_32338,N_32075);
or U36336 (N_36336,N_33753,N_30915);
and U36337 (N_36337,N_31339,N_34835);
and U36338 (N_36338,N_34497,N_31351);
and U36339 (N_36339,N_30041,N_32532);
nand U36340 (N_36340,N_34231,N_33971);
nand U36341 (N_36341,N_33204,N_32406);
and U36342 (N_36342,N_32476,N_33845);
or U36343 (N_36343,N_34471,N_34814);
xnor U36344 (N_36344,N_30778,N_32483);
xor U36345 (N_36345,N_32546,N_30333);
xor U36346 (N_36346,N_34055,N_31710);
or U36347 (N_36347,N_31889,N_32636);
or U36348 (N_36348,N_31120,N_33515);
nand U36349 (N_36349,N_32494,N_32313);
and U36350 (N_36350,N_30716,N_31452);
nor U36351 (N_36351,N_31436,N_32644);
or U36352 (N_36352,N_32950,N_30166);
and U36353 (N_36353,N_30876,N_31441);
or U36354 (N_36354,N_34921,N_30355);
nor U36355 (N_36355,N_34132,N_32674);
and U36356 (N_36356,N_30311,N_32056);
nor U36357 (N_36357,N_31136,N_31173);
xnor U36358 (N_36358,N_34826,N_33345);
nand U36359 (N_36359,N_34620,N_33343);
and U36360 (N_36360,N_32517,N_32716);
and U36361 (N_36361,N_31589,N_30597);
nor U36362 (N_36362,N_32765,N_33065);
xnor U36363 (N_36363,N_32050,N_34692);
or U36364 (N_36364,N_31992,N_31602);
nor U36365 (N_36365,N_30682,N_34672);
or U36366 (N_36366,N_32864,N_34433);
and U36367 (N_36367,N_31158,N_33733);
xnor U36368 (N_36368,N_34453,N_34881);
and U36369 (N_36369,N_34125,N_31448);
or U36370 (N_36370,N_32581,N_30787);
nand U36371 (N_36371,N_33526,N_32698);
xor U36372 (N_36372,N_30956,N_34020);
or U36373 (N_36373,N_30646,N_34628);
nor U36374 (N_36374,N_30659,N_33239);
nor U36375 (N_36375,N_34413,N_31322);
nor U36376 (N_36376,N_32614,N_31228);
nor U36377 (N_36377,N_32967,N_34451);
and U36378 (N_36378,N_31520,N_32995);
nor U36379 (N_36379,N_32029,N_33227);
and U36380 (N_36380,N_31194,N_33390);
xor U36381 (N_36381,N_34833,N_34196);
and U36382 (N_36382,N_32088,N_31186);
nand U36383 (N_36383,N_30306,N_33628);
xnor U36384 (N_36384,N_30529,N_31883);
and U36385 (N_36385,N_30059,N_30464);
or U36386 (N_36386,N_31285,N_30576);
xor U36387 (N_36387,N_33779,N_33764);
or U36388 (N_36388,N_32202,N_33395);
or U36389 (N_36389,N_34506,N_34583);
xnor U36390 (N_36390,N_31895,N_34543);
xnor U36391 (N_36391,N_30187,N_32681);
and U36392 (N_36392,N_32610,N_31386);
nand U36393 (N_36393,N_31645,N_31881);
xnor U36394 (N_36394,N_31524,N_31901);
and U36395 (N_36395,N_30540,N_32819);
or U36396 (N_36396,N_30649,N_33505);
or U36397 (N_36397,N_34854,N_30370);
xor U36398 (N_36398,N_34660,N_30389);
xnor U36399 (N_36399,N_33744,N_31369);
xnor U36400 (N_36400,N_30163,N_34219);
xnor U36401 (N_36401,N_33840,N_30132);
or U36402 (N_36402,N_32862,N_31433);
or U36403 (N_36403,N_31903,N_33593);
nor U36404 (N_36404,N_30825,N_32477);
nor U36405 (N_36405,N_31730,N_31691);
or U36406 (N_36406,N_32233,N_32832);
or U36407 (N_36407,N_31629,N_33525);
nand U36408 (N_36408,N_30502,N_31378);
xnor U36409 (N_36409,N_33800,N_32730);
xor U36410 (N_36410,N_34355,N_30452);
and U36411 (N_36411,N_33256,N_34386);
xor U36412 (N_36412,N_32980,N_33611);
nand U36413 (N_36413,N_33798,N_32452);
nand U36414 (N_36414,N_30346,N_31622);
or U36415 (N_36415,N_31481,N_34092);
nor U36416 (N_36416,N_33596,N_32871);
nand U36417 (N_36417,N_30727,N_33013);
nand U36418 (N_36418,N_31621,N_31558);
or U36419 (N_36419,N_34993,N_33506);
nor U36420 (N_36420,N_33347,N_31546);
and U36421 (N_36421,N_34548,N_30852);
xor U36422 (N_36422,N_33834,N_33814);
nor U36423 (N_36423,N_34562,N_34752);
xor U36424 (N_36424,N_32456,N_33810);
and U36425 (N_36425,N_31206,N_30291);
nand U36426 (N_36426,N_34980,N_32580);
xnor U36427 (N_36427,N_34490,N_33467);
nor U36428 (N_36428,N_32331,N_31461);
nand U36429 (N_36429,N_34295,N_30519);
and U36430 (N_36430,N_33054,N_34248);
xor U36431 (N_36431,N_31510,N_34964);
and U36432 (N_36432,N_34817,N_31823);
xor U36433 (N_36433,N_33238,N_30289);
and U36434 (N_36434,N_34142,N_34759);
nand U36435 (N_36435,N_34376,N_30215);
nor U36436 (N_36436,N_34041,N_34546);
or U36437 (N_36437,N_34024,N_30832);
or U36438 (N_36438,N_32091,N_34186);
xor U36439 (N_36439,N_32623,N_31023);
or U36440 (N_36440,N_33132,N_30203);
or U36441 (N_36441,N_31040,N_31146);
or U36442 (N_36442,N_32544,N_34280);
nand U36443 (N_36443,N_34671,N_32105);
nand U36444 (N_36444,N_31836,N_32299);
xnor U36445 (N_36445,N_33534,N_33905);
nor U36446 (N_36446,N_32058,N_30495);
or U36447 (N_36447,N_30864,N_30221);
nand U36448 (N_36448,N_30710,N_30877);
and U36449 (N_36449,N_31226,N_32982);
xor U36450 (N_36450,N_31848,N_32143);
nor U36451 (N_36451,N_33235,N_32365);
and U36452 (N_36452,N_30974,N_34037);
or U36453 (N_36453,N_34215,N_33313);
or U36454 (N_36454,N_30092,N_32811);
nand U36455 (N_36455,N_34637,N_30551);
and U36456 (N_36456,N_33449,N_30893);
and U36457 (N_36457,N_31141,N_30523);
and U36458 (N_36458,N_31344,N_30377);
or U36459 (N_36459,N_34369,N_32291);
nand U36460 (N_36460,N_32377,N_30158);
xor U36461 (N_36461,N_30010,N_30543);
nand U36462 (N_36462,N_33980,N_32865);
and U36463 (N_36463,N_34645,N_32172);
nor U36464 (N_36464,N_31469,N_30183);
or U36465 (N_36465,N_30001,N_32806);
nand U36466 (N_36466,N_34986,N_33292);
nor U36467 (N_36467,N_31372,N_30371);
nand U36468 (N_36468,N_32335,N_32305);
nand U36469 (N_36469,N_30674,N_30695);
nor U36470 (N_36470,N_30842,N_32109);
nand U36471 (N_36471,N_33742,N_33535);
and U36472 (N_36472,N_31366,N_30304);
and U36473 (N_36473,N_32275,N_30780);
xor U36474 (N_36474,N_32199,N_31359);
nand U36475 (N_36475,N_31615,N_31012);
or U36476 (N_36476,N_31532,N_33575);
xor U36477 (N_36477,N_34296,N_32118);
and U36478 (N_36478,N_30921,N_33530);
or U36479 (N_36479,N_31277,N_34118);
nor U36480 (N_36480,N_34594,N_30961);
xnor U36481 (N_36481,N_33369,N_31581);
nor U36482 (N_36482,N_31209,N_30299);
or U36483 (N_36483,N_31219,N_31723);
and U36484 (N_36484,N_30581,N_31098);
xnor U36485 (N_36485,N_30279,N_34860);
nand U36486 (N_36486,N_32040,N_30593);
or U36487 (N_36487,N_32578,N_33306);
xnor U36488 (N_36488,N_32937,N_34912);
or U36489 (N_36489,N_30496,N_32015);
and U36490 (N_36490,N_32595,N_32917);
nor U36491 (N_36491,N_31772,N_33244);
nand U36492 (N_36492,N_31483,N_31443);
nand U36493 (N_36493,N_30582,N_31238);
xnor U36494 (N_36494,N_33559,N_30774);
or U36495 (N_36495,N_31939,N_34518);
and U36496 (N_36496,N_32837,N_31963);
and U36497 (N_36497,N_31863,N_33047);
or U36498 (N_36498,N_33268,N_34128);
xnor U36499 (N_36499,N_32577,N_34403);
nand U36500 (N_36500,N_30900,N_33164);
nor U36501 (N_36501,N_31102,N_33308);
xnor U36502 (N_36502,N_33867,N_30796);
or U36503 (N_36503,N_33317,N_30336);
and U36504 (N_36504,N_30926,N_34053);
nor U36505 (N_36505,N_31722,N_34728);
nand U36506 (N_36506,N_34062,N_32621);
and U36507 (N_36507,N_33600,N_32981);
xor U36508 (N_36508,N_33234,N_30869);
nor U36509 (N_36509,N_32175,N_31989);
nor U36510 (N_36510,N_32079,N_34785);
or U36511 (N_36511,N_32880,N_30442);
or U36512 (N_36512,N_34899,N_30914);
nor U36513 (N_36513,N_32234,N_32236);
xnor U36514 (N_36514,N_31806,N_31827);
xnor U36515 (N_36515,N_32989,N_32124);
or U36516 (N_36516,N_32422,N_32717);
and U36517 (N_36517,N_31495,N_30937);
xor U36518 (N_36518,N_33005,N_33321);
xnor U36519 (N_36519,N_30373,N_30619);
xor U36520 (N_36520,N_32005,N_31547);
and U36521 (N_36521,N_30712,N_31005);
nand U36522 (N_36522,N_32324,N_33081);
and U36523 (N_36523,N_31814,N_34792);
and U36524 (N_36524,N_31682,N_31956);
or U36525 (N_36525,N_32991,N_34761);
and U36526 (N_36526,N_30402,N_34313);
nand U36527 (N_36527,N_30626,N_30636);
nand U36528 (N_36528,N_34970,N_32238);
or U36529 (N_36529,N_30325,N_32182);
nand U36530 (N_36530,N_33230,N_32498);
or U36531 (N_36531,N_34431,N_31354);
xnor U36532 (N_36532,N_30388,N_31950);
xor U36533 (N_36533,N_31058,N_33088);
or U36534 (N_36534,N_31793,N_32616);
and U36535 (N_36535,N_30671,N_34420);
and U36536 (N_36536,N_32479,N_33651);
nor U36537 (N_36537,N_30023,N_30168);
xnor U36538 (N_36538,N_30427,N_33349);
or U36539 (N_36539,N_32553,N_33966);
and U36540 (N_36540,N_32447,N_33875);
nand U36541 (N_36541,N_33803,N_34885);
nand U36542 (N_36542,N_34646,N_33301);
nor U36543 (N_36543,N_32312,N_34458);
or U36544 (N_36544,N_30839,N_32003);
nor U36545 (N_36545,N_30824,N_33738);
and U36546 (N_36546,N_31267,N_32220);
xor U36547 (N_36547,N_32246,N_33855);
nand U36548 (N_36548,N_33015,N_31318);
and U36549 (N_36549,N_30323,N_32592);
or U36550 (N_36550,N_34239,N_32515);
or U36551 (N_36551,N_30513,N_34076);
xnor U36552 (N_36552,N_33111,N_34563);
or U36553 (N_36553,N_30463,N_31505);
or U36554 (N_36554,N_30802,N_30454);
or U36555 (N_36555,N_32810,N_34547);
and U36556 (N_36556,N_33758,N_30713);
xnor U36557 (N_36557,N_32006,N_30967);
xnor U36558 (N_36558,N_33532,N_33756);
or U36559 (N_36559,N_31640,N_33189);
nor U36560 (N_36560,N_30939,N_30726);
xor U36561 (N_36561,N_34884,N_30488);
or U36562 (N_36562,N_34730,N_33565);
nand U36563 (N_36563,N_33174,N_31398);
or U36564 (N_36564,N_31446,N_34544);
nand U36565 (N_36565,N_31712,N_32992);
xor U36566 (N_36566,N_34049,N_32624);
nor U36567 (N_36567,N_30021,N_30256);
nand U36568 (N_36568,N_34727,N_30738);
xnor U36569 (N_36569,N_30691,N_32830);
xnor U36570 (N_36570,N_33215,N_33045);
and U36571 (N_36571,N_31016,N_33195);
nor U36572 (N_36572,N_32382,N_33226);
or U36573 (N_36573,N_32164,N_33960);
and U36574 (N_36574,N_30942,N_30692);
and U36575 (N_36575,N_33775,N_32201);
xor U36576 (N_36576,N_34615,N_31470);
or U36577 (N_36577,N_34678,N_32113);
xnor U36578 (N_36578,N_32480,N_30561);
and U36579 (N_36579,N_34658,N_34077);
xnor U36580 (N_36580,N_34649,N_31118);
and U36581 (N_36581,N_34931,N_33127);
nor U36582 (N_36582,N_32352,N_32820);
xnor U36583 (N_36583,N_30736,N_30437);
or U36584 (N_36584,N_34371,N_33972);
and U36585 (N_36585,N_34455,N_33622);
xnor U36586 (N_36586,N_31242,N_31412);
nand U36587 (N_36587,N_32714,N_34491);
nand U36588 (N_36588,N_30287,N_30799);
xor U36589 (N_36589,N_31695,N_31336);
nand U36590 (N_36590,N_33028,N_31744);
xor U36591 (N_36591,N_33918,N_31991);
nand U36592 (N_36592,N_34338,N_32214);
or U36593 (N_36593,N_31103,N_34277);
and U36594 (N_36594,N_34940,N_30733);
xnor U36595 (N_36595,N_33871,N_32943);
nor U36596 (N_36596,N_34208,N_32330);
nor U36597 (N_36597,N_31498,N_33223);
nand U36598 (N_36598,N_32527,N_32676);
nand U36599 (N_36599,N_34130,N_30906);
nand U36600 (N_36600,N_33780,N_30770);
and U36601 (N_36601,N_31896,N_30806);
nand U36602 (N_36602,N_31247,N_32513);
nor U36603 (N_36603,N_31759,N_31878);
xnor U36604 (N_36604,N_31365,N_34264);
xnor U36605 (N_36605,N_31456,N_34104);
nor U36606 (N_36606,N_32213,N_32044);
xnor U36607 (N_36607,N_32123,N_34365);
nor U36608 (N_36608,N_34307,N_34306);
and U36609 (N_36609,N_30664,N_33954);
nand U36610 (N_36610,N_32975,N_34149);
and U36611 (N_36611,N_31262,N_34182);
xnor U36612 (N_36612,N_33294,N_31548);
nor U36613 (N_36613,N_33736,N_30459);
or U36614 (N_36614,N_30590,N_33922);
nor U36615 (N_36615,N_30762,N_34276);
nor U36616 (N_36616,N_32686,N_33115);
and U36617 (N_36617,N_33462,N_33701);
and U36618 (N_36618,N_30443,N_31462);
xnor U36619 (N_36619,N_33709,N_32420);
xnor U36620 (N_36620,N_31932,N_32219);
or U36621 (N_36621,N_31450,N_30332);
nand U36622 (N_36622,N_31252,N_33374);
nand U36623 (N_36623,N_34841,N_32274);
or U36624 (N_36624,N_30647,N_34425);
or U36625 (N_36625,N_31002,N_32994);
nand U36626 (N_36626,N_34746,N_33342);
xnor U36627 (N_36627,N_34454,N_31183);
nor U36628 (N_36628,N_30037,N_34743);
xor U36629 (N_36629,N_31914,N_30315);
nor U36630 (N_36630,N_30535,N_31687);
nand U36631 (N_36631,N_33415,N_31327);
or U36632 (N_36632,N_31473,N_31748);
nand U36633 (N_36633,N_31970,N_34250);
nor U36634 (N_36634,N_34786,N_34180);
and U36635 (N_36635,N_33816,N_30148);
nand U36636 (N_36636,N_32988,N_31960);
nor U36637 (N_36637,N_30335,N_33371);
nor U36638 (N_36638,N_34888,N_31192);
xnor U36639 (N_36639,N_31501,N_31750);
nand U36640 (N_36640,N_32363,N_30526);
xnor U36641 (N_36641,N_30804,N_32166);
xnor U36642 (N_36642,N_34674,N_34767);
or U36643 (N_36643,N_32473,N_34698);
nand U36644 (N_36644,N_31151,N_30687);
nand U36645 (N_36645,N_32222,N_34567);
nor U36646 (N_36646,N_33357,N_33551);
and U36647 (N_36647,N_33110,N_33550);
nor U36648 (N_36648,N_34778,N_32725);
nand U36649 (N_36649,N_33829,N_32729);
xor U36650 (N_36650,N_30968,N_32055);
nand U36651 (N_36651,N_33206,N_30607);
xnor U36652 (N_36652,N_32542,N_32339);
or U36653 (N_36653,N_30002,N_32803);
and U36654 (N_36654,N_34642,N_34395);
or U36655 (N_36655,N_34093,N_33678);
xor U36656 (N_36656,N_30969,N_33255);
and U36657 (N_36657,N_34189,N_31507);
nor U36658 (N_36658,N_33276,N_34706);
nand U36659 (N_36659,N_33432,N_31097);
nor U36660 (N_36660,N_34154,N_30201);
or U36661 (N_36661,N_31225,N_32566);
xnor U36662 (N_36662,N_33945,N_30345);
nand U36663 (N_36663,N_31171,N_32813);
nor U36664 (N_36664,N_32688,N_33458);
xnor U36665 (N_36665,N_31816,N_34479);
and U36666 (N_36666,N_31007,N_32918);
xor U36667 (N_36667,N_30174,N_31459);
nand U36668 (N_36668,N_30392,N_30193);
xnor U36669 (N_36669,N_32574,N_34266);
nand U36670 (N_36670,N_33455,N_34126);
or U36671 (N_36671,N_33214,N_33386);
nand U36672 (N_36672,N_32986,N_30349);
nor U36673 (N_36673,N_30580,N_30458);
nor U36674 (N_36674,N_33170,N_33331);
nand U36675 (N_36675,N_32138,N_31223);
and U36676 (N_36676,N_32599,N_34827);
nor U36677 (N_36677,N_32173,N_34829);
nand U36678 (N_36678,N_32543,N_30932);
nand U36679 (N_36679,N_33655,N_31074);
xnor U36680 (N_36680,N_30152,N_32017);
nand U36681 (N_36681,N_33411,N_30775);
and U36682 (N_36682,N_33940,N_32846);
and U36683 (N_36683,N_34704,N_32337);
and U36684 (N_36684,N_34004,N_31807);
nor U36685 (N_36685,N_32682,N_33865);
nand U36686 (N_36686,N_30748,N_30887);
and U36687 (N_36687,N_34039,N_32264);
nor U36688 (N_36688,N_30999,N_31587);
xor U36689 (N_36689,N_31770,N_34610);
nor U36690 (N_36690,N_30996,N_33266);
nor U36691 (N_36691,N_34948,N_30173);
or U36692 (N_36692,N_33160,N_34078);
and U36693 (N_36693,N_34599,N_32052);
nand U36694 (N_36694,N_30833,N_30501);
and U36695 (N_36695,N_30899,N_34508);
xor U36696 (N_36696,N_30977,N_33717);
and U36697 (N_36697,N_32329,N_31134);
xnor U36698 (N_36698,N_31755,N_34133);
nand U36699 (N_36699,N_33074,N_32554);
xor U36700 (N_36700,N_32664,N_31590);
xnor U36701 (N_36701,N_32443,N_32776);
and U36702 (N_36702,N_30357,N_32740);
xnor U36703 (N_36703,N_30997,N_30940);
or U36704 (N_36704,N_33976,N_31298);
and U36705 (N_36705,N_34667,N_31115);
or U36706 (N_36706,N_34828,N_30761);
nor U36707 (N_36707,N_30369,N_32448);
or U36708 (N_36708,N_32344,N_34143);
and U36709 (N_36709,N_31514,N_34865);
and U36710 (N_36710,N_30469,N_33683);
xnor U36711 (N_36711,N_34337,N_34908);
nor U36712 (N_36712,N_33968,N_34535);
and U36713 (N_36713,N_31894,N_31815);
or U36714 (N_36714,N_32241,N_33202);
nand U36715 (N_36715,N_33049,N_34274);
xor U36716 (N_36716,N_33916,N_30620);
xor U36717 (N_36717,N_33060,N_33413);
or U36718 (N_36718,N_30709,N_33435);
or U36719 (N_36719,N_32860,N_32545);
and U36720 (N_36720,N_34923,N_33383);
and U36721 (N_36721,N_33992,N_32286);
and U36722 (N_36722,N_34867,N_31334);
nand U36723 (N_36723,N_30393,N_32481);
xnor U36724 (N_36724,N_32384,N_34124);
xnor U36725 (N_36725,N_32444,N_30208);
xnor U36726 (N_36726,N_33365,N_31188);
or U36727 (N_36727,N_31785,N_32700);
and U36728 (N_36728,N_32585,N_33791);
or U36729 (N_36729,N_32204,N_31157);
nor U36730 (N_36730,N_34323,N_30891);
nand U36731 (N_36731,N_31675,N_33826);
nand U36732 (N_36732,N_33269,N_31037);
and U36733 (N_36733,N_30145,N_33409);
xor U36734 (N_36734,N_34305,N_31773);
nor U36735 (N_36735,N_34852,N_33305);
nand U36736 (N_36736,N_33598,N_34793);
or U36737 (N_36737,N_33533,N_32958);
and U36738 (N_36738,N_33589,N_34254);
nor U36739 (N_36739,N_33687,N_30861);
and U36740 (N_36740,N_32807,N_30933);
nor U36741 (N_36741,N_30522,N_32804);
nor U36742 (N_36742,N_31993,N_31405);
nor U36743 (N_36743,N_30871,N_34247);
or U36744 (N_36744,N_32319,N_33366);
or U36745 (N_36745,N_30397,N_30960);
and U36746 (N_36746,N_30072,N_32601);
or U36747 (N_36747,N_33879,N_34446);
nor U36748 (N_36748,N_33773,N_32952);
nand U36749 (N_36749,N_32586,N_32885);
or U36750 (N_36750,N_34900,N_33430);
or U36751 (N_36751,N_32168,N_34849);
nand U36752 (N_36752,N_33973,N_30819);
and U36753 (N_36753,N_31052,N_32897);
nand U36754 (N_36754,N_31078,N_30556);
nor U36755 (N_36755,N_32067,N_30018);
nor U36756 (N_36756,N_34939,N_34842);
and U36757 (N_36757,N_32046,N_31783);
or U36758 (N_36758,N_30875,N_30759);
nand U36759 (N_36759,N_34025,N_34871);
and U36760 (N_36760,N_32370,N_33728);
nor U36761 (N_36761,N_31535,N_33509);
and U36762 (N_36762,N_32849,N_34059);
or U36763 (N_36763,N_30938,N_34360);
nor U36764 (N_36764,N_30728,N_33346);
nor U36765 (N_36765,N_31375,N_32126);
or U36766 (N_36766,N_32959,N_34162);
nor U36767 (N_36767,N_32271,N_33441);
nor U36768 (N_36768,N_31453,N_32392);
nand U36769 (N_36769,N_34974,N_34644);
nor U36770 (N_36770,N_34736,N_30424);
nor U36771 (N_36771,N_30245,N_32341);
and U36772 (N_36772,N_33417,N_33172);
or U36773 (N_36773,N_34659,N_32857);
nor U36774 (N_36774,N_30248,N_30473);
and U36775 (N_36775,N_32393,N_33137);
or U36776 (N_36776,N_33538,N_32488);
xor U36777 (N_36777,N_30308,N_30706);
or U36778 (N_36778,N_30744,N_34263);
or U36779 (N_36779,N_30497,N_34909);
nor U36780 (N_36780,N_32719,N_32868);
and U36781 (N_36781,N_30462,N_33545);
and U36782 (N_36782,N_32745,N_33656);
nor U36783 (N_36783,N_31690,N_33258);
nor U36784 (N_36784,N_32464,N_32499);
xor U36785 (N_36785,N_31902,N_34339);
xor U36786 (N_36786,N_33032,N_33394);
nor U36787 (N_36787,N_30782,N_32770);
nor U36788 (N_36788,N_34732,N_34839);
nor U36789 (N_36789,N_30579,N_32183);
nor U36790 (N_36790,N_34589,N_31969);
nand U36791 (N_36791,N_32742,N_33967);
nand U36792 (N_36792,N_33772,N_34441);
nor U36793 (N_36793,N_30234,N_34265);
and U36794 (N_36794,N_33895,N_30076);
nand U36795 (N_36795,N_31135,N_34507);
xor U36796 (N_36796,N_31222,N_33071);
and U36797 (N_36797,N_34155,N_33461);
and U36798 (N_36798,N_33494,N_34929);
xor U36799 (N_36799,N_30863,N_32047);
and U36800 (N_36800,N_30913,N_33176);
xnor U36801 (N_36801,N_33086,N_31818);
or U36802 (N_36802,N_33835,N_34702);
or U36803 (N_36803,N_31955,N_31699);
and U36804 (N_36804,N_34686,N_34236);
xnor U36805 (N_36805,N_34944,N_31274);
and U36806 (N_36806,N_30385,N_31232);
nor U36807 (N_36807,N_33055,N_30017);
nor U36808 (N_36808,N_34898,N_33874);
and U36809 (N_36809,N_30764,N_32936);
nor U36810 (N_36810,N_30603,N_32177);
xor U36811 (N_36811,N_30200,N_31810);
or U36812 (N_36812,N_33815,N_33300);
nor U36813 (N_36813,N_31904,N_31030);
and U36814 (N_36814,N_33491,N_34539);
nor U36815 (N_36815,N_30457,N_33429);
nor U36816 (N_36816,N_34936,N_34170);
xnor U36817 (N_36817,N_30492,N_33126);
nor U36818 (N_36818,N_33522,N_33765);
or U36819 (N_36819,N_32419,N_30721);
and U36820 (N_36820,N_33493,N_32002);
and U36821 (N_36821,N_33739,N_34999);
or U36822 (N_36822,N_31616,N_34613);
nor U36823 (N_36823,N_30378,N_31287);
nand U36824 (N_36824,N_31090,N_32539);
nor U36825 (N_36825,N_33218,N_31060);
or U36826 (N_36826,N_33858,N_30401);
xor U36827 (N_36827,N_31482,N_31126);
or U36828 (N_36828,N_31213,N_31174);
or U36829 (N_36829,N_34385,N_31066);
or U36830 (N_36830,N_30058,N_34788);
and U36831 (N_36831,N_32663,N_33207);
or U36832 (N_36832,N_34398,N_30011);
or U36833 (N_36833,N_34082,N_32099);
nand U36834 (N_36834,N_34878,N_32245);
or U36835 (N_36835,N_34348,N_31243);
nor U36836 (N_36836,N_34894,N_31879);
or U36837 (N_36837,N_32102,N_33685);
and U36838 (N_36838,N_30587,N_32431);
nand U36839 (N_36839,N_33665,N_32254);
nand U36840 (N_36840,N_33280,N_30505);
nor U36841 (N_36841,N_34091,N_33889);
and U36842 (N_36842,N_32087,N_34963);
or U36843 (N_36843,N_33105,N_32879);
or U36844 (N_36844,N_30376,N_31559);
or U36845 (N_36845,N_31143,N_33393);
nor U36846 (N_36846,N_33199,N_31383);
or U36847 (N_36847,N_30889,N_31196);
and U36848 (N_36848,N_33627,N_30879);
and U36849 (N_36849,N_30134,N_30305);
xnor U36850 (N_36850,N_33302,N_31488);
xor U36851 (N_36851,N_33724,N_34315);
and U36852 (N_36852,N_30729,N_32696);
nand U36853 (N_36853,N_34903,N_32520);
xor U36854 (N_36854,N_32340,N_31341);
or U36855 (N_36855,N_30849,N_31389);
nand U36856 (N_36856,N_32358,N_30412);
nand U36857 (N_36857,N_33169,N_33938);
xnor U36858 (N_36858,N_33057,N_30362);
and U36859 (N_36859,N_32903,N_30159);
or U36860 (N_36860,N_33418,N_32556);
nand U36861 (N_36861,N_30048,N_31019);
nand U36862 (N_36862,N_30490,N_34905);
nor U36863 (N_36863,N_30013,N_31304);
or U36864 (N_36864,N_30319,N_34445);
and U36865 (N_36865,N_31170,N_33402);
xnor U36866 (N_36866,N_30752,N_31649);
and U36867 (N_36867,N_30838,N_32287);
nor U36868 (N_36868,N_30123,N_31585);
xnor U36869 (N_36869,N_30928,N_33314);
nor U36870 (N_36870,N_33384,N_32761);
or U36871 (N_36871,N_32475,N_33518);
nor U36872 (N_36872,N_31688,N_34495);
nor U36873 (N_36873,N_32185,N_33624);
xor U36874 (N_36874,N_32768,N_33171);
or U36875 (N_36875,N_34401,N_31966);
xnor U36876 (N_36876,N_32266,N_32292);
nand U36877 (N_36877,N_33745,N_32260);
and U36878 (N_36878,N_33382,N_32038);
and U36879 (N_36879,N_32705,N_32095);
and U36880 (N_36880,N_30063,N_34534);
xor U36881 (N_36881,N_30426,N_34879);
nand U36882 (N_36882,N_31526,N_31630);
nand U36883 (N_36883,N_33544,N_33483);
and U36884 (N_36884,N_30624,N_33893);
xnor U36885 (N_36885,N_31337,N_33872);
nor U36886 (N_36886,N_33883,N_34735);
nor U36887 (N_36887,N_33232,N_30422);
nor U36888 (N_36888,N_30677,N_32662);
nand U36889 (N_36889,N_32021,N_30188);
xor U36890 (N_36890,N_32373,N_30116);
nor U36891 (N_36891,N_30831,N_33549);
nand U36892 (N_36892,N_33524,N_30467);
or U36893 (N_36893,N_34934,N_32560);
nor U36894 (N_36894,N_34018,N_32429);
nor U36895 (N_36895,N_32540,N_33741);
nand U36896 (N_36896,N_31951,N_31401);
nand U36897 (N_36897,N_34643,N_34256);
xnor U36898 (N_36898,N_33262,N_33251);
or U36899 (N_36899,N_34210,N_33630);
xor U36900 (N_36900,N_31718,N_34988);
nor U36901 (N_36901,N_33711,N_32225);
nand U36902 (N_36902,N_33192,N_32115);
nor U36903 (N_36903,N_30404,N_34135);
nor U36904 (N_36904,N_30080,N_30689);
xnor U36905 (N_36905,N_34462,N_31664);
nand U36906 (N_36906,N_33514,N_33396);
nand U36907 (N_36907,N_33618,N_33075);
xor U36908 (N_36908,N_30417,N_33786);
nand U36909 (N_36909,N_34034,N_34043);
nor U36910 (N_36910,N_31741,N_33663);
and U36911 (N_36911,N_33264,N_32149);
xor U36912 (N_36912,N_30484,N_34629);
nand U36913 (N_36913,N_31564,N_31536);
nand U36914 (N_36914,N_33599,N_33167);
and U36915 (N_36915,N_33444,N_31475);
or U36916 (N_36916,N_34358,N_30609);
xor U36917 (N_36917,N_34558,N_34473);
xor U36918 (N_36918,N_33018,N_32839);
xnor U36919 (N_36919,N_32786,N_31635);
nor U36920 (N_36920,N_33323,N_31681);
or U36921 (N_36921,N_31260,N_33686);
or U36922 (N_36922,N_32771,N_32085);
nor U36923 (N_36923,N_34217,N_30359);
or U36924 (N_36924,N_30230,N_32243);
nor U36925 (N_36925,N_34444,N_33372);
nor U36926 (N_36926,N_30075,N_31571);
xnor U36927 (N_36927,N_30790,N_31994);
and U36928 (N_36928,N_33900,N_33812);
and U36929 (N_36929,N_34382,N_33691);
or U36930 (N_36930,N_30813,N_32472);
xor U36931 (N_36931,N_32985,N_31311);
nand U36932 (N_36932,N_30167,N_33716);
xnor U36933 (N_36933,N_32441,N_32445);
nor U36934 (N_36934,N_30088,N_30054);
xor U36935 (N_36935,N_33144,N_32916);
or U36936 (N_36936,N_31644,N_33863);
xnor U36937 (N_36937,N_32600,N_34720);
or U36938 (N_36938,N_32174,N_32764);
and U36939 (N_36939,N_34158,N_32380);
nor U36940 (N_36940,N_34499,N_34758);
nand U36941 (N_36941,N_30964,N_30192);
xnor U36942 (N_36942,N_33749,N_33853);
or U36943 (N_36943,N_30638,N_32747);
nand U36944 (N_36944,N_31769,N_30077);
nor U36945 (N_36945,N_30344,N_32816);
xor U36946 (N_36946,N_30083,N_33362);
xnor U36947 (N_36947,N_32405,N_34057);
xor U36948 (N_36948,N_33823,N_30005);
or U36949 (N_36949,N_31637,N_34942);
or U36950 (N_36950,N_30949,N_34361);
and U36951 (N_36951,N_30994,N_33987);
nand U36952 (N_36952,N_32550,N_30098);
or U36953 (N_36953,N_34764,N_34027);
and U36954 (N_36954,N_30874,N_31340);
and U36955 (N_36955,N_30541,N_30416);
xor U36956 (N_36956,N_30253,N_31923);
or U36957 (N_36957,N_34745,N_30957);
nand U36958 (N_36958,N_34047,N_30460);
nand U36959 (N_36959,N_31128,N_33862);
or U36960 (N_36960,N_33587,N_31221);
or U36961 (N_36961,N_32822,N_34701);
and U36962 (N_36962,N_32829,N_31485);
xnor U36963 (N_36963,N_30032,N_33719);
nor U36964 (N_36964,N_32670,N_34240);
and U36965 (N_36965,N_34202,N_33209);
nor U36966 (N_36966,N_34601,N_34866);
xor U36967 (N_36967,N_34893,N_32232);
xor U36968 (N_36968,N_30074,N_34815);
nor U36969 (N_36969,N_33790,N_33951);
xnor U36970 (N_36970,N_33576,N_34843);
or U36971 (N_36971,N_34725,N_34891);
or U36972 (N_36972,N_31211,N_30331);
nor U36973 (N_36973,N_32956,N_30792);
and U36974 (N_36974,N_33876,N_30061);
xnor U36975 (N_36975,N_32597,N_31486);
or U36976 (N_36976,N_31374,N_30282);
nor U36977 (N_36977,N_32634,N_31368);
nand U36978 (N_36978,N_30562,N_31850);
nand U36979 (N_36979,N_30894,N_30881);
nor U36980 (N_36980,N_32825,N_32146);
xnor U36981 (N_36981,N_32843,N_31271);
nand U36982 (N_36982,N_30328,N_30115);
and U36983 (N_36983,N_32976,N_31162);
or U36984 (N_36984,N_34188,N_33211);
and U36985 (N_36985,N_32589,N_32216);
or U36986 (N_36986,N_33438,N_32847);
nor U36987 (N_36987,N_31079,N_33824);
nor U36988 (N_36988,N_33718,N_30227);
nor U36989 (N_36989,N_34918,N_31362);
nor U36990 (N_36990,N_30108,N_30314);
nor U36991 (N_36991,N_32374,N_31984);
or U36992 (N_36992,N_30195,N_31419);
nand U36993 (N_36993,N_30420,N_30053);
and U36994 (N_36994,N_31594,N_33404);
nor U36995 (N_36995,N_33328,N_33116);
or U36996 (N_36996,N_33759,N_33221);
nor U36997 (N_36997,N_34780,N_32584);
xnor U36998 (N_36998,N_32497,N_30004);
and U36999 (N_36999,N_31739,N_33977);
or U37000 (N_37000,N_33339,N_31534);
and U37001 (N_37001,N_32137,N_31537);
xnor U37002 (N_37002,N_34058,N_33712);
xor U37003 (N_37003,N_32576,N_31306);
or U37004 (N_37004,N_31205,N_34687);
nand U37005 (N_37005,N_34090,N_30578);
nor U37006 (N_37006,N_34693,N_33249);
nand U37007 (N_37007,N_31395,N_31839);
nor U37008 (N_37008,N_33318,N_34630);
and U37009 (N_37009,N_32797,N_32983);
or U37010 (N_37010,N_31159,N_31257);
or U37011 (N_37011,N_30800,N_33648);
nand U37012 (N_37012,N_33450,N_32570);
or U37013 (N_37013,N_33482,N_34976);
nand U37014 (N_37014,N_32996,N_30560);
or U37015 (N_37015,N_31217,N_32394);
and U37016 (N_37016,N_32536,N_30296);
or U37017 (N_37017,N_30418,N_32735);
nand U37018 (N_37018,N_30106,N_34966);
nand U37019 (N_37019,N_32012,N_33605);
xor U37020 (N_37020,N_30604,N_34357);
and U37021 (N_37021,N_33503,N_34904);
or U37022 (N_37022,N_31349,N_31513);
nor U37023 (N_37023,N_32541,N_31658);
and U37024 (N_37024,N_31921,N_31728);
and U37025 (N_37025,N_31013,N_30294);
or U37026 (N_37026,N_34007,N_32551);
xor U37027 (N_37027,N_34873,N_34938);
nor U37028 (N_37028,N_33903,N_32754);
nand U37029 (N_37029,N_30661,N_33080);
xor U37030 (N_37030,N_32427,N_31808);
xnor U37031 (N_37031,N_30235,N_31497);
and U37032 (N_37032,N_32455,N_32369);
and U37033 (N_37033,N_33096,N_30850);
nor U37034 (N_37034,N_30572,N_33743);
and U37035 (N_37035,N_34968,N_30266);
nor U37036 (N_37036,N_31215,N_33996);
xnor U37037 (N_37037,N_32629,N_31619);
or U37038 (N_37038,N_31958,N_32277);
nor U37039 (N_37039,N_33841,N_33781);
or U37040 (N_37040,N_31714,N_31123);
or U37041 (N_37041,N_34694,N_32152);
and U37042 (N_37042,N_31422,N_34679);
and U37043 (N_37043,N_33389,N_33668);
nor U37044 (N_37044,N_30558,N_31725);
or U37045 (N_37045,N_32861,N_33451);
xor U37046 (N_37046,N_30573,N_34960);
nor U37047 (N_37047,N_31316,N_34840);
nand U37048 (N_37048,N_31983,N_32023);
nand U37049 (N_37049,N_31583,N_32509);
xnor U37050 (N_37050,N_30112,N_31129);
nand U37051 (N_37051,N_30340,N_33487);
or U37052 (N_37052,N_33159,N_31822);
nor U37053 (N_37053,N_34498,N_33008);
nor U37054 (N_37054,N_30275,N_34631);
xnor U37055 (N_37055,N_34955,N_34187);
xor U37056 (N_37056,N_30407,N_30241);
or U37057 (N_37057,N_33056,N_30481);
xnor U37058 (N_37058,N_30904,N_31847);
nand U37059 (N_37059,N_30126,N_31297);
nand U37060 (N_37060,N_34652,N_30699);
nand U37061 (N_37061,N_32253,N_33564);
nand U37062 (N_37062,N_33363,N_30498);
and U37063 (N_37063,N_32789,N_34541);
nor U37064 (N_37064,N_34008,N_33092);
or U37065 (N_37065,N_30260,N_32653);
or U37066 (N_37066,N_30886,N_31155);
xnor U37067 (N_37067,N_32709,N_32627);
nor U37068 (N_37068,N_30396,N_31235);
and U37069 (N_37069,N_30419,N_32364);
nor U37070 (N_37070,N_30767,N_31666);
xnor U37071 (N_37071,N_34665,N_30006);
and U37072 (N_37072,N_32179,N_32881);
and U37073 (N_37073,N_34528,N_32077);
nor U37074 (N_37074,N_31166,N_34807);
or U37075 (N_37075,N_34517,N_31737);
nor U37076 (N_37076,N_34291,N_34916);
xor U37077 (N_37077,N_34412,N_31676);
nand U37078 (N_37078,N_34930,N_30042);
and U37079 (N_37079,N_33542,N_32802);
nand U37080 (N_37080,N_33844,N_34002);
or U37081 (N_37081,N_34596,N_34777);
nand U37082 (N_37082,N_31648,N_34896);
nand U37083 (N_37083,N_31121,N_32826);
and U37084 (N_37084,N_31429,N_33616);
nor U37085 (N_37085,N_30178,N_30815);
nand U37086 (N_37086,N_32571,N_34819);
xor U37087 (N_37087,N_34712,N_32408);
xor U37088 (N_37088,N_31189,N_33768);
nor U37089 (N_37089,N_32289,N_34394);
xor U37090 (N_37090,N_33379,N_33846);
nand U37091 (N_37091,N_32390,N_33252);
xor U37092 (N_37092,N_32894,N_30670);
nor U37093 (N_37093,N_32836,N_30654);
xor U37094 (N_37094,N_30008,N_30574);
xnor U37095 (N_37095,N_34638,N_34026);
nand U37096 (N_37096,N_33785,N_33263);
nor U37097 (N_37097,N_30623,N_31715);
nand U37098 (N_37098,N_31618,N_33439);
nor U37099 (N_37099,N_34193,N_31055);
and U37100 (N_37100,N_32263,N_34179);
nand U37101 (N_37101,N_32048,N_30601);
nor U37102 (N_37102,N_32641,N_33446);
or U37103 (N_37103,N_30143,N_33465);
nand U37104 (N_37104,N_32057,N_30599);
nand U37105 (N_37105,N_33797,N_31442);
nor U37106 (N_37106,N_30528,N_33904);
nand U37107 (N_37107,N_32904,N_33367);
xnor U37108 (N_37108,N_30917,N_32176);
xor U37109 (N_37109,N_31720,N_31663);
nand U37110 (N_37110,N_32613,N_31385);
xor U37111 (N_37111,N_33101,N_30662);
xnor U37112 (N_37112,N_32303,N_34227);
xnor U37113 (N_37113,N_34379,N_33673);
or U37114 (N_37114,N_32221,N_34303);
and U37115 (N_37115,N_33007,N_34994);
nand U37116 (N_37116,N_34723,N_31971);
nand U37117 (N_37117,N_34399,N_31660);
or U37118 (N_37118,N_30732,N_34349);
and U37119 (N_37119,N_30945,N_33722);
xnor U37120 (N_37120,N_33019,N_30386);
nand U37121 (N_37121,N_34270,N_30537);
nor U37122 (N_37122,N_32438,N_32689);
nand U37123 (N_37123,N_31444,N_33708);
xnor U37124 (N_37124,N_33818,N_32961);
and U37125 (N_37125,N_34001,N_31595);
nor U37126 (N_37126,N_31938,N_31812);
nor U37127 (N_37127,N_34032,N_34363);
xnor U37128 (N_37128,N_31139,N_32766);
and U37129 (N_37129,N_34000,N_34019);
and U37130 (N_37130,N_34972,N_31312);
or U37131 (N_37131,N_34461,N_33311);
nor U37132 (N_37132,N_34805,N_31218);
or U37133 (N_37133,N_33142,N_33121);
and U37134 (N_37134,N_31533,N_33093);
nand U37135 (N_37135,N_30552,N_33129);
xor U37136 (N_37136,N_32911,N_34533);
xnor U37137 (N_37137,N_30226,N_34070);
nor U37138 (N_37138,N_34022,N_33952);
or U37139 (N_37139,N_31415,N_30525);
nand U37140 (N_37140,N_32418,N_34690);
or U37141 (N_37141,N_32568,N_33140);
or U37142 (N_37142,N_30916,N_33061);
nand U37143 (N_37143,N_32333,N_32256);
and U37144 (N_37144,N_34503,N_30448);
nor U37145 (N_37145,N_32375,N_33997);
xor U37146 (N_37146,N_34442,N_33769);
nor U37147 (N_37147,N_34430,N_31096);
nor U37148 (N_37148,N_30743,N_32376);
nand U37149 (N_37149,N_32368,N_34779);
or U37150 (N_37150,N_32939,N_33058);
xor U37151 (N_37151,N_31634,N_30205);
or U37152 (N_37152,N_32502,N_33299);
and U37153 (N_37153,N_30113,N_34176);
and U37154 (N_37154,N_34485,N_33869);
or U37155 (N_37155,N_34957,N_34396);
nor U37156 (N_37156,N_32134,N_34632);
nor U37157 (N_37157,N_34060,N_33937);
nor U37158 (N_37158,N_30051,N_31704);
nand U37159 (N_37159,N_31916,N_33674);
and U37160 (N_37160,N_31877,N_31854);
xor U37161 (N_37161,N_33041,N_30724);
and U37162 (N_37162,N_31197,N_33155);
xnor U37163 (N_37163,N_31599,N_34316);
or U37164 (N_37164,N_32037,N_33003);
nor U37165 (N_37165,N_31251,N_32661);
and U37166 (N_37166,N_30559,N_33723);
nor U37167 (N_37167,N_34926,N_30923);
and U37168 (N_37168,N_32687,N_30896);
nor U37169 (N_37169,N_31919,N_30067);
or U37170 (N_37170,N_34390,N_31947);
xor U37171 (N_37171,N_33489,N_31373);
or U37172 (N_37172,N_31363,N_31926);
and U37173 (N_37173,N_30432,N_32684);
xor U37174 (N_37174,N_31460,N_31560);
nand U37175 (N_37175,N_34220,N_33536);
nand U37176 (N_37176,N_31014,N_30546);
and U37177 (N_37177,N_34172,N_31029);
xnor U37178 (N_37178,N_30667,N_32529);
and U37179 (N_37179,N_30684,N_30970);
and U37180 (N_37180,N_30232,N_34914);
xor U37181 (N_37181,N_34782,N_32642);
xor U37182 (N_37182,N_34268,N_31967);
nor U37183 (N_37183,N_33799,N_32343);
and U37184 (N_37184,N_32014,N_32454);
nand U37185 (N_37185,N_34586,N_30614);
xor U37186 (N_37186,N_31880,N_30024);
nand U37187 (N_37187,N_31761,N_34203);
xnor U37188 (N_37188,N_33507,N_31575);
and U37189 (N_37189,N_31108,N_32239);
or U37190 (N_37190,N_30637,N_32387);
nor U37191 (N_37191,N_31765,N_33580);
and U37192 (N_37192,N_30925,N_34489);
or U37193 (N_37193,N_33606,N_30811);
nor U37194 (N_37194,N_34377,N_34911);
nand U37195 (N_37195,N_32272,N_33802);
nor U37196 (N_37196,N_32414,N_33957);
nor U37197 (N_37197,N_33421,N_30033);
and U37198 (N_37198,N_31809,N_30244);
or U37199 (N_37199,N_33084,N_30628);
or U37200 (N_37200,N_33484,N_32658);
and U37201 (N_37201,N_30563,N_32084);
or U37202 (N_37202,N_30391,N_30660);
nor U37203 (N_37203,N_34588,N_31047);
or U37204 (N_37204,N_33399,N_32315);
and U37205 (N_37205,N_30924,N_31729);
xor U37206 (N_37206,N_30486,N_30060);
nand U37207 (N_37207,N_30617,N_31837);
nor U37208 (N_37208,N_30348,N_34483);
xnor U37209 (N_37209,N_30177,N_30972);
nand U37210 (N_37210,N_31091,N_33881);
xor U37211 (N_37211,N_30150,N_32605);
or U37212 (N_37212,N_34703,N_33378);
xnor U37213 (N_37213,N_33706,N_30031);
nor U37214 (N_37214,N_30105,N_31321);
nor U37215 (N_37215,N_33330,N_32925);
xor U37216 (N_37216,N_33118,N_30007);
nand U37217 (N_37217,N_31282,N_30856);
or U37218 (N_37218,N_33730,N_31124);
nand U37219 (N_37219,N_30823,N_33247);
nor U37220 (N_37220,N_34319,N_34088);
or U37221 (N_37221,N_33325,N_30690);
nand U37222 (N_37222,N_30600,N_34087);
nor U37223 (N_37223,N_32302,N_30771);
or U37224 (N_37224,N_31053,N_34238);
xor U37225 (N_37225,N_32855,N_30993);
nand U37226 (N_37226,N_33748,N_30538);
nor U37227 (N_37227,N_34023,N_30902);
and U37228 (N_37228,N_32270,N_34524);
nor U37229 (N_37229,N_33516,N_32278);
xor U37230 (N_37230,N_33629,N_31977);
or U37231 (N_37231,N_31198,N_30803);
xnor U37232 (N_37232,N_32931,N_32148);
nand U37233 (N_37233,N_30438,N_31181);
and U37234 (N_37234,N_31399,N_32963);
and U37235 (N_37235,N_32336,N_34576);
nor U37236 (N_37236,N_33353,N_31551);
and U37237 (N_37237,N_30504,N_30826);
nor U37238 (N_37238,N_34587,N_33762);
or U37239 (N_37239,N_33257,N_31684);
or U37240 (N_37240,N_32141,N_33640);
nand U37241 (N_37241,N_31900,N_31948);
nand U37242 (N_37242,N_34275,N_32361);
and U37243 (N_37243,N_30430,N_30506);
xor U37244 (N_37244,N_31876,N_34954);
nand U37245 (N_37245,N_31432,N_31231);
nor U37246 (N_37246,N_31177,N_30530);
or U37247 (N_37247,N_32231,N_30720);
nor U37248 (N_37248,N_33859,N_34343);
or U37249 (N_37249,N_32465,N_31538);
xor U37250 (N_37250,N_31531,N_31867);
nor U37251 (N_37251,N_31276,N_33529);
or U37252 (N_37252,N_31152,N_30700);
nand U37253 (N_37253,N_32787,N_33475);
and U37254 (N_37254,N_31468,N_30341);
xor U37255 (N_37255,N_33376,N_33072);
and U37256 (N_37256,N_32267,N_31601);
xor U37257 (N_37257,N_34500,N_33434);
nor U37258 (N_37258,N_32080,N_32351);
nor U37259 (N_37259,N_34438,N_34325);
nand U37260 (N_37260,N_30655,N_32391);
and U37261 (N_37261,N_31786,N_32192);
nand U37262 (N_37262,N_34464,N_32034);
nor U37263 (N_37263,N_30971,N_33094);
xnor U37264 (N_37264,N_33403,N_30987);
or U37265 (N_37265,N_31673,N_34978);
nand U37266 (N_37266,N_31050,N_34685);
nand U37267 (N_37267,N_33179,N_30493);
xnor U37268 (N_37268,N_32814,N_33634);
and U37269 (N_37269,N_33681,N_31357);
nor U37270 (N_37270,N_33527,N_34449);
nor U37271 (N_37271,N_33165,N_34591);
and U37272 (N_37272,N_31697,N_34328);
xnor U37273 (N_37273,N_31065,N_32557);
xor U37274 (N_37274,N_33886,N_33720);
or U37275 (N_37275,N_30797,N_31936);
or U37276 (N_37276,N_33117,N_33684);
nor U37277 (N_37277,N_33870,N_34740);
xnor U37278 (N_37278,N_30086,N_30930);
and U37279 (N_37279,N_32821,N_32815);
xnor U37280 (N_37280,N_30209,N_34579);
and U37281 (N_37281,N_31972,N_32947);
and U37282 (N_37282,N_34640,N_30474);
nand U37283 (N_37283,N_32076,N_32500);
and U37284 (N_37284,N_32492,N_34864);
nand U37285 (N_37285,N_30642,N_32665);
or U37286 (N_37286,N_31627,N_31245);
and U37287 (N_37287,N_33574,N_32573);
nor U37288 (N_37288,N_31355,N_33757);
nor U37289 (N_37289,N_33412,N_31698);
and U37290 (N_37290,N_31540,N_31724);
and U37291 (N_37291,N_33737,N_30676);
nand U37292 (N_37292,N_30739,N_32812);
or U37293 (N_37293,N_32485,N_33135);
and U37294 (N_37294,N_31457,N_30441);
or U37295 (N_37295,N_34152,N_30478);
or U37296 (N_37296,N_30087,N_32417);
or U37297 (N_37297,N_30351,N_33500);
nand U37298 (N_37298,N_32749,N_34131);
and U37299 (N_37299,N_32852,N_33006);
nand U37300 (N_37300,N_33831,N_33295);
nand U37301 (N_37301,N_30730,N_34768);
nand U37302 (N_37302,N_32772,N_30747);
or U37303 (N_37303,N_30675,N_31480);
nand U37304 (N_37304,N_33463,N_31776);
or U37305 (N_37305,N_34476,N_33423);
xnor U37306 (N_37306,N_32875,N_34086);
nor U37307 (N_37307,N_34169,N_33219);
nand U37308 (N_37308,N_31360,N_33822);
and U37309 (N_37309,N_33123,N_33040);
xnor U37310 (N_37310,N_34474,N_33669);
and U37311 (N_37311,N_34260,N_32737);
nand U37312 (N_37312,N_32434,N_31964);
nor U37313 (N_37313,N_32195,N_32615);
nor U37314 (N_37314,N_34437,N_32151);
and U37315 (N_37315,N_30131,N_34818);
xnor U37316 (N_37316,N_34982,N_30998);
and U37317 (N_37317,N_30240,N_33679);
or U37318 (N_37318,N_34424,N_32831);
and U37319 (N_37319,N_32510,N_33899);
xor U37320 (N_37320,N_31353,N_34990);
or U37321 (N_37321,N_31516,N_32680);
nor U37322 (N_37322,N_32654,N_34432);
nor U37323 (N_37323,N_33136,N_31679);
and U37324 (N_37324,N_33887,N_30934);
nor U37325 (N_37325,N_30950,N_32877);
and U37326 (N_37326,N_33751,N_34289);
or U37327 (N_37327,N_32598,N_33603);
nor U37328 (N_37328,N_30632,N_30943);
and U37329 (N_37329,N_34061,N_34809);
nand U37330 (N_37330,N_31626,N_33794);
and U37331 (N_37331,N_32645,N_31411);
or U37332 (N_37332,N_32892,N_31119);
and U37333 (N_37333,N_33750,N_34943);
nand U37334 (N_37334,N_30616,N_33324);
nand U37335 (N_37335,N_30550,N_34183);
or U37336 (N_37336,N_33607,N_33274);
and U37337 (N_37337,N_30668,N_31458);
and U37338 (N_37338,N_34109,N_32739);
and U37339 (N_37339,N_32522,N_32432);
nor U37340 (N_37340,N_34230,N_34922);
or U37341 (N_37341,N_34762,N_31865);
xor U37342 (N_37342,N_32878,N_33154);
xor U37343 (N_37343,N_33770,N_34870);
xnor U37344 (N_37344,N_33184,N_30104);
or U37345 (N_37345,N_31184,N_34850);
or U37346 (N_37346,N_34068,N_32252);
or U37347 (N_37347,N_31623,N_34181);
xnor U37348 (N_37348,N_30499,N_32323);
nor U37349 (N_37349,N_31979,N_32565);
or U37350 (N_37350,N_31388,N_34682);
xor U37351 (N_37351,N_30297,N_31195);
nor U37352 (N_37352,N_32157,N_34724);
xnor U37353 (N_37353,N_33152,N_30536);
xor U37354 (N_37354,N_33427,N_32593);
nor U37355 (N_37355,N_32799,N_30779);
or U37356 (N_37356,N_34353,N_32160);
nor U37357 (N_37357,N_34261,N_31117);
or U37358 (N_37358,N_33440,N_30449);
xor U37359 (N_37359,N_30817,N_31727);
or U37360 (N_37360,N_33198,N_34869);
or U37361 (N_37361,N_33572,N_30980);
nor U37362 (N_37362,N_33273,N_32873);
nand U37363 (N_37363,N_31127,N_33643);
nor U37364 (N_37364,N_33531,N_32031);
and U37365 (N_37365,N_31506,N_31328);
nor U37366 (N_37366,N_34856,N_32938);
xnor U37367 (N_37367,N_30435,N_30184);
nor U37368 (N_37368,N_34201,N_31075);
or U37369 (N_37369,N_34515,N_31647);
nand U37370 (N_37370,N_31842,N_31749);
xor U37371 (N_37371,N_31320,N_30237);
or U37372 (N_37372,N_31545,N_34100);
nand U37373 (N_37373,N_32564,N_32534);
and U37374 (N_37374,N_32724,N_31841);
and U37375 (N_37375,N_34171,N_34177);
nor U37376 (N_37376,N_32840,N_30251);
and U37377 (N_37377,N_33710,N_33381);
nand U37378 (N_37378,N_31578,N_32889);
nor U37379 (N_37379,N_31185,N_32657);
xnor U37380 (N_37380,N_31549,N_32998);
xor U37381 (N_37381,N_30324,N_34400);
or U37382 (N_37382,N_31745,N_34113);
xnor U37383 (N_37383,N_31496,N_30012);
or U37384 (N_37384,N_32235,N_31239);
nand U37385 (N_37385,N_30583,N_31265);
xor U37386 (N_37386,N_31086,N_30612);
or U37387 (N_37387,N_34243,N_33070);
and U37388 (N_37388,N_31738,N_33288);
and U37389 (N_37389,N_32007,N_31832);
and U37390 (N_37390,N_31020,N_33125);
xor U37391 (N_37391,N_33190,N_34387);
xnor U37392 (N_37392,N_31541,N_33391);
xnor U37393 (N_37393,N_32611,N_32224);
nand U37394 (N_37394,N_33555,N_30491);
and U37395 (N_37395,N_31279,N_32457);
nand U37396 (N_37396,N_33666,N_30320);
or U37397 (N_37397,N_34050,N_32693);
and U37398 (N_37398,N_32999,N_32297);
xor U37399 (N_37399,N_34411,N_33095);
xor U37400 (N_37400,N_32965,N_30828);
or U37401 (N_37401,N_32436,N_34616);
xnor U37402 (N_37402,N_30555,N_32794);
and U37403 (N_37403,N_30608,N_30309);
nor U37404 (N_37404,N_32167,N_30705);
nor U37405 (N_37405,N_30553,N_34722);
and U37406 (N_37406,N_31036,N_32257);
nor U37407 (N_37407,N_31025,N_30694);
and U37408 (N_37408,N_34981,N_33847);
nand U37409 (N_37409,N_34089,N_32990);
xor U37410 (N_37410,N_33035,N_31006);
nor U37411 (N_37411,N_32941,N_32851);
xnor U37412 (N_37412,N_32558,N_33866);
nand U37413 (N_37413,N_33447,N_32094);
xor U37414 (N_37414,N_34457,N_34928);
nor U37415 (N_37415,N_34783,N_33181);
nor U37416 (N_37416,N_34427,N_33293);
nor U37417 (N_37417,N_30322,N_30872);
or U37418 (N_37418,N_30982,N_31169);
nor U37419 (N_37419,N_33036,N_34519);
nand U37420 (N_37420,N_33864,N_31416);
nor U37421 (N_37421,N_33490,N_33466);
or U37422 (N_37422,N_30395,N_34556);
and U37423 (N_37423,N_31299,N_34521);
nand U37424 (N_37424,N_31707,N_32129);
xnor U37425 (N_37425,N_32273,N_32993);
or U37426 (N_37426,N_34967,N_32746);
or U37427 (N_37427,N_34655,N_33470);
or U37428 (N_37428,N_30818,N_31382);
or U37429 (N_37429,N_31112,N_31489);
and U37430 (N_37430,N_30285,N_32635);
nand U37431 (N_37431,N_30785,N_32486);
nand U37432 (N_37432,N_33619,N_33210);
or U37433 (N_37433,N_30715,N_31529);
xor U37434 (N_37434,N_30157,N_31044);
xnor U37435 (N_37435,N_32774,N_32858);
nor U37436 (N_37436,N_32606,N_32751);
nor U37437 (N_37437,N_33947,N_30302);
and U37438 (N_37438,N_31568,N_31779);
xnor U37439 (N_37439,N_34150,N_33597);
and U37440 (N_37440,N_33236,N_32083);
nor U37441 (N_37441,N_32066,N_31105);
or U37442 (N_37442,N_33919,N_31689);
xnor U37443 (N_37443,N_31752,N_31831);
nor U37444 (N_37444,N_34447,N_30249);
xor U37445 (N_37445,N_32450,N_32962);
nor U37446 (N_37446,N_33452,N_31624);
or U37447 (N_37447,N_34612,N_33361);
and U37448 (N_37448,N_32205,N_34209);
nand U37449 (N_37449,N_34095,N_31503);
nor U37450 (N_37450,N_34410,N_32024);
and U37451 (N_37451,N_32249,N_32069);
nor U37452 (N_37452,N_34707,N_32926);
or U37453 (N_37453,N_31586,N_30089);
nand U37454 (N_37454,N_31799,N_34294);
and U37455 (N_37455,N_30479,N_32518);
and U37456 (N_37456,N_34030,N_34416);
nand U37457 (N_37457,N_34381,N_32955);
nor U37458 (N_37458,N_30966,N_31294);
nor U37459 (N_37459,N_31763,N_34114);
nand U37460 (N_37460,N_31204,N_31021);
xnor U37461 (N_37461,N_32884,N_34467);
or U37462 (N_37462,N_34097,N_33014);
nor U37463 (N_37463,N_34675,N_31350);
and U37464 (N_37464,N_33082,N_30570);
and U37465 (N_37465,N_33637,N_30814);
or U37466 (N_37466,N_30910,N_34804);
or U37467 (N_37467,N_31574,N_34886);
or U37468 (N_37468,N_31138,N_30278);
xnor U37469 (N_37469,N_33340,N_33194);
nand U37470 (N_37470,N_32325,N_30963);
xor U37471 (N_37471,N_34836,N_31868);
and U37472 (N_37472,N_31920,N_31845);
nand U37473 (N_37473,N_30640,N_30621);
nor U37474 (N_37474,N_32474,N_32462);
or U37475 (N_37475,N_31199,N_33796);
or U37476 (N_37476,N_31210,N_31190);
and U37477 (N_37477,N_34373,N_34066);
and U37478 (N_37478,N_34750,N_34514);
or U37479 (N_37479,N_33012,N_34664);
or U37480 (N_37480,N_31144,N_30000);
nor U37481 (N_37481,N_33926,N_33320);
or U37482 (N_37482,N_32346,N_32367);
xor U37483 (N_37483,N_32914,N_34145);
xnor U37484 (N_37484,N_32942,N_33676);
xnor U37485 (N_37485,N_33917,N_31946);
and U37486 (N_37486,N_31941,N_32638);
xnor U37487 (N_37487,N_32930,N_30290);
nor U37488 (N_37488,N_32025,N_33066);
nand U37489 (N_37489,N_30888,N_33224);
nor U37490 (N_37490,N_31760,N_30358);
nor U37491 (N_37491,N_34094,N_32155);
nor U37492 (N_37492,N_34127,N_32269);
and U37493 (N_37493,N_31032,N_33454);
xnor U37494 (N_37494,N_32893,N_34593);
or U37495 (N_37495,N_33586,N_30976);
nor U37496 (N_37496,N_31233,N_30383);
xnor U37497 (N_37497,N_30326,N_30207);
nand U37498 (N_37498,N_32128,N_34014);
xnor U37499 (N_37499,N_31509,N_32572);
and U37500 (N_37500,N_30054,N_30443);
and U37501 (N_37501,N_30913,N_30813);
or U37502 (N_37502,N_34241,N_30972);
nor U37503 (N_37503,N_31515,N_34853);
or U37504 (N_37504,N_34830,N_31021);
or U37505 (N_37505,N_32031,N_33433);
nand U37506 (N_37506,N_30598,N_33208);
or U37507 (N_37507,N_34868,N_30553);
nor U37508 (N_37508,N_31162,N_32628);
xnor U37509 (N_37509,N_33283,N_33337);
xor U37510 (N_37510,N_32660,N_33250);
or U37511 (N_37511,N_32737,N_31377);
or U37512 (N_37512,N_30978,N_32635);
xor U37513 (N_37513,N_33417,N_33478);
and U37514 (N_37514,N_34628,N_33067);
or U37515 (N_37515,N_32051,N_33911);
nand U37516 (N_37516,N_31781,N_31415);
xnor U37517 (N_37517,N_31204,N_30407);
or U37518 (N_37518,N_32092,N_33702);
nand U37519 (N_37519,N_31094,N_34349);
nand U37520 (N_37520,N_34497,N_32100);
xor U37521 (N_37521,N_31948,N_34171);
nor U37522 (N_37522,N_33084,N_33125);
nor U37523 (N_37523,N_32000,N_33150);
nor U37524 (N_37524,N_33989,N_34121);
nand U37525 (N_37525,N_32750,N_32245);
nand U37526 (N_37526,N_31460,N_30383);
nor U37527 (N_37527,N_33140,N_31781);
nor U37528 (N_37528,N_32444,N_30661);
and U37529 (N_37529,N_32446,N_33280);
or U37530 (N_37530,N_30604,N_30564);
or U37531 (N_37531,N_34716,N_33343);
nand U37532 (N_37532,N_31103,N_34745);
and U37533 (N_37533,N_30667,N_31059);
nor U37534 (N_37534,N_34531,N_32135);
and U37535 (N_37535,N_30707,N_30559);
and U37536 (N_37536,N_31319,N_30648);
nand U37537 (N_37537,N_33235,N_31799);
nand U37538 (N_37538,N_32780,N_33109);
xnor U37539 (N_37539,N_34876,N_34136);
and U37540 (N_37540,N_32225,N_33456);
nor U37541 (N_37541,N_34353,N_31994);
nor U37542 (N_37542,N_34340,N_32613);
nor U37543 (N_37543,N_30408,N_32572);
xnor U37544 (N_37544,N_34168,N_33792);
nand U37545 (N_37545,N_33531,N_34998);
and U37546 (N_37546,N_33018,N_30229);
and U37547 (N_37547,N_32824,N_30713);
xnor U37548 (N_37548,N_33579,N_32122);
or U37549 (N_37549,N_32067,N_33133);
and U37550 (N_37550,N_30856,N_31628);
nand U37551 (N_37551,N_33406,N_32000);
nand U37552 (N_37552,N_32767,N_31537);
nor U37553 (N_37553,N_31401,N_31514);
nand U37554 (N_37554,N_34479,N_33810);
nand U37555 (N_37555,N_30986,N_33585);
nor U37556 (N_37556,N_31855,N_30763);
or U37557 (N_37557,N_31585,N_32245);
nor U37558 (N_37558,N_34947,N_32978);
or U37559 (N_37559,N_30102,N_34927);
nand U37560 (N_37560,N_33899,N_31428);
or U37561 (N_37561,N_31675,N_34014);
nand U37562 (N_37562,N_31371,N_34203);
nor U37563 (N_37563,N_31986,N_34558);
nand U37564 (N_37564,N_33268,N_31120);
xnor U37565 (N_37565,N_32347,N_31847);
nand U37566 (N_37566,N_34329,N_33405);
nor U37567 (N_37567,N_30533,N_30288);
and U37568 (N_37568,N_32032,N_32728);
nand U37569 (N_37569,N_31232,N_32396);
or U37570 (N_37570,N_30543,N_30081);
nor U37571 (N_37571,N_30987,N_34641);
nor U37572 (N_37572,N_31372,N_31221);
or U37573 (N_37573,N_34850,N_33212);
xnor U37574 (N_37574,N_32572,N_31252);
xnor U37575 (N_37575,N_32980,N_31524);
and U37576 (N_37576,N_30747,N_30332);
nand U37577 (N_37577,N_31960,N_30720);
nor U37578 (N_37578,N_30393,N_34863);
xor U37579 (N_37579,N_34259,N_34253);
or U37580 (N_37580,N_34186,N_34792);
and U37581 (N_37581,N_30681,N_30618);
and U37582 (N_37582,N_33768,N_32719);
or U37583 (N_37583,N_33392,N_30181);
nor U37584 (N_37584,N_33662,N_31473);
and U37585 (N_37585,N_30702,N_32798);
or U37586 (N_37586,N_34227,N_30066);
nor U37587 (N_37587,N_34163,N_30131);
nor U37588 (N_37588,N_31060,N_30755);
and U37589 (N_37589,N_31799,N_31930);
nand U37590 (N_37590,N_33300,N_31856);
nand U37591 (N_37591,N_31008,N_34122);
or U37592 (N_37592,N_31777,N_32140);
nor U37593 (N_37593,N_31843,N_31792);
and U37594 (N_37594,N_33703,N_30089);
and U37595 (N_37595,N_32300,N_32216);
nand U37596 (N_37596,N_33387,N_30145);
xnor U37597 (N_37597,N_32411,N_31670);
and U37598 (N_37598,N_31042,N_34611);
or U37599 (N_37599,N_33297,N_33445);
or U37600 (N_37600,N_34129,N_32979);
nor U37601 (N_37601,N_30026,N_30896);
xor U37602 (N_37602,N_31238,N_32749);
and U37603 (N_37603,N_31033,N_34095);
or U37604 (N_37604,N_32027,N_30951);
nor U37605 (N_37605,N_34100,N_31593);
or U37606 (N_37606,N_33796,N_30351);
nor U37607 (N_37607,N_30637,N_34084);
nor U37608 (N_37608,N_33292,N_33430);
or U37609 (N_37609,N_32627,N_31709);
xnor U37610 (N_37610,N_31133,N_34179);
and U37611 (N_37611,N_34635,N_31229);
nor U37612 (N_37612,N_34645,N_32772);
xnor U37613 (N_37613,N_32091,N_32115);
nand U37614 (N_37614,N_33182,N_31081);
and U37615 (N_37615,N_30218,N_32563);
nor U37616 (N_37616,N_34530,N_34847);
nand U37617 (N_37617,N_34555,N_30155);
nor U37618 (N_37618,N_34605,N_31057);
nor U37619 (N_37619,N_30284,N_34925);
and U37620 (N_37620,N_32786,N_31225);
nand U37621 (N_37621,N_31370,N_33688);
and U37622 (N_37622,N_34123,N_30760);
or U37623 (N_37623,N_32412,N_30532);
and U37624 (N_37624,N_33564,N_30034);
or U37625 (N_37625,N_30688,N_33843);
and U37626 (N_37626,N_32273,N_34575);
nand U37627 (N_37627,N_33085,N_30067);
nand U37628 (N_37628,N_32676,N_31079);
nand U37629 (N_37629,N_31137,N_30888);
nand U37630 (N_37630,N_32623,N_32198);
and U37631 (N_37631,N_32200,N_33801);
or U37632 (N_37632,N_30740,N_31643);
or U37633 (N_37633,N_34451,N_32029);
nand U37634 (N_37634,N_30460,N_30650);
nand U37635 (N_37635,N_30273,N_32360);
and U37636 (N_37636,N_31426,N_34865);
nor U37637 (N_37637,N_31363,N_32802);
or U37638 (N_37638,N_31220,N_34051);
and U37639 (N_37639,N_31115,N_33622);
xnor U37640 (N_37640,N_32122,N_31269);
and U37641 (N_37641,N_31418,N_33873);
and U37642 (N_37642,N_32606,N_34508);
and U37643 (N_37643,N_34264,N_32674);
xnor U37644 (N_37644,N_31496,N_32610);
nand U37645 (N_37645,N_33503,N_30890);
nor U37646 (N_37646,N_31988,N_32735);
nand U37647 (N_37647,N_33854,N_30393);
nand U37648 (N_37648,N_30047,N_32593);
xnor U37649 (N_37649,N_31038,N_32084);
xnor U37650 (N_37650,N_30978,N_31284);
nor U37651 (N_37651,N_34518,N_30479);
and U37652 (N_37652,N_30914,N_34779);
nor U37653 (N_37653,N_33840,N_33407);
and U37654 (N_37654,N_34506,N_30797);
nand U37655 (N_37655,N_31404,N_31201);
or U37656 (N_37656,N_33002,N_32417);
and U37657 (N_37657,N_33729,N_34543);
nor U37658 (N_37658,N_33461,N_31625);
nor U37659 (N_37659,N_34974,N_32130);
or U37660 (N_37660,N_34113,N_32172);
nor U37661 (N_37661,N_32744,N_33075);
xnor U37662 (N_37662,N_31462,N_33715);
xnor U37663 (N_37663,N_32001,N_32339);
nand U37664 (N_37664,N_34139,N_33765);
and U37665 (N_37665,N_32186,N_33067);
nand U37666 (N_37666,N_30471,N_31110);
nand U37667 (N_37667,N_33238,N_33540);
nand U37668 (N_37668,N_31480,N_30771);
nand U37669 (N_37669,N_33483,N_34135);
nand U37670 (N_37670,N_31438,N_31615);
and U37671 (N_37671,N_30895,N_32926);
nand U37672 (N_37672,N_30557,N_33997);
nor U37673 (N_37673,N_31617,N_30038);
nor U37674 (N_37674,N_33173,N_31193);
and U37675 (N_37675,N_34706,N_31743);
nand U37676 (N_37676,N_32526,N_32144);
nor U37677 (N_37677,N_34447,N_32663);
nor U37678 (N_37678,N_31875,N_33953);
nand U37679 (N_37679,N_31394,N_31808);
nor U37680 (N_37680,N_30728,N_34975);
and U37681 (N_37681,N_30351,N_30006);
nand U37682 (N_37682,N_31549,N_34520);
nand U37683 (N_37683,N_34813,N_32980);
nand U37684 (N_37684,N_31197,N_32253);
xnor U37685 (N_37685,N_34476,N_32343);
or U37686 (N_37686,N_30380,N_32459);
nor U37687 (N_37687,N_31544,N_32323);
xor U37688 (N_37688,N_30226,N_30731);
nor U37689 (N_37689,N_30707,N_31278);
nand U37690 (N_37690,N_32684,N_32905);
and U37691 (N_37691,N_31585,N_31730);
nor U37692 (N_37692,N_32771,N_31679);
and U37693 (N_37693,N_30511,N_34989);
nand U37694 (N_37694,N_33542,N_30289);
nor U37695 (N_37695,N_34706,N_33333);
xor U37696 (N_37696,N_30280,N_33859);
and U37697 (N_37697,N_32395,N_33766);
and U37698 (N_37698,N_34072,N_32345);
or U37699 (N_37699,N_32248,N_31957);
nor U37700 (N_37700,N_33718,N_32422);
xor U37701 (N_37701,N_34185,N_31154);
or U37702 (N_37702,N_30055,N_31009);
nor U37703 (N_37703,N_32880,N_34072);
xor U37704 (N_37704,N_32084,N_31439);
nor U37705 (N_37705,N_33318,N_34249);
or U37706 (N_37706,N_32313,N_30709);
or U37707 (N_37707,N_33247,N_32370);
and U37708 (N_37708,N_33948,N_34116);
nand U37709 (N_37709,N_30694,N_32272);
nor U37710 (N_37710,N_34124,N_31401);
and U37711 (N_37711,N_34945,N_34434);
xor U37712 (N_37712,N_34077,N_34004);
nor U37713 (N_37713,N_32594,N_30469);
xnor U37714 (N_37714,N_34469,N_34286);
or U37715 (N_37715,N_32712,N_33213);
and U37716 (N_37716,N_33726,N_34063);
and U37717 (N_37717,N_32961,N_34379);
nand U37718 (N_37718,N_32640,N_34911);
or U37719 (N_37719,N_30824,N_34520);
nand U37720 (N_37720,N_34800,N_31461);
and U37721 (N_37721,N_33767,N_33813);
xor U37722 (N_37722,N_31485,N_33674);
and U37723 (N_37723,N_34872,N_31191);
xnor U37724 (N_37724,N_31459,N_31767);
or U37725 (N_37725,N_32494,N_34212);
xnor U37726 (N_37726,N_31792,N_30308);
or U37727 (N_37727,N_31826,N_32061);
xor U37728 (N_37728,N_33712,N_31068);
nor U37729 (N_37729,N_30606,N_33398);
nand U37730 (N_37730,N_31727,N_31447);
and U37731 (N_37731,N_30490,N_31159);
or U37732 (N_37732,N_31855,N_33652);
or U37733 (N_37733,N_34796,N_33716);
nor U37734 (N_37734,N_31512,N_30097);
or U37735 (N_37735,N_30121,N_30481);
xnor U37736 (N_37736,N_30539,N_31385);
nor U37737 (N_37737,N_32802,N_33464);
nand U37738 (N_37738,N_30703,N_34446);
nor U37739 (N_37739,N_32446,N_33200);
xnor U37740 (N_37740,N_34967,N_33633);
nand U37741 (N_37741,N_31872,N_30214);
and U37742 (N_37742,N_32887,N_34485);
xor U37743 (N_37743,N_33795,N_32613);
xor U37744 (N_37744,N_32220,N_32380);
and U37745 (N_37745,N_32949,N_34367);
xor U37746 (N_37746,N_33890,N_32175);
and U37747 (N_37747,N_33017,N_33868);
or U37748 (N_37748,N_32818,N_31793);
xor U37749 (N_37749,N_32280,N_30064);
xor U37750 (N_37750,N_31494,N_33190);
nand U37751 (N_37751,N_31034,N_30223);
nor U37752 (N_37752,N_34546,N_31695);
and U37753 (N_37753,N_32409,N_30486);
xnor U37754 (N_37754,N_31659,N_31851);
nand U37755 (N_37755,N_34712,N_30194);
nand U37756 (N_37756,N_30049,N_34188);
nand U37757 (N_37757,N_30240,N_34015);
xor U37758 (N_37758,N_30128,N_32413);
nor U37759 (N_37759,N_32976,N_32635);
or U37760 (N_37760,N_31362,N_30900);
nand U37761 (N_37761,N_30679,N_33065);
and U37762 (N_37762,N_30208,N_32800);
xnor U37763 (N_37763,N_33692,N_34868);
nand U37764 (N_37764,N_31011,N_32468);
xnor U37765 (N_37765,N_30093,N_32625);
and U37766 (N_37766,N_33758,N_32387);
xor U37767 (N_37767,N_30314,N_34779);
or U37768 (N_37768,N_30581,N_32934);
nand U37769 (N_37769,N_32612,N_30271);
xor U37770 (N_37770,N_33889,N_31578);
nand U37771 (N_37771,N_31212,N_30680);
and U37772 (N_37772,N_31036,N_30517);
xnor U37773 (N_37773,N_33779,N_30142);
and U37774 (N_37774,N_33864,N_34697);
nor U37775 (N_37775,N_33493,N_32196);
nand U37776 (N_37776,N_34474,N_34141);
and U37777 (N_37777,N_31490,N_33166);
nor U37778 (N_37778,N_32369,N_31774);
nand U37779 (N_37779,N_31416,N_30037);
xnor U37780 (N_37780,N_31458,N_32731);
or U37781 (N_37781,N_33437,N_33667);
or U37782 (N_37782,N_33098,N_31757);
or U37783 (N_37783,N_32143,N_34411);
nand U37784 (N_37784,N_34681,N_31432);
and U37785 (N_37785,N_31173,N_33613);
nor U37786 (N_37786,N_31532,N_30210);
nand U37787 (N_37787,N_30200,N_34402);
nand U37788 (N_37788,N_34266,N_33422);
nor U37789 (N_37789,N_33624,N_31229);
nor U37790 (N_37790,N_31071,N_31483);
or U37791 (N_37791,N_34942,N_33570);
nor U37792 (N_37792,N_33417,N_31191);
or U37793 (N_37793,N_34648,N_30031);
nor U37794 (N_37794,N_33367,N_33503);
or U37795 (N_37795,N_31573,N_31606);
nor U37796 (N_37796,N_34251,N_33587);
xnor U37797 (N_37797,N_34472,N_34119);
nand U37798 (N_37798,N_30956,N_33226);
and U37799 (N_37799,N_31458,N_33386);
nor U37800 (N_37800,N_31037,N_34922);
nand U37801 (N_37801,N_31874,N_32785);
nand U37802 (N_37802,N_30080,N_31344);
xor U37803 (N_37803,N_33667,N_30714);
xnor U37804 (N_37804,N_34345,N_32347);
or U37805 (N_37805,N_32758,N_34882);
and U37806 (N_37806,N_31339,N_31728);
xor U37807 (N_37807,N_31926,N_34890);
xor U37808 (N_37808,N_33122,N_32357);
nor U37809 (N_37809,N_32521,N_31050);
nor U37810 (N_37810,N_30794,N_31028);
nand U37811 (N_37811,N_33073,N_31030);
nand U37812 (N_37812,N_34975,N_34202);
and U37813 (N_37813,N_34321,N_31497);
and U37814 (N_37814,N_34620,N_31953);
nor U37815 (N_37815,N_31706,N_32741);
xnor U37816 (N_37816,N_30110,N_30790);
nor U37817 (N_37817,N_31664,N_33991);
or U37818 (N_37818,N_31483,N_33597);
nor U37819 (N_37819,N_31312,N_34628);
or U37820 (N_37820,N_30320,N_33728);
nor U37821 (N_37821,N_30462,N_33926);
and U37822 (N_37822,N_32890,N_33524);
and U37823 (N_37823,N_33672,N_33468);
nand U37824 (N_37824,N_34131,N_34914);
or U37825 (N_37825,N_30156,N_32713);
nand U37826 (N_37826,N_34440,N_31122);
and U37827 (N_37827,N_33129,N_34934);
and U37828 (N_37828,N_30771,N_31565);
and U37829 (N_37829,N_31897,N_31217);
xnor U37830 (N_37830,N_31946,N_31860);
nand U37831 (N_37831,N_30668,N_32350);
nor U37832 (N_37832,N_30118,N_30653);
and U37833 (N_37833,N_30226,N_33698);
or U37834 (N_37834,N_33352,N_32506);
nor U37835 (N_37835,N_31368,N_30017);
and U37836 (N_37836,N_32245,N_31165);
xor U37837 (N_37837,N_34848,N_32039);
nor U37838 (N_37838,N_30015,N_31571);
nand U37839 (N_37839,N_31137,N_34310);
nor U37840 (N_37840,N_30275,N_34180);
or U37841 (N_37841,N_33172,N_34234);
xor U37842 (N_37842,N_34619,N_30585);
or U37843 (N_37843,N_31617,N_31453);
nor U37844 (N_37844,N_33941,N_31803);
xor U37845 (N_37845,N_34028,N_34103);
xnor U37846 (N_37846,N_31375,N_33082);
nand U37847 (N_37847,N_30697,N_31322);
nor U37848 (N_37848,N_30112,N_33019);
and U37849 (N_37849,N_32327,N_33108);
nor U37850 (N_37850,N_34417,N_34285);
and U37851 (N_37851,N_32714,N_34689);
or U37852 (N_37852,N_31649,N_32915);
and U37853 (N_37853,N_32773,N_33637);
nor U37854 (N_37854,N_32018,N_30453);
xnor U37855 (N_37855,N_32658,N_33942);
nand U37856 (N_37856,N_33797,N_33513);
nand U37857 (N_37857,N_30816,N_33147);
or U37858 (N_37858,N_34361,N_33414);
and U37859 (N_37859,N_30868,N_33610);
xor U37860 (N_37860,N_30669,N_32779);
nand U37861 (N_37861,N_30589,N_30734);
or U37862 (N_37862,N_31480,N_32623);
nand U37863 (N_37863,N_31778,N_33735);
and U37864 (N_37864,N_32055,N_31999);
xnor U37865 (N_37865,N_30878,N_31649);
xor U37866 (N_37866,N_33958,N_33576);
nor U37867 (N_37867,N_31611,N_30901);
xnor U37868 (N_37868,N_32351,N_32086);
and U37869 (N_37869,N_33456,N_33771);
or U37870 (N_37870,N_32422,N_31367);
nor U37871 (N_37871,N_31148,N_30028);
and U37872 (N_37872,N_31374,N_31759);
xnor U37873 (N_37873,N_33689,N_34209);
and U37874 (N_37874,N_32786,N_31513);
nor U37875 (N_37875,N_33056,N_32497);
xnor U37876 (N_37876,N_32806,N_32755);
nor U37877 (N_37877,N_34139,N_30861);
or U37878 (N_37878,N_30419,N_34293);
nand U37879 (N_37879,N_33766,N_30396);
or U37880 (N_37880,N_33887,N_32947);
nor U37881 (N_37881,N_34121,N_30448);
xnor U37882 (N_37882,N_34769,N_30648);
xnor U37883 (N_37883,N_30940,N_31478);
xnor U37884 (N_37884,N_34686,N_33093);
nand U37885 (N_37885,N_34677,N_32519);
or U37886 (N_37886,N_30922,N_31299);
xor U37887 (N_37887,N_31893,N_33445);
nand U37888 (N_37888,N_30741,N_34911);
xnor U37889 (N_37889,N_33579,N_33431);
xnor U37890 (N_37890,N_32594,N_34360);
and U37891 (N_37891,N_31735,N_32383);
nand U37892 (N_37892,N_33718,N_30366);
nor U37893 (N_37893,N_32621,N_31728);
and U37894 (N_37894,N_34308,N_33885);
and U37895 (N_37895,N_34393,N_31674);
nand U37896 (N_37896,N_33807,N_30918);
nor U37897 (N_37897,N_30355,N_32340);
and U37898 (N_37898,N_31926,N_31970);
or U37899 (N_37899,N_33444,N_34348);
nand U37900 (N_37900,N_34446,N_31879);
xor U37901 (N_37901,N_34181,N_34444);
and U37902 (N_37902,N_30221,N_33667);
and U37903 (N_37903,N_33228,N_30057);
and U37904 (N_37904,N_32538,N_34516);
xnor U37905 (N_37905,N_33208,N_31591);
or U37906 (N_37906,N_32673,N_33980);
xnor U37907 (N_37907,N_33029,N_31045);
xor U37908 (N_37908,N_30337,N_34025);
nor U37909 (N_37909,N_30759,N_33601);
and U37910 (N_37910,N_32529,N_33894);
nor U37911 (N_37911,N_32626,N_34674);
xor U37912 (N_37912,N_32924,N_34792);
nand U37913 (N_37913,N_30600,N_30501);
nor U37914 (N_37914,N_31073,N_30620);
and U37915 (N_37915,N_30716,N_30693);
nand U37916 (N_37916,N_31314,N_30343);
nor U37917 (N_37917,N_34944,N_34019);
xor U37918 (N_37918,N_30673,N_31731);
or U37919 (N_37919,N_32523,N_30380);
nand U37920 (N_37920,N_33873,N_32191);
or U37921 (N_37921,N_34983,N_30999);
nand U37922 (N_37922,N_32573,N_30005);
and U37923 (N_37923,N_33293,N_34141);
nand U37924 (N_37924,N_32748,N_33514);
xor U37925 (N_37925,N_34036,N_31131);
xor U37926 (N_37926,N_34208,N_31404);
nor U37927 (N_37927,N_31390,N_33120);
and U37928 (N_37928,N_30839,N_33370);
nor U37929 (N_37929,N_31439,N_31211);
nor U37930 (N_37930,N_31762,N_30346);
and U37931 (N_37931,N_30854,N_33712);
xnor U37932 (N_37932,N_32407,N_33523);
nor U37933 (N_37933,N_31858,N_30177);
xor U37934 (N_37934,N_34467,N_31807);
and U37935 (N_37935,N_34642,N_34344);
or U37936 (N_37936,N_32534,N_31796);
or U37937 (N_37937,N_32314,N_33268);
nand U37938 (N_37938,N_30681,N_31041);
xnor U37939 (N_37939,N_33413,N_31015);
nand U37940 (N_37940,N_34821,N_34773);
nor U37941 (N_37941,N_30037,N_32919);
nor U37942 (N_37942,N_31003,N_32349);
and U37943 (N_37943,N_31459,N_31308);
or U37944 (N_37944,N_34543,N_31877);
or U37945 (N_37945,N_32250,N_33245);
nor U37946 (N_37946,N_33678,N_31059);
nor U37947 (N_37947,N_31969,N_32264);
xnor U37948 (N_37948,N_34475,N_33037);
nor U37949 (N_37949,N_30255,N_32273);
xnor U37950 (N_37950,N_32894,N_32317);
nand U37951 (N_37951,N_30011,N_33895);
nor U37952 (N_37952,N_32693,N_31486);
nand U37953 (N_37953,N_33021,N_33407);
and U37954 (N_37954,N_31568,N_33464);
and U37955 (N_37955,N_34144,N_30188);
nand U37956 (N_37956,N_31816,N_32267);
xnor U37957 (N_37957,N_30475,N_30841);
nor U37958 (N_37958,N_33245,N_30995);
nand U37959 (N_37959,N_30401,N_32866);
nor U37960 (N_37960,N_31587,N_32544);
xnor U37961 (N_37961,N_34712,N_31563);
and U37962 (N_37962,N_34220,N_31843);
and U37963 (N_37963,N_32870,N_33886);
xnor U37964 (N_37964,N_33821,N_34448);
or U37965 (N_37965,N_33942,N_30466);
or U37966 (N_37966,N_32391,N_33373);
nor U37967 (N_37967,N_33810,N_34186);
and U37968 (N_37968,N_31951,N_34687);
nand U37969 (N_37969,N_31953,N_33856);
xor U37970 (N_37970,N_32608,N_34372);
xnor U37971 (N_37971,N_33198,N_32332);
xor U37972 (N_37972,N_30530,N_31122);
nand U37973 (N_37973,N_30007,N_33557);
or U37974 (N_37974,N_31905,N_33153);
xnor U37975 (N_37975,N_32502,N_34698);
or U37976 (N_37976,N_30435,N_34872);
nor U37977 (N_37977,N_31351,N_32359);
or U37978 (N_37978,N_30299,N_31260);
nand U37979 (N_37979,N_33985,N_33241);
nand U37980 (N_37980,N_33206,N_30567);
xor U37981 (N_37981,N_30533,N_31529);
and U37982 (N_37982,N_32136,N_33171);
xnor U37983 (N_37983,N_31795,N_34353);
xor U37984 (N_37984,N_34879,N_30136);
nand U37985 (N_37985,N_32981,N_34701);
or U37986 (N_37986,N_32092,N_33732);
and U37987 (N_37987,N_32847,N_30370);
nand U37988 (N_37988,N_31051,N_34128);
nor U37989 (N_37989,N_30307,N_34282);
xnor U37990 (N_37990,N_31391,N_34191);
nand U37991 (N_37991,N_34691,N_34750);
xor U37992 (N_37992,N_31441,N_32042);
nor U37993 (N_37993,N_33842,N_30444);
xor U37994 (N_37994,N_33748,N_32643);
nand U37995 (N_37995,N_31698,N_32559);
and U37996 (N_37996,N_33169,N_31829);
xnor U37997 (N_37997,N_30264,N_30141);
and U37998 (N_37998,N_34119,N_30122);
xor U37999 (N_37999,N_34963,N_32665);
or U38000 (N_38000,N_34052,N_31592);
xor U38001 (N_38001,N_34128,N_32562);
nor U38002 (N_38002,N_30854,N_34350);
or U38003 (N_38003,N_31683,N_34713);
nor U38004 (N_38004,N_32358,N_34615);
nand U38005 (N_38005,N_34623,N_31968);
xnor U38006 (N_38006,N_33091,N_33453);
or U38007 (N_38007,N_31764,N_33182);
nand U38008 (N_38008,N_30215,N_33506);
and U38009 (N_38009,N_34226,N_32069);
or U38010 (N_38010,N_30241,N_30655);
nand U38011 (N_38011,N_32325,N_30206);
and U38012 (N_38012,N_31266,N_31969);
and U38013 (N_38013,N_32672,N_31934);
xnor U38014 (N_38014,N_32661,N_33149);
and U38015 (N_38015,N_32861,N_33869);
nor U38016 (N_38016,N_32112,N_30072);
nand U38017 (N_38017,N_31211,N_33572);
nor U38018 (N_38018,N_31881,N_32979);
and U38019 (N_38019,N_31072,N_33779);
nor U38020 (N_38020,N_32919,N_33308);
xnor U38021 (N_38021,N_33958,N_34182);
xor U38022 (N_38022,N_30792,N_34267);
nor U38023 (N_38023,N_32787,N_31111);
nand U38024 (N_38024,N_34441,N_31802);
xor U38025 (N_38025,N_34714,N_34197);
nor U38026 (N_38026,N_30801,N_32764);
xor U38027 (N_38027,N_30750,N_30723);
xnor U38028 (N_38028,N_33787,N_32558);
xor U38029 (N_38029,N_32827,N_32341);
xor U38030 (N_38030,N_31868,N_33287);
nand U38031 (N_38031,N_31850,N_31982);
nand U38032 (N_38032,N_32378,N_32861);
nand U38033 (N_38033,N_33588,N_33841);
and U38034 (N_38034,N_30221,N_33693);
nand U38035 (N_38035,N_32344,N_32520);
and U38036 (N_38036,N_30622,N_32723);
xor U38037 (N_38037,N_30248,N_31948);
nand U38038 (N_38038,N_31017,N_32323);
nor U38039 (N_38039,N_33019,N_34763);
and U38040 (N_38040,N_34112,N_32513);
xor U38041 (N_38041,N_30294,N_33120);
and U38042 (N_38042,N_34220,N_34502);
and U38043 (N_38043,N_34791,N_32469);
or U38044 (N_38044,N_30095,N_33419);
and U38045 (N_38045,N_32495,N_30581);
and U38046 (N_38046,N_32794,N_34786);
nor U38047 (N_38047,N_31350,N_30415);
and U38048 (N_38048,N_33477,N_31656);
and U38049 (N_38049,N_32354,N_32795);
xnor U38050 (N_38050,N_32364,N_32811);
and U38051 (N_38051,N_32494,N_30780);
nor U38052 (N_38052,N_30760,N_33345);
nor U38053 (N_38053,N_31453,N_31384);
xor U38054 (N_38054,N_32333,N_31389);
nand U38055 (N_38055,N_34204,N_32341);
and U38056 (N_38056,N_30810,N_30491);
xor U38057 (N_38057,N_31141,N_31258);
nand U38058 (N_38058,N_32619,N_31390);
or U38059 (N_38059,N_31964,N_32654);
nand U38060 (N_38060,N_34696,N_33168);
or U38061 (N_38061,N_33884,N_32172);
nand U38062 (N_38062,N_30797,N_33074);
and U38063 (N_38063,N_30197,N_33454);
xnor U38064 (N_38064,N_33605,N_30940);
and U38065 (N_38065,N_31711,N_34709);
or U38066 (N_38066,N_31370,N_33631);
nor U38067 (N_38067,N_31580,N_32380);
and U38068 (N_38068,N_33535,N_32868);
or U38069 (N_38069,N_34268,N_32249);
nand U38070 (N_38070,N_32557,N_34286);
nand U38071 (N_38071,N_34815,N_32525);
and U38072 (N_38072,N_32089,N_34245);
nand U38073 (N_38073,N_34380,N_31503);
nor U38074 (N_38074,N_34298,N_32993);
xnor U38075 (N_38075,N_31753,N_34937);
nor U38076 (N_38076,N_33037,N_34162);
and U38077 (N_38077,N_33691,N_31471);
and U38078 (N_38078,N_34693,N_30456);
and U38079 (N_38079,N_34108,N_32945);
nand U38080 (N_38080,N_34070,N_33694);
or U38081 (N_38081,N_32865,N_33100);
xnor U38082 (N_38082,N_33067,N_34895);
and U38083 (N_38083,N_30059,N_34307);
and U38084 (N_38084,N_33911,N_34076);
nor U38085 (N_38085,N_34269,N_34368);
nand U38086 (N_38086,N_33251,N_33693);
xor U38087 (N_38087,N_32165,N_33312);
or U38088 (N_38088,N_34008,N_32458);
and U38089 (N_38089,N_30786,N_31623);
nand U38090 (N_38090,N_31166,N_31457);
and U38091 (N_38091,N_31206,N_34741);
or U38092 (N_38092,N_34193,N_32900);
and U38093 (N_38093,N_32694,N_30146);
xor U38094 (N_38094,N_33396,N_30117);
and U38095 (N_38095,N_34022,N_32109);
nand U38096 (N_38096,N_30672,N_33363);
nor U38097 (N_38097,N_32032,N_34187);
xnor U38098 (N_38098,N_31207,N_34792);
xnor U38099 (N_38099,N_32706,N_31085);
and U38100 (N_38100,N_33943,N_32220);
or U38101 (N_38101,N_32154,N_32822);
nor U38102 (N_38102,N_31303,N_34479);
or U38103 (N_38103,N_33409,N_32597);
xnor U38104 (N_38104,N_32416,N_32994);
xor U38105 (N_38105,N_32391,N_31084);
nand U38106 (N_38106,N_31289,N_31918);
nand U38107 (N_38107,N_30883,N_33786);
nor U38108 (N_38108,N_30347,N_32851);
xor U38109 (N_38109,N_34407,N_30215);
and U38110 (N_38110,N_33297,N_34398);
xnor U38111 (N_38111,N_30724,N_30234);
and U38112 (N_38112,N_34837,N_31445);
xnor U38113 (N_38113,N_32762,N_33296);
xor U38114 (N_38114,N_34478,N_31659);
and U38115 (N_38115,N_34618,N_32883);
and U38116 (N_38116,N_32375,N_31416);
nor U38117 (N_38117,N_32370,N_33753);
nor U38118 (N_38118,N_34783,N_31015);
and U38119 (N_38119,N_33790,N_33059);
and U38120 (N_38120,N_33446,N_33119);
nor U38121 (N_38121,N_31349,N_30464);
xnor U38122 (N_38122,N_30396,N_30843);
nor U38123 (N_38123,N_32666,N_31160);
and U38124 (N_38124,N_31646,N_30747);
or U38125 (N_38125,N_34488,N_32530);
nor U38126 (N_38126,N_30759,N_30007);
nor U38127 (N_38127,N_33643,N_32750);
or U38128 (N_38128,N_32723,N_32386);
nor U38129 (N_38129,N_30448,N_33416);
nor U38130 (N_38130,N_32780,N_32141);
xnor U38131 (N_38131,N_30212,N_34755);
and U38132 (N_38132,N_31227,N_34003);
nor U38133 (N_38133,N_31486,N_30385);
and U38134 (N_38134,N_33376,N_31575);
xor U38135 (N_38135,N_34081,N_33387);
nor U38136 (N_38136,N_30320,N_32564);
nand U38137 (N_38137,N_31957,N_34997);
xor U38138 (N_38138,N_31968,N_33589);
or U38139 (N_38139,N_32114,N_31055);
and U38140 (N_38140,N_34821,N_33972);
or U38141 (N_38141,N_30595,N_30226);
nor U38142 (N_38142,N_32451,N_31336);
xnor U38143 (N_38143,N_30220,N_32222);
xnor U38144 (N_38144,N_32461,N_32477);
nand U38145 (N_38145,N_32380,N_34032);
xnor U38146 (N_38146,N_32557,N_31796);
nand U38147 (N_38147,N_33176,N_34420);
xor U38148 (N_38148,N_32267,N_30098);
and U38149 (N_38149,N_32202,N_30013);
or U38150 (N_38150,N_34117,N_34926);
and U38151 (N_38151,N_34950,N_34236);
nor U38152 (N_38152,N_31591,N_32550);
or U38153 (N_38153,N_30882,N_30194);
nand U38154 (N_38154,N_31445,N_34431);
or U38155 (N_38155,N_31398,N_33700);
nor U38156 (N_38156,N_30602,N_31825);
and U38157 (N_38157,N_30324,N_33553);
nand U38158 (N_38158,N_31769,N_33685);
nand U38159 (N_38159,N_30077,N_34067);
nand U38160 (N_38160,N_32887,N_30409);
xnor U38161 (N_38161,N_31519,N_33339);
nand U38162 (N_38162,N_31964,N_32407);
xnor U38163 (N_38163,N_32125,N_34676);
and U38164 (N_38164,N_31864,N_34027);
xor U38165 (N_38165,N_34627,N_31173);
nor U38166 (N_38166,N_34417,N_30835);
or U38167 (N_38167,N_34510,N_30300);
or U38168 (N_38168,N_34922,N_30980);
xnor U38169 (N_38169,N_32757,N_32901);
and U38170 (N_38170,N_33132,N_31452);
xnor U38171 (N_38171,N_32999,N_32419);
nand U38172 (N_38172,N_31059,N_32115);
and U38173 (N_38173,N_32103,N_33518);
and U38174 (N_38174,N_32079,N_30496);
xnor U38175 (N_38175,N_31979,N_31359);
nor U38176 (N_38176,N_34690,N_31083);
and U38177 (N_38177,N_33148,N_32362);
nor U38178 (N_38178,N_33786,N_32041);
or U38179 (N_38179,N_33575,N_34947);
xor U38180 (N_38180,N_31916,N_34386);
nand U38181 (N_38181,N_34685,N_34825);
nor U38182 (N_38182,N_34593,N_33737);
nor U38183 (N_38183,N_34778,N_33493);
or U38184 (N_38184,N_34564,N_34185);
and U38185 (N_38185,N_32890,N_33853);
or U38186 (N_38186,N_32649,N_34480);
and U38187 (N_38187,N_30348,N_33499);
nand U38188 (N_38188,N_31913,N_31170);
nor U38189 (N_38189,N_34810,N_31711);
or U38190 (N_38190,N_33064,N_30959);
or U38191 (N_38191,N_34719,N_34238);
nor U38192 (N_38192,N_33415,N_31383);
nor U38193 (N_38193,N_32412,N_34934);
nand U38194 (N_38194,N_32011,N_31815);
and U38195 (N_38195,N_30691,N_33840);
nor U38196 (N_38196,N_32420,N_31588);
or U38197 (N_38197,N_31606,N_30374);
nor U38198 (N_38198,N_34716,N_31558);
nor U38199 (N_38199,N_31284,N_30330);
and U38200 (N_38200,N_30337,N_30738);
nand U38201 (N_38201,N_30310,N_32901);
or U38202 (N_38202,N_30952,N_30761);
xor U38203 (N_38203,N_30244,N_32230);
and U38204 (N_38204,N_32454,N_33253);
or U38205 (N_38205,N_32164,N_32021);
xor U38206 (N_38206,N_31912,N_31512);
and U38207 (N_38207,N_34547,N_33500);
xor U38208 (N_38208,N_33984,N_34099);
and U38209 (N_38209,N_32738,N_33669);
xor U38210 (N_38210,N_30700,N_34696);
or U38211 (N_38211,N_32036,N_33852);
or U38212 (N_38212,N_33957,N_32436);
and U38213 (N_38213,N_31541,N_30025);
xnor U38214 (N_38214,N_30767,N_30835);
and U38215 (N_38215,N_32982,N_33264);
nor U38216 (N_38216,N_31882,N_32014);
xnor U38217 (N_38217,N_33143,N_34035);
nor U38218 (N_38218,N_32957,N_31553);
and U38219 (N_38219,N_33223,N_32319);
xnor U38220 (N_38220,N_30077,N_34811);
nor U38221 (N_38221,N_30464,N_33427);
xnor U38222 (N_38222,N_34605,N_34049);
xor U38223 (N_38223,N_31619,N_32610);
nand U38224 (N_38224,N_33283,N_33906);
nor U38225 (N_38225,N_33931,N_33368);
xor U38226 (N_38226,N_30528,N_30874);
and U38227 (N_38227,N_30186,N_31072);
nand U38228 (N_38228,N_34907,N_30104);
and U38229 (N_38229,N_32473,N_30706);
nor U38230 (N_38230,N_33982,N_32800);
or U38231 (N_38231,N_34963,N_30425);
or U38232 (N_38232,N_30853,N_31616);
or U38233 (N_38233,N_32896,N_33657);
nand U38234 (N_38234,N_32515,N_34581);
nor U38235 (N_38235,N_30240,N_34934);
and U38236 (N_38236,N_31060,N_33192);
xnor U38237 (N_38237,N_33700,N_31847);
nor U38238 (N_38238,N_31014,N_34125);
xnor U38239 (N_38239,N_31368,N_30618);
xor U38240 (N_38240,N_32638,N_32086);
or U38241 (N_38241,N_33561,N_31950);
nor U38242 (N_38242,N_31098,N_30742);
and U38243 (N_38243,N_30302,N_33403);
and U38244 (N_38244,N_32188,N_34820);
nor U38245 (N_38245,N_33864,N_33168);
xnor U38246 (N_38246,N_34675,N_30703);
and U38247 (N_38247,N_33289,N_33233);
and U38248 (N_38248,N_34514,N_30957);
and U38249 (N_38249,N_31812,N_30835);
xnor U38250 (N_38250,N_34506,N_31938);
nand U38251 (N_38251,N_32336,N_32565);
and U38252 (N_38252,N_32227,N_32289);
and U38253 (N_38253,N_31668,N_33347);
nor U38254 (N_38254,N_31355,N_30141);
nand U38255 (N_38255,N_30000,N_34305);
nor U38256 (N_38256,N_30454,N_34268);
and U38257 (N_38257,N_34334,N_30255);
nor U38258 (N_38258,N_31436,N_33976);
xor U38259 (N_38259,N_30128,N_32134);
nand U38260 (N_38260,N_32091,N_31335);
and U38261 (N_38261,N_33414,N_32762);
and U38262 (N_38262,N_30319,N_31395);
xor U38263 (N_38263,N_33940,N_31742);
xor U38264 (N_38264,N_33451,N_33312);
and U38265 (N_38265,N_33299,N_30288);
and U38266 (N_38266,N_33838,N_33179);
nand U38267 (N_38267,N_31554,N_33452);
and U38268 (N_38268,N_30013,N_31101);
and U38269 (N_38269,N_33298,N_33386);
nor U38270 (N_38270,N_32324,N_31420);
nand U38271 (N_38271,N_31985,N_34807);
nand U38272 (N_38272,N_33882,N_34336);
nor U38273 (N_38273,N_30564,N_33789);
and U38274 (N_38274,N_31124,N_30193);
nor U38275 (N_38275,N_32433,N_32787);
and U38276 (N_38276,N_33446,N_31113);
or U38277 (N_38277,N_30963,N_33279);
nor U38278 (N_38278,N_33129,N_32956);
xnor U38279 (N_38279,N_30612,N_32740);
and U38280 (N_38280,N_32653,N_34772);
nor U38281 (N_38281,N_33625,N_30858);
nor U38282 (N_38282,N_30033,N_34413);
or U38283 (N_38283,N_34651,N_33409);
nor U38284 (N_38284,N_33827,N_31661);
xor U38285 (N_38285,N_34841,N_31841);
xnor U38286 (N_38286,N_31827,N_32840);
and U38287 (N_38287,N_33613,N_30582);
and U38288 (N_38288,N_30677,N_30999);
nor U38289 (N_38289,N_32427,N_31386);
or U38290 (N_38290,N_31826,N_33610);
or U38291 (N_38291,N_33812,N_34702);
xnor U38292 (N_38292,N_31073,N_34420);
nand U38293 (N_38293,N_31062,N_30368);
and U38294 (N_38294,N_32366,N_34237);
nand U38295 (N_38295,N_31173,N_31864);
nand U38296 (N_38296,N_34474,N_33945);
and U38297 (N_38297,N_34887,N_30937);
nor U38298 (N_38298,N_32372,N_31361);
nand U38299 (N_38299,N_32665,N_33502);
xnor U38300 (N_38300,N_33976,N_32483);
xnor U38301 (N_38301,N_33136,N_31155);
or U38302 (N_38302,N_31298,N_31251);
or U38303 (N_38303,N_34500,N_32059);
nand U38304 (N_38304,N_31126,N_34951);
nand U38305 (N_38305,N_31158,N_33559);
and U38306 (N_38306,N_31553,N_33367);
or U38307 (N_38307,N_30958,N_33491);
or U38308 (N_38308,N_34537,N_30163);
and U38309 (N_38309,N_32044,N_32440);
nor U38310 (N_38310,N_31668,N_34069);
xor U38311 (N_38311,N_33965,N_30452);
xor U38312 (N_38312,N_30494,N_33266);
xnor U38313 (N_38313,N_33299,N_34115);
nor U38314 (N_38314,N_33193,N_32766);
nand U38315 (N_38315,N_33661,N_33915);
nand U38316 (N_38316,N_34364,N_30409);
nor U38317 (N_38317,N_31662,N_30114);
xnor U38318 (N_38318,N_34933,N_34524);
and U38319 (N_38319,N_32254,N_33386);
nor U38320 (N_38320,N_34151,N_30601);
nand U38321 (N_38321,N_30816,N_32176);
and U38322 (N_38322,N_34655,N_32740);
xnor U38323 (N_38323,N_31606,N_30660);
xor U38324 (N_38324,N_32250,N_31225);
nand U38325 (N_38325,N_30963,N_32510);
and U38326 (N_38326,N_30562,N_33362);
xnor U38327 (N_38327,N_30621,N_30858);
nor U38328 (N_38328,N_30266,N_30898);
or U38329 (N_38329,N_33677,N_34049);
or U38330 (N_38330,N_30950,N_33209);
nor U38331 (N_38331,N_30209,N_34511);
and U38332 (N_38332,N_32384,N_30919);
and U38333 (N_38333,N_34425,N_32099);
xor U38334 (N_38334,N_33901,N_30230);
nand U38335 (N_38335,N_31105,N_31807);
or U38336 (N_38336,N_33327,N_31027);
nand U38337 (N_38337,N_30077,N_32190);
and U38338 (N_38338,N_33588,N_31756);
and U38339 (N_38339,N_31738,N_33249);
nor U38340 (N_38340,N_30345,N_31601);
or U38341 (N_38341,N_30848,N_30747);
xor U38342 (N_38342,N_32257,N_32447);
nand U38343 (N_38343,N_32725,N_32184);
and U38344 (N_38344,N_34906,N_30261);
nand U38345 (N_38345,N_33560,N_32624);
and U38346 (N_38346,N_31263,N_33696);
nand U38347 (N_38347,N_31021,N_32566);
or U38348 (N_38348,N_34028,N_30215);
nand U38349 (N_38349,N_32553,N_30187);
and U38350 (N_38350,N_33609,N_34708);
nand U38351 (N_38351,N_32538,N_34173);
nand U38352 (N_38352,N_31703,N_32253);
or U38353 (N_38353,N_34775,N_33346);
and U38354 (N_38354,N_31347,N_34230);
nand U38355 (N_38355,N_32015,N_32805);
or U38356 (N_38356,N_33863,N_30961);
nand U38357 (N_38357,N_33385,N_31469);
and U38358 (N_38358,N_34973,N_34246);
xor U38359 (N_38359,N_33279,N_34007);
nor U38360 (N_38360,N_30940,N_31567);
and U38361 (N_38361,N_33290,N_31931);
and U38362 (N_38362,N_32357,N_33751);
and U38363 (N_38363,N_31992,N_34271);
xor U38364 (N_38364,N_32048,N_34042);
and U38365 (N_38365,N_31150,N_30167);
nor U38366 (N_38366,N_34367,N_30111);
nor U38367 (N_38367,N_32170,N_30038);
nand U38368 (N_38368,N_33551,N_34483);
or U38369 (N_38369,N_34928,N_30989);
nand U38370 (N_38370,N_34776,N_31612);
and U38371 (N_38371,N_31500,N_31841);
xor U38372 (N_38372,N_34166,N_32590);
xor U38373 (N_38373,N_30843,N_30418);
xor U38374 (N_38374,N_30964,N_30012);
nand U38375 (N_38375,N_30255,N_30762);
xnor U38376 (N_38376,N_31373,N_33315);
nand U38377 (N_38377,N_34765,N_33681);
and U38378 (N_38378,N_30477,N_32529);
or U38379 (N_38379,N_33400,N_32391);
and U38380 (N_38380,N_30199,N_34816);
nor U38381 (N_38381,N_34922,N_34827);
nand U38382 (N_38382,N_34740,N_33582);
or U38383 (N_38383,N_33282,N_31865);
nor U38384 (N_38384,N_32803,N_32242);
nor U38385 (N_38385,N_33811,N_34754);
xnor U38386 (N_38386,N_31926,N_31715);
nand U38387 (N_38387,N_32844,N_30928);
nor U38388 (N_38388,N_31870,N_32587);
nor U38389 (N_38389,N_30875,N_31949);
nor U38390 (N_38390,N_34475,N_30707);
and U38391 (N_38391,N_32659,N_32907);
and U38392 (N_38392,N_34867,N_33882);
xnor U38393 (N_38393,N_34922,N_30107);
or U38394 (N_38394,N_34236,N_33362);
xor U38395 (N_38395,N_30943,N_34577);
or U38396 (N_38396,N_31359,N_31761);
xnor U38397 (N_38397,N_32747,N_34829);
or U38398 (N_38398,N_31644,N_30699);
nand U38399 (N_38399,N_33213,N_31542);
and U38400 (N_38400,N_34857,N_34730);
and U38401 (N_38401,N_31002,N_32230);
nor U38402 (N_38402,N_34447,N_32803);
or U38403 (N_38403,N_31571,N_30990);
nor U38404 (N_38404,N_31725,N_32663);
or U38405 (N_38405,N_33272,N_34273);
or U38406 (N_38406,N_34281,N_32587);
xor U38407 (N_38407,N_33867,N_34291);
nand U38408 (N_38408,N_32905,N_34582);
xor U38409 (N_38409,N_30965,N_31777);
or U38410 (N_38410,N_31164,N_33293);
xor U38411 (N_38411,N_32170,N_31524);
nor U38412 (N_38412,N_30782,N_31496);
xnor U38413 (N_38413,N_34810,N_30685);
or U38414 (N_38414,N_34879,N_32711);
or U38415 (N_38415,N_33175,N_34469);
nand U38416 (N_38416,N_32184,N_33920);
nor U38417 (N_38417,N_32921,N_31867);
nand U38418 (N_38418,N_32986,N_31913);
nor U38419 (N_38419,N_32536,N_32448);
and U38420 (N_38420,N_33179,N_34009);
and U38421 (N_38421,N_34231,N_34950);
nand U38422 (N_38422,N_31656,N_34832);
or U38423 (N_38423,N_34155,N_34817);
xor U38424 (N_38424,N_31009,N_32477);
and U38425 (N_38425,N_31670,N_34317);
nor U38426 (N_38426,N_30948,N_30013);
and U38427 (N_38427,N_33950,N_31759);
nand U38428 (N_38428,N_32173,N_34389);
or U38429 (N_38429,N_34063,N_34527);
nor U38430 (N_38430,N_31583,N_32968);
nor U38431 (N_38431,N_31971,N_30572);
nor U38432 (N_38432,N_31250,N_33274);
nor U38433 (N_38433,N_33713,N_30349);
nand U38434 (N_38434,N_33543,N_31563);
or U38435 (N_38435,N_33860,N_31505);
or U38436 (N_38436,N_34163,N_33810);
nand U38437 (N_38437,N_30605,N_30442);
xnor U38438 (N_38438,N_32049,N_32030);
and U38439 (N_38439,N_31125,N_33677);
and U38440 (N_38440,N_32725,N_32279);
and U38441 (N_38441,N_30347,N_34089);
or U38442 (N_38442,N_30633,N_33245);
or U38443 (N_38443,N_30555,N_30492);
or U38444 (N_38444,N_34605,N_34186);
xor U38445 (N_38445,N_31408,N_30315);
nor U38446 (N_38446,N_32578,N_30805);
nor U38447 (N_38447,N_30595,N_30945);
or U38448 (N_38448,N_31486,N_30831);
and U38449 (N_38449,N_30398,N_30453);
nand U38450 (N_38450,N_33830,N_34947);
or U38451 (N_38451,N_32743,N_31492);
nand U38452 (N_38452,N_32616,N_33254);
nand U38453 (N_38453,N_34374,N_30057);
or U38454 (N_38454,N_33378,N_32968);
and U38455 (N_38455,N_33967,N_34481);
xnor U38456 (N_38456,N_32048,N_32217);
nor U38457 (N_38457,N_32549,N_34028);
and U38458 (N_38458,N_30872,N_34682);
nand U38459 (N_38459,N_32311,N_31480);
and U38460 (N_38460,N_34536,N_32155);
xnor U38461 (N_38461,N_32307,N_34631);
and U38462 (N_38462,N_30202,N_30839);
nor U38463 (N_38463,N_34259,N_32384);
xnor U38464 (N_38464,N_32495,N_33601);
and U38465 (N_38465,N_30673,N_31453);
and U38466 (N_38466,N_31244,N_33856);
and U38467 (N_38467,N_30059,N_30155);
or U38468 (N_38468,N_33222,N_32732);
xor U38469 (N_38469,N_30772,N_30368);
nand U38470 (N_38470,N_33813,N_30764);
nor U38471 (N_38471,N_30082,N_30805);
xnor U38472 (N_38472,N_31878,N_34589);
nor U38473 (N_38473,N_31806,N_30887);
or U38474 (N_38474,N_30924,N_31157);
nand U38475 (N_38475,N_33154,N_30783);
nor U38476 (N_38476,N_34819,N_32203);
nand U38477 (N_38477,N_30845,N_32770);
or U38478 (N_38478,N_34466,N_30132);
and U38479 (N_38479,N_31245,N_31929);
xnor U38480 (N_38480,N_30079,N_31602);
nor U38481 (N_38481,N_31086,N_30618);
or U38482 (N_38482,N_33622,N_30842);
nor U38483 (N_38483,N_32294,N_30092);
xor U38484 (N_38484,N_33588,N_34047);
or U38485 (N_38485,N_30237,N_32589);
nand U38486 (N_38486,N_33219,N_34885);
nor U38487 (N_38487,N_31317,N_32448);
nand U38488 (N_38488,N_30213,N_34155);
nor U38489 (N_38489,N_33505,N_31875);
xnor U38490 (N_38490,N_31551,N_34897);
xor U38491 (N_38491,N_31894,N_34455);
nor U38492 (N_38492,N_32820,N_33526);
nor U38493 (N_38493,N_34198,N_31259);
xor U38494 (N_38494,N_31934,N_33824);
xnor U38495 (N_38495,N_33102,N_31666);
or U38496 (N_38496,N_34247,N_32326);
xnor U38497 (N_38497,N_34133,N_31306);
or U38498 (N_38498,N_30736,N_34163);
nor U38499 (N_38499,N_31120,N_34932);
xnor U38500 (N_38500,N_33221,N_34679);
nand U38501 (N_38501,N_30167,N_32103);
or U38502 (N_38502,N_34990,N_30840);
xor U38503 (N_38503,N_32237,N_33171);
xor U38504 (N_38504,N_33579,N_33937);
nor U38505 (N_38505,N_30874,N_33521);
and U38506 (N_38506,N_33917,N_31246);
nand U38507 (N_38507,N_31955,N_30857);
nor U38508 (N_38508,N_31465,N_30068);
or U38509 (N_38509,N_31778,N_31305);
xnor U38510 (N_38510,N_34122,N_32010);
nand U38511 (N_38511,N_32863,N_30801);
or U38512 (N_38512,N_32809,N_34823);
and U38513 (N_38513,N_31111,N_33405);
xor U38514 (N_38514,N_31757,N_30771);
or U38515 (N_38515,N_33102,N_32840);
nor U38516 (N_38516,N_31757,N_33392);
and U38517 (N_38517,N_32529,N_31939);
and U38518 (N_38518,N_31219,N_32578);
and U38519 (N_38519,N_32051,N_32731);
nor U38520 (N_38520,N_32687,N_30535);
and U38521 (N_38521,N_32213,N_33396);
or U38522 (N_38522,N_30014,N_33655);
xor U38523 (N_38523,N_32579,N_33973);
or U38524 (N_38524,N_31249,N_33471);
and U38525 (N_38525,N_31914,N_34693);
and U38526 (N_38526,N_33936,N_33444);
and U38527 (N_38527,N_30485,N_32847);
or U38528 (N_38528,N_34930,N_32540);
or U38529 (N_38529,N_33592,N_33602);
and U38530 (N_38530,N_30702,N_30818);
nor U38531 (N_38531,N_30603,N_34804);
or U38532 (N_38532,N_31021,N_31146);
xnor U38533 (N_38533,N_30137,N_30378);
nor U38534 (N_38534,N_32316,N_34775);
nand U38535 (N_38535,N_34630,N_34164);
nand U38536 (N_38536,N_33428,N_34161);
or U38537 (N_38537,N_34980,N_32684);
xnor U38538 (N_38538,N_33716,N_30173);
and U38539 (N_38539,N_33000,N_32169);
nor U38540 (N_38540,N_30417,N_31489);
and U38541 (N_38541,N_30054,N_34264);
nand U38542 (N_38542,N_34318,N_32391);
xor U38543 (N_38543,N_33654,N_34757);
and U38544 (N_38544,N_30272,N_32256);
or U38545 (N_38545,N_34838,N_31299);
xor U38546 (N_38546,N_34651,N_31086);
nor U38547 (N_38547,N_32819,N_34140);
and U38548 (N_38548,N_30554,N_31677);
nor U38549 (N_38549,N_34345,N_33067);
or U38550 (N_38550,N_32001,N_30693);
or U38551 (N_38551,N_31047,N_34728);
nor U38552 (N_38552,N_34281,N_33191);
and U38553 (N_38553,N_31147,N_30575);
nor U38554 (N_38554,N_34738,N_32262);
xor U38555 (N_38555,N_31031,N_32891);
and U38556 (N_38556,N_33480,N_31221);
xnor U38557 (N_38557,N_30448,N_33604);
xor U38558 (N_38558,N_34005,N_30795);
nand U38559 (N_38559,N_31020,N_34166);
xnor U38560 (N_38560,N_33786,N_34411);
xor U38561 (N_38561,N_34021,N_32085);
or U38562 (N_38562,N_33389,N_30460);
and U38563 (N_38563,N_30420,N_31795);
xor U38564 (N_38564,N_30102,N_33132);
and U38565 (N_38565,N_30889,N_34386);
xnor U38566 (N_38566,N_33813,N_34335);
nand U38567 (N_38567,N_32134,N_31105);
or U38568 (N_38568,N_30875,N_33287);
nand U38569 (N_38569,N_30610,N_34494);
xnor U38570 (N_38570,N_32860,N_30653);
xnor U38571 (N_38571,N_34576,N_30606);
nand U38572 (N_38572,N_33307,N_32378);
xnor U38573 (N_38573,N_33397,N_33422);
or U38574 (N_38574,N_30105,N_33563);
and U38575 (N_38575,N_30819,N_33853);
nand U38576 (N_38576,N_32675,N_34165);
nor U38577 (N_38577,N_31307,N_31766);
xnor U38578 (N_38578,N_31685,N_30608);
or U38579 (N_38579,N_30352,N_30357);
nand U38580 (N_38580,N_32450,N_34693);
or U38581 (N_38581,N_34296,N_32132);
xnor U38582 (N_38582,N_33050,N_34268);
or U38583 (N_38583,N_33432,N_34901);
or U38584 (N_38584,N_32878,N_30283);
or U38585 (N_38585,N_31548,N_34164);
or U38586 (N_38586,N_31553,N_32658);
or U38587 (N_38587,N_33325,N_34161);
or U38588 (N_38588,N_31612,N_33096);
xnor U38589 (N_38589,N_31254,N_34439);
and U38590 (N_38590,N_31417,N_34838);
nor U38591 (N_38591,N_33472,N_31331);
nor U38592 (N_38592,N_30576,N_34616);
nor U38593 (N_38593,N_31517,N_33338);
nand U38594 (N_38594,N_30899,N_30667);
nand U38595 (N_38595,N_34187,N_30361);
xnor U38596 (N_38596,N_32476,N_33821);
nand U38597 (N_38597,N_32509,N_33435);
xnor U38598 (N_38598,N_34199,N_31583);
or U38599 (N_38599,N_32090,N_34063);
and U38600 (N_38600,N_34599,N_32959);
nor U38601 (N_38601,N_34001,N_30493);
and U38602 (N_38602,N_32102,N_32885);
or U38603 (N_38603,N_34078,N_33662);
xnor U38604 (N_38604,N_30370,N_31345);
or U38605 (N_38605,N_30933,N_31357);
and U38606 (N_38606,N_32020,N_32952);
and U38607 (N_38607,N_34287,N_33409);
xor U38608 (N_38608,N_31060,N_30498);
xor U38609 (N_38609,N_32999,N_31125);
or U38610 (N_38610,N_32318,N_34829);
or U38611 (N_38611,N_34830,N_31627);
xnor U38612 (N_38612,N_34429,N_30804);
xor U38613 (N_38613,N_33124,N_34566);
nor U38614 (N_38614,N_30316,N_32112);
and U38615 (N_38615,N_33568,N_32467);
or U38616 (N_38616,N_32385,N_34940);
xor U38617 (N_38617,N_31624,N_34891);
nor U38618 (N_38618,N_34435,N_34984);
xnor U38619 (N_38619,N_30494,N_30397);
nand U38620 (N_38620,N_31045,N_34945);
and U38621 (N_38621,N_33995,N_31748);
xnor U38622 (N_38622,N_32700,N_32475);
or U38623 (N_38623,N_33280,N_31311);
and U38624 (N_38624,N_30855,N_30597);
xnor U38625 (N_38625,N_31342,N_30481);
nand U38626 (N_38626,N_30101,N_31609);
nand U38627 (N_38627,N_34308,N_30430);
or U38628 (N_38628,N_34478,N_30793);
and U38629 (N_38629,N_33678,N_33030);
xnor U38630 (N_38630,N_32756,N_32672);
xnor U38631 (N_38631,N_34312,N_34125);
nor U38632 (N_38632,N_32355,N_33887);
nand U38633 (N_38633,N_32458,N_31271);
or U38634 (N_38634,N_31392,N_30974);
nor U38635 (N_38635,N_30246,N_32745);
or U38636 (N_38636,N_34233,N_31068);
xor U38637 (N_38637,N_34364,N_30812);
or U38638 (N_38638,N_30786,N_30044);
or U38639 (N_38639,N_33758,N_30983);
nor U38640 (N_38640,N_33491,N_31904);
xor U38641 (N_38641,N_33043,N_30695);
and U38642 (N_38642,N_31595,N_32504);
nor U38643 (N_38643,N_31970,N_32723);
xor U38644 (N_38644,N_33117,N_31491);
or U38645 (N_38645,N_30632,N_32625);
or U38646 (N_38646,N_33998,N_33052);
or U38647 (N_38647,N_31681,N_31060);
or U38648 (N_38648,N_32833,N_34029);
and U38649 (N_38649,N_33567,N_30228);
nand U38650 (N_38650,N_33230,N_33011);
nor U38651 (N_38651,N_31366,N_32412);
xor U38652 (N_38652,N_32860,N_30056);
and U38653 (N_38653,N_32543,N_34442);
nor U38654 (N_38654,N_34648,N_30487);
and U38655 (N_38655,N_32690,N_33068);
nand U38656 (N_38656,N_34865,N_32439);
xnor U38657 (N_38657,N_32863,N_32574);
or U38658 (N_38658,N_34379,N_32319);
and U38659 (N_38659,N_30316,N_34796);
or U38660 (N_38660,N_34825,N_34518);
nor U38661 (N_38661,N_30588,N_31897);
xor U38662 (N_38662,N_33589,N_33967);
and U38663 (N_38663,N_34024,N_30141);
nand U38664 (N_38664,N_33295,N_32927);
and U38665 (N_38665,N_32605,N_33520);
xor U38666 (N_38666,N_32420,N_31538);
and U38667 (N_38667,N_34786,N_31132);
or U38668 (N_38668,N_31347,N_30684);
and U38669 (N_38669,N_34032,N_30836);
nor U38670 (N_38670,N_30341,N_31657);
or U38671 (N_38671,N_30728,N_34367);
nor U38672 (N_38672,N_32736,N_32152);
xor U38673 (N_38673,N_30544,N_33330);
or U38674 (N_38674,N_30920,N_30982);
xnor U38675 (N_38675,N_34661,N_34584);
nor U38676 (N_38676,N_30513,N_32924);
nor U38677 (N_38677,N_33618,N_33800);
xor U38678 (N_38678,N_31697,N_33930);
and U38679 (N_38679,N_34821,N_34103);
nor U38680 (N_38680,N_30310,N_32714);
or U38681 (N_38681,N_34703,N_32121);
nand U38682 (N_38682,N_30385,N_31965);
xor U38683 (N_38683,N_34996,N_32232);
xnor U38684 (N_38684,N_33766,N_34729);
xnor U38685 (N_38685,N_33494,N_34779);
nand U38686 (N_38686,N_32938,N_32510);
nand U38687 (N_38687,N_30658,N_34952);
nor U38688 (N_38688,N_32441,N_31581);
nor U38689 (N_38689,N_31652,N_30521);
xor U38690 (N_38690,N_33464,N_34581);
or U38691 (N_38691,N_32802,N_30010);
nor U38692 (N_38692,N_30209,N_31428);
xor U38693 (N_38693,N_33481,N_32308);
nor U38694 (N_38694,N_33654,N_33715);
or U38695 (N_38695,N_30950,N_32744);
and U38696 (N_38696,N_34645,N_32930);
nor U38697 (N_38697,N_30210,N_33219);
nor U38698 (N_38698,N_33400,N_34873);
nor U38699 (N_38699,N_31159,N_33027);
nand U38700 (N_38700,N_31978,N_31447);
nor U38701 (N_38701,N_31650,N_34378);
nor U38702 (N_38702,N_34813,N_30863);
or U38703 (N_38703,N_32832,N_34859);
or U38704 (N_38704,N_32366,N_32611);
and U38705 (N_38705,N_34465,N_32032);
and U38706 (N_38706,N_33820,N_30997);
or U38707 (N_38707,N_31684,N_31039);
xor U38708 (N_38708,N_31779,N_34153);
nand U38709 (N_38709,N_30367,N_30903);
or U38710 (N_38710,N_31162,N_30359);
nand U38711 (N_38711,N_33184,N_32973);
or U38712 (N_38712,N_32005,N_32283);
nand U38713 (N_38713,N_32706,N_32149);
nand U38714 (N_38714,N_30769,N_32194);
xnor U38715 (N_38715,N_34310,N_32358);
xnor U38716 (N_38716,N_34770,N_31014);
xor U38717 (N_38717,N_30316,N_34110);
xor U38718 (N_38718,N_31154,N_34752);
nor U38719 (N_38719,N_34261,N_30842);
and U38720 (N_38720,N_31463,N_33021);
nor U38721 (N_38721,N_31676,N_34233);
xnor U38722 (N_38722,N_33794,N_32550);
and U38723 (N_38723,N_31167,N_32184);
nand U38724 (N_38724,N_30696,N_31360);
and U38725 (N_38725,N_30546,N_33657);
nand U38726 (N_38726,N_32174,N_33120);
or U38727 (N_38727,N_31178,N_30908);
xnor U38728 (N_38728,N_31012,N_33161);
and U38729 (N_38729,N_34433,N_33375);
or U38730 (N_38730,N_32185,N_31448);
nor U38731 (N_38731,N_34843,N_30733);
nor U38732 (N_38732,N_34790,N_31232);
or U38733 (N_38733,N_31424,N_33853);
nor U38734 (N_38734,N_30751,N_34860);
xnor U38735 (N_38735,N_34965,N_34379);
or U38736 (N_38736,N_32362,N_31693);
or U38737 (N_38737,N_33555,N_31261);
nor U38738 (N_38738,N_34737,N_30808);
nand U38739 (N_38739,N_33842,N_30025);
xor U38740 (N_38740,N_34038,N_34545);
nand U38741 (N_38741,N_33308,N_34404);
or U38742 (N_38742,N_34947,N_30368);
xor U38743 (N_38743,N_30111,N_34685);
nand U38744 (N_38744,N_31421,N_30119);
or U38745 (N_38745,N_32888,N_31494);
xor U38746 (N_38746,N_30152,N_34341);
xor U38747 (N_38747,N_31223,N_34285);
nand U38748 (N_38748,N_34582,N_31239);
xnor U38749 (N_38749,N_30585,N_31524);
xnor U38750 (N_38750,N_31667,N_31012);
nand U38751 (N_38751,N_33077,N_34115);
nand U38752 (N_38752,N_32642,N_34584);
or U38753 (N_38753,N_33936,N_30198);
xor U38754 (N_38754,N_34155,N_32197);
nor U38755 (N_38755,N_33989,N_34496);
xnor U38756 (N_38756,N_30827,N_34630);
and U38757 (N_38757,N_34262,N_34279);
nand U38758 (N_38758,N_30872,N_31454);
nand U38759 (N_38759,N_34138,N_31554);
xnor U38760 (N_38760,N_34560,N_33322);
nand U38761 (N_38761,N_30625,N_30476);
nand U38762 (N_38762,N_32277,N_31367);
and U38763 (N_38763,N_32839,N_30505);
and U38764 (N_38764,N_30605,N_31396);
nor U38765 (N_38765,N_30845,N_32157);
nor U38766 (N_38766,N_33331,N_33426);
xnor U38767 (N_38767,N_30045,N_32899);
nor U38768 (N_38768,N_34621,N_32587);
and U38769 (N_38769,N_32745,N_34506);
xnor U38770 (N_38770,N_31612,N_34534);
or U38771 (N_38771,N_31043,N_31342);
nor U38772 (N_38772,N_31009,N_30850);
nor U38773 (N_38773,N_33636,N_33542);
nand U38774 (N_38774,N_31648,N_34849);
nand U38775 (N_38775,N_32722,N_34629);
and U38776 (N_38776,N_34782,N_31413);
and U38777 (N_38777,N_31998,N_32414);
nand U38778 (N_38778,N_31341,N_30032);
nor U38779 (N_38779,N_30617,N_33626);
and U38780 (N_38780,N_32766,N_32613);
and U38781 (N_38781,N_33749,N_31717);
xnor U38782 (N_38782,N_32132,N_31120);
and U38783 (N_38783,N_32192,N_32327);
nor U38784 (N_38784,N_33161,N_34251);
or U38785 (N_38785,N_30196,N_34132);
and U38786 (N_38786,N_33416,N_31507);
nand U38787 (N_38787,N_33167,N_33605);
or U38788 (N_38788,N_33330,N_32225);
nand U38789 (N_38789,N_34933,N_31193);
or U38790 (N_38790,N_34646,N_31286);
nor U38791 (N_38791,N_31215,N_30919);
nor U38792 (N_38792,N_32854,N_30720);
or U38793 (N_38793,N_32563,N_31864);
nand U38794 (N_38794,N_33160,N_34598);
nor U38795 (N_38795,N_33860,N_32072);
nor U38796 (N_38796,N_34689,N_33860);
or U38797 (N_38797,N_33345,N_32487);
nor U38798 (N_38798,N_33357,N_31410);
and U38799 (N_38799,N_31282,N_30206);
and U38800 (N_38800,N_34790,N_34234);
xor U38801 (N_38801,N_32737,N_31418);
xnor U38802 (N_38802,N_34250,N_34834);
or U38803 (N_38803,N_31508,N_33469);
xor U38804 (N_38804,N_34033,N_34434);
nor U38805 (N_38805,N_34015,N_33193);
nand U38806 (N_38806,N_30148,N_34274);
nand U38807 (N_38807,N_34086,N_34830);
nand U38808 (N_38808,N_33678,N_31871);
nor U38809 (N_38809,N_33404,N_32757);
nand U38810 (N_38810,N_32035,N_31412);
xnor U38811 (N_38811,N_30551,N_34727);
xor U38812 (N_38812,N_31317,N_31401);
xnor U38813 (N_38813,N_33378,N_34137);
nand U38814 (N_38814,N_31029,N_32143);
and U38815 (N_38815,N_34013,N_30409);
nand U38816 (N_38816,N_34245,N_33332);
xor U38817 (N_38817,N_32980,N_33502);
or U38818 (N_38818,N_33681,N_30053);
nand U38819 (N_38819,N_30240,N_30053);
nand U38820 (N_38820,N_33693,N_30313);
nor U38821 (N_38821,N_31756,N_33799);
nor U38822 (N_38822,N_30343,N_34309);
nor U38823 (N_38823,N_30512,N_30052);
nand U38824 (N_38824,N_33359,N_32804);
nand U38825 (N_38825,N_30074,N_32752);
xnor U38826 (N_38826,N_33859,N_31172);
xor U38827 (N_38827,N_31913,N_30570);
nor U38828 (N_38828,N_31439,N_32059);
and U38829 (N_38829,N_31663,N_30848);
xnor U38830 (N_38830,N_33267,N_34964);
nor U38831 (N_38831,N_30629,N_32721);
xnor U38832 (N_38832,N_31969,N_33402);
xnor U38833 (N_38833,N_32640,N_31504);
nor U38834 (N_38834,N_33397,N_31340);
and U38835 (N_38835,N_32858,N_34129);
nor U38836 (N_38836,N_34911,N_30967);
and U38837 (N_38837,N_34358,N_31766);
xnor U38838 (N_38838,N_32774,N_34135);
or U38839 (N_38839,N_30569,N_32999);
nand U38840 (N_38840,N_32785,N_33817);
and U38841 (N_38841,N_32106,N_32973);
xor U38842 (N_38842,N_34633,N_30297);
xnor U38843 (N_38843,N_32638,N_32347);
or U38844 (N_38844,N_31333,N_30343);
nor U38845 (N_38845,N_30312,N_33296);
or U38846 (N_38846,N_31329,N_33606);
or U38847 (N_38847,N_32838,N_33637);
xnor U38848 (N_38848,N_30270,N_30833);
nor U38849 (N_38849,N_32644,N_33241);
and U38850 (N_38850,N_31322,N_30017);
nor U38851 (N_38851,N_33808,N_30774);
and U38852 (N_38852,N_34531,N_33957);
xor U38853 (N_38853,N_31933,N_30758);
nor U38854 (N_38854,N_30750,N_34591);
nor U38855 (N_38855,N_31484,N_32989);
or U38856 (N_38856,N_30005,N_33102);
xnor U38857 (N_38857,N_32347,N_32940);
nor U38858 (N_38858,N_31367,N_34998);
and U38859 (N_38859,N_30794,N_30036);
or U38860 (N_38860,N_32810,N_32744);
nand U38861 (N_38861,N_33761,N_33841);
or U38862 (N_38862,N_33948,N_31416);
or U38863 (N_38863,N_30607,N_32211);
and U38864 (N_38864,N_31496,N_31124);
nor U38865 (N_38865,N_34331,N_30536);
nor U38866 (N_38866,N_30397,N_34746);
or U38867 (N_38867,N_31322,N_33754);
nand U38868 (N_38868,N_33556,N_34496);
or U38869 (N_38869,N_32651,N_32969);
nor U38870 (N_38870,N_30465,N_33047);
xnor U38871 (N_38871,N_33259,N_31123);
xor U38872 (N_38872,N_30994,N_30440);
or U38873 (N_38873,N_33636,N_31815);
xnor U38874 (N_38874,N_33193,N_34994);
and U38875 (N_38875,N_32599,N_33077);
xnor U38876 (N_38876,N_32075,N_32231);
nor U38877 (N_38877,N_33295,N_31597);
nand U38878 (N_38878,N_34528,N_30804);
nor U38879 (N_38879,N_33418,N_34001);
or U38880 (N_38880,N_33085,N_34308);
nor U38881 (N_38881,N_33641,N_33851);
xnor U38882 (N_38882,N_31284,N_30550);
xnor U38883 (N_38883,N_31369,N_34781);
nand U38884 (N_38884,N_33315,N_30234);
or U38885 (N_38885,N_34696,N_31870);
and U38886 (N_38886,N_33784,N_34879);
nand U38887 (N_38887,N_34938,N_30403);
xor U38888 (N_38888,N_32587,N_31903);
or U38889 (N_38889,N_33433,N_34151);
or U38890 (N_38890,N_34974,N_32668);
nor U38891 (N_38891,N_32334,N_34946);
or U38892 (N_38892,N_33951,N_31350);
or U38893 (N_38893,N_31927,N_33940);
nor U38894 (N_38894,N_32900,N_32279);
nand U38895 (N_38895,N_31281,N_32140);
nand U38896 (N_38896,N_33486,N_32044);
and U38897 (N_38897,N_30982,N_34336);
nor U38898 (N_38898,N_30475,N_30913);
nor U38899 (N_38899,N_33325,N_32693);
nor U38900 (N_38900,N_32313,N_34126);
xor U38901 (N_38901,N_31787,N_31204);
nor U38902 (N_38902,N_30816,N_34664);
nor U38903 (N_38903,N_34697,N_30926);
xor U38904 (N_38904,N_30921,N_32983);
and U38905 (N_38905,N_34844,N_33443);
or U38906 (N_38906,N_33792,N_30348);
xnor U38907 (N_38907,N_34151,N_31069);
or U38908 (N_38908,N_30767,N_31326);
xor U38909 (N_38909,N_33923,N_33238);
and U38910 (N_38910,N_32695,N_32920);
and U38911 (N_38911,N_32282,N_30059);
nor U38912 (N_38912,N_30047,N_32396);
nand U38913 (N_38913,N_34031,N_31979);
xor U38914 (N_38914,N_33674,N_34983);
or U38915 (N_38915,N_33562,N_31045);
nand U38916 (N_38916,N_32967,N_33626);
xor U38917 (N_38917,N_31090,N_33946);
nand U38918 (N_38918,N_33017,N_33021);
nand U38919 (N_38919,N_31837,N_31989);
or U38920 (N_38920,N_31415,N_34181);
nand U38921 (N_38921,N_34861,N_33343);
nand U38922 (N_38922,N_31798,N_30546);
or U38923 (N_38923,N_32882,N_32282);
nand U38924 (N_38924,N_34895,N_30422);
nor U38925 (N_38925,N_31479,N_34412);
nor U38926 (N_38926,N_31763,N_32189);
xnor U38927 (N_38927,N_32263,N_31840);
nand U38928 (N_38928,N_33309,N_32148);
or U38929 (N_38929,N_34013,N_34381);
nor U38930 (N_38930,N_30144,N_34931);
and U38931 (N_38931,N_33059,N_30114);
or U38932 (N_38932,N_30917,N_30593);
xor U38933 (N_38933,N_32781,N_34097);
and U38934 (N_38934,N_30057,N_31170);
and U38935 (N_38935,N_33010,N_34342);
xor U38936 (N_38936,N_32752,N_32040);
nor U38937 (N_38937,N_31202,N_31061);
and U38938 (N_38938,N_32391,N_34996);
xnor U38939 (N_38939,N_31881,N_32300);
or U38940 (N_38940,N_31820,N_32377);
or U38941 (N_38941,N_33402,N_30492);
nor U38942 (N_38942,N_34556,N_34318);
xnor U38943 (N_38943,N_31539,N_30975);
or U38944 (N_38944,N_31875,N_31761);
nand U38945 (N_38945,N_31783,N_34861);
nand U38946 (N_38946,N_30338,N_33324);
or U38947 (N_38947,N_33461,N_32707);
or U38948 (N_38948,N_33156,N_30586);
or U38949 (N_38949,N_30406,N_30627);
and U38950 (N_38950,N_33036,N_31983);
or U38951 (N_38951,N_31748,N_33668);
nor U38952 (N_38952,N_32048,N_34692);
and U38953 (N_38953,N_34592,N_31930);
nand U38954 (N_38954,N_33487,N_34479);
and U38955 (N_38955,N_33674,N_30422);
and U38956 (N_38956,N_33090,N_31232);
and U38957 (N_38957,N_31777,N_30570);
nand U38958 (N_38958,N_30068,N_33326);
xnor U38959 (N_38959,N_32772,N_31291);
xor U38960 (N_38960,N_33906,N_31315);
and U38961 (N_38961,N_34608,N_31361);
xnor U38962 (N_38962,N_30434,N_32404);
nor U38963 (N_38963,N_32650,N_33040);
nand U38964 (N_38964,N_32446,N_31013);
and U38965 (N_38965,N_30445,N_30263);
nor U38966 (N_38966,N_30803,N_34362);
or U38967 (N_38967,N_33692,N_31762);
nand U38968 (N_38968,N_34536,N_32507);
nor U38969 (N_38969,N_31004,N_31080);
xor U38970 (N_38970,N_30908,N_31251);
xor U38971 (N_38971,N_32439,N_34095);
nand U38972 (N_38972,N_31865,N_30257);
nand U38973 (N_38973,N_34716,N_34613);
nor U38974 (N_38974,N_34384,N_33177);
nor U38975 (N_38975,N_32096,N_31338);
nor U38976 (N_38976,N_31317,N_31414);
or U38977 (N_38977,N_30094,N_34525);
or U38978 (N_38978,N_34377,N_31374);
nand U38979 (N_38979,N_34224,N_33091);
and U38980 (N_38980,N_32538,N_32270);
and U38981 (N_38981,N_31563,N_33426);
nor U38982 (N_38982,N_33347,N_33844);
or U38983 (N_38983,N_34412,N_32586);
nand U38984 (N_38984,N_34320,N_33484);
xor U38985 (N_38985,N_33501,N_30329);
xor U38986 (N_38986,N_34778,N_34527);
nand U38987 (N_38987,N_30120,N_34632);
nand U38988 (N_38988,N_31552,N_31134);
and U38989 (N_38989,N_33278,N_30168);
nand U38990 (N_38990,N_34016,N_30154);
nand U38991 (N_38991,N_30032,N_30372);
nor U38992 (N_38992,N_33053,N_31394);
and U38993 (N_38993,N_33575,N_30270);
nand U38994 (N_38994,N_33582,N_34275);
xnor U38995 (N_38995,N_32062,N_32253);
or U38996 (N_38996,N_30479,N_30836);
or U38997 (N_38997,N_31976,N_34228);
or U38998 (N_38998,N_32803,N_34827);
or U38999 (N_38999,N_34724,N_33984);
or U39000 (N_39000,N_30384,N_31893);
xnor U39001 (N_39001,N_34291,N_34681);
xor U39002 (N_39002,N_34306,N_33463);
xor U39003 (N_39003,N_32228,N_31897);
or U39004 (N_39004,N_31750,N_30339);
nand U39005 (N_39005,N_31331,N_32266);
nor U39006 (N_39006,N_31876,N_33522);
xor U39007 (N_39007,N_30832,N_34652);
nand U39008 (N_39008,N_33173,N_31017);
nor U39009 (N_39009,N_32759,N_32924);
or U39010 (N_39010,N_31717,N_33327);
or U39011 (N_39011,N_31489,N_32444);
nand U39012 (N_39012,N_32471,N_31564);
nand U39013 (N_39013,N_32763,N_34252);
nor U39014 (N_39014,N_30116,N_30486);
xor U39015 (N_39015,N_33157,N_31897);
nand U39016 (N_39016,N_32689,N_32114);
or U39017 (N_39017,N_34565,N_33947);
nand U39018 (N_39018,N_34100,N_33423);
nor U39019 (N_39019,N_32908,N_33780);
and U39020 (N_39020,N_34523,N_33600);
xor U39021 (N_39021,N_32594,N_33660);
nand U39022 (N_39022,N_33341,N_30752);
nand U39023 (N_39023,N_32620,N_30680);
and U39024 (N_39024,N_32218,N_33467);
nand U39025 (N_39025,N_33086,N_30336);
and U39026 (N_39026,N_32885,N_34117);
xnor U39027 (N_39027,N_34184,N_32643);
or U39028 (N_39028,N_33361,N_30592);
and U39029 (N_39029,N_32832,N_30653);
and U39030 (N_39030,N_33439,N_31747);
nand U39031 (N_39031,N_32808,N_31483);
xor U39032 (N_39032,N_34540,N_30880);
nor U39033 (N_39033,N_32246,N_30223);
or U39034 (N_39034,N_34235,N_33319);
nand U39035 (N_39035,N_31321,N_30981);
and U39036 (N_39036,N_31121,N_32940);
and U39037 (N_39037,N_30000,N_30333);
and U39038 (N_39038,N_31998,N_33125);
nand U39039 (N_39039,N_31715,N_32762);
nand U39040 (N_39040,N_30386,N_34475);
and U39041 (N_39041,N_32882,N_32800);
nand U39042 (N_39042,N_32028,N_30893);
or U39043 (N_39043,N_34768,N_33325);
xnor U39044 (N_39044,N_32289,N_33256);
or U39045 (N_39045,N_34178,N_33798);
xnor U39046 (N_39046,N_32604,N_30592);
xnor U39047 (N_39047,N_31182,N_31649);
or U39048 (N_39048,N_31655,N_32142);
nor U39049 (N_39049,N_34906,N_33489);
nor U39050 (N_39050,N_30611,N_34181);
nand U39051 (N_39051,N_32974,N_30958);
xor U39052 (N_39052,N_30375,N_31096);
nand U39053 (N_39053,N_32325,N_33420);
nand U39054 (N_39054,N_32735,N_34087);
xnor U39055 (N_39055,N_34428,N_32138);
nand U39056 (N_39056,N_34075,N_31861);
and U39057 (N_39057,N_32661,N_33848);
nor U39058 (N_39058,N_32363,N_31475);
nand U39059 (N_39059,N_34995,N_32864);
nand U39060 (N_39060,N_32272,N_31187);
or U39061 (N_39061,N_31453,N_31510);
and U39062 (N_39062,N_30018,N_33274);
nand U39063 (N_39063,N_34447,N_33017);
and U39064 (N_39064,N_34092,N_31150);
xnor U39065 (N_39065,N_33432,N_30985);
and U39066 (N_39066,N_32280,N_31369);
and U39067 (N_39067,N_33796,N_34996);
and U39068 (N_39068,N_32324,N_31124);
xor U39069 (N_39069,N_32626,N_30104);
or U39070 (N_39070,N_33713,N_30049);
nor U39071 (N_39071,N_32197,N_32724);
and U39072 (N_39072,N_31913,N_32764);
nand U39073 (N_39073,N_33074,N_32999);
or U39074 (N_39074,N_31625,N_31496);
or U39075 (N_39075,N_31650,N_31206);
nor U39076 (N_39076,N_31761,N_32631);
or U39077 (N_39077,N_34257,N_33783);
nor U39078 (N_39078,N_30761,N_32213);
or U39079 (N_39079,N_31385,N_30095);
and U39080 (N_39080,N_32634,N_32080);
xor U39081 (N_39081,N_30513,N_31334);
and U39082 (N_39082,N_31648,N_32131);
and U39083 (N_39083,N_30894,N_30981);
nand U39084 (N_39084,N_30584,N_34561);
xor U39085 (N_39085,N_33333,N_31591);
nand U39086 (N_39086,N_31577,N_30968);
nor U39087 (N_39087,N_34533,N_31815);
xnor U39088 (N_39088,N_30805,N_33231);
or U39089 (N_39089,N_32361,N_34636);
or U39090 (N_39090,N_30386,N_30965);
and U39091 (N_39091,N_31810,N_32850);
xor U39092 (N_39092,N_31938,N_31057);
or U39093 (N_39093,N_30215,N_33843);
nand U39094 (N_39094,N_34168,N_32899);
and U39095 (N_39095,N_32285,N_33807);
or U39096 (N_39096,N_32606,N_33585);
nand U39097 (N_39097,N_32023,N_32326);
and U39098 (N_39098,N_33969,N_30018);
nor U39099 (N_39099,N_31544,N_33955);
and U39100 (N_39100,N_33223,N_32941);
xnor U39101 (N_39101,N_31656,N_33067);
and U39102 (N_39102,N_32254,N_31042);
nor U39103 (N_39103,N_32032,N_31716);
nor U39104 (N_39104,N_30738,N_32165);
xor U39105 (N_39105,N_34306,N_32769);
or U39106 (N_39106,N_30427,N_34884);
or U39107 (N_39107,N_32254,N_32401);
and U39108 (N_39108,N_31799,N_34154);
nor U39109 (N_39109,N_30521,N_34718);
xnor U39110 (N_39110,N_34209,N_30226);
nor U39111 (N_39111,N_32951,N_30887);
nor U39112 (N_39112,N_32554,N_32818);
xnor U39113 (N_39113,N_34246,N_31590);
or U39114 (N_39114,N_32819,N_33801);
nand U39115 (N_39115,N_33849,N_32794);
nand U39116 (N_39116,N_31462,N_31180);
nor U39117 (N_39117,N_31568,N_31468);
and U39118 (N_39118,N_33301,N_32576);
or U39119 (N_39119,N_33495,N_30449);
and U39120 (N_39120,N_31005,N_34727);
or U39121 (N_39121,N_33918,N_31205);
xor U39122 (N_39122,N_33866,N_34575);
nand U39123 (N_39123,N_31798,N_31657);
nand U39124 (N_39124,N_33052,N_31513);
or U39125 (N_39125,N_30310,N_34959);
nor U39126 (N_39126,N_32970,N_32682);
and U39127 (N_39127,N_30533,N_33975);
xor U39128 (N_39128,N_30726,N_32799);
nand U39129 (N_39129,N_33956,N_31734);
nor U39130 (N_39130,N_31470,N_33681);
nand U39131 (N_39131,N_34300,N_31614);
nand U39132 (N_39132,N_34420,N_32225);
and U39133 (N_39133,N_31307,N_30348);
nand U39134 (N_39134,N_31435,N_33803);
nand U39135 (N_39135,N_31388,N_30951);
or U39136 (N_39136,N_31451,N_33996);
nor U39137 (N_39137,N_30994,N_32338);
nand U39138 (N_39138,N_32742,N_33543);
and U39139 (N_39139,N_33364,N_32415);
nand U39140 (N_39140,N_30415,N_32984);
nor U39141 (N_39141,N_30389,N_30310);
or U39142 (N_39142,N_31046,N_30001);
nor U39143 (N_39143,N_32437,N_34603);
nand U39144 (N_39144,N_30478,N_31660);
nand U39145 (N_39145,N_32339,N_30257);
or U39146 (N_39146,N_30459,N_33304);
nand U39147 (N_39147,N_30459,N_33851);
and U39148 (N_39148,N_33318,N_33600);
or U39149 (N_39149,N_33395,N_30349);
and U39150 (N_39150,N_31133,N_32083);
xnor U39151 (N_39151,N_33586,N_32580);
and U39152 (N_39152,N_33986,N_33365);
nor U39153 (N_39153,N_32242,N_31174);
nand U39154 (N_39154,N_34336,N_31104);
or U39155 (N_39155,N_33254,N_32652);
nor U39156 (N_39156,N_31230,N_34834);
nand U39157 (N_39157,N_31663,N_34167);
or U39158 (N_39158,N_30929,N_31765);
nor U39159 (N_39159,N_31709,N_31838);
and U39160 (N_39160,N_34634,N_30613);
nor U39161 (N_39161,N_32752,N_33872);
or U39162 (N_39162,N_33113,N_33130);
nor U39163 (N_39163,N_30009,N_34991);
or U39164 (N_39164,N_33831,N_34592);
and U39165 (N_39165,N_33628,N_34380);
xnor U39166 (N_39166,N_34518,N_33711);
nor U39167 (N_39167,N_34105,N_34242);
nand U39168 (N_39168,N_32248,N_32290);
xor U39169 (N_39169,N_33548,N_32571);
xnor U39170 (N_39170,N_34491,N_32155);
xnor U39171 (N_39171,N_32002,N_34111);
and U39172 (N_39172,N_31322,N_33204);
nor U39173 (N_39173,N_34232,N_31789);
and U39174 (N_39174,N_33958,N_30040);
nand U39175 (N_39175,N_34161,N_32355);
xnor U39176 (N_39176,N_32087,N_32874);
and U39177 (N_39177,N_33367,N_34352);
and U39178 (N_39178,N_33983,N_30976);
xnor U39179 (N_39179,N_34521,N_31039);
nor U39180 (N_39180,N_32178,N_34829);
nor U39181 (N_39181,N_33763,N_32002);
xor U39182 (N_39182,N_32086,N_32936);
nor U39183 (N_39183,N_33358,N_34026);
nor U39184 (N_39184,N_30184,N_34988);
and U39185 (N_39185,N_33271,N_34935);
xor U39186 (N_39186,N_34192,N_30090);
nor U39187 (N_39187,N_31754,N_34034);
or U39188 (N_39188,N_32281,N_32618);
xnor U39189 (N_39189,N_31125,N_30835);
nand U39190 (N_39190,N_33398,N_31327);
and U39191 (N_39191,N_30867,N_33139);
nor U39192 (N_39192,N_30915,N_33420);
nor U39193 (N_39193,N_33465,N_30174);
and U39194 (N_39194,N_33047,N_34656);
xnor U39195 (N_39195,N_32706,N_34282);
or U39196 (N_39196,N_31686,N_33294);
nor U39197 (N_39197,N_34365,N_33302);
or U39198 (N_39198,N_33864,N_30137);
xnor U39199 (N_39199,N_34477,N_30444);
or U39200 (N_39200,N_33605,N_34216);
or U39201 (N_39201,N_31237,N_33515);
or U39202 (N_39202,N_34221,N_31437);
xor U39203 (N_39203,N_33755,N_32973);
nor U39204 (N_39204,N_32131,N_30429);
nand U39205 (N_39205,N_33515,N_31154);
nor U39206 (N_39206,N_34575,N_32431);
nor U39207 (N_39207,N_32011,N_31468);
nand U39208 (N_39208,N_31466,N_32080);
nor U39209 (N_39209,N_34122,N_32218);
nand U39210 (N_39210,N_34152,N_31132);
xor U39211 (N_39211,N_30156,N_34349);
xor U39212 (N_39212,N_31487,N_34794);
and U39213 (N_39213,N_32344,N_32499);
nand U39214 (N_39214,N_30699,N_31956);
or U39215 (N_39215,N_33786,N_34011);
and U39216 (N_39216,N_34635,N_34029);
nor U39217 (N_39217,N_32442,N_33948);
xor U39218 (N_39218,N_30175,N_32548);
nand U39219 (N_39219,N_31582,N_32721);
nand U39220 (N_39220,N_30802,N_34774);
nor U39221 (N_39221,N_32299,N_30564);
nor U39222 (N_39222,N_32010,N_33002);
nor U39223 (N_39223,N_31703,N_31265);
xor U39224 (N_39224,N_32613,N_30963);
nand U39225 (N_39225,N_30862,N_32075);
xor U39226 (N_39226,N_33660,N_30307);
nand U39227 (N_39227,N_31289,N_34084);
xnor U39228 (N_39228,N_30237,N_33697);
nor U39229 (N_39229,N_32060,N_32160);
nand U39230 (N_39230,N_32272,N_34703);
nand U39231 (N_39231,N_32246,N_34336);
or U39232 (N_39232,N_31297,N_32172);
or U39233 (N_39233,N_30168,N_32547);
nor U39234 (N_39234,N_30650,N_33297);
xor U39235 (N_39235,N_33488,N_33614);
nor U39236 (N_39236,N_31484,N_30332);
or U39237 (N_39237,N_33580,N_31622);
or U39238 (N_39238,N_30941,N_34033);
or U39239 (N_39239,N_33826,N_34898);
nor U39240 (N_39240,N_31414,N_30734);
xor U39241 (N_39241,N_32008,N_34232);
xor U39242 (N_39242,N_31528,N_32204);
nor U39243 (N_39243,N_30592,N_33586);
and U39244 (N_39244,N_34852,N_34948);
nand U39245 (N_39245,N_34056,N_34215);
nor U39246 (N_39246,N_34319,N_30188);
or U39247 (N_39247,N_33232,N_30290);
or U39248 (N_39248,N_31095,N_32994);
nor U39249 (N_39249,N_30602,N_30606);
and U39250 (N_39250,N_31286,N_33375);
or U39251 (N_39251,N_30999,N_32015);
or U39252 (N_39252,N_33091,N_32149);
nor U39253 (N_39253,N_31881,N_31096);
nand U39254 (N_39254,N_31264,N_33823);
and U39255 (N_39255,N_31626,N_32167);
or U39256 (N_39256,N_34142,N_34592);
xnor U39257 (N_39257,N_32506,N_32208);
and U39258 (N_39258,N_34987,N_30562);
xnor U39259 (N_39259,N_32894,N_32039);
xnor U39260 (N_39260,N_31230,N_32288);
and U39261 (N_39261,N_30140,N_32619);
nor U39262 (N_39262,N_32614,N_31134);
and U39263 (N_39263,N_34556,N_30096);
or U39264 (N_39264,N_31853,N_34017);
or U39265 (N_39265,N_32953,N_33374);
xnor U39266 (N_39266,N_33163,N_31271);
nand U39267 (N_39267,N_32468,N_33458);
and U39268 (N_39268,N_31408,N_31510);
and U39269 (N_39269,N_33138,N_34162);
nand U39270 (N_39270,N_31283,N_30883);
and U39271 (N_39271,N_34064,N_32556);
or U39272 (N_39272,N_33841,N_33820);
nand U39273 (N_39273,N_33740,N_30202);
nand U39274 (N_39274,N_32377,N_32901);
xor U39275 (N_39275,N_32033,N_30802);
and U39276 (N_39276,N_32459,N_34413);
xor U39277 (N_39277,N_31446,N_32411);
and U39278 (N_39278,N_32960,N_31709);
nand U39279 (N_39279,N_31852,N_34272);
nor U39280 (N_39280,N_33027,N_31734);
nand U39281 (N_39281,N_33699,N_30498);
xnor U39282 (N_39282,N_30129,N_31746);
nand U39283 (N_39283,N_31611,N_34992);
or U39284 (N_39284,N_32086,N_31034);
xnor U39285 (N_39285,N_34139,N_34882);
xor U39286 (N_39286,N_30647,N_33736);
nor U39287 (N_39287,N_31681,N_32243);
nor U39288 (N_39288,N_33116,N_33532);
xor U39289 (N_39289,N_33642,N_32412);
or U39290 (N_39290,N_33659,N_31786);
nand U39291 (N_39291,N_30634,N_31522);
and U39292 (N_39292,N_32272,N_33921);
xnor U39293 (N_39293,N_32703,N_31554);
xnor U39294 (N_39294,N_30015,N_33643);
nor U39295 (N_39295,N_30223,N_30534);
or U39296 (N_39296,N_30986,N_32958);
xnor U39297 (N_39297,N_31204,N_34794);
and U39298 (N_39298,N_30627,N_31966);
or U39299 (N_39299,N_33116,N_32649);
or U39300 (N_39300,N_34743,N_31445);
nand U39301 (N_39301,N_30878,N_34575);
nor U39302 (N_39302,N_32081,N_32968);
nand U39303 (N_39303,N_32373,N_30388);
xor U39304 (N_39304,N_30593,N_32947);
or U39305 (N_39305,N_33474,N_31786);
and U39306 (N_39306,N_30040,N_30368);
nor U39307 (N_39307,N_31030,N_34762);
and U39308 (N_39308,N_34065,N_34561);
or U39309 (N_39309,N_30013,N_33809);
nor U39310 (N_39310,N_31073,N_34363);
and U39311 (N_39311,N_33055,N_33091);
and U39312 (N_39312,N_32859,N_33279);
nand U39313 (N_39313,N_32146,N_34303);
nor U39314 (N_39314,N_33234,N_31549);
nand U39315 (N_39315,N_34088,N_30450);
xnor U39316 (N_39316,N_32729,N_30674);
and U39317 (N_39317,N_32659,N_32862);
nor U39318 (N_39318,N_32984,N_31457);
and U39319 (N_39319,N_34111,N_34538);
nand U39320 (N_39320,N_30334,N_32727);
nand U39321 (N_39321,N_31710,N_34494);
and U39322 (N_39322,N_34709,N_31123);
xor U39323 (N_39323,N_32446,N_33834);
nor U39324 (N_39324,N_30708,N_33898);
or U39325 (N_39325,N_31270,N_32041);
nor U39326 (N_39326,N_33234,N_32600);
and U39327 (N_39327,N_31059,N_30015);
nor U39328 (N_39328,N_31871,N_32041);
nand U39329 (N_39329,N_33317,N_30570);
xnor U39330 (N_39330,N_32310,N_34328);
or U39331 (N_39331,N_31472,N_30389);
or U39332 (N_39332,N_34439,N_34543);
and U39333 (N_39333,N_31526,N_34689);
nand U39334 (N_39334,N_30750,N_33288);
nand U39335 (N_39335,N_31420,N_32042);
xor U39336 (N_39336,N_30620,N_34081);
and U39337 (N_39337,N_31618,N_34870);
nand U39338 (N_39338,N_34716,N_30633);
xnor U39339 (N_39339,N_33330,N_34505);
and U39340 (N_39340,N_31464,N_33284);
nand U39341 (N_39341,N_30445,N_30671);
nand U39342 (N_39342,N_33004,N_33562);
and U39343 (N_39343,N_30881,N_32236);
nor U39344 (N_39344,N_31789,N_31883);
nand U39345 (N_39345,N_30705,N_34810);
and U39346 (N_39346,N_33820,N_32597);
nand U39347 (N_39347,N_31031,N_34348);
nand U39348 (N_39348,N_32568,N_32085);
xnor U39349 (N_39349,N_32512,N_32750);
nor U39350 (N_39350,N_33308,N_32631);
nand U39351 (N_39351,N_31867,N_30446);
and U39352 (N_39352,N_34954,N_32920);
or U39353 (N_39353,N_32168,N_30682);
nor U39354 (N_39354,N_33747,N_34491);
xor U39355 (N_39355,N_31605,N_34111);
nor U39356 (N_39356,N_32189,N_32588);
nor U39357 (N_39357,N_34716,N_32480);
or U39358 (N_39358,N_32585,N_33301);
xor U39359 (N_39359,N_30436,N_32887);
xor U39360 (N_39360,N_32842,N_31653);
xnor U39361 (N_39361,N_31792,N_34512);
nand U39362 (N_39362,N_33780,N_32179);
xor U39363 (N_39363,N_30821,N_33919);
nand U39364 (N_39364,N_34849,N_33733);
nor U39365 (N_39365,N_30929,N_32887);
xor U39366 (N_39366,N_32360,N_32992);
or U39367 (N_39367,N_30018,N_34955);
xnor U39368 (N_39368,N_34296,N_34291);
xnor U39369 (N_39369,N_31838,N_32764);
or U39370 (N_39370,N_31804,N_30445);
nor U39371 (N_39371,N_33881,N_30136);
nand U39372 (N_39372,N_34992,N_34890);
nor U39373 (N_39373,N_30484,N_31527);
xor U39374 (N_39374,N_31433,N_32940);
nand U39375 (N_39375,N_30953,N_30190);
xnor U39376 (N_39376,N_33023,N_32266);
nand U39377 (N_39377,N_34223,N_33908);
or U39378 (N_39378,N_34559,N_32807);
xor U39379 (N_39379,N_34606,N_32797);
nand U39380 (N_39380,N_34039,N_33898);
nand U39381 (N_39381,N_33854,N_34808);
and U39382 (N_39382,N_33902,N_34252);
and U39383 (N_39383,N_34978,N_33317);
nor U39384 (N_39384,N_34023,N_30651);
and U39385 (N_39385,N_30140,N_34459);
nand U39386 (N_39386,N_32051,N_32565);
xor U39387 (N_39387,N_33203,N_33664);
or U39388 (N_39388,N_34417,N_33121);
or U39389 (N_39389,N_31367,N_34058);
and U39390 (N_39390,N_31025,N_33589);
nand U39391 (N_39391,N_33562,N_31247);
nand U39392 (N_39392,N_33881,N_31953);
and U39393 (N_39393,N_31464,N_30759);
nor U39394 (N_39394,N_30835,N_32947);
or U39395 (N_39395,N_30740,N_33816);
nor U39396 (N_39396,N_32248,N_30150);
or U39397 (N_39397,N_31039,N_30330);
nand U39398 (N_39398,N_33564,N_33847);
nand U39399 (N_39399,N_30380,N_30365);
nand U39400 (N_39400,N_33746,N_34768);
or U39401 (N_39401,N_32064,N_34830);
nand U39402 (N_39402,N_30587,N_30877);
and U39403 (N_39403,N_34123,N_31171);
and U39404 (N_39404,N_32422,N_31253);
nand U39405 (N_39405,N_33112,N_34602);
nand U39406 (N_39406,N_33640,N_31216);
and U39407 (N_39407,N_33530,N_30647);
or U39408 (N_39408,N_32804,N_30554);
xor U39409 (N_39409,N_31866,N_32646);
nand U39410 (N_39410,N_32094,N_32872);
or U39411 (N_39411,N_34943,N_34808);
and U39412 (N_39412,N_32947,N_31779);
nand U39413 (N_39413,N_34395,N_31364);
or U39414 (N_39414,N_30619,N_34636);
and U39415 (N_39415,N_32051,N_31076);
xnor U39416 (N_39416,N_31326,N_33136);
nor U39417 (N_39417,N_34603,N_34117);
nor U39418 (N_39418,N_32590,N_33223);
and U39419 (N_39419,N_30161,N_33077);
nand U39420 (N_39420,N_34341,N_30675);
or U39421 (N_39421,N_33599,N_32639);
nand U39422 (N_39422,N_33808,N_31712);
or U39423 (N_39423,N_33700,N_30620);
or U39424 (N_39424,N_30353,N_33292);
xnor U39425 (N_39425,N_34479,N_30748);
and U39426 (N_39426,N_34320,N_32806);
and U39427 (N_39427,N_34693,N_31826);
and U39428 (N_39428,N_34268,N_30446);
nor U39429 (N_39429,N_30653,N_33535);
nor U39430 (N_39430,N_31510,N_34369);
nand U39431 (N_39431,N_34304,N_33897);
nor U39432 (N_39432,N_32738,N_30603);
xor U39433 (N_39433,N_30222,N_30074);
nand U39434 (N_39434,N_32406,N_30496);
and U39435 (N_39435,N_34075,N_33174);
nand U39436 (N_39436,N_31815,N_33250);
nor U39437 (N_39437,N_32093,N_30666);
nor U39438 (N_39438,N_33277,N_31521);
or U39439 (N_39439,N_31550,N_30248);
nor U39440 (N_39440,N_33862,N_33839);
nor U39441 (N_39441,N_32906,N_30187);
nor U39442 (N_39442,N_33034,N_34440);
xnor U39443 (N_39443,N_32074,N_32094);
or U39444 (N_39444,N_31642,N_33861);
nor U39445 (N_39445,N_32223,N_33508);
and U39446 (N_39446,N_30289,N_34120);
nand U39447 (N_39447,N_34739,N_32690);
nor U39448 (N_39448,N_31280,N_30840);
and U39449 (N_39449,N_30665,N_33970);
nand U39450 (N_39450,N_34719,N_32786);
or U39451 (N_39451,N_32977,N_33006);
or U39452 (N_39452,N_33088,N_34009);
or U39453 (N_39453,N_33326,N_31787);
or U39454 (N_39454,N_33312,N_33834);
xor U39455 (N_39455,N_32599,N_33211);
and U39456 (N_39456,N_31178,N_31551);
xor U39457 (N_39457,N_30042,N_31299);
xor U39458 (N_39458,N_30219,N_33405);
nor U39459 (N_39459,N_30062,N_32898);
nor U39460 (N_39460,N_30194,N_33558);
and U39461 (N_39461,N_34612,N_32860);
or U39462 (N_39462,N_34000,N_31298);
and U39463 (N_39463,N_33354,N_31853);
and U39464 (N_39464,N_30076,N_31065);
and U39465 (N_39465,N_34963,N_33262);
nand U39466 (N_39466,N_34430,N_32736);
xnor U39467 (N_39467,N_30487,N_34630);
and U39468 (N_39468,N_30204,N_32582);
or U39469 (N_39469,N_30040,N_33441);
xnor U39470 (N_39470,N_32920,N_33930);
or U39471 (N_39471,N_34296,N_32149);
xnor U39472 (N_39472,N_33180,N_30013);
xor U39473 (N_39473,N_30084,N_33061);
nand U39474 (N_39474,N_31096,N_31896);
nand U39475 (N_39475,N_31150,N_32101);
nor U39476 (N_39476,N_32381,N_32636);
or U39477 (N_39477,N_31120,N_33947);
xor U39478 (N_39478,N_30673,N_33239);
nand U39479 (N_39479,N_33837,N_31588);
nor U39480 (N_39480,N_31560,N_31336);
and U39481 (N_39481,N_33821,N_30276);
nand U39482 (N_39482,N_32914,N_34256);
xnor U39483 (N_39483,N_31742,N_32693);
or U39484 (N_39484,N_32914,N_33283);
nand U39485 (N_39485,N_33052,N_31810);
and U39486 (N_39486,N_34518,N_32132);
or U39487 (N_39487,N_32414,N_32915);
xor U39488 (N_39488,N_34306,N_31493);
or U39489 (N_39489,N_32524,N_30257);
or U39490 (N_39490,N_32245,N_34414);
and U39491 (N_39491,N_31661,N_32740);
or U39492 (N_39492,N_34148,N_31838);
nor U39493 (N_39493,N_34344,N_33345);
xor U39494 (N_39494,N_30915,N_32783);
or U39495 (N_39495,N_30787,N_34943);
or U39496 (N_39496,N_31865,N_32982);
and U39497 (N_39497,N_34680,N_32934);
or U39498 (N_39498,N_32629,N_30139);
xnor U39499 (N_39499,N_32230,N_30334);
nand U39500 (N_39500,N_33719,N_31133);
xnor U39501 (N_39501,N_34174,N_31425);
nor U39502 (N_39502,N_34412,N_34178);
and U39503 (N_39503,N_30360,N_32981);
nand U39504 (N_39504,N_33155,N_30355);
nand U39505 (N_39505,N_34161,N_31184);
and U39506 (N_39506,N_30726,N_34000);
xnor U39507 (N_39507,N_34696,N_31455);
nand U39508 (N_39508,N_31711,N_33182);
nand U39509 (N_39509,N_30789,N_31035);
nor U39510 (N_39510,N_33449,N_31767);
or U39511 (N_39511,N_32186,N_32349);
xor U39512 (N_39512,N_30865,N_32816);
nand U39513 (N_39513,N_33681,N_31697);
nor U39514 (N_39514,N_33319,N_31561);
and U39515 (N_39515,N_32669,N_32955);
nor U39516 (N_39516,N_30084,N_31662);
and U39517 (N_39517,N_31853,N_31626);
nor U39518 (N_39518,N_32326,N_32648);
xor U39519 (N_39519,N_31271,N_34006);
or U39520 (N_39520,N_34018,N_31675);
nor U39521 (N_39521,N_34774,N_34557);
nor U39522 (N_39522,N_34389,N_30218);
or U39523 (N_39523,N_30960,N_33654);
nand U39524 (N_39524,N_30151,N_33233);
nand U39525 (N_39525,N_30844,N_31492);
nor U39526 (N_39526,N_34052,N_30723);
nor U39527 (N_39527,N_32666,N_34076);
or U39528 (N_39528,N_31030,N_33085);
nand U39529 (N_39529,N_30686,N_34032);
nand U39530 (N_39530,N_31756,N_31646);
nand U39531 (N_39531,N_33454,N_34665);
xnor U39532 (N_39532,N_32533,N_30534);
nand U39533 (N_39533,N_33386,N_32411);
and U39534 (N_39534,N_33873,N_31141);
or U39535 (N_39535,N_30676,N_33118);
or U39536 (N_39536,N_30802,N_32100);
nor U39537 (N_39537,N_34091,N_31452);
and U39538 (N_39538,N_30173,N_34160);
and U39539 (N_39539,N_34175,N_32105);
nor U39540 (N_39540,N_31875,N_32001);
nor U39541 (N_39541,N_32816,N_30128);
nor U39542 (N_39542,N_32404,N_32006);
or U39543 (N_39543,N_31405,N_31362);
and U39544 (N_39544,N_33067,N_30125);
or U39545 (N_39545,N_32734,N_32616);
and U39546 (N_39546,N_32020,N_33585);
nor U39547 (N_39547,N_31925,N_31774);
or U39548 (N_39548,N_33883,N_32953);
and U39549 (N_39549,N_31998,N_30968);
nand U39550 (N_39550,N_34877,N_32663);
xnor U39551 (N_39551,N_32479,N_31042);
or U39552 (N_39552,N_33222,N_32377);
nor U39553 (N_39553,N_30953,N_30727);
nand U39554 (N_39554,N_31936,N_33862);
nand U39555 (N_39555,N_31337,N_33180);
nand U39556 (N_39556,N_32273,N_34107);
and U39557 (N_39557,N_32105,N_30784);
xor U39558 (N_39558,N_31368,N_34013);
nor U39559 (N_39559,N_34747,N_34818);
and U39560 (N_39560,N_30595,N_33331);
nor U39561 (N_39561,N_34431,N_32693);
nor U39562 (N_39562,N_33836,N_33654);
nand U39563 (N_39563,N_34001,N_33794);
xnor U39564 (N_39564,N_32066,N_30184);
nor U39565 (N_39565,N_31488,N_33414);
nor U39566 (N_39566,N_33476,N_34039);
and U39567 (N_39567,N_33226,N_34433);
xor U39568 (N_39568,N_33341,N_32643);
xor U39569 (N_39569,N_32951,N_32259);
nand U39570 (N_39570,N_31553,N_31844);
nor U39571 (N_39571,N_30343,N_32410);
and U39572 (N_39572,N_30151,N_31547);
or U39573 (N_39573,N_31518,N_33691);
xor U39574 (N_39574,N_31045,N_32470);
or U39575 (N_39575,N_30820,N_34802);
nand U39576 (N_39576,N_30385,N_31755);
nor U39577 (N_39577,N_33524,N_32149);
xor U39578 (N_39578,N_33920,N_34878);
and U39579 (N_39579,N_32035,N_34011);
xor U39580 (N_39580,N_34344,N_31176);
and U39581 (N_39581,N_31559,N_34412);
xor U39582 (N_39582,N_33562,N_32770);
or U39583 (N_39583,N_34125,N_32397);
or U39584 (N_39584,N_32411,N_32003);
xor U39585 (N_39585,N_30394,N_30870);
xnor U39586 (N_39586,N_30080,N_32827);
nor U39587 (N_39587,N_30198,N_30511);
xor U39588 (N_39588,N_32973,N_32488);
and U39589 (N_39589,N_31419,N_30850);
or U39590 (N_39590,N_33653,N_34773);
and U39591 (N_39591,N_31399,N_30546);
xor U39592 (N_39592,N_34360,N_31486);
nor U39593 (N_39593,N_34583,N_33118);
or U39594 (N_39594,N_31834,N_30816);
and U39595 (N_39595,N_30820,N_30430);
xor U39596 (N_39596,N_34596,N_34263);
xnor U39597 (N_39597,N_31956,N_31645);
and U39598 (N_39598,N_34669,N_33005);
and U39599 (N_39599,N_30453,N_33032);
and U39600 (N_39600,N_34326,N_34722);
xor U39601 (N_39601,N_34777,N_30913);
or U39602 (N_39602,N_34798,N_33455);
nor U39603 (N_39603,N_31412,N_31170);
xnor U39604 (N_39604,N_31818,N_33525);
nor U39605 (N_39605,N_34044,N_33608);
and U39606 (N_39606,N_34735,N_31999);
nand U39607 (N_39607,N_32092,N_33513);
xnor U39608 (N_39608,N_32428,N_31340);
and U39609 (N_39609,N_32985,N_31609);
or U39610 (N_39610,N_32253,N_34918);
nand U39611 (N_39611,N_31365,N_30134);
and U39612 (N_39612,N_34070,N_30480);
xnor U39613 (N_39613,N_32121,N_31574);
or U39614 (N_39614,N_30552,N_31336);
nor U39615 (N_39615,N_31492,N_33508);
nor U39616 (N_39616,N_32579,N_30816);
nor U39617 (N_39617,N_32529,N_30731);
and U39618 (N_39618,N_31135,N_33178);
nor U39619 (N_39619,N_32949,N_30995);
nand U39620 (N_39620,N_30367,N_30825);
nand U39621 (N_39621,N_34508,N_32212);
xnor U39622 (N_39622,N_31422,N_32004);
xor U39623 (N_39623,N_32032,N_30648);
or U39624 (N_39624,N_34750,N_33548);
or U39625 (N_39625,N_32882,N_32558);
nand U39626 (N_39626,N_34176,N_32906);
nand U39627 (N_39627,N_32677,N_32733);
and U39628 (N_39628,N_33345,N_30663);
xor U39629 (N_39629,N_30672,N_30224);
and U39630 (N_39630,N_31330,N_34297);
xnor U39631 (N_39631,N_34427,N_33473);
or U39632 (N_39632,N_32723,N_34966);
nor U39633 (N_39633,N_31607,N_31010);
nand U39634 (N_39634,N_33546,N_33400);
nand U39635 (N_39635,N_34235,N_33728);
and U39636 (N_39636,N_30521,N_32665);
or U39637 (N_39637,N_30953,N_30813);
nor U39638 (N_39638,N_32373,N_30423);
or U39639 (N_39639,N_32358,N_30239);
and U39640 (N_39640,N_32948,N_34560);
xnor U39641 (N_39641,N_33611,N_31997);
xor U39642 (N_39642,N_34929,N_33209);
nor U39643 (N_39643,N_32692,N_32219);
nor U39644 (N_39644,N_34203,N_34958);
nand U39645 (N_39645,N_31879,N_32011);
or U39646 (N_39646,N_31806,N_32255);
nor U39647 (N_39647,N_34332,N_34665);
nor U39648 (N_39648,N_34569,N_33784);
or U39649 (N_39649,N_34138,N_31966);
nor U39650 (N_39650,N_32840,N_31305);
nand U39651 (N_39651,N_32668,N_31008);
xor U39652 (N_39652,N_31003,N_30812);
xnor U39653 (N_39653,N_32936,N_33434);
and U39654 (N_39654,N_33910,N_34757);
nor U39655 (N_39655,N_33882,N_32026);
or U39656 (N_39656,N_30702,N_32415);
xor U39657 (N_39657,N_30401,N_31850);
xnor U39658 (N_39658,N_33331,N_32263);
xnor U39659 (N_39659,N_30375,N_32736);
and U39660 (N_39660,N_32457,N_33638);
or U39661 (N_39661,N_30005,N_30841);
nor U39662 (N_39662,N_30743,N_32130);
and U39663 (N_39663,N_31421,N_30891);
xnor U39664 (N_39664,N_33619,N_30489);
nand U39665 (N_39665,N_30807,N_34983);
or U39666 (N_39666,N_32166,N_31682);
nand U39667 (N_39667,N_30468,N_31608);
or U39668 (N_39668,N_34724,N_30935);
nor U39669 (N_39669,N_32539,N_32477);
nor U39670 (N_39670,N_32545,N_32366);
and U39671 (N_39671,N_32843,N_31405);
nand U39672 (N_39672,N_32949,N_31136);
nor U39673 (N_39673,N_33442,N_31686);
xor U39674 (N_39674,N_33450,N_32333);
nand U39675 (N_39675,N_32657,N_30338);
xnor U39676 (N_39676,N_32707,N_34007);
nor U39677 (N_39677,N_33889,N_34678);
and U39678 (N_39678,N_33883,N_32153);
nand U39679 (N_39679,N_31163,N_34548);
or U39680 (N_39680,N_31641,N_34860);
xor U39681 (N_39681,N_31604,N_30599);
or U39682 (N_39682,N_30650,N_31817);
and U39683 (N_39683,N_33347,N_31265);
nor U39684 (N_39684,N_33241,N_34408);
xnor U39685 (N_39685,N_32247,N_30039);
nor U39686 (N_39686,N_30458,N_30121);
and U39687 (N_39687,N_34385,N_31651);
nor U39688 (N_39688,N_31553,N_33541);
or U39689 (N_39689,N_31112,N_30154);
and U39690 (N_39690,N_30001,N_31017);
nand U39691 (N_39691,N_32543,N_31752);
xnor U39692 (N_39692,N_34164,N_32300);
xnor U39693 (N_39693,N_31348,N_30531);
or U39694 (N_39694,N_32899,N_33411);
and U39695 (N_39695,N_30200,N_34991);
nor U39696 (N_39696,N_34498,N_32437);
or U39697 (N_39697,N_34883,N_34265);
nor U39698 (N_39698,N_34959,N_31188);
and U39699 (N_39699,N_32483,N_31232);
nor U39700 (N_39700,N_30895,N_32271);
and U39701 (N_39701,N_30386,N_34772);
nand U39702 (N_39702,N_31217,N_32706);
or U39703 (N_39703,N_33366,N_34699);
nand U39704 (N_39704,N_34912,N_34515);
nand U39705 (N_39705,N_34112,N_30065);
nor U39706 (N_39706,N_34511,N_31186);
nand U39707 (N_39707,N_32762,N_30584);
and U39708 (N_39708,N_34702,N_31879);
nand U39709 (N_39709,N_34724,N_31736);
nor U39710 (N_39710,N_32314,N_31992);
nor U39711 (N_39711,N_32428,N_33713);
or U39712 (N_39712,N_34080,N_34443);
or U39713 (N_39713,N_34047,N_30361);
or U39714 (N_39714,N_33473,N_31172);
and U39715 (N_39715,N_30042,N_31469);
or U39716 (N_39716,N_33109,N_31703);
and U39717 (N_39717,N_30257,N_30692);
xor U39718 (N_39718,N_30909,N_34658);
nor U39719 (N_39719,N_33875,N_30550);
or U39720 (N_39720,N_32097,N_31448);
and U39721 (N_39721,N_33560,N_30264);
or U39722 (N_39722,N_31806,N_34960);
xor U39723 (N_39723,N_33456,N_34905);
or U39724 (N_39724,N_34210,N_33404);
and U39725 (N_39725,N_31857,N_33833);
or U39726 (N_39726,N_31955,N_32217);
or U39727 (N_39727,N_32125,N_31783);
or U39728 (N_39728,N_30319,N_33911);
xnor U39729 (N_39729,N_34182,N_32061);
nor U39730 (N_39730,N_32156,N_33766);
nor U39731 (N_39731,N_34454,N_33648);
xnor U39732 (N_39732,N_30851,N_34555);
xnor U39733 (N_39733,N_32335,N_33842);
or U39734 (N_39734,N_33733,N_32553);
and U39735 (N_39735,N_33538,N_31355);
xor U39736 (N_39736,N_31890,N_32562);
nor U39737 (N_39737,N_32546,N_32230);
or U39738 (N_39738,N_30692,N_32854);
nand U39739 (N_39739,N_34823,N_31935);
nor U39740 (N_39740,N_33051,N_34211);
and U39741 (N_39741,N_31192,N_33663);
and U39742 (N_39742,N_32616,N_32405);
and U39743 (N_39743,N_33345,N_32440);
and U39744 (N_39744,N_30178,N_33898);
nor U39745 (N_39745,N_32228,N_32879);
and U39746 (N_39746,N_32397,N_32702);
and U39747 (N_39747,N_33509,N_34001);
nor U39748 (N_39748,N_30498,N_33596);
xor U39749 (N_39749,N_33690,N_32143);
and U39750 (N_39750,N_30238,N_32303);
nor U39751 (N_39751,N_33383,N_30713);
nand U39752 (N_39752,N_31358,N_33280);
nor U39753 (N_39753,N_30959,N_30116);
nor U39754 (N_39754,N_31707,N_34658);
nand U39755 (N_39755,N_30291,N_33928);
nand U39756 (N_39756,N_34878,N_32543);
and U39757 (N_39757,N_30467,N_31411);
and U39758 (N_39758,N_32642,N_31342);
and U39759 (N_39759,N_32220,N_34462);
and U39760 (N_39760,N_33961,N_30892);
nand U39761 (N_39761,N_33495,N_33062);
nor U39762 (N_39762,N_30570,N_33826);
or U39763 (N_39763,N_33239,N_31532);
xnor U39764 (N_39764,N_31889,N_34667);
nand U39765 (N_39765,N_32967,N_30547);
nand U39766 (N_39766,N_33604,N_32819);
and U39767 (N_39767,N_30918,N_33735);
and U39768 (N_39768,N_33786,N_31768);
nand U39769 (N_39769,N_31666,N_34356);
nor U39770 (N_39770,N_30729,N_31463);
nor U39771 (N_39771,N_30256,N_32709);
or U39772 (N_39772,N_30101,N_31907);
nand U39773 (N_39773,N_34350,N_34150);
or U39774 (N_39774,N_30050,N_32463);
nand U39775 (N_39775,N_33798,N_34506);
nor U39776 (N_39776,N_32628,N_34613);
and U39777 (N_39777,N_31469,N_33476);
or U39778 (N_39778,N_31613,N_30657);
nor U39779 (N_39779,N_34301,N_34012);
xor U39780 (N_39780,N_33066,N_34691);
xnor U39781 (N_39781,N_34955,N_32445);
or U39782 (N_39782,N_34039,N_32163);
nor U39783 (N_39783,N_30811,N_30605);
nor U39784 (N_39784,N_31927,N_31131);
or U39785 (N_39785,N_33586,N_34386);
or U39786 (N_39786,N_30203,N_32279);
and U39787 (N_39787,N_32271,N_33140);
or U39788 (N_39788,N_31078,N_33624);
or U39789 (N_39789,N_33115,N_33967);
or U39790 (N_39790,N_32011,N_31461);
or U39791 (N_39791,N_30641,N_33585);
nand U39792 (N_39792,N_31530,N_32731);
or U39793 (N_39793,N_30030,N_32464);
xnor U39794 (N_39794,N_31397,N_32428);
nand U39795 (N_39795,N_30560,N_33444);
nand U39796 (N_39796,N_30334,N_32938);
xnor U39797 (N_39797,N_34080,N_33917);
nor U39798 (N_39798,N_34020,N_33845);
nand U39799 (N_39799,N_33283,N_31282);
and U39800 (N_39800,N_34361,N_31585);
nand U39801 (N_39801,N_34306,N_31946);
or U39802 (N_39802,N_33839,N_31217);
nand U39803 (N_39803,N_30834,N_34955);
xor U39804 (N_39804,N_34638,N_32890);
or U39805 (N_39805,N_30758,N_31606);
xor U39806 (N_39806,N_34955,N_32006);
nor U39807 (N_39807,N_32451,N_31317);
and U39808 (N_39808,N_33408,N_32646);
or U39809 (N_39809,N_34529,N_30129);
or U39810 (N_39810,N_32279,N_33811);
or U39811 (N_39811,N_34503,N_32620);
and U39812 (N_39812,N_30970,N_32976);
xnor U39813 (N_39813,N_34834,N_32744);
or U39814 (N_39814,N_32301,N_33109);
or U39815 (N_39815,N_33237,N_30145);
and U39816 (N_39816,N_34987,N_30730);
xnor U39817 (N_39817,N_31248,N_32241);
xnor U39818 (N_39818,N_34874,N_30051);
nor U39819 (N_39819,N_30845,N_34261);
xnor U39820 (N_39820,N_30114,N_30406);
and U39821 (N_39821,N_30549,N_32046);
nor U39822 (N_39822,N_34360,N_30028);
xnor U39823 (N_39823,N_31265,N_32887);
nor U39824 (N_39824,N_33376,N_30583);
xor U39825 (N_39825,N_34588,N_30704);
nand U39826 (N_39826,N_30957,N_33300);
xor U39827 (N_39827,N_32861,N_31836);
xor U39828 (N_39828,N_31904,N_33269);
and U39829 (N_39829,N_34021,N_30854);
and U39830 (N_39830,N_33226,N_33261);
nand U39831 (N_39831,N_32872,N_33337);
xor U39832 (N_39832,N_30257,N_31525);
xnor U39833 (N_39833,N_34207,N_32149);
xor U39834 (N_39834,N_31583,N_30048);
nor U39835 (N_39835,N_33758,N_34865);
and U39836 (N_39836,N_33251,N_32121);
xor U39837 (N_39837,N_31138,N_31358);
xor U39838 (N_39838,N_30625,N_30811);
xnor U39839 (N_39839,N_34906,N_32876);
xor U39840 (N_39840,N_33560,N_34632);
and U39841 (N_39841,N_33530,N_30552);
xnor U39842 (N_39842,N_34084,N_34213);
nand U39843 (N_39843,N_30446,N_30249);
nand U39844 (N_39844,N_32955,N_33565);
or U39845 (N_39845,N_30277,N_32789);
nor U39846 (N_39846,N_33309,N_32226);
and U39847 (N_39847,N_31992,N_31902);
or U39848 (N_39848,N_31645,N_32812);
nor U39849 (N_39849,N_30258,N_31929);
nand U39850 (N_39850,N_33057,N_30345);
and U39851 (N_39851,N_33951,N_30783);
nand U39852 (N_39852,N_32983,N_34417);
or U39853 (N_39853,N_33369,N_34333);
or U39854 (N_39854,N_31464,N_32778);
and U39855 (N_39855,N_33451,N_33947);
nor U39856 (N_39856,N_30159,N_30888);
and U39857 (N_39857,N_33325,N_32896);
or U39858 (N_39858,N_34529,N_32925);
nand U39859 (N_39859,N_30805,N_30612);
and U39860 (N_39860,N_31251,N_30296);
nor U39861 (N_39861,N_31037,N_32128);
nor U39862 (N_39862,N_33162,N_32371);
nand U39863 (N_39863,N_32233,N_30734);
nor U39864 (N_39864,N_34213,N_33290);
or U39865 (N_39865,N_32397,N_30196);
or U39866 (N_39866,N_32415,N_30974);
nand U39867 (N_39867,N_33310,N_31468);
nand U39868 (N_39868,N_30798,N_34657);
nand U39869 (N_39869,N_33815,N_32783);
nor U39870 (N_39870,N_33548,N_31380);
and U39871 (N_39871,N_33226,N_32848);
or U39872 (N_39872,N_30091,N_30852);
and U39873 (N_39873,N_32629,N_33897);
or U39874 (N_39874,N_33411,N_32751);
xor U39875 (N_39875,N_31726,N_32895);
nor U39876 (N_39876,N_34232,N_33616);
and U39877 (N_39877,N_32003,N_34360);
nor U39878 (N_39878,N_34195,N_32158);
nor U39879 (N_39879,N_33342,N_31703);
and U39880 (N_39880,N_31886,N_30382);
and U39881 (N_39881,N_34763,N_34181);
nor U39882 (N_39882,N_33321,N_34920);
nand U39883 (N_39883,N_34756,N_33786);
and U39884 (N_39884,N_34053,N_31703);
nor U39885 (N_39885,N_33289,N_34507);
xor U39886 (N_39886,N_32161,N_34118);
or U39887 (N_39887,N_30421,N_30445);
nor U39888 (N_39888,N_31632,N_32616);
xnor U39889 (N_39889,N_30950,N_30465);
nor U39890 (N_39890,N_30031,N_34605);
nand U39891 (N_39891,N_34738,N_30908);
nand U39892 (N_39892,N_30380,N_32649);
xnor U39893 (N_39893,N_30299,N_30070);
or U39894 (N_39894,N_31400,N_33053);
and U39895 (N_39895,N_34045,N_31550);
nor U39896 (N_39896,N_34484,N_34856);
and U39897 (N_39897,N_30683,N_33740);
nand U39898 (N_39898,N_33590,N_33566);
nand U39899 (N_39899,N_31414,N_34558);
nand U39900 (N_39900,N_34252,N_31323);
nand U39901 (N_39901,N_31341,N_34047);
nand U39902 (N_39902,N_32456,N_33408);
nor U39903 (N_39903,N_31972,N_32755);
nor U39904 (N_39904,N_33077,N_33334);
and U39905 (N_39905,N_31893,N_34947);
nand U39906 (N_39906,N_31487,N_33734);
nand U39907 (N_39907,N_30635,N_32208);
or U39908 (N_39908,N_34715,N_34173);
and U39909 (N_39909,N_31474,N_31721);
or U39910 (N_39910,N_32541,N_34271);
or U39911 (N_39911,N_33504,N_30943);
xnor U39912 (N_39912,N_33032,N_30573);
or U39913 (N_39913,N_32759,N_33715);
nor U39914 (N_39914,N_30557,N_32562);
or U39915 (N_39915,N_33570,N_31857);
and U39916 (N_39916,N_34437,N_33666);
nand U39917 (N_39917,N_34004,N_33385);
or U39918 (N_39918,N_31956,N_31507);
xnor U39919 (N_39919,N_32214,N_32402);
nor U39920 (N_39920,N_31991,N_30318);
or U39921 (N_39921,N_30666,N_30790);
nand U39922 (N_39922,N_33194,N_33259);
xor U39923 (N_39923,N_34846,N_34932);
xor U39924 (N_39924,N_33420,N_30553);
nand U39925 (N_39925,N_33649,N_30889);
or U39926 (N_39926,N_31826,N_32734);
or U39927 (N_39927,N_32460,N_31724);
nand U39928 (N_39928,N_31248,N_31461);
nor U39929 (N_39929,N_33685,N_33424);
xnor U39930 (N_39930,N_31413,N_30110);
nand U39931 (N_39931,N_33275,N_34311);
nand U39932 (N_39932,N_34784,N_30275);
or U39933 (N_39933,N_32558,N_32388);
or U39934 (N_39934,N_33564,N_34677);
and U39935 (N_39935,N_30086,N_34075);
and U39936 (N_39936,N_31714,N_30019);
nor U39937 (N_39937,N_34484,N_31075);
and U39938 (N_39938,N_34806,N_32693);
xnor U39939 (N_39939,N_31150,N_34213);
or U39940 (N_39940,N_31998,N_34346);
and U39941 (N_39941,N_32333,N_32904);
or U39942 (N_39942,N_33562,N_30916);
nor U39943 (N_39943,N_34862,N_33234);
xnor U39944 (N_39944,N_30415,N_31414);
nor U39945 (N_39945,N_34686,N_30536);
xnor U39946 (N_39946,N_30426,N_33824);
xor U39947 (N_39947,N_30262,N_33139);
nor U39948 (N_39948,N_34823,N_30143);
xnor U39949 (N_39949,N_30773,N_34468);
or U39950 (N_39950,N_32944,N_31478);
xnor U39951 (N_39951,N_30651,N_32640);
xor U39952 (N_39952,N_30620,N_31952);
and U39953 (N_39953,N_34300,N_32030);
nand U39954 (N_39954,N_34737,N_30153);
and U39955 (N_39955,N_30628,N_32560);
and U39956 (N_39956,N_32753,N_33266);
nand U39957 (N_39957,N_33668,N_30946);
xor U39958 (N_39958,N_32535,N_32438);
nand U39959 (N_39959,N_33049,N_33398);
nor U39960 (N_39960,N_33482,N_33849);
and U39961 (N_39961,N_32291,N_31699);
or U39962 (N_39962,N_30371,N_30960);
nand U39963 (N_39963,N_33721,N_33536);
xnor U39964 (N_39964,N_32656,N_33056);
nand U39965 (N_39965,N_31302,N_32061);
and U39966 (N_39966,N_33842,N_34440);
and U39967 (N_39967,N_30892,N_32567);
and U39968 (N_39968,N_34407,N_32161);
and U39969 (N_39969,N_31496,N_30036);
and U39970 (N_39970,N_34681,N_30808);
and U39971 (N_39971,N_33944,N_32633);
or U39972 (N_39972,N_30618,N_33346);
or U39973 (N_39973,N_30662,N_31371);
or U39974 (N_39974,N_31552,N_30401);
nand U39975 (N_39975,N_34386,N_30344);
or U39976 (N_39976,N_30606,N_34426);
nand U39977 (N_39977,N_31117,N_34722);
nor U39978 (N_39978,N_32791,N_33907);
xnor U39979 (N_39979,N_30456,N_34310);
xor U39980 (N_39980,N_30830,N_32106);
and U39981 (N_39981,N_34861,N_32932);
or U39982 (N_39982,N_31889,N_32030);
nand U39983 (N_39983,N_30293,N_31064);
and U39984 (N_39984,N_33583,N_33227);
or U39985 (N_39985,N_34081,N_32345);
nand U39986 (N_39986,N_33852,N_32686);
xor U39987 (N_39987,N_33865,N_31633);
and U39988 (N_39988,N_34174,N_34570);
nor U39989 (N_39989,N_30785,N_30841);
or U39990 (N_39990,N_30311,N_34826);
and U39991 (N_39991,N_33685,N_33503);
nor U39992 (N_39992,N_32017,N_32670);
nor U39993 (N_39993,N_34685,N_34281);
nor U39994 (N_39994,N_32326,N_30981);
and U39995 (N_39995,N_33234,N_32855);
and U39996 (N_39996,N_33178,N_34393);
xor U39997 (N_39997,N_31099,N_31534);
nor U39998 (N_39998,N_33246,N_32692);
nor U39999 (N_39999,N_30648,N_31683);
or U40000 (N_40000,N_38401,N_39917);
or U40001 (N_40001,N_39431,N_37893);
nor U40002 (N_40002,N_35035,N_39781);
nand U40003 (N_40003,N_37161,N_39971);
or U40004 (N_40004,N_38523,N_37702);
and U40005 (N_40005,N_35521,N_35566);
xnor U40006 (N_40006,N_39119,N_35995);
and U40007 (N_40007,N_36004,N_37971);
and U40008 (N_40008,N_37026,N_36246);
nand U40009 (N_40009,N_37583,N_39098);
xor U40010 (N_40010,N_35022,N_35003);
nand U40011 (N_40011,N_39452,N_39738);
or U40012 (N_40012,N_37946,N_38159);
xor U40013 (N_40013,N_36235,N_35222);
and U40014 (N_40014,N_39358,N_38054);
or U40015 (N_40015,N_36305,N_37945);
nand U40016 (N_40016,N_37638,N_35043);
or U40017 (N_40017,N_36698,N_36466);
nor U40018 (N_40018,N_36750,N_36752);
and U40019 (N_40019,N_38620,N_37829);
nand U40020 (N_40020,N_37754,N_35607);
and U40021 (N_40021,N_37028,N_38173);
nand U40022 (N_40022,N_37207,N_37392);
nor U40023 (N_40023,N_37200,N_36574);
nand U40024 (N_40024,N_37813,N_38410);
xnor U40025 (N_40025,N_39132,N_36505);
or U40026 (N_40026,N_38970,N_37628);
and U40027 (N_40027,N_36947,N_36177);
xor U40028 (N_40028,N_39699,N_38567);
nor U40029 (N_40029,N_36497,N_37598);
nand U40030 (N_40030,N_38099,N_37578);
xnor U40031 (N_40031,N_39862,N_36735);
xor U40032 (N_40032,N_38486,N_36333);
nor U40033 (N_40033,N_39664,N_35723);
nor U40034 (N_40034,N_36804,N_37494);
xor U40035 (N_40035,N_39476,N_37928);
nor U40036 (N_40036,N_35650,N_36648);
and U40037 (N_40037,N_39042,N_39133);
or U40038 (N_40038,N_37532,N_36686);
and U40039 (N_40039,N_39461,N_37184);
and U40040 (N_40040,N_38751,N_36808);
nor U40041 (N_40041,N_39574,N_38538);
nor U40042 (N_40042,N_39730,N_39182);
nor U40043 (N_40043,N_39618,N_36137);
xor U40044 (N_40044,N_37199,N_39563);
or U40045 (N_40045,N_36167,N_37958);
nor U40046 (N_40046,N_35265,N_36352);
nor U40047 (N_40047,N_35688,N_39253);
nor U40048 (N_40048,N_37349,N_35161);
nand U40049 (N_40049,N_35441,N_37544);
nand U40050 (N_40050,N_35407,N_37446);
nor U40051 (N_40051,N_35060,N_39580);
and U40052 (N_40052,N_36168,N_35386);
or U40053 (N_40053,N_37575,N_36579);
and U40054 (N_40054,N_39802,N_35643);
nor U40055 (N_40055,N_37197,N_36222);
and U40056 (N_40056,N_39866,N_39824);
nor U40057 (N_40057,N_36960,N_35203);
and U40058 (N_40058,N_38740,N_38676);
xnor U40059 (N_40059,N_35131,N_39295);
nor U40060 (N_40060,N_35352,N_36549);
and U40061 (N_40061,N_36530,N_38644);
nand U40062 (N_40062,N_36240,N_38507);
nor U40063 (N_40063,N_39659,N_38650);
and U40064 (N_40064,N_35534,N_37175);
nand U40065 (N_40065,N_36276,N_39887);
xnor U40066 (N_40066,N_37972,N_36347);
and U40067 (N_40067,N_35246,N_37894);
nand U40068 (N_40068,N_39684,N_35686);
or U40069 (N_40069,N_35026,N_37925);
nand U40070 (N_40070,N_38298,N_35269);
nor U40071 (N_40071,N_36714,N_37097);
and U40072 (N_40072,N_35991,N_36248);
xnor U40073 (N_40073,N_39875,N_37570);
and U40074 (N_40074,N_36994,N_37213);
xnor U40075 (N_40075,N_37084,N_36812);
or U40076 (N_40076,N_36557,N_38016);
and U40077 (N_40077,N_35618,N_36899);
or U40078 (N_40078,N_36626,N_37872);
nor U40079 (N_40079,N_39316,N_35539);
xor U40080 (N_40080,N_35801,N_39255);
or U40081 (N_40081,N_37183,N_38842);
nand U40082 (N_40082,N_35102,N_35389);
and U40083 (N_40083,N_36535,N_36928);
nor U40084 (N_40084,N_36744,N_39429);
nor U40085 (N_40085,N_36763,N_38284);
and U40086 (N_40086,N_39005,N_36067);
or U40087 (N_40087,N_36739,N_35829);
or U40088 (N_40088,N_39660,N_36609);
nor U40089 (N_40089,N_39625,N_36554);
nand U40090 (N_40090,N_38420,N_35355);
xor U40091 (N_40091,N_39127,N_38922);
xnor U40092 (N_40092,N_38807,N_38626);
and U40093 (N_40093,N_38301,N_35239);
or U40094 (N_40094,N_39532,N_35270);
nand U40095 (N_40095,N_37838,N_38886);
or U40096 (N_40096,N_37630,N_38458);
or U40097 (N_40097,N_38382,N_37879);
nand U40098 (N_40098,N_36369,N_37451);
or U40099 (N_40099,N_38192,N_36071);
and U40100 (N_40100,N_35624,N_39650);
xor U40101 (N_40101,N_38815,N_38830);
nand U40102 (N_40102,N_39187,N_37779);
and U40103 (N_40103,N_36601,N_39202);
and U40104 (N_40104,N_39487,N_36701);
or U40105 (N_40105,N_37492,N_35195);
nor U40106 (N_40106,N_39050,N_39726);
or U40107 (N_40107,N_36644,N_38134);
xnor U40108 (N_40108,N_37165,N_35007);
nand U40109 (N_40109,N_36874,N_38964);
and U40110 (N_40110,N_38417,N_39921);
nor U40111 (N_40111,N_37013,N_35636);
xor U40112 (N_40112,N_38406,N_39195);
nor U40113 (N_40113,N_36399,N_39078);
nand U40114 (N_40114,N_39721,N_39791);
nand U40115 (N_40115,N_39756,N_39405);
xor U40116 (N_40116,N_38639,N_38975);
nand U40117 (N_40117,N_39914,N_35617);
or U40118 (N_40118,N_37358,N_38371);
or U40119 (N_40119,N_38914,N_35054);
and U40120 (N_40120,N_39116,N_36537);
xnor U40121 (N_40121,N_35588,N_36160);
xor U40122 (N_40122,N_39986,N_37616);
nor U40123 (N_40123,N_35567,N_35240);
nand U40124 (N_40124,N_35317,N_35740);
and U40125 (N_40125,N_38221,N_35721);
nor U40126 (N_40126,N_35464,N_39249);
nand U40127 (N_40127,N_38439,N_37997);
nor U40128 (N_40128,N_35076,N_37102);
or U40129 (N_40129,N_35635,N_38863);
nor U40130 (N_40130,N_35308,N_39273);
and U40131 (N_40131,N_35509,N_37642);
nand U40132 (N_40132,N_38461,N_39038);
and U40133 (N_40133,N_35393,N_38230);
or U40134 (N_40134,N_39286,N_39442);
nand U40135 (N_40135,N_36014,N_35287);
or U40136 (N_40136,N_36524,N_37366);
xnor U40137 (N_40137,N_36597,N_38643);
and U40138 (N_40138,N_36077,N_38231);
xor U40139 (N_40139,N_35209,N_36787);
or U40140 (N_40140,N_38011,N_39617);
and U40141 (N_40141,N_38725,N_39562);
or U40142 (N_40142,N_36542,N_36925);
and U40143 (N_40143,N_39221,N_35546);
xnor U40144 (N_40144,N_38154,N_36835);
and U40145 (N_40145,N_39833,N_39216);
xor U40146 (N_40146,N_35787,N_37874);
or U40147 (N_40147,N_35877,N_39670);
xor U40148 (N_40148,N_36000,N_38541);
or U40149 (N_40149,N_38068,N_38570);
or U40150 (N_40150,N_38573,N_36506);
nand U40151 (N_40151,N_35281,N_37311);
or U40152 (N_40152,N_36564,N_37514);
nor U40153 (N_40153,N_36128,N_39878);
and U40154 (N_40154,N_35793,N_37363);
nor U40155 (N_40155,N_35250,N_39736);
nor U40156 (N_40156,N_38803,N_38973);
and U40157 (N_40157,N_36274,N_39123);
nand U40158 (N_40158,N_37671,N_37901);
or U40159 (N_40159,N_39997,N_36978);
nand U40160 (N_40160,N_39616,N_35337);
and U40161 (N_40161,N_36913,N_35694);
nand U40162 (N_40162,N_35581,N_37976);
or U40163 (N_40163,N_39830,N_38312);
nor U40164 (N_40164,N_37303,N_36334);
nand U40165 (N_40165,N_36610,N_36003);
nor U40166 (N_40166,N_38108,N_37924);
and U40167 (N_40167,N_38217,N_39524);
nand U40168 (N_40168,N_36461,N_35145);
and U40169 (N_40169,N_38252,N_36845);
nand U40170 (N_40170,N_36007,N_36640);
or U40171 (N_40171,N_37182,N_38208);
and U40172 (N_40172,N_37788,N_39855);
nand U40173 (N_40173,N_39918,N_37468);
xor U40174 (N_40174,N_36694,N_38675);
xor U40175 (N_40175,N_35728,N_37239);
nor U40176 (N_40176,N_38880,N_35395);
or U40177 (N_40177,N_38754,N_39526);
xnor U40178 (N_40178,N_38520,N_38519);
nand U40179 (N_40179,N_38606,N_35558);
or U40180 (N_40180,N_35971,N_38913);
xnor U40181 (N_40181,N_38015,N_36754);
and U40182 (N_40182,N_36885,N_38818);
nor U40183 (N_40183,N_38462,N_37194);
and U40184 (N_40184,N_37409,N_39085);
nor U40185 (N_40185,N_36513,N_36230);
or U40186 (N_40186,N_35612,N_38105);
nor U40187 (N_40187,N_37826,N_38107);
nand U40188 (N_40188,N_35548,N_37274);
or U40189 (N_40189,N_37969,N_38492);
and U40190 (N_40190,N_38269,N_35847);
and U40191 (N_40191,N_36290,N_37321);
and U40192 (N_40192,N_37320,N_36409);
xor U40193 (N_40193,N_35127,N_37342);
xnor U40194 (N_40194,N_35059,N_35514);
nand U40195 (N_40195,N_36050,N_37775);
xor U40196 (N_40196,N_35266,N_38408);
xnor U40197 (N_40197,N_35837,N_37648);
and U40198 (N_40198,N_39139,N_36327);
or U40199 (N_40199,N_38843,N_35183);
nor U40200 (N_40200,N_35247,N_36487);
nand U40201 (N_40201,N_37498,N_36367);
nand U40202 (N_40202,N_35681,N_35870);
and U40203 (N_40203,N_36591,N_36786);
nand U40204 (N_40204,N_35196,N_36291);
xnor U40205 (N_40205,N_39317,N_38524);
nor U40206 (N_40206,N_35890,N_36691);
or U40207 (N_40207,N_39185,N_35319);
or U40208 (N_40208,N_36257,N_35443);
xor U40209 (N_40209,N_37094,N_38082);
or U40210 (N_40210,N_36410,N_38767);
or U40211 (N_40211,N_35606,N_37278);
or U40212 (N_40212,N_37109,N_35353);
xnor U40213 (N_40213,N_35100,N_39895);
and U40214 (N_40214,N_35782,N_36187);
and U40215 (N_40215,N_36232,N_35487);
and U40216 (N_40216,N_35638,N_37131);
nor U40217 (N_40217,N_35419,N_35188);
xnor U40218 (N_40218,N_37679,N_39981);
and U40219 (N_40219,N_38790,N_36558);
nand U40220 (N_40220,N_39382,N_35347);
nand U40221 (N_40221,N_38587,N_36769);
or U40222 (N_40222,N_39779,N_38473);
xor U40223 (N_40223,N_39517,N_35537);
nor U40224 (N_40224,N_39138,N_38579);
xor U40225 (N_40225,N_36243,N_39033);
and U40226 (N_40226,N_39937,N_38533);
or U40227 (N_40227,N_38188,N_37685);
and U40228 (N_40228,N_38129,N_36238);
xnor U40229 (N_40229,N_35673,N_35707);
or U40230 (N_40230,N_36104,N_36272);
nor U40231 (N_40231,N_38812,N_39019);
nor U40232 (N_40232,N_35243,N_35506);
and U40233 (N_40233,N_35577,N_36553);
nor U40234 (N_40234,N_39144,N_36432);
nor U40235 (N_40235,N_35106,N_39677);
and U40236 (N_40236,N_39632,N_36414);
and U40237 (N_40237,N_36527,N_35794);
nor U40238 (N_40238,N_39312,N_36278);
or U40239 (N_40239,N_35055,N_39229);
or U40240 (N_40240,N_38680,N_38045);
nand U40241 (N_40241,N_37836,N_35743);
nor U40242 (N_40242,N_38512,N_36565);
nor U40243 (N_40243,N_35949,N_35160);
and U40244 (N_40244,N_37626,N_39759);
xor U40245 (N_40245,N_37063,N_36285);
nor U40246 (N_40246,N_37079,N_38562);
nand U40247 (N_40247,N_36357,N_37567);
or U40248 (N_40248,N_36148,N_35118);
nor U40249 (N_40249,N_38804,N_35150);
nor U40250 (N_40250,N_35500,N_37588);
nor U40251 (N_40251,N_35712,N_35073);
or U40252 (N_40252,N_38900,N_38387);
nand U40253 (N_40253,N_36783,N_37231);
xnor U40254 (N_40254,N_37371,N_35963);
or U40255 (N_40255,N_35220,N_35855);
nor U40256 (N_40256,N_35955,N_38633);
xor U40257 (N_40257,N_35024,N_38870);
or U40258 (N_40258,N_35553,N_39264);
or U40259 (N_40259,N_35872,N_37335);
and U40260 (N_40260,N_37238,N_35025);
nor U40261 (N_40261,N_39439,N_39327);
nor U40262 (N_40262,N_37686,N_39766);
nand U40263 (N_40263,N_35988,N_35415);
and U40264 (N_40264,N_36470,N_35111);
and U40265 (N_40265,N_36952,N_37756);
or U40266 (N_40266,N_35279,N_37748);
and U40267 (N_40267,N_39846,N_37908);
nand U40268 (N_40268,N_38490,N_35057);
xnor U40269 (N_40269,N_38614,N_38747);
and U40270 (N_40270,N_35138,N_38048);
and U40271 (N_40271,N_39374,N_37364);
nor U40272 (N_40272,N_36029,N_35212);
and U40273 (N_40273,N_38474,N_36094);
nand U40274 (N_40274,N_37017,N_35820);
nor U40275 (N_40275,N_39930,N_38086);
nand U40276 (N_40276,N_35267,N_39115);
nand U40277 (N_40277,N_39941,N_36185);
xnor U40278 (N_40278,N_38278,N_38619);
xnor U40279 (N_40279,N_38187,N_38356);
nand U40280 (N_40280,N_36732,N_38789);
nor U40281 (N_40281,N_36719,N_36528);
and U40282 (N_40282,N_35310,N_35392);
or U40283 (N_40283,N_36927,N_35591);
nand U40284 (N_40284,N_39148,N_37062);
and U40285 (N_40285,N_36970,N_39266);
nand U40286 (N_40286,N_39949,N_38228);
or U40287 (N_40287,N_39772,N_37055);
and U40288 (N_40288,N_39992,N_35677);
or U40289 (N_40289,N_37739,N_39534);
or U40290 (N_40290,N_37328,N_38896);
nor U40291 (N_40291,N_38243,N_36018);
or U40292 (N_40292,N_38019,N_35357);
xnor U40293 (N_40293,N_35187,N_35678);
nor U40294 (N_40294,N_35658,N_38700);
xnor U40295 (N_40295,N_39473,N_37999);
xor U40296 (N_40296,N_37898,N_37794);
nand U40297 (N_40297,N_35140,N_35552);
nor U40298 (N_40298,N_37235,N_37961);
or U40299 (N_40299,N_39268,N_36297);
nor U40300 (N_40300,N_35826,N_36270);
and U40301 (N_40301,N_39210,N_38687);
nor U40302 (N_40302,N_39121,N_37220);
or U40303 (N_40303,N_35403,N_39274);
nand U40304 (N_40304,N_38345,N_36482);
or U40305 (N_40305,N_37133,N_37499);
nor U40306 (N_40306,N_36522,N_36267);
xnor U40307 (N_40307,N_37761,N_37649);
nor U40308 (N_40308,N_36888,N_38427);
nor U40309 (N_40309,N_39716,N_36995);
and U40310 (N_40310,N_35792,N_38209);
and U40311 (N_40311,N_39365,N_37887);
xnor U40312 (N_40312,N_38906,N_35065);
nand U40313 (N_40313,N_39798,N_38165);
nand U40314 (N_40314,N_38733,N_39719);
xor U40315 (N_40315,N_39252,N_37764);
and U40316 (N_40316,N_39842,N_39776);
nor U40317 (N_40317,N_37413,N_38918);
nor U40318 (N_40318,N_37652,N_39635);
and U40319 (N_40319,N_39117,N_36634);
nand U40320 (N_40320,N_38211,N_36159);
xor U40321 (N_40321,N_39882,N_37608);
and U40322 (N_40322,N_39678,N_39602);
or U40323 (N_40323,N_39044,N_36164);
nor U40324 (N_40324,N_39111,N_38861);
nand U40325 (N_40325,N_37509,N_36818);
nand U40326 (N_40326,N_37024,N_36780);
nand U40327 (N_40327,N_36452,N_37839);
nor U40328 (N_40328,N_38442,N_39811);
or U40329 (N_40329,N_38374,N_35486);
nor U40330 (N_40330,N_38858,N_39960);
nand U40331 (N_40331,N_39886,N_37793);
xnor U40332 (N_40332,N_37272,N_35844);
or U40333 (N_40333,N_37439,N_36480);
xnor U40334 (N_40334,N_39926,N_37645);
nor U40335 (N_40335,N_36517,N_39275);
or U40336 (N_40336,N_35962,N_39692);
nor U40337 (N_40337,N_37340,N_37751);
nand U40338 (N_40338,N_35046,N_39606);
or U40339 (N_40339,N_35732,N_37404);
nor U40340 (N_40340,N_38666,N_36226);
and U40341 (N_40341,N_37438,N_37932);
and U40342 (N_40342,N_35238,N_39145);
and U40343 (N_40343,N_36448,N_35812);
xnor U40344 (N_40344,N_36262,N_39901);
and U40345 (N_40345,N_35050,N_38132);
xor U40346 (N_40346,N_38325,N_36412);
and U40347 (N_40347,N_39440,N_38398);
and U40348 (N_40348,N_37688,N_36456);
nor U40349 (N_40349,N_36075,N_39894);
nand U40350 (N_40350,N_38953,N_38544);
or U40351 (N_40351,N_37986,N_39474);
or U40352 (N_40352,N_39634,N_39159);
or U40353 (N_40353,N_36912,N_38407);
xor U40354 (N_40354,N_39100,N_37001);
xnor U40355 (N_40355,N_37500,N_35797);
nor U40356 (N_40356,N_35155,N_38043);
xor U40357 (N_40357,N_38480,N_39934);
xor U40358 (N_40358,N_36473,N_38779);
or U40359 (N_40359,N_38856,N_35502);
nand U40360 (N_40360,N_35735,N_37581);
xnor U40361 (N_40361,N_37218,N_35582);
nor U40362 (N_40362,N_39828,N_38518);
or U40363 (N_40363,N_38600,N_35058);
nor U40364 (N_40364,N_36125,N_37611);
or U40365 (N_40365,N_36551,N_35571);
xnor U40366 (N_40366,N_35460,N_36241);
or U40367 (N_40367,N_36523,N_36606);
and U40368 (N_40368,N_35072,N_38076);
and U40369 (N_40369,N_38470,N_37146);
nand U40370 (N_40370,N_36051,N_38169);
nor U40371 (N_40371,N_39970,N_39432);
nor U40372 (N_40372,N_39092,N_37115);
nor U40373 (N_40373,N_38229,N_37457);
nor U40374 (N_40374,N_38389,N_37141);
and U40375 (N_40375,N_35978,N_38218);
or U40376 (N_40376,N_36598,N_36492);
nand U40377 (N_40377,N_35153,N_39987);
nand U40378 (N_40378,N_39447,N_35147);
nand U40379 (N_40379,N_38203,N_35687);
nand U40380 (N_40380,N_39484,N_39646);
nand U40381 (N_40381,N_39430,N_38758);
xor U40382 (N_40382,N_37354,N_36881);
nor U40383 (N_40383,N_39610,N_35229);
or U40384 (N_40384,N_39137,N_39453);
nor U40385 (N_40385,N_38051,N_36814);
and U40386 (N_40386,N_39865,N_38942);
nand U40387 (N_40387,N_39998,N_39805);
or U40388 (N_40388,N_39568,N_35470);
nand U40389 (N_40389,N_38826,N_39978);
nand U40390 (N_40390,N_39276,N_39064);
and U40391 (N_40391,N_37066,N_35613);
and U40392 (N_40392,N_38359,N_38884);
xnor U40393 (N_40393,N_36911,N_39489);
nor U40394 (N_40394,N_39792,N_37797);
nand U40395 (N_40395,N_36548,N_35103);
and U40396 (N_40396,N_38664,N_36219);
or U40397 (N_40397,N_39188,N_39774);
nand U40398 (N_40398,N_37855,N_38276);
nand U40399 (N_40399,N_36063,N_36775);
nand U40400 (N_40400,N_38331,N_37444);
nor U40401 (N_40401,N_36649,N_37253);
or U40402 (N_40402,N_36115,N_39906);
or U40403 (N_40403,N_35384,N_37193);
nand U40404 (N_40404,N_39108,N_35597);
xnor U40405 (N_40405,N_35236,N_37139);
xor U40406 (N_40406,N_39032,N_37112);
or U40407 (N_40407,N_35904,N_38588);
xor U40408 (N_40408,N_39293,N_35090);
xor U40409 (N_40409,N_35587,N_39357);
or U40410 (N_40410,N_36762,N_37281);
or U40411 (N_40411,N_37978,N_37100);
nor U40412 (N_40412,N_39378,N_35302);
or U40413 (N_40413,N_37860,N_37584);
xnor U40414 (N_40414,N_38075,N_38501);
nand U40415 (N_40415,N_38934,N_36277);
nand U40416 (N_40416,N_39521,N_35718);
and U40417 (N_40417,N_35334,N_39289);
and U40418 (N_40418,N_35724,N_35562);
or U40419 (N_40419,N_38267,N_35123);
xor U40420 (N_40420,N_36580,N_36990);
or U40421 (N_40421,N_39333,N_36467);
or U40422 (N_40422,N_37279,N_39336);
or U40423 (N_40423,N_37546,N_37460);
nand U40424 (N_40424,N_38287,N_39558);
nor U40425 (N_40425,N_37891,N_35030);
nor U40426 (N_40426,N_37568,N_36503);
and U40427 (N_40427,N_38665,N_37562);
nor U40428 (N_40428,N_38277,N_35016);
or U40429 (N_40429,N_39419,N_37866);
nand U40430 (N_40430,N_39816,N_39239);
xor U40431 (N_40431,N_35888,N_38852);
xnor U40432 (N_40432,N_37244,N_35508);
and U40433 (N_40433,N_35023,N_38696);
nor U40434 (N_40434,N_39813,N_37655);
and U40435 (N_40435,N_38987,N_38049);
xnor U40436 (N_40436,N_36603,N_38311);
xor U40437 (N_40437,N_38118,N_38008);
and U40438 (N_40438,N_37657,N_38605);
nor U40439 (N_40439,N_36657,N_38364);
nor U40440 (N_40440,N_39656,N_37510);
nand U40441 (N_40441,N_35853,N_36204);
nor U40442 (N_40442,N_36544,N_36855);
and U40443 (N_40443,N_37130,N_36864);
xnor U40444 (N_40444,N_38855,N_38923);
nor U40445 (N_40445,N_39368,N_36013);
or U40446 (N_40446,N_37323,N_39283);
nand U40447 (N_40447,N_38543,N_38303);
or U40448 (N_40448,N_36950,N_36733);
and U40449 (N_40449,N_36875,N_35856);
nand U40450 (N_40450,N_37482,N_37059);
or U40451 (N_40451,N_39871,N_38613);
or U40452 (N_40452,N_36633,N_39778);
nor U40453 (N_40453,N_38199,N_37664);
nor U40454 (N_40454,N_37663,N_39152);
or U40455 (N_40455,N_38152,N_36441);
and U40456 (N_40456,N_35146,N_37540);
nand U40457 (N_40457,N_37044,N_37952);
or U40458 (N_40458,N_36022,N_37036);
and U40459 (N_40459,N_39297,N_38965);
xor U40460 (N_40460,N_36669,N_39714);
xor U40461 (N_40461,N_37089,N_38875);
or U40462 (N_40462,N_37827,N_36258);
nand U40463 (N_40463,N_39945,N_38956);
xor U40464 (N_40464,N_38095,N_38743);
xor U40465 (N_40465,N_38808,N_35533);
xnor U40466 (N_40466,N_36728,N_37283);
or U40467 (N_40467,N_37766,N_39101);
nand U40468 (N_40468,N_37099,N_38877);
and U40469 (N_40469,N_39400,N_36491);
nor U40470 (N_40470,N_35725,N_37357);
nor U40471 (N_40471,N_37774,N_39136);
nand U40472 (N_40472,N_36652,N_35373);
nor U40473 (N_40473,N_35101,N_36992);
nor U40474 (N_40474,N_36759,N_37390);
and U40475 (N_40475,N_39248,N_36433);
and U40476 (N_40476,N_38888,N_37505);
nor U40477 (N_40477,N_39463,N_37005);
nor U40478 (N_40478,N_35843,N_36585);
nand U40479 (N_40479,N_38582,N_38242);
or U40480 (N_40480,N_37951,N_38106);
nor U40481 (N_40481,N_37268,N_37796);
or U40482 (N_40482,N_35432,N_36890);
xnor U40483 (N_40483,N_36683,N_38655);
nand U40484 (N_40484,N_36102,N_38745);
xor U40485 (N_40485,N_37612,N_39796);
or U40486 (N_40486,N_35727,N_38793);
and U40487 (N_40487,N_36791,N_36302);
and U40488 (N_40488,N_37569,N_36010);
nor U40489 (N_40489,N_36996,N_37658);
nand U40490 (N_40490,N_37296,N_39310);
or U40491 (N_40491,N_38444,N_35189);
and U40492 (N_40492,N_37917,N_37786);
or U40493 (N_40493,N_37890,N_38727);
nand U40494 (N_40494,N_35859,N_38575);
or U40495 (N_40495,N_38440,N_36504);
nand U40496 (N_40496,N_37959,N_36655);
nand U40497 (N_40497,N_38977,N_36035);
or U40498 (N_40498,N_37769,N_38894);
and U40499 (N_40499,N_39782,N_39306);
nand U40500 (N_40500,N_38527,N_38098);
and U40501 (N_40501,N_39915,N_39794);
nand U40502 (N_40502,N_36709,N_37267);
xnor U40503 (N_40503,N_36109,N_35202);
xor U40504 (N_40504,N_39550,N_37844);
xor U40505 (N_40505,N_37832,N_36173);
nand U40506 (N_40506,N_36617,N_37497);
and U40507 (N_40507,N_35081,N_36514);
nand U40508 (N_40508,N_36821,N_36275);
xnor U40509 (N_40509,N_39244,N_36483);
xor U40510 (N_40510,N_35559,N_35703);
xnor U40511 (N_40511,N_37157,N_36364);
or U40512 (N_40512,N_37729,N_39868);
nor U40513 (N_40513,N_39321,N_37464);
xnor U40514 (N_40514,N_38599,N_39457);
and U40515 (N_40515,N_38400,N_39911);
nand U40516 (N_40516,N_37561,N_37129);
or U40517 (N_40517,N_38525,N_38021);
nand U40518 (N_40518,N_36011,N_36702);
xor U40519 (N_40519,N_37933,N_37177);
nor U40520 (N_40520,N_37247,N_36622);
nor U40521 (N_40521,N_38213,N_37654);
or U40522 (N_40522,N_36566,N_36449);
and U40523 (N_40523,N_38206,N_39503);
or U40524 (N_40524,N_38453,N_35771);
xor U40525 (N_40525,N_35488,N_39315);
or U40526 (N_40526,N_38678,N_38306);
and U40527 (N_40527,N_39854,N_38963);
or U40528 (N_40528,N_39931,N_39449);
or U40529 (N_40529,N_35752,N_36930);
or U40530 (N_40530,N_38185,N_37892);
nand U40531 (N_40531,N_38763,N_37515);
xor U40532 (N_40532,N_37957,N_39478);
nand U40533 (N_40533,N_38640,N_35726);
or U40534 (N_40534,N_35832,N_36895);
xor U40535 (N_40535,N_39840,N_39370);
nand U40536 (N_40536,N_35485,N_38550);
nor U40537 (N_40537,N_36203,N_36854);
or U40538 (N_40538,N_39410,N_36319);
and U40539 (N_40539,N_39544,N_36047);
or U40540 (N_40540,N_35009,N_35863);
nor U40541 (N_40541,N_35993,N_38648);
nand U40542 (N_40542,N_38872,N_37249);
xor U40543 (N_40543,N_37833,N_35950);
xor U40544 (N_40544,N_36228,N_37566);
or U40545 (N_40545,N_38198,N_35852);
nor U40546 (N_40546,N_36858,N_38566);
nand U40547 (N_40547,N_38334,N_39807);
nor U40548 (N_40548,N_36853,N_39748);
or U40549 (N_40549,N_35901,N_37542);
nand U40550 (N_40550,N_38383,N_37824);
or U40551 (N_40551,N_37299,N_39755);
nor U40552 (N_40552,N_35551,N_36176);
xor U40553 (N_40553,N_36440,N_37983);
nand U40554 (N_40554,N_39636,N_36103);
nand U40555 (N_40555,N_36917,N_38263);
xor U40556 (N_40556,N_39600,N_35167);
nor U40557 (N_40557,N_37709,N_37308);
and U40558 (N_40558,N_38632,N_39342);
nand U40559 (N_40559,N_36098,N_37302);
nand U40560 (N_40560,N_36974,N_38919);
nand U40561 (N_40561,N_38931,N_35960);
xnor U40562 (N_40562,N_35303,N_37362);
or U40563 (N_40563,N_37254,N_37644);
xor U40564 (N_40564,N_35784,N_35342);
xnor U40565 (N_40565,N_36149,N_38085);
xnor U40566 (N_40566,N_36829,N_38974);
or U40567 (N_40567,N_38433,N_36112);
nor U40568 (N_40568,N_36442,N_39902);
xnor U40569 (N_40569,N_39469,N_36040);
nand U40570 (N_40570,N_38369,N_36194);
and U40571 (N_40571,N_38580,N_38347);
or U40572 (N_40572,N_35258,N_38522);
and U40573 (N_40573,N_36348,N_37718);
or U40574 (N_40574,N_36457,N_36740);
and U40575 (N_40575,N_36065,N_36678);
nand U40576 (N_40576,N_37307,N_37852);
nand U40577 (N_40577,N_39924,N_35776);
xor U40578 (N_40578,N_38916,N_37294);
and U40579 (N_40579,N_36313,N_37212);
nand U40580 (N_40580,N_37518,N_35605);
nand U40581 (N_40581,N_38716,N_37900);
xor U40582 (N_40582,N_36172,N_36923);
xnor U40583 (N_40583,N_35555,N_38805);
nor U40584 (N_40584,N_36183,N_39788);
or U40585 (N_40585,N_38241,N_36959);
nand U40586 (N_40586,N_39711,N_36170);
and U40587 (N_40587,N_38636,N_35014);
nor U40588 (N_40588,N_35578,N_37553);
nor U40589 (N_40589,N_35799,N_35093);
or U40590 (N_40590,N_35614,N_35252);
or U40591 (N_40591,N_36929,N_35828);
and U40592 (N_40592,N_37742,N_39737);
nor U40593 (N_40593,N_38898,N_35881);
and U40594 (N_40594,N_39348,N_39879);
or U40595 (N_40595,N_36146,N_37989);
and U40596 (N_40596,N_39839,N_36190);
nor U40597 (N_40597,N_36420,N_35294);
nand U40598 (N_40598,N_37339,N_39196);
nor U40599 (N_40599,N_38403,N_38849);
or U40600 (N_40600,N_36977,N_39933);
nor U40601 (N_40601,N_39569,N_35122);
nand U40602 (N_40602,N_35857,N_35833);
and U40603 (N_40603,N_37563,N_39060);
nor U40604 (N_40604,N_38847,N_38517);
nand U40605 (N_40605,N_36967,N_37487);
nor U40606 (N_40606,N_38876,N_39674);
and U40607 (N_40607,N_39643,N_36345);
nor U40608 (N_40608,N_38646,N_35184);
xnor U40609 (N_40609,N_36700,N_38908);
or U40610 (N_40610,N_35976,N_38038);
xor U40611 (N_40611,N_39752,N_37186);
nand U40612 (N_40612,N_37064,N_37441);
xor U40613 (N_40613,N_37417,N_37293);
and U40614 (N_40614,N_35747,N_37954);
nand U40615 (N_40615,N_38983,N_36620);
and U40616 (N_40616,N_35656,N_39071);
or U40617 (N_40617,N_36301,N_37110);
nor U40618 (N_40618,N_36163,N_35616);
nand U40619 (N_40619,N_39880,N_39793);
or U40620 (N_40620,N_35417,N_36199);
and U40621 (N_40621,N_37502,N_37975);
and U40622 (N_40622,N_38530,N_35323);
or U40623 (N_40623,N_36245,N_36113);
xor U40624 (N_40624,N_36532,N_37173);
and U40625 (N_40625,N_36849,N_38094);
nor U40626 (N_40626,N_36584,N_36918);
and U40627 (N_40627,N_39039,N_36935);
or U40628 (N_40628,N_36255,N_35659);
nand U40629 (N_40629,N_39505,N_37406);
xor U40630 (N_40630,N_39860,N_38910);
xnor U40631 (N_40631,N_36559,N_36026);
nor U40632 (N_40632,N_38717,N_35702);
and U40633 (N_40633,N_38386,N_38984);
or U40634 (N_40634,N_36726,N_35943);
nand U40635 (N_40635,N_39178,N_35216);
nand U40636 (N_40636,N_35113,N_37019);
nand U40637 (N_40637,N_38264,N_36872);
and U40638 (N_40638,N_38262,N_35152);
nor U40639 (N_40639,N_35610,N_36811);
nor U40640 (N_40640,N_37937,N_38989);
xor U40641 (N_40641,N_37991,N_36322);
and U40642 (N_40642,N_37048,N_36256);
nand U40643 (N_40643,N_38191,N_35800);
xnor U40644 (N_40644,N_36496,N_35313);
nand U40645 (N_40645,N_39329,N_36227);
nor U40646 (N_40646,N_37984,N_39102);
xor U40647 (N_40647,N_39284,N_39607);
nor U40648 (N_40648,N_39750,N_37437);
or U40649 (N_40649,N_38370,N_37621);
nand U40650 (N_40650,N_38324,N_38271);
nand U40651 (N_40651,N_38031,N_38653);
and U40652 (N_40652,N_39227,N_36749);
xor U40653 (N_40653,N_36605,N_39657);
nand U40654 (N_40654,N_36001,N_38576);
or U40655 (N_40655,N_36017,N_37158);
and U40656 (N_40656,N_35503,N_35368);
nand U40657 (N_40657,N_35777,N_39120);
nand U40658 (N_40658,N_38300,N_38866);
and U40659 (N_40659,N_35010,N_37203);
nor U40660 (N_40660,N_38892,N_36903);
and U40661 (N_40661,N_38147,N_37378);
nor U40662 (N_40662,N_36295,N_37703);
and U40663 (N_40663,N_36942,N_37780);
and U40664 (N_40664,N_37585,N_36981);
nand U40665 (N_40665,N_36209,N_36096);
nand U40666 (N_40666,N_36857,N_38176);
nand U40667 (N_40667,N_37572,N_39967);
nor U40668 (N_40668,N_39034,N_38336);
and U40669 (N_40669,N_37043,N_39974);
and U40670 (N_40670,N_36436,N_37528);
or U40671 (N_40671,N_38968,N_35177);
or U40672 (N_40672,N_38484,N_38109);
xor U40673 (N_40673,N_38927,N_36915);
nand U40674 (N_40674,N_39977,N_38366);
nand U40675 (N_40675,N_35922,N_37687);
xor U40676 (N_40676,N_35637,N_39282);
and U40677 (N_40677,N_37940,N_35245);
nand U40678 (N_40678,N_35811,N_38090);
nand U40679 (N_40679,N_36798,N_39096);
xor U40680 (N_40680,N_37674,N_35965);
and U40681 (N_40681,N_38719,N_39556);
or U40682 (N_40682,N_37728,N_36676);
nor U40683 (N_40683,N_36489,N_36865);
nor U40684 (N_40684,N_37237,N_35471);
xnor U40685 (N_40685,N_37206,N_37276);
nor U40686 (N_40686,N_36856,N_39377);
or U40687 (N_40687,N_36233,N_37070);
nand U40688 (N_40688,N_36595,N_35914);
nor U40689 (N_40689,N_38783,N_35737);
xor U40690 (N_40690,N_38961,N_38377);
xor U40691 (N_40691,N_39332,N_39609);
and U40692 (N_40692,N_35554,N_38949);
nand U40693 (N_40693,N_36339,N_38339);
and U40694 (N_40694,N_39628,N_36687);
nor U40695 (N_40695,N_39943,N_38946);
nor U40696 (N_40696,N_38411,N_35742);
xnor U40697 (N_40697,N_39773,N_35312);
xor U40698 (N_40698,N_39953,N_37250);
or U40699 (N_40699,N_36807,N_38657);
nor U40700 (N_40700,N_35087,N_38445);
nor U40701 (N_40701,N_39604,N_38791);
nand U40702 (N_40702,N_38196,N_36932);
xor U40703 (N_40703,N_36156,N_35894);
xnor U40704 (N_40704,N_38756,N_39648);
and U40705 (N_40705,N_38286,N_37704);
xor U40706 (N_40706,N_35354,N_37755);
or U40707 (N_40707,N_37057,N_36625);
or U40708 (N_40708,N_39443,N_39825);
xnor U40709 (N_40709,N_39313,N_39359);
and U40710 (N_40710,N_38033,N_38479);
or U40711 (N_40711,N_37734,N_38593);
nand U40712 (N_40712,N_35505,N_38634);
xor U40713 (N_40713,N_39641,N_36810);
and U40714 (N_40714,N_36129,N_35583);
and U40715 (N_40715,N_36383,N_35037);
nand U40716 (N_40716,N_38673,N_35008);
and U40717 (N_40717,N_38124,N_39211);
nor U40718 (N_40718,N_35402,N_38222);
xnor U40719 (N_40719,N_39508,N_37749);
nor U40720 (N_40720,N_38917,N_35274);
xor U40721 (N_40721,N_38911,N_37436);
nor U40722 (N_40722,N_37741,N_39162);
nor U40723 (N_40723,N_37071,N_38732);
or U40724 (N_40724,N_39661,N_37074);
or U40725 (N_40725,N_37134,N_39920);
or U40726 (N_40726,N_37154,N_35497);
nand U40727 (N_40727,N_39486,N_36827);
and U40728 (N_40728,N_38496,N_36223);
nand U40729 (N_40729,N_37633,N_38988);
nand U40730 (N_40730,N_38215,N_35215);
nor U40731 (N_40731,N_36848,N_37124);
nor U40732 (N_40732,N_35191,N_36926);
or U40733 (N_40733,N_37108,N_35321);
nor U40734 (N_40734,N_38930,N_37440);
nor U40735 (N_40735,N_39049,N_35911);
nand U40736 (N_40736,N_35526,N_39973);
nand U40737 (N_40737,N_39361,N_35538);
nand U40738 (N_40738,N_39090,N_37705);
xor U40739 (N_40739,N_39451,N_37577);
or U40740 (N_40740,N_39080,N_38692);
and U40741 (N_40741,N_35944,N_39712);
or U40742 (N_40742,N_37910,N_37604);
and U40743 (N_40743,N_38160,N_38041);
nand U40744 (N_40744,N_38735,N_36121);
and U40745 (N_40745,N_36737,N_37230);
nand U40746 (N_40746,N_39649,N_38000);
and U40747 (N_40747,N_37907,N_37670);
and U40748 (N_40748,N_36373,N_35541);
nand U40749 (N_40749,N_39620,N_35192);
xor U40750 (N_40750,N_39222,N_36359);
nand U40751 (N_40751,N_38869,N_35969);
xnor U40752 (N_40752,N_35778,N_39968);
or U40753 (N_40753,N_38951,N_36802);
and U40754 (N_40754,N_38476,N_36546);
or U40755 (N_40755,N_39954,N_38029);
nand U40756 (N_40756,N_38955,N_36477);
and U40757 (N_40757,N_37501,N_39308);
nand U40758 (N_40758,N_37045,N_38698);
or U40759 (N_40759,N_38649,N_35455);
nor U40760 (N_40760,N_37519,N_39589);
nor U40761 (N_40761,N_35126,N_36662);
and U40762 (N_40762,N_35271,N_35091);
and U40763 (N_40763,N_37263,N_39157);
nand U40764 (N_40764,N_38873,N_36880);
nand U40765 (N_40765,N_37333,N_35224);
nand U40766 (N_40766,N_38214,N_37571);
and U40767 (N_40767,N_39859,N_36839);
nor U40768 (N_40768,N_37753,N_35835);
nor U40769 (N_40769,N_39339,N_39403);
nor U40770 (N_40770,N_39768,N_38901);
nand U40771 (N_40771,N_37018,N_38889);
xnor U40772 (N_40772,N_39826,N_36150);
or U40773 (N_40773,N_37373,N_35079);
and U40774 (N_40774,N_37516,N_37429);
xor U40775 (N_40775,N_36840,N_37977);
or U40776 (N_40776,N_39619,N_38548);
nor U40777 (N_40777,N_37521,N_37914);
xnor U40778 (N_40778,N_39820,N_35217);
or U40779 (N_40779,N_35946,N_38388);
nor U40780 (N_40780,N_35753,N_37830);
nor U40781 (N_40781,N_39498,N_38851);
or U40782 (N_40782,N_39198,N_39304);
xor U40783 (N_40783,N_38660,N_37737);
nand U40784 (N_40784,N_37309,N_38255);
nand U40785 (N_40785,N_37326,N_35275);
and U40786 (N_40786,N_37489,N_39338);
and U40787 (N_40787,N_37993,N_38455);
nor U40788 (N_40788,N_38895,N_38225);
and U40789 (N_40789,N_35322,N_36083);
xor U40790 (N_40790,N_36361,N_35549);
or U40791 (N_40791,N_35825,N_36570);
xnor U40792 (N_40792,N_35382,N_36421);
nand U40793 (N_40793,N_38357,N_35661);
nor U40794 (N_40794,N_36188,N_36736);
xor U40795 (N_40795,N_37646,N_36922);
nor U40796 (N_40796,N_38450,N_35720);
xor U40797 (N_40797,N_36613,N_38466);
xor U40798 (N_40798,N_38893,N_37968);
nor U40799 (N_40799,N_38990,N_38177);
and U40800 (N_40800,N_35596,N_38608);
nor U40801 (N_40801,N_37421,N_37798);
xnor U40802 (N_40802,N_37095,N_36973);
nand U40803 (N_40803,N_36438,N_38101);
nor U40804 (N_40804,N_39233,N_36667);
nor U40805 (N_40805,N_37472,N_39631);
and U40806 (N_40806,N_38210,N_37778);
nand U40807 (N_40807,N_37629,N_35430);
nor U40808 (N_40808,N_36988,N_37418);
nand U40809 (N_40809,N_38103,N_39169);
and U40810 (N_40810,N_37162,N_35849);
and U40811 (N_40811,N_37287,N_35830);
xor U40812 (N_40812,N_39396,N_38125);
nand U40813 (N_40813,N_36685,N_39905);
nor U40814 (N_40814,N_36501,N_35627);
nor U40815 (N_40815,N_35990,N_37153);
or U40816 (N_40816,N_38618,N_39309);
xor U40817 (N_40817,N_35754,N_37352);
xnor U40818 (N_40818,N_36600,N_37701);
xnor U40819 (N_40819,N_39020,N_35532);
xnor U40820 (N_40820,N_38155,N_35935);
nand U40821 (N_40821,N_36213,N_38583);
or U40822 (N_40822,N_35755,N_35498);
or U40823 (N_40823,N_37719,N_35595);
and U40824 (N_40824,N_38441,N_36502);
or U40825 (N_40825,N_38498,N_39022);
xnor U40826 (N_40826,N_35557,N_38452);
xnor U40827 (N_40827,N_35385,N_37428);
and U40828 (N_40828,N_38368,N_37229);
and U40829 (N_40829,N_35084,N_35149);
xor U40830 (N_40830,N_39236,N_36124);
nor U40831 (N_40831,N_38865,N_35483);
nor U40832 (N_40832,N_38776,N_35339);
and U40833 (N_40833,N_38604,N_39425);
nor U40834 (N_40834,N_39154,N_38253);
or U40835 (N_40835,N_36877,N_37122);
nor U40836 (N_40836,N_35098,N_35983);
xor U40837 (N_40837,N_38536,N_38402);
nand U40838 (N_40838,N_36423,N_36842);
xnor U40839 (N_40839,N_37828,N_39588);
and U40840 (N_40840,N_39581,N_37396);
nor U40841 (N_40841,N_39409,N_39161);
nor U40842 (N_40842,N_36611,N_35672);
xnor U40843 (N_40843,N_39493,N_35645);
nand U40844 (N_40844,N_39829,N_39398);
nand U40845 (N_40845,N_37624,N_37720);
and U40846 (N_40846,N_37330,N_36443);
and U40847 (N_40847,N_36938,N_39645);
nor U40848 (N_40848,N_37490,N_38111);
and U40849 (N_40849,N_37201,N_35651);
or U40850 (N_40850,N_38731,N_36193);
xnor U40851 (N_40851,N_38957,N_39801);
xor U40852 (N_40852,N_35186,N_36898);
and U40853 (N_40853,N_35710,N_39891);
and U40854 (N_40854,N_39935,N_39733);
nor U40855 (N_40855,N_37668,N_35880);
and U40856 (N_40856,N_35733,N_38891);
and U40857 (N_40857,N_38430,N_38239);
nand U40858 (N_40858,N_39002,N_39834);
nand U40859 (N_40859,N_39175,N_35947);
nor U40860 (N_40860,N_39366,N_35685);
xor U40861 (N_40861,N_37762,N_35414);
nand U40862 (N_40862,N_38488,N_35437);
and U40863 (N_40863,N_37121,N_35320);
or U40864 (N_40864,N_36140,N_39243);
or U40865 (N_40865,N_38868,N_37077);
xnor U40866 (N_40866,N_36266,N_35295);
and U40867 (N_40867,N_37367,N_38493);
xor U40868 (N_40868,N_39066,N_36999);
xnor U40869 (N_40869,N_35851,N_36181);
xor U40870 (N_40870,N_38943,N_35422);
or U40871 (N_40871,N_38161,N_38510);
nand U40872 (N_40872,N_38995,N_35137);
xnor U40873 (N_40873,N_36468,N_39330);
xor U40874 (N_40874,N_36020,N_37883);
or U40875 (N_40875,N_37426,N_35985);
nand U40876 (N_40876,N_35518,N_35640);
xor U40877 (N_40877,N_38742,N_38318);
or U40878 (N_40878,N_38083,N_36822);
nor U40879 (N_40879,N_37353,N_38405);
xor U40880 (N_40880,N_37763,N_37431);
and U40881 (N_40881,N_38091,N_36582);
or U40882 (N_40882,N_35306,N_35766);
or U40883 (N_40883,N_39570,N_37987);
nor U40884 (N_40884,N_36893,N_36824);
nor U40885 (N_40885,N_35064,N_36910);
or U40886 (N_40886,N_36309,N_39540);
xor U40887 (N_40887,N_37248,N_37202);
or U40888 (N_40888,N_38506,N_38136);
xor U40889 (N_40889,N_37590,N_38037);
xnor U40890 (N_40890,N_38998,N_36249);
nand U40891 (N_40891,N_38817,N_38078);
or U40892 (N_40892,N_37673,N_39220);
xnor U40893 (N_40893,N_39889,N_39373);
xnor U40894 (N_40894,N_39975,N_39519);
nor U40895 (N_40895,N_36866,N_38612);
or U40896 (N_40896,N_39126,N_36422);
nand U40897 (N_40897,N_35398,N_35958);
or U40898 (N_40898,N_36437,N_39903);
nor U40899 (N_40899,N_36378,N_39549);
nor U40900 (N_40900,N_39345,N_38741);
nor U40901 (N_40901,N_36120,N_35631);
and U40902 (N_40902,N_38394,N_36398);
or U40903 (N_40903,N_35940,N_37610);
nand U40904 (N_40904,N_35952,N_36314);
nand U40905 (N_40905,N_37049,N_38545);
and U40906 (N_40906,N_38677,N_35573);
nand U40907 (N_40907,N_37329,N_36954);
nand U40908 (N_40908,N_39392,N_35892);
or U40909 (N_40909,N_37346,N_35543);
nor U40910 (N_40910,N_36138,N_35094);
and U40911 (N_40911,N_36368,N_39751);
nand U40912 (N_40912,N_36868,N_38003);
or U40913 (N_40913,N_35006,N_37656);
nand U40914 (N_40914,N_37453,N_36186);
xnor U40915 (N_40915,N_38539,N_39292);
nand U40916 (N_40916,N_39261,N_35951);
xnor U40917 (N_40917,N_36573,N_38967);
xor U40918 (N_40918,N_35066,N_37939);
and U40919 (N_40919,N_35621,N_36237);
nor U40920 (N_40920,N_37579,N_38879);
or U40921 (N_40921,N_39206,N_38354);
xnor U40922 (N_40922,N_36039,N_36545);
nand U40923 (N_40923,N_35779,N_37190);
xor U40924 (N_40924,N_35139,N_38219);
xor U40925 (N_40925,N_39324,N_39585);
or U40926 (N_40926,N_36425,N_36965);
nand U40927 (N_40927,N_35997,N_37132);
xnor U40928 (N_40928,N_35699,N_35805);
and U40929 (N_40929,N_38712,N_39655);
nand U40930 (N_40930,N_35036,N_39929);
xor U40931 (N_40931,N_36526,N_36518);
nor U40932 (N_40932,N_35086,N_38044);
nor U40933 (N_40933,N_38346,N_39561);
nor U40934 (N_40934,N_36006,N_38449);
nand U40935 (N_40935,N_37548,N_38234);
xor U40936 (N_40936,N_37730,N_35927);
and U40937 (N_40937,N_38978,N_39271);
and U40938 (N_40938,N_38755,N_38158);
xnor U40939 (N_40939,N_35749,N_39597);
xnor U40940 (N_40940,N_36538,N_37384);
or U40941 (N_40941,N_37039,N_37348);
nand U40942 (N_40942,N_36268,N_39741);
xor U40943 (N_40943,N_36751,N_35482);
nor U40944 (N_40944,N_38066,N_36005);
and U40945 (N_40945,N_39173,N_38883);
or U40946 (N_40946,N_36725,N_35698);
nand U40947 (N_40947,N_37455,N_36049);
nor U40948 (N_40948,N_37144,N_35164);
nand U40949 (N_40949,N_37559,N_38821);
xor U40950 (N_40950,N_38175,N_39421);
nor U40951 (N_40951,N_39932,N_37615);
and U40952 (N_40952,N_36321,N_38909);
nor U40953 (N_40953,N_36292,N_37149);
or U40954 (N_40954,N_35989,N_38351);
xnor U40955 (N_40955,N_35524,N_37752);
and U40956 (N_40956,N_35501,N_37913);
and U40957 (N_40957,N_36078,N_37475);
and U40958 (N_40958,N_37034,N_39110);
or U40959 (N_40959,N_38065,N_36229);
nor U40960 (N_40960,N_39696,N_38753);
and U40961 (N_40961,N_39472,N_35012);
or U40962 (N_40962,N_35063,N_39219);
nand U40963 (N_40963,N_39654,N_38947);
xor U40964 (N_40964,N_35404,N_36239);
and U40965 (N_40965,N_38704,N_36788);
xnor U40966 (N_40966,N_38515,N_36589);
or U40967 (N_40967,N_35473,N_38690);
and U40968 (N_40968,N_35148,N_38996);
nand U40969 (N_40969,N_36777,N_36637);
xnor U40970 (N_40970,N_39477,N_35351);
and U40971 (N_40971,N_35889,N_36599);
xnor U40972 (N_40972,N_38540,N_39114);
xor U40973 (N_40973,N_35162,N_37745);
and U40974 (N_40974,N_39936,N_38723);
xor U40975 (N_40975,N_35071,N_37027);
nor U40976 (N_40976,N_35869,N_35620);
and U40977 (N_40977,N_37849,N_38059);
nand U40978 (N_40978,N_38806,N_36499);
or U40979 (N_40979,N_39151,N_38034);
or U40980 (N_40980,N_38846,N_36162);
nand U40981 (N_40981,N_35999,N_35647);
xnor U40982 (N_40982,N_37964,N_38860);
xor U40983 (N_40983,N_38596,N_38195);
nand U40984 (N_40984,N_38532,N_39051);
and U40985 (N_40985,N_36028,N_38039);
xor U40986 (N_40986,N_36365,N_35062);
nand U40987 (N_40987,N_35589,N_38323);
xor U40988 (N_40988,N_39725,N_38148);
or U40989 (N_40989,N_39350,N_38088);
or U40990 (N_40990,N_39727,N_35201);
nor U40991 (N_40991,N_39910,N_38897);
nor U40992 (N_40992,N_35325,N_36216);
and U40993 (N_40993,N_39837,N_38739);
xnor U40994 (N_40994,N_35418,N_39785);
and U40995 (N_40995,N_37189,N_38272);
xnor U40996 (N_40996,N_35848,N_35436);
and U40997 (N_40997,N_37314,N_38017);
or U40998 (N_40998,N_37573,N_37935);
or U40999 (N_40999,N_35143,N_35604);
or U41000 (N_41000,N_35774,N_39325);
or U41001 (N_41001,N_35428,N_38071);
or U41002 (N_41002,N_38785,N_36271);
nand U41003 (N_41003,N_35530,N_39724);
nor U41004 (N_41004,N_39279,N_39769);
and U41005 (N_41005,N_38294,N_39043);
xnor U41006 (N_41006,N_35982,N_35547);
and U41007 (N_41007,N_38316,N_37614);
or U41008 (N_41008,N_39518,N_35585);
xor U41009 (N_41009,N_35067,N_37923);
or U41010 (N_41010,N_38902,N_35758);
xor U41011 (N_41011,N_39731,N_38100);
nor U41012 (N_41012,N_35746,N_37551);
nand U41013 (N_41013,N_35689,N_36878);
nand U41014 (N_41014,N_37963,N_37061);
and U41015 (N_41015,N_35013,N_37277);
or U41016 (N_41016,N_37180,N_35515);
nor U41017 (N_41017,N_36572,N_38845);
xnor U41018 (N_41018,N_37355,N_39165);
nand U41019 (N_41019,N_37547,N_38113);
and U41020 (N_41020,N_39947,N_36490);
nor U41021 (N_41021,N_35507,N_36286);
or U41022 (N_41022,N_39369,N_39037);
or U41023 (N_41023,N_39058,N_36315);
nand U41024 (N_41024,N_38765,N_39909);
or U41025 (N_41025,N_36344,N_37381);
and U41026 (N_41026,N_38749,N_36876);
xnor U41027 (N_41027,N_36068,N_36638);
nand U41028 (N_41028,N_38063,N_36675);
xor U41029 (N_41029,N_37462,N_37090);
nand U41030 (N_41030,N_36666,N_37313);
nor U41031 (N_41031,N_35513,N_38820);
nor U41032 (N_41032,N_35846,N_38053);
xnor U41033 (N_41033,N_37527,N_39372);
xnor U41034 (N_41034,N_39530,N_35569);
or U41035 (N_41035,N_36031,N_36571);
xor U41036 (N_41036,N_39168,N_39000);
xor U41037 (N_41037,N_36371,N_38722);
nor U41038 (N_41038,N_39640,N_35264);
xnor U41039 (N_41039,N_35156,N_39097);
or U41040 (N_41040,N_35748,N_37955);
and U41041 (N_41041,N_38572,N_35761);
or U41042 (N_41042,N_37397,N_37641);
or U41043 (N_41043,N_37470,N_35798);
xnor U41044 (N_41044,N_36884,N_35448);
and U41045 (N_41045,N_38027,N_39323);
and U41046 (N_41046,N_37106,N_38683);
nand U41047 (N_41047,N_38651,N_36370);
or U41048 (N_41048,N_35691,N_39638);
nor U41049 (N_41049,N_38310,N_37873);
xnor U41050 (N_41050,N_39337,N_36462);
xor U41051 (N_41051,N_38642,N_36299);
xor U41052 (N_41052,N_38265,N_36293);
xnor U41053 (N_41053,N_36058,N_37700);
or U41054 (N_41054,N_37152,N_36459);
nand U41055 (N_41055,N_38289,N_37690);
and U41056 (N_41056,N_38592,N_38313);
nand U41057 (N_41057,N_39510,N_39416);
and U41058 (N_41058,N_35427,N_37262);
nand U41059 (N_41059,N_38102,N_38694);
xor U41060 (N_41060,N_35114,N_36012);
and U41061 (N_41061,N_38454,N_39415);
xor U41062 (N_41062,N_39059,N_38577);
or U41063 (N_41063,N_39946,N_35783);
nor U41064 (N_41064,N_39301,N_38617);
xor U41065 (N_41065,N_36748,N_36653);
nor U41066 (N_41066,N_37192,N_37785);
xnor U41067 (N_41067,N_35803,N_36715);
or U41068 (N_41068,N_37047,N_39448);
and U41069 (N_41069,N_37619,N_39106);
nor U41070 (N_41070,N_38864,N_39072);
and U41071 (N_41071,N_38670,N_38502);
or U41072 (N_41072,N_39506,N_35912);
nor U41073 (N_41073,N_37234,N_35966);
nor U41074 (N_41074,N_38451,N_35910);
nand U41075 (N_41075,N_36196,N_35472);
or U41076 (N_41076,N_39787,N_38322);
xnor U41077 (N_41077,N_38131,N_35343);
nor U41078 (N_41078,N_35185,N_36407);
nor U41079 (N_41079,N_35529,N_39107);
or U41080 (N_41080,N_39475,N_37650);
or U41081 (N_41081,N_37513,N_37205);
nand U41082 (N_41082,N_36629,N_37867);
nor U41083 (N_41083,N_35329,N_36046);
nand U41084 (N_41084,N_37902,N_37042);
xnor U41085 (N_41085,N_37927,N_39497);
xnor U41086 (N_41086,N_36376,N_37419);
and U41087 (N_41087,N_37713,N_35850);
nand U41088 (N_41088,N_35915,N_37715);
nor U41089 (N_41089,N_37988,N_36820);
xnor U41090 (N_41090,N_35667,N_38637);
and U41091 (N_41091,N_39939,N_35017);
or U41092 (N_41092,N_38133,N_36394);
or U41093 (N_41093,N_36349,N_38296);
nand U41094 (N_41094,N_39667,N_35244);
xor U41095 (N_41095,N_39988,N_36713);
xnor U41096 (N_41096,N_36155,N_38139);
nand U41097 (N_41097,N_39467,N_37286);
xnor U41098 (N_41098,N_39083,N_36165);
or U41099 (N_41099,N_35262,N_35356);
and U41100 (N_41100,N_38774,N_37842);
xnor U41101 (N_41101,N_35625,N_39979);
nor U41102 (N_41102,N_39679,N_35481);
nor U41103 (N_41103,N_39991,N_39514);
or U41104 (N_41104,N_35235,N_38121);
or U41105 (N_41105,N_38555,N_35981);
nand U41106 (N_41106,N_38422,N_37772);
and U41107 (N_41107,N_37862,N_37252);
or U41108 (N_41108,N_38960,N_38822);
or U41109 (N_41109,N_35104,N_36281);
nor U41110 (N_41110,N_35477,N_39984);
xor U41111 (N_41111,N_39592,N_36642);
or U41112 (N_41112,N_35845,N_36201);
nand U41113 (N_41113,N_35041,N_35957);
nor U41114 (N_41114,N_38332,N_36434);
nor U41115 (N_41115,N_35193,N_38721);
nor U41116 (N_41116,N_36785,N_38149);
xor U41117 (N_41117,N_37114,N_39408);
nand U41118 (N_41118,N_39225,N_36741);
or U41119 (N_41119,N_35544,N_36654);
and U41120 (N_41120,N_35630,N_37240);
nor U41121 (N_41121,N_36831,N_38317);
xnor U41122 (N_41122,N_35675,N_35372);
nor U41123 (N_41123,N_39166,N_38130);
xnor U41124 (N_41124,N_38467,N_39758);
nor U41125 (N_41125,N_39662,N_37481);
nand U41126 (N_41126,N_37564,N_36122);
nand U41127 (N_41127,N_36417,N_35070);
nor U41128 (N_41128,N_39200,N_38126);
nor U41129 (N_41129,N_36900,N_35080);
xor U41130 (N_41130,N_35840,N_36090);
xor U41131 (N_41131,N_35042,N_39395);
nor U41132 (N_41132,N_39515,N_37574);
and U41133 (N_41133,N_38117,N_39923);
nor U41134 (N_41134,N_38503,N_38788);
or U41135 (N_41135,N_38280,N_37038);
nor U41136 (N_41136,N_36197,N_36377);
nor U41137 (N_41137,N_38744,N_35994);
nor U41138 (N_41138,N_36215,N_38709);
or U41139 (N_41139,N_37275,N_37520);
nand U41140 (N_41140,N_36583,N_36110);
xnor U41141 (N_41141,N_38962,N_38104);
or U41142 (N_41142,N_37868,N_38330);
xnor U41143 (N_41143,N_38244,N_39030);
xnor U41144 (N_41144,N_37853,N_38882);
nor U41145 (N_41145,N_39613,N_35401);
nand U41146 (N_41146,N_35467,N_38397);
nand U41147 (N_41147,N_37447,N_36710);
nor U41148 (N_41148,N_36569,N_35525);
nor U41149 (N_41149,N_39197,N_39267);
nand U41150 (N_41150,N_38144,N_35682);
xnor U41151 (N_41151,N_38834,N_35465);
and U41152 (N_41152,N_35905,N_39231);
nor U41153 (N_41153,N_38150,N_35154);
and U41154 (N_41154,N_37389,N_36805);
xnor U41155 (N_41155,N_37990,N_39594);
xnor U41156 (N_41156,N_37743,N_38937);
nor U41157 (N_41157,N_37593,N_38991);
and U41158 (N_41158,N_38780,N_35556);
nand U41159 (N_41159,N_36887,N_37710);
and U41160 (N_41160,N_37962,N_37942);
and U41161 (N_41161,N_39951,N_38581);
nand U41162 (N_41162,N_39399,N_35141);
nor U41163 (N_41163,N_38412,N_39056);
and U41164 (N_41164,N_37773,N_36123);
nor U41165 (N_41165,N_35964,N_38658);
nand U41166 (N_41166,N_35693,N_37840);
nor U41167 (N_41167,N_39732,N_38969);
nor U41168 (N_41168,N_38933,N_36265);
or U41169 (N_41169,N_36403,N_38958);
and U41170 (N_41170,N_36289,N_38691);
nor U41171 (N_41171,N_38899,N_35251);
xnor U41172 (N_41172,N_35242,N_35061);
xor U41173 (N_41173,N_38489,N_39529);
nand U41174 (N_41174,N_39789,N_35770);
or U41175 (N_41175,N_35165,N_37298);
nand U41176 (N_41176,N_37712,N_37714);
nor U41177 (N_41177,N_37473,N_37488);
xor U41178 (N_41178,N_38950,N_35788);
nor U41179 (N_41179,N_35130,N_35674);
nand U41180 (N_41180,N_37733,N_39204);
xnor U41181 (N_41181,N_38799,N_38814);
and U41182 (N_41182,N_38752,N_38338);
and U41183 (N_41183,N_39522,N_37678);
and U41184 (N_41184,N_36411,N_37432);
xor U41185 (N_41185,N_37317,N_36485);
or U41186 (N_41186,N_35564,N_39844);
xor U41187 (N_41187,N_39363,N_36696);
nor U41188 (N_41188,N_37783,N_38077);
or U41189 (N_41189,N_37792,N_38119);
xnor U41190 (N_41190,N_37760,N_35813);
and U41191 (N_41191,N_37050,N_35730);
nor U41192 (N_41192,N_38042,N_38436);
nand U41193 (N_41193,N_35574,N_35511);
and U41194 (N_41194,N_36578,N_38784);
and U41195 (N_41195,N_36916,N_38797);
nand U41196 (N_41196,N_38654,N_38928);
nand U41197 (N_41197,N_39904,N_38122);
nor U41198 (N_41198,N_39614,N_37801);
nor U41199 (N_41199,N_39328,N_36453);
or U41200 (N_41200,N_35097,N_36086);
nand U41201 (N_41201,N_37467,N_36174);
xnor U41202 (N_41202,N_38457,N_35027);
or U41203 (N_41203,N_35223,N_39547);
nand U41204 (N_41204,N_37143,N_36782);
xnor U41205 (N_41205,N_37301,N_36355);
and U41206 (N_41206,N_39459,N_38841);
nand U41207 (N_41207,N_35775,N_36142);
nor U41208 (N_41208,N_36328,N_37884);
xor U41209 (N_41209,N_38293,N_38926);
nand U41210 (N_41210,N_38838,N_37382);
or U41211 (N_41211,N_38375,N_39352);
nand U41212 (N_41212,N_36087,N_36636);
nand U41213 (N_41213,N_35397,N_36360);
or U41214 (N_41214,N_35744,N_36730);
nor U41215 (N_41215,N_39963,N_35704);
nor U41216 (N_41216,N_39334,N_38656);
or U41217 (N_41217,N_38352,N_37814);
and U41218 (N_41218,N_37920,N_39543);
nor U41219 (N_41219,N_36795,N_39852);
nand U41220 (N_41220,N_39583,N_39956);
nand U41221 (N_41221,N_35974,N_37740);
nand U41222 (N_41222,N_38766,N_38684);
and U41223 (N_41223,N_39087,N_36846);
xor U41224 (N_41224,N_37195,N_36332);
and U41225 (N_41225,N_37950,N_39688);
and U41226 (N_41226,N_36547,N_38413);
nor U41227 (N_41227,N_37697,N_39009);
nor U41228 (N_41228,N_37434,N_38602);
nand U41229 (N_41229,N_36826,N_36933);
or U41230 (N_41230,N_39565,N_37435);
xnor U41231 (N_41231,N_39384,N_39870);
xor U41232 (N_41232,N_35657,N_39023);
or U41233 (N_41233,N_35701,N_38800);
and U41234 (N_41234,N_38114,N_37405);
nand U41235 (N_41235,N_39849,N_37944);
nand U41236 (N_41236,N_36052,N_35230);
or U41237 (N_41237,N_38465,N_35176);
nand U41238 (N_41238,N_37822,N_38871);
nand U41239 (N_41239,N_35979,N_38030);
and U41240 (N_41240,N_38542,N_35048);
nor U41241 (N_41241,N_35433,N_35499);
nand U41242 (N_41242,N_37854,N_38535);
nand U41243 (N_41243,N_37609,N_37886);
and U41244 (N_41244,N_37665,N_37214);
and U41245 (N_41245,N_36089,N_36247);
nand U41246 (N_41246,N_36269,N_37370);
nor U41247 (N_41247,N_37008,N_37172);
or U41248 (N_41248,N_36147,N_36158);
and U41249 (N_41249,N_39627,N_37531);
nand U41250 (N_41250,N_38835,N_35696);
or U41251 (N_41251,N_36906,N_38273);
and U41252 (N_41252,N_39958,N_37261);
xnor U41253 (N_41253,N_39735,N_36191);
nor U41254 (N_41254,N_36670,N_39024);
nor U41255 (N_41255,N_35411,N_35773);
nor U41256 (N_41256,N_35254,N_38288);
and U41257 (N_41257,N_37861,N_37414);
nand U41258 (N_41258,N_35615,N_39504);
nor U41259 (N_41259,N_35272,N_38853);
nor U41260 (N_41260,N_39193,N_39771);
or U41261 (N_41261,N_37463,N_38268);
xnor U41262 (N_41262,N_36520,N_36852);
or U41263 (N_41263,N_35786,N_38035);
xnor U41264 (N_41264,N_36072,N_37041);
or U41265 (N_41265,N_35391,N_36830);
and U41266 (N_41266,N_37336,N_39260);
xor U41267 (N_41267,N_35237,N_39579);
nand U41268 (N_41268,N_39464,N_38689);
nand U41269 (N_41269,N_35288,N_39622);
xor U41270 (N_41270,N_39541,N_36495);
xor U41271 (N_41271,N_37091,N_35296);
xnor U41272 (N_41272,N_35626,N_38414);
or U41273 (N_41273,N_39605,N_35956);
nor U41274 (N_41274,N_39743,N_37602);
nand U41275 (N_41275,N_36794,N_36400);
nand U41276 (N_41276,N_37622,N_37466);
nor U41277 (N_41277,N_39246,N_37260);
nand U41278 (N_41278,N_36873,N_39360);
nand U41279 (N_41279,N_36404,N_39455);
nand U41280 (N_41280,N_37236,N_38343);
nand U41281 (N_41281,N_38378,N_35038);
nand U41282 (N_41282,N_36475,N_37800);
nor U41283 (N_41283,N_36639,N_35299);
nand U41284 (N_41284,N_38250,N_35980);
or U41285 (N_41285,N_35021,N_39017);
nor U41286 (N_41286,N_35205,N_36531);
or U41287 (N_41287,N_35494,N_36500);
or U41288 (N_41288,N_38976,N_39881);
xor U41289 (N_41289,N_36326,N_39707);
xnor U41290 (N_41290,N_35535,N_37676);
xnor U41291 (N_41291,N_39761,N_39125);
and U41292 (N_41292,N_37677,N_35286);
xnor U41293 (N_41293,N_39863,N_39172);
xor U41294 (N_41294,N_37864,N_39364);
xnor U41295 (N_41295,N_36055,N_39029);
or U41296 (N_41296,N_37040,N_38904);
xor U41297 (N_41297,N_36793,N_35899);
or U41298 (N_41298,N_39669,N_38787);
and U41299 (N_41299,N_35572,N_36931);
and U41300 (N_41300,N_38014,N_39262);
or U41301 (N_41301,N_37576,N_36288);
xor U41302 (N_41302,N_35968,N_38703);
nand U41303 (N_41303,N_38796,N_35818);
and U41304 (N_41304,N_37142,N_39533);
and U41305 (N_41305,N_38459,N_39858);
or U41306 (N_41306,N_37522,N_37875);
or U41307 (N_41307,N_38380,N_38002);
nor U41308 (N_41308,N_36205,N_37266);
nand U41309 (N_41309,N_35580,N_36391);
and U41310 (N_41310,N_35865,N_38477);
nor U41311 (N_41311,N_37280,N_36166);
xnor U41312 (N_41312,N_38565,N_38256);
nand U41313 (N_41313,N_37653,N_35874);
nor U41314 (N_41314,N_35301,N_36879);
and U41315 (N_41315,N_38304,N_37549);
nand U41316 (N_41316,N_39990,N_39784);
xor U41317 (N_41317,N_36478,N_38980);
and U41318 (N_41318,N_39422,N_39940);
and U41319 (N_41319,N_35360,N_38110);
nand U41320 (N_41320,N_35434,N_37587);
and U41321 (N_41321,N_38509,N_37675);
or U41322 (N_41322,N_35860,N_39224);
or U41323 (N_41323,N_36335,N_36680);
nor U41324 (N_41324,N_38328,N_37185);
xnor U41325 (N_41325,N_36834,N_38381);
or U41326 (N_41326,N_39174,N_37485);
nand U41327 (N_41327,N_35044,N_36936);
or U41328 (N_41328,N_38672,N_35887);
or U41329 (N_41329,N_39251,N_35309);
nand U41330 (N_41330,N_38715,N_38179);
nor U41331 (N_41331,N_39513,N_38777);
xnor U41332 (N_41332,N_38390,N_38421);
nor U41333 (N_41333,N_39907,N_36445);
xnor U41334 (N_41334,N_37312,N_39128);
and U41335 (N_41335,N_39705,N_37424);
or U41336 (N_41336,N_39747,N_37680);
and U41337 (N_41337,N_36341,N_37053);
and U41338 (N_41338,N_35934,N_38275);
nor U41339 (N_41339,N_35906,N_39147);
xor U41340 (N_41340,N_38809,N_39695);
nand U41341 (N_41341,N_35492,N_39444);
or U41342 (N_41342,N_39509,N_35603);
xor U41343 (N_41343,N_35083,N_35371);
or U41344 (N_41344,N_36415,N_38434);
and U41345 (N_41345,N_36095,N_35469);
and U41346 (N_41346,N_35125,N_35823);
and U41347 (N_41347,N_39426,N_37383);
and U41348 (N_41348,N_37877,N_37031);
nor U41349 (N_41349,N_38184,N_38259);
xnor U41350 (N_41350,N_38052,N_36590);
nor U41351 (N_41351,N_38905,N_35029);
xor U41352 (N_41352,N_36130,N_37787);
and U41353 (N_41353,N_35211,N_35942);
or U41354 (N_41354,N_35416,N_36948);
and U41355 (N_41355,N_35449,N_37947);
nor U41356 (N_41356,N_39821,N_37217);
or U41357 (N_41357,N_39961,N_36914);
or U41358 (N_41358,N_38072,N_35000);
nand U41359 (N_41359,N_36030,N_37850);
or U41360 (N_41360,N_36202,N_36779);
or U41361 (N_41361,N_39353,N_38659);
or U41362 (N_41362,N_37620,N_38084);
nand U41363 (N_41363,N_38004,N_39598);
and U41364 (N_41364,N_39070,N_38925);
nand U41365 (N_41365,N_37747,N_35134);
nor U41366 (N_41366,N_39723,N_38283);
nor U41367 (N_41367,N_36464,N_35099);
nor U41368 (N_41368,N_37717,N_37398);
xnor U41369 (N_41369,N_38428,N_38178);
xor U41370 (N_41370,N_37337,N_37869);
or U41371 (N_41371,N_35124,N_35163);
nor U41372 (N_41372,N_36939,N_38291);
or U41373 (N_41373,N_35878,N_35210);
nand U41374 (N_41374,N_36705,N_37241);
nand U41375 (N_41375,N_36632,N_38813);
xor U41376 (N_41376,N_35396,N_39081);
nand U41377 (N_41377,N_35913,N_37707);
xnor U41378 (N_41378,N_39675,N_35622);
or U41379 (N_41379,N_38944,N_37511);
and U41380 (N_41380,N_35170,N_38251);
or U41381 (N_41381,N_38240,N_39103);
xor U41382 (N_41382,N_35268,N_36225);
nor U41383 (N_41383,N_38207,N_37159);
and U41384 (N_41384,N_36139,N_35697);
and U41385 (N_41385,N_36317,N_38772);
nor U41386 (N_41386,N_35219,N_39925);
and U41387 (N_41387,N_38707,N_36384);
and U41388 (N_41388,N_39205,N_38610);
or U41389 (N_41389,N_35791,N_37118);
nor U41390 (N_41390,N_39676,N_36949);
or U41391 (N_41391,N_38281,N_39008);
xor U41392 (N_41392,N_35836,N_39146);
xor U41393 (N_41393,N_39698,N_39471);
nand U41394 (N_41394,N_38140,N_35925);
xor U41395 (N_41395,N_36563,N_37119);
and U41396 (N_41396,N_35713,N_37004);
nor U41397 (N_41397,N_36817,N_35814);
nand U41398 (N_41398,N_35231,N_35954);
nor U41399 (N_41399,N_39993,N_39075);
or U41400 (N_41400,N_35117,N_39913);
and U41401 (N_41401,N_36766,N_35563);
xor U41402 (N_41402,N_35327,N_37391);
xnor U41403 (N_41403,N_38824,N_37379);
nor U41404 (N_41404,N_39441,N_36250);
or U41405 (N_41405,N_35179,N_35439);
and U41406 (N_41406,N_39468,N_37056);
nor U41407 (N_41407,N_39300,N_39192);
xnor U41408 (N_41408,N_39982,N_37906);
nand U41409 (N_41409,N_36616,N_37699);
xor U41410 (N_41410,N_37445,N_39088);
nor U41411 (N_41411,N_39851,N_39567);
xor U41412 (N_41412,N_39516,N_38190);
or U41413 (N_41413,N_36066,N_38981);
and U41414 (N_41414,N_35491,N_36847);
or U41415 (N_41415,N_35316,N_35827);
xnor U41416 (N_41416,N_37223,N_37782);
and U41417 (N_41417,N_37054,N_39672);
nand U41418 (N_41418,N_37101,N_35121);
nand U41419 (N_41419,N_35109,N_36106);
xor U41420 (N_41420,N_39603,N_36476);
nor U41421 (N_41421,N_36064,N_39827);
or U41422 (N_41422,N_38396,N_36408);
nor U41423 (N_41423,N_38220,N_37105);
or U41424 (N_41424,N_36770,N_35641);
nor U41425 (N_41425,N_39601,N_37092);
or U41426 (N_41426,N_35105,N_38999);
xnor U41427 (N_41427,N_35429,N_39311);
nor U41428 (N_41428,N_35652,N_37222);
and U41429 (N_41429,N_35256,N_39460);
or U41430 (N_41430,N_36641,N_35669);
xor U41431 (N_41431,N_35765,N_36387);
xor U41432 (N_41432,N_37325,N_39015);
and U41433 (N_41433,N_39591,N_39052);
xnor U41434 (N_41434,N_37736,N_37126);
nand U41435 (N_41435,N_38079,N_35676);
nand U41436 (N_41436,N_39890,N_35668);
xnor U41437 (N_41437,N_36175,N_36093);
xnor U41438 (N_41438,N_36964,N_35891);
and U41439 (N_41439,N_37243,N_38475);
and U41440 (N_41440,N_35377,N_39994);
or U41441 (N_41441,N_36036,N_36968);
or U41442 (N_41442,N_37233,N_39069);
xnor U41443 (N_41443,N_35722,N_38652);
or U41444 (N_41444,N_38859,N_36838);
and U41445 (N_41445,N_36366,N_39091);
or U41446 (N_41446,N_39349,N_36471);
xor U41447 (N_41447,N_38839,N_36937);
or U41448 (N_41448,N_38801,N_38662);
nor U41449 (N_41449,N_39089,N_37459);
nor U41450 (N_41450,N_39240,N_39340);
or U41451 (N_41451,N_35623,N_36100);
and U41452 (N_41452,N_35200,N_38093);
and U41453 (N_41453,N_35592,N_37164);
or U41454 (N_41454,N_35390,N_36984);
or U41455 (N_41455,N_37543,N_38770);
nor U41456 (N_41456,N_38006,N_37896);
xor U41457 (N_41457,N_37319,N_36704);
xnor U41458 (N_41458,N_39254,N_35263);
or U41459 (N_41459,N_36663,N_36135);
and U41460 (N_41460,N_39952,N_39242);
or U41461 (N_41461,N_39571,N_36560);
nor U41462 (N_41462,N_39158,N_36612);
nand U41463 (N_41463,N_37387,N_37820);
nand U41464 (N_41464,N_37808,N_37758);
xor U41465 (N_41465,N_37145,N_39433);
nor U41466 (N_41466,N_39691,N_38635);
nand U41467 (N_41467,N_37930,N_37083);
xor U41468 (N_41468,N_38393,N_37271);
and U41469 (N_41469,N_38425,N_38551);
nand U41470 (N_41470,N_36991,N_39835);
xnor U41471 (N_41471,N_36016,N_36602);
nand U41472 (N_41472,N_35173,N_35260);
and U41473 (N_41473,N_37613,N_37111);
and U41474 (N_41474,N_38333,N_35410);
nor U41475 (N_41475,N_38138,N_39001);
nand U41476 (N_41476,N_39320,N_39777);
nand U41477 (N_41477,N_37535,N_39864);
nand U41478 (N_41478,N_38628,N_39046);
nand U41479 (N_41479,N_38025,N_38391);
or U41480 (N_41480,N_36809,N_35479);
xnor U41481 (N_41481,N_39528,N_39838);
nor U41482 (N_41482,N_37805,N_35442);
xnor U41483 (N_41483,N_39438,N_37224);
nor U41484 (N_41484,N_36379,N_37306);
and U41485 (N_41485,N_35917,N_37731);
nand U41486 (N_41486,N_38050,N_38032);
and U41487 (N_41487,N_38936,N_39411);
and U41488 (N_41488,N_38945,N_35424);
xor U41489 (N_41489,N_36351,N_35047);
and U41490 (N_41490,N_37174,N_38997);
or U41491 (N_41491,N_37744,N_37334);
and U41492 (N_41492,N_36943,N_35305);
nor U41493 (N_41493,N_37076,N_38762);
nor U41494 (N_41494,N_37065,N_37804);
nor U41495 (N_41495,N_35206,N_39318);
and U41496 (N_41496,N_36987,N_37394);
xnor U41497 (N_41497,N_39270,N_37603);
xnor U41498 (N_41498,N_39584,N_39806);
or U41499 (N_41499,N_35074,N_38557);
xor U41500 (N_41500,N_39938,N_36859);
nand U41501 (N_41501,N_37215,N_38308);
and U41502 (N_41502,N_36776,N_35077);
and U41503 (N_41503,N_39140,N_36254);
or U41504 (N_41504,N_37395,N_39203);
nand U41505 (N_41505,N_39258,N_36706);
xor U41506 (N_41506,N_36727,N_39869);
and U41507 (N_41507,N_36451,N_38340);
nor U41508 (N_41508,N_36533,N_39626);
xor U41509 (N_41509,N_37881,N_38625);
and U41510 (N_41510,N_35931,N_35655);
and U41511 (N_41511,N_37635,N_35249);
nand U41512 (N_41512,N_38001,N_36356);
and U41513 (N_41513,N_39259,N_39296);
nor U41514 (N_41514,N_36658,N_35440);
xor U41515 (N_41515,N_39393,N_37086);
nand U41516 (N_41516,N_37721,N_39841);
and U41517 (N_41517,N_37080,N_37368);
nand U41518 (N_41518,N_35664,N_36521);
and U41519 (N_41519,N_38511,N_39153);
nand U41520 (N_41520,N_35089,N_37681);
or U41521 (N_41521,N_35919,N_36307);
or U41522 (N_41522,N_38903,N_35804);
xor U41523 (N_41523,N_37504,N_37332);
nand U41524 (N_41524,N_37555,N_37825);
nand U41525 (N_41525,N_36843,N_38070);
or U41526 (N_41526,N_36141,N_39790);
and U41527 (N_41527,N_39130,N_38163);
xnor U41528 (N_41528,N_39014,N_36048);
nand U41529 (N_41529,N_37726,N_37033);
or U41530 (N_41530,N_35049,N_38631);
or U41531 (N_41531,N_35190,N_39593);
xnor U41532 (N_41532,N_37784,N_35883);
nor U41533 (N_41533,N_35133,N_37858);
nor U41534 (N_41534,N_38463,N_35897);
and U41535 (N_41535,N_39720,N_39213);
nand U41536 (N_41536,N_37903,N_36427);
xnor U41537 (N_41537,N_35453,N_38335);
nand U41538 (N_41538,N_36320,N_39031);
nor U41539 (N_41539,N_36588,N_39290);
and U41540 (N_41540,N_36889,N_36813);
or U41541 (N_41541,N_37771,N_37338);
and U41542 (N_41542,N_36792,N_38429);
nor U41543 (N_41543,N_36206,N_36318);
nand U41544 (N_41544,N_37128,N_36796);
nand U41545 (N_41545,N_37067,N_37484);
and U41546 (N_41546,N_35324,N_36576);
or U41547 (N_41547,N_38232,N_35450);
or U41548 (N_41548,N_36023,N_39666);
xor U41549 (N_41549,N_37631,N_39893);
nor U41550 (N_41550,N_39356,N_36806);
nor U41551 (N_41551,N_38064,N_38811);
and U41552 (N_41552,N_37606,N_39996);
or U41553 (N_41553,N_37166,N_35734);
and U41554 (N_41554,N_35593,N_36871);
and U41555 (N_41555,N_37295,N_39762);
xor U41556 (N_41556,N_35001,N_36474);
and U41557 (N_41557,N_38235,N_38447);
or U41558 (N_41558,N_36516,N_38571);
or U41559 (N_41559,N_35854,N_38885);
or U41560 (N_41560,N_39948,N_38685);
nand U41561 (N_41561,N_37911,N_37871);
or U41562 (N_41562,N_35359,N_35466);
and U41563 (N_41563,N_38491,N_39129);
nor U41564 (N_41564,N_36426,N_38327);
xnor U41565 (N_41565,N_37273,N_39214);
nor U41566 (N_41566,N_37478,N_37560);
or U41567 (N_41567,N_39681,N_39057);
nand U41568 (N_41568,N_35642,N_39035);
or U41569 (N_41569,N_38424,N_39749);
nand U41570 (N_41570,N_38392,N_35182);
xor U41571 (N_41571,N_39595,N_37245);
xnor U41572 (N_41572,N_38423,N_36695);
xnor U41573 (N_41573,N_35446,N_38431);
xnor U41574 (N_41574,N_37536,N_37125);
xor U41575 (N_41575,N_35986,N_35654);
and U41576 (N_41576,N_36886,N_39718);
nor U41577 (N_41577,N_36444,N_37171);
and U41578 (N_41578,N_35807,N_37178);
nand U41579 (N_41579,N_39552,N_36019);
nand U41580 (N_41580,N_36062,N_35116);
and U41581 (N_41581,N_39553,N_38686);
or U41582 (N_41582,N_39795,N_35120);
and U41583 (N_41583,N_37347,N_37085);
nor U41584 (N_41584,N_35095,N_38438);
or U41585 (N_41585,N_38775,N_36723);
nand U41586 (N_41586,N_36961,N_35882);
nor U41587 (N_41587,N_37995,N_36105);
xor U41588 (N_41588,N_39689,N_35019);
nand U41589 (N_41589,N_36099,N_39966);
xor U41590 (N_41590,N_36816,N_39757);
nor U41591 (N_41591,N_37789,N_39149);
xor U41592 (N_41592,N_36192,N_37979);
nor U41593 (N_41593,N_36593,N_36708);
nor U41594 (N_41594,N_37816,N_36656);
nor U41595 (N_41595,N_36338,N_38260);
nand U41596 (N_41596,N_36828,N_37232);
nor U41597 (N_41597,N_36946,N_39199);
xnor U41598 (N_41598,N_39575,N_39744);
and U41599 (N_41599,N_35336,N_38771);
and U41600 (N_41600,N_35421,N_39223);
and U41601 (N_41601,N_37407,N_36760);
nor U41602 (N_41602,N_37967,N_39226);
nor U41603 (N_41603,N_38840,N_38615);
nor U41604 (N_41604,N_39808,N_35444);
nor U41605 (N_41605,N_35108,N_38833);
nor U41606 (N_41606,N_36747,N_36742);
and U41607 (N_41607,N_36153,N_37899);
nand U41608 (N_41608,N_38630,N_35208);
and U41609 (N_41609,N_36756,N_36717);
and U41610 (N_41610,N_37289,N_35255);
xnor U41611 (N_41611,N_36214,N_39016);
nand U41612 (N_41612,N_37454,N_37331);
xnor U41613 (N_41613,N_38363,N_37904);
nand U41614 (N_41614,N_36684,N_39435);
nor U41615 (N_41615,N_37282,N_38710);
nand U41616 (N_41616,N_36015,N_37343);
xor U41617 (N_41617,N_38005,N_39287);
xnor U41618 (N_41618,N_35331,N_35907);
nor U41619 (N_41619,N_36430,N_38641);
and U41620 (N_41620,N_38560,N_38183);
and U41621 (N_41621,N_35218,N_35474);
nand U41622 (N_41622,N_38786,N_39888);
xor U41623 (N_41623,N_36116,N_36883);
xnor U41624 (N_41624,N_38724,N_37416);
or U41625 (N_41625,N_36862,N_36405);
nor U41626 (N_41626,N_35088,N_36919);
nand U41627 (N_41627,N_39590,N_37011);
nor U41628 (N_41628,N_35729,N_35536);
nand U41629 (N_41629,N_35790,N_37000);
nor U41630 (N_41630,N_36510,N_36388);
and U41631 (N_41631,N_35328,N_39215);
nand U41632 (N_41632,N_37476,N_39305);
nor U41633 (N_41633,N_35468,N_37592);
xnor U41634 (N_41634,N_37107,N_35760);
nor U41635 (N_41635,N_35789,N_38534);
and U41636 (N_41636,N_36618,N_38040);
nor U41637 (N_41637,N_38127,N_35495);
or U41638 (N_41638,N_35346,N_39663);
and U41639 (N_41639,N_36659,N_37693);
or U41640 (N_41640,N_39599,N_36765);
or U41641 (N_41641,N_37365,N_39234);
nand U41642 (N_41642,N_36358,N_36550);
and U41643 (N_41643,N_35570,N_37926);
and U41644 (N_41644,N_35276,N_35634);
nor U41645 (N_41645,N_35885,N_38061);
and U41646 (N_41646,N_39899,N_38266);
or U41647 (N_41647,N_36920,N_35565);
xnor U41648 (N_41648,N_39786,N_38047);
nand U41649 (N_41649,N_36665,N_39269);
nand U41650 (N_41650,N_36803,N_36664);
nand U41651 (N_41651,N_38750,N_35575);
nor U41652 (N_41652,N_37722,N_39143);
nand U41653 (N_41653,N_36406,N_35738);
nor U41654 (N_41654,N_36033,N_36252);
xnor U41655 (N_41655,N_36397,N_35670);
or U41656 (N_41656,N_37324,N_37981);
or U41657 (N_41657,N_35886,N_35700);
xnor U41658 (N_41658,N_39390,N_36819);
nor U41659 (N_41659,N_35898,N_39479);
nor U41660 (N_41660,N_35527,N_37623);
or U41661 (N_41661,N_36841,N_38116);
nand U41662 (N_41662,N_35056,N_36986);
nor U41663 (N_41663,N_39652,N_37292);
or U41664 (N_41664,N_36189,N_39375);
nand U41665 (N_41665,N_38825,N_35599);
and U41666 (N_41666,N_37759,N_36529);
and U41667 (N_41667,N_35660,N_35378);
nor U41668 (N_41668,N_35918,N_38115);
xor U41669 (N_41669,N_39896,N_39861);
nand U41670 (N_41670,N_35908,N_38120);
or U41671 (N_41671,N_39615,N_38695);
and U41672 (N_41672,N_37512,N_38816);
nor U41673 (N_41673,N_35374,N_38718);
and U41674 (N_41674,N_38290,N_38504);
xor U41675 (N_41675,N_36221,N_36894);
or U41676 (N_41676,N_38180,N_36200);
nor U41677 (N_41677,N_35388,N_35520);
or U41678 (N_41678,N_38607,N_37356);
nor U41679 (N_41679,N_36212,N_37812);
xnor U41680 (N_41680,N_39067,N_37525);
and U41681 (N_41681,N_39367,N_38746);
or U41682 (N_41682,N_39170,N_39483);
or U41683 (N_41683,N_38948,N_38181);
and U41684 (N_41684,N_39989,N_36624);
or U41685 (N_41685,N_37666,N_39542);
nand U41686 (N_41686,N_38513,N_39331);
or U41687 (N_41687,N_38026,N_36673);
xor U41688 (N_41688,N_37691,N_36161);
nor U41689 (N_41689,N_37290,N_39217);
and U41690 (N_41690,N_39298,N_35680);
nor U41691 (N_41691,N_39495,N_36070);
and U41692 (N_41692,N_36008,N_39394);
or U41693 (N_41693,N_35383,N_36892);
xor U41694 (N_41694,N_39885,N_38971);
nor U41695 (N_41695,N_35706,N_36294);
nor U41696 (N_41696,N_35750,N_35817);
nor U41697 (N_41697,N_39729,N_35785);
and U41698 (N_41698,N_38985,N_36778);
xnor U41699 (N_41699,N_36279,N_39512);
or U41700 (N_41700,N_37069,N_37150);
xnor U41701 (N_41701,N_37469,N_39171);
or U41702 (N_41702,N_37809,N_35998);
and U41703 (N_41703,N_39073,N_38092);
xor U41704 (N_41704,N_38186,N_39263);
xor U41705 (N_41705,N_37496,N_36401);
xnor U41706 (N_41706,N_38384,N_38471);
xnor U41707 (N_41707,N_35051,N_38939);
and U41708 (N_41708,N_36897,N_38701);
or U41709 (N_41709,N_37427,N_38142);
and U41710 (N_41710,N_39702,N_35884);
nand U41711 (N_41711,N_35939,N_38682);
xor U41712 (N_41712,N_36182,N_38629);
and U41713 (N_41713,N_36298,N_37672);
or U41714 (N_41714,N_37068,N_35052);
or U41715 (N_41715,N_36061,N_38558);
nor U41716 (N_41716,N_39456,N_36385);
and U41717 (N_41717,N_39164,N_39754);
or U41718 (N_41718,N_38881,N_36382);
xor U41719 (N_41719,N_36389,N_35400);
and U41720 (N_41720,N_35297,N_36479);
and U41721 (N_41721,N_39815,N_36041);
nor U41722 (N_41722,N_35174,N_39247);
and U41723 (N_41723,N_38623,N_35092);
xnor U41724 (N_41724,N_37667,N_37138);
or U41725 (N_41725,N_37477,N_35408);
nor U41726 (N_41726,N_37380,N_38584);
or U41727 (N_41727,N_35484,N_36594);
nand U41728 (N_41728,N_38729,N_35510);
and U41729 (N_41729,N_36081,N_35282);
nand U41730 (N_41730,N_35228,N_37541);
and U41731 (N_41731,N_38282,N_39962);
and U41732 (N_41732,N_36337,N_39344);
nor U41733 (N_41733,N_36983,N_39068);
nand U41734 (N_41734,N_36693,N_36924);
xor U41735 (N_41735,N_36512,N_39760);
xnor U41736 (N_41736,N_37479,N_37344);
and U41737 (N_41737,N_38714,N_36746);
nand U41738 (N_41738,N_36721,N_39134);
or U41739 (N_41739,N_39303,N_37768);
or U41740 (N_41740,N_35875,N_36745);
nand U41741 (N_41741,N_37305,N_38193);
nand U41742 (N_41742,N_39401,N_38862);
nand U41743 (N_41743,N_39814,N_36324);
xor U41744 (N_41744,N_37725,N_36234);
or U41745 (N_41745,N_37974,N_36073);
or U41746 (N_41746,N_39764,N_39566);
nor U41747 (N_41747,N_38285,N_38986);
nand U41748 (N_41748,N_39680,N_37711);
xor U41749 (N_41749,N_39013,N_39351);
xor U41750 (N_41750,N_36844,N_35298);
and U41751 (N_41751,N_35144,N_36541);
xor U41752 (N_41752,N_35461,N_36958);
or U41753 (N_41753,N_39257,N_37443);
nor U41754 (N_41754,N_39983,N_36619);
xnor U41755 (N_41755,N_35806,N_37304);
and U41756 (N_41756,N_35975,N_37878);
and U41757 (N_41757,N_35291,N_36231);
nor U41758 (N_41758,N_35576,N_36424);
nand U41759 (N_41759,N_38437,N_36689);
or U41760 (N_41760,N_36833,N_35602);
xnor U41761 (N_41761,N_36901,N_36481);
nand U41762 (N_41762,N_35716,N_38069);
nand U41763 (N_41763,N_36236,N_38305);
nor U41764 (N_41764,N_35078,N_39490);
nor U41765 (N_41765,N_37351,N_37552);
or U41766 (N_41766,N_35423,N_38292);
nor U41767 (N_41767,N_36261,N_37265);
nand U41768 (N_41768,N_39857,N_39025);
or U41769 (N_41769,N_35763,N_37449);
xor U41770 (N_41770,N_39995,N_38123);
nand U41771 (N_41771,N_37360,N_39548);
or U41772 (N_41772,N_36282,N_39156);
nand U41773 (N_41773,N_37204,N_39867);
nand U41774 (N_41774,N_36363,N_36645);
xor U41775 (N_41775,N_35405,N_37888);
and U41776 (N_41776,N_39853,N_35695);
xnor U41777 (N_41777,N_35033,N_35225);
xnor U41778 (N_41778,N_39877,N_36561);
nor U41779 (N_41779,N_37087,N_38464);
xor U41780 (N_41780,N_37136,N_36870);
nand U41781 (N_41781,N_39715,N_37738);
nor U41782 (N_41782,N_35364,N_39388);
or U41783 (N_41783,N_35842,N_35178);
nor U41784 (N_41784,N_39957,N_39485);
xor U41785 (N_41785,N_36169,N_36107);
nor U41786 (N_41786,N_39884,N_37818);
nand U41787 (N_41787,N_38938,N_38781);
or U41788 (N_41788,N_36979,N_37135);
nand U41789 (N_41789,N_37037,N_39465);
nand U41790 (N_41790,N_38137,N_35349);
nand U41791 (N_41791,N_36343,N_38350);
nand U41792 (N_41792,N_39687,N_37627);
xor U41793 (N_41793,N_37167,N_37104);
xor U41794 (N_41794,N_37155,N_37526);
xor U41795 (N_41795,N_35128,N_39385);
nand U41796 (N_41796,N_36042,N_35665);
nor U41797 (N_41797,N_39201,N_36734);
nor U41798 (N_41798,N_38315,N_36447);
and U41799 (N_41799,N_39491,N_39573);
xor U41800 (N_41800,N_35011,N_36525);
nor U41801 (N_41801,N_38295,N_35767);
or U41802 (N_41802,N_35809,N_39560);
xor U41803 (N_41803,N_36353,N_39658);
and U41804 (N_41804,N_39612,N_36450);
nor U41805 (N_41805,N_36211,N_37403);
and U41806 (N_41806,N_35909,N_39965);
nand U41807 (N_41807,N_35900,N_35757);
nand U41808 (N_41808,N_39546,N_39482);
xor U41809 (N_41809,N_36738,N_39488);
nor U41810 (N_41810,N_35348,N_39190);
nand U41811 (N_41811,N_37724,N_36896);
and U41812 (N_41812,N_36154,N_39181);
nor U41813 (N_41813,N_37637,N_39810);
and U41814 (N_41814,N_35489,N_36672);
and U41815 (N_41815,N_35560,N_39578);
and U41816 (N_41816,N_36647,N_38529);
nor U41817 (N_41817,N_36108,N_38416);
and U41818 (N_41818,N_36699,N_37020);
nand U41819 (N_41819,N_36057,N_36145);
nor U41820 (N_41820,N_36439,N_37557);
or U41821 (N_41821,N_38726,N_37727);
and U41822 (N_41822,N_38212,N_37255);
nor U41823 (N_41823,N_39026,N_35769);
xnor U41824 (N_41824,N_39799,N_35151);
nor U41825 (N_41825,N_39704,N_36329);
xor U41826 (N_41826,N_38202,N_37558);
nand U41827 (N_41827,N_36681,N_37251);
nand U41828 (N_41828,N_39587,N_37010);
and U41829 (N_41829,N_37811,N_35253);
nand U41830 (N_41830,N_37915,N_36509);
or U41831 (N_41831,N_37817,N_39230);
nor U41832 (N_41832,N_36688,N_36198);
and U41833 (N_41833,N_38966,N_39639);
and U41834 (N_41834,N_35893,N_37596);
nand U41835 (N_41835,N_38734,N_37093);
nor U41836 (N_41836,N_38373,N_36045);
nor U41837 (N_41837,N_35839,N_39507);
or U41838 (N_41838,N_38358,N_39074);
nand U41839 (N_41839,N_36390,N_36428);
xor U41840 (N_41840,N_36957,N_36731);
nor U41841 (N_41841,N_37506,N_36643);
and U41842 (N_41842,N_37486,N_37909);
nor U41843 (N_41843,N_37374,N_35751);
nand U41844 (N_41844,N_37916,N_38062);
or U41845 (N_41845,N_38448,N_38993);
nand U41846 (N_41846,N_37113,N_35365);
nor U41847 (N_41847,N_39742,N_39545);
nand U41848 (N_41848,N_37259,N_38058);
nor U41849 (N_41849,N_35476,N_36815);
xor U41850 (N_41850,N_39637,N_39964);
nor U41851 (N_41851,N_38172,N_38500);
nand U41852 (N_41852,N_35315,N_38344);
xnor U41853 (N_41853,N_36539,N_35311);
nand U41854 (N_41854,N_35523,N_36891);
and U41855 (N_41855,N_36002,N_38249);
xnor U41856 (N_41856,N_39576,N_37770);
nor U41857 (N_41857,N_39160,N_36454);
nor U41858 (N_41858,N_37030,N_35376);
xor U41859 (N_41859,N_39892,N_37634);
xor U41860 (N_41860,N_35862,N_37246);
or U41861 (N_41861,N_35926,N_36998);
xor U41862 (N_41862,N_35112,N_38590);
and U41863 (N_41863,N_36118,N_37669);
and U41864 (N_41864,N_36021,N_37651);
and U41865 (N_41865,N_38456,N_37052);
and U41866 (N_41866,N_38761,N_38237);
xnor U41867 (N_41867,N_37985,N_39179);
nand U41868 (N_41868,N_39437,N_38081);
or U41869 (N_41869,N_38624,N_36562);
nand U41870 (N_41870,N_39346,N_37538);
nor U41871 (N_41871,N_36431,N_37750);
or U41872 (N_41872,N_35075,N_38248);
xnor U41873 (N_41873,N_35018,N_38982);
xnor U41874 (N_41874,N_36677,N_39406);
nor U41875 (N_41875,N_36126,N_36724);
and U41876 (N_41876,N_35921,N_38128);
or U41877 (N_41877,N_35361,N_37350);
nand U41878 (N_41878,N_38823,N_37361);
and U41879 (N_41879,N_36082,N_35930);
xnor U41880 (N_41880,N_39701,N_38223);
nor U41881 (N_41881,N_35938,N_39086);
and U41882 (N_41882,N_37082,N_37523);
and U41883 (N_41883,N_37625,N_37662);
xnor U41884 (N_41884,N_39112,N_35924);
or U41885 (N_41885,N_39142,N_39458);
or U41886 (N_41886,N_37799,N_39208);
nand U41887 (N_41887,N_39397,N_37607);
and U41888 (N_41888,N_39062,N_38337);
nand U41889 (N_41889,N_38994,N_35663);
xnor U41890 (N_41890,N_37269,N_39061);
and U41891 (N_41891,N_35034,N_37480);
nand U41892 (N_41892,N_36074,N_36244);
nor U41893 (N_41893,N_38302,N_37388);
nor U41894 (N_41894,N_37851,N_35861);
and U41895 (N_41895,N_36346,N_37698);
or U41896 (N_41896,N_37966,N_35257);
nand U41897 (N_41897,N_39856,N_38764);
xnor U41898 (N_41898,N_36300,N_39703);
nor U41899 (N_41899,N_38367,N_39511);
and U41900 (N_41900,N_39077,N_36712);
or U41901 (N_41901,N_36143,N_36540);
or U41902 (N_41902,N_39873,N_38151);
nand U41903 (N_41903,N_39623,N_39105);
nand U41904 (N_41904,N_39450,N_38153);
nor U41905 (N_41905,N_38706,N_37327);
nor U41906 (N_41906,N_38497,N_35895);
nor U41907 (N_41907,N_37960,N_37931);
and U41908 (N_41908,N_38748,N_38395);
nor U41909 (N_41909,N_37412,N_37035);
or U41910 (N_41910,N_38929,N_36682);
nand U41911 (N_41911,N_35409,N_38320);
xnor U41912 (N_41912,N_37016,N_37046);
or U41913 (N_41913,N_37643,N_37684);
xor U41914 (N_41914,N_37605,N_39007);
and U41915 (N_41915,N_36034,N_38096);
xor U41916 (N_41916,N_36908,N_39919);
nor U41917 (N_41917,N_39250,N_36180);
xnor U41918 (N_41918,N_38074,N_37889);
and U41919 (N_41919,N_35731,N_38559);
nand U41920 (N_41920,N_39502,N_37491);
xor U41921 (N_41921,N_36308,N_38361);
nand U41922 (N_41922,N_38171,N_36044);
or U41923 (N_41923,N_35002,N_35933);
or U41924 (N_41924,N_37226,N_38728);
or U41925 (N_41925,N_36850,N_36534);
nand U41926 (N_41926,N_39184,N_37014);
or U41927 (N_41927,N_38591,N_39436);
and U41928 (N_41928,N_35278,N_38197);
nor U41929 (N_41929,N_36152,N_36171);
and U41930 (N_41930,N_37918,N_36905);
and U41931 (N_41931,N_36552,N_36697);
and U41932 (N_41932,N_39535,N_37430);
or U41933 (N_41933,N_38609,N_37776);
nand U41934 (N_41934,N_37452,N_39927);
xnor U41935 (N_41935,N_36488,N_37401);
nand U41936 (N_41936,N_36784,N_39713);
xnor U41937 (N_41937,N_39307,N_39424);
or U41938 (N_41938,N_38226,N_38521);
or U41939 (N_41939,N_39831,N_35493);
xor U41940 (N_41940,N_36587,N_37137);
nor U41941 (N_41941,N_36283,N_38528);
xnor U41942 (N_41942,N_36133,N_37375);
xor U41943 (N_41943,N_36304,N_36260);
nor U41944 (N_41944,N_37003,N_37007);
nor U41945 (N_41945,N_39076,N_39413);
xor U41946 (N_41946,N_35690,N_37863);
nand U41947 (N_41947,N_35714,N_37219);
or U41948 (N_41948,N_39955,N_38819);
or U41949 (N_41949,N_38598,N_38143);
and U41950 (N_41950,N_39596,N_39241);
or U41951 (N_41951,N_36084,N_38341);
nand U41952 (N_41952,N_38531,N_38135);
nand U41953 (N_41953,N_37140,N_38556);
xor U41954 (N_41954,N_35972,N_35586);
nand U41955 (N_41955,N_35475,N_39322);
nor U41956 (N_41956,N_39470,N_38844);
xor U41957 (N_41957,N_36761,N_36092);
nor U41958 (N_41958,N_37372,N_38711);
nand U41959 (N_41959,N_36303,N_38508);
and U41960 (N_41960,N_36631,N_39180);
nand U41961 (N_41961,N_37636,N_39564);
nand U41962 (N_41962,N_36184,N_37781);
nand U41963 (N_41963,N_36507,N_38611);
or U41964 (N_41964,N_39063,N_39228);
nand U41965 (N_41965,N_37399,N_38597);
and U41966 (N_41966,N_39653,N_39010);
and U41967 (N_41967,N_37450,N_39651);
nor U41968 (N_41968,N_35107,N_38516);
nor U41969 (N_41969,N_35157,N_36997);
nand U41970 (N_41970,N_39555,N_38782);
nand U41971 (N_41971,N_37537,N_36381);
or U41972 (N_41972,N_35756,N_38055);
xor U41973 (N_41973,N_38418,N_36975);
and U41974 (N_41974,N_37591,N_39272);
and U41975 (N_41975,N_36429,N_39847);
nand U41976 (N_41976,N_36661,N_39402);
nand U41977 (N_41977,N_38245,N_38216);
nand U41978 (N_41978,N_35480,N_39775);
and U41979 (N_41979,N_36080,N_37597);
nor U41980 (N_41980,N_35135,N_36316);
nor U41981 (N_41981,N_39095,N_38810);
xor U41982 (N_41982,N_37837,N_37706);
or U41983 (N_41983,N_36330,N_35283);
nor U41984 (N_41984,N_38258,N_37843);
xnor U41985 (N_41985,N_35719,N_37857);
xnor U41986 (N_41986,N_37545,N_37369);
or U41987 (N_41987,N_39302,N_36956);
nor U41988 (N_41988,N_35967,N_39985);
xnor U41989 (N_41989,N_37170,N_39207);
xor U41990 (N_41990,N_39898,N_39872);
nand U41991 (N_41991,N_36720,N_35452);
nand U41992 (N_41992,N_39341,N_39163);
and U41993 (N_41993,N_35936,N_37209);
nor U41994 (N_41994,N_36581,N_36823);
or U41995 (N_41995,N_37088,N_35350);
and U41996 (N_41996,N_36455,N_37524);
nor U41997 (N_41997,N_35873,N_39551);
and U41998 (N_41998,N_35736,N_35961);
and U41999 (N_41999,N_36419,N_36218);
nand U42000 (N_42000,N_39708,N_37941);
or U42001 (N_42001,N_38616,N_36781);
nor U42002 (N_42002,N_37163,N_38067);
or U42003 (N_42003,N_36722,N_39186);
xnor U42004 (N_42004,N_37723,N_35838);
nor U42005 (N_42005,N_37980,N_37400);
or U42006 (N_42006,N_35937,N_37176);
nor U42007 (N_42007,N_36650,N_35110);
nand U42008 (N_42008,N_39036,N_39288);
and U42009 (N_42009,N_35594,N_37402);
nor U42010 (N_42010,N_38419,N_36743);
xor U42011 (N_42011,N_38468,N_39093);
and U42012 (N_42012,N_35032,N_36195);
xnor U42013 (N_42013,N_39874,N_39819);
nor U42014 (N_42014,N_38874,N_39150);
nor U42015 (N_42015,N_37965,N_35338);
and U42016 (N_42016,N_36264,N_38007);
nor U42017 (N_42017,N_36955,N_39812);
nand U42018 (N_42018,N_39209,N_38162);
nand U42019 (N_42019,N_35977,N_36630);
nor U42020 (N_42020,N_38060,N_39693);
xor U42021 (N_42021,N_35199,N_38757);
and U42022 (N_42022,N_38915,N_39836);
nor U42023 (N_42023,N_37618,N_37586);
or U42024 (N_42024,N_39265,N_37632);
or U42025 (N_42025,N_39462,N_37103);
xnor U42026 (N_42026,N_38935,N_35824);
nor U42027 (N_42027,N_35300,N_35344);
nor U42028 (N_42028,N_37503,N_38887);
or U42029 (N_42029,N_36386,N_36151);
or U42030 (N_42030,N_37410,N_36646);
xnor U42031 (N_42031,N_39668,N_35399);
or U42032 (N_42032,N_35318,N_37938);
xnor U42033 (N_42033,N_37458,N_39189);
and U42034 (N_42034,N_38773,N_39817);
and U42035 (N_42035,N_36774,N_37865);
or U42036 (N_42036,N_38432,N_39155);
nand U42037 (N_42037,N_39922,N_36980);
nor U42038 (N_42038,N_35456,N_37228);
nand U42039 (N_42039,N_36799,N_39850);
nand U42040 (N_42040,N_36340,N_39520);
and U42041 (N_42041,N_35375,N_35457);
nand U42042 (N_42042,N_37456,N_39976);
nand U42043 (N_42043,N_35045,N_37529);
or U42044 (N_42044,N_37795,N_35039);
xor U42045 (N_42045,N_36907,N_36596);
nand U42046 (N_42046,N_37746,N_36009);
xor U42047 (N_42047,N_36757,N_37422);
xor U42048 (N_42048,N_39630,N_39235);
or U42049 (N_42049,N_36079,N_39277);
xnor U42050 (N_42050,N_38097,N_37594);
and U42051 (N_42051,N_38174,N_36758);
xnor U42052 (N_42052,N_36660,N_35406);
or U42053 (N_42053,N_38482,N_38920);
nor U42054 (N_42054,N_39383,N_37695);
xnor U42055 (N_42055,N_35290,N_39047);
nand U42056 (N_42056,N_38603,N_37032);
xor U42057 (N_42057,N_39804,N_38443);
nand U42058 (N_42058,N_35379,N_38829);
xor U42059 (N_42059,N_38854,N_35053);
xnor U42060 (N_42060,N_38145,N_39314);
nor U42061 (N_42061,N_39055,N_39041);
xnor U42062 (N_42062,N_37123,N_37539);
or U42063 (N_42063,N_35879,N_37058);
nand U42064 (N_42064,N_35867,N_39104);
or U42065 (N_42065,N_35213,N_37208);
and U42066 (N_42066,N_39045,N_39706);
xnor U42067 (N_42067,N_36032,N_35762);
xnor U42068 (N_42068,N_37078,N_36091);
nor U42069 (N_42069,N_39004,N_35866);
and U42070 (N_42070,N_39611,N_38627);
nand U42071 (N_42071,N_36962,N_35705);
nand U42072 (N_42072,N_38674,N_39218);
xor U42073 (N_42073,N_35633,N_37876);
and U42074 (N_42074,N_37807,N_38563);
xnor U42075 (N_42075,N_35454,N_37689);
xnor U42076 (N_42076,N_36703,N_36718);
nor U42077 (N_42077,N_35550,N_39212);
nor U42078 (N_42078,N_37856,N_38020);
nor U42079 (N_42079,N_38028,N_39280);
and U42080 (N_42080,N_38564,N_36764);
nand U42081 (N_42081,N_39686,N_37148);
nand U42082 (N_42082,N_37803,N_35568);
xnor U42083 (N_42083,N_35293,N_37291);
and U42084 (N_42084,N_36463,N_36469);
nor U42085 (N_42085,N_36494,N_36902);
nor U42086 (N_42086,N_37423,N_35445);
xor U42087 (N_42087,N_39500,N_35031);
or U42088 (N_42088,N_36037,N_39527);
nand U42089 (N_42089,N_37885,N_36690);
xor U42090 (N_42090,N_39355,N_37806);
xor U42091 (N_42091,N_36627,N_38907);
nor U42092 (N_42092,N_36097,N_38204);
or U42093 (N_42093,N_36119,N_37284);
xor U42094 (N_42094,N_37316,N_36614);
nor U42095 (N_42095,N_36555,N_36224);
or U42096 (N_42096,N_35822,N_35987);
xnor U42097 (N_42097,N_35040,N_36921);
or U42098 (N_42098,N_36059,N_39797);
nand U42099 (N_42099,N_39843,N_35628);
nand U42100 (N_42100,N_37188,N_35387);
xnor U42101 (N_42101,N_35261,N_36797);
nor U42102 (N_42102,N_36934,N_37953);
xor U42103 (N_42103,N_35795,N_37386);
nand U42104 (N_42104,N_35172,N_37660);
and U42105 (N_42105,N_39525,N_37589);
or U42106 (N_42106,N_38435,N_35871);
and U42107 (N_42107,N_36458,N_37433);
or U42108 (N_42108,N_36651,N_39671);
nor U42109 (N_42109,N_39048,N_37847);
xnor U42110 (N_42110,N_37264,N_38247);
nand U42111 (N_42111,N_35129,N_35632);
nor U42112 (N_42112,N_37345,N_37735);
nand U42113 (N_42113,N_37859,N_38499);
or U42114 (N_42114,N_35198,N_38254);
xnor U42115 (N_42115,N_39006,N_38737);
or U42116 (N_42116,N_37696,N_39135);
nor U42117 (N_42117,N_38156,N_38270);
or U42118 (N_42118,N_35248,N_36393);
xor U42119 (N_42119,N_35345,N_35970);
nand U42120 (N_42120,N_37973,N_38505);
nor U42121 (N_42121,N_38979,N_36621);
nand U42122 (N_42122,N_38478,N_39428);
xor U42123 (N_42123,N_38850,N_35815);
and U42124 (N_42124,N_39335,N_35683);
nand U42125 (N_42125,N_35490,N_38828);
and U42126 (N_42126,N_39021,N_35768);
nor U42127 (N_42127,N_38848,N_38912);
xor U42128 (N_42128,N_36380,N_39823);
and U42129 (N_42129,N_36280,N_37534);
nand U42130 (N_42130,N_35609,N_39644);
and U42131 (N_42131,N_36772,N_38309);
or U42132 (N_42132,N_37012,N_35598);
and U42133 (N_42133,N_38601,N_38379);
nand U42134 (N_42134,N_37411,N_37002);
nand U42135 (N_42135,N_38549,N_37420);
xnor U42136 (N_42136,N_36575,N_38372);
xnor U42137 (N_42137,N_38552,N_37310);
nor U42138 (N_42138,N_35169,N_38360);
nand U42139 (N_42139,N_38569,N_37009);
nor U42140 (N_42140,N_38769,N_38705);
xnor U42141 (N_42141,N_37461,N_39124);
and U42142 (N_42142,N_36941,N_35522);
nor U42143 (N_42143,N_37442,N_38167);
nand U42144 (N_42144,N_38594,N_36053);
nor U42145 (N_42145,N_36635,N_35412);
or U42146 (N_42146,N_39291,N_38553);
and U42147 (N_42147,N_39690,N_35367);
xnor U42148 (N_42148,N_36043,N_37533);
xnor U42149 (N_42149,N_39848,N_39018);
and U42150 (N_42150,N_39281,N_38342);
or U42151 (N_42151,N_35772,N_38679);
or U42152 (N_42152,N_37970,N_38736);
nor U42153 (N_42153,N_38485,N_35876);
or U42154 (N_42154,N_35159,N_37471);
nor U42155 (N_42155,N_37385,N_38472);
nor U42156 (N_42156,N_38802,N_36904);
nand U42157 (N_42157,N_35381,N_37025);
nor U42158 (N_42158,N_39900,N_35545);
nor U42159 (N_42159,N_35745,N_38688);
nor U42160 (N_42160,N_37936,N_36287);
and U42161 (N_42161,N_36484,N_35370);
xnor U42162 (N_42162,N_37196,N_36716);
and U42163 (N_42163,N_38236,N_35896);
nand U42164 (N_42164,N_38730,N_37956);
and U42165 (N_42165,N_35273,N_39845);
nand U42166 (N_42166,N_36114,N_36259);
xnor U42167 (N_42167,N_38622,N_38526);
or U42168 (N_42168,N_38494,N_36982);
or U42169 (N_42169,N_39531,N_37897);
nand U42170 (N_42170,N_35903,N_38233);
or U42171 (N_42171,N_39167,N_36971);
nand U42172 (N_42172,N_36768,N_35158);
or U42173 (N_42173,N_36284,N_39094);
xnor U42174 (N_42174,N_39347,N_38697);
nor U42175 (N_42175,N_37495,N_38547);
xor U42176 (N_42176,N_39763,N_36671);
xnor U42177 (N_42177,N_35781,N_36800);
nor U42178 (N_42178,N_36395,N_39783);
xnor U42179 (N_42179,N_39722,N_35280);
xnor U42180 (N_42180,N_39586,N_36375);
or U42181 (N_42181,N_35653,N_36416);
nor U42182 (N_42182,N_38932,N_37393);
or U42183 (N_42183,N_36296,N_37315);
or U42184 (N_42184,N_39876,N_39109);
or U42185 (N_42185,N_37242,N_36711);
xor U42186 (N_42186,N_39294,N_35227);
nand U42187 (N_42187,N_38404,N_37376);
nor U42188 (N_42188,N_38514,N_36976);
or U42189 (N_42189,N_36076,N_39557);
nor U42190 (N_42190,N_39700,N_35692);
nor U42191 (N_42191,N_37415,N_35608);
nor U42192 (N_42192,N_37257,N_35358);
nor U42193 (N_42193,N_37191,N_35226);
nor U42194 (N_42194,N_36767,N_35841);
or U42195 (N_42195,N_39980,N_35973);
xor U42196 (N_42196,N_35462,N_35136);
nand U42197 (N_42197,N_39682,N_35330);
and U42198 (N_42198,N_36311,N_36837);
or U42199 (N_42199,N_35234,N_37949);
xor U42200 (N_42200,N_37116,N_36217);
and U42201 (N_42201,N_38355,N_37791);
or U42202 (N_42202,N_36220,N_36372);
or U42203 (N_42203,N_38399,N_35289);
nand U42204 (N_42204,N_36969,N_36608);
xor U42205 (N_42205,N_37821,N_36207);
nor U42206 (N_42206,N_36729,N_35600);
and U42207 (N_42207,N_35764,N_38760);
nor U42208 (N_42208,N_35197,N_36088);
or U42209 (N_42209,N_39040,N_37994);
and U42210 (N_42210,N_38009,N_35068);
and U42211 (N_42211,N_37377,N_35181);
and U42212 (N_42212,N_35834,N_38671);
or U42213 (N_42213,N_38297,N_35463);
xnor U42214 (N_42214,N_39494,N_35096);
xnor U42215 (N_42215,N_35540,N_37659);
and U42216 (N_42216,N_35941,N_35819);
and U42217 (N_42217,N_36604,N_39739);
nand U42218 (N_42218,N_36413,N_38415);
nand U42219 (N_42219,N_35496,N_37015);
xor U42220 (N_42220,N_39572,N_36882);
and U42221 (N_42221,N_37934,N_36989);
or U42222 (N_42222,N_35579,N_35333);
xor U42223 (N_42223,N_35644,N_39466);
nor U42224 (N_42224,N_39194,N_35380);
nor U42225 (N_42225,N_39745,N_35611);
nor U42226 (N_42226,N_37996,N_39376);
or U42227 (N_42227,N_36801,N_37297);
and U42228 (N_42228,N_39770,N_37151);
nor U42229 (N_42229,N_37929,N_37507);
xor U42230 (N_42230,N_35517,N_37600);
or U42231 (N_42231,N_37757,N_39238);
xor U42232 (N_42232,N_37300,N_36832);
xnor U42233 (N_42233,N_37716,N_35292);
and U42234 (N_42234,N_37982,N_35601);
or U42235 (N_42235,N_39999,N_37617);
nor U42236 (N_42236,N_39803,N_38080);
nand U42237 (N_42237,N_37517,N_35085);
and U42238 (N_42238,N_37096,N_37227);
and U42239 (N_42239,N_35335,N_39371);
xnor U42240 (N_42240,N_35639,N_36508);
or U42241 (N_42241,N_35671,N_37556);
nand U42242 (N_42242,N_39362,N_35233);
nand U42243 (N_42243,N_37117,N_38182);
nor U42244 (N_42244,N_39326,N_38205);
nand U42245 (N_42245,N_37051,N_36418);
nor U42246 (N_42246,N_38798,N_36771);
xor U42247 (N_42247,N_38693,N_38554);
and U42248 (N_42248,N_36263,N_39728);
nor U42249 (N_42249,N_39278,N_38941);
xnor U42250 (N_42250,N_37815,N_35561);
xor U42251 (N_42251,N_38647,N_35115);
and U42252 (N_42252,N_37647,N_39480);
nor U42253 (N_42253,N_37601,N_37565);
or U42254 (N_42254,N_36350,N_39387);
or U42255 (N_42255,N_38837,N_39237);
nor U42256 (N_42256,N_35953,N_36435);
xor U42257 (N_42257,N_38954,N_38992);
or U42258 (N_42258,N_38036,N_35916);
nand U42259 (N_42259,N_35119,N_39523);
and U42260 (N_42260,N_35132,N_36707);
nand U42261 (N_42261,N_36323,N_37216);
and U42262 (N_42262,N_35684,N_35142);
or U42263 (N_42263,N_38224,N_35082);
nand U42264 (N_42264,N_39959,N_37870);
and U42265 (N_42265,N_37483,N_39818);
nor U42266 (N_42266,N_36511,N_39582);
nor U42267 (N_42267,N_36056,N_37408);
and U42268 (N_42268,N_36692,N_35069);
nand U42269 (N_42269,N_39418,N_36944);
nand U42270 (N_42270,N_37210,N_39003);
and U42271 (N_42271,N_38201,N_39916);
and U42272 (N_42272,N_37692,N_37765);
xnor U42273 (N_42273,N_38759,N_37120);
and U42274 (N_42274,N_36836,N_36446);
xnor U42275 (N_42275,N_35858,N_39683);
and U42276 (N_42276,N_35519,N_35504);
nand U42277 (N_42277,N_37661,N_36567);
xnor U42278 (N_42278,N_39183,N_39928);
nand U42279 (N_42279,N_36909,N_38469);
nor U42280 (N_42280,N_36396,N_38663);
nand U42281 (N_42281,N_37256,N_35996);
or U42282 (N_42282,N_36127,N_35204);
xor U42283 (N_42283,N_36060,N_36519);
and U42284 (N_42284,N_39245,N_35194);
nor U42285 (N_42285,N_39822,N_39809);
nand U42286 (N_42286,N_36985,N_36966);
nand U42287 (N_42287,N_35542,N_39685);
nor U42288 (N_42288,N_37943,N_38713);
or U42289 (N_42289,N_37777,N_38362);
or U42290 (N_42290,N_36679,N_35284);
nor U42291 (N_42291,N_37169,N_37639);
and U42292 (N_42292,N_38668,N_38568);
xor U42293 (N_42293,N_35413,N_36460);
or U42294 (N_42294,N_38321,N_37694);
nor U42295 (N_42295,N_37448,N_38426);
nand U42296 (N_42296,N_39386,N_37127);
or U42297 (N_42297,N_39354,N_35831);
xnor U42298 (N_42298,N_35326,N_39883);
or U42299 (N_42299,N_38073,N_38589);
and U42300 (N_42300,N_36325,N_36607);
xnor U42301 (N_42301,N_35868,N_35649);
nand U42302 (N_42302,N_35458,N_36131);
and U42303 (N_42303,N_35516,N_35816);
xor U42304 (N_42304,N_39908,N_35932);
and U42305 (N_42305,N_39082,N_39131);
nor U42306 (N_42306,N_36861,N_38667);
or U42307 (N_42307,N_39027,N_36085);
nand U42308 (N_42308,N_37831,N_37682);
xor U42309 (N_42309,N_39379,N_37580);
or U42310 (N_42310,N_37081,N_35447);
nand U42311 (N_42311,N_35426,N_37168);
or U42312 (N_42312,N_39404,N_36101);
nor U42313 (N_42313,N_35180,N_39629);
and U42314 (N_42314,N_36623,N_36362);
or U42315 (N_42315,N_37098,N_39944);
xnor U42316 (N_42316,N_36027,N_38681);
xor U42317 (N_42317,N_39445,N_39912);
xor U42318 (N_42318,N_37882,N_35920);
or U42319 (N_42319,N_35864,N_36536);
xnor U42320 (N_42320,N_36136,N_36753);
xor U42321 (N_42321,N_36354,N_36117);
nand U42322 (N_42322,N_35341,N_39734);
or U42323 (N_42323,N_37285,N_35984);
xnor U42324 (N_42324,N_38921,N_38487);
or U42325 (N_42325,N_35662,N_37905);
and U42326 (N_42326,N_38832,N_38574);
or U42327 (N_42327,N_36331,N_36025);
xnor U42328 (N_42328,N_39647,N_35802);
xor U42329 (N_42329,N_39391,N_39950);
nor U42330 (N_42330,N_37835,N_39554);
nor U42331 (N_42331,N_35020,N_38959);
xnor U42332 (N_42332,N_38778,N_36773);
or U42333 (N_42333,N_39740,N_38495);
nor U42334 (N_42334,N_36867,N_38561);
and U42335 (N_42335,N_35646,N_36273);
nand U42336 (N_42336,N_39537,N_35277);
xor U42337 (N_42337,N_38141,N_39642);
or U42338 (N_42338,N_37072,N_35528);
or U42339 (N_42339,N_39414,N_35821);
nand U42340 (N_42340,N_37425,N_38146);
and U42341 (N_42341,N_35959,N_39412);
nand U42342 (N_42342,N_37073,N_36940);
or U42343 (N_42343,N_37465,N_38326);
nand U42344 (N_42344,N_36586,N_39538);
nor U42345 (N_42345,N_38022,N_36210);
and U42346 (N_42346,N_35304,N_39099);
nand U42347 (N_42347,N_39113,N_38200);
and U42348 (N_42348,N_35992,N_37023);
and U42349 (N_42349,N_36069,N_37790);
nand U42350 (N_42350,N_38940,N_38261);
nor U42351 (N_42351,N_36179,N_36515);
or U42352 (N_42352,N_37708,N_38023);
and U42353 (N_42353,N_39753,N_38585);
and U42354 (N_42354,N_39832,N_39407);
nand U42355 (N_42355,N_39709,N_37493);
or U42356 (N_42356,N_35207,N_38348);
and U42357 (N_42357,N_37599,N_38595);
nand U42358 (N_42358,N_37595,N_38329);
or U42359 (N_42359,N_38702,N_35717);
or U42360 (N_42360,N_38720,N_39299);
nand U42361 (N_42361,N_38057,N_36392);
xnor U42362 (N_42362,N_39012,N_39499);
xnor U42363 (N_42363,N_38018,N_38365);
and U42364 (N_42364,N_37841,N_39232);
nand U42365 (N_42365,N_35438,N_39665);
nor U42366 (N_42366,N_38166,N_39343);
and U42367 (N_42367,N_38586,N_35629);
nand U42368 (N_42368,N_38046,N_35478);
xnor U42369 (N_42369,N_37921,N_37322);
nor U42370 (N_42370,N_35923,N_39765);
or U42371 (N_42371,N_38189,N_38010);
or U42372 (N_42372,N_37530,N_36486);
and U42373 (N_42373,N_35711,N_38708);
xor U42374 (N_42374,N_38795,N_36556);
nand U42375 (N_42375,N_35902,N_38164);
or U42376 (N_42376,N_39496,N_39079);
xor U42377 (N_42377,N_39717,N_36972);
xor U42378 (N_42378,N_39897,N_35307);
and U42379 (N_42379,N_35715,N_35810);
xnor U42380 (N_42380,N_39380,N_36568);
nor U42381 (N_42381,N_35166,N_39053);
nand U42382 (N_42382,N_35232,N_37912);
or U42383 (N_42383,N_38238,N_35214);
nor U42384 (N_42384,N_35928,N_36310);
nor U42385 (N_42385,N_39481,N_38227);
nand U42386 (N_42386,N_39011,N_37895);
nand U42387 (N_42387,N_36024,N_36869);
or U42388 (N_42388,N_38972,N_35332);
and U42389 (N_42389,N_37211,N_35780);
nand U42390 (N_42390,N_39176,N_38867);
xor U42391 (N_42391,N_37998,N_36157);
nor U42392 (N_42392,N_37880,N_35004);
nand U42393 (N_42393,N_35314,N_39800);
nand U42394 (N_42394,N_39673,N_35708);
nor U42395 (N_42395,N_38089,N_38274);
nand U42396 (N_42396,N_36253,N_35948);
xor U42397 (N_42397,N_39065,N_35929);
nor U42398 (N_42398,N_36178,N_39621);
nor U42399 (N_42399,N_38012,N_38307);
and U42400 (N_42400,N_37474,N_38170);
or U42401 (N_42401,N_35648,N_37848);
nor U42402 (N_42402,N_36336,N_36615);
or U42403 (N_42403,N_38836,N_39710);
nor U42404 (N_42404,N_37823,N_35366);
nor U42405 (N_42405,N_35739,N_36342);
xnor U42406 (N_42406,N_37179,N_37160);
nand U42407 (N_42407,N_38924,N_38013);
or U42408 (N_42408,N_37258,N_39624);
xnor U42409 (N_42409,N_36860,N_38661);
nor U42410 (N_42410,N_37359,N_35171);
nor U42411 (N_42411,N_37767,N_38621);
nor U42412 (N_42412,N_37922,N_38157);
nor U42413 (N_42413,N_39319,N_38112);
or U42414 (N_42414,N_36851,N_35945);
nor U42415 (N_42415,N_36993,N_39389);
nor U42416 (N_42416,N_35531,N_37187);
xnor U42417 (N_42417,N_35168,N_39420);
nand U42418 (N_42418,N_35590,N_39559);
and U42419 (N_42419,N_37060,N_38385);
nor U42420 (N_42420,N_37845,N_37550);
or U42421 (N_42421,N_38546,N_38645);
nand U42422 (N_42422,N_35512,N_35285);
nand U42423 (N_42423,N_38087,N_36963);
nor U42424 (N_42424,N_38831,N_35796);
and U42425 (N_42425,N_38890,N_39694);
and U42426 (N_42426,N_35741,N_36374);
or U42427 (N_42427,N_35619,N_38578);
nand U42428 (N_42428,N_38699,N_36144);
nand U42429 (N_42429,N_36674,N_39972);
or U42430 (N_42430,N_37810,N_36953);
and U42431 (N_42431,N_36577,N_37992);
nor U42432 (N_42432,N_37270,N_38056);
nand U42433 (N_42433,N_37147,N_39122);
or U42434 (N_42434,N_37554,N_38246);
or U42435 (N_42435,N_38768,N_35584);
nor U42436 (N_42436,N_38353,N_39423);
nand U42437 (N_42437,N_39942,N_37198);
nand U42438 (N_42438,N_39028,N_39191);
and U42439 (N_42439,N_37341,N_37022);
and U42440 (N_42440,N_37288,N_35005);
xor U42441 (N_42441,N_38460,N_37075);
and U42442 (N_42442,N_37508,N_38279);
xnor U42443 (N_42443,N_36472,N_35340);
xor U42444 (N_42444,N_38669,N_37683);
xnor U42445 (N_42445,N_35679,N_39084);
or U42446 (N_42446,N_36493,N_39697);
nor U42447 (N_42447,N_35709,N_35394);
xnor U42448 (N_42448,N_38376,N_38299);
xnor U42449 (N_42449,N_37225,N_36306);
xor U42450 (N_42450,N_36242,N_36312);
xnor U42451 (N_42451,N_35459,N_38319);
or U42452 (N_42452,N_38878,N_39492);
and U42453 (N_42453,N_39539,N_37006);
and U42454 (N_42454,N_35362,N_37819);
and U42455 (N_42455,N_35435,N_39501);
nand U42456 (N_42456,N_39969,N_37156);
xnor U42457 (N_42457,N_38827,N_37948);
nand U42458 (N_42458,N_36755,N_38738);
nand U42459 (N_42459,N_38952,N_39446);
and U42460 (N_42460,N_39536,N_36543);
nand U42461 (N_42461,N_39417,N_36208);
nor U42462 (N_42462,N_36592,N_37846);
nand U42463 (N_42463,N_37919,N_39177);
and U42464 (N_42464,N_36668,N_36498);
or U42465 (N_42465,N_36790,N_38314);
nand U42466 (N_42466,N_36251,N_38257);
nor U42467 (N_42467,N_38349,N_35431);
nand U42468 (N_42468,N_38194,N_37318);
or U42469 (N_42469,N_39608,N_39454);
or U42470 (N_42470,N_35015,N_36054);
xor U42471 (N_42471,N_39054,N_35808);
or U42472 (N_42472,N_35028,N_39633);
nand U42473 (N_42473,N_36038,N_39746);
and U42474 (N_42474,N_36132,N_39780);
and U42475 (N_42475,N_39285,N_37021);
xor U42476 (N_42476,N_35759,N_36789);
nand U42477 (N_42477,N_38168,N_35666);
nor U42478 (N_42478,N_37834,N_36945);
or U42479 (N_42479,N_35175,N_37732);
nand U42480 (N_42480,N_39256,N_38792);
nand U42481 (N_42481,N_38537,N_35259);
xnor U42482 (N_42482,N_37640,N_39381);
xnor U42483 (N_42483,N_39427,N_38024);
and U42484 (N_42484,N_35221,N_37221);
nor U42485 (N_42485,N_38481,N_35369);
and U42486 (N_42486,N_35451,N_36111);
nor U42487 (N_42487,N_36825,N_38857);
nor U42488 (N_42488,N_37802,N_39577);
nor U42489 (N_42489,N_38794,N_38409);
and U42490 (N_42490,N_39434,N_35420);
or U42491 (N_42491,N_35363,N_36628);
or U42492 (N_42492,N_37029,N_38638);
nor U42493 (N_42493,N_36465,N_36951);
and U42494 (N_42494,N_39141,N_39118);
nor U42495 (N_42495,N_37181,N_39767);
nand U42496 (N_42496,N_36863,N_36402);
xor U42497 (N_42497,N_37582,N_38483);
nor U42498 (N_42498,N_38446,N_35241);
and U42499 (N_42499,N_36134,N_35425);
xnor U42500 (N_42500,N_35792,N_39709);
or U42501 (N_42501,N_38098,N_35794);
or U42502 (N_42502,N_39522,N_36095);
xnor U42503 (N_42503,N_38914,N_39325);
nor U42504 (N_42504,N_37441,N_39157);
xnor U42505 (N_42505,N_38959,N_35505);
nand U42506 (N_42506,N_35834,N_37991);
nand U42507 (N_42507,N_35366,N_37958);
xor U42508 (N_42508,N_37844,N_35892);
or U42509 (N_42509,N_37523,N_38664);
xnor U42510 (N_42510,N_35725,N_35277);
and U42511 (N_42511,N_37000,N_38998);
and U42512 (N_42512,N_39925,N_37315);
nor U42513 (N_42513,N_36981,N_36239);
and U42514 (N_42514,N_38296,N_39014);
and U42515 (N_42515,N_38612,N_39516);
nor U42516 (N_42516,N_35440,N_36572);
nand U42517 (N_42517,N_37247,N_36447);
nand U42518 (N_42518,N_39604,N_38796);
nand U42519 (N_42519,N_38377,N_37275);
nor U42520 (N_42520,N_36453,N_39958);
and U42521 (N_42521,N_36366,N_36393);
and U42522 (N_42522,N_37928,N_36376);
and U42523 (N_42523,N_35501,N_38272);
nor U42524 (N_42524,N_38279,N_35919);
or U42525 (N_42525,N_36721,N_37979);
and U42526 (N_42526,N_35346,N_36254);
nor U42527 (N_42527,N_36875,N_38626);
nand U42528 (N_42528,N_39007,N_39896);
nand U42529 (N_42529,N_37573,N_35798);
or U42530 (N_42530,N_39836,N_36048);
and U42531 (N_42531,N_39807,N_35710);
xnor U42532 (N_42532,N_38365,N_38782);
nand U42533 (N_42533,N_35232,N_37857);
and U42534 (N_42534,N_39615,N_36311);
xor U42535 (N_42535,N_38203,N_36893);
or U42536 (N_42536,N_39639,N_36701);
and U42537 (N_42537,N_37840,N_36407);
and U42538 (N_42538,N_36828,N_38308);
xor U42539 (N_42539,N_37206,N_37168);
and U42540 (N_42540,N_37710,N_35236);
nor U42541 (N_42541,N_38013,N_35418);
and U42542 (N_42542,N_35416,N_38995);
and U42543 (N_42543,N_36227,N_39518);
and U42544 (N_42544,N_38603,N_36633);
xor U42545 (N_42545,N_38020,N_38181);
and U42546 (N_42546,N_35781,N_35264);
or U42547 (N_42547,N_36372,N_36145);
xor U42548 (N_42548,N_38358,N_36200);
nor U42549 (N_42549,N_37058,N_39410);
and U42550 (N_42550,N_38737,N_39734);
nor U42551 (N_42551,N_35045,N_35414);
xor U42552 (N_42552,N_36610,N_36459);
and U42553 (N_42553,N_37668,N_38964);
nand U42554 (N_42554,N_35822,N_39381);
or U42555 (N_42555,N_37908,N_37524);
xor U42556 (N_42556,N_35187,N_37480);
nor U42557 (N_42557,N_38332,N_36674);
xor U42558 (N_42558,N_38478,N_36507);
nand U42559 (N_42559,N_36101,N_38999);
nor U42560 (N_42560,N_35450,N_35858);
nand U42561 (N_42561,N_36531,N_39528);
nand U42562 (N_42562,N_38327,N_39056);
and U42563 (N_42563,N_36824,N_35194);
xnor U42564 (N_42564,N_39029,N_37506);
or U42565 (N_42565,N_38244,N_35673);
nand U42566 (N_42566,N_39243,N_38036);
xor U42567 (N_42567,N_35761,N_35465);
nor U42568 (N_42568,N_35373,N_38565);
or U42569 (N_42569,N_38618,N_37508);
xor U42570 (N_42570,N_39370,N_38571);
and U42571 (N_42571,N_36992,N_38965);
or U42572 (N_42572,N_38336,N_36469);
nand U42573 (N_42573,N_38656,N_36504);
or U42574 (N_42574,N_36975,N_36959);
xor U42575 (N_42575,N_37309,N_39102);
nand U42576 (N_42576,N_39392,N_38007);
nand U42577 (N_42577,N_37850,N_36101);
or U42578 (N_42578,N_39037,N_37913);
and U42579 (N_42579,N_37348,N_35810);
nand U42580 (N_42580,N_37143,N_38574);
nor U42581 (N_42581,N_39928,N_37920);
and U42582 (N_42582,N_39147,N_37746);
and U42583 (N_42583,N_37471,N_36827);
xor U42584 (N_42584,N_35088,N_37970);
xor U42585 (N_42585,N_36453,N_38296);
nand U42586 (N_42586,N_37127,N_38437);
and U42587 (N_42587,N_38319,N_39870);
xnor U42588 (N_42588,N_37361,N_39453);
or U42589 (N_42589,N_35591,N_38277);
nor U42590 (N_42590,N_36159,N_36198);
xnor U42591 (N_42591,N_39671,N_38903);
nand U42592 (N_42592,N_37386,N_38305);
and U42593 (N_42593,N_35537,N_39635);
and U42594 (N_42594,N_36222,N_39287);
nor U42595 (N_42595,N_36319,N_36305);
and U42596 (N_42596,N_39409,N_36469);
xnor U42597 (N_42597,N_38366,N_36357);
nand U42598 (N_42598,N_38011,N_35716);
nand U42599 (N_42599,N_35117,N_35827);
nor U42600 (N_42600,N_36508,N_37859);
xor U42601 (N_42601,N_36170,N_38146);
and U42602 (N_42602,N_36370,N_38785);
xor U42603 (N_42603,N_36469,N_37573);
xnor U42604 (N_42604,N_39873,N_37705);
and U42605 (N_42605,N_39533,N_38614);
and U42606 (N_42606,N_36259,N_39333);
nor U42607 (N_42607,N_36585,N_36234);
xor U42608 (N_42608,N_35762,N_35964);
xnor U42609 (N_42609,N_36528,N_36282);
and U42610 (N_42610,N_36343,N_36884);
nand U42611 (N_42611,N_36609,N_37004);
nor U42612 (N_42612,N_36577,N_39480);
nor U42613 (N_42613,N_36125,N_38695);
nand U42614 (N_42614,N_38360,N_35981);
nand U42615 (N_42615,N_37160,N_36045);
xnor U42616 (N_42616,N_38144,N_38840);
xor U42617 (N_42617,N_37020,N_37886);
and U42618 (N_42618,N_36160,N_36751);
and U42619 (N_42619,N_37133,N_39209);
nor U42620 (N_42620,N_36739,N_37601);
nor U42621 (N_42621,N_37544,N_38820);
and U42622 (N_42622,N_36164,N_35531);
nand U42623 (N_42623,N_35840,N_37763);
nand U42624 (N_42624,N_38287,N_35925);
nand U42625 (N_42625,N_38639,N_37493);
nand U42626 (N_42626,N_36511,N_36596);
xor U42627 (N_42627,N_35403,N_39772);
and U42628 (N_42628,N_36877,N_35421);
nor U42629 (N_42629,N_38751,N_36333);
xnor U42630 (N_42630,N_38337,N_38576);
or U42631 (N_42631,N_35569,N_37852);
xnor U42632 (N_42632,N_39962,N_39767);
or U42633 (N_42633,N_37345,N_39645);
xor U42634 (N_42634,N_37769,N_38054);
and U42635 (N_42635,N_37989,N_35791);
and U42636 (N_42636,N_39232,N_36225);
nor U42637 (N_42637,N_39949,N_37293);
or U42638 (N_42638,N_38524,N_39756);
nor U42639 (N_42639,N_37294,N_35698);
nand U42640 (N_42640,N_38437,N_39756);
nand U42641 (N_42641,N_35486,N_36235);
and U42642 (N_42642,N_36174,N_39122);
nand U42643 (N_42643,N_38642,N_36798);
nor U42644 (N_42644,N_36575,N_39133);
and U42645 (N_42645,N_39455,N_38834);
xnor U42646 (N_42646,N_39016,N_37627);
nor U42647 (N_42647,N_37023,N_37199);
nor U42648 (N_42648,N_37155,N_39787);
or U42649 (N_42649,N_36957,N_36309);
and U42650 (N_42650,N_36290,N_36738);
and U42651 (N_42651,N_37144,N_35430);
nor U42652 (N_42652,N_39736,N_36101);
nand U42653 (N_42653,N_36440,N_38630);
nor U42654 (N_42654,N_37533,N_36810);
and U42655 (N_42655,N_37449,N_37894);
nand U42656 (N_42656,N_36312,N_35506);
xnor U42657 (N_42657,N_36667,N_36811);
nor U42658 (N_42658,N_39955,N_39060);
or U42659 (N_42659,N_39390,N_39059);
nand U42660 (N_42660,N_38374,N_39807);
nor U42661 (N_42661,N_35723,N_39697);
xnor U42662 (N_42662,N_39706,N_37192);
and U42663 (N_42663,N_37382,N_39310);
and U42664 (N_42664,N_38653,N_38436);
or U42665 (N_42665,N_39264,N_37977);
nor U42666 (N_42666,N_36787,N_39851);
nand U42667 (N_42667,N_36499,N_39776);
nand U42668 (N_42668,N_37350,N_36109);
or U42669 (N_42669,N_39256,N_39816);
nor U42670 (N_42670,N_38118,N_36674);
and U42671 (N_42671,N_35601,N_36160);
nand U42672 (N_42672,N_36126,N_38874);
nor U42673 (N_42673,N_35931,N_35822);
nor U42674 (N_42674,N_37034,N_36989);
or U42675 (N_42675,N_38531,N_36967);
nand U42676 (N_42676,N_39660,N_35459);
or U42677 (N_42677,N_37153,N_39745);
nand U42678 (N_42678,N_36411,N_39703);
or U42679 (N_42679,N_38727,N_38396);
or U42680 (N_42680,N_37611,N_37299);
or U42681 (N_42681,N_36642,N_38548);
and U42682 (N_42682,N_37739,N_38401);
nor U42683 (N_42683,N_37628,N_35277);
xnor U42684 (N_42684,N_36940,N_38351);
nor U42685 (N_42685,N_37128,N_37370);
or U42686 (N_42686,N_36640,N_38793);
xnor U42687 (N_42687,N_38727,N_36113);
and U42688 (N_42688,N_35019,N_37003);
and U42689 (N_42689,N_36056,N_38208);
or U42690 (N_42690,N_39755,N_35171);
xor U42691 (N_42691,N_39955,N_38728);
nand U42692 (N_42692,N_36484,N_35523);
and U42693 (N_42693,N_39719,N_37776);
xnor U42694 (N_42694,N_36745,N_35211);
or U42695 (N_42695,N_38518,N_35188);
or U42696 (N_42696,N_39091,N_37481);
nand U42697 (N_42697,N_36331,N_39848);
xnor U42698 (N_42698,N_37829,N_35044);
nand U42699 (N_42699,N_37954,N_36501);
nand U42700 (N_42700,N_35047,N_39425);
or U42701 (N_42701,N_36726,N_36780);
or U42702 (N_42702,N_38957,N_37849);
xnor U42703 (N_42703,N_37777,N_35993);
nor U42704 (N_42704,N_38909,N_37640);
or U42705 (N_42705,N_35899,N_37057);
or U42706 (N_42706,N_39454,N_36624);
and U42707 (N_42707,N_36044,N_37325);
nor U42708 (N_42708,N_37165,N_39642);
xnor U42709 (N_42709,N_38069,N_35854);
or U42710 (N_42710,N_37747,N_37615);
xnor U42711 (N_42711,N_38685,N_39823);
xnor U42712 (N_42712,N_37283,N_38076);
xor U42713 (N_42713,N_37550,N_35936);
nor U42714 (N_42714,N_37028,N_37272);
and U42715 (N_42715,N_39455,N_39178);
nand U42716 (N_42716,N_37334,N_38680);
xor U42717 (N_42717,N_39762,N_39196);
xnor U42718 (N_42718,N_38320,N_38468);
or U42719 (N_42719,N_37045,N_36952);
xor U42720 (N_42720,N_37502,N_36237);
nor U42721 (N_42721,N_38633,N_37060);
nor U42722 (N_42722,N_38558,N_37892);
or U42723 (N_42723,N_37816,N_35027);
nor U42724 (N_42724,N_39522,N_39495);
or U42725 (N_42725,N_39291,N_35971);
or U42726 (N_42726,N_35872,N_38314);
and U42727 (N_42727,N_39051,N_36622);
xnor U42728 (N_42728,N_35518,N_38099);
nor U42729 (N_42729,N_39093,N_35473);
xor U42730 (N_42730,N_35625,N_37748);
and U42731 (N_42731,N_37614,N_38162);
nand U42732 (N_42732,N_39202,N_38858);
nand U42733 (N_42733,N_37806,N_36679);
nand U42734 (N_42734,N_38032,N_39658);
nor U42735 (N_42735,N_39087,N_37444);
and U42736 (N_42736,N_36272,N_38536);
and U42737 (N_42737,N_35900,N_35872);
nand U42738 (N_42738,N_35269,N_36032);
nor U42739 (N_42739,N_35352,N_37633);
xnor U42740 (N_42740,N_39688,N_37778);
or U42741 (N_42741,N_39725,N_39569);
or U42742 (N_42742,N_38287,N_35918);
nand U42743 (N_42743,N_37013,N_39016);
xnor U42744 (N_42744,N_39497,N_36727);
or U42745 (N_42745,N_35995,N_35072);
nor U42746 (N_42746,N_38034,N_36112);
xor U42747 (N_42747,N_35897,N_37139);
nand U42748 (N_42748,N_35454,N_35993);
nand U42749 (N_42749,N_39416,N_35160);
or U42750 (N_42750,N_38650,N_38464);
nand U42751 (N_42751,N_37449,N_37049);
nor U42752 (N_42752,N_38651,N_38003);
and U42753 (N_42753,N_39357,N_38157);
or U42754 (N_42754,N_35822,N_39972);
xnor U42755 (N_42755,N_36414,N_38239);
nor U42756 (N_42756,N_38954,N_38944);
nor U42757 (N_42757,N_36233,N_39286);
or U42758 (N_42758,N_35939,N_36854);
and U42759 (N_42759,N_37483,N_38112);
nor U42760 (N_42760,N_35570,N_38795);
nand U42761 (N_42761,N_38797,N_38076);
nand U42762 (N_42762,N_39299,N_36092);
xnor U42763 (N_42763,N_39009,N_35861);
or U42764 (N_42764,N_35838,N_36754);
or U42765 (N_42765,N_35482,N_37283);
and U42766 (N_42766,N_36381,N_35272);
xnor U42767 (N_42767,N_35820,N_38344);
or U42768 (N_42768,N_35253,N_37271);
and U42769 (N_42769,N_35257,N_36447);
xnor U42770 (N_42770,N_35515,N_35612);
nor U42771 (N_42771,N_36043,N_38658);
and U42772 (N_42772,N_35746,N_37145);
or U42773 (N_42773,N_37749,N_35078);
and U42774 (N_42774,N_38705,N_36208);
and U42775 (N_42775,N_38215,N_35098);
xnor U42776 (N_42776,N_36994,N_39874);
or U42777 (N_42777,N_35833,N_36663);
or U42778 (N_42778,N_38827,N_38758);
nand U42779 (N_42779,N_38905,N_36795);
and U42780 (N_42780,N_37807,N_35978);
nand U42781 (N_42781,N_37798,N_38773);
nor U42782 (N_42782,N_36619,N_39936);
nand U42783 (N_42783,N_39498,N_39508);
nor U42784 (N_42784,N_36769,N_35136);
or U42785 (N_42785,N_37264,N_37624);
or U42786 (N_42786,N_39712,N_39114);
nor U42787 (N_42787,N_39616,N_36679);
or U42788 (N_42788,N_38975,N_39108);
nand U42789 (N_42789,N_37233,N_36981);
xor U42790 (N_42790,N_37560,N_36525);
or U42791 (N_42791,N_35119,N_36111);
and U42792 (N_42792,N_35771,N_36191);
or U42793 (N_42793,N_36253,N_39340);
or U42794 (N_42794,N_39946,N_38690);
or U42795 (N_42795,N_36032,N_39293);
and U42796 (N_42796,N_38416,N_39660);
xor U42797 (N_42797,N_35072,N_36589);
nor U42798 (N_42798,N_37754,N_36001);
xnor U42799 (N_42799,N_39416,N_36935);
and U42800 (N_42800,N_39091,N_39578);
and U42801 (N_42801,N_37531,N_39686);
or U42802 (N_42802,N_36230,N_38509);
nor U42803 (N_42803,N_39608,N_37219);
nand U42804 (N_42804,N_38268,N_39098);
xnor U42805 (N_42805,N_35183,N_35631);
xor U42806 (N_42806,N_37339,N_35116);
or U42807 (N_42807,N_36559,N_36977);
nand U42808 (N_42808,N_39784,N_37379);
nor U42809 (N_42809,N_39611,N_36169);
or U42810 (N_42810,N_38131,N_35016);
nand U42811 (N_42811,N_37540,N_39783);
nand U42812 (N_42812,N_39370,N_39818);
and U42813 (N_42813,N_36547,N_37448);
or U42814 (N_42814,N_36305,N_39095);
xnor U42815 (N_42815,N_36577,N_37804);
or U42816 (N_42816,N_39235,N_37896);
and U42817 (N_42817,N_39457,N_38898);
nor U42818 (N_42818,N_35746,N_35281);
or U42819 (N_42819,N_39415,N_39573);
nand U42820 (N_42820,N_37737,N_39022);
xor U42821 (N_42821,N_39022,N_38797);
nor U42822 (N_42822,N_37475,N_36968);
or U42823 (N_42823,N_37746,N_38390);
xor U42824 (N_42824,N_36005,N_37384);
xnor U42825 (N_42825,N_38682,N_37887);
nand U42826 (N_42826,N_38950,N_35838);
nor U42827 (N_42827,N_37665,N_36262);
or U42828 (N_42828,N_38914,N_37283);
nand U42829 (N_42829,N_39386,N_36187);
xor U42830 (N_42830,N_39485,N_39791);
xor U42831 (N_42831,N_39610,N_35143);
and U42832 (N_42832,N_39568,N_37035);
or U42833 (N_42833,N_35021,N_35253);
xnor U42834 (N_42834,N_39004,N_36084);
or U42835 (N_42835,N_38023,N_38987);
xor U42836 (N_42836,N_39922,N_38747);
xor U42837 (N_42837,N_37491,N_38111);
xnor U42838 (N_42838,N_35307,N_36745);
or U42839 (N_42839,N_39165,N_36809);
or U42840 (N_42840,N_36612,N_36369);
or U42841 (N_42841,N_37292,N_39459);
nand U42842 (N_42842,N_36104,N_37093);
xnor U42843 (N_42843,N_37736,N_38946);
nor U42844 (N_42844,N_36299,N_36909);
nor U42845 (N_42845,N_38266,N_39304);
nor U42846 (N_42846,N_38936,N_37189);
nand U42847 (N_42847,N_35455,N_37373);
nand U42848 (N_42848,N_38689,N_37670);
or U42849 (N_42849,N_37339,N_38046);
nand U42850 (N_42850,N_37276,N_39369);
and U42851 (N_42851,N_37676,N_35428);
nor U42852 (N_42852,N_38463,N_36816);
xor U42853 (N_42853,N_36218,N_36189);
and U42854 (N_42854,N_35953,N_39122);
and U42855 (N_42855,N_39382,N_38241);
and U42856 (N_42856,N_35362,N_38371);
or U42857 (N_42857,N_35943,N_39608);
and U42858 (N_42858,N_35582,N_36250);
nor U42859 (N_42859,N_38965,N_36025);
and U42860 (N_42860,N_39292,N_38300);
nor U42861 (N_42861,N_39459,N_39933);
nand U42862 (N_42862,N_37659,N_37575);
and U42863 (N_42863,N_37353,N_36031);
nor U42864 (N_42864,N_35388,N_37120);
or U42865 (N_42865,N_36341,N_38718);
nor U42866 (N_42866,N_36458,N_36146);
or U42867 (N_42867,N_37126,N_39963);
nand U42868 (N_42868,N_37893,N_36679);
nor U42869 (N_42869,N_37868,N_36966);
xor U42870 (N_42870,N_36785,N_36600);
or U42871 (N_42871,N_37447,N_38575);
nor U42872 (N_42872,N_35191,N_35273);
xnor U42873 (N_42873,N_36988,N_35226);
nor U42874 (N_42874,N_38791,N_35619);
and U42875 (N_42875,N_35117,N_39018);
nand U42876 (N_42876,N_36355,N_38121);
nor U42877 (N_42877,N_38914,N_39441);
nand U42878 (N_42878,N_39852,N_38963);
and U42879 (N_42879,N_37099,N_35843);
and U42880 (N_42880,N_39106,N_38670);
or U42881 (N_42881,N_36462,N_37633);
and U42882 (N_42882,N_37617,N_36909);
and U42883 (N_42883,N_38394,N_35614);
and U42884 (N_42884,N_36180,N_35861);
and U42885 (N_42885,N_35870,N_38096);
and U42886 (N_42886,N_39904,N_39833);
and U42887 (N_42887,N_35568,N_35411);
nand U42888 (N_42888,N_39218,N_37851);
nand U42889 (N_42889,N_37329,N_35772);
nor U42890 (N_42890,N_39791,N_39853);
and U42891 (N_42891,N_36973,N_36188);
nand U42892 (N_42892,N_37836,N_37213);
or U42893 (N_42893,N_35263,N_37826);
nand U42894 (N_42894,N_39154,N_37301);
xnor U42895 (N_42895,N_37244,N_36554);
nor U42896 (N_42896,N_37452,N_37557);
or U42897 (N_42897,N_37544,N_35724);
nand U42898 (N_42898,N_39588,N_36246);
or U42899 (N_42899,N_37360,N_35120);
and U42900 (N_42900,N_37831,N_39026);
nor U42901 (N_42901,N_39244,N_35034);
nor U42902 (N_42902,N_35074,N_39601);
nor U42903 (N_42903,N_39247,N_39147);
nand U42904 (N_42904,N_37889,N_36470);
nor U42905 (N_42905,N_39017,N_38925);
nor U42906 (N_42906,N_38776,N_36107);
xnor U42907 (N_42907,N_35670,N_37299);
nor U42908 (N_42908,N_37722,N_37700);
nor U42909 (N_42909,N_39774,N_38490);
and U42910 (N_42910,N_35709,N_36576);
and U42911 (N_42911,N_37408,N_35745);
xnor U42912 (N_42912,N_38246,N_39889);
nor U42913 (N_42913,N_38293,N_38261);
nor U42914 (N_42914,N_38752,N_39662);
or U42915 (N_42915,N_37053,N_35014);
and U42916 (N_42916,N_35148,N_37962);
and U42917 (N_42917,N_36907,N_36024);
nor U42918 (N_42918,N_39117,N_35798);
xor U42919 (N_42919,N_35490,N_37298);
and U42920 (N_42920,N_35820,N_35030);
and U42921 (N_42921,N_38209,N_36727);
xnor U42922 (N_42922,N_39506,N_36863);
and U42923 (N_42923,N_38955,N_35521);
xor U42924 (N_42924,N_35197,N_38183);
nand U42925 (N_42925,N_36218,N_39472);
xnor U42926 (N_42926,N_38802,N_37506);
nand U42927 (N_42927,N_38360,N_39899);
nand U42928 (N_42928,N_36091,N_36921);
or U42929 (N_42929,N_37266,N_39203);
or U42930 (N_42930,N_37857,N_39268);
or U42931 (N_42931,N_38427,N_37308);
nand U42932 (N_42932,N_37139,N_38324);
xnor U42933 (N_42933,N_35438,N_38932);
nor U42934 (N_42934,N_38760,N_35556);
or U42935 (N_42935,N_35798,N_39830);
nor U42936 (N_42936,N_39211,N_37419);
and U42937 (N_42937,N_38218,N_36698);
xor U42938 (N_42938,N_35761,N_39322);
or U42939 (N_42939,N_37541,N_36497);
nand U42940 (N_42940,N_35215,N_37963);
or U42941 (N_42941,N_36903,N_37129);
nand U42942 (N_42942,N_37352,N_36033);
nor U42943 (N_42943,N_39121,N_37323);
and U42944 (N_42944,N_39308,N_39166);
nand U42945 (N_42945,N_38084,N_35469);
or U42946 (N_42946,N_36407,N_35070);
and U42947 (N_42947,N_35212,N_38621);
and U42948 (N_42948,N_37537,N_36876);
or U42949 (N_42949,N_36648,N_38914);
nor U42950 (N_42950,N_36067,N_35658);
xor U42951 (N_42951,N_35755,N_39840);
or U42952 (N_42952,N_35479,N_39539);
and U42953 (N_42953,N_39819,N_35822);
nor U42954 (N_42954,N_38457,N_36166);
nand U42955 (N_42955,N_38749,N_37536);
nor U42956 (N_42956,N_35895,N_35478);
or U42957 (N_42957,N_37606,N_35931);
xnor U42958 (N_42958,N_36305,N_36700);
nor U42959 (N_42959,N_35199,N_35024);
or U42960 (N_42960,N_38728,N_37417);
xnor U42961 (N_42961,N_39638,N_39467);
nor U42962 (N_42962,N_37077,N_37803);
and U42963 (N_42963,N_38523,N_35779);
nor U42964 (N_42964,N_36135,N_39285);
xnor U42965 (N_42965,N_38697,N_39860);
nand U42966 (N_42966,N_39503,N_38908);
nand U42967 (N_42967,N_36678,N_35315);
nand U42968 (N_42968,N_39537,N_36353);
nand U42969 (N_42969,N_37800,N_38444);
or U42970 (N_42970,N_38867,N_38240);
xor U42971 (N_42971,N_37270,N_37212);
nor U42972 (N_42972,N_35505,N_37999);
nor U42973 (N_42973,N_39903,N_35253);
or U42974 (N_42974,N_39149,N_39443);
or U42975 (N_42975,N_39256,N_35465);
or U42976 (N_42976,N_39363,N_37433);
xor U42977 (N_42977,N_37743,N_35432);
xor U42978 (N_42978,N_37872,N_38930);
nand U42979 (N_42979,N_38314,N_39069);
xnor U42980 (N_42980,N_39947,N_35146);
or U42981 (N_42981,N_36291,N_37959);
nor U42982 (N_42982,N_37424,N_35270);
nor U42983 (N_42983,N_38435,N_38852);
nor U42984 (N_42984,N_37741,N_36397);
nor U42985 (N_42985,N_36163,N_36020);
nor U42986 (N_42986,N_36276,N_37021);
nand U42987 (N_42987,N_37569,N_38934);
xnor U42988 (N_42988,N_37843,N_36347);
nor U42989 (N_42989,N_37744,N_35881);
nand U42990 (N_42990,N_37276,N_39390);
and U42991 (N_42991,N_35729,N_39114);
xor U42992 (N_42992,N_37174,N_38753);
or U42993 (N_42993,N_38950,N_37179);
nor U42994 (N_42994,N_38084,N_36702);
nand U42995 (N_42995,N_39854,N_36455);
or U42996 (N_42996,N_35284,N_35092);
nand U42997 (N_42997,N_37412,N_37158);
xor U42998 (N_42998,N_35431,N_39816);
nand U42999 (N_42999,N_37929,N_38335);
nand U43000 (N_43000,N_38322,N_38694);
and U43001 (N_43001,N_37135,N_38112);
nor U43002 (N_43002,N_35012,N_39332);
xor U43003 (N_43003,N_38543,N_38123);
nor U43004 (N_43004,N_35835,N_35374);
nor U43005 (N_43005,N_37007,N_38019);
nand U43006 (N_43006,N_35595,N_37732);
or U43007 (N_43007,N_37903,N_36473);
and U43008 (N_43008,N_37806,N_36897);
and U43009 (N_43009,N_39451,N_36365);
or U43010 (N_43010,N_35404,N_35007);
or U43011 (N_43011,N_39836,N_38878);
nand U43012 (N_43012,N_35745,N_37394);
nand U43013 (N_43013,N_36246,N_39051);
nand U43014 (N_43014,N_39578,N_36923);
nor U43015 (N_43015,N_38309,N_35629);
or U43016 (N_43016,N_35279,N_38441);
and U43017 (N_43017,N_35275,N_35158);
and U43018 (N_43018,N_37075,N_37215);
or U43019 (N_43019,N_36538,N_36435);
nor U43020 (N_43020,N_35625,N_36699);
nor U43021 (N_43021,N_38581,N_38435);
or U43022 (N_43022,N_36947,N_38719);
xnor U43023 (N_43023,N_35395,N_37910);
nand U43024 (N_43024,N_39188,N_37937);
or U43025 (N_43025,N_36923,N_36516);
nand U43026 (N_43026,N_39055,N_35447);
xor U43027 (N_43027,N_36518,N_37857);
xnor U43028 (N_43028,N_35627,N_37156);
and U43029 (N_43029,N_38963,N_37026);
nor U43030 (N_43030,N_36514,N_36819);
nor U43031 (N_43031,N_38799,N_38009);
or U43032 (N_43032,N_35957,N_37146);
nor U43033 (N_43033,N_35770,N_39104);
xnor U43034 (N_43034,N_38432,N_35688);
nand U43035 (N_43035,N_37451,N_36978);
or U43036 (N_43036,N_39970,N_35451);
xnor U43037 (N_43037,N_39825,N_38524);
and U43038 (N_43038,N_39171,N_36320);
and U43039 (N_43039,N_36200,N_35504);
xnor U43040 (N_43040,N_35593,N_36259);
and U43041 (N_43041,N_37374,N_38023);
and U43042 (N_43042,N_38113,N_39632);
xnor U43043 (N_43043,N_38821,N_37067);
and U43044 (N_43044,N_35970,N_36462);
nor U43045 (N_43045,N_35319,N_35194);
xnor U43046 (N_43046,N_36770,N_35308);
nor U43047 (N_43047,N_35986,N_39375);
and U43048 (N_43048,N_35583,N_36337);
or U43049 (N_43049,N_35449,N_35973);
or U43050 (N_43050,N_38710,N_37724);
and U43051 (N_43051,N_38507,N_35917);
nand U43052 (N_43052,N_38830,N_38828);
or U43053 (N_43053,N_38164,N_38385);
and U43054 (N_43054,N_35226,N_39921);
nor U43055 (N_43055,N_36366,N_39920);
and U43056 (N_43056,N_36804,N_38268);
nand U43057 (N_43057,N_37715,N_39848);
and U43058 (N_43058,N_39274,N_39788);
or U43059 (N_43059,N_39814,N_37843);
nand U43060 (N_43060,N_35720,N_38131);
nor U43061 (N_43061,N_39609,N_35182);
or U43062 (N_43062,N_36884,N_38893);
nand U43063 (N_43063,N_35296,N_36123);
or U43064 (N_43064,N_37835,N_38065);
nand U43065 (N_43065,N_35630,N_37527);
nor U43066 (N_43066,N_35991,N_35646);
nor U43067 (N_43067,N_36543,N_38666);
and U43068 (N_43068,N_37942,N_37691);
nand U43069 (N_43069,N_39635,N_37146);
and U43070 (N_43070,N_36525,N_38406);
and U43071 (N_43071,N_36831,N_39738);
xnor U43072 (N_43072,N_35272,N_38102);
and U43073 (N_43073,N_36064,N_35326);
nor U43074 (N_43074,N_39776,N_37077);
nand U43075 (N_43075,N_36838,N_39929);
and U43076 (N_43076,N_39154,N_39773);
xnor U43077 (N_43077,N_37471,N_38743);
or U43078 (N_43078,N_36543,N_38484);
or U43079 (N_43079,N_35886,N_36040);
nand U43080 (N_43080,N_37836,N_36698);
nand U43081 (N_43081,N_39697,N_35819);
xor U43082 (N_43082,N_39687,N_38125);
nand U43083 (N_43083,N_39015,N_38154);
xor U43084 (N_43084,N_36160,N_39482);
nand U43085 (N_43085,N_36004,N_36457);
and U43086 (N_43086,N_36108,N_35649);
nand U43087 (N_43087,N_35278,N_35325);
and U43088 (N_43088,N_37427,N_35947);
nand U43089 (N_43089,N_37071,N_39893);
nor U43090 (N_43090,N_39751,N_36101);
and U43091 (N_43091,N_35344,N_38121);
xnor U43092 (N_43092,N_39274,N_38248);
nor U43093 (N_43093,N_35224,N_35599);
nand U43094 (N_43094,N_37659,N_38804);
nor U43095 (N_43095,N_35410,N_36524);
and U43096 (N_43096,N_35401,N_39582);
nand U43097 (N_43097,N_37720,N_39139);
or U43098 (N_43098,N_35253,N_36538);
nor U43099 (N_43099,N_39359,N_37311);
or U43100 (N_43100,N_38080,N_35554);
xnor U43101 (N_43101,N_38975,N_39043);
xor U43102 (N_43102,N_36160,N_37338);
xnor U43103 (N_43103,N_39062,N_37533);
nor U43104 (N_43104,N_39762,N_35889);
xor U43105 (N_43105,N_38552,N_35789);
nand U43106 (N_43106,N_39049,N_36489);
nor U43107 (N_43107,N_38128,N_38777);
nor U43108 (N_43108,N_36502,N_35858);
nand U43109 (N_43109,N_38381,N_39282);
nand U43110 (N_43110,N_38005,N_36307);
or U43111 (N_43111,N_38895,N_38345);
or U43112 (N_43112,N_39557,N_38832);
xor U43113 (N_43113,N_36348,N_36482);
nor U43114 (N_43114,N_39153,N_38667);
nor U43115 (N_43115,N_35081,N_36708);
xor U43116 (N_43116,N_35273,N_39742);
and U43117 (N_43117,N_36849,N_35088);
and U43118 (N_43118,N_39812,N_39395);
nor U43119 (N_43119,N_37739,N_39001);
xor U43120 (N_43120,N_38181,N_36656);
or U43121 (N_43121,N_35606,N_35079);
and U43122 (N_43122,N_39601,N_37350);
xnor U43123 (N_43123,N_36756,N_37737);
and U43124 (N_43124,N_39878,N_35053);
xnor U43125 (N_43125,N_38017,N_37811);
nand U43126 (N_43126,N_35938,N_39577);
nand U43127 (N_43127,N_37284,N_38819);
nor U43128 (N_43128,N_37482,N_36788);
nor U43129 (N_43129,N_38841,N_39931);
or U43130 (N_43130,N_36716,N_36024);
or U43131 (N_43131,N_36748,N_37698);
xnor U43132 (N_43132,N_38920,N_35164);
nand U43133 (N_43133,N_36815,N_39511);
nand U43134 (N_43134,N_37338,N_38875);
xnor U43135 (N_43135,N_37028,N_36829);
xor U43136 (N_43136,N_36182,N_39135);
nor U43137 (N_43137,N_35368,N_38756);
nand U43138 (N_43138,N_35365,N_38251);
xor U43139 (N_43139,N_38929,N_39890);
xor U43140 (N_43140,N_39771,N_37268);
nor U43141 (N_43141,N_35082,N_39194);
xor U43142 (N_43142,N_37307,N_36607);
xor U43143 (N_43143,N_37817,N_36086);
and U43144 (N_43144,N_38092,N_35907);
and U43145 (N_43145,N_37925,N_39247);
xnor U43146 (N_43146,N_36982,N_36254);
and U43147 (N_43147,N_37990,N_35193);
nor U43148 (N_43148,N_37144,N_37270);
nor U43149 (N_43149,N_36923,N_37679);
and U43150 (N_43150,N_37272,N_38702);
nand U43151 (N_43151,N_36739,N_37769);
nor U43152 (N_43152,N_38101,N_39332);
nor U43153 (N_43153,N_38166,N_36604);
nor U43154 (N_43154,N_38371,N_37598);
or U43155 (N_43155,N_39394,N_37282);
nor U43156 (N_43156,N_39102,N_36703);
or U43157 (N_43157,N_39633,N_35389);
and U43158 (N_43158,N_39631,N_38136);
and U43159 (N_43159,N_35488,N_35802);
nor U43160 (N_43160,N_37513,N_39340);
or U43161 (N_43161,N_39516,N_38751);
xnor U43162 (N_43162,N_35899,N_37309);
nand U43163 (N_43163,N_39616,N_37913);
nand U43164 (N_43164,N_38300,N_37773);
xnor U43165 (N_43165,N_36015,N_35840);
and U43166 (N_43166,N_35548,N_37819);
nand U43167 (N_43167,N_38575,N_38322);
nand U43168 (N_43168,N_38921,N_39512);
or U43169 (N_43169,N_35822,N_38087);
nand U43170 (N_43170,N_39378,N_36396);
nand U43171 (N_43171,N_37414,N_38603);
xnor U43172 (N_43172,N_39942,N_39802);
or U43173 (N_43173,N_38625,N_39965);
or U43174 (N_43174,N_39730,N_37344);
nor U43175 (N_43175,N_35515,N_37524);
or U43176 (N_43176,N_38299,N_39600);
nand U43177 (N_43177,N_38722,N_38834);
and U43178 (N_43178,N_37323,N_35294);
or U43179 (N_43179,N_39833,N_37145);
nand U43180 (N_43180,N_37071,N_39523);
nor U43181 (N_43181,N_38839,N_39575);
and U43182 (N_43182,N_38209,N_36563);
xor U43183 (N_43183,N_37961,N_36795);
and U43184 (N_43184,N_35273,N_36827);
or U43185 (N_43185,N_39379,N_39166);
xnor U43186 (N_43186,N_37886,N_39194);
xor U43187 (N_43187,N_36566,N_36439);
or U43188 (N_43188,N_37922,N_35660);
and U43189 (N_43189,N_35732,N_37264);
nand U43190 (N_43190,N_38763,N_36287);
and U43191 (N_43191,N_38290,N_36264);
nor U43192 (N_43192,N_35291,N_36443);
and U43193 (N_43193,N_35754,N_35098);
nand U43194 (N_43194,N_35953,N_35107);
nor U43195 (N_43195,N_37057,N_37272);
xor U43196 (N_43196,N_38593,N_35222);
xor U43197 (N_43197,N_38461,N_38707);
nand U43198 (N_43198,N_35588,N_38339);
nand U43199 (N_43199,N_37099,N_39212);
xor U43200 (N_43200,N_35673,N_39360);
or U43201 (N_43201,N_36181,N_37539);
xnor U43202 (N_43202,N_36991,N_37272);
and U43203 (N_43203,N_35093,N_35802);
nor U43204 (N_43204,N_36136,N_37312);
nand U43205 (N_43205,N_35709,N_38315);
nor U43206 (N_43206,N_37428,N_37381);
nand U43207 (N_43207,N_38583,N_39186);
nor U43208 (N_43208,N_37182,N_38170);
nor U43209 (N_43209,N_37548,N_39887);
nand U43210 (N_43210,N_37420,N_38755);
or U43211 (N_43211,N_37227,N_35895);
nand U43212 (N_43212,N_35476,N_38011);
and U43213 (N_43213,N_37870,N_39482);
or U43214 (N_43214,N_39790,N_35728);
nand U43215 (N_43215,N_38468,N_38334);
nor U43216 (N_43216,N_35694,N_35407);
nor U43217 (N_43217,N_37867,N_39876);
xnor U43218 (N_43218,N_37917,N_38359);
xor U43219 (N_43219,N_36546,N_37891);
and U43220 (N_43220,N_38295,N_39861);
nor U43221 (N_43221,N_36729,N_36035);
nand U43222 (N_43222,N_35364,N_35511);
nand U43223 (N_43223,N_36517,N_37553);
xnor U43224 (N_43224,N_37668,N_38887);
and U43225 (N_43225,N_37568,N_39751);
xnor U43226 (N_43226,N_37832,N_35530);
nand U43227 (N_43227,N_37071,N_37078);
xnor U43228 (N_43228,N_36681,N_36922);
or U43229 (N_43229,N_35211,N_36062);
nand U43230 (N_43230,N_35525,N_39998);
nor U43231 (N_43231,N_35503,N_38243);
or U43232 (N_43232,N_35260,N_39601);
nand U43233 (N_43233,N_35548,N_39844);
nor U43234 (N_43234,N_35629,N_38412);
nand U43235 (N_43235,N_36637,N_39658);
nand U43236 (N_43236,N_35719,N_37355);
nand U43237 (N_43237,N_35635,N_39305);
nor U43238 (N_43238,N_37003,N_39147);
xnor U43239 (N_43239,N_38426,N_36128);
nor U43240 (N_43240,N_37041,N_37923);
nand U43241 (N_43241,N_39139,N_37881);
xnor U43242 (N_43242,N_36121,N_36247);
nor U43243 (N_43243,N_39641,N_38999);
and U43244 (N_43244,N_36803,N_37346);
nor U43245 (N_43245,N_35125,N_38582);
nor U43246 (N_43246,N_36499,N_36848);
xnor U43247 (N_43247,N_38191,N_39976);
nand U43248 (N_43248,N_35586,N_35681);
or U43249 (N_43249,N_37398,N_38334);
or U43250 (N_43250,N_37151,N_37374);
xnor U43251 (N_43251,N_36528,N_39663);
xnor U43252 (N_43252,N_38716,N_38399);
nor U43253 (N_43253,N_37251,N_35624);
nor U43254 (N_43254,N_37722,N_39302);
nand U43255 (N_43255,N_35092,N_38755);
nand U43256 (N_43256,N_35198,N_38501);
and U43257 (N_43257,N_38605,N_39092);
and U43258 (N_43258,N_37329,N_37070);
nand U43259 (N_43259,N_35389,N_37795);
nand U43260 (N_43260,N_35236,N_36191);
and U43261 (N_43261,N_39706,N_38727);
and U43262 (N_43262,N_35866,N_36790);
nor U43263 (N_43263,N_37911,N_37129);
and U43264 (N_43264,N_38117,N_37632);
or U43265 (N_43265,N_35966,N_38314);
nand U43266 (N_43266,N_37612,N_38755);
or U43267 (N_43267,N_37547,N_36495);
and U43268 (N_43268,N_38644,N_39876);
and U43269 (N_43269,N_36037,N_39133);
xnor U43270 (N_43270,N_35783,N_35360);
xor U43271 (N_43271,N_39423,N_35658);
and U43272 (N_43272,N_39257,N_36342);
or U43273 (N_43273,N_39808,N_36011);
xor U43274 (N_43274,N_38664,N_38170);
nand U43275 (N_43275,N_35440,N_35370);
and U43276 (N_43276,N_37634,N_38479);
or U43277 (N_43277,N_37516,N_35496);
xnor U43278 (N_43278,N_35548,N_35775);
and U43279 (N_43279,N_38362,N_35648);
or U43280 (N_43280,N_39593,N_36002);
nor U43281 (N_43281,N_35334,N_35528);
nand U43282 (N_43282,N_35203,N_35429);
and U43283 (N_43283,N_37619,N_35928);
or U43284 (N_43284,N_38803,N_37614);
nand U43285 (N_43285,N_37086,N_38399);
or U43286 (N_43286,N_35446,N_38569);
nor U43287 (N_43287,N_39473,N_36347);
or U43288 (N_43288,N_36725,N_35756);
and U43289 (N_43289,N_39529,N_35401);
nor U43290 (N_43290,N_35886,N_36778);
nor U43291 (N_43291,N_35918,N_35993);
nor U43292 (N_43292,N_38052,N_36930);
xnor U43293 (N_43293,N_37908,N_38122);
and U43294 (N_43294,N_38451,N_39953);
xor U43295 (N_43295,N_35869,N_39398);
nor U43296 (N_43296,N_36594,N_38923);
or U43297 (N_43297,N_35862,N_35542);
nor U43298 (N_43298,N_35174,N_39028);
or U43299 (N_43299,N_37458,N_37484);
or U43300 (N_43300,N_39173,N_38601);
or U43301 (N_43301,N_38202,N_39360);
nand U43302 (N_43302,N_36520,N_39142);
xnor U43303 (N_43303,N_38295,N_39934);
and U43304 (N_43304,N_39020,N_35745);
xor U43305 (N_43305,N_39901,N_37965);
nor U43306 (N_43306,N_37589,N_39534);
nand U43307 (N_43307,N_36847,N_38428);
xor U43308 (N_43308,N_39112,N_35672);
xnor U43309 (N_43309,N_39283,N_36550);
xnor U43310 (N_43310,N_37579,N_37512);
xor U43311 (N_43311,N_39782,N_36038);
or U43312 (N_43312,N_38180,N_35801);
xor U43313 (N_43313,N_36853,N_35370);
or U43314 (N_43314,N_35094,N_36740);
xor U43315 (N_43315,N_37622,N_36321);
and U43316 (N_43316,N_36813,N_37497);
nor U43317 (N_43317,N_39720,N_36901);
nand U43318 (N_43318,N_38174,N_38481);
xor U43319 (N_43319,N_39494,N_36020);
nand U43320 (N_43320,N_35682,N_36549);
nand U43321 (N_43321,N_36393,N_39761);
nor U43322 (N_43322,N_39382,N_36152);
xnor U43323 (N_43323,N_37297,N_38945);
xor U43324 (N_43324,N_38604,N_38913);
nor U43325 (N_43325,N_37837,N_39899);
xor U43326 (N_43326,N_36534,N_39274);
xnor U43327 (N_43327,N_37528,N_35449);
xor U43328 (N_43328,N_37373,N_39825);
nand U43329 (N_43329,N_36012,N_36267);
xor U43330 (N_43330,N_37535,N_38773);
and U43331 (N_43331,N_36911,N_35658);
and U43332 (N_43332,N_38384,N_36417);
nand U43333 (N_43333,N_38435,N_36545);
or U43334 (N_43334,N_36166,N_39762);
nand U43335 (N_43335,N_37401,N_38591);
nor U43336 (N_43336,N_35396,N_37880);
nor U43337 (N_43337,N_36300,N_39366);
nand U43338 (N_43338,N_37907,N_37691);
and U43339 (N_43339,N_39062,N_36511);
or U43340 (N_43340,N_38504,N_39518);
xnor U43341 (N_43341,N_36283,N_35254);
nand U43342 (N_43342,N_36890,N_37770);
and U43343 (N_43343,N_36579,N_38901);
nand U43344 (N_43344,N_35682,N_36265);
or U43345 (N_43345,N_35760,N_37906);
nand U43346 (N_43346,N_39239,N_39000);
nor U43347 (N_43347,N_36004,N_38941);
nand U43348 (N_43348,N_35912,N_38021);
xnor U43349 (N_43349,N_36319,N_36349);
and U43350 (N_43350,N_36110,N_39585);
or U43351 (N_43351,N_37506,N_38368);
nor U43352 (N_43352,N_38728,N_39296);
or U43353 (N_43353,N_37794,N_38771);
xor U43354 (N_43354,N_35338,N_36859);
or U43355 (N_43355,N_38513,N_37605);
nand U43356 (N_43356,N_35950,N_39866);
nand U43357 (N_43357,N_35967,N_35108);
xnor U43358 (N_43358,N_39609,N_37474);
or U43359 (N_43359,N_37661,N_35596);
or U43360 (N_43360,N_36721,N_39065);
nand U43361 (N_43361,N_35051,N_39802);
or U43362 (N_43362,N_38351,N_37175);
nor U43363 (N_43363,N_38627,N_35636);
xnor U43364 (N_43364,N_37467,N_36125);
xor U43365 (N_43365,N_35284,N_37611);
and U43366 (N_43366,N_39756,N_37881);
xnor U43367 (N_43367,N_36061,N_38188);
nor U43368 (N_43368,N_39062,N_38607);
nor U43369 (N_43369,N_39937,N_39686);
and U43370 (N_43370,N_36036,N_38289);
xnor U43371 (N_43371,N_36851,N_39843);
xnor U43372 (N_43372,N_37771,N_38607);
and U43373 (N_43373,N_39982,N_35489);
or U43374 (N_43374,N_35735,N_37262);
nand U43375 (N_43375,N_38810,N_38982);
or U43376 (N_43376,N_38731,N_36385);
xnor U43377 (N_43377,N_36957,N_38414);
or U43378 (N_43378,N_38357,N_38154);
xor U43379 (N_43379,N_39027,N_35265);
nand U43380 (N_43380,N_37381,N_37698);
nor U43381 (N_43381,N_38442,N_37792);
or U43382 (N_43382,N_36632,N_38240);
xnor U43383 (N_43383,N_35175,N_38934);
nand U43384 (N_43384,N_38826,N_37452);
or U43385 (N_43385,N_37299,N_36370);
nor U43386 (N_43386,N_38553,N_39521);
and U43387 (N_43387,N_37444,N_39972);
nand U43388 (N_43388,N_36090,N_37161);
nor U43389 (N_43389,N_36395,N_35619);
nand U43390 (N_43390,N_38358,N_38521);
nor U43391 (N_43391,N_36985,N_37886);
xnor U43392 (N_43392,N_35119,N_35294);
and U43393 (N_43393,N_36796,N_38690);
nand U43394 (N_43394,N_39662,N_35030);
or U43395 (N_43395,N_35327,N_38380);
nor U43396 (N_43396,N_36176,N_37520);
nor U43397 (N_43397,N_36755,N_38395);
nor U43398 (N_43398,N_38980,N_37133);
nor U43399 (N_43399,N_35703,N_36904);
or U43400 (N_43400,N_35360,N_36981);
nand U43401 (N_43401,N_36422,N_39196);
or U43402 (N_43402,N_39345,N_35524);
and U43403 (N_43403,N_35379,N_35348);
nor U43404 (N_43404,N_38443,N_37258);
nor U43405 (N_43405,N_38597,N_35680);
or U43406 (N_43406,N_38037,N_37842);
or U43407 (N_43407,N_35926,N_36162);
or U43408 (N_43408,N_39677,N_38484);
and U43409 (N_43409,N_37257,N_38505);
nor U43410 (N_43410,N_36972,N_36364);
nor U43411 (N_43411,N_38658,N_36630);
nand U43412 (N_43412,N_38020,N_39147);
nand U43413 (N_43413,N_36946,N_36938);
nand U43414 (N_43414,N_36987,N_36546);
xor U43415 (N_43415,N_39842,N_36681);
nand U43416 (N_43416,N_37162,N_38103);
and U43417 (N_43417,N_35771,N_36931);
and U43418 (N_43418,N_37038,N_38185);
xnor U43419 (N_43419,N_35042,N_37213);
and U43420 (N_43420,N_35708,N_39026);
nor U43421 (N_43421,N_36169,N_39036);
xor U43422 (N_43422,N_38965,N_38632);
or U43423 (N_43423,N_39781,N_35871);
nand U43424 (N_43424,N_37514,N_35579);
nand U43425 (N_43425,N_38682,N_35628);
nand U43426 (N_43426,N_37142,N_38413);
nor U43427 (N_43427,N_35709,N_37595);
or U43428 (N_43428,N_39491,N_35701);
nor U43429 (N_43429,N_39047,N_39520);
nor U43430 (N_43430,N_35757,N_37619);
nor U43431 (N_43431,N_35618,N_36497);
xor U43432 (N_43432,N_36740,N_35955);
nand U43433 (N_43433,N_38085,N_36587);
and U43434 (N_43434,N_39846,N_39178);
nor U43435 (N_43435,N_35779,N_35599);
xnor U43436 (N_43436,N_39710,N_36395);
nand U43437 (N_43437,N_37551,N_35897);
nor U43438 (N_43438,N_35138,N_39905);
nor U43439 (N_43439,N_38011,N_35037);
and U43440 (N_43440,N_35125,N_38885);
or U43441 (N_43441,N_39831,N_36165);
and U43442 (N_43442,N_38946,N_38268);
nand U43443 (N_43443,N_38584,N_36287);
nand U43444 (N_43444,N_36617,N_35918);
xnor U43445 (N_43445,N_36391,N_39540);
nor U43446 (N_43446,N_37488,N_39008);
nor U43447 (N_43447,N_36070,N_38238);
nor U43448 (N_43448,N_38129,N_37834);
and U43449 (N_43449,N_39446,N_38966);
nor U43450 (N_43450,N_35666,N_38205);
xor U43451 (N_43451,N_35641,N_38178);
or U43452 (N_43452,N_35387,N_35345);
or U43453 (N_43453,N_39530,N_39415);
nor U43454 (N_43454,N_37356,N_35784);
xor U43455 (N_43455,N_36990,N_38024);
nand U43456 (N_43456,N_35116,N_38950);
nor U43457 (N_43457,N_38058,N_36378);
xor U43458 (N_43458,N_35401,N_38997);
xnor U43459 (N_43459,N_35780,N_39606);
xor U43460 (N_43460,N_37595,N_37991);
xor U43461 (N_43461,N_37487,N_38158);
or U43462 (N_43462,N_37621,N_38071);
xor U43463 (N_43463,N_35035,N_38571);
or U43464 (N_43464,N_38823,N_39975);
or U43465 (N_43465,N_39243,N_37679);
and U43466 (N_43466,N_39471,N_36185);
or U43467 (N_43467,N_36497,N_39912);
nand U43468 (N_43468,N_39746,N_39072);
nor U43469 (N_43469,N_35548,N_37700);
nand U43470 (N_43470,N_37058,N_35311);
or U43471 (N_43471,N_39981,N_36288);
xor U43472 (N_43472,N_35970,N_37822);
xnor U43473 (N_43473,N_37863,N_38639);
and U43474 (N_43474,N_38623,N_37361);
or U43475 (N_43475,N_39763,N_38357);
nand U43476 (N_43476,N_38289,N_35097);
nor U43477 (N_43477,N_35305,N_35204);
nor U43478 (N_43478,N_36933,N_37058);
and U43479 (N_43479,N_39667,N_39586);
nand U43480 (N_43480,N_35389,N_39512);
nor U43481 (N_43481,N_36591,N_38050);
and U43482 (N_43482,N_36366,N_35819);
nor U43483 (N_43483,N_36344,N_38577);
or U43484 (N_43484,N_36524,N_39664);
xnor U43485 (N_43485,N_35854,N_37457);
or U43486 (N_43486,N_36566,N_39070);
nor U43487 (N_43487,N_35719,N_37680);
nand U43488 (N_43488,N_35908,N_38010);
and U43489 (N_43489,N_38702,N_35598);
xnor U43490 (N_43490,N_37279,N_37115);
and U43491 (N_43491,N_36941,N_35051);
nor U43492 (N_43492,N_37507,N_37262);
or U43493 (N_43493,N_38987,N_37185);
nand U43494 (N_43494,N_35205,N_36183);
or U43495 (N_43495,N_36202,N_36178);
nor U43496 (N_43496,N_38445,N_35252);
xor U43497 (N_43497,N_35031,N_38695);
or U43498 (N_43498,N_36938,N_35353);
nand U43499 (N_43499,N_37173,N_39480);
nor U43500 (N_43500,N_38727,N_37396);
and U43501 (N_43501,N_38514,N_36885);
nor U43502 (N_43502,N_35813,N_38776);
or U43503 (N_43503,N_36134,N_39853);
nor U43504 (N_43504,N_37318,N_38569);
xnor U43505 (N_43505,N_35015,N_38704);
and U43506 (N_43506,N_38125,N_35247);
and U43507 (N_43507,N_37784,N_36717);
and U43508 (N_43508,N_35567,N_37196);
xnor U43509 (N_43509,N_39125,N_39948);
and U43510 (N_43510,N_35816,N_39721);
and U43511 (N_43511,N_36669,N_35012);
or U43512 (N_43512,N_37109,N_37362);
xnor U43513 (N_43513,N_38581,N_36887);
nor U43514 (N_43514,N_36260,N_37878);
nor U43515 (N_43515,N_35936,N_35771);
or U43516 (N_43516,N_37449,N_36886);
nor U43517 (N_43517,N_37219,N_38636);
nor U43518 (N_43518,N_39588,N_38168);
nand U43519 (N_43519,N_37003,N_38100);
nand U43520 (N_43520,N_36230,N_37855);
nand U43521 (N_43521,N_36885,N_39390);
or U43522 (N_43522,N_38954,N_36079);
and U43523 (N_43523,N_36862,N_35264);
nor U43524 (N_43524,N_35724,N_39271);
or U43525 (N_43525,N_36965,N_39197);
or U43526 (N_43526,N_37033,N_37204);
or U43527 (N_43527,N_36692,N_38671);
xnor U43528 (N_43528,N_35515,N_36580);
nor U43529 (N_43529,N_38354,N_38798);
nand U43530 (N_43530,N_37802,N_39562);
nand U43531 (N_43531,N_38065,N_35375);
xnor U43532 (N_43532,N_38774,N_36025);
nor U43533 (N_43533,N_36365,N_37214);
nor U43534 (N_43534,N_36407,N_37319);
or U43535 (N_43535,N_35136,N_38006);
xor U43536 (N_43536,N_39899,N_39768);
or U43537 (N_43537,N_38109,N_35247);
or U43538 (N_43538,N_39593,N_39357);
nor U43539 (N_43539,N_39724,N_37424);
and U43540 (N_43540,N_36799,N_38985);
or U43541 (N_43541,N_36230,N_35682);
or U43542 (N_43542,N_37221,N_37866);
nor U43543 (N_43543,N_36126,N_38285);
nor U43544 (N_43544,N_38788,N_35615);
xnor U43545 (N_43545,N_36271,N_35180);
nand U43546 (N_43546,N_36785,N_38889);
or U43547 (N_43547,N_35901,N_37403);
and U43548 (N_43548,N_36525,N_39048);
xor U43549 (N_43549,N_35030,N_39982);
xor U43550 (N_43550,N_38413,N_37734);
nor U43551 (N_43551,N_35310,N_36299);
or U43552 (N_43552,N_38708,N_39524);
xor U43553 (N_43553,N_37489,N_39233);
or U43554 (N_43554,N_39167,N_35937);
nor U43555 (N_43555,N_35561,N_36314);
nor U43556 (N_43556,N_36791,N_38257);
xnor U43557 (N_43557,N_37389,N_35387);
xnor U43558 (N_43558,N_37998,N_37858);
nor U43559 (N_43559,N_38376,N_36312);
xor U43560 (N_43560,N_35726,N_38964);
xor U43561 (N_43561,N_35294,N_38477);
nand U43562 (N_43562,N_35259,N_36335);
nand U43563 (N_43563,N_36947,N_38289);
nand U43564 (N_43564,N_39063,N_37467);
nand U43565 (N_43565,N_38022,N_35510);
nand U43566 (N_43566,N_37276,N_39777);
or U43567 (N_43567,N_39226,N_38446);
or U43568 (N_43568,N_39276,N_35980);
and U43569 (N_43569,N_36953,N_35947);
xnor U43570 (N_43570,N_36538,N_35040);
xnor U43571 (N_43571,N_36814,N_38629);
or U43572 (N_43572,N_39916,N_39884);
and U43573 (N_43573,N_35613,N_38694);
or U43574 (N_43574,N_36426,N_36110);
and U43575 (N_43575,N_37699,N_39233);
xnor U43576 (N_43576,N_36935,N_35430);
and U43577 (N_43577,N_36998,N_37233);
and U43578 (N_43578,N_37387,N_38907);
nand U43579 (N_43579,N_38048,N_35972);
xnor U43580 (N_43580,N_38439,N_38994);
xor U43581 (N_43581,N_37875,N_36441);
nand U43582 (N_43582,N_38462,N_36482);
nand U43583 (N_43583,N_39352,N_36675);
xnor U43584 (N_43584,N_39223,N_38237);
or U43585 (N_43585,N_36905,N_39588);
and U43586 (N_43586,N_37737,N_36780);
nand U43587 (N_43587,N_37822,N_37909);
xor U43588 (N_43588,N_39485,N_35367);
nor U43589 (N_43589,N_37981,N_37228);
nor U43590 (N_43590,N_38433,N_36940);
or U43591 (N_43591,N_39833,N_35159);
and U43592 (N_43592,N_39992,N_36447);
nand U43593 (N_43593,N_37111,N_36708);
nor U43594 (N_43594,N_38794,N_38345);
and U43595 (N_43595,N_37160,N_38740);
xor U43596 (N_43596,N_37587,N_37438);
xor U43597 (N_43597,N_37090,N_37837);
xnor U43598 (N_43598,N_39366,N_39673);
or U43599 (N_43599,N_35248,N_36251);
or U43600 (N_43600,N_38141,N_37389);
nand U43601 (N_43601,N_36831,N_37850);
and U43602 (N_43602,N_35221,N_37547);
nor U43603 (N_43603,N_35914,N_36042);
or U43604 (N_43604,N_35334,N_36004);
xnor U43605 (N_43605,N_37236,N_35953);
or U43606 (N_43606,N_36234,N_39056);
nor U43607 (N_43607,N_36661,N_39229);
or U43608 (N_43608,N_39847,N_37297);
nor U43609 (N_43609,N_37165,N_38947);
and U43610 (N_43610,N_36064,N_36023);
or U43611 (N_43611,N_35431,N_39933);
nand U43612 (N_43612,N_37852,N_38286);
nand U43613 (N_43613,N_39947,N_35477);
and U43614 (N_43614,N_39466,N_39490);
nand U43615 (N_43615,N_39847,N_38526);
nand U43616 (N_43616,N_37326,N_36528);
xor U43617 (N_43617,N_36882,N_37055);
and U43618 (N_43618,N_37246,N_36422);
nand U43619 (N_43619,N_37995,N_37795);
nor U43620 (N_43620,N_39448,N_37981);
nand U43621 (N_43621,N_38715,N_36061);
xnor U43622 (N_43622,N_36448,N_37234);
xnor U43623 (N_43623,N_35030,N_39144);
and U43624 (N_43624,N_36423,N_35740);
xor U43625 (N_43625,N_35934,N_37111);
nand U43626 (N_43626,N_39047,N_36242);
nor U43627 (N_43627,N_38919,N_36946);
xnor U43628 (N_43628,N_39071,N_38231);
nand U43629 (N_43629,N_36454,N_38132);
nor U43630 (N_43630,N_35230,N_37301);
and U43631 (N_43631,N_36779,N_35163);
xnor U43632 (N_43632,N_37990,N_35365);
and U43633 (N_43633,N_36770,N_36168);
xnor U43634 (N_43634,N_35810,N_37075);
nor U43635 (N_43635,N_36190,N_35033);
and U43636 (N_43636,N_37790,N_37680);
xnor U43637 (N_43637,N_35708,N_37724);
nand U43638 (N_43638,N_37200,N_37327);
xor U43639 (N_43639,N_36710,N_36955);
or U43640 (N_43640,N_38339,N_39837);
xor U43641 (N_43641,N_39024,N_37651);
or U43642 (N_43642,N_37045,N_39976);
and U43643 (N_43643,N_35712,N_37626);
and U43644 (N_43644,N_36246,N_35852);
nor U43645 (N_43645,N_37553,N_35780);
or U43646 (N_43646,N_36324,N_38679);
nand U43647 (N_43647,N_38721,N_38110);
or U43648 (N_43648,N_37027,N_39307);
or U43649 (N_43649,N_39846,N_35696);
xor U43650 (N_43650,N_36668,N_36296);
xor U43651 (N_43651,N_39786,N_39713);
nor U43652 (N_43652,N_36974,N_36987);
or U43653 (N_43653,N_36097,N_39580);
nor U43654 (N_43654,N_36186,N_36951);
nand U43655 (N_43655,N_39905,N_35725);
and U43656 (N_43656,N_38354,N_39210);
or U43657 (N_43657,N_38732,N_39142);
nand U43658 (N_43658,N_36063,N_38352);
xnor U43659 (N_43659,N_35025,N_39512);
xor U43660 (N_43660,N_36456,N_35985);
nor U43661 (N_43661,N_37125,N_37368);
nand U43662 (N_43662,N_36939,N_36379);
xnor U43663 (N_43663,N_35922,N_37811);
or U43664 (N_43664,N_37523,N_37371);
and U43665 (N_43665,N_37900,N_36595);
and U43666 (N_43666,N_36306,N_36469);
nor U43667 (N_43667,N_36214,N_39368);
nor U43668 (N_43668,N_39876,N_38550);
or U43669 (N_43669,N_37772,N_35953);
nor U43670 (N_43670,N_38955,N_36628);
nor U43671 (N_43671,N_35014,N_37688);
xor U43672 (N_43672,N_37913,N_37875);
nor U43673 (N_43673,N_38518,N_36414);
and U43674 (N_43674,N_35348,N_36440);
nor U43675 (N_43675,N_37885,N_37932);
nand U43676 (N_43676,N_38265,N_39849);
nor U43677 (N_43677,N_37681,N_38958);
and U43678 (N_43678,N_37131,N_36912);
or U43679 (N_43679,N_38154,N_39512);
or U43680 (N_43680,N_36053,N_36861);
and U43681 (N_43681,N_39579,N_36351);
nor U43682 (N_43682,N_38764,N_36577);
nor U43683 (N_43683,N_37299,N_36811);
nand U43684 (N_43684,N_35886,N_38531);
and U43685 (N_43685,N_35578,N_37156);
or U43686 (N_43686,N_39616,N_37643);
xnor U43687 (N_43687,N_38785,N_38169);
or U43688 (N_43688,N_35024,N_39373);
and U43689 (N_43689,N_37132,N_38513);
and U43690 (N_43690,N_36414,N_38680);
xor U43691 (N_43691,N_36158,N_35433);
xnor U43692 (N_43692,N_36983,N_39731);
xor U43693 (N_43693,N_35644,N_35045);
and U43694 (N_43694,N_36877,N_37518);
nor U43695 (N_43695,N_37432,N_37719);
nor U43696 (N_43696,N_37684,N_35186);
or U43697 (N_43697,N_38385,N_37885);
and U43698 (N_43698,N_36666,N_35702);
nand U43699 (N_43699,N_35694,N_38436);
and U43700 (N_43700,N_36978,N_37726);
xor U43701 (N_43701,N_35970,N_38667);
or U43702 (N_43702,N_37464,N_38489);
nor U43703 (N_43703,N_39988,N_37146);
or U43704 (N_43704,N_36693,N_36698);
nand U43705 (N_43705,N_35029,N_36699);
or U43706 (N_43706,N_38343,N_35561);
nor U43707 (N_43707,N_35030,N_35300);
nand U43708 (N_43708,N_39870,N_37910);
xnor U43709 (N_43709,N_38709,N_39899);
or U43710 (N_43710,N_38544,N_36137);
nand U43711 (N_43711,N_37652,N_38469);
and U43712 (N_43712,N_38845,N_38886);
nand U43713 (N_43713,N_39956,N_37063);
or U43714 (N_43714,N_39187,N_39856);
xnor U43715 (N_43715,N_36332,N_37225);
nand U43716 (N_43716,N_37320,N_35720);
xnor U43717 (N_43717,N_37114,N_37514);
and U43718 (N_43718,N_35703,N_35540);
or U43719 (N_43719,N_35911,N_35328);
or U43720 (N_43720,N_37466,N_37831);
or U43721 (N_43721,N_37462,N_36526);
nand U43722 (N_43722,N_35114,N_39927);
xnor U43723 (N_43723,N_35637,N_37191);
xor U43724 (N_43724,N_35007,N_35197);
nand U43725 (N_43725,N_39728,N_38864);
nor U43726 (N_43726,N_35785,N_39134);
or U43727 (N_43727,N_35965,N_37146);
or U43728 (N_43728,N_36624,N_35587);
and U43729 (N_43729,N_35407,N_39767);
nand U43730 (N_43730,N_38254,N_38648);
xor U43731 (N_43731,N_36025,N_36838);
xor U43732 (N_43732,N_35175,N_38348);
nand U43733 (N_43733,N_36675,N_38760);
xor U43734 (N_43734,N_37401,N_36907);
nor U43735 (N_43735,N_36816,N_36717);
nand U43736 (N_43736,N_37932,N_38245);
and U43737 (N_43737,N_36952,N_36358);
xnor U43738 (N_43738,N_38430,N_36572);
and U43739 (N_43739,N_36689,N_37458);
nand U43740 (N_43740,N_36670,N_35865);
nand U43741 (N_43741,N_38423,N_39548);
and U43742 (N_43742,N_38551,N_37807);
nor U43743 (N_43743,N_36741,N_37187);
and U43744 (N_43744,N_38349,N_36832);
nand U43745 (N_43745,N_37563,N_38978);
nand U43746 (N_43746,N_36453,N_35686);
nor U43747 (N_43747,N_37864,N_38260);
nor U43748 (N_43748,N_36053,N_39192);
or U43749 (N_43749,N_36890,N_35439);
and U43750 (N_43750,N_35370,N_39980);
xor U43751 (N_43751,N_38062,N_37458);
xnor U43752 (N_43752,N_35713,N_38236);
or U43753 (N_43753,N_36606,N_37876);
xor U43754 (N_43754,N_38651,N_36273);
xor U43755 (N_43755,N_36951,N_39679);
nand U43756 (N_43756,N_37562,N_39610);
or U43757 (N_43757,N_36902,N_36632);
or U43758 (N_43758,N_39893,N_36464);
nand U43759 (N_43759,N_37224,N_38377);
nand U43760 (N_43760,N_36118,N_37537);
xnor U43761 (N_43761,N_39947,N_36327);
or U43762 (N_43762,N_37275,N_38855);
nor U43763 (N_43763,N_36935,N_35184);
xor U43764 (N_43764,N_39967,N_38946);
and U43765 (N_43765,N_39344,N_35600);
xor U43766 (N_43766,N_35537,N_36436);
and U43767 (N_43767,N_35518,N_36690);
nor U43768 (N_43768,N_39552,N_39326);
nor U43769 (N_43769,N_39104,N_39389);
nand U43770 (N_43770,N_37953,N_36236);
nand U43771 (N_43771,N_38009,N_36068);
xnor U43772 (N_43772,N_37635,N_37481);
or U43773 (N_43773,N_37683,N_39874);
xnor U43774 (N_43774,N_39765,N_36537);
nor U43775 (N_43775,N_35480,N_37889);
and U43776 (N_43776,N_36150,N_35806);
nand U43777 (N_43777,N_36173,N_37760);
nor U43778 (N_43778,N_35311,N_39512);
or U43779 (N_43779,N_36953,N_36908);
nand U43780 (N_43780,N_37582,N_38166);
xnor U43781 (N_43781,N_35247,N_35475);
nor U43782 (N_43782,N_35238,N_38934);
xor U43783 (N_43783,N_39960,N_35541);
nor U43784 (N_43784,N_35105,N_38182);
xnor U43785 (N_43785,N_39758,N_36621);
or U43786 (N_43786,N_35454,N_38214);
nor U43787 (N_43787,N_37403,N_36269);
xnor U43788 (N_43788,N_36066,N_37906);
nor U43789 (N_43789,N_39817,N_38142);
nor U43790 (N_43790,N_36292,N_38753);
and U43791 (N_43791,N_39202,N_39960);
or U43792 (N_43792,N_36785,N_36525);
nor U43793 (N_43793,N_37770,N_38235);
nor U43794 (N_43794,N_38318,N_35017);
nor U43795 (N_43795,N_38530,N_37505);
nand U43796 (N_43796,N_38382,N_35260);
or U43797 (N_43797,N_39982,N_36081);
or U43798 (N_43798,N_38693,N_36409);
xor U43799 (N_43799,N_35203,N_38106);
nor U43800 (N_43800,N_35377,N_39756);
and U43801 (N_43801,N_38053,N_39377);
xnor U43802 (N_43802,N_38915,N_39460);
xnor U43803 (N_43803,N_38780,N_35232);
xor U43804 (N_43804,N_39788,N_35472);
or U43805 (N_43805,N_39000,N_36058);
nand U43806 (N_43806,N_39896,N_36897);
nor U43807 (N_43807,N_38620,N_37344);
xnor U43808 (N_43808,N_36569,N_35990);
nand U43809 (N_43809,N_38718,N_39033);
or U43810 (N_43810,N_39763,N_38475);
or U43811 (N_43811,N_37888,N_36431);
and U43812 (N_43812,N_36925,N_38806);
or U43813 (N_43813,N_39143,N_37037);
xor U43814 (N_43814,N_38419,N_37818);
and U43815 (N_43815,N_36383,N_38619);
nor U43816 (N_43816,N_37787,N_36973);
nand U43817 (N_43817,N_39600,N_35058);
nand U43818 (N_43818,N_36718,N_38242);
xnor U43819 (N_43819,N_37888,N_36525);
and U43820 (N_43820,N_35178,N_38575);
xor U43821 (N_43821,N_37457,N_38240);
nand U43822 (N_43822,N_38846,N_35800);
nor U43823 (N_43823,N_36920,N_35519);
and U43824 (N_43824,N_37349,N_39662);
or U43825 (N_43825,N_37465,N_39315);
and U43826 (N_43826,N_39970,N_36571);
nand U43827 (N_43827,N_38764,N_38403);
xor U43828 (N_43828,N_39217,N_37097);
nand U43829 (N_43829,N_39597,N_39010);
nand U43830 (N_43830,N_35365,N_35540);
xnor U43831 (N_43831,N_39043,N_36402);
xnor U43832 (N_43832,N_38073,N_36505);
xnor U43833 (N_43833,N_35132,N_38605);
nor U43834 (N_43834,N_35693,N_38007);
nor U43835 (N_43835,N_38340,N_38423);
or U43836 (N_43836,N_39216,N_38824);
nor U43837 (N_43837,N_36027,N_35301);
nand U43838 (N_43838,N_38252,N_36208);
and U43839 (N_43839,N_38815,N_35001);
nor U43840 (N_43840,N_35788,N_38261);
xnor U43841 (N_43841,N_37924,N_36651);
or U43842 (N_43842,N_36087,N_37529);
or U43843 (N_43843,N_39304,N_35877);
and U43844 (N_43844,N_38688,N_39572);
nor U43845 (N_43845,N_38044,N_38647);
xor U43846 (N_43846,N_36899,N_36135);
and U43847 (N_43847,N_37979,N_38988);
nor U43848 (N_43848,N_35886,N_36143);
and U43849 (N_43849,N_37791,N_39940);
nand U43850 (N_43850,N_39622,N_35939);
nand U43851 (N_43851,N_38158,N_35271);
nor U43852 (N_43852,N_37842,N_38733);
nor U43853 (N_43853,N_37120,N_38191);
xnor U43854 (N_43854,N_35549,N_36566);
xor U43855 (N_43855,N_39392,N_39032);
or U43856 (N_43856,N_35280,N_39284);
nand U43857 (N_43857,N_37982,N_39724);
nand U43858 (N_43858,N_36364,N_35441);
and U43859 (N_43859,N_36239,N_35810);
and U43860 (N_43860,N_35072,N_35110);
and U43861 (N_43861,N_36301,N_38447);
nor U43862 (N_43862,N_35455,N_39616);
and U43863 (N_43863,N_36708,N_35827);
and U43864 (N_43864,N_35384,N_38848);
nand U43865 (N_43865,N_35691,N_37296);
xnor U43866 (N_43866,N_39635,N_38777);
xnor U43867 (N_43867,N_38168,N_38460);
xnor U43868 (N_43868,N_36739,N_35485);
and U43869 (N_43869,N_38763,N_36828);
or U43870 (N_43870,N_35212,N_39708);
or U43871 (N_43871,N_36360,N_38223);
nor U43872 (N_43872,N_38073,N_37783);
xnor U43873 (N_43873,N_36357,N_35567);
nand U43874 (N_43874,N_37285,N_36570);
and U43875 (N_43875,N_39433,N_36176);
or U43876 (N_43876,N_35199,N_35904);
or U43877 (N_43877,N_35099,N_36300);
nand U43878 (N_43878,N_39035,N_38571);
xor U43879 (N_43879,N_35929,N_35160);
nor U43880 (N_43880,N_35708,N_35199);
and U43881 (N_43881,N_38121,N_36341);
xnor U43882 (N_43882,N_39207,N_36260);
nand U43883 (N_43883,N_39732,N_39310);
nor U43884 (N_43884,N_38744,N_37000);
nor U43885 (N_43885,N_35832,N_39220);
xor U43886 (N_43886,N_38744,N_35865);
nor U43887 (N_43887,N_35894,N_36045);
or U43888 (N_43888,N_35367,N_38922);
and U43889 (N_43889,N_35574,N_35665);
xor U43890 (N_43890,N_38729,N_36124);
or U43891 (N_43891,N_35129,N_39318);
nor U43892 (N_43892,N_39454,N_39418);
or U43893 (N_43893,N_36562,N_38536);
xor U43894 (N_43894,N_36045,N_39810);
nand U43895 (N_43895,N_38008,N_39703);
and U43896 (N_43896,N_39627,N_36372);
and U43897 (N_43897,N_35671,N_37102);
nor U43898 (N_43898,N_38650,N_37461);
nand U43899 (N_43899,N_37243,N_36323);
or U43900 (N_43900,N_38718,N_37279);
nor U43901 (N_43901,N_39744,N_36263);
nor U43902 (N_43902,N_39621,N_37643);
nor U43903 (N_43903,N_36358,N_36909);
or U43904 (N_43904,N_37091,N_36497);
and U43905 (N_43905,N_35227,N_39411);
nor U43906 (N_43906,N_37518,N_36027);
nand U43907 (N_43907,N_37712,N_38532);
xor U43908 (N_43908,N_38761,N_38474);
or U43909 (N_43909,N_39210,N_39895);
or U43910 (N_43910,N_36934,N_38006);
nand U43911 (N_43911,N_38403,N_38620);
nand U43912 (N_43912,N_36517,N_36398);
xor U43913 (N_43913,N_36540,N_38560);
xor U43914 (N_43914,N_37699,N_35303);
nor U43915 (N_43915,N_38022,N_37341);
xor U43916 (N_43916,N_35321,N_37002);
nor U43917 (N_43917,N_39170,N_38128);
nor U43918 (N_43918,N_38902,N_35670);
nand U43919 (N_43919,N_35057,N_38642);
or U43920 (N_43920,N_35332,N_39413);
or U43921 (N_43921,N_38363,N_39240);
nor U43922 (N_43922,N_36226,N_38943);
nand U43923 (N_43923,N_39808,N_38328);
and U43924 (N_43924,N_39962,N_38746);
nor U43925 (N_43925,N_39310,N_36640);
xor U43926 (N_43926,N_37984,N_36048);
xnor U43927 (N_43927,N_39273,N_36655);
nand U43928 (N_43928,N_39551,N_36046);
or U43929 (N_43929,N_36440,N_39170);
nor U43930 (N_43930,N_37576,N_39807);
and U43931 (N_43931,N_39841,N_38790);
and U43932 (N_43932,N_35886,N_36054);
xor U43933 (N_43933,N_38417,N_39238);
nand U43934 (N_43934,N_38206,N_36400);
nand U43935 (N_43935,N_37904,N_36713);
or U43936 (N_43936,N_35416,N_35123);
nand U43937 (N_43937,N_38559,N_37920);
or U43938 (N_43938,N_39563,N_36723);
xnor U43939 (N_43939,N_38918,N_36269);
nor U43940 (N_43940,N_35234,N_35068);
or U43941 (N_43941,N_39504,N_35814);
xnor U43942 (N_43942,N_35012,N_35982);
nor U43943 (N_43943,N_36779,N_38644);
or U43944 (N_43944,N_37095,N_35786);
nand U43945 (N_43945,N_38614,N_38102);
xnor U43946 (N_43946,N_39650,N_37376);
xnor U43947 (N_43947,N_37985,N_36693);
and U43948 (N_43948,N_37486,N_36579);
nand U43949 (N_43949,N_37150,N_37106);
and U43950 (N_43950,N_39224,N_38351);
nand U43951 (N_43951,N_37467,N_39288);
nand U43952 (N_43952,N_38520,N_36584);
xor U43953 (N_43953,N_39763,N_35786);
and U43954 (N_43954,N_35163,N_38841);
xor U43955 (N_43955,N_36187,N_35633);
or U43956 (N_43956,N_38358,N_39442);
or U43957 (N_43957,N_38840,N_38639);
or U43958 (N_43958,N_39567,N_36800);
nand U43959 (N_43959,N_38622,N_36009);
and U43960 (N_43960,N_39111,N_39920);
xor U43961 (N_43961,N_36019,N_39518);
xnor U43962 (N_43962,N_39863,N_37517);
xor U43963 (N_43963,N_36367,N_39428);
nor U43964 (N_43964,N_35877,N_37764);
and U43965 (N_43965,N_38186,N_36860);
nand U43966 (N_43966,N_39294,N_36984);
and U43967 (N_43967,N_37762,N_38874);
or U43968 (N_43968,N_39447,N_38533);
and U43969 (N_43969,N_39432,N_39278);
nor U43970 (N_43970,N_37843,N_37602);
or U43971 (N_43971,N_36534,N_37325);
nor U43972 (N_43972,N_37687,N_36107);
or U43973 (N_43973,N_37553,N_37029);
or U43974 (N_43974,N_39678,N_37376);
or U43975 (N_43975,N_37482,N_38115);
xor U43976 (N_43976,N_35839,N_39847);
nand U43977 (N_43977,N_35464,N_36871);
xnor U43978 (N_43978,N_38352,N_35621);
xnor U43979 (N_43979,N_35099,N_36688);
nor U43980 (N_43980,N_38359,N_38312);
xor U43981 (N_43981,N_37804,N_35232);
xor U43982 (N_43982,N_36833,N_36951);
and U43983 (N_43983,N_38759,N_37746);
nor U43984 (N_43984,N_38516,N_37033);
or U43985 (N_43985,N_38233,N_37483);
and U43986 (N_43986,N_36024,N_39461);
nand U43987 (N_43987,N_37136,N_39660);
and U43988 (N_43988,N_38680,N_37570);
and U43989 (N_43989,N_35066,N_35349);
xor U43990 (N_43990,N_35916,N_37029);
nand U43991 (N_43991,N_37764,N_36124);
and U43992 (N_43992,N_39957,N_35006);
or U43993 (N_43993,N_35827,N_36410);
nor U43994 (N_43994,N_36111,N_36157);
nand U43995 (N_43995,N_39348,N_35159);
and U43996 (N_43996,N_35997,N_36923);
nand U43997 (N_43997,N_39117,N_38702);
and U43998 (N_43998,N_37482,N_35298);
xnor U43999 (N_43999,N_39338,N_35826);
or U44000 (N_44000,N_35157,N_39697);
xnor U44001 (N_44001,N_35625,N_38474);
and U44002 (N_44002,N_36710,N_38884);
xnor U44003 (N_44003,N_36603,N_38271);
and U44004 (N_44004,N_37792,N_37993);
xor U44005 (N_44005,N_37888,N_38627);
or U44006 (N_44006,N_39612,N_37861);
xnor U44007 (N_44007,N_38959,N_38544);
xor U44008 (N_44008,N_36356,N_38811);
nand U44009 (N_44009,N_37533,N_35660);
nor U44010 (N_44010,N_37263,N_38490);
nand U44011 (N_44011,N_36685,N_39107);
nor U44012 (N_44012,N_38300,N_35214);
or U44013 (N_44013,N_37668,N_37227);
or U44014 (N_44014,N_35516,N_36045);
nor U44015 (N_44015,N_39445,N_37865);
xor U44016 (N_44016,N_37139,N_37193);
or U44017 (N_44017,N_36358,N_37849);
nor U44018 (N_44018,N_39543,N_38673);
xnor U44019 (N_44019,N_37217,N_36033);
and U44020 (N_44020,N_37821,N_37448);
nor U44021 (N_44021,N_39618,N_37434);
nand U44022 (N_44022,N_36096,N_38658);
and U44023 (N_44023,N_37820,N_39232);
and U44024 (N_44024,N_35598,N_39155);
nand U44025 (N_44025,N_35822,N_37205);
and U44026 (N_44026,N_37342,N_35025);
nand U44027 (N_44027,N_35877,N_39944);
nor U44028 (N_44028,N_36913,N_38997);
nand U44029 (N_44029,N_38638,N_36117);
and U44030 (N_44030,N_35037,N_37909);
or U44031 (N_44031,N_37233,N_35949);
xor U44032 (N_44032,N_35427,N_37005);
and U44033 (N_44033,N_38224,N_37362);
or U44034 (N_44034,N_39849,N_36750);
or U44035 (N_44035,N_35813,N_35176);
and U44036 (N_44036,N_37088,N_35848);
and U44037 (N_44037,N_38797,N_38949);
nand U44038 (N_44038,N_37087,N_35066);
and U44039 (N_44039,N_37935,N_37146);
and U44040 (N_44040,N_36520,N_38940);
or U44041 (N_44041,N_35092,N_36719);
xor U44042 (N_44042,N_38537,N_37625);
nor U44043 (N_44043,N_36483,N_37099);
nand U44044 (N_44044,N_39651,N_38891);
nor U44045 (N_44045,N_38886,N_38226);
nor U44046 (N_44046,N_36194,N_39956);
and U44047 (N_44047,N_39777,N_36404);
xnor U44048 (N_44048,N_39077,N_37082);
nor U44049 (N_44049,N_38506,N_38619);
or U44050 (N_44050,N_37862,N_39909);
nor U44051 (N_44051,N_38942,N_39633);
and U44052 (N_44052,N_35432,N_36345);
xnor U44053 (N_44053,N_38105,N_37241);
and U44054 (N_44054,N_36475,N_38312);
or U44055 (N_44055,N_35908,N_38668);
and U44056 (N_44056,N_35472,N_39278);
and U44057 (N_44057,N_36453,N_39869);
and U44058 (N_44058,N_37204,N_38981);
xnor U44059 (N_44059,N_39100,N_39863);
nand U44060 (N_44060,N_38120,N_38770);
or U44061 (N_44061,N_39457,N_37000);
and U44062 (N_44062,N_39489,N_36592);
nand U44063 (N_44063,N_37101,N_35983);
and U44064 (N_44064,N_36854,N_37923);
or U44065 (N_44065,N_35702,N_35377);
or U44066 (N_44066,N_36891,N_37109);
nand U44067 (N_44067,N_35609,N_38060);
and U44068 (N_44068,N_35586,N_37694);
nand U44069 (N_44069,N_39140,N_37990);
nand U44070 (N_44070,N_38675,N_37497);
and U44071 (N_44071,N_36519,N_36629);
or U44072 (N_44072,N_35036,N_38280);
nor U44073 (N_44073,N_38972,N_35593);
xnor U44074 (N_44074,N_35593,N_39756);
nand U44075 (N_44075,N_39634,N_37659);
nand U44076 (N_44076,N_35558,N_38247);
xnor U44077 (N_44077,N_36778,N_35673);
or U44078 (N_44078,N_37671,N_37465);
nor U44079 (N_44079,N_38239,N_35058);
or U44080 (N_44080,N_39382,N_35702);
or U44081 (N_44081,N_37920,N_38084);
or U44082 (N_44082,N_38953,N_37442);
and U44083 (N_44083,N_38430,N_36795);
or U44084 (N_44084,N_39940,N_38114);
or U44085 (N_44085,N_39556,N_35916);
nor U44086 (N_44086,N_35687,N_39270);
nand U44087 (N_44087,N_39857,N_38352);
or U44088 (N_44088,N_36912,N_35847);
nand U44089 (N_44089,N_36015,N_35081);
xnor U44090 (N_44090,N_37551,N_35492);
nor U44091 (N_44091,N_37924,N_35828);
xnor U44092 (N_44092,N_35467,N_35732);
nand U44093 (N_44093,N_37497,N_36290);
or U44094 (N_44094,N_39484,N_39464);
nor U44095 (N_44095,N_35402,N_38827);
and U44096 (N_44096,N_35119,N_36110);
xnor U44097 (N_44097,N_36361,N_37754);
xnor U44098 (N_44098,N_37278,N_37355);
nor U44099 (N_44099,N_36447,N_38359);
nor U44100 (N_44100,N_38865,N_36690);
xnor U44101 (N_44101,N_38533,N_35478);
nor U44102 (N_44102,N_36450,N_37239);
and U44103 (N_44103,N_37277,N_36229);
and U44104 (N_44104,N_36756,N_36200);
xor U44105 (N_44105,N_37515,N_38909);
nand U44106 (N_44106,N_39152,N_37577);
or U44107 (N_44107,N_35057,N_39206);
and U44108 (N_44108,N_38328,N_37461);
nand U44109 (N_44109,N_38590,N_39638);
nand U44110 (N_44110,N_36310,N_38535);
or U44111 (N_44111,N_36935,N_38935);
nand U44112 (N_44112,N_36997,N_39682);
nand U44113 (N_44113,N_37755,N_36315);
nor U44114 (N_44114,N_39173,N_38503);
nand U44115 (N_44115,N_37395,N_39426);
and U44116 (N_44116,N_35956,N_38181);
or U44117 (N_44117,N_39463,N_37096);
or U44118 (N_44118,N_38493,N_38082);
xor U44119 (N_44119,N_35043,N_37357);
nor U44120 (N_44120,N_38872,N_37990);
nor U44121 (N_44121,N_37323,N_37747);
nand U44122 (N_44122,N_35186,N_35009);
xor U44123 (N_44123,N_38722,N_38070);
or U44124 (N_44124,N_35917,N_35845);
xor U44125 (N_44125,N_38102,N_37287);
nand U44126 (N_44126,N_38675,N_37468);
nand U44127 (N_44127,N_36977,N_38695);
and U44128 (N_44128,N_38664,N_37426);
nand U44129 (N_44129,N_37020,N_35968);
and U44130 (N_44130,N_36971,N_35544);
nor U44131 (N_44131,N_38524,N_35395);
nor U44132 (N_44132,N_35849,N_37447);
nand U44133 (N_44133,N_36383,N_36509);
nand U44134 (N_44134,N_37448,N_38990);
and U44135 (N_44135,N_36658,N_35902);
and U44136 (N_44136,N_36457,N_37117);
nand U44137 (N_44137,N_39918,N_39202);
nor U44138 (N_44138,N_39710,N_35514);
or U44139 (N_44139,N_39921,N_39666);
or U44140 (N_44140,N_36378,N_35447);
nand U44141 (N_44141,N_39096,N_35080);
nor U44142 (N_44142,N_39885,N_36460);
nand U44143 (N_44143,N_37010,N_38913);
or U44144 (N_44144,N_36796,N_35386);
and U44145 (N_44145,N_35082,N_37333);
or U44146 (N_44146,N_37409,N_37745);
or U44147 (N_44147,N_35324,N_35738);
nor U44148 (N_44148,N_37984,N_37391);
or U44149 (N_44149,N_38156,N_37166);
or U44150 (N_44150,N_36150,N_39511);
and U44151 (N_44151,N_39868,N_38196);
and U44152 (N_44152,N_39339,N_37533);
or U44153 (N_44153,N_35299,N_35961);
nor U44154 (N_44154,N_36736,N_38173);
xnor U44155 (N_44155,N_38739,N_39777);
nor U44156 (N_44156,N_35515,N_38505);
nand U44157 (N_44157,N_38944,N_36540);
and U44158 (N_44158,N_35026,N_36668);
xor U44159 (N_44159,N_37571,N_36499);
nor U44160 (N_44160,N_37489,N_37175);
xnor U44161 (N_44161,N_35281,N_36176);
nand U44162 (N_44162,N_38601,N_35461);
nor U44163 (N_44163,N_36493,N_35045);
nand U44164 (N_44164,N_36146,N_39555);
xor U44165 (N_44165,N_37331,N_35892);
or U44166 (N_44166,N_38619,N_39137);
nor U44167 (N_44167,N_39260,N_36631);
and U44168 (N_44168,N_36610,N_37131);
nor U44169 (N_44169,N_35541,N_35853);
nand U44170 (N_44170,N_37310,N_38421);
and U44171 (N_44171,N_35368,N_39240);
and U44172 (N_44172,N_39578,N_37648);
nor U44173 (N_44173,N_37023,N_35750);
or U44174 (N_44174,N_35889,N_39939);
or U44175 (N_44175,N_36669,N_38544);
nor U44176 (N_44176,N_35205,N_37483);
and U44177 (N_44177,N_39593,N_39206);
xor U44178 (N_44178,N_36176,N_37271);
and U44179 (N_44179,N_36745,N_35927);
xor U44180 (N_44180,N_38118,N_36981);
or U44181 (N_44181,N_39750,N_36428);
or U44182 (N_44182,N_37686,N_37408);
nor U44183 (N_44183,N_38086,N_38517);
and U44184 (N_44184,N_36111,N_38056);
nor U44185 (N_44185,N_37713,N_39408);
nand U44186 (N_44186,N_36325,N_38124);
or U44187 (N_44187,N_39901,N_37948);
or U44188 (N_44188,N_38772,N_39622);
and U44189 (N_44189,N_39773,N_36115);
nand U44190 (N_44190,N_38633,N_36772);
and U44191 (N_44191,N_35071,N_37259);
nand U44192 (N_44192,N_36830,N_36938);
nor U44193 (N_44193,N_37732,N_36298);
xor U44194 (N_44194,N_38100,N_38127);
nor U44195 (N_44195,N_37753,N_39582);
nand U44196 (N_44196,N_36837,N_36320);
and U44197 (N_44197,N_35227,N_39879);
nor U44198 (N_44198,N_36585,N_36816);
nor U44199 (N_44199,N_37867,N_39067);
nand U44200 (N_44200,N_39807,N_37317);
and U44201 (N_44201,N_36483,N_37690);
and U44202 (N_44202,N_37084,N_37357);
xnor U44203 (N_44203,N_36904,N_39125);
nor U44204 (N_44204,N_36397,N_35557);
nand U44205 (N_44205,N_35731,N_37223);
or U44206 (N_44206,N_36398,N_36749);
nor U44207 (N_44207,N_39621,N_36360);
nor U44208 (N_44208,N_39968,N_38725);
or U44209 (N_44209,N_39301,N_37441);
or U44210 (N_44210,N_37575,N_39108);
or U44211 (N_44211,N_36283,N_36913);
nand U44212 (N_44212,N_36252,N_36535);
or U44213 (N_44213,N_39400,N_37136);
or U44214 (N_44214,N_39953,N_36725);
xor U44215 (N_44215,N_39753,N_37759);
nand U44216 (N_44216,N_36368,N_35774);
and U44217 (N_44217,N_36266,N_37204);
nor U44218 (N_44218,N_39887,N_36585);
or U44219 (N_44219,N_38518,N_37698);
nand U44220 (N_44220,N_38698,N_35827);
or U44221 (N_44221,N_38728,N_38270);
nor U44222 (N_44222,N_35864,N_35468);
xor U44223 (N_44223,N_35410,N_39466);
and U44224 (N_44224,N_35548,N_36599);
nand U44225 (N_44225,N_39706,N_36110);
or U44226 (N_44226,N_37155,N_39710);
or U44227 (N_44227,N_39966,N_35028);
or U44228 (N_44228,N_36270,N_36553);
and U44229 (N_44229,N_39064,N_39050);
nand U44230 (N_44230,N_35775,N_35023);
nand U44231 (N_44231,N_35504,N_38078);
nand U44232 (N_44232,N_37421,N_37935);
xor U44233 (N_44233,N_36671,N_37593);
and U44234 (N_44234,N_36062,N_39319);
or U44235 (N_44235,N_37524,N_38719);
or U44236 (N_44236,N_37291,N_35837);
and U44237 (N_44237,N_36329,N_38584);
nor U44238 (N_44238,N_36397,N_36944);
nor U44239 (N_44239,N_38540,N_37710);
xor U44240 (N_44240,N_35292,N_35705);
xnor U44241 (N_44241,N_38181,N_37215);
or U44242 (N_44242,N_35288,N_39840);
xor U44243 (N_44243,N_37188,N_35844);
and U44244 (N_44244,N_37094,N_39206);
or U44245 (N_44245,N_36353,N_39681);
or U44246 (N_44246,N_36509,N_35942);
xor U44247 (N_44247,N_36194,N_39089);
xnor U44248 (N_44248,N_39818,N_39634);
or U44249 (N_44249,N_36347,N_37290);
xnor U44250 (N_44250,N_35394,N_36700);
nor U44251 (N_44251,N_39802,N_37783);
nor U44252 (N_44252,N_36888,N_35751);
or U44253 (N_44253,N_36378,N_35150);
or U44254 (N_44254,N_39973,N_36928);
or U44255 (N_44255,N_39028,N_37572);
nand U44256 (N_44256,N_36420,N_37491);
nor U44257 (N_44257,N_36617,N_36286);
nor U44258 (N_44258,N_36873,N_36983);
nor U44259 (N_44259,N_39719,N_39983);
or U44260 (N_44260,N_36663,N_37892);
nor U44261 (N_44261,N_37501,N_37097);
nor U44262 (N_44262,N_35249,N_39611);
nor U44263 (N_44263,N_35494,N_39303);
xor U44264 (N_44264,N_39025,N_36929);
or U44265 (N_44265,N_38588,N_37312);
xnor U44266 (N_44266,N_36416,N_35836);
or U44267 (N_44267,N_35442,N_36069);
nor U44268 (N_44268,N_39441,N_35374);
nand U44269 (N_44269,N_39016,N_36325);
nand U44270 (N_44270,N_38480,N_35663);
or U44271 (N_44271,N_35099,N_35751);
nand U44272 (N_44272,N_39131,N_38517);
xnor U44273 (N_44273,N_37714,N_38374);
xor U44274 (N_44274,N_35796,N_36799);
nor U44275 (N_44275,N_37088,N_36707);
or U44276 (N_44276,N_39140,N_37550);
xor U44277 (N_44277,N_35103,N_36689);
xnor U44278 (N_44278,N_39898,N_39026);
xor U44279 (N_44279,N_38056,N_37972);
xor U44280 (N_44280,N_38322,N_39661);
or U44281 (N_44281,N_37841,N_37787);
or U44282 (N_44282,N_36110,N_36778);
nand U44283 (N_44283,N_37115,N_37559);
or U44284 (N_44284,N_37807,N_38252);
nand U44285 (N_44285,N_37829,N_35435);
xnor U44286 (N_44286,N_38227,N_38753);
nand U44287 (N_44287,N_39946,N_39372);
nand U44288 (N_44288,N_38199,N_36139);
nand U44289 (N_44289,N_36908,N_38858);
nand U44290 (N_44290,N_35731,N_35097);
nand U44291 (N_44291,N_38540,N_35107);
or U44292 (N_44292,N_38502,N_38180);
and U44293 (N_44293,N_39944,N_35205);
nand U44294 (N_44294,N_37867,N_35963);
and U44295 (N_44295,N_39168,N_38093);
nor U44296 (N_44296,N_36915,N_37074);
or U44297 (N_44297,N_36847,N_35992);
and U44298 (N_44298,N_35931,N_38842);
and U44299 (N_44299,N_38510,N_36528);
xnor U44300 (N_44300,N_37108,N_38318);
or U44301 (N_44301,N_36464,N_36714);
and U44302 (N_44302,N_38295,N_39580);
nand U44303 (N_44303,N_38556,N_38349);
nand U44304 (N_44304,N_38081,N_37044);
nand U44305 (N_44305,N_39968,N_37355);
xor U44306 (N_44306,N_36586,N_39969);
xor U44307 (N_44307,N_38523,N_37715);
nor U44308 (N_44308,N_35133,N_37755);
or U44309 (N_44309,N_39298,N_39080);
and U44310 (N_44310,N_37913,N_37117);
xnor U44311 (N_44311,N_36942,N_37427);
and U44312 (N_44312,N_36200,N_38273);
xor U44313 (N_44313,N_37839,N_37610);
or U44314 (N_44314,N_38451,N_38780);
nor U44315 (N_44315,N_37990,N_39256);
nand U44316 (N_44316,N_38804,N_38656);
or U44317 (N_44317,N_36516,N_35078);
or U44318 (N_44318,N_36800,N_39194);
nor U44319 (N_44319,N_39715,N_38485);
xor U44320 (N_44320,N_37414,N_39780);
nor U44321 (N_44321,N_38684,N_36968);
or U44322 (N_44322,N_35292,N_37594);
or U44323 (N_44323,N_35314,N_38541);
and U44324 (N_44324,N_38852,N_38848);
xor U44325 (N_44325,N_38856,N_36255);
or U44326 (N_44326,N_37144,N_39227);
xnor U44327 (N_44327,N_36342,N_38127);
nand U44328 (N_44328,N_37099,N_38756);
nand U44329 (N_44329,N_39577,N_37458);
and U44330 (N_44330,N_39828,N_37887);
or U44331 (N_44331,N_37254,N_37768);
nor U44332 (N_44332,N_37044,N_39711);
and U44333 (N_44333,N_36850,N_38718);
nand U44334 (N_44334,N_39025,N_37904);
or U44335 (N_44335,N_38747,N_37130);
xnor U44336 (N_44336,N_35234,N_36113);
nor U44337 (N_44337,N_36496,N_35710);
xor U44338 (N_44338,N_36516,N_37689);
nand U44339 (N_44339,N_35832,N_35043);
nor U44340 (N_44340,N_39693,N_35793);
nand U44341 (N_44341,N_38261,N_38154);
or U44342 (N_44342,N_35347,N_39793);
or U44343 (N_44343,N_35222,N_38375);
nor U44344 (N_44344,N_35948,N_35787);
or U44345 (N_44345,N_37468,N_36584);
nand U44346 (N_44346,N_36842,N_36938);
nand U44347 (N_44347,N_35218,N_36384);
and U44348 (N_44348,N_39271,N_35371);
or U44349 (N_44349,N_35167,N_36494);
xnor U44350 (N_44350,N_38834,N_38627);
nor U44351 (N_44351,N_37539,N_37190);
xor U44352 (N_44352,N_35107,N_38989);
nor U44353 (N_44353,N_36398,N_37782);
nor U44354 (N_44354,N_39757,N_36391);
nor U44355 (N_44355,N_39184,N_38984);
xnor U44356 (N_44356,N_37864,N_35786);
xor U44357 (N_44357,N_36608,N_35559);
and U44358 (N_44358,N_35931,N_37762);
and U44359 (N_44359,N_35386,N_39507);
or U44360 (N_44360,N_38342,N_35717);
or U44361 (N_44361,N_36619,N_37274);
or U44362 (N_44362,N_36065,N_39172);
nor U44363 (N_44363,N_35090,N_37845);
nand U44364 (N_44364,N_35260,N_36210);
nand U44365 (N_44365,N_38155,N_37161);
or U44366 (N_44366,N_36408,N_37506);
xnor U44367 (N_44367,N_36770,N_39172);
xor U44368 (N_44368,N_39590,N_37666);
or U44369 (N_44369,N_35765,N_39847);
or U44370 (N_44370,N_36351,N_37515);
and U44371 (N_44371,N_35319,N_37222);
xor U44372 (N_44372,N_37324,N_36512);
nor U44373 (N_44373,N_35857,N_39860);
nand U44374 (N_44374,N_35907,N_35075);
or U44375 (N_44375,N_39113,N_38179);
nand U44376 (N_44376,N_36885,N_38292);
nand U44377 (N_44377,N_38364,N_37340);
and U44378 (N_44378,N_39257,N_38788);
nand U44379 (N_44379,N_37764,N_36228);
or U44380 (N_44380,N_38290,N_35690);
or U44381 (N_44381,N_36573,N_37263);
and U44382 (N_44382,N_39434,N_38876);
and U44383 (N_44383,N_38598,N_36407);
nand U44384 (N_44384,N_39243,N_36893);
nand U44385 (N_44385,N_38277,N_37659);
xnor U44386 (N_44386,N_38275,N_39860);
xnor U44387 (N_44387,N_37925,N_37245);
or U44388 (N_44388,N_38066,N_39254);
nand U44389 (N_44389,N_37123,N_35529);
nand U44390 (N_44390,N_37545,N_39556);
nand U44391 (N_44391,N_35283,N_35377);
nor U44392 (N_44392,N_37323,N_36464);
and U44393 (N_44393,N_38132,N_35416);
or U44394 (N_44394,N_35719,N_39473);
nor U44395 (N_44395,N_39463,N_36903);
or U44396 (N_44396,N_36714,N_35239);
or U44397 (N_44397,N_38879,N_37036);
and U44398 (N_44398,N_37456,N_35134);
nor U44399 (N_44399,N_37376,N_35398);
or U44400 (N_44400,N_37070,N_38227);
nor U44401 (N_44401,N_39326,N_38719);
or U44402 (N_44402,N_39333,N_35817);
nor U44403 (N_44403,N_36707,N_39492);
and U44404 (N_44404,N_37732,N_35822);
xor U44405 (N_44405,N_39073,N_39475);
nor U44406 (N_44406,N_38403,N_36755);
nor U44407 (N_44407,N_36720,N_39544);
and U44408 (N_44408,N_38841,N_35833);
xor U44409 (N_44409,N_36029,N_35635);
xnor U44410 (N_44410,N_36261,N_39170);
or U44411 (N_44411,N_36830,N_38831);
and U44412 (N_44412,N_39302,N_38912);
and U44413 (N_44413,N_35739,N_35806);
nor U44414 (N_44414,N_39480,N_35367);
or U44415 (N_44415,N_39196,N_37096);
nor U44416 (N_44416,N_35242,N_38629);
or U44417 (N_44417,N_37057,N_37998);
and U44418 (N_44418,N_36560,N_39082);
xnor U44419 (N_44419,N_37491,N_35518);
nor U44420 (N_44420,N_36964,N_38023);
nand U44421 (N_44421,N_36672,N_35030);
xnor U44422 (N_44422,N_38153,N_35258);
nor U44423 (N_44423,N_36772,N_36247);
and U44424 (N_44424,N_38357,N_35742);
nand U44425 (N_44425,N_36744,N_39430);
or U44426 (N_44426,N_38789,N_37386);
nand U44427 (N_44427,N_36867,N_38361);
or U44428 (N_44428,N_37006,N_37803);
xor U44429 (N_44429,N_36127,N_38354);
nand U44430 (N_44430,N_37032,N_36833);
nand U44431 (N_44431,N_39068,N_38534);
nand U44432 (N_44432,N_39422,N_36065);
nor U44433 (N_44433,N_35419,N_38121);
nand U44434 (N_44434,N_36463,N_39222);
xor U44435 (N_44435,N_38849,N_38998);
and U44436 (N_44436,N_36134,N_38892);
or U44437 (N_44437,N_37619,N_36469);
xor U44438 (N_44438,N_38819,N_39468);
xnor U44439 (N_44439,N_39133,N_39322);
nor U44440 (N_44440,N_39225,N_36472);
and U44441 (N_44441,N_36066,N_35648);
nor U44442 (N_44442,N_35178,N_39229);
nor U44443 (N_44443,N_37793,N_39923);
or U44444 (N_44444,N_35072,N_38553);
nor U44445 (N_44445,N_35106,N_38338);
or U44446 (N_44446,N_39662,N_35970);
nand U44447 (N_44447,N_36626,N_39072);
and U44448 (N_44448,N_36863,N_36421);
nor U44449 (N_44449,N_38331,N_36243);
and U44450 (N_44450,N_36675,N_36495);
nor U44451 (N_44451,N_35235,N_36093);
or U44452 (N_44452,N_38665,N_37894);
and U44453 (N_44453,N_36194,N_35180);
and U44454 (N_44454,N_35097,N_37298);
or U44455 (N_44455,N_37394,N_36655);
xnor U44456 (N_44456,N_37345,N_38157);
xor U44457 (N_44457,N_35272,N_35211);
nand U44458 (N_44458,N_37938,N_36527);
nor U44459 (N_44459,N_38727,N_36721);
nand U44460 (N_44460,N_37865,N_35732);
or U44461 (N_44461,N_35814,N_39065);
or U44462 (N_44462,N_37895,N_37445);
or U44463 (N_44463,N_35826,N_39753);
and U44464 (N_44464,N_38874,N_38124);
nor U44465 (N_44465,N_36293,N_38244);
nand U44466 (N_44466,N_38612,N_39127);
nor U44467 (N_44467,N_38604,N_36863);
nor U44468 (N_44468,N_38585,N_36932);
xnor U44469 (N_44469,N_37906,N_35673);
nor U44470 (N_44470,N_37075,N_37832);
nand U44471 (N_44471,N_36244,N_38071);
xor U44472 (N_44472,N_39565,N_37289);
xor U44473 (N_44473,N_38894,N_36203);
and U44474 (N_44474,N_38468,N_36113);
and U44475 (N_44475,N_38218,N_38473);
nand U44476 (N_44476,N_35833,N_35443);
nand U44477 (N_44477,N_38484,N_38688);
xor U44478 (N_44478,N_38501,N_39461);
nand U44479 (N_44479,N_35450,N_37140);
or U44480 (N_44480,N_35802,N_39241);
or U44481 (N_44481,N_37938,N_36089);
xnor U44482 (N_44482,N_36670,N_36022);
nand U44483 (N_44483,N_39486,N_36615);
and U44484 (N_44484,N_37918,N_37956);
nand U44485 (N_44485,N_38709,N_39345);
xor U44486 (N_44486,N_37058,N_35419);
or U44487 (N_44487,N_37506,N_35330);
nor U44488 (N_44488,N_36723,N_36934);
or U44489 (N_44489,N_37847,N_38423);
xnor U44490 (N_44490,N_38544,N_37114);
nor U44491 (N_44491,N_36530,N_38233);
nand U44492 (N_44492,N_38757,N_38875);
xor U44493 (N_44493,N_37672,N_35134);
nor U44494 (N_44494,N_38265,N_39257);
or U44495 (N_44495,N_38108,N_36748);
nand U44496 (N_44496,N_37693,N_35846);
or U44497 (N_44497,N_38544,N_36278);
or U44498 (N_44498,N_36636,N_37422);
nand U44499 (N_44499,N_35180,N_35079);
xor U44500 (N_44500,N_35874,N_35722);
or U44501 (N_44501,N_35908,N_36934);
and U44502 (N_44502,N_37406,N_37481);
nor U44503 (N_44503,N_35690,N_36004);
nor U44504 (N_44504,N_37719,N_36751);
nor U44505 (N_44505,N_35765,N_37504);
nand U44506 (N_44506,N_37630,N_38675);
or U44507 (N_44507,N_38622,N_36111);
xor U44508 (N_44508,N_36193,N_39090);
nor U44509 (N_44509,N_38271,N_35480);
nor U44510 (N_44510,N_35334,N_38884);
and U44511 (N_44511,N_36986,N_38244);
nor U44512 (N_44512,N_36596,N_35050);
nand U44513 (N_44513,N_35843,N_39465);
and U44514 (N_44514,N_35707,N_36810);
nand U44515 (N_44515,N_39868,N_38077);
and U44516 (N_44516,N_36405,N_38023);
and U44517 (N_44517,N_37005,N_35918);
and U44518 (N_44518,N_39076,N_39749);
and U44519 (N_44519,N_38615,N_39814);
nor U44520 (N_44520,N_35553,N_35160);
or U44521 (N_44521,N_35924,N_38133);
and U44522 (N_44522,N_35896,N_36460);
or U44523 (N_44523,N_38331,N_39825);
or U44524 (N_44524,N_39903,N_36899);
nand U44525 (N_44525,N_37182,N_37176);
nor U44526 (N_44526,N_36718,N_35381);
nand U44527 (N_44527,N_35303,N_38831);
or U44528 (N_44528,N_35653,N_37163);
nor U44529 (N_44529,N_38418,N_37345);
xnor U44530 (N_44530,N_38640,N_39898);
and U44531 (N_44531,N_35688,N_35790);
xnor U44532 (N_44532,N_39432,N_37728);
and U44533 (N_44533,N_36211,N_36899);
or U44534 (N_44534,N_36793,N_36973);
and U44535 (N_44535,N_36120,N_39575);
nand U44536 (N_44536,N_38315,N_38819);
or U44537 (N_44537,N_39993,N_39032);
nor U44538 (N_44538,N_39315,N_38509);
nor U44539 (N_44539,N_39149,N_37837);
xor U44540 (N_44540,N_38903,N_36256);
nor U44541 (N_44541,N_36353,N_39962);
and U44542 (N_44542,N_39305,N_38528);
nand U44543 (N_44543,N_39017,N_36619);
and U44544 (N_44544,N_35421,N_39102);
or U44545 (N_44545,N_35543,N_35802);
and U44546 (N_44546,N_39811,N_38418);
and U44547 (N_44547,N_36926,N_38291);
or U44548 (N_44548,N_36061,N_39654);
or U44549 (N_44549,N_35124,N_36611);
nand U44550 (N_44550,N_35683,N_35443);
xnor U44551 (N_44551,N_38905,N_39625);
or U44552 (N_44552,N_39613,N_38577);
and U44553 (N_44553,N_39760,N_37322);
nand U44554 (N_44554,N_36520,N_35408);
and U44555 (N_44555,N_39141,N_36646);
or U44556 (N_44556,N_38364,N_37039);
nor U44557 (N_44557,N_39550,N_37681);
nor U44558 (N_44558,N_39147,N_35323);
or U44559 (N_44559,N_37546,N_37504);
and U44560 (N_44560,N_37049,N_38537);
or U44561 (N_44561,N_39571,N_39806);
nor U44562 (N_44562,N_39326,N_36816);
nor U44563 (N_44563,N_36887,N_39484);
or U44564 (N_44564,N_35393,N_35478);
nand U44565 (N_44565,N_37511,N_37279);
nand U44566 (N_44566,N_35037,N_38537);
or U44567 (N_44567,N_39412,N_39869);
or U44568 (N_44568,N_35292,N_35531);
nand U44569 (N_44569,N_35541,N_38875);
nor U44570 (N_44570,N_35594,N_36581);
or U44571 (N_44571,N_35271,N_36559);
xnor U44572 (N_44572,N_37510,N_35640);
nand U44573 (N_44573,N_38630,N_37237);
nand U44574 (N_44574,N_35188,N_38740);
xnor U44575 (N_44575,N_37839,N_38726);
or U44576 (N_44576,N_38776,N_38051);
nor U44577 (N_44577,N_39427,N_37447);
and U44578 (N_44578,N_37121,N_38586);
nand U44579 (N_44579,N_36452,N_37698);
nor U44580 (N_44580,N_37656,N_38623);
nand U44581 (N_44581,N_35695,N_37188);
or U44582 (N_44582,N_39145,N_38914);
nand U44583 (N_44583,N_35291,N_38962);
or U44584 (N_44584,N_37567,N_39635);
nand U44585 (N_44585,N_38603,N_39582);
or U44586 (N_44586,N_36679,N_36969);
nand U44587 (N_44587,N_35235,N_37420);
and U44588 (N_44588,N_39546,N_35364);
and U44589 (N_44589,N_39216,N_37293);
nor U44590 (N_44590,N_39898,N_38432);
and U44591 (N_44591,N_38843,N_38139);
nand U44592 (N_44592,N_39949,N_39441);
nor U44593 (N_44593,N_35294,N_35404);
nor U44594 (N_44594,N_38242,N_35410);
nor U44595 (N_44595,N_39470,N_39636);
or U44596 (N_44596,N_36490,N_38044);
xnor U44597 (N_44597,N_38548,N_38702);
nor U44598 (N_44598,N_36545,N_35755);
xor U44599 (N_44599,N_38293,N_38457);
and U44600 (N_44600,N_38111,N_39727);
or U44601 (N_44601,N_38351,N_35571);
or U44602 (N_44602,N_35027,N_36142);
nand U44603 (N_44603,N_39973,N_39928);
and U44604 (N_44604,N_37932,N_37606);
nand U44605 (N_44605,N_38983,N_38752);
nor U44606 (N_44606,N_37552,N_36376);
and U44607 (N_44607,N_36660,N_37092);
xnor U44608 (N_44608,N_37370,N_39035);
or U44609 (N_44609,N_36498,N_35844);
nor U44610 (N_44610,N_38835,N_37544);
and U44611 (N_44611,N_39305,N_36749);
nand U44612 (N_44612,N_37879,N_35373);
nand U44613 (N_44613,N_36804,N_35580);
nor U44614 (N_44614,N_38320,N_37626);
nand U44615 (N_44615,N_38782,N_38061);
or U44616 (N_44616,N_38874,N_35502);
nor U44617 (N_44617,N_37763,N_38519);
nor U44618 (N_44618,N_37794,N_36348);
nor U44619 (N_44619,N_37058,N_39387);
xor U44620 (N_44620,N_39301,N_38390);
or U44621 (N_44621,N_35540,N_36772);
or U44622 (N_44622,N_38057,N_39563);
nand U44623 (N_44623,N_39745,N_36461);
or U44624 (N_44624,N_38768,N_37141);
nand U44625 (N_44625,N_38065,N_37908);
nand U44626 (N_44626,N_37490,N_35071);
nor U44627 (N_44627,N_37193,N_36406);
or U44628 (N_44628,N_35426,N_38108);
nand U44629 (N_44629,N_37656,N_35301);
xor U44630 (N_44630,N_36167,N_39519);
nand U44631 (N_44631,N_36761,N_38464);
nand U44632 (N_44632,N_39792,N_35604);
or U44633 (N_44633,N_38556,N_38821);
or U44634 (N_44634,N_35445,N_35142);
xor U44635 (N_44635,N_35608,N_36281);
nor U44636 (N_44636,N_39410,N_36137);
or U44637 (N_44637,N_38128,N_39064);
nor U44638 (N_44638,N_37088,N_35286);
or U44639 (N_44639,N_36879,N_39547);
xor U44640 (N_44640,N_39088,N_39426);
nand U44641 (N_44641,N_38219,N_39514);
nand U44642 (N_44642,N_39649,N_36285);
and U44643 (N_44643,N_37360,N_39640);
xnor U44644 (N_44644,N_38259,N_38471);
or U44645 (N_44645,N_38007,N_39698);
nor U44646 (N_44646,N_35868,N_35063);
nand U44647 (N_44647,N_38401,N_38526);
or U44648 (N_44648,N_39708,N_35721);
nand U44649 (N_44649,N_38975,N_38421);
or U44650 (N_44650,N_37045,N_37150);
nor U44651 (N_44651,N_38132,N_38221);
xor U44652 (N_44652,N_36660,N_36392);
or U44653 (N_44653,N_39511,N_38707);
xnor U44654 (N_44654,N_35075,N_38167);
xnor U44655 (N_44655,N_39676,N_39996);
and U44656 (N_44656,N_38466,N_38662);
nor U44657 (N_44657,N_36326,N_37894);
nor U44658 (N_44658,N_39779,N_39064);
nand U44659 (N_44659,N_37327,N_35825);
nand U44660 (N_44660,N_36910,N_38968);
xnor U44661 (N_44661,N_36114,N_36051);
or U44662 (N_44662,N_38835,N_39213);
and U44663 (N_44663,N_39551,N_35970);
or U44664 (N_44664,N_35968,N_36770);
or U44665 (N_44665,N_35897,N_39287);
or U44666 (N_44666,N_38421,N_38071);
nor U44667 (N_44667,N_38095,N_36866);
or U44668 (N_44668,N_38996,N_39969);
nand U44669 (N_44669,N_37475,N_37795);
and U44670 (N_44670,N_39844,N_38587);
nor U44671 (N_44671,N_35590,N_36562);
or U44672 (N_44672,N_38483,N_38899);
and U44673 (N_44673,N_36011,N_35952);
xor U44674 (N_44674,N_39848,N_38557);
or U44675 (N_44675,N_35982,N_38449);
xor U44676 (N_44676,N_39982,N_36926);
nor U44677 (N_44677,N_38501,N_36776);
xnor U44678 (N_44678,N_38585,N_39563);
nor U44679 (N_44679,N_35965,N_37249);
and U44680 (N_44680,N_38197,N_37931);
and U44681 (N_44681,N_38656,N_38186);
or U44682 (N_44682,N_37438,N_36562);
xnor U44683 (N_44683,N_37821,N_37835);
nand U44684 (N_44684,N_37924,N_35408);
xnor U44685 (N_44685,N_37370,N_36814);
and U44686 (N_44686,N_37667,N_38087);
and U44687 (N_44687,N_39416,N_36124);
nand U44688 (N_44688,N_36237,N_37461);
or U44689 (N_44689,N_35231,N_38694);
and U44690 (N_44690,N_35835,N_37413);
and U44691 (N_44691,N_38358,N_38885);
nor U44692 (N_44692,N_39443,N_37869);
xnor U44693 (N_44693,N_37179,N_38620);
and U44694 (N_44694,N_38980,N_39564);
nand U44695 (N_44695,N_35466,N_39957);
and U44696 (N_44696,N_38148,N_37067);
xnor U44697 (N_44697,N_35530,N_36663);
nand U44698 (N_44698,N_36645,N_37481);
nand U44699 (N_44699,N_39205,N_36870);
and U44700 (N_44700,N_36164,N_37992);
and U44701 (N_44701,N_35685,N_37490);
or U44702 (N_44702,N_38061,N_36341);
xor U44703 (N_44703,N_38419,N_39170);
or U44704 (N_44704,N_38584,N_38891);
nor U44705 (N_44705,N_36041,N_39315);
nor U44706 (N_44706,N_35089,N_39250);
and U44707 (N_44707,N_38078,N_39621);
and U44708 (N_44708,N_36626,N_37799);
xnor U44709 (N_44709,N_35057,N_39799);
or U44710 (N_44710,N_39099,N_38090);
and U44711 (N_44711,N_37075,N_37204);
nand U44712 (N_44712,N_39282,N_36786);
or U44713 (N_44713,N_39939,N_39057);
or U44714 (N_44714,N_37582,N_37874);
xor U44715 (N_44715,N_37867,N_35660);
xnor U44716 (N_44716,N_37499,N_39582);
xor U44717 (N_44717,N_37378,N_38491);
or U44718 (N_44718,N_37684,N_35689);
or U44719 (N_44719,N_38761,N_36503);
nand U44720 (N_44720,N_35575,N_35693);
nand U44721 (N_44721,N_39030,N_35399);
nor U44722 (N_44722,N_38832,N_39143);
xor U44723 (N_44723,N_35572,N_37626);
or U44724 (N_44724,N_37884,N_35067);
nor U44725 (N_44725,N_37196,N_38486);
xnor U44726 (N_44726,N_37168,N_39151);
xnor U44727 (N_44727,N_39157,N_39519);
xor U44728 (N_44728,N_36304,N_36661);
and U44729 (N_44729,N_39638,N_39340);
nor U44730 (N_44730,N_35226,N_38576);
nand U44731 (N_44731,N_38737,N_37432);
xor U44732 (N_44732,N_35406,N_35343);
or U44733 (N_44733,N_37506,N_35466);
nor U44734 (N_44734,N_35563,N_39370);
nor U44735 (N_44735,N_39389,N_36837);
xnor U44736 (N_44736,N_39327,N_35773);
nand U44737 (N_44737,N_39733,N_37390);
nand U44738 (N_44738,N_38870,N_38692);
xnor U44739 (N_44739,N_37934,N_37778);
nor U44740 (N_44740,N_37064,N_37999);
nor U44741 (N_44741,N_37608,N_39238);
nor U44742 (N_44742,N_39120,N_38269);
nor U44743 (N_44743,N_36584,N_36488);
nand U44744 (N_44744,N_35007,N_37545);
or U44745 (N_44745,N_35543,N_38711);
and U44746 (N_44746,N_35357,N_39787);
or U44747 (N_44747,N_37005,N_38382);
nand U44748 (N_44748,N_38094,N_38401);
and U44749 (N_44749,N_35618,N_36202);
nor U44750 (N_44750,N_35970,N_38788);
nand U44751 (N_44751,N_37528,N_36596);
xnor U44752 (N_44752,N_39283,N_37817);
and U44753 (N_44753,N_35887,N_35309);
xor U44754 (N_44754,N_35514,N_39802);
nor U44755 (N_44755,N_38153,N_38697);
and U44756 (N_44756,N_38815,N_39399);
or U44757 (N_44757,N_36385,N_37119);
and U44758 (N_44758,N_37524,N_39043);
nor U44759 (N_44759,N_38284,N_36519);
xor U44760 (N_44760,N_39441,N_39941);
nand U44761 (N_44761,N_39670,N_35220);
xnor U44762 (N_44762,N_37917,N_35669);
nor U44763 (N_44763,N_36961,N_38686);
and U44764 (N_44764,N_35792,N_39789);
and U44765 (N_44765,N_36553,N_38429);
xor U44766 (N_44766,N_39432,N_36234);
and U44767 (N_44767,N_38226,N_35970);
nand U44768 (N_44768,N_39178,N_35726);
nand U44769 (N_44769,N_35661,N_39454);
xor U44770 (N_44770,N_37221,N_39770);
nand U44771 (N_44771,N_37225,N_37655);
nand U44772 (N_44772,N_37644,N_38493);
nor U44773 (N_44773,N_38428,N_38232);
nand U44774 (N_44774,N_38942,N_36198);
xnor U44775 (N_44775,N_38801,N_38794);
nor U44776 (N_44776,N_37824,N_39851);
and U44777 (N_44777,N_37084,N_36705);
nand U44778 (N_44778,N_38997,N_36189);
nor U44779 (N_44779,N_38599,N_35161);
xor U44780 (N_44780,N_35718,N_38080);
or U44781 (N_44781,N_37611,N_39075);
nor U44782 (N_44782,N_35487,N_36650);
or U44783 (N_44783,N_38947,N_37905);
xnor U44784 (N_44784,N_39004,N_38300);
nor U44785 (N_44785,N_37313,N_37740);
and U44786 (N_44786,N_39404,N_39814);
and U44787 (N_44787,N_36337,N_36647);
nor U44788 (N_44788,N_35632,N_38976);
nor U44789 (N_44789,N_36346,N_35455);
nor U44790 (N_44790,N_39130,N_38587);
nor U44791 (N_44791,N_35491,N_38275);
nor U44792 (N_44792,N_37984,N_37722);
xor U44793 (N_44793,N_38299,N_36809);
nand U44794 (N_44794,N_36148,N_37601);
and U44795 (N_44795,N_38496,N_35740);
nor U44796 (N_44796,N_38961,N_36828);
xnor U44797 (N_44797,N_39758,N_36476);
nor U44798 (N_44798,N_38769,N_35301);
or U44799 (N_44799,N_36576,N_38636);
xor U44800 (N_44800,N_37364,N_39371);
nand U44801 (N_44801,N_38176,N_36308);
xnor U44802 (N_44802,N_39136,N_38341);
nor U44803 (N_44803,N_35674,N_36657);
or U44804 (N_44804,N_39599,N_37679);
and U44805 (N_44805,N_37532,N_38458);
nand U44806 (N_44806,N_39834,N_36389);
xor U44807 (N_44807,N_38194,N_36905);
and U44808 (N_44808,N_39912,N_39903);
or U44809 (N_44809,N_35639,N_36835);
nor U44810 (N_44810,N_35055,N_35293);
nand U44811 (N_44811,N_35561,N_38750);
nand U44812 (N_44812,N_36653,N_38820);
nor U44813 (N_44813,N_37348,N_36840);
or U44814 (N_44814,N_35916,N_39074);
and U44815 (N_44815,N_35752,N_37083);
nand U44816 (N_44816,N_36231,N_37195);
and U44817 (N_44817,N_38299,N_39676);
xnor U44818 (N_44818,N_35025,N_35682);
nand U44819 (N_44819,N_35276,N_37748);
or U44820 (N_44820,N_37679,N_36903);
or U44821 (N_44821,N_38965,N_37072);
or U44822 (N_44822,N_37674,N_36309);
and U44823 (N_44823,N_35500,N_35573);
or U44824 (N_44824,N_35788,N_36182);
or U44825 (N_44825,N_38858,N_38399);
xor U44826 (N_44826,N_36880,N_35083);
nor U44827 (N_44827,N_37534,N_38592);
xnor U44828 (N_44828,N_36880,N_39445);
nor U44829 (N_44829,N_37563,N_39138);
nor U44830 (N_44830,N_39623,N_36054);
and U44831 (N_44831,N_38620,N_35498);
nor U44832 (N_44832,N_37371,N_39520);
nand U44833 (N_44833,N_35092,N_39957);
xor U44834 (N_44834,N_38115,N_39248);
nor U44835 (N_44835,N_36153,N_38032);
nand U44836 (N_44836,N_37117,N_39931);
nor U44837 (N_44837,N_38286,N_36121);
xor U44838 (N_44838,N_39402,N_36866);
nand U44839 (N_44839,N_36054,N_39075);
xnor U44840 (N_44840,N_36427,N_37977);
nor U44841 (N_44841,N_36396,N_38621);
nor U44842 (N_44842,N_38847,N_38602);
xor U44843 (N_44843,N_35747,N_37437);
or U44844 (N_44844,N_35589,N_39973);
xor U44845 (N_44845,N_38496,N_37113);
nand U44846 (N_44846,N_39805,N_39862);
xor U44847 (N_44847,N_38804,N_36130);
xor U44848 (N_44848,N_38289,N_35383);
and U44849 (N_44849,N_37738,N_38692);
xnor U44850 (N_44850,N_39284,N_38554);
xnor U44851 (N_44851,N_39246,N_37784);
nor U44852 (N_44852,N_38239,N_36715);
and U44853 (N_44853,N_37110,N_39698);
nand U44854 (N_44854,N_35109,N_38172);
or U44855 (N_44855,N_39498,N_38289);
nand U44856 (N_44856,N_39924,N_37726);
xor U44857 (N_44857,N_39689,N_39867);
xor U44858 (N_44858,N_38745,N_38952);
nand U44859 (N_44859,N_39375,N_39876);
or U44860 (N_44860,N_35787,N_39727);
xnor U44861 (N_44861,N_39998,N_39610);
nand U44862 (N_44862,N_38573,N_39854);
or U44863 (N_44863,N_39719,N_35278);
xor U44864 (N_44864,N_37396,N_37147);
nand U44865 (N_44865,N_37820,N_37197);
and U44866 (N_44866,N_35049,N_37889);
xnor U44867 (N_44867,N_37787,N_36719);
and U44868 (N_44868,N_39884,N_36369);
and U44869 (N_44869,N_37444,N_36545);
and U44870 (N_44870,N_39062,N_36689);
and U44871 (N_44871,N_37304,N_35072);
or U44872 (N_44872,N_38664,N_38663);
and U44873 (N_44873,N_36719,N_35647);
and U44874 (N_44874,N_39165,N_35846);
xor U44875 (N_44875,N_36203,N_35956);
and U44876 (N_44876,N_35265,N_38499);
xor U44877 (N_44877,N_35629,N_36890);
or U44878 (N_44878,N_35311,N_37898);
and U44879 (N_44879,N_38149,N_38977);
or U44880 (N_44880,N_37876,N_37894);
xor U44881 (N_44881,N_35433,N_38611);
and U44882 (N_44882,N_35620,N_37809);
xor U44883 (N_44883,N_36419,N_35569);
nor U44884 (N_44884,N_36394,N_39951);
or U44885 (N_44885,N_35423,N_38647);
and U44886 (N_44886,N_39810,N_39498);
xor U44887 (N_44887,N_36268,N_39616);
nor U44888 (N_44888,N_37647,N_38487);
or U44889 (N_44889,N_39460,N_38437);
and U44890 (N_44890,N_37660,N_37374);
nor U44891 (N_44891,N_39449,N_38982);
and U44892 (N_44892,N_36208,N_37342);
xor U44893 (N_44893,N_37212,N_38555);
nor U44894 (N_44894,N_38247,N_38010);
and U44895 (N_44895,N_38513,N_38334);
nor U44896 (N_44896,N_37812,N_36521);
or U44897 (N_44897,N_38517,N_38775);
nor U44898 (N_44898,N_39523,N_38708);
xor U44899 (N_44899,N_39425,N_35403);
and U44900 (N_44900,N_37402,N_35539);
and U44901 (N_44901,N_36062,N_38350);
xnor U44902 (N_44902,N_39993,N_37937);
or U44903 (N_44903,N_37115,N_37915);
or U44904 (N_44904,N_35947,N_38000);
xnor U44905 (N_44905,N_38959,N_37016);
and U44906 (N_44906,N_38076,N_39988);
or U44907 (N_44907,N_36658,N_36567);
and U44908 (N_44908,N_38509,N_38168);
nand U44909 (N_44909,N_38471,N_39816);
or U44910 (N_44910,N_38108,N_36906);
nand U44911 (N_44911,N_38766,N_37672);
xnor U44912 (N_44912,N_36823,N_35167);
xor U44913 (N_44913,N_37019,N_39283);
and U44914 (N_44914,N_35383,N_36060);
and U44915 (N_44915,N_36212,N_35929);
nor U44916 (N_44916,N_36202,N_39129);
nor U44917 (N_44917,N_37658,N_37174);
and U44918 (N_44918,N_39836,N_37578);
or U44919 (N_44919,N_36907,N_35927);
or U44920 (N_44920,N_39205,N_36390);
and U44921 (N_44921,N_35615,N_39372);
and U44922 (N_44922,N_37185,N_39357);
xor U44923 (N_44923,N_37677,N_39798);
and U44924 (N_44924,N_36000,N_35373);
xor U44925 (N_44925,N_38880,N_37417);
xor U44926 (N_44926,N_37307,N_37367);
nand U44927 (N_44927,N_35765,N_38588);
nand U44928 (N_44928,N_37225,N_36129);
nor U44929 (N_44929,N_38014,N_36104);
and U44930 (N_44930,N_36868,N_38340);
xnor U44931 (N_44931,N_38532,N_37696);
xor U44932 (N_44932,N_36017,N_36460);
nand U44933 (N_44933,N_35088,N_39856);
or U44934 (N_44934,N_39249,N_37431);
nand U44935 (N_44935,N_35042,N_35682);
nor U44936 (N_44936,N_35729,N_36975);
or U44937 (N_44937,N_38704,N_38529);
xnor U44938 (N_44938,N_39403,N_35983);
xor U44939 (N_44939,N_38937,N_38978);
xnor U44940 (N_44940,N_39264,N_36864);
nor U44941 (N_44941,N_38059,N_36737);
or U44942 (N_44942,N_39320,N_38977);
nor U44943 (N_44943,N_39541,N_38330);
nand U44944 (N_44944,N_38918,N_38769);
and U44945 (N_44945,N_35609,N_36257);
nor U44946 (N_44946,N_39834,N_39609);
and U44947 (N_44947,N_37216,N_39690);
xnor U44948 (N_44948,N_35452,N_38178);
or U44949 (N_44949,N_35519,N_35146);
nor U44950 (N_44950,N_37462,N_37275);
and U44951 (N_44951,N_35113,N_39065);
or U44952 (N_44952,N_39700,N_38065);
and U44953 (N_44953,N_36230,N_37316);
xnor U44954 (N_44954,N_36778,N_39339);
nor U44955 (N_44955,N_38381,N_37393);
nor U44956 (N_44956,N_38292,N_39809);
nand U44957 (N_44957,N_37440,N_36783);
nand U44958 (N_44958,N_38918,N_36116);
and U44959 (N_44959,N_38016,N_37924);
nand U44960 (N_44960,N_36002,N_39941);
or U44961 (N_44961,N_39416,N_39569);
and U44962 (N_44962,N_36347,N_39314);
or U44963 (N_44963,N_36831,N_35049);
and U44964 (N_44964,N_39322,N_36778);
nand U44965 (N_44965,N_38820,N_36387);
nor U44966 (N_44966,N_37109,N_35693);
or U44967 (N_44967,N_37611,N_38912);
xnor U44968 (N_44968,N_35784,N_35997);
nor U44969 (N_44969,N_37080,N_38792);
xor U44970 (N_44970,N_36141,N_39067);
or U44971 (N_44971,N_35643,N_38303);
nor U44972 (N_44972,N_38832,N_35089);
and U44973 (N_44973,N_35415,N_38220);
nor U44974 (N_44974,N_38472,N_37629);
nor U44975 (N_44975,N_36353,N_38868);
nand U44976 (N_44976,N_35448,N_38999);
nand U44977 (N_44977,N_38323,N_37432);
nor U44978 (N_44978,N_39167,N_38007);
nand U44979 (N_44979,N_39929,N_35322);
nand U44980 (N_44980,N_39763,N_36583);
xor U44981 (N_44981,N_35018,N_37293);
and U44982 (N_44982,N_36430,N_38229);
nand U44983 (N_44983,N_37994,N_36834);
or U44984 (N_44984,N_35237,N_36864);
nor U44985 (N_44985,N_36904,N_36581);
nand U44986 (N_44986,N_39696,N_36740);
xor U44987 (N_44987,N_38636,N_37991);
xor U44988 (N_44988,N_35249,N_36465);
or U44989 (N_44989,N_36409,N_37611);
nor U44990 (N_44990,N_38763,N_36398);
or U44991 (N_44991,N_36718,N_36239);
nand U44992 (N_44992,N_38528,N_36032);
nand U44993 (N_44993,N_35585,N_35935);
xnor U44994 (N_44994,N_37011,N_37808);
nand U44995 (N_44995,N_35152,N_39997);
or U44996 (N_44996,N_37293,N_38252);
xnor U44997 (N_44997,N_38219,N_37906);
xnor U44998 (N_44998,N_37312,N_37589);
nand U44999 (N_44999,N_35953,N_35230);
or U45000 (N_45000,N_41935,N_43130);
nor U45001 (N_45001,N_40688,N_44716);
nand U45002 (N_45002,N_42675,N_44620);
nor U45003 (N_45003,N_40921,N_43730);
xor U45004 (N_45004,N_40054,N_41054);
or U45005 (N_45005,N_42658,N_40948);
or U45006 (N_45006,N_44154,N_40458);
or U45007 (N_45007,N_41702,N_44452);
nand U45008 (N_45008,N_42041,N_42730);
and U45009 (N_45009,N_44350,N_40372);
nand U45010 (N_45010,N_42492,N_43751);
xor U45011 (N_45011,N_40530,N_40312);
nor U45012 (N_45012,N_42136,N_41226);
nor U45013 (N_45013,N_42363,N_44582);
or U45014 (N_45014,N_44299,N_44641);
nor U45015 (N_45015,N_44071,N_42765);
or U45016 (N_45016,N_44816,N_41997);
xnor U45017 (N_45017,N_40701,N_43807);
and U45018 (N_45018,N_41932,N_41814);
and U45019 (N_45019,N_43257,N_42021);
nand U45020 (N_45020,N_43221,N_42143);
xor U45021 (N_45021,N_44461,N_42903);
xnor U45022 (N_45022,N_41843,N_40851);
and U45023 (N_45023,N_40428,N_44510);
or U45024 (N_45024,N_43554,N_41560);
xor U45025 (N_45025,N_41206,N_40708);
or U45026 (N_45026,N_43036,N_44355);
or U45027 (N_45027,N_41175,N_40098);
nand U45028 (N_45028,N_40734,N_41886);
xnor U45029 (N_45029,N_43777,N_41679);
nor U45030 (N_45030,N_44965,N_41030);
nor U45031 (N_45031,N_44194,N_42076);
nand U45032 (N_45032,N_42277,N_42800);
nor U45033 (N_45033,N_41233,N_42617);
and U45034 (N_45034,N_43517,N_41671);
nor U45035 (N_45035,N_43499,N_41251);
nor U45036 (N_45036,N_42378,N_42390);
xnor U45037 (N_45037,N_41516,N_43229);
and U45038 (N_45038,N_44607,N_43564);
nor U45039 (N_45039,N_40060,N_42005);
or U45040 (N_45040,N_40581,N_43561);
nor U45041 (N_45041,N_42388,N_42811);
nand U45042 (N_45042,N_41334,N_42276);
nor U45043 (N_45043,N_42508,N_42635);
nand U45044 (N_45044,N_42497,N_42734);
or U45045 (N_45045,N_41165,N_44920);
or U45046 (N_45046,N_44183,N_40801);
or U45047 (N_45047,N_41195,N_42458);
nor U45048 (N_45048,N_43496,N_42840);
or U45049 (N_45049,N_42036,N_44746);
or U45050 (N_45050,N_43988,N_43833);
nand U45051 (N_45051,N_42343,N_41669);
xnor U45052 (N_45052,N_44516,N_44706);
and U45053 (N_45053,N_43811,N_41704);
nor U45054 (N_45054,N_41009,N_43659);
or U45055 (N_45055,N_44980,N_42769);
or U45056 (N_45056,N_42216,N_40025);
and U45057 (N_45057,N_40517,N_43260);
and U45058 (N_45058,N_44542,N_41210);
xnor U45059 (N_45059,N_44743,N_43521);
nor U45060 (N_45060,N_42274,N_41387);
or U45061 (N_45061,N_42038,N_42100);
xnor U45062 (N_45062,N_43658,N_41230);
or U45063 (N_45063,N_43198,N_42318);
nor U45064 (N_45064,N_40214,N_43228);
or U45065 (N_45065,N_41551,N_44683);
nand U45066 (N_45066,N_44229,N_40467);
nor U45067 (N_45067,N_43901,N_43971);
or U45068 (N_45068,N_41207,N_40176);
nand U45069 (N_45069,N_42472,N_42908);
xnor U45070 (N_45070,N_42962,N_41020);
xnor U45071 (N_45071,N_40862,N_40969);
or U45072 (N_45072,N_40356,N_43821);
and U45073 (N_45073,N_44069,N_40845);
nand U45074 (N_45074,N_44223,N_42651);
nor U45075 (N_45075,N_44755,N_43645);
nand U45076 (N_45076,N_42562,N_40953);
nor U45077 (N_45077,N_42251,N_43979);
or U45078 (N_45078,N_41014,N_42348);
nor U45079 (N_45079,N_41635,N_41940);
and U45080 (N_45080,N_40813,N_43592);
nor U45081 (N_45081,N_43143,N_41043);
or U45082 (N_45082,N_42961,N_41696);
nand U45083 (N_45083,N_44158,N_43154);
nand U45084 (N_45084,N_44102,N_42434);
xor U45085 (N_45085,N_44500,N_44916);
nand U45086 (N_45086,N_43794,N_42055);
nand U45087 (N_45087,N_43982,N_41055);
nor U45088 (N_45088,N_43851,N_42245);
nand U45089 (N_45089,N_40295,N_43675);
nor U45090 (N_45090,N_40123,N_41513);
xor U45091 (N_45091,N_42873,N_44244);
nor U45092 (N_45092,N_43177,N_40896);
or U45093 (N_45093,N_41307,N_42052);
xor U45094 (N_45094,N_43921,N_41095);
xnor U45095 (N_45095,N_40716,N_40571);
nor U45096 (N_45096,N_40736,N_42542);
or U45097 (N_45097,N_40313,N_41688);
or U45098 (N_45098,N_43339,N_44023);
and U45099 (N_45099,N_42965,N_43701);
nor U45100 (N_45100,N_40051,N_40446);
nor U45101 (N_45101,N_43719,N_41653);
and U45102 (N_45102,N_41885,N_43743);
nand U45103 (N_45103,N_40799,N_44002);
and U45104 (N_45104,N_42269,N_40362);
or U45105 (N_45105,N_43171,N_44742);
and U45106 (N_45106,N_40925,N_43184);
xnor U45107 (N_45107,N_41205,N_44204);
nand U45108 (N_45108,N_41336,N_43467);
nor U45109 (N_45109,N_40516,N_40271);
nor U45110 (N_45110,N_44935,N_40396);
nand U45111 (N_45111,N_40836,N_41778);
and U45112 (N_45112,N_41752,N_41735);
nand U45113 (N_45113,N_42056,N_44533);
nand U45114 (N_45114,N_44873,N_44674);
or U45115 (N_45115,N_41673,N_40321);
nand U45116 (N_45116,N_43938,N_41450);
nand U45117 (N_45117,N_42945,N_42547);
or U45118 (N_45118,N_43056,N_41874);
xnor U45119 (N_45119,N_40623,N_42719);
or U45120 (N_45120,N_44958,N_40785);
nor U45121 (N_45121,N_42892,N_43937);
nand U45122 (N_45122,N_41304,N_41581);
nor U45123 (N_45123,N_41798,N_43041);
and U45124 (N_45124,N_43981,N_42273);
or U45125 (N_45125,N_43599,N_42009);
nand U45126 (N_45126,N_42357,N_42128);
nor U45127 (N_45127,N_42196,N_42422);
nor U45128 (N_45128,N_42219,N_43071);
or U45129 (N_45129,N_42202,N_41291);
nor U45130 (N_45130,N_42442,N_43200);
and U45131 (N_45131,N_42834,N_44015);
and U45132 (N_45132,N_42333,N_40773);
nor U45133 (N_45133,N_40478,N_44250);
or U45134 (N_45134,N_42950,N_42159);
nor U45135 (N_45135,N_44235,N_41637);
or U45136 (N_45136,N_43435,N_41512);
nand U45137 (N_45137,N_41375,N_42450);
nand U45138 (N_45138,N_44831,N_44814);
and U45139 (N_45139,N_40498,N_42370);
xor U45140 (N_45140,N_44687,N_40594);
or U45141 (N_45141,N_40565,N_44179);
or U45142 (N_45142,N_43123,N_44526);
or U45143 (N_45143,N_40730,N_41829);
nand U45144 (N_45144,N_43250,N_44891);
nor U45145 (N_45145,N_41571,N_44342);
nand U45146 (N_45146,N_44583,N_41625);
or U45147 (N_45147,N_44029,N_40911);
nor U45148 (N_45148,N_41302,N_44850);
xnor U45149 (N_45149,N_44281,N_43356);
nand U45150 (N_45150,N_42307,N_42500);
nor U45151 (N_45151,N_44415,N_40535);
and U45152 (N_45152,N_43300,N_41572);
xor U45153 (N_45153,N_44495,N_42411);
and U45154 (N_45154,N_42167,N_42369);
nand U45155 (N_45155,N_41805,N_43026);
or U45156 (N_45156,N_41996,N_42032);
nor U45157 (N_45157,N_43654,N_43954);
or U45158 (N_45158,N_40908,N_44326);
and U45159 (N_45159,N_44626,N_40978);
xnor U45160 (N_45160,N_42035,N_43651);
or U45161 (N_45161,N_43740,N_44453);
nor U45162 (N_45162,N_44243,N_40027);
nor U45163 (N_45163,N_40946,N_43600);
nand U45164 (N_45164,N_43519,N_43380);
xor U45165 (N_45165,N_44210,N_44983);
xor U45166 (N_45166,N_42392,N_44982);
nand U45167 (N_45167,N_41909,N_40551);
or U45168 (N_45168,N_42376,N_43135);
nand U45169 (N_45169,N_43082,N_40547);
nand U45170 (N_45170,N_42365,N_40979);
xnor U45171 (N_45171,N_40369,N_40602);
or U45172 (N_45172,N_44203,N_44829);
xor U45173 (N_45173,N_42158,N_42573);
or U45174 (N_45174,N_41786,N_40455);
nor U45175 (N_45175,N_42499,N_40126);
or U45176 (N_45176,N_40032,N_42090);
nor U45177 (N_45177,N_44178,N_43692);
nand U45178 (N_45178,N_43349,N_43239);
nand U45179 (N_45179,N_43681,N_44788);
nor U45180 (N_45180,N_44538,N_41577);
nand U45181 (N_45181,N_41739,N_42859);
or U45182 (N_45182,N_42067,N_40501);
and U45183 (N_45183,N_42698,N_44307);
or U45184 (N_45184,N_44662,N_40273);
nor U45185 (N_45185,N_44792,N_40844);
nor U45186 (N_45186,N_44425,N_44368);
or U45187 (N_45187,N_41860,N_44142);
nor U45188 (N_45188,N_43949,N_44637);
xnor U45189 (N_45189,N_43573,N_41189);
and U45190 (N_45190,N_44185,N_40666);
nand U45191 (N_45191,N_44314,N_43422);
xnor U45192 (N_45192,N_41119,N_42105);
nand U45193 (N_45193,N_41140,N_44907);
and U45194 (N_45194,N_41758,N_41089);
and U45195 (N_45195,N_40834,N_43855);
and U45196 (N_45196,N_44460,N_44991);
and U45197 (N_45197,N_42642,N_43650);
and U45198 (N_45198,N_40597,N_44233);
or U45199 (N_45199,N_40213,N_44752);
xnor U45200 (N_45200,N_40926,N_43662);
xnor U45201 (N_45201,N_42132,N_44031);
nand U45202 (N_45202,N_41204,N_44602);
nand U45203 (N_45203,N_43014,N_40221);
xnor U45204 (N_45204,N_43428,N_40513);
xnor U45205 (N_45205,N_44430,N_41453);
and U45206 (N_45206,N_43567,N_42759);
or U45207 (N_45207,N_40608,N_40936);
nand U45208 (N_45208,N_43503,N_42728);
xnor U45209 (N_45209,N_40584,N_43501);
nand U45210 (N_45210,N_40725,N_44987);
nand U45211 (N_45211,N_42043,N_40550);
and U45212 (N_45212,N_41836,N_43776);
nor U45213 (N_45213,N_42410,N_42352);
nand U45214 (N_45214,N_44310,N_43414);
xor U45215 (N_45215,N_40359,N_40249);
or U45216 (N_45216,N_44232,N_44875);
and U45217 (N_45217,N_42987,N_42096);
nand U45218 (N_45218,N_42576,N_44170);
and U45219 (N_45219,N_42327,N_44475);
and U45220 (N_45220,N_44544,N_44159);
xor U45221 (N_45221,N_40185,N_43731);
or U45222 (N_45222,N_43125,N_44643);
nor U45223 (N_45223,N_44758,N_42594);
and U45224 (N_45224,N_44981,N_41213);
nor U45225 (N_45225,N_43138,N_43936);
or U45226 (N_45226,N_40409,N_44024);
or U45227 (N_45227,N_43323,N_43585);
or U45228 (N_45228,N_40568,N_41167);
and U45229 (N_45229,N_41761,N_41182);
nand U45230 (N_45230,N_42874,N_41612);
or U45231 (N_45231,N_41993,N_43310);
or U45232 (N_45232,N_43950,N_42663);
xor U45233 (N_45233,N_41595,N_40100);
xnor U45234 (N_45234,N_43879,N_41854);
and U45235 (N_45235,N_43488,N_40430);
xor U45236 (N_45236,N_42853,N_41051);
xor U45237 (N_45237,N_44364,N_43589);
nand U45238 (N_45238,N_43736,N_42204);
nor U45239 (N_45239,N_43185,N_42498);
nor U45240 (N_45240,N_44843,N_43845);
nand U45241 (N_45241,N_44613,N_44195);
and U45242 (N_45242,N_40089,N_44611);
or U45243 (N_45243,N_42195,N_44714);
or U45244 (N_45244,N_44008,N_44554);
xor U45245 (N_45245,N_44793,N_40385);
nand U45246 (N_45246,N_40552,N_42176);
and U45247 (N_45247,N_40744,N_41824);
and U45248 (N_45248,N_44269,N_41289);
and U45249 (N_45249,N_44412,N_42374);
or U45250 (N_45250,N_44764,N_44512);
and U45251 (N_45251,N_43984,N_41025);
nand U45252 (N_45252,N_42290,N_43986);
or U45253 (N_45253,N_44937,N_44664);
nand U45254 (N_45254,N_41142,N_40915);
and U45255 (N_45255,N_41478,N_41105);
xnor U45256 (N_45256,N_42944,N_42194);
or U45257 (N_45257,N_43848,N_43825);
nor U45258 (N_45258,N_44035,N_41700);
or U45259 (N_45259,N_42483,N_43305);
and U45260 (N_45260,N_43085,N_41587);
xnor U45261 (N_45261,N_41217,N_42708);
or U45262 (N_45262,N_44395,N_43684);
nor U45263 (N_45263,N_40819,N_44367);
xnor U45264 (N_45264,N_42943,N_44389);
or U45265 (N_45265,N_44869,N_40743);
and U45266 (N_45266,N_41744,N_42014);
nor U45267 (N_45267,N_44592,N_44696);
nor U45268 (N_45268,N_42402,N_42074);
xnor U45269 (N_45269,N_44379,N_44330);
xor U45270 (N_45270,N_40417,N_42782);
nor U45271 (N_45271,N_42806,N_44836);
or U45272 (N_45272,N_43044,N_43612);
and U45273 (N_45273,N_41792,N_41769);
or U45274 (N_45274,N_40558,N_42791);
and U45275 (N_45275,N_43957,N_44635);
or U45276 (N_45276,N_40986,N_40152);
nor U45277 (N_45277,N_40404,N_43399);
nor U45278 (N_45278,N_41593,N_40425);
and U45279 (N_45279,N_41227,N_40999);
nor U45280 (N_45280,N_41393,N_40325);
nand U45281 (N_45281,N_41951,N_40363);
and U45282 (N_45282,N_44969,N_41785);
and U45283 (N_45283,N_40657,N_42662);
nor U45284 (N_45284,N_44551,N_40745);
and U45285 (N_45285,N_40655,N_40869);
nor U45286 (N_45286,N_40504,N_44865);
and U45287 (N_45287,N_44226,N_42565);
and U45288 (N_45288,N_41211,N_44870);
xnor U45289 (N_45289,N_42579,N_43121);
nor U45290 (N_45290,N_40483,N_43906);
nor U45291 (N_45291,N_43073,N_43856);
and U45292 (N_45292,N_40172,N_44098);
nor U45293 (N_45293,N_44694,N_43314);
nand U45294 (N_45294,N_43023,N_44313);
nand U45295 (N_45295,N_41665,N_41208);
or U45296 (N_45296,N_41479,N_40416);
or U45297 (N_45297,N_43758,N_41942);
xor U45298 (N_45298,N_43420,N_40639);
xor U45299 (N_45299,N_43820,N_40237);
nand U45300 (N_45300,N_40858,N_44278);
xor U45301 (N_45301,N_43775,N_43116);
nand U45302 (N_45302,N_41172,N_40143);
nand U45303 (N_45303,N_41121,N_44832);
nor U45304 (N_45304,N_41346,N_44537);
nand U45305 (N_45305,N_44082,N_43141);
xnor U45306 (N_45306,N_44862,N_43598);
or U45307 (N_45307,N_40320,N_43463);
or U45308 (N_45308,N_42625,N_44563);
or U45309 (N_45309,N_43273,N_42033);
and U45310 (N_45310,N_42780,N_41876);
xnor U45311 (N_45311,N_43887,N_43985);
nor U45312 (N_45312,N_40304,N_44092);
nand U45313 (N_45313,N_40793,N_44219);
xor U45314 (N_45314,N_44847,N_43225);
xor U45315 (N_45315,N_43169,N_41071);
xor U45316 (N_45316,N_42353,N_41098);
or U45317 (N_45317,N_43159,N_44901);
xor U45318 (N_45318,N_43858,N_43369);
nor U45319 (N_45319,N_44550,N_40491);
nand U45320 (N_45320,N_44316,N_44036);
nand U45321 (N_45321,N_42350,N_43261);
xnor U45322 (N_45322,N_40660,N_44094);
nand U45323 (N_45323,N_43477,N_43993);
nand U45324 (N_45324,N_40528,N_43571);
or U45325 (N_45325,N_41008,N_43557);
nand U45326 (N_45326,N_42454,N_40252);
nand U45327 (N_45327,N_41952,N_40088);
nand U45328 (N_45328,N_42308,N_43417);
and U45329 (N_45329,N_40019,N_40916);
and U45330 (N_45330,N_43570,N_42334);
nand U45331 (N_45331,N_43699,N_41272);
nor U45332 (N_45332,N_43466,N_44954);
and U45333 (N_45333,N_43452,N_43952);
or U45334 (N_45334,N_42201,N_41856);
nand U45335 (N_45335,N_44397,N_43223);
xor U45336 (N_45336,N_42699,N_42137);
and U45337 (N_45337,N_42300,N_43508);
and U45338 (N_45338,N_44892,N_41762);
nand U45339 (N_45339,N_42464,N_42119);
or U45340 (N_45340,N_41928,N_41736);
xor U45341 (N_45341,N_43388,N_40894);
or U45342 (N_45342,N_40265,N_44441);
and U45343 (N_45343,N_43375,N_40135);
or U45344 (N_45344,N_43390,N_44328);
or U45345 (N_45345,N_43386,N_40183);
and U45346 (N_45346,N_40975,N_41549);
xor U45347 (N_45347,N_44797,N_42440);
nand U45348 (N_45348,N_41701,N_41046);
and U45349 (N_45349,N_41955,N_41707);
xor U45350 (N_45350,N_41490,N_41618);
or U45351 (N_45351,N_41040,N_42200);
nand U45352 (N_45352,N_42424,N_42523);
nor U45353 (N_45353,N_44349,N_40354);
and U45354 (N_45354,N_43810,N_41435);
and U45355 (N_45355,N_40515,N_40593);
or U45356 (N_45356,N_42895,N_42910);
nor U45357 (N_45357,N_40297,N_40180);
xor U45358 (N_45358,N_43733,N_40073);
or U45359 (N_45359,N_40493,N_40559);
nor U45360 (N_45360,N_42248,N_43511);
nor U45361 (N_45361,N_43755,N_42823);
nand U45362 (N_45362,N_43972,N_44467);
nor U45363 (N_45363,N_42799,N_40949);
and U45364 (N_45364,N_43498,N_43366);
and U45365 (N_45365,N_41371,N_40873);
or U45366 (N_45366,N_41573,N_40033);
xnor U45367 (N_45367,N_43707,N_44523);
nand U45368 (N_45368,N_41883,N_42437);
nor U45369 (N_45369,N_40792,N_42963);
and U45370 (N_45370,N_42985,N_40284);
nor U45371 (N_45371,N_41884,N_42827);
and U45372 (N_45372,N_41062,N_44234);
nor U45373 (N_45373,N_40360,N_43661);
and U45374 (N_45374,N_41525,N_43092);
and U45375 (N_45375,N_43129,N_42608);
and U45376 (N_45376,N_44091,N_44568);
nor U45377 (N_45377,N_41579,N_42710);
nor U45378 (N_45378,N_44414,N_40110);
or U45379 (N_45379,N_42537,N_43107);
xor U45380 (N_45380,N_44302,N_43964);
or U45381 (N_45381,N_41651,N_44319);
or U45382 (N_45382,N_40216,N_42757);
and U45383 (N_45383,N_42380,N_40093);
nand U45384 (N_45384,N_44841,N_43621);
nand U45385 (N_45385,N_42724,N_43882);
xnor U45386 (N_45386,N_42727,N_40720);
and U45387 (N_45387,N_44534,N_41488);
nand U45388 (N_45388,N_42400,N_43437);
nor U45389 (N_45389,N_44573,N_42828);
xor U45390 (N_45390,N_40058,N_41599);
nor U45391 (N_45391,N_40775,N_44005);
nand U45392 (N_45392,N_44486,N_44188);
nand U45393 (N_45393,N_40454,N_41541);
nor U45394 (N_45394,N_41862,N_44724);
and U45395 (N_45395,N_44013,N_43543);
xor U45396 (N_45396,N_44236,N_43847);
or U45397 (N_45397,N_41586,N_42170);
or U45398 (N_45398,N_40103,N_41646);
nor U45399 (N_45399,N_42741,N_44051);
and U45400 (N_45400,N_40595,N_42126);
xor U45401 (N_45401,N_40543,N_40804);
nand U45402 (N_45402,N_43226,N_41292);
nand U45403 (N_45403,N_44259,N_42817);
or U45404 (N_45404,N_44025,N_41399);
and U45405 (N_45405,N_42496,N_41898);
nand U45406 (N_45406,N_43162,N_43943);
nand U45407 (N_45407,N_40957,N_42210);
nor U45408 (N_45408,N_42198,N_44206);
nand U45409 (N_45409,N_44921,N_43165);
or U45410 (N_45410,N_44168,N_40330);
xor U45411 (N_45411,N_43320,N_40275);
nor U45412 (N_45412,N_40236,N_42085);
nor U45413 (N_45413,N_42818,N_42815);
or U45414 (N_45414,N_43105,N_42923);
or U45415 (N_45415,N_43577,N_40193);
nor U45416 (N_45416,N_44230,N_43338);
and U45417 (N_45417,N_40939,N_41921);
xnor U45418 (N_45418,N_43240,N_44738);
xor U45419 (N_45419,N_43786,N_41104);
xnor U45420 (N_45420,N_41415,N_41994);
xor U45421 (N_45421,N_42089,N_42669);
or U45422 (N_45422,N_44353,N_42439);
and U45423 (N_45423,N_44298,N_40053);
and U45424 (N_45424,N_42181,N_42484);
and U45425 (N_45425,N_42125,N_41806);
xor U45426 (N_45426,N_42025,N_44134);
or U45427 (N_45427,N_40930,N_44042);
xnor U45428 (N_45428,N_42495,N_42849);
and U45429 (N_45429,N_43487,N_44491);
and U45430 (N_45430,N_40596,N_40147);
xor U45431 (N_45431,N_44589,N_43728);
xor U45432 (N_45432,N_44945,N_44595);
and U45433 (N_45433,N_43854,N_42754);
nand U45434 (N_45434,N_40310,N_40879);
nor U45435 (N_45435,N_41042,N_43181);
or U45436 (N_45436,N_43020,N_44936);
or U45437 (N_45437,N_41750,N_41088);
and U45438 (N_45438,N_40522,N_40373);
and U45439 (N_45439,N_42763,N_41097);
and U45440 (N_45440,N_43447,N_44050);
and U45441 (N_45441,N_43371,N_41832);
or U45442 (N_45442,N_41357,N_40452);
xor U45443 (N_45443,N_42104,N_40769);
xnor U45444 (N_45444,N_42024,N_43419);
nand U45445 (N_45445,N_44772,N_42952);
or U45446 (N_45446,N_41911,N_41622);
and U45447 (N_45447,N_41539,N_43611);
or U45448 (N_45448,N_41457,N_44262);
nor U45449 (N_45449,N_40825,N_40561);
nor U45450 (N_45450,N_43899,N_41929);
nor U45451 (N_45451,N_41144,N_41675);
and U45452 (N_45452,N_41661,N_40765);
nand U45453 (N_45453,N_40514,N_44133);
or U45454 (N_45454,N_41392,N_40675);
xor U45455 (N_45455,N_43760,N_41420);
nand U45456 (N_45456,N_41975,N_42093);
and U45457 (N_45457,N_44681,N_43485);
nand U45458 (N_45458,N_40338,N_44290);
and U45459 (N_45459,N_44968,N_43966);
xor U45460 (N_45460,N_42525,N_40820);
xor U45461 (N_45461,N_41831,N_40508);
nand U45462 (N_45462,N_41363,N_44143);
xor U45463 (N_45463,N_40636,N_44722);
xor U45464 (N_45464,N_42505,N_44735);
nor U45465 (N_45465,N_44539,N_43762);
nand U45466 (N_45466,N_40267,N_43110);
or U45467 (N_45467,N_41359,N_42094);
nand U45468 (N_45468,N_40258,N_40263);
xnor U45469 (N_45469,N_43407,N_43377);
or U45470 (N_45470,N_40826,N_41995);
nand U45471 (N_45471,N_44868,N_43316);
nand U45472 (N_45472,N_42742,N_43358);
xnor U45473 (N_45473,N_44341,N_40062);
xnor U45474 (N_45474,N_42890,N_40523);
nand U45475 (N_45475,N_41096,N_40342);
or U45476 (N_45476,N_43510,N_44088);
nor U45477 (N_45477,N_41428,N_44360);
and U45478 (N_45478,N_43559,N_42426);
and U45479 (N_45479,N_42417,N_42443);
or U45480 (N_45480,N_40621,N_41076);
nand U45481 (N_45481,N_44402,N_42623);
nor U45482 (N_45482,N_44605,N_40182);
or U45483 (N_45483,N_42364,N_41601);
xnor U45484 (N_45484,N_42648,N_41328);
nand U45485 (N_45485,N_43333,N_44241);
and U45486 (N_45486,N_44707,N_44727);
xnor U45487 (N_45487,N_41780,N_40272);
nor U45488 (N_45488,N_41880,N_44803);
and U45489 (N_45489,N_40861,N_41753);
and U45490 (N_45490,N_40337,N_40822);
nor U45491 (N_45491,N_40470,N_40629);
nand U45492 (N_45492,N_41694,N_41250);
nor U45493 (N_45493,N_43902,N_40931);
nand U45494 (N_45494,N_43471,N_42467);
and U45495 (N_45495,N_43078,N_43195);
nand U45496 (N_45496,N_42820,N_40790);
or U45497 (N_45497,N_41575,N_42556);
xor U45498 (N_45498,N_41748,N_44795);
nand U45499 (N_45499,N_41636,N_41633);
nor U45500 (N_45500,N_41544,N_42079);
nor U45501 (N_45501,N_40131,N_43969);
and U45502 (N_45502,N_40780,N_42491);
nor U45503 (N_45503,N_44576,N_40546);
nor U45504 (N_45504,N_42755,N_44636);
xnor U45505 (N_45505,N_40071,N_40802);
nand U45506 (N_45506,N_44628,N_41664);
xor U45507 (N_45507,N_41396,N_43441);
nand U45508 (N_45508,N_40566,N_40013);
nand U45509 (N_45509,N_41000,N_41828);
or U45510 (N_45510,N_42826,N_44910);
xnor U45511 (N_45511,N_41582,N_44939);
xor U45512 (N_45512,N_40282,N_41436);
nor U45513 (N_45513,N_42331,N_40302);
xnor U45514 (N_45514,N_42580,N_43977);
and U45515 (N_45515,N_40798,N_44854);
nor U45516 (N_45516,N_41235,N_42445);
xnor U45517 (N_45517,N_42435,N_41990);
nor U45518 (N_45518,N_44303,N_44767);
nor U45519 (N_45519,N_44952,N_40431);
and U45520 (N_45520,N_42722,N_43489);
nand U45521 (N_45521,N_40411,N_44199);
nor U45522 (N_45522,N_43066,N_41959);
or U45523 (N_45523,N_42684,N_43624);
nor U45524 (N_45524,N_42156,N_43513);
and U45525 (N_45525,N_43623,N_40256);
nand U45526 (N_45526,N_43394,N_40889);
xor U45527 (N_45527,N_41214,N_43756);
nor U45528 (N_45528,N_43789,N_44334);
nand U45529 (N_45529,N_43846,N_41520);
xnor U45530 (N_45530,N_42151,N_41446);
xor U45531 (N_45531,N_44496,N_43294);
xor U45532 (N_45532,N_43667,N_40917);
and U45533 (N_45533,N_40192,N_41710);
xor U45534 (N_45534,N_42877,N_41306);
and U45535 (N_45535,N_41944,N_44697);
and U45536 (N_45536,N_41706,N_44749);
nand U45537 (N_45537,N_43885,N_43389);
and U45538 (N_45538,N_42661,N_41181);
nand U45539 (N_45539,N_40965,N_41931);
xor U45540 (N_45540,N_42524,N_42012);
nor U45541 (N_45541,N_42612,N_44630);
or U45542 (N_45542,N_42183,N_42184);
nand U45543 (N_45543,N_40173,N_40057);
nand U45544 (N_45544,N_40296,N_43607);
nor U45545 (N_45545,N_44080,N_43630);
and U45546 (N_45546,N_42883,N_42106);
nand U45547 (N_45547,N_41894,N_41329);
or U45548 (N_45548,N_40408,N_44086);
nor U45549 (N_45549,N_43830,N_42456);
nor U45550 (N_45550,N_40164,N_41811);
xor U45551 (N_45551,N_44712,N_40778);
or U45552 (N_45552,N_43739,N_41261);
or U45553 (N_45553,N_42027,N_40784);
and U45554 (N_45554,N_43889,N_44273);
and U45555 (N_45555,N_40007,N_43581);
xnor U45556 (N_45556,N_43759,N_40770);
and U45557 (N_45557,N_42848,N_41099);
nand U45558 (N_45558,N_44480,N_42477);
and U45559 (N_45559,N_44710,N_42960);
nor U45560 (N_45560,N_40381,N_42061);
and U45561 (N_45561,N_44137,N_44161);
nand U45562 (N_45562,N_41402,N_40717);
nand U45563 (N_45563,N_40521,N_42432);
or U45564 (N_45564,N_44530,N_43941);
nand U45565 (N_45565,N_41864,N_43266);
nand U45566 (N_45566,N_42165,N_43364);
xnor U45567 (N_45567,N_44631,N_43063);
xor U45568 (N_45568,N_43813,N_40210);
and U45569 (N_45569,N_40968,N_41906);
nand U45570 (N_45570,N_41655,N_40043);
or U45571 (N_45571,N_42783,N_43426);
nor U45572 (N_45572,N_41045,N_43872);
nand U45573 (N_45573,N_41937,N_43047);
nor U45574 (N_45574,N_43955,N_41029);
nand U45575 (N_45575,N_42372,N_40161);
xor U45576 (N_45576,N_41789,N_40850);
xnor U45577 (N_45577,N_42825,N_42482);
nand U45578 (N_45578,N_40641,N_41125);
and U45579 (N_45579,N_40293,N_41965);
and U45580 (N_45580,N_41791,N_43208);
nor U45581 (N_45581,N_40171,N_42681);
and U45582 (N_45582,N_41281,N_44196);
nor U45583 (N_45583,N_41794,N_43318);
or U45584 (N_45584,N_43241,N_42218);
and U45585 (N_45585,N_43686,N_43244);
nor U45586 (N_45586,N_41841,N_41687);
or U45587 (N_45587,N_42639,N_42260);
and U45588 (N_45588,N_44352,N_40349);
nand U45589 (N_45589,N_42286,N_43823);
nand U45590 (N_45590,N_44409,N_40626);
nor U45591 (N_45591,N_43771,N_42063);
nor U45592 (N_45592,N_43814,N_40964);
or U45593 (N_45593,N_41135,N_43395);
and U45594 (N_45594,N_43412,N_40423);
nor U45595 (N_45595,N_43303,N_41763);
or U45596 (N_45596,N_44129,N_41743);
nor U45597 (N_45597,N_41145,N_43252);
or U45598 (N_45598,N_43072,N_41440);
nand U45599 (N_45599,N_43657,N_43413);
xor U45600 (N_45600,N_42948,N_43163);
nand U45601 (N_45601,N_43343,N_43022);
and U45602 (N_45602,N_41903,N_43824);
xnor U45603 (N_45603,N_40881,N_41659);
xor U45604 (N_45604,N_42855,N_40632);
and U45605 (N_45605,N_44215,N_44345);
xnor U45606 (N_45606,N_43627,N_41493);
nor U45607 (N_45607,N_43212,N_44986);
nand U45608 (N_45608,N_43722,N_42473);
nand U45609 (N_45609,N_43282,N_41215);
nand U45610 (N_45610,N_44371,N_42678);
nand U45611 (N_45611,N_44603,N_44827);
nor U45612 (N_45612,N_41968,N_40562);
and U45613 (N_45613,N_40913,N_44872);
nor U45614 (N_45614,N_44659,N_44114);
xnor U45615 (N_45615,N_44704,N_44717);
xnor U45616 (N_45616,N_42522,N_44165);
nor U45617 (N_45617,N_40622,N_44315);
nand U45618 (N_45618,N_41245,N_44173);
nand U45619 (N_45619,N_41893,N_40482);
and U45620 (N_45620,N_41683,N_44541);
nor U45621 (N_45621,N_41362,N_42550);
xnor U45622 (N_45622,N_42753,N_43500);
nand U45623 (N_45623,N_43669,N_40886);
xnor U45624 (N_45624,N_41550,N_44721);
nand U45625 (N_45625,N_40752,N_42809);
and U45626 (N_45626,N_42084,N_43174);
nor U45627 (N_45627,N_42384,N_44505);
xnor U45628 (N_45628,N_40899,N_43490);
and U45629 (N_45629,N_43724,N_43263);
or U45630 (N_45630,N_44619,N_41823);
nor U45631 (N_45631,N_44009,N_44494);
nand U45632 (N_45632,N_42835,N_42141);
nor U45633 (N_45633,N_43462,N_43748);
xnor U45634 (N_45634,N_41534,N_44699);
xor U45635 (N_45635,N_44923,N_41383);
or U45636 (N_45636,N_44388,N_43469);
and U45637 (N_45637,N_41374,N_41641);
xnor U45638 (N_45638,N_44656,N_44182);
and U45639 (N_45639,N_44692,N_40351);
nor U45640 (N_45640,N_43695,N_44740);
and U45641 (N_45641,N_44107,N_42515);
xor U45642 (N_45642,N_44846,N_41150);
and U45643 (N_45643,N_42743,N_44141);
nor U45644 (N_45644,N_42004,N_43553);
and U45645 (N_45645,N_42714,N_41048);
nand U45646 (N_45646,N_40394,N_42224);
and U45647 (N_45647,N_41391,N_42302);
nand U45648 (N_45648,N_43342,N_43815);
and U45649 (N_45649,N_41159,N_43336);
xnor U45650 (N_45650,N_40091,N_41180);
nor U45651 (N_45651,N_41455,N_44900);
xnor U45652 (N_45652,N_42601,N_42017);
nor U45653 (N_45653,N_40668,N_40395);
xnor U45654 (N_45654,N_43502,N_43363);
nor U45655 (N_45655,N_44566,N_44004);
xor U45656 (N_45656,N_44190,N_40995);
xor U45657 (N_45657,N_42843,N_42915);
nand U45658 (N_45658,N_43296,N_40120);
nand U45659 (N_45659,N_42660,N_43634);
or U45660 (N_45660,N_40205,N_40086);
xnor U45661 (N_45661,N_41416,N_43655);
xor U45662 (N_45662,N_43151,N_41279);
nor U45663 (N_45663,N_40564,N_41768);
or U45664 (N_45664,N_41709,N_44301);
nand U45665 (N_45665,N_42620,N_41034);
nor U45666 (N_45666,N_40787,N_40653);
and U45667 (N_45667,N_41692,N_40727);
nand U45668 (N_45668,N_43905,N_40524);
xor U45669 (N_45669,N_42455,N_44919);
or U45670 (N_45670,N_43232,N_42589);
nor U45671 (N_45671,N_40162,N_42254);
xor U45672 (N_45672,N_42964,N_44416);
and U45673 (N_45673,N_40006,N_43738);
xor U45674 (N_45674,N_41366,N_42053);
nand U45675 (N_45675,N_42653,N_40614);
nor U45676 (N_45676,N_42549,N_41007);
and U45677 (N_45677,N_43700,N_44560);
nand U45678 (N_45678,N_44623,N_41857);
xor U45679 (N_45679,N_42711,N_44120);
xnor U45680 (N_45680,N_44556,N_42957);
xnor U45681 (N_45681,N_44956,N_43486);
xnor U45682 (N_45682,N_42163,N_43840);
or U45683 (N_45683,N_41989,N_42229);
nand U45684 (N_45684,N_43242,N_40156);
xnor U45685 (N_45685,N_43796,N_40365);
or U45686 (N_45686,N_44074,N_40040);
nor U45687 (N_45687,N_41360,N_41764);
or U45688 (N_45688,N_41578,N_44208);
nor U45689 (N_45689,N_41984,N_42112);
nor U45690 (N_45690,N_40364,N_41093);
nor U45691 (N_45691,N_41576,N_44715);
nor U45692 (N_45692,N_44796,N_42805);
xnor U45693 (N_45693,N_43281,N_40034);
nor U45694 (N_45694,N_42936,N_40031);
and U45695 (N_45695,N_42355,N_41855);
and U45696 (N_45696,N_44027,N_41741);
or U45697 (N_45697,N_43913,N_40989);
nand U45698 (N_45698,N_43387,N_43891);
xor U45699 (N_45699,N_44588,N_44076);
nand U45700 (N_45700,N_40980,N_44736);
nor U45701 (N_45701,N_42314,N_41776);
and U45702 (N_45702,N_43322,N_43808);
nand U45703 (N_45703,N_44765,N_44852);
and U45704 (N_45704,N_43011,N_41722);
xnor U45705 (N_45705,N_43480,N_40035);
and U45706 (N_45706,N_44468,N_43525);
xnor U45707 (N_45707,N_40096,N_43103);
xor U45708 (N_45708,N_43334,N_42989);
or U45709 (N_45709,N_43613,N_41718);
or U45710 (N_45710,N_41154,N_42829);
nor U45711 (N_45711,N_41426,N_43983);
or U45712 (N_45712,N_44131,N_43919);
xor U45713 (N_45713,N_43246,N_40499);
nor U45714 (N_45714,N_41102,N_43908);
and U45715 (N_45715,N_44451,N_40791);
nand U45716 (N_45716,N_44449,N_40697);
or U45717 (N_45717,N_40811,N_41069);
xor U45718 (N_45718,N_40305,N_41265);
nand U45719 (N_45719,N_44929,N_44897);
or U45720 (N_45720,N_43933,N_42544);
or U45721 (N_45721,N_43584,N_41032);
nand U45722 (N_45722,N_40011,N_41826);
or U45723 (N_45723,N_44511,N_41680);
nand U45724 (N_45724,N_41187,N_41114);
xnor U45725 (N_45725,N_40574,N_42263);
and U45726 (N_45726,N_43397,N_44904);
nor U45727 (N_45727,N_41255,N_40474);
and U45728 (N_45728,N_42264,N_43290);
nor U45729 (N_45729,N_43867,N_42108);
and U45730 (N_45730,N_41219,N_41406);
and U45731 (N_45731,N_41452,N_41535);
nand U45732 (N_45732,N_43046,N_41358);
nand U45733 (N_45733,N_41244,N_40082);
nor U45734 (N_45734,N_43631,N_43190);
nand U45735 (N_45735,N_40656,N_40842);
xnor U45736 (N_45736,N_41130,N_41058);
nor U45737 (N_45737,N_43404,N_43852);
xor U45738 (N_45738,N_44055,N_40805);
xnor U45739 (N_45739,N_40977,N_42250);
nand U45740 (N_45740,N_40492,N_44113);
nor U45741 (N_45741,N_44401,N_41492);
nor U45742 (N_45742,N_42468,N_44709);
xor U45743 (N_45743,N_40669,N_41026);
or U45744 (N_45744,N_42396,N_44493);
and U45745 (N_45745,N_44679,N_42969);
xnor U45746 (N_45746,N_42771,N_41199);
or U45747 (N_45747,N_42320,N_42377);
and U45748 (N_45748,N_42846,N_42168);
or U45749 (N_45749,N_44934,N_40000);
or U45750 (N_45750,N_42404,N_44543);
or U45751 (N_45751,N_42740,N_41355);
and U45752 (N_45752,N_40510,N_43126);
nand U45753 (N_45753,N_44172,N_43528);
or U45754 (N_45754,N_42836,N_43685);
nor U45755 (N_45755,N_41247,N_44810);
nand U45756 (N_45756,N_42744,N_41538);
nand U45757 (N_45757,N_41946,N_43024);
xor U45758 (N_45758,N_40068,N_42569);
or U45759 (N_45759,N_41608,N_42186);
nor U45760 (N_45760,N_40418,N_42955);
nand U45761 (N_45761,N_40796,N_40649);
nand U45762 (N_45762,N_41902,N_44443);
and U45763 (N_45763,N_44590,N_41129);
nor U45764 (N_45764,N_41938,N_44485);
nand U45765 (N_45765,N_43583,N_40700);
xor U45766 (N_45766,N_42670,N_40971);
and U45767 (N_45767,N_43626,N_44633);
and U45768 (N_45768,N_41605,N_40829);
or U45769 (N_45769,N_44338,N_44213);
and U45770 (N_45770,N_44472,N_44487);
nand U45771 (N_45771,N_43182,N_41727);
or U45772 (N_45772,N_40081,N_44524);
nor U45773 (N_45773,N_40827,N_43052);
or U45774 (N_45774,N_44046,N_40625);
nor U45775 (N_45775,N_40997,N_43051);
or U45776 (N_45776,N_43315,N_42275);
and U45777 (N_45777,N_43507,N_43313);
nor U45778 (N_45778,N_41693,N_41717);
nor U45779 (N_45779,N_44366,N_41297);
and U45780 (N_45780,N_42344,N_40662);
and U45781 (N_45781,N_43666,N_42080);
nor U45782 (N_45782,N_40115,N_43838);
xor U45783 (N_45783,N_41755,N_44162);
or U45784 (N_45784,N_44757,N_42029);
or U45785 (N_45785,N_44205,N_40026);
nand U45786 (N_45786,N_42566,N_40419);
and U45787 (N_45787,N_40613,N_40270);
nand U45788 (N_45788,N_44799,N_43091);
xor U45789 (N_45789,N_42382,N_40627);
nor U45790 (N_45790,N_44476,N_41985);
nor U45791 (N_45791,N_42921,N_40664);
or U45792 (N_45792,N_41319,N_42593);
nor U45793 (N_45793,N_41731,N_42602);
or U45794 (N_45794,N_40534,N_44197);
nand U45795 (N_45795,N_42626,N_40719);
nand U45796 (N_45796,N_41332,N_40463);
nor U45797 (N_45797,N_43094,N_41670);
or U45798 (N_45798,N_40893,N_40429);
xor U45799 (N_45799,N_41128,N_40286);
or U45800 (N_45800,N_41859,N_44571);
nand U45801 (N_45801,N_42792,N_42230);
or U45802 (N_45802,N_41705,N_43383);
or U45803 (N_45803,N_41286,N_42228);
nand U45804 (N_45804,N_44953,N_41602);
xnor U45805 (N_45805,N_44711,N_40102);
xor U45806 (N_45806,N_44362,N_41947);
nor U45807 (N_45807,N_44423,N_44501);
nand U45808 (N_45808,N_42527,N_40303);
or U45809 (N_45809,N_42366,N_43111);
and U45810 (N_45810,N_43258,N_41915);
nand U45811 (N_45811,N_44729,N_42124);
nand U45812 (N_45812,N_40713,N_41317);
xor U45813 (N_45813,N_40215,N_42768);
and U45814 (N_45814,N_41248,N_44064);
xor U45815 (N_45815,N_44007,N_42360);
nor U45816 (N_45816,N_41388,N_41606);
xnor U45817 (N_45817,N_40658,N_40934);
nand U45818 (N_45818,N_40702,N_43558);
and U45819 (N_45819,N_40764,N_40129);
nand U45820 (N_45820,N_42644,N_41417);
or U45821 (N_45821,N_42238,N_41514);
xor U45822 (N_45822,N_43043,N_43470);
and U45823 (N_45823,N_40484,N_43278);
xor U45824 (N_45824,N_42760,N_44180);
nor U45825 (N_45825,N_42489,N_41724);
and U45826 (N_45826,N_44555,N_42148);
or U45827 (N_45827,N_40943,N_43080);
nor U45828 (N_45828,N_41574,N_40695);
nand U45829 (N_45829,N_40382,N_44432);
and U45830 (N_45830,N_41260,N_42193);
xnor U45831 (N_45831,N_40466,N_41131);
nand U45832 (N_45832,N_44581,N_42325);
nand U45833 (N_45833,N_41472,N_42283);
xor U45834 (N_45834,N_40726,N_43603);
nand U45835 (N_45835,N_41979,N_43641);
or U45836 (N_45836,N_40866,N_41390);
nand U45837 (N_45837,N_44063,N_43897);
and U45838 (N_45838,N_42289,N_40245);
and U45839 (N_45839,N_41331,N_42519);
nor U45840 (N_45840,N_40224,N_40127);
nand U45841 (N_45841,N_42702,N_43773);
and U45842 (N_45842,N_41006,N_41691);
or U45843 (N_45843,N_40410,N_43715);
nand U45844 (N_45844,N_41504,N_44741);
nand U45845 (N_45845,N_44998,N_41547);
nand U45846 (N_45846,N_40731,N_41137);
nand U45847 (N_45847,N_42359,N_40868);
or U45848 (N_45848,N_40541,N_41770);
and U45849 (N_45849,N_41865,N_41558);
or U45850 (N_45850,N_42879,N_41948);
nand U45851 (N_45851,N_41340,N_44531);
and U45852 (N_45852,N_40240,N_42501);
or U45853 (N_45853,N_40261,N_44373);
nor U45854 (N_45854,N_42346,N_43928);
nor U45855 (N_45855,N_44079,N_43353);
xnor U45856 (N_45856,N_43183,N_40107);
nor U45857 (N_45857,N_43311,N_43900);
nor U45858 (N_45858,N_42413,N_44011);
nand U45859 (N_45859,N_42570,N_41505);
and U45860 (N_45860,N_44690,N_43832);
and U45861 (N_45861,N_43438,N_43865);
xor U45862 (N_45862,N_42717,N_41132);
xor U45863 (N_45863,N_40650,N_41460);
nor U45864 (N_45864,N_43670,N_41201);
nor U45865 (N_45865,N_44876,N_41031);
xnor U45866 (N_45866,N_44492,N_43444);
nor U45867 (N_45867,N_42406,N_42572);
and U45868 (N_45868,N_40644,N_41958);
nor U45869 (N_45869,N_42504,N_40202);
nand U45870 (N_45870,N_40795,N_42790);
xor U45871 (N_45871,N_44504,N_40548);
nor U45872 (N_45872,N_41537,N_43678);
xnor U45873 (N_45873,N_40847,N_42309);
or U45874 (N_45874,N_41275,N_44207);
or U45875 (N_45875,N_41740,N_41650);
xnor U45876 (N_45876,N_43990,N_40991);
or U45877 (N_45877,N_41896,N_43100);
nor U45878 (N_45878,N_44340,N_44737);
nor U45879 (N_45879,N_40289,N_42804);
nor U45880 (N_45880,N_44448,N_43035);
xnor U45881 (N_45881,N_41961,N_40075);
nand U45882 (N_45882,N_41924,N_44222);
xor U45883 (N_45883,N_40352,N_41846);
nand U45884 (N_45884,N_43698,N_42752);
or U45885 (N_45885,N_41751,N_40711);
nor U45886 (N_45886,N_42226,N_43822);
nor U45887 (N_45887,N_44126,N_44578);
nand U45888 (N_45888,N_40380,N_42951);
and U45889 (N_45889,N_40509,N_43451);
nor U45890 (N_45890,N_42381,N_44759);
nand U45891 (N_45891,N_41681,N_43774);
nand U45892 (N_45892,N_42946,N_41370);
nand U45893 (N_45893,N_41925,N_41759);
or U45894 (N_45894,N_42718,N_43827);
nand U45895 (N_45895,N_42461,N_43069);
or U45896 (N_45896,N_43586,N_40198);
and U45897 (N_45897,N_43432,N_43608);
or U45898 (N_45898,N_41458,N_44672);
or U45899 (N_45899,N_43060,N_43534);
and U45900 (N_45900,N_42373,N_42745);
nand U45901 (N_45901,N_41439,N_40121);
nor U45902 (N_45902,N_40407,N_41269);
xnor U45903 (N_45903,N_42864,N_41238);
nor U45904 (N_45904,N_41352,N_42779);
xnor U45905 (N_45905,N_40922,N_44992);
xor U45906 (N_45906,N_41178,N_41239);
nor U45907 (N_45907,N_44944,N_40747);
xor U45908 (N_45908,N_40742,N_42914);
nand U45909 (N_45909,N_44293,N_40387);
nor U45910 (N_45910,N_42116,N_44358);
nand U45911 (N_45911,N_44597,N_41822);
or U45912 (N_45912,N_41486,N_42841);
nand U45913 (N_45913,N_41987,N_43870);
nand U45914 (N_45914,N_42010,N_42657);
nand U45915 (N_45915,N_43302,N_42207);
xor U45916 (N_45916,N_44762,N_40654);
nand U45917 (N_45917,N_43893,N_44489);
xnor U45918 (N_45918,N_42690,N_43620);
nor U45919 (N_45919,N_40090,N_42814);
nand U45920 (N_45920,N_42172,N_41588);
or U45921 (N_45921,N_40334,N_41229);
nor U45922 (N_45922,N_43099,N_41870);
or U45923 (N_45923,N_41980,N_40432);
and U45924 (N_45924,N_40923,N_43594);
nor U45925 (N_45925,N_42428,N_41982);
or U45926 (N_45926,N_41003,N_40553);
xnor U45927 (N_45927,N_42403,N_42668);
nor U45928 (N_45928,N_42123,N_44775);
nor U45929 (N_45929,N_40652,N_41333);
nor U45930 (N_45930,N_41293,N_41960);
nor U45931 (N_45931,N_40447,N_41888);
nor U45932 (N_45932,N_41853,N_43245);
and U45933 (N_45933,N_43875,N_40518);
xnor U45934 (N_45934,N_41697,N_40287);
and U45935 (N_45935,N_42142,N_40199);
and U45936 (N_45936,N_43243,N_40583);
or U45937 (N_45937,N_43978,N_44201);
nor U45938 (N_45938,N_40145,N_42016);
xnor U45939 (N_45939,N_41350,N_43999);
nor U45940 (N_45940,N_42553,N_40472);
or U45941 (N_45941,N_44519,N_41991);
nor U45942 (N_45942,N_44284,N_43203);
and U45943 (N_45943,N_40637,N_44606);
or U45944 (N_45944,N_44627,N_41930);
nor U45945 (N_45945,N_44436,N_40376);
nand U45946 (N_45946,N_42875,N_41904);
nand U45947 (N_45947,N_44372,N_42977);
nor U45948 (N_45948,N_41495,N_44978);
xnor U45949 (N_45949,N_42932,N_40497);
or U45950 (N_45950,N_42407,N_42991);
nor U45951 (N_45951,N_42862,N_40177);
or U45952 (N_45952,N_44853,N_43497);
xnor U45953 (N_45953,N_40788,N_41424);
nor U45954 (N_45954,N_41540,N_44127);
nor U45955 (N_45955,N_44917,N_44105);
nand U45956 (N_45956,N_40004,N_42259);
or U45957 (N_45957,N_42301,N_40355);
xor U45958 (N_45958,N_43193,N_44691);
nand U45959 (N_45959,N_43455,N_43265);
or U45960 (N_45960,N_41548,N_42984);
and U45961 (N_45961,N_40434,N_44317);
nand U45962 (N_45962,N_43545,N_44288);
and U45963 (N_45963,N_44995,N_43574);
nor U45964 (N_45964,N_42169,N_43601);
or U45965 (N_45965,N_40902,N_43693);
and U45966 (N_45966,N_40206,N_42838);
or U45967 (N_45967,N_43951,N_43861);
and U45968 (N_45968,N_44610,N_41285);
nand U45969 (N_45969,N_41369,N_43209);
or U45970 (N_45970,N_42786,N_44768);
nand U45971 (N_45971,N_43109,N_41345);
or U45972 (N_45972,N_43269,N_42341);
nor U45973 (N_45973,N_41277,N_43219);
xnor U45974 (N_45974,N_43025,N_41337);
nand U45975 (N_45975,N_41028,N_44258);
xor U45976 (N_45976,N_42912,N_43831);
or U45977 (N_45977,N_43550,N_44844);
or U45978 (N_45978,N_43888,N_42415);
or U45979 (N_45979,N_40634,N_44251);
and U45980 (N_45980,N_43713,N_41470);
xor U45981 (N_45981,N_43704,N_44771);
nor U45982 (N_45982,N_43575,N_43459);
and U45983 (N_45983,N_42585,N_44994);
nor U45984 (N_45984,N_43248,N_43946);
xor U45985 (N_45985,N_43560,N_43536);
nand U45986 (N_45986,N_41627,N_42996);
nor U45987 (N_45987,N_43454,N_41073);
and U45988 (N_45988,N_42534,N_42383);
or U45989 (N_45989,N_44279,N_41640);
nand U45990 (N_45990,N_41974,N_42685);
nand U45991 (N_45991,N_43335,N_43711);
and U45992 (N_45992,N_41296,N_40159);
nand U45993 (N_45993,N_44407,N_41773);
xor U45994 (N_45994,N_40928,N_42688);
xnor U45995 (N_45995,N_41567,N_43196);
xnor U45996 (N_45996,N_40616,N_41908);
nor U45997 (N_45997,N_41148,N_41839);
or U45998 (N_45998,N_44561,N_41628);
and U45999 (N_45999,N_44864,N_40314);
nand U46000 (N_46000,N_44351,N_40837);
or U46001 (N_46001,N_43595,N_44928);
or U46002 (N_46002,N_44049,N_41116);
or U46003 (N_46003,N_44861,N_40307);
nor U46004 (N_46004,N_42916,N_41747);
nand U46005 (N_46005,N_41613,N_44867);
and U46006 (N_46006,N_43068,N_40166);
and U46007 (N_46007,N_42312,N_40984);
or U46008 (N_46008,N_40544,N_44933);
and U46009 (N_46009,N_40774,N_42317);
or U46010 (N_46010,N_42619,N_43799);
or U46011 (N_46011,N_41280,N_41818);
and U46012 (N_46012,N_44227,N_42737);
nand U46013 (N_46013,N_43725,N_44579);
xnor U46014 (N_46014,N_41781,N_43295);
nor U46015 (N_46015,N_42637,N_42507);
xnor U46016 (N_46016,N_42000,N_44237);
nor U46017 (N_46017,N_44522,N_40448);
nor U46018 (N_46018,N_41259,N_42607);
or U46019 (N_46019,N_43649,N_41973);
or U46020 (N_46020,N_43515,N_41344);
nand U46021 (N_46021,N_42356,N_40954);
nor U46022 (N_46022,N_42577,N_42882);
nor U46023 (N_46023,N_42031,N_44988);
nand U46024 (N_46024,N_40181,N_41431);
nor U46025 (N_46025,N_44649,N_40972);
or U46026 (N_46026,N_43062,N_40998);
nor U46027 (N_46027,N_44457,N_44651);
nor U46028 (N_46028,N_40165,N_42444);
or U46029 (N_46029,N_41604,N_44271);
nand U46030 (N_46030,N_43836,N_41309);
and U46031 (N_46031,N_43945,N_40426);
nor U46032 (N_46032,N_44570,N_43160);
and U46033 (N_46033,N_43639,N_43224);
nor U46034 (N_46034,N_44377,N_41326);
nor U46035 (N_46035,N_40157,N_44596);
nand U46036 (N_46036,N_44751,N_42528);
nand U46037 (N_46037,N_40174,N_43609);
nor U46038 (N_46038,N_43652,N_40420);
nand U46039 (N_46039,N_43391,N_40887);
and U46040 (N_46040,N_42222,N_41494);
and U46041 (N_46041,N_43723,N_40855);
nor U46042 (N_46042,N_42894,N_42712);
or U46043 (N_46043,N_42433,N_43541);
xor U46044 (N_46044,N_42423,N_44421);
nand U46045 (N_46045,N_43878,N_41449);
and U46046 (N_46046,N_42789,N_44695);
and U46047 (N_46047,N_40318,N_43877);
nand U46048 (N_46048,N_44224,N_40449);
or U46049 (N_46049,N_40050,N_42488);
or U46050 (N_46050,N_44866,N_43277);
nand U46051 (N_46051,N_44296,N_40078);
and U46052 (N_46052,N_44383,N_44384);
nor U46053 (N_46053,N_42022,N_40353);
nand U46054 (N_46054,N_42164,N_41237);
or U46055 (N_46055,N_43961,N_42837);
nor U46056 (N_46056,N_44096,N_41021);
nand U46057 (N_46057,N_40709,N_40651);
xor U46058 (N_46058,N_42682,N_40397);
nand U46059 (N_46059,N_42231,N_41631);
or U46060 (N_46060,N_42266,N_42284);
nand U46061 (N_46061,N_40970,N_42028);
nand U46062 (N_46062,N_44665,N_40909);
and U46063 (N_46063,N_44426,N_40072);
and U46064 (N_46064,N_42502,N_40683);
nand U46065 (N_46065,N_41209,N_42993);
or U46066 (N_46066,N_43142,N_44405);
nor U46067 (N_46067,N_40577,N_40190);
nand U46068 (N_46068,N_43074,N_44150);
or U46069 (N_46069,N_40118,N_43134);
nor U46070 (N_46070,N_42975,N_40831);
xor U46071 (N_46071,N_43769,N_43117);
nor U46072 (N_46072,N_41812,N_41609);
xnor U46073 (N_46073,N_40048,N_42867);
xor U46074 (N_46074,N_40670,N_40319);
or U46075 (N_46075,N_40220,N_41410);
or U46076 (N_46076,N_43689,N_43939);
and U46077 (N_46077,N_40610,N_42347);
or U46078 (N_46078,N_41174,N_41120);
or U46079 (N_46079,N_44077,N_41986);
or U46080 (N_46080,N_42101,N_40424);
or U46081 (N_46081,N_43045,N_40692);
or U46082 (N_46082,N_42155,N_44473);
or U46083 (N_46083,N_44268,N_42003);
and U46084 (N_46084,N_40280,N_42643);
nor U46085 (N_46085,N_40238,N_42922);
and U46086 (N_46086,N_41879,N_41033);
or U46087 (N_46087,N_41294,N_41521);
nand U46088 (N_46088,N_44536,N_42285);
xnor U46089 (N_46089,N_42705,N_42399);
xnor U46090 (N_46090,N_42558,N_44776);
nor U46091 (N_46091,N_40900,N_40646);
or U46092 (N_46092,N_43802,N_44663);
and U46093 (N_46093,N_41316,N_40153);
xor U46094 (N_46094,N_42139,N_43819);
or U46095 (N_46095,N_40768,N_42070);
and U46096 (N_46096,N_41036,N_43368);
nand U46097 (N_46097,N_42918,N_44103);
xnor U46098 (N_46098,N_44927,N_44167);
nor U46099 (N_46099,N_41614,N_40870);
or U46100 (N_46100,N_44068,N_42114);
nor U46101 (N_46101,N_41467,N_43148);
nor U46102 (N_46102,N_40901,N_44884);
nor U46103 (N_46103,N_41445,N_40846);
nor U46104 (N_46104,N_41621,N_42693);
nor U46105 (N_46105,N_43124,N_40807);
or U46106 (N_46106,N_42161,N_42447);
and U46107 (N_46107,N_42037,N_40149);
xnor U46108 (N_46108,N_40776,N_44548);
nand U46109 (N_46109,N_44399,N_44658);
or U46110 (N_46110,N_40327,N_41851);
nand U46111 (N_46111,N_43168,N_40575);
or U46112 (N_46112,N_43914,N_40441);
or U46113 (N_46113,N_44774,N_43809);
nand U46114 (N_46114,N_43003,N_43492);
nor U46115 (N_46115,N_40545,N_44734);
nor U46116 (N_46116,N_40277,N_41966);
and U46117 (N_46117,N_41283,N_43800);
nand U46118 (N_46118,N_42858,N_43844);
or U46119 (N_46119,N_40063,N_43274);
and U46120 (N_46120,N_41695,N_41179);
or U46121 (N_46121,N_40754,N_41666);
xor U46122 (N_46122,N_44686,N_44609);
or U46123 (N_46123,N_43482,N_40883);
or U46124 (N_46124,N_42618,N_40328);
xor U46125 (N_46125,N_40138,N_43804);
nand U46126 (N_46126,N_44335,N_44000);
nor U46127 (N_46127,N_43175,N_40952);
xor U46128 (N_46128,N_42420,N_43785);
xnor U46129 (N_46129,N_44529,N_40370);
nand U46130 (N_46130,N_42262,N_44239);
nor U46131 (N_46131,N_42133,N_43284);
or U46132 (N_46132,N_42747,N_44058);
nand U46133 (N_46133,N_44871,N_43098);
or U46134 (N_46134,N_40440,N_43691);
nor U46135 (N_46135,N_42214,N_40117);
nand U46136 (N_46136,N_42700,N_41873);
or U46137 (N_46137,N_44484,N_43017);
nor U46138 (N_46138,N_41877,N_41437);
or U46139 (N_46139,N_41339,N_43133);
nand U46140 (N_46140,N_40036,N_44857);
nand U46141 (N_46141,N_42622,N_43593);
nand U46142 (N_46142,N_42592,N_42798);
nor U46143 (N_46143,N_41108,N_41796);
or U46144 (N_46144,N_41784,N_41267);
or U46145 (N_46145,N_42931,N_40003);
nor U46146 (N_46146,N_42587,N_44181);
xor U46147 (N_46147,N_44608,N_44783);
xnor U46148 (N_46148,N_44363,N_41464);
xor U46149 (N_46149,N_43494,N_41298);
xnor U46150 (N_46150,N_44502,N_40457);
and U46151 (N_46151,N_42598,N_43214);
or U46152 (N_46152,N_42311,N_42246);
nor U46153 (N_46153,N_42296,N_41531);
nand U46154 (N_46154,N_44123,N_43067);
xnor U46155 (N_46155,N_43816,N_40783);
xor U46156 (N_46156,N_44466,N_40549);
and U46157 (N_46157,N_43340,N_43734);
or U46158 (N_46158,N_44528,N_42758);
nor U46159 (N_46159,N_44445,N_42857);
and U46160 (N_46160,N_43696,N_44574);
nor U46161 (N_46161,N_41110,N_44787);
and U46162 (N_46162,N_43237,N_43672);
nor U46163 (N_46163,N_44673,N_44274);
nand U46164 (N_46164,N_43079,N_40507);
or U46165 (N_46165,N_41086,N_41162);
or U46166 (N_46166,N_44601,N_40291);
or U46167 (N_46167,N_43995,N_41191);
nor U46168 (N_46168,N_41421,N_42310);
nand U46169 (N_46169,N_40037,N_43604);
nand U46170 (N_46170,N_41964,N_42127);
nand U46171 (N_46171,N_41242,N_44782);
and U46172 (N_46172,N_43104,N_42280);
nor U46173 (N_46173,N_44903,N_43090);
or U46174 (N_46174,N_40055,N_41852);
nor U46175 (N_46175,N_40039,N_43582);
nand U46176 (N_46176,N_42182,N_41553);
nand U46177 (N_46177,N_43572,N_41591);
or U46178 (N_46178,N_41522,N_44375);
and U46179 (N_46179,N_44811,N_41303);
xnor U46180 (N_46180,N_44348,N_44503);
nand U46181 (N_46181,N_44446,N_44940);
xnor U46182 (N_46182,N_41024,N_43153);
and U46183 (N_46183,N_41430,N_44357);
or U46184 (N_46184,N_44010,N_43768);
and U46185 (N_46185,N_44336,N_41517);
and U46186 (N_46186,N_43926,N_41868);
nor U46187 (N_46187,N_40208,N_43210);
xnor U46188 (N_46188,N_43309,N_41063);
nor U46189 (N_46189,N_43264,N_44498);
nand U46190 (N_46190,N_43357,N_41198);
nor U46191 (N_46191,N_40609,N_44254);
nor U46192 (N_46192,N_40520,N_40336);
or U46193 (N_46193,N_40993,N_42057);
or U46194 (N_46194,N_43396,N_42640);
nand U46195 (N_46195,N_41820,N_42887);
nand U46196 (N_46196,N_42235,N_43167);
nor U46197 (N_46197,N_44324,N_42267);
or U46198 (N_46198,N_40366,N_42990);
or U46199 (N_46199,N_42162,N_42909);
nand U46200 (N_46200,N_40244,N_44331);
or U46201 (N_46201,N_43456,N_42192);
nor U46202 (N_46202,N_44078,N_42405);
nand U46203 (N_46203,N_44376,N_43189);
nor U46204 (N_46204,N_44835,N_44545);
xnor U46205 (N_46205,N_42288,N_40592);
and U46206 (N_46206,N_41434,N_40460);
nor U46207 (N_46207,N_42917,N_42704);
xnor U46208 (N_46208,N_44859,N_40487);
nand U46209 (N_46209,N_40746,N_43299);
nand U46210 (N_46210,N_42013,N_42401);
and U46211 (N_46211,N_44931,N_40377);
nand U46212 (N_46212,N_43155,N_42077);
nand U46213 (N_46213,N_40134,N_43597);
nand U46214 (N_46214,N_41783,N_44849);
nand U46215 (N_46215,N_41438,N_41394);
or U46216 (N_46216,N_40459,N_43871);
and U46217 (N_46217,N_43526,N_43077);
nand U46218 (N_46218,N_41916,N_43619);
and U46219 (N_46219,N_43088,N_42521);
xor U46220 (N_46220,N_42797,N_42054);
xnor U46221 (N_46221,N_42110,N_44977);
nand U46222 (N_46222,N_40241,N_44599);
xnor U46223 (N_46223,N_42062,N_43179);
nor U46224 (N_46224,N_41663,N_44553);
nand U46225 (N_46225,N_40281,N_44946);
or U46226 (N_46226,N_42065,N_40473);
or U46227 (N_46227,N_40150,N_42981);
xnor U46228 (N_46228,N_43565,N_41320);
nor U46229 (N_46229,N_44462,N_40710);
and U46230 (N_46230,N_42122,N_42540);
nand U46231 (N_46231,N_42379,N_40586);
or U46232 (N_46232,N_43676,N_41327);
xnor U46233 (N_46233,N_40052,N_42175);
or U46234 (N_46234,N_41016,N_40555);
nor U46235 (N_46235,N_44176,N_42281);
or U46236 (N_46236,N_43410,N_41090);
nand U46237 (N_46237,N_44761,N_41569);
or U46238 (N_46238,N_43251,N_44902);
xor U46239 (N_46239,N_41527,N_41648);
or U46240 (N_46240,N_40828,N_44842);
or U46241 (N_46241,N_40148,N_40200);
and U46242 (N_46242,N_43828,N_43849);
xor U46243 (N_46243,N_40163,N_41308);
xor U46244 (N_46244,N_44930,N_43409);
xor U46245 (N_46245,N_44720,N_41585);
nor U46246 (N_46246,N_40712,N_41963);
nor U46247 (N_46247,N_40160,N_42199);
nand U46248 (N_46248,N_44125,N_44766);
nor U46249 (N_46249,N_41592,N_43166);
nand U46250 (N_46250,N_42371,N_43886);
or U46251 (N_46251,N_40906,N_42866);
and U46252 (N_46252,N_41737,N_40402);
nand U46253 (N_46253,N_43001,N_40378);
or U46254 (N_46254,N_43671,N_44688);
and U46255 (N_46255,N_40422,N_42531);
or U46256 (N_46256,N_43618,N_41202);
nand U46257 (N_46257,N_44558,N_44108);
or U46258 (N_46258,N_40136,N_43948);
nand U46259 (N_46259,N_42888,N_43122);
and U46260 (N_46260,N_40872,N_42243);
xnor U46261 (N_46261,N_41186,N_44186);
and U46262 (N_46262,N_44594,N_41561);
nand U46263 (N_46263,N_42906,N_41085);
xor U46264 (N_46264,N_41155,N_44572);
or U46265 (N_46265,N_44464,N_40630);
xnor U46266 (N_46266,N_41367,N_44657);
xor U46267 (N_46267,N_44708,N_41404);
nand U46268 (N_46268,N_42543,N_43746);
nor U46269 (N_46269,N_43319,N_42529);
nor U46270 (N_46270,N_41223,N_40735);
nor U46271 (N_46271,N_43029,N_43569);
nand U46272 (N_46272,N_42131,N_43782);
nor U46273 (N_46273,N_43434,N_41715);
and U46274 (N_46274,N_41061,N_44833);
xor U46275 (N_46275,N_41545,N_42107);
and U46276 (N_46276,N_44828,N_43587);
nand U46277 (N_46277,N_41972,N_40611);
xor U46278 (N_46278,N_41461,N_42088);
and U46279 (N_46279,N_41645,N_40648);
nand U46280 (N_46280,N_40891,N_42253);
and U46281 (N_46281,N_40967,N_42777);
or U46282 (N_46282,N_40676,N_40758);
nor U46283 (N_46283,N_42393,N_44497);
or U46284 (N_46284,N_40502,N_44719);
xor U46285 (N_46285,N_41690,N_44642);
nor U46286 (N_46286,N_43347,N_41962);
nand U46287 (N_46287,N_42933,N_44261);
nand U46288 (N_46288,N_44702,N_44276);
xor U46289 (N_46289,N_42713,N_41484);
or U46290 (N_46290,N_42756,N_43403);
nand U46291 (N_46291,N_42583,N_41365);
nand U46292 (N_46292,N_43524,N_42436);
nor U46293 (N_46293,N_42796,N_41934);
or U46294 (N_46294,N_41184,N_41677);
nand U46295 (N_46295,N_42696,N_42586);
xor U46296 (N_46296,N_40015,N_41564);
and U46297 (N_46297,N_44212,N_44322);
or U46298 (N_46298,N_43703,N_44139);
nand U46299 (N_46299,N_42732,N_40912);
nor U46300 (N_46300,N_44062,N_40099);
xor U46301 (N_46301,N_44979,N_44217);
or U46302 (N_46302,N_41918,N_43576);
and U46303 (N_46303,N_44117,N_42947);
xor U46304 (N_46304,N_40763,N_41790);
xnor U46305 (N_46305,N_40335,N_40572);
and U46306 (N_46306,N_41524,N_44908);
nor U46307 (N_46307,N_40598,N_41222);
xor U46308 (N_46308,N_44056,N_42513);
nand U46309 (N_46309,N_41160,N_44295);
and U46310 (N_46310,N_43958,N_43797);
nand U46311 (N_46311,N_41787,N_40757);
or U46312 (N_46312,N_43101,N_44380);
xnor U46313 (N_46313,N_43894,N_42414);
nor U46314 (N_46314,N_44270,N_41300);
nand U46315 (N_46315,N_43236,N_43801);
or U46316 (N_46316,N_41668,N_42774);
or U46317 (N_46317,N_42138,N_44732);
and U46318 (N_46318,N_43445,N_42463);
and U46319 (N_46319,N_40772,N_42239);
nand U46320 (N_46320,N_40722,N_43917);
nor U46321 (N_46321,N_42980,N_43359);
or U46322 (N_46322,N_42335,N_44506);
nor U46323 (N_46323,N_41264,N_43663);
and U46324 (N_46324,N_41891,N_41501);
xnor U46325 (N_46325,N_40907,N_41377);
nor U46326 (N_46326,N_43653,N_40001);
or U46327 (N_46327,N_42913,N_42709);
and U46328 (N_46328,N_40111,N_41619);
and U46329 (N_46329,N_42091,N_41258);
nor U46330 (N_46330,N_44655,N_43965);
and U46331 (N_46331,N_43004,N_43164);
and U46332 (N_46332,N_43362,N_40803);
or U46333 (N_46333,N_42323,N_42294);
or U46334 (N_46334,N_40699,N_42876);
nand U46335 (N_46335,N_42546,N_42538);
nand U46336 (N_46336,N_43275,N_42548);
or U46337 (N_46337,N_42485,N_41977);
nand U46338 (N_46338,N_44638,N_42135);
or U46339 (N_46339,N_40808,N_40823);
nand U46340 (N_46340,N_40714,N_40083);
nand U46341 (N_46341,N_41667,N_41324);
xnor U46342 (N_46342,N_41249,N_40511);
xnor U46343 (N_46343,N_40830,N_40927);
and U46344 (N_46344,N_42532,N_42451);
nand U46345 (N_46345,N_42466,N_40737);
nor U46346 (N_46346,N_43457,N_42092);
nor U46347 (N_46347,N_44914,N_40642);
xnor U46348 (N_46348,N_44115,N_41408);
or U46349 (N_46349,N_41256,N_44518);
nand U46350 (N_46350,N_41765,N_40195);
nand U46351 (N_46351,N_44756,N_43448);
or U46352 (N_46352,N_44095,N_40771);
xor U46353 (N_46353,N_44569,N_40988);
or U46354 (N_46354,N_41100,N_42872);
nor U46355 (N_46355,N_41067,N_40259);
xnor U46356 (N_46356,N_42058,N_40848);
or U46357 (N_46357,N_43039,N_43665);
and U46358 (N_46358,N_43694,N_44618);
xnor U46359 (N_46359,N_43304,N_44101);
nand U46360 (N_46360,N_44427,N_42632);
nand U46361 (N_46361,N_43970,N_44640);
xnor U46362 (N_46362,N_43566,N_42039);
nor U46363 (N_46363,N_41122,N_40228);
or U46364 (N_46364,N_42788,N_44488);
and U46365 (N_46365,N_44109,N_43254);
xor U46366 (N_46366,N_40814,N_41109);
and U46367 (N_46367,N_42973,N_40169);
nor U46368 (N_46368,N_41882,N_43772);
xor U46369 (N_46369,N_43927,N_43055);
xor U46370 (N_46370,N_43440,N_40105);
nor U46371 (N_46371,N_42470,N_41610);
xnor U46372 (N_46372,N_44580,N_44240);
nand U46373 (N_46373,N_43042,N_41804);
xor U46374 (N_46374,N_41465,N_41079);
and U46375 (N_46375,N_42236,N_41815);
nor U46376 (N_46376,N_42621,N_41094);
and U46377 (N_46377,N_44997,N_42506);
or U46378 (N_46378,N_41487,N_40905);
xnor U46379 (N_46379,N_44343,N_43220);
nor U46380 (N_46380,N_40170,N_43192);
or U46381 (N_46381,N_41624,N_43960);
and U46382 (N_46382,N_44780,N_41107);
and U46383 (N_46383,N_43539,N_41282);
xnor U46384 (N_46384,N_43227,N_42045);
nand U46385 (N_46385,N_42563,N_44521);
and U46386 (N_46386,N_40012,N_40231);
nand U46387 (N_46387,N_43270,N_42098);
and U46388 (N_46388,N_43114,N_44177);
nor U46389 (N_46389,N_44993,N_42655);
nand U46390 (N_46390,N_40849,N_43674);
or U46391 (N_46391,N_43547,N_41788);
nand U46392 (N_46392,N_42145,N_44818);
xnor U46393 (N_46393,N_41318,N_41197);
or U46394 (N_46394,N_40488,N_41945);
xnor U46395 (N_46395,N_40750,N_43102);
nor U46396 (N_46396,N_44283,N_41216);
xor U46397 (N_46397,N_40268,N_43718);
nand U46398 (N_46398,N_44169,N_43418);
nor U46399 (N_46399,N_42487,N_43008);
nand U46400 (N_46400,N_42624,N_44110);
nand U46401 (N_46401,N_42860,N_42146);
nor U46402 (N_46402,N_42069,N_40065);
and U46403 (N_46403,N_41176,N_41835);
and U46404 (N_46404,N_42008,N_40506);
nor U46405 (N_46405,N_42206,N_44231);
nor U46406 (N_46406,N_44465,N_42490);
xnor U46407 (N_46407,N_44812,N_44406);
nand U46408 (N_46408,N_44410,N_43453);
xor U46409 (N_46409,N_40140,N_42157);
nand U46410 (N_46410,N_41526,N_40079);
nand U46411 (N_46411,N_42261,N_44575);
and U46412 (N_46412,N_44156,N_44394);
and U46413 (N_46413,N_43433,N_40020);
or U46414 (N_46414,N_40056,N_41998);
or U46415 (N_46415,N_43158,N_40253);
xor U46416 (N_46416,N_43202,N_41017);
xor U46417 (N_46417,N_42904,N_42115);
or U46418 (N_46418,N_43912,N_44047);
nand U46419 (N_46419,N_44855,N_42095);
and U46420 (N_46420,N_40741,N_43896);
or U46421 (N_46421,N_44970,N_44976);
xnor U46422 (N_46422,N_41347,N_44438);
nand U46423 (N_46423,N_41170,N_42884);
or U46424 (N_46424,N_41348,N_42075);
xor U46425 (N_46425,N_42595,N_41243);
nor U46426 (N_46426,N_44616,N_43798);
or U46427 (N_46427,N_42613,N_41295);
nor U46428 (N_46428,N_40008,N_42958);
or U46429 (N_46429,N_41481,N_43084);
or U46430 (N_46430,N_40496,N_41271);
and U46431 (N_46431,N_43267,N_42179);
nor U46432 (N_46432,N_41803,N_42590);
nor U46433 (N_46433,N_40343,N_43753);
nand U46434 (N_46434,N_41732,N_42197);
or U46435 (N_46435,N_43617,N_43683);
or U46436 (N_46436,N_40230,N_42571);
xor U46437 (N_46437,N_44654,N_41173);
nor U46438 (N_46438,N_40374,N_40643);
xor U46439 (N_46439,N_40860,N_44300);
or U46440 (N_46440,N_41830,N_40531);
nand U46441 (N_46441,N_41078,N_40667);
nor U46442 (N_46442,N_42615,N_44941);
and U46443 (N_46443,N_44450,N_42211);
xor U46444 (N_46444,N_43450,N_40179);
xnor U46445 (N_46445,N_44135,N_40255);
or U46446 (N_46446,N_44955,N_40186);
xnor U46447 (N_46447,N_40112,N_43625);
and U46448 (N_46448,N_43018,N_41443);
and U46449 (N_46449,N_40767,N_42898);
or U46450 (N_46450,N_43726,N_44730);
or U46451 (N_46451,N_41842,N_43732);
and U46452 (N_46452,N_42596,N_44974);
xor U46453 (N_46453,N_41543,N_44634);
and U46454 (N_46454,N_41771,N_42011);
and U46455 (N_46455,N_44971,N_43075);
nand U46456 (N_46456,N_41920,N_42938);
or U46457 (N_46457,N_43835,N_41077);
nand U46458 (N_46458,N_42329,N_41503);
nand U46459 (N_46459,N_40877,N_41866);
or U46460 (N_46460,N_41500,N_40503);
or U46461 (N_46461,N_42793,N_43998);
nor U46462 (N_46462,N_40226,N_43215);
nand U46463 (N_46463,N_40705,N_43188);
xor U46464 (N_46464,N_44984,N_43710);
or U46465 (N_46465,N_44053,N_41157);
nor U46466 (N_46466,N_43279,N_41489);
nor U46467 (N_46467,N_44889,N_44038);
nand U46468 (N_46468,N_40580,N_41169);
and U46469 (N_46469,N_42536,N_44639);
or U46470 (N_46470,N_41236,N_44418);
nand U46471 (N_46471,N_40406,N_40465);
nor U46472 (N_46472,N_40132,N_43370);
and U46473 (N_46473,N_41194,N_42679);
nand U46474 (N_46474,N_42907,N_40393);
or U46475 (N_46475,N_44515,N_40178);
nand U46476 (N_46476,N_42306,N_40706);
nor U46477 (N_46477,N_41011,N_41546);
or U46478 (N_46478,N_43568,N_43962);
xnor U46479 (N_46479,N_43416,N_40196);
and U46480 (N_46480,N_40703,N_42225);
or U46481 (N_46481,N_44147,N_41065);
nand U46482 (N_46482,N_41603,N_41473);
nand U46483 (N_46483,N_43152,N_41674);
or U46484 (N_46484,N_44604,N_42153);
nor U46485 (N_46485,N_40456,N_44499);
and U46486 (N_46486,N_40219,N_44424);
and U46487 (N_46487,N_41146,N_42205);
nand U46488 (N_46488,N_42552,N_44680);
nand U46489 (N_46489,N_41459,N_42257);
or U46490 (N_46490,N_43720,N_40444);
and U46491 (N_46491,N_42928,N_41617);
and U46492 (N_46492,N_41922,N_40990);
nand U46493 (N_46493,N_42140,N_42736);
nand U46494 (N_46494,N_40794,N_41728);
and U46495 (N_46495,N_44507,N_41012);
or U46496 (N_46496,N_43070,N_42784);
xor U46497 (N_46497,N_40624,N_40412);
nor U46498 (N_46498,N_41188,N_44253);
nand U46499 (N_46499,N_41196,N_43216);
or U46500 (N_46500,N_42603,N_42901);
nor U46501 (N_46501,N_43139,N_40864);
or U46502 (N_46502,N_44678,N_43792);
or U46503 (N_46503,N_44896,N_41038);
nor U46504 (N_46504,N_42656,N_40266);
nor U46505 (N_46505,N_40612,N_44286);
or U46506 (N_46506,N_40239,N_40346);
xor U46507 (N_46507,N_44030,N_41310);
xor U46508 (N_46508,N_41623,N_44459);
and U46509 (N_46509,N_44060,N_43911);
nor U46510 (N_46510,N_44339,N_43157);
or U46511 (N_46511,N_41498,N_43687);
and U46512 (N_46512,N_44434,N_44191);
xor U46513 (N_46513,N_43918,N_43664);
nor U46514 (N_46514,N_42324,N_43783);
nand U46515 (N_46515,N_41556,N_40810);
or U46516 (N_46516,N_40815,N_41228);
nor U46517 (N_46517,N_41889,N_42889);
xor U46518 (N_46518,N_40130,N_41502);
and U46519 (N_46519,N_41384,N_44684);
nor U46520 (N_46520,N_44155,N_43272);
or U46521 (N_46521,N_42535,N_40109);
nand U46522 (N_46522,N_44547,N_43131);
nand U46523 (N_46523,N_40821,N_43520);
and U46524 (N_46524,N_40074,N_41448);
nand U46525 (N_46525,N_44805,N_40880);
nand U46526 (N_46526,N_42994,N_42588);
xnor U46527 (N_46527,N_42812,N_40061);
or U46528 (N_46528,N_41511,N_44567);
nor U46529 (N_46529,N_42611,N_44037);
and U46530 (N_46530,N_44791,N_43916);
nand U46531 (N_46531,N_44893,N_43468);
nand U46532 (N_46532,N_43709,N_43430);
or U46533 (N_46533,N_40982,N_43714);
nor U46534 (N_46534,N_43910,N_44878);
and U46535 (N_46535,N_44932,N_40292);
nor U46536 (N_46536,N_44099,N_40607);
xor U46537 (N_46537,N_42475,N_42652);
nand U46538 (N_46538,N_40707,N_44989);
xnor U46539 (N_46539,N_44926,N_42252);
or U46540 (N_46540,N_40937,N_40070);
xor U46541 (N_46541,N_43449,N_41314);
nand U46542 (N_46542,N_40839,N_41583);
and U46543 (N_46543,N_40756,N_43546);
xnor U46544 (N_46544,N_43259,N_40833);
and U46545 (N_46545,N_42015,N_41401);
nor U46546 (N_46546,N_42941,N_44151);
or U46547 (N_46547,N_41910,N_40461);
nand U46548 (N_46548,N_43255,N_42545);
nor U46549 (N_46549,N_40890,N_44584);
and U46550 (N_46550,N_40095,N_42801);
nand U46551 (N_46551,N_42650,N_43425);
or U46552 (N_46552,N_40671,N_40184);
or U46553 (N_46553,N_40002,N_41480);
nor U46554 (N_46554,N_42533,N_42362);
or U46555 (N_46555,N_43427,N_43518);
nand U46556 (N_46556,N_44809,N_40532);
nor U46557 (N_46557,N_41570,N_40679);
and U46558 (N_46558,N_40490,N_40191);
nor U46559 (N_46559,N_44291,N_44565);
nor U46560 (N_46560,N_42020,N_42776);
nor U46561 (N_46561,N_41278,N_41954);
nor U46562 (N_46562,N_41518,N_44220);
or U46563 (N_46563,N_40665,N_44540);
nor U46564 (N_46564,N_40262,N_40673);
xor U46565 (N_46565,N_43869,N_40326);
or U46566 (N_46566,N_42919,N_42351);
nor U46567 (N_46567,N_40437,N_41476);
nor U46568 (N_46568,N_44164,N_43744);
and U46569 (N_46569,N_42083,N_44806);
or U46570 (N_46570,N_43841,N_41288);
xor U46571 (N_46571,N_40315,N_43280);
nor U46572 (N_46572,N_43330,N_43868);
nor U46573 (N_46573,N_40677,N_41050);
and U46574 (N_46574,N_40500,N_42180);
nor U46575 (N_46575,N_40897,N_44369);
or U46576 (N_46576,N_41290,N_40197);
xnor U46577 (N_46577,N_42358,N_44149);
or U46578 (N_46578,N_43765,N_42486);
nor U46579 (N_46579,N_43944,N_43636);
and U46580 (N_46580,N_40840,N_44386);
xnor U46581 (N_46581,N_44189,N_44121);
nor U46582 (N_46582,N_41220,N_44483);
nor U46583 (N_46583,N_43947,N_42234);
xor U46584 (N_46584,N_41647,N_44157);
or U46585 (N_46585,N_43745,N_44733);
nand U46586 (N_46586,N_40139,N_40144);
nor U46587 (N_46587,N_41257,N_43161);
xnor U46588 (N_46588,N_43968,N_40782);
or U46589 (N_46589,N_40047,N_42878);
nand U46590 (N_46590,N_42630,N_43034);
or U46591 (N_46591,N_40857,N_40142);
xor U46592 (N_46592,N_44003,N_40167);
or U46593 (N_46593,N_40966,N_44021);
nor U46594 (N_46594,N_44701,N_44557);
xnor U46595 (N_46595,N_41957,N_42287);
or U46596 (N_46596,N_40589,N_42514);
nor U46597 (N_46597,N_42939,N_41386);
or U46598 (N_46598,N_42481,N_41497);
and U46599 (N_46599,N_41035,N_44629);
nor U46600 (N_46600,N_40471,N_43925);
nand U46601 (N_46601,N_42361,N_42217);
and U46602 (N_46602,N_44773,N_40391);
or U46603 (N_46603,N_44807,N_42278);
xnor U46604 (N_46604,N_44413,N_44906);
xor U46605 (N_46605,N_44826,N_43145);
and U46606 (N_46606,N_42471,N_43379);
and U46607 (N_46607,N_44661,N_44040);
and U46608 (N_46608,N_42839,N_41499);
nor U46609 (N_46609,N_41087,N_40341);
xnor U46610 (N_46610,N_44272,N_44192);
nand U46611 (N_46611,N_41530,N_42256);
nand U46612 (N_46612,N_41907,N_41456);
xnor U46613 (N_46613,N_42150,N_41639);
xnor U46614 (N_46614,N_41409,N_40992);
xor U46615 (N_46615,N_43530,N_43907);
and U46616 (N_46616,N_40843,N_42869);
nor U46617 (N_46617,N_42368,N_44808);
nand U46618 (N_46618,N_44802,N_40601);
nor U46619 (N_46619,N_43890,N_41626);
or U46620 (N_46620,N_41354,N_43472);
or U46621 (N_46621,N_42983,N_41115);
xnor U46622 (N_46622,N_43205,N_44481);
nand U46623 (N_46623,N_44959,N_40246);
and U46624 (N_46624,N_41733,N_41817);
xnor U46625 (N_46625,N_43010,N_41441);
and U46626 (N_46626,N_44477,N_41005);
nand U46627 (N_46627,N_42807,N_44769);
nor U46628 (N_46628,N_41976,N_44677);
and U46629 (N_46629,N_43283,N_44748);
and U46630 (N_46630,N_42102,N_41466);
or U46631 (N_46631,N_42479,N_41049);
nand U46632 (N_46632,N_41468,N_42268);
nor U46633 (N_46633,N_41138,N_40951);
or U46634 (N_46634,N_44975,N_43750);
xor U46635 (N_46635,N_44152,N_43614);
xor U46636 (N_46636,N_40903,N_41074);
xnor U46637 (N_46637,N_43361,N_40367);
and U46638 (N_46638,N_43793,N_44564);
nand U46639 (N_46639,N_40932,N_43128);
nand U46640 (N_46640,N_44187,N_40021);
xnor U46641 (N_46641,N_41471,N_40405);
nand U46642 (N_46642,N_40888,N_44332);
nand U46643 (N_46643,N_43012,N_41562);
and U46644 (N_46644,N_40413,N_43360);
or U46645 (N_46645,N_40749,N_43113);
or U46646 (N_46646,N_42701,N_40910);
and U46647 (N_46647,N_42995,N_40981);
nor U46648 (N_46648,N_40227,N_44017);
nand U46649 (N_46649,N_44132,N_40576);
nor U46650 (N_46650,N_42117,N_44671);
and U46651 (N_46651,N_42510,N_40680);
or U46652 (N_46652,N_44225,N_44598);
or U46653 (N_46653,N_41881,N_41185);
nor U46654 (N_46654,N_43863,N_41118);
or U46655 (N_46655,N_43615,N_43643);
xor U46656 (N_46656,N_44246,N_44214);
or U46657 (N_46657,N_44052,N_40285);
xor U46658 (N_46658,N_42129,N_41833);
nand U46659 (N_46659,N_44419,N_40945);
or U46660 (N_46660,N_40542,N_42634);
nand U46661 (N_46661,N_42935,N_44922);
or U46662 (N_46662,N_41598,N_40693);
nor U46663 (N_46663,N_44894,N_43996);
and U46664 (N_46664,N_44646,N_41596);
or U46665 (N_46665,N_44118,N_40041);
nand U46666 (N_46666,N_44821,N_43556);
xor U46667 (N_46667,N_40950,N_44256);
nand U46668 (N_46668,N_41642,N_40863);
nand U46669 (N_46669,N_41698,N_40587);
xnor U46670 (N_46670,N_41725,N_40960);
or U46671 (N_46671,N_44041,N_44760);
or U46672 (N_46672,N_44066,N_41597);
nand U46673 (N_46673,N_42900,N_44951);
nor U46674 (N_46674,N_43610,N_40128);
nand U46675 (N_46675,N_43616,N_41117);
nor U46676 (N_46676,N_44408,N_42896);
and U46677 (N_46677,N_43400,N_41802);
or U46678 (N_46678,N_43656,N_44912);
nand U46679 (N_46679,N_42416,N_44260);
xnor U46680 (N_46680,N_41284,N_41066);
nor U46681 (N_46681,N_43373,N_40898);
xnor U46682 (N_46682,N_42551,N_40933);
nand U46683 (N_46683,N_44285,N_42419);
nor U46684 (N_46684,N_42920,N_41475);
xnor U46685 (N_46685,N_41797,N_43013);
xnor U46686 (N_46686,N_41738,N_42691);
or U46687 (N_46687,N_42868,N_42733);
xor U46688 (N_46688,N_44625,N_42188);
or U46689 (N_46689,N_40087,N_40914);
and U46690 (N_46690,N_41153,N_44083);
nor U46691 (N_46691,N_43784,N_42970);
nor U46692 (N_46692,N_40188,N_42773);
nor U46693 (N_46693,N_41212,N_43992);
nand U46694 (N_46694,N_43021,N_44967);
xnor U46695 (N_46695,N_41469,N_44264);
nand U46696 (N_46696,N_41057,N_43859);
and U46697 (N_46697,N_44883,N_40203);
xnor U46698 (N_46698,N_42078,N_41594);
nor U46699 (N_46699,N_44925,N_43081);
or U46700 (N_46700,N_44789,N_43401);
or U46701 (N_46701,N_41506,N_44026);
nand U46702 (N_46702,N_43345,N_41349);
or U46703 (N_46703,N_40124,N_41563);
or U46704 (N_46704,N_42232,N_40046);
or U46705 (N_46705,N_44043,N_43147);
nand U46706 (N_46706,N_41405,N_41630);
or U46707 (N_46707,N_44885,N_41052);
nand U46708 (N_46708,N_44731,N_44073);
xor U46709 (N_46709,N_41568,N_41192);
or U46710 (N_46710,N_40919,N_42469);
xor U46711 (N_46711,N_44615,N_41654);
nand U46712 (N_46712,N_43976,N_43474);
or U46713 (N_46713,N_44378,N_44374);
or U46714 (N_46714,N_40696,N_43931);
xor U46715 (N_46715,N_43384,N_40537);
and U46716 (N_46716,N_43761,N_40505);
nor U46717 (N_46717,N_42081,N_40229);
and U46718 (N_46718,N_40257,N_44359);
or U46719 (N_46719,N_40962,N_40789);
or U46720 (N_46720,N_44785,N_41253);
and U46721 (N_46721,N_44392,N_40080);
nand U46722 (N_46722,N_43864,N_44104);
or U46723 (N_46723,N_44136,N_42305);
xor U46724 (N_46724,N_42597,N_41113);
nand U46725 (N_46725,N_41554,N_42808);
nand U46726 (N_46726,N_42249,N_40439);
nand U46727 (N_46727,N_42897,N_41845);
nor U46728 (N_46728,N_41809,N_43579);
nor U46729 (N_46729,N_41825,N_42833);
nand U46730 (N_46730,N_44509,N_44148);
nor U46731 (N_46731,N_44106,N_40904);
nor U46732 (N_46732,N_40066,N_40486);
or U46733 (N_46733,N_44800,N_42654);
xor U46734 (N_46734,N_40871,N_41141);
nand U46735 (N_46735,N_42659,N_43895);
nand U46736 (N_46736,N_42272,N_43540);
or U46737 (N_46737,N_40254,N_42221);
nand U46738 (N_46738,N_42046,N_41041);
xnor U46739 (N_46739,N_40014,N_44356);
nor U46740 (N_46740,N_42395,N_41477);
or U46741 (N_46741,N_40686,N_44700);
and U46742 (N_46742,N_44621,N_44267);
and U46743 (N_46743,N_44514,N_42560);
nor U46744 (N_46744,N_40947,N_42338);
or U46745 (N_46745,N_44470,N_40242);
xor U46746 (N_46746,N_42387,N_43176);
nand U46747 (N_46747,N_41064,N_43204);
nor U46748 (N_46748,N_44815,N_44400);
or U46749 (N_46749,N_42446,N_40269);
or U46750 (N_46750,N_44577,N_41330);
and U46751 (N_46751,N_40462,N_41092);
and U46752 (N_46752,N_41772,N_42645);
xnor U46753 (N_46753,N_42795,N_40663);
nand U46754 (N_46754,N_41425,N_42770);
or U46755 (N_46755,N_41678,N_44962);
xor U46756 (N_46756,N_42664,N_42418);
nand U46757 (N_46757,N_44957,N_40874);
and U46758 (N_46758,N_42956,N_42998);
and U46759 (N_46759,N_44713,N_43086);
or U46760 (N_46760,N_41913,N_40955);
or U46761 (N_46761,N_40283,N_44779);
or U46762 (N_46762,N_43201,N_43551);
nand U46763 (N_46763,N_41397,N_44337);
and U46764 (N_46764,N_41726,N_40739);
and U46765 (N_46765,N_44200,N_43533);
nand U46766 (N_46766,N_43120,N_41800);
xor U46767 (N_46767,N_44116,N_41936);
or U46768 (N_46768,N_42408,N_43940);
xnor U46769 (N_46769,N_43942,N_41287);
xnor U46770 (N_46770,N_41270,N_42649);
nor U46771 (N_46771,N_42354,N_42715);
nand U46772 (N_46772,N_43065,N_43256);
or U46773 (N_46773,N_40973,N_42871);
nor U46774 (N_46774,N_43331,N_41897);
xnor U46775 (N_46775,N_44404,N_42103);
xor U46776 (N_46776,N_41933,N_40212);
xor U46777 (N_46777,N_42223,N_44918);
nand U46778 (N_46778,N_40204,N_42721);
or U46779 (N_46779,N_44242,N_42134);
or U46780 (N_46780,N_43987,N_40647);
nor U46781 (N_46781,N_42394,N_43721);
nor U46782 (N_46782,N_43767,N_42629);
nand U46783 (N_46783,N_42191,N_42441);
nor U46784 (N_46784,N_42255,N_42821);
nor U46785 (N_46785,N_42750,N_42516);
and U46786 (N_46786,N_42431,N_43475);
nor U46787 (N_46787,N_44329,N_43191);
xnor U46788 (N_46788,N_42212,N_44950);
and U46789 (N_46789,N_40029,N_41407);
or U46790 (N_46790,N_41039,N_41361);
and U46791 (N_46791,N_44666,N_43635);
xor U46792 (N_46792,N_42924,N_41491);
nand U46793 (N_46793,N_43591,N_44163);
or U46794 (N_46794,N_40704,N_41158);
nor U46795 (N_46795,N_44075,N_43795);
nand U46796 (N_46796,N_41254,N_40698);
and U46797 (N_46797,N_43431,N_43481);
and U46798 (N_46798,N_41779,N_42295);
xor U46799 (N_46799,N_43588,N_43903);
nand U46800 (N_46800,N_43076,N_42494);
or U46801 (N_46801,N_43262,N_41956);
nor U46802 (N_46802,N_43006,N_43132);
or U46803 (N_46803,N_42899,N_40786);
xnor U46804 (N_46804,N_42610,N_44390);
and U46805 (N_46805,N_42526,N_44085);
and U46806 (N_46806,N_42729,N_44819);
xor U46807 (N_46807,N_41372,N_44863);
nor U46808 (N_46808,N_42775,N_42213);
nand U46809 (N_46809,N_40097,N_44044);
xnor U46810 (N_46810,N_42697,N_41381);
or U46811 (N_46811,N_40064,N_43989);
xnor U46812 (N_46812,N_40985,N_40976);
nand U46813 (N_46813,N_41001,N_40617);
nand U46814 (N_46814,N_43032,N_42778);
and U46815 (N_46815,N_41084,N_40684);
nand U46816 (N_46816,N_44057,N_42683);
and U46817 (N_46817,N_42761,N_42856);
or U46818 (N_46818,N_43461,N_40398);
nand U46819 (N_46819,N_40421,N_40659);
nor U46820 (N_46820,N_42927,N_42279);
or U46821 (N_46821,N_41847,N_40533);
or U46822 (N_46822,N_41368,N_41656);
xor U46823 (N_46823,N_44670,N_44938);
or U46824 (N_46824,N_42999,N_40495);
nor U46825 (N_46825,N_40681,N_43381);
nand U46826 (N_46826,N_41509,N_42292);
or U46827 (N_46827,N_44728,N_43235);
nor U46828 (N_46828,N_40306,N_42342);
nor U46829 (N_46829,N_41901,N_40018);
nor U46830 (N_46830,N_44097,N_40005);
xor U46831 (N_46831,N_40225,N_42040);
nor U46832 (N_46832,N_41451,N_41447);
nand U46833 (N_46833,N_43920,N_41686);
or U46834 (N_46834,N_42762,N_43590);
xnor U46835 (N_46835,N_43097,N_43406);
xnor U46836 (N_46836,N_40567,N_41507);
xnor U46837 (N_46837,N_40603,N_40201);
or U46838 (N_46838,N_44822,N_42633);
nor U46839 (N_46839,N_44145,N_42448);
xor U46840 (N_46840,N_40961,N_43230);
nand U46841 (N_46841,N_41652,N_42453);
nand U46842 (N_46842,N_44915,N_41634);
nor U46843 (N_46843,N_44648,N_42541);
nand U46844 (N_46844,N_40761,N_41777);
and U46845 (N_46845,N_44745,N_43234);
and U46846 (N_46846,N_41418,N_40605);
and U46847 (N_46847,N_40235,N_43033);
xnor U46848 (N_46848,N_42881,N_41939);
and U46849 (N_46849,N_40400,N_43787);
or U46850 (N_46850,N_42852,N_41774);
xor U46851 (N_46851,N_42398,N_42339);
nand U46852 (N_46852,N_43915,N_42880);
and U46853 (N_46853,N_41496,N_41711);
nor U46854 (N_46854,N_43337,N_42049);
xnor U46855 (N_46855,N_40974,N_42189);
and U46856 (N_46856,N_40590,N_40875);
nand U46857 (N_46857,N_41152,N_41714);
nand U46858 (N_46858,N_41060,N_44840);
nand U46859 (N_46859,N_44898,N_40935);
nand U46860 (N_46860,N_40724,N_43367);
and U46861 (N_46861,N_42672,N_40384);
or U46862 (N_46862,N_43563,N_41423);
and U46863 (N_46863,N_40345,N_41221);
nor U46864 (N_46864,N_40194,N_43544);
nand U46865 (N_46865,N_41412,N_41742);
nand U46866 (N_46866,N_42677,N_44211);
nand U46867 (N_46867,N_43717,N_40045);
xnor U46868 (N_46868,N_40094,N_41719);
nor U46869 (N_46869,N_43648,N_43959);
xnor U46870 (N_46870,N_41112,N_42480);
and U46871 (N_46871,N_40557,N_42209);
nand U46872 (N_46872,N_43271,N_42030);
or U46873 (N_46873,N_44387,N_41123);
and U46874 (N_46874,N_43050,N_43705);
or U46875 (N_46875,N_42178,N_43763);
nand U46876 (N_46876,N_42687,N_44265);
or U46877 (N_46877,N_40733,N_44146);
and U46878 (N_46878,N_41083,N_43535);
and U46879 (N_46879,N_42971,N_43935);
nor U46880 (N_46880,N_44667,N_44255);
or U46881 (N_46881,N_44354,N_43839);
nor U46882 (N_46882,N_43194,N_43424);
nor U46883 (N_46883,N_41557,N_40309);
or U46884 (N_46884,N_42911,N_41010);
or U46885 (N_46885,N_44786,N_43332);
nand U46886 (N_46886,N_43712,N_42389);
xnor U46887 (N_46887,N_40588,N_41580);
and U46888 (N_46888,N_40329,N_40678);
nor U46889 (N_46889,N_43994,N_43506);
and U46890 (N_46890,N_40691,N_41143);
and U46891 (N_46891,N_43697,N_43975);
nand U46892 (N_46892,N_42530,N_40853);
nor U46893 (N_46893,N_42220,N_44845);
and U46894 (N_46894,N_42641,N_40316);
or U46895 (N_46895,N_40718,N_43285);
and U46896 (N_46896,N_40856,N_43439);
xnor U46897 (N_46897,N_42386,N_43178);
or U46898 (N_46898,N_42493,N_44645);
xor U46899 (N_46899,N_42270,N_41127);
or U46900 (N_46900,N_42555,N_42966);
or U46901 (N_46901,N_41981,N_40604);
xor U46902 (N_46902,N_41385,N_40207);
nor U46903 (N_46903,N_41508,N_43058);
nand U46904 (N_46904,N_40895,N_41684);
or U46905 (N_46905,N_40732,N_40924);
nand U46906 (N_46906,N_42190,N_44361);
nand U46907 (N_46907,N_42666,N_42227);
and U46908 (N_46908,N_44895,N_42561);
or U46909 (N_46909,N_44128,N_43382);
nand U46910 (N_46910,N_42581,N_42723);
and U46911 (N_46911,N_44006,N_40234);
or U46912 (N_46912,N_40331,N_41246);
nor U46913 (N_46913,N_40570,N_41978);
nand U46914 (N_46914,N_43352,N_40941);
nand U46915 (N_46915,N_44585,N_44675);
and U46916 (N_46916,N_40777,N_41821);
xnor U46917 (N_46917,N_41059,N_44012);
nor U46918 (N_46918,N_43881,N_44698);
and U46919 (N_46919,N_44888,N_44318);
xor U46920 (N_46920,N_43000,N_41444);
xnor U46921 (N_46921,N_41325,N_40635);
nor U46922 (N_46922,N_44312,N_42459);
xnor U46923 (N_46923,N_44653,N_42154);
and U46924 (N_46924,N_40748,N_44546);
nand U46925 (N_46925,N_44482,N_43892);
xnor U46926 (N_46926,N_40383,N_44282);
or U46927 (N_46927,N_41927,N_40375);
or U46928 (N_46928,N_44202,N_43880);
and U46929 (N_46929,N_43679,N_44964);
xnor U46930 (N_46930,N_41134,N_41379);
and U46931 (N_46931,N_41782,N_44032);
or U46932 (N_46932,N_42646,N_41872);
nor U46933 (N_46933,N_44381,N_44245);
nand U46934 (N_46934,N_42671,N_42425);
or U46935 (N_46935,N_44093,N_43028);
nand U46936 (N_46936,N_41023,N_43505);
and U46937 (N_46937,N_41827,N_41395);
xor U46938 (N_46938,N_42614,N_44587);
nor U46939 (N_46939,N_44851,N_44823);
nor U46940 (N_46940,N_43268,N_44442);
nand U46941 (N_46941,N_42706,N_44001);
or U46942 (N_46942,N_42113,N_41793);
xnor U46943 (N_46943,N_41156,N_43429);
or U46944 (N_46944,N_43253,N_44084);
nor U46945 (N_46945,N_42111,N_43967);
and U46946 (N_46946,N_43344,N_43690);
and U46947 (N_46947,N_40918,N_42578);
nand U46948 (N_46948,N_41161,N_41133);
or U46949 (N_46949,N_43549,N_43973);
nor U46950 (N_46950,N_40619,N_42940);
xnor U46951 (N_46951,N_41869,N_40022);
nor U46952 (N_46952,N_41442,N_42452);
nor U46953 (N_46953,N_40554,N_44382);
and U46954 (N_46954,N_40573,N_40606);
and U46955 (N_46955,N_40433,N_42764);
nand U46956 (N_46956,N_42819,N_44297);
or U46957 (N_46957,N_44059,N_42905);
and U46958 (N_46958,N_43532,N_42925);
and U46959 (N_46959,N_41422,N_44990);
or U46960 (N_46960,N_43812,N_40260);
or U46961 (N_46961,N_42707,N_43061);
xor U46962 (N_46962,N_42018,N_41799);
or U46963 (N_46963,N_42885,N_43980);
xor U46964 (N_46964,N_42171,N_40489);
nand U46965 (N_46965,N_43372,N_41941);
nor U46966 (N_46966,N_42582,N_44881);
or U46967 (N_46967,N_41970,N_43341);
nor U46968 (N_46968,N_43436,N_41775);
nand U46969 (N_46969,N_43997,N_42297);
and U46970 (N_46970,N_41419,N_42725);
xnor U46971 (N_46971,N_44130,N_43037);
nand U46972 (N_46972,N_42177,N_40892);
nand U46973 (N_46973,N_43805,N_40264);
nand U46974 (N_46974,N_44184,N_44016);
or U46975 (N_46975,N_44517,N_43932);
or U46976 (N_46976,N_40987,N_44090);
nor U46977 (N_46977,N_44370,N_44794);
and U46978 (N_46978,N_44669,N_43108);
and U46979 (N_46979,N_40854,N_40232);
nor U46980 (N_46980,N_41662,N_43146);
or U46981 (N_46981,N_42591,N_40512);
nor U46982 (N_46982,N_44458,N_41075);
and U46983 (N_46983,N_41949,N_42731);
xnor U46984 (N_46984,N_41983,N_42185);
nand U46985 (N_46985,N_44804,N_44422);
and U46986 (N_46986,N_41139,N_44882);
nor U46987 (N_46987,N_41528,N_43473);
nor U46988 (N_46988,N_43297,N_43884);
or U46989 (N_46989,N_40274,N_40469);
nand U46990 (N_46990,N_40223,N_42997);
nor U46991 (N_46991,N_42822,N_43974);
nor U46992 (N_46992,N_42599,N_40715);
xor U46993 (N_46993,N_42982,N_40468);
nand U46994 (N_46994,N_41013,N_40044);
or U46995 (N_46995,N_44054,N_41729);
xor U46996 (N_46996,N_41483,N_42638);
nor U46997 (N_46997,N_42609,N_41912);
and U46998 (N_46998,N_40251,N_43408);
nand U46999 (N_46999,N_40538,N_43934);
and U47000 (N_47000,N_40085,N_42144);
nand U47001 (N_47001,N_43874,N_44263);
or U47002 (N_47002,N_40451,N_42291);
nor U47003 (N_47003,N_40682,N_43286);
xor U47004 (N_47004,N_43850,N_40485);
and U47005 (N_47005,N_44435,N_44325);
nor U47006 (N_47006,N_42767,N_44999);
xnor U47007 (N_47007,N_41890,N_41600);
xor U47008 (N_47008,N_43276,N_44856);
nand U47009 (N_47009,N_42787,N_43764);
nor U47010 (N_47010,N_44065,N_43478);
or U47011 (N_47011,N_42802,N_44469);
nor U47012 (N_47012,N_43218,N_41044);
xor U47013 (N_47013,N_40299,N_43860);
and U47014 (N_47014,N_41047,N_41685);
nand U47015 (N_47015,N_44209,N_44398);
xnor U47016 (N_47016,N_44320,N_42749);
nor U47017 (N_47017,N_43504,N_43199);
xnor U47018 (N_47018,N_43790,N_44943);
and U47019 (N_47019,N_40920,N_40443);
xor U47020 (N_47020,N_42321,N_43292);
nand U47021 (N_47021,N_40759,N_44726);
nor U47022 (N_47022,N_42567,N_44647);
xnor U47023 (N_47023,N_41225,N_40010);
nor U47024 (N_47024,N_43680,N_40940);
and U47025 (N_47025,N_44456,N_41905);
nor U47026 (N_47026,N_41203,N_44801);
nor U47027 (N_47027,N_43150,N_42735);
nor U47028 (N_47028,N_40133,N_40556);
nand U47029 (N_47029,N_42627,N_44479);
nand U47030 (N_47030,N_44218,N_40324);
or U47031 (N_47031,N_41863,N_43064);
or U47032 (N_47032,N_42850,N_41106);
nor U47033 (N_47033,N_41322,N_42072);
nor U47034 (N_47034,N_42557,N_40114);
nand U47035 (N_47035,N_43350,N_41953);
nor U47036 (N_47036,N_40620,N_42686);
nor U47037 (N_47037,N_40753,N_43834);
nand U47038 (N_47038,N_43629,N_41411);
nor U47039 (N_47039,N_42099,N_41068);
nand U47040 (N_47040,N_40243,N_44111);
xnor U47041 (N_47041,N_42460,N_42087);
and U47042 (N_47042,N_41532,N_41590);
xnor U47043 (N_47043,N_42968,N_43929);
and U47044 (N_47044,N_40116,N_43476);
nand U47045 (N_47045,N_43628,N_41413);
xnor U47046 (N_47046,N_42130,N_42244);
nand U47047 (N_47047,N_44160,N_44292);
or U47048 (N_47048,N_41072,N_42665);
and U47049 (N_47049,N_42160,N_42034);
xnor U47050 (N_47050,N_43555,N_44072);
xnor U47051 (N_47051,N_43803,N_41111);
or U47052 (N_47052,N_42349,N_42720);
or U47053 (N_47053,N_42949,N_41795);
nor U47054 (N_47054,N_43963,N_40399);
nor U47055 (N_47055,N_43415,N_41323);
and U47056 (N_47056,N_40809,N_40187);
xor U47057 (N_47057,N_43512,N_42832);
nor U47058 (N_47058,N_40217,N_42845);
and U47059 (N_47059,N_41263,N_44216);
or U47060 (N_47060,N_43637,N_44417);
xnor U47061 (N_47061,N_40357,N_43325);
or U47062 (N_47062,N_41749,N_41616);
and U47063 (N_47063,N_43057,N_43747);
nand U47064 (N_47064,N_41454,N_41510);
nor U47065 (N_47065,N_42391,N_41615);
and U47066 (N_47066,N_41734,N_41533);
xnor U47067 (N_47067,N_40276,N_43837);
xnor U47068 (N_47068,N_40638,N_42631);
or U47069 (N_47069,N_44048,N_41555);
xor U47070 (N_47070,N_43328,N_43644);
nand U47071 (N_47071,N_42474,N_41022);
nand U47072 (N_47072,N_44622,N_41536);
nand U47073 (N_47073,N_44652,N_43376);
xor U47074 (N_47074,N_41240,N_44347);
or U47075 (N_47075,N_43206,N_42606);
nor U47076 (N_47076,N_44112,N_44632);
or U47077 (N_47077,N_41766,N_41080);
and U47078 (N_47078,N_43509,N_41299);
nor U47079 (N_47079,N_44963,N_40519);
xor U47080 (N_47080,N_40464,N_43053);
or U47081 (N_47081,N_43119,N_41124);
and U47082 (N_47082,N_42293,N_44685);
xnor U47083 (N_47083,N_43289,N_42332);
xnor U47084 (N_47084,N_44763,N_44087);
nor U47085 (N_47085,N_41682,N_40540);
or U47086 (N_47086,N_44174,N_43857);
or U47087 (N_47087,N_40392,N_40631);
or U47088 (N_47088,N_43673,N_42258);
nand U47089 (N_47089,N_40403,N_43180);
nand U47090 (N_47090,N_42187,N_41620);
nand U47091 (N_47091,N_42886,N_42893);
xnor U47092 (N_47092,N_41892,N_41037);
and U47093 (N_47093,N_44559,N_42397);
nand U47094 (N_47094,N_43923,N_40740);
xor U47095 (N_47095,N_44153,N_42203);
nor U47096 (N_47096,N_43633,N_43040);
and U47097 (N_47097,N_43829,N_43826);
nand U47098 (N_47098,N_42208,N_40779);
nor U47099 (N_47099,N_40956,N_42298);
nor U47100 (N_47100,N_41632,N_43446);
and U47101 (N_47101,N_40738,N_43173);
nand U47102 (N_47102,N_43222,N_42942);
nand U47103 (N_47103,N_43605,N_40996);
or U47104 (N_47104,N_42503,N_43708);
and U47105 (N_47105,N_41427,N_40209);
nor U47106 (N_47106,N_43578,N_40028);
xnor U47107 (N_47107,N_41756,N_41895);
nand U47108 (N_47108,N_40125,N_42689);
nand U47109 (N_47109,N_44175,N_40401);
nand U47110 (N_47110,N_42509,N_40092);
nand U47111 (N_47111,N_43247,N_41315);
nand U47112 (N_47112,N_44277,N_42680);
xnor U47113 (N_47113,N_40119,N_40042);
nor U47114 (N_47114,N_40476,N_43402);
or U47115 (N_47115,N_40189,N_42367);
and U47116 (N_47116,N_40645,N_43465);
and U47117 (N_47117,N_40578,N_40248);
or U47118 (N_47118,N_42831,N_40690);
nand U47119 (N_47119,N_44961,N_42322);
and U47120 (N_47120,N_43329,N_44257);
or U47121 (N_47121,N_44586,N_42073);
and U47122 (N_47122,N_41382,N_40929);
nor U47123 (N_47123,N_40766,N_41356);
and U47124 (N_47124,N_42584,N_41321);
or U47125 (N_47125,N_42674,N_44393);
nor U47126 (N_47126,N_42430,N_44886);
and U47127 (N_47127,N_44198,N_41241);
nand U47128 (N_47128,N_42972,N_44600);
and U47129 (N_47129,N_41380,N_40290);
nand U47130 (N_47130,N_44973,N_41716);
or U47131 (N_47131,N_42237,N_40760);
and U47132 (N_47132,N_41712,N_40672);
nand U47133 (N_47133,N_43083,N_41070);
nor U47134 (N_47134,N_40755,N_42992);
and U47135 (N_47135,N_41611,N_40628);
or U47136 (N_47136,N_43646,N_44824);
or U47137 (N_47137,N_41126,N_43287);
nor U47138 (N_47138,N_43516,N_41266);
nor U47139 (N_47139,N_42520,N_42851);
nand U47140 (N_47140,N_43956,N_42147);
and U47141 (N_47141,N_40453,N_40311);
nand U47142 (N_47142,N_41589,N_44124);
nand U47143 (N_47143,N_44668,N_41462);
nand U47144 (N_47144,N_40308,N_41584);
nand U47145 (N_47145,N_43781,N_44532);
or U47146 (N_47146,N_43421,N_40350);
nand U47147 (N_47147,N_41529,N_40806);
nor U47148 (N_47148,N_44905,N_42953);
and U47149 (N_47149,N_44403,N_41305);
and U47150 (N_47150,N_43327,N_40247);
xor U47151 (N_47151,N_42042,N_41482);
nand U47152 (N_47152,N_44682,N_42738);
nor U47153 (N_47153,N_43059,N_41999);
and U47154 (N_47154,N_43355,N_41754);
nor U47155 (N_47155,N_43922,N_43464);
xnor U47156 (N_47156,N_43737,N_44391);
xor U47157 (N_47157,N_40339,N_41644);
xnor U47158 (N_47158,N_43324,N_43791);
nor U47159 (N_47159,N_41268,N_44014);
or U47160 (N_47160,N_40030,N_44593);
xnor U47161 (N_47161,N_40069,N_42068);
nand U47162 (N_47162,N_43862,N_40560);
xor U47163 (N_47163,N_44166,N_42242);
and U47164 (N_47164,N_42929,N_42539);
xnor U47165 (N_47165,N_43095,N_43291);
or U47166 (N_47166,N_43602,N_44739);
xnor U47167 (N_47167,N_44899,N_40817);
or U47168 (N_47168,N_40983,N_43930);
nand U47169 (N_47169,N_41101,N_40218);
or U47170 (N_47170,N_44718,N_40963);
or U47171 (N_47171,N_42986,N_43002);
nand U47172 (N_47172,N_42478,N_43479);
nor U47173 (N_47173,N_44960,N_42409);
or U47174 (N_47174,N_43883,N_43351);
xnor U47175 (N_47175,N_43817,N_40348);
xor U47176 (N_47176,N_44020,N_40582);
nor U47177 (N_47177,N_43156,N_40279);
nand U47178 (N_47178,N_41018,N_44860);
or U47179 (N_47179,N_41848,N_40841);
nor U47180 (N_47180,N_41875,N_42023);
xnor U47181 (N_47181,N_41485,N_43531);
nor U47182 (N_47182,N_43632,N_41463);
nand U47183 (N_47183,N_40108,N_44327);
and U47184 (N_47184,N_41676,N_42616);
nand U47185 (N_47185,N_44428,N_43354);
nand U47186 (N_47186,N_44266,N_41992);
and U47187 (N_47187,N_43757,N_41027);
xor U47188 (N_47188,N_41878,N_40867);
nand U47189 (N_47189,N_40049,N_44305);
nand U47190 (N_47190,N_41840,N_42930);
and U47191 (N_47191,N_44848,N_40728);
nand U47192 (N_47192,N_41819,N_43346);
and U47193 (N_47193,N_42694,N_42438);
or U47194 (N_47194,N_43186,N_43443);
xor U47195 (N_47195,N_41871,N_41335);
nand U47196 (N_47196,N_42830,N_41376);
nand U47197 (N_47197,N_44790,N_43137);
xnor U47198 (N_47198,N_43606,N_43172);
xnor U47199 (N_47199,N_42330,N_42739);
and U47200 (N_47200,N_40481,N_42457);
or U47201 (N_47201,N_44411,N_40436);
xor U47202 (N_47202,N_40388,N_42517);
nand U47203 (N_47203,N_44508,N_42781);
nor U47204 (N_47204,N_41943,N_44490);
and U47205 (N_47205,N_42673,N_40386);
xor U47206 (N_47206,N_40038,N_43093);
or U47207 (N_47207,N_41849,N_43495);
nor U47208 (N_47208,N_43405,N_40615);
nor U47209 (N_47209,N_43904,N_44911);
nor U47210 (N_47210,N_41056,N_43538);
xor U47211 (N_47211,N_43668,N_44431);
nand U47212 (N_47212,N_42048,N_40832);
nand U47213 (N_47213,N_43378,N_40347);
nor U47214 (N_47214,N_42692,N_40865);
xor U47215 (N_47215,N_41629,N_43197);
nor U47216 (N_47216,N_41136,N_44228);
and U47217 (N_47217,N_42628,N_42152);
and U47218 (N_47218,N_41311,N_41164);
nor U47219 (N_47219,N_40332,N_42328);
or U47220 (N_47220,N_43706,N_41746);
nor U47221 (N_47221,N_43529,N_43866);
nand U47222 (N_47222,N_40361,N_42060);
or U47223 (N_47223,N_41559,N_40527);
nand U47224 (N_47224,N_43527,N_42518);
nor U47225 (N_47225,N_44396,N_44306);
nor U47226 (N_47226,N_40379,N_41400);
xnor U47227 (N_47227,N_43779,N_44346);
nand U47228 (N_47228,N_43048,N_44996);
and U47229 (N_47229,N_43207,N_43460);
nand U47230 (N_47230,N_43009,N_42449);
nor U47231 (N_47231,N_40633,N_43735);
xnor U47232 (N_47232,N_41838,N_42118);
and U47233 (N_47233,N_41917,N_41552);
or U47234 (N_47234,N_40818,N_40151);
and U47235 (N_47235,N_43484,N_43423);
xor U47236 (N_47236,N_44705,N_43542);
xor U47237 (N_47237,N_44676,N_43312);
and U47238 (N_47238,N_43647,N_41002);
and U47239 (N_47239,N_44744,N_40751);
or U47240 (N_47240,N_43398,N_43766);
nor U47241 (N_47241,N_44948,N_43211);
or U47242 (N_47242,N_40882,N_44067);
and U47243 (N_47243,N_42066,N_40294);
nand U47244 (N_47244,N_41378,N_44034);
and U47245 (N_47245,N_40427,N_40494);
and U47246 (N_47246,N_43876,N_42751);
or U47247 (N_47247,N_40154,N_44784);
and U47248 (N_47248,N_40450,N_42001);
and U47249 (N_47249,N_44535,N_42564);
and U47250 (N_47250,N_44834,N_44880);
and U47251 (N_47251,N_41103,N_43393);
nand U47252 (N_47252,N_40389,N_42794);
xor U47253 (N_47253,N_42271,N_44612);
nor U47254 (N_47254,N_41657,N_43231);
and U47255 (N_47255,N_44323,N_43853);
xor U47256 (N_47256,N_43307,N_42976);
or U47257 (N_47257,N_43019,N_43522);
nor U47258 (N_47258,N_40640,N_41338);
or U47259 (N_47259,N_42427,N_44247);
or U47260 (N_47260,N_44238,N_40368);
nor U47261 (N_47261,N_42173,N_44119);
nor U47262 (N_47262,N_43638,N_43780);
nand U47263 (N_47263,N_44624,N_41403);
nand U47264 (N_47264,N_40585,N_42816);
and U47265 (N_47265,N_40800,N_44913);
nor U47266 (N_47266,N_44061,N_43788);
or U47267 (N_47267,N_43552,N_41474);
xor U47268 (N_47268,N_40480,N_41699);
nand U47269 (N_47269,N_42937,N_43843);
and U47270 (N_47270,N_40958,N_44122);
nand U47271 (N_47271,N_42465,N_42044);
nor U47272 (N_47272,N_42636,N_43298);
and U47273 (N_47273,N_42282,N_44033);
or U47274 (N_47274,N_42978,N_42215);
xnor U47275 (N_47275,N_40944,N_41919);
or U47276 (N_47276,N_44440,N_40076);
or U47277 (N_47277,N_41967,N_42575);
nor U47278 (N_47278,N_40122,N_43249);
or U47279 (N_47279,N_40084,N_43170);
xor U47280 (N_47280,N_44365,N_43005);
and U47281 (N_47281,N_43308,N_40340);
or U47282 (N_47282,N_43049,N_43007);
xnor U47283 (N_47283,N_43688,N_40059);
nor U47284 (N_47284,N_43317,N_44689);
xnor U47285 (N_47285,N_43483,N_40158);
nand U47286 (N_47286,N_42865,N_43030);
xor U47287 (N_47287,N_40344,N_42605);
and U47288 (N_47288,N_44171,N_40721);
and U47289 (N_47289,N_41004,N_43548);
and U47290 (N_47290,N_42772,N_41723);
or U47291 (N_47291,N_42462,N_42047);
or U47292 (N_47292,N_41899,N_42785);
nand U47293 (N_47293,N_44513,N_40016);
or U47294 (N_47294,N_40729,N_43112);
xnor U47295 (N_47295,N_42926,N_44527);
nand U47296 (N_47296,N_40536,N_41720);
and U47297 (N_47297,N_43537,N_44248);
and U47298 (N_47298,N_43749,N_44144);
nand U47299 (N_47299,N_41658,N_41801);
or U47300 (N_47300,N_41730,N_44770);
or U47301 (N_47301,N_42934,N_42902);
or U47302 (N_47302,N_43596,N_44471);
and U47303 (N_47303,N_41262,N_42315);
nor U47304 (N_47304,N_44825,N_41414);
nor U47305 (N_47305,N_44308,N_40884);
xor U47306 (N_47306,N_40390,N_42421);
xnor U47307 (N_47307,N_44703,N_43326);
xnor U47308 (N_47308,N_43442,N_40539);
xnor U47309 (N_47309,N_44644,N_42412);
nor U47310 (N_47310,N_40525,N_43392);
or U47311 (N_47311,N_42316,N_40250);
nor U47312 (N_47312,N_40838,N_40942);
and U47313 (N_47313,N_43640,N_41151);
and U47314 (N_47314,N_44437,N_41200);
xnor U47315 (N_47315,N_41807,N_40137);
xnor U47316 (N_47316,N_40824,N_44309);
or U47317 (N_47317,N_41276,N_44439);
and U47318 (N_47318,N_44591,N_43306);
nor U47319 (N_47319,N_44830,N_41301);
xnor U47320 (N_47320,N_44660,N_42967);
nand U47321 (N_47321,N_44280,N_43806);
xnor U47322 (N_47322,N_41672,N_40723);
and U47323 (N_47323,N_40104,N_43301);
nor U47324 (N_47324,N_43660,N_41313);
or U47325 (N_47325,N_41312,N_41252);
or U47326 (N_47326,N_40211,N_44838);
and U47327 (N_47327,N_42026,N_41923);
and U47328 (N_47328,N_41351,N_43514);
nor U47329 (N_47329,N_43411,N_41193);
or U47330 (N_47330,N_41019,N_40023);
xnor U47331 (N_47331,N_42337,N_40835);
and U47332 (N_47332,N_43385,N_43770);
xor U47333 (N_47333,N_43493,N_43752);
nand U47334 (N_47334,N_42954,N_40475);
xor U47335 (N_47335,N_44287,N_42891);
nand U47336 (N_47336,N_42512,N_43031);
xor U47337 (N_47337,N_40442,N_43727);
nor U47338 (N_47338,N_44333,N_41607);
or U47339 (N_47339,N_42703,N_43909);
or U47340 (N_47340,N_44813,N_44877);
nor U47341 (N_47341,N_41168,N_44321);
nor U47342 (N_47342,N_40852,N_44549);
and U47343 (N_47343,N_44028,N_43288);
nor U47344 (N_47344,N_40106,N_42050);
or U47345 (N_47345,N_43149,N_41163);
nor U47346 (N_47346,N_44429,N_43016);
and U47347 (N_47347,N_41926,N_42844);
xor U47348 (N_47348,N_41638,N_41523);
nor U47349 (N_47349,N_41566,N_44614);
nand U47350 (N_47350,N_40067,N_42247);
xnor U47351 (N_47351,N_44966,N_44221);
nor U47352 (N_47352,N_43038,N_44455);
and U47353 (N_47353,N_44650,N_42265);
nand U47354 (N_47354,N_40938,N_41231);
nand U47355 (N_47355,N_43089,N_40435);
and U47356 (N_47356,N_42149,N_43622);
xor U47357 (N_47357,N_41081,N_44385);
and U47358 (N_47358,N_43742,N_43741);
and U47359 (N_47359,N_41649,N_44972);
or U47360 (N_47360,N_42847,N_40333);
and U47361 (N_47361,N_44887,N_44478);
xnor U47362 (N_47362,N_43118,N_43580);
or U47363 (N_47363,N_41703,N_42002);
nand U47364 (N_47364,N_43106,N_42375);
and U47365 (N_47365,N_44552,N_41341);
and U47366 (N_47366,N_41900,N_41353);
nand U47367 (N_47367,N_40591,N_42007);
and U47368 (N_47368,N_41389,N_44817);
and U47369 (N_47369,N_42746,N_41971);
nand U47370 (N_47370,N_40878,N_44753);
xor U47371 (N_47371,N_41343,N_44193);
xnor U47372 (N_47372,N_40298,N_44444);
nand U47373 (N_47373,N_43778,N_44474);
nand U47374 (N_47374,N_40529,N_40661);
or U47375 (N_47375,N_44089,N_40175);
xor U47376 (N_47376,N_44039,N_44879);
or U47377 (N_47377,N_44942,N_41274);
and U47378 (N_47378,N_43642,N_44820);
or U47379 (N_47379,N_43365,N_40781);
nand U47380 (N_47380,N_40876,N_42429);
and U47381 (N_47381,N_42959,N_40358);
xnor U47382 (N_47382,N_42974,N_41190);
and U47383 (N_47383,N_41183,N_41858);
nand U47384 (N_47384,N_41914,N_44520);
or U47385 (N_47385,N_41988,N_40579);
xor U47386 (N_47386,N_40222,N_44019);
or U47387 (N_47387,N_42059,N_44750);
nor U47388 (N_47388,N_44693,N_42120);
or U47389 (N_47389,N_41708,N_40141);
nand U47390 (N_47390,N_41171,N_40233);
or U47391 (N_47391,N_40816,N_41844);
nor U47392 (N_47392,N_43374,N_41767);
and U47393 (N_47393,N_44275,N_44924);
or U47394 (N_47394,N_41053,N_44045);
and U47395 (N_47395,N_40477,N_44617);
nand U47396 (N_47396,N_40885,N_44249);
or U47397 (N_47397,N_42824,N_42726);
nor U47398 (N_47398,N_42097,N_44289);
nor U47399 (N_47399,N_43015,N_42511);
or U47400 (N_47400,N_44909,N_41224);
nand U47401 (N_47401,N_44778,N_42476);
nand U47402 (N_47402,N_44304,N_40414);
nand U47403 (N_47403,N_40101,N_42813);
nand U47404 (N_47404,N_40017,N_41234);
nand U47405 (N_47405,N_40168,N_43523);
or U47406 (N_47406,N_40812,N_43953);
and U47407 (N_47407,N_44985,N_41166);
xnor U47408 (N_47408,N_42695,N_44839);
xor U47409 (N_47409,N_42870,N_44781);
xnor U47410 (N_47410,N_42667,N_43087);
nand U47411 (N_47411,N_41542,N_42803);
nor U47412 (N_47412,N_40371,N_43348);
nand U47413 (N_47413,N_40415,N_42313);
nor U47414 (N_47414,N_42340,N_40687);
nor U47415 (N_47415,N_41342,N_41218);
nand U47416 (N_47416,N_41398,N_42071);
nor U47417 (N_47417,N_42304,N_41813);
xor U47418 (N_47418,N_43136,N_42854);
xnor U47419 (N_47419,N_44138,N_40278);
xor U47420 (N_47420,N_42647,N_44525);
xnor U47421 (N_47421,N_42064,N_44081);
nor U47422 (N_47422,N_41429,N_44454);
and U47423 (N_47423,N_41643,N_42241);
and U47424 (N_47424,N_40146,N_44070);
nor U47425 (N_47425,N_42336,N_43458);
and U47426 (N_47426,N_43924,N_40762);
xnor U47427 (N_47427,N_41861,N_44890);
xor U47428 (N_47428,N_42121,N_43238);
nor U47429 (N_47429,N_44798,N_44252);
or U47430 (N_47430,N_40859,N_40288);
xor U47431 (N_47431,N_42748,N_44140);
nand U47432 (N_47432,N_41433,N_42086);
nor U47433 (N_47433,N_41373,N_43233);
xnor U47434 (N_47434,N_40599,N_42019);
nor U47435 (N_47435,N_40155,N_42303);
or U47436 (N_47436,N_41816,N_43716);
or U47437 (N_47437,N_42716,N_40300);
nand U47438 (N_47438,N_42174,N_40024);
nand U47439 (N_47439,N_42166,N_44562);
and U47440 (N_47440,N_43321,N_44777);
xnor U47441 (N_47441,N_40113,N_40563);
or U47442 (N_47442,N_40445,N_40569);
and U47443 (N_47443,N_40479,N_43562);
and U47444 (N_47444,N_40689,N_41177);
nor U47445 (N_47445,N_41565,N_41721);
or U47446 (N_47446,N_44874,N_43682);
xnor U47447 (N_47447,N_42676,N_42766);
or U47448 (N_47448,N_40994,N_41837);
and U47449 (N_47449,N_41091,N_40694);
nand U47450 (N_47450,N_43754,N_42299);
and U47451 (N_47451,N_44747,N_40526);
nand U47452 (N_47452,N_43054,N_43702);
xnor U47453 (N_47453,N_42604,N_44725);
xnor U47454 (N_47454,N_42842,N_41515);
nand U47455 (N_47455,N_43677,N_41015);
xnor U47456 (N_47456,N_44447,N_41834);
nor U47457 (N_47457,N_41808,N_40618);
and U47458 (N_47458,N_44949,N_40797);
nor U47459 (N_47459,N_42568,N_42988);
and U47460 (N_47460,N_42810,N_41969);
or U47461 (N_47461,N_40438,N_41082);
or U47462 (N_47462,N_42600,N_42559);
xor U47463 (N_47463,N_40959,N_43187);
or U47464 (N_47464,N_41810,N_40323);
nand U47465 (N_47465,N_44433,N_42051);
nor U47466 (N_47466,N_43873,N_42979);
nor U47467 (N_47467,N_43898,N_41364);
nor U47468 (N_47468,N_44344,N_41867);
nand U47469 (N_47469,N_43144,N_44723);
xor U47470 (N_47470,N_43140,N_41432);
xor U47471 (N_47471,N_44463,N_41745);
nor U47472 (N_47472,N_41232,N_43991);
xor U47473 (N_47473,N_40009,N_43096);
xnor U47474 (N_47474,N_44858,N_42006);
or U47475 (N_47475,N_41147,N_44837);
nor U47476 (N_47476,N_43127,N_43027);
xnor U47477 (N_47477,N_40685,N_40301);
nor U47478 (N_47478,N_41149,N_44294);
or U47479 (N_47479,N_40317,N_44754);
nor U47480 (N_47480,N_44947,N_42861);
or U47481 (N_47481,N_43491,N_40674);
nand U47482 (N_47482,N_42863,N_42109);
nor U47483 (N_47483,N_41519,N_42233);
or U47484 (N_47484,N_41689,N_42319);
and U47485 (N_47485,N_44420,N_41760);
nor U47486 (N_47486,N_42082,N_41713);
and U47487 (N_47487,N_44100,N_43213);
xnor U47488 (N_47488,N_40600,N_44018);
nor U47489 (N_47489,N_41660,N_42240);
xnor U47490 (N_47490,N_41950,N_44022);
or U47491 (N_47491,N_41273,N_41887);
or U47492 (N_47492,N_41757,N_40077);
nand U47493 (N_47493,N_43293,N_43217);
xnor U47494 (N_47494,N_42574,N_43842);
and U47495 (N_47495,N_42345,N_42554);
and U47496 (N_47496,N_43115,N_41850);
xnor U47497 (N_47497,N_40322,N_42385);
nand U47498 (N_47498,N_43818,N_43729);
or U47499 (N_47499,N_42326,N_44311);
nand U47500 (N_47500,N_42825,N_42253);
nand U47501 (N_47501,N_41319,N_44822);
nand U47502 (N_47502,N_44847,N_43996);
and U47503 (N_47503,N_40259,N_42397);
xnor U47504 (N_47504,N_40501,N_41454);
nand U47505 (N_47505,N_40197,N_44206);
nor U47506 (N_47506,N_40880,N_40252);
or U47507 (N_47507,N_42406,N_42966);
nand U47508 (N_47508,N_43273,N_41006);
xor U47509 (N_47509,N_44552,N_42653);
xor U47510 (N_47510,N_44460,N_41747);
or U47511 (N_47511,N_40308,N_44902);
and U47512 (N_47512,N_43461,N_41831);
xor U47513 (N_47513,N_41616,N_44402);
or U47514 (N_47514,N_43087,N_41708);
nand U47515 (N_47515,N_43057,N_40191);
nand U47516 (N_47516,N_41404,N_40355);
xnor U47517 (N_47517,N_41480,N_40615);
xor U47518 (N_47518,N_40743,N_40756);
nor U47519 (N_47519,N_41190,N_44503);
xnor U47520 (N_47520,N_44641,N_44716);
nor U47521 (N_47521,N_40583,N_44281);
nor U47522 (N_47522,N_43696,N_42686);
nor U47523 (N_47523,N_41482,N_44834);
xor U47524 (N_47524,N_44658,N_44528);
nor U47525 (N_47525,N_43005,N_43115);
and U47526 (N_47526,N_44735,N_41455);
or U47527 (N_47527,N_43985,N_40943);
and U47528 (N_47528,N_44708,N_40760);
and U47529 (N_47529,N_43994,N_44727);
xor U47530 (N_47530,N_43658,N_42766);
nor U47531 (N_47531,N_42189,N_42503);
nand U47532 (N_47532,N_44016,N_41894);
nor U47533 (N_47533,N_41575,N_40075);
xor U47534 (N_47534,N_40236,N_43594);
xnor U47535 (N_47535,N_42316,N_43769);
nor U47536 (N_47536,N_41304,N_43888);
or U47537 (N_47537,N_43459,N_40112);
xnor U47538 (N_47538,N_41062,N_44812);
or U47539 (N_47539,N_43310,N_40206);
and U47540 (N_47540,N_41587,N_42384);
nand U47541 (N_47541,N_41346,N_43761);
xnor U47542 (N_47542,N_43888,N_44924);
and U47543 (N_47543,N_43366,N_40148);
nor U47544 (N_47544,N_43704,N_40023);
xnor U47545 (N_47545,N_41924,N_40949);
nand U47546 (N_47546,N_44496,N_44614);
or U47547 (N_47547,N_42395,N_42243);
nand U47548 (N_47548,N_41878,N_44874);
and U47549 (N_47549,N_40280,N_44698);
xor U47550 (N_47550,N_42698,N_43899);
or U47551 (N_47551,N_40659,N_41300);
or U47552 (N_47552,N_43538,N_42725);
nand U47553 (N_47553,N_40934,N_40543);
and U47554 (N_47554,N_40064,N_42353);
nand U47555 (N_47555,N_42145,N_41615);
xnor U47556 (N_47556,N_44079,N_40488);
and U47557 (N_47557,N_44170,N_41698);
nor U47558 (N_47558,N_44293,N_41676);
nand U47559 (N_47559,N_43951,N_40383);
nand U47560 (N_47560,N_42196,N_41022);
nand U47561 (N_47561,N_43109,N_40610);
and U47562 (N_47562,N_43327,N_43545);
nand U47563 (N_47563,N_42548,N_43606);
xnor U47564 (N_47564,N_44475,N_42374);
or U47565 (N_47565,N_41796,N_43659);
xor U47566 (N_47566,N_42260,N_40009);
nand U47567 (N_47567,N_44893,N_41192);
nor U47568 (N_47568,N_42158,N_41168);
or U47569 (N_47569,N_40778,N_41932);
or U47570 (N_47570,N_43617,N_41871);
xor U47571 (N_47571,N_40533,N_43180);
or U47572 (N_47572,N_44348,N_41412);
nand U47573 (N_47573,N_42076,N_43681);
nand U47574 (N_47574,N_42531,N_44663);
or U47575 (N_47575,N_41942,N_44699);
nand U47576 (N_47576,N_43123,N_42546);
nand U47577 (N_47577,N_42682,N_42831);
nand U47578 (N_47578,N_43059,N_43252);
xor U47579 (N_47579,N_41415,N_43051);
nand U47580 (N_47580,N_41556,N_40876);
nor U47581 (N_47581,N_41154,N_40942);
nand U47582 (N_47582,N_44467,N_43056);
or U47583 (N_47583,N_42404,N_41856);
and U47584 (N_47584,N_42544,N_44397);
and U47585 (N_47585,N_43081,N_41950);
nor U47586 (N_47586,N_42652,N_42315);
nand U47587 (N_47587,N_40788,N_41713);
or U47588 (N_47588,N_44405,N_42833);
xnor U47589 (N_47589,N_41620,N_41887);
xor U47590 (N_47590,N_44654,N_44907);
and U47591 (N_47591,N_40497,N_43316);
or U47592 (N_47592,N_43379,N_43470);
and U47593 (N_47593,N_44557,N_44104);
and U47594 (N_47594,N_40344,N_43302);
or U47595 (N_47595,N_44778,N_44095);
xor U47596 (N_47596,N_41616,N_42619);
nor U47597 (N_47597,N_41017,N_40381);
nand U47598 (N_47598,N_41233,N_40684);
nand U47599 (N_47599,N_40569,N_41534);
and U47600 (N_47600,N_41421,N_40482);
nor U47601 (N_47601,N_40901,N_41477);
or U47602 (N_47602,N_44301,N_41971);
xnor U47603 (N_47603,N_43134,N_40059);
and U47604 (N_47604,N_42862,N_40596);
nand U47605 (N_47605,N_42247,N_44031);
and U47606 (N_47606,N_44766,N_43125);
and U47607 (N_47607,N_44500,N_44895);
xnor U47608 (N_47608,N_41443,N_40050);
and U47609 (N_47609,N_44306,N_43576);
and U47610 (N_47610,N_41203,N_41146);
or U47611 (N_47611,N_42913,N_41778);
or U47612 (N_47612,N_43256,N_43381);
xor U47613 (N_47613,N_41375,N_41021);
nand U47614 (N_47614,N_43492,N_40039);
nor U47615 (N_47615,N_40970,N_43350);
nand U47616 (N_47616,N_44720,N_42603);
xor U47617 (N_47617,N_43510,N_40282);
xor U47618 (N_47618,N_41278,N_43032);
nand U47619 (N_47619,N_42003,N_42718);
or U47620 (N_47620,N_41991,N_42301);
nand U47621 (N_47621,N_44690,N_43524);
nor U47622 (N_47622,N_42191,N_43179);
nand U47623 (N_47623,N_41145,N_41391);
nand U47624 (N_47624,N_44889,N_40283);
or U47625 (N_47625,N_44477,N_44287);
nand U47626 (N_47626,N_40236,N_42546);
nand U47627 (N_47627,N_41637,N_41838);
nand U47628 (N_47628,N_44556,N_42402);
xnor U47629 (N_47629,N_41316,N_41907);
or U47630 (N_47630,N_42716,N_40715);
or U47631 (N_47631,N_40748,N_43913);
nor U47632 (N_47632,N_41299,N_42709);
or U47633 (N_47633,N_42574,N_42862);
xnor U47634 (N_47634,N_43777,N_41320);
or U47635 (N_47635,N_44654,N_40767);
and U47636 (N_47636,N_40377,N_43997);
and U47637 (N_47637,N_41979,N_41017);
nor U47638 (N_47638,N_43107,N_41850);
xor U47639 (N_47639,N_41822,N_44185);
and U47640 (N_47640,N_40247,N_44314);
or U47641 (N_47641,N_44801,N_42545);
and U47642 (N_47642,N_43563,N_42912);
or U47643 (N_47643,N_44846,N_42528);
nand U47644 (N_47644,N_43307,N_42470);
nand U47645 (N_47645,N_42078,N_42922);
nand U47646 (N_47646,N_41288,N_43550);
nor U47647 (N_47647,N_42789,N_43694);
xnor U47648 (N_47648,N_40112,N_43686);
or U47649 (N_47649,N_41622,N_41163);
xor U47650 (N_47650,N_43212,N_40131);
nor U47651 (N_47651,N_44130,N_41362);
xor U47652 (N_47652,N_43855,N_42552);
nor U47653 (N_47653,N_44232,N_40830);
nand U47654 (N_47654,N_40660,N_41139);
nand U47655 (N_47655,N_40847,N_44918);
nor U47656 (N_47656,N_41684,N_40761);
nand U47657 (N_47657,N_41753,N_43657);
nand U47658 (N_47658,N_44135,N_40415);
nand U47659 (N_47659,N_43167,N_41340);
xor U47660 (N_47660,N_40011,N_42704);
nand U47661 (N_47661,N_41939,N_40260);
nand U47662 (N_47662,N_42123,N_44830);
nand U47663 (N_47663,N_44353,N_44456);
nand U47664 (N_47664,N_43684,N_40607);
nor U47665 (N_47665,N_40613,N_41354);
or U47666 (N_47666,N_44929,N_40469);
nand U47667 (N_47667,N_42141,N_43305);
nor U47668 (N_47668,N_43839,N_40996);
nand U47669 (N_47669,N_40511,N_43817);
nand U47670 (N_47670,N_42734,N_44931);
nor U47671 (N_47671,N_44566,N_43052);
or U47672 (N_47672,N_40921,N_40492);
nor U47673 (N_47673,N_41242,N_41456);
xor U47674 (N_47674,N_41571,N_42699);
and U47675 (N_47675,N_43183,N_42001);
xnor U47676 (N_47676,N_40907,N_42757);
nand U47677 (N_47677,N_43607,N_42973);
or U47678 (N_47678,N_40334,N_42651);
xor U47679 (N_47679,N_42012,N_40970);
xnor U47680 (N_47680,N_42246,N_44325);
nor U47681 (N_47681,N_44111,N_44010);
and U47682 (N_47682,N_43585,N_43606);
or U47683 (N_47683,N_42400,N_43023);
nand U47684 (N_47684,N_43471,N_44953);
nand U47685 (N_47685,N_42772,N_44861);
nand U47686 (N_47686,N_42234,N_41170);
xnor U47687 (N_47687,N_42182,N_41014);
and U47688 (N_47688,N_41707,N_44402);
or U47689 (N_47689,N_42300,N_42228);
and U47690 (N_47690,N_40198,N_41593);
nand U47691 (N_47691,N_43664,N_44370);
xor U47692 (N_47692,N_44681,N_42905);
and U47693 (N_47693,N_42062,N_40405);
and U47694 (N_47694,N_42497,N_40321);
nand U47695 (N_47695,N_44978,N_44531);
xor U47696 (N_47696,N_43811,N_40030);
nand U47697 (N_47697,N_41954,N_44992);
nor U47698 (N_47698,N_42998,N_44414);
and U47699 (N_47699,N_40580,N_40327);
and U47700 (N_47700,N_44176,N_41181);
or U47701 (N_47701,N_43133,N_41373);
nor U47702 (N_47702,N_41412,N_44371);
nand U47703 (N_47703,N_42198,N_40047);
or U47704 (N_47704,N_42695,N_40269);
or U47705 (N_47705,N_43231,N_44506);
nor U47706 (N_47706,N_44571,N_43020);
nand U47707 (N_47707,N_41784,N_43436);
xor U47708 (N_47708,N_42768,N_42079);
xor U47709 (N_47709,N_44797,N_40177);
xnor U47710 (N_47710,N_41980,N_43499);
and U47711 (N_47711,N_44815,N_42248);
nand U47712 (N_47712,N_42437,N_43538);
xor U47713 (N_47713,N_40738,N_41633);
nor U47714 (N_47714,N_41667,N_43727);
xor U47715 (N_47715,N_42273,N_44876);
nor U47716 (N_47716,N_40399,N_42264);
nand U47717 (N_47717,N_40414,N_41137);
nand U47718 (N_47718,N_41272,N_42336);
nand U47719 (N_47719,N_43680,N_41091);
and U47720 (N_47720,N_40826,N_44664);
nand U47721 (N_47721,N_41142,N_42443);
nand U47722 (N_47722,N_42715,N_40163);
and U47723 (N_47723,N_44015,N_42125);
xnor U47724 (N_47724,N_40279,N_40356);
and U47725 (N_47725,N_43401,N_40584);
and U47726 (N_47726,N_42038,N_44067);
nor U47727 (N_47727,N_43620,N_40557);
and U47728 (N_47728,N_41417,N_43501);
xnor U47729 (N_47729,N_42812,N_43093);
xnor U47730 (N_47730,N_40093,N_44652);
nand U47731 (N_47731,N_42382,N_43271);
xor U47732 (N_47732,N_41982,N_41329);
nand U47733 (N_47733,N_41696,N_43642);
or U47734 (N_47734,N_40494,N_40963);
nand U47735 (N_47735,N_44183,N_41695);
xnor U47736 (N_47736,N_44620,N_42452);
nand U47737 (N_47737,N_44023,N_42974);
nand U47738 (N_47738,N_43816,N_43964);
or U47739 (N_47739,N_40625,N_41089);
and U47740 (N_47740,N_40147,N_44073);
xnor U47741 (N_47741,N_44761,N_40862);
nand U47742 (N_47742,N_43743,N_43991);
nor U47743 (N_47743,N_44068,N_42317);
or U47744 (N_47744,N_42082,N_42281);
xor U47745 (N_47745,N_42391,N_41955);
and U47746 (N_47746,N_41138,N_43703);
nand U47747 (N_47747,N_44663,N_43141);
and U47748 (N_47748,N_44811,N_43297);
and U47749 (N_47749,N_42957,N_42316);
nor U47750 (N_47750,N_41510,N_44569);
or U47751 (N_47751,N_40911,N_43357);
or U47752 (N_47752,N_40513,N_44643);
or U47753 (N_47753,N_43035,N_43520);
xnor U47754 (N_47754,N_40694,N_40081);
nor U47755 (N_47755,N_42396,N_43874);
and U47756 (N_47756,N_43496,N_44898);
and U47757 (N_47757,N_44461,N_40596);
xor U47758 (N_47758,N_40124,N_42586);
or U47759 (N_47759,N_44612,N_44423);
or U47760 (N_47760,N_43246,N_42947);
and U47761 (N_47761,N_42987,N_42091);
and U47762 (N_47762,N_44131,N_40226);
nor U47763 (N_47763,N_41058,N_43332);
or U47764 (N_47764,N_44510,N_43409);
xnor U47765 (N_47765,N_40171,N_42766);
nor U47766 (N_47766,N_44685,N_43594);
xor U47767 (N_47767,N_42941,N_43524);
and U47768 (N_47768,N_40480,N_42480);
xnor U47769 (N_47769,N_41648,N_41271);
nand U47770 (N_47770,N_40714,N_42800);
nand U47771 (N_47771,N_42434,N_40572);
nand U47772 (N_47772,N_44149,N_42596);
or U47773 (N_47773,N_43839,N_40742);
nand U47774 (N_47774,N_41739,N_40360);
or U47775 (N_47775,N_40273,N_41731);
or U47776 (N_47776,N_43079,N_40477);
xnor U47777 (N_47777,N_42345,N_43396);
or U47778 (N_47778,N_44499,N_42259);
and U47779 (N_47779,N_43440,N_43536);
nand U47780 (N_47780,N_44890,N_44800);
and U47781 (N_47781,N_41203,N_43691);
xor U47782 (N_47782,N_43980,N_44284);
or U47783 (N_47783,N_43061,N_40401);
nor U47784 (N_47784,N_41008,N_43482);
and U47785 (N_47785,N_44698,N_40975);
xor U47786 (N_47786,N_40752,N_44185);
nand U47787 (N_47787,N_44098,N_42345);
or U47788 (N_47788,N_41005,N_44798);
nand U47789 (N_47789,N_40063,N_42171);
nand U47790 (N_47790,N_43717,N_43471);
or U47791 (N_47791,N_44296,N_42483);
nand U47792 (N_47792,N_44590,N_44969);
and U47793 (N_47793,N_40413,N_44148);
nor U47794 (N_47794,N_41070,N_41775);
xor U47795 (N_47795,N_44164,N_40889);
and U47796 (N_47796,N_41042,N_43201);
nand U47797 (N_47797,N_44620,N_43494);
and U47798 (N_47798,N_42962,N_43043);
nor U47799 (N_47799,N_40859,N_43894);
and U47800 (N_47800,N_44388,N_42044);
nor U47801 (N_47801,N_42226,N_41751);
nand U47802 (N_47802,N_44813,N_40193);
xor U47803 (N_47803,N_43418,N_42718);
and U47804 (N_47804,N_43786,N_44684);
nand U47805 (N_47805,N_43341,N_42829);
nand U47806 (N_47806,N_42585,N_43401);
or U47807 (N_47807,N_40504,N_42181);
nand U47808 (N_47808,N_40442,N_40485);
nand U47809 (N_47809,N_44606,N_43514);
or U47810 (N_47810,N_41915,N_41456);
and U47811 (N_47811,N_40860,N_40215);
nor U47812 (N_47812,N_41354,N_40880);
xor U47813 (N_47813,N_42511,N_43602);
nor U47814 (N_47814,N_40204,N_41563);
or U47815 (N_47815,N_42319,N_43201);
nor U47816 (N_47816,N_40086,N_44006);
or U47817 (N_47817,N_43262,N_42877);
and U47818 (N_47818,N_42277,N_42645);
and U47819 (N_47819,N_42191,N_40626);
and U47820 (N_47820,N_42679,N_42280);
or U47821 (N_47821,N_41018,N_44921);
nor U47822 (N_47822,N_43039,N_42371);
xnor U47823 (N_47823,N_40798,N_42282);
nor U47824 (N_47824,N_43142,N_40614);
nand U47825 (N_47825,N_44171,N_44599);
nand U47826 (N_47826,N_41941,N_40145);
nor U47827 (N_47827,N_43607,N_40364);
xor U47828 (N_47828,N_43920,N_41102);
or U47829 (N_47829,N_43455,N_42783);
xor U47830 (N_47830,N_44727,N_42500);
nand U47831 (N_47831,N_42019,N_41872);
xor U47832 (N_47832,N_42407,N_43200);
xnor U47833 (N_47833,N_42411,N_40729);
xnor U47834 (N_47834,N_41850,N_44351);
xnor U47835 (N_47835,N_40087,N_44200);
nand U47836 (N_47836,N_41169,N_44187);
and U47837 (N_47837,N_41129,N_41863);
or U47838 (N_47838,N_40966,N_44683);
nand U47839 (N_47839,N_40682,N_43170);
nor U47840 (N_47840,N_43056,N_42040);
nand U47841 (N_47841,N_41340,N_44529);
and U47842 (N_47842,N_44865,N_44445);
xor U47843 (N_47843,N_43215,N_44815);
or U47844 (N_47844,N_42708,N_43119);
xor U47845 (N_47845,N_41854,N_42834);
and U47846 (N_47846,N_41603,N_44137);
and U47847 (N_47847,N_44514,N_40220);
nor U47848 (N_47848,N_43137,N_40608);
or U47849 (N_47849,N_40109,N_43233);
nand U47850 (N_47850,N_41474,N_42417);
nand U47851 (N_47851,N_42480,N_41574);
nand U47852 (N_47852,N_41552,N_40504);
nor U47853 (N_47853,N_41733,N_44139);
nor U47854 (N_47854,N_44232,N_44353);
nor U47855 (N_47855,N_44752,N_44059);
xnor U47856 (N_47856,N_42912,N_41625);
or U47857 (N_47857,N_43478,N_42346);
nor U47858 (N_47858,N_42597,N_42989);
and U47859 (N_47859,N_44515,N_43152);
or U47860 (N_47860,N_43838,N_44343);
xor U47861 (N_47861,N_41927,N_43066);
nor U47862 (N_47862,N_44092,N_42901);
or U47863 (N_47863,N_43641,N_42196);
and U47864 (N_47864,N_42298,N_43353);
nor U47865 (N_47865,N_40455,N_41693);
xor U47866 (N_47866,N_42034,N_43072);
and U47867 (N_47867,N_40543,N_44292);
and U47868 (N_47868,N_40438,N_44467);
or U47869 (N_47869,N_42766,N_43389);
nor U47870 (N_47870,N_41324,N_40049);
xor U47871 (N_47871,N_42044,N_44124);
nor U47872 (N_47872,N_41918,N_44632);
xor U47873 (N_47873,N_44203,N_42841);
and U47874 (N_47874,N_41536,N_44569);
xnor U47875 (N_47875,N_42550,N_41019);
or U47876 (N_47876,N_42083,N_44555);
and U47877 (N_47877,N_43654,N_40693);
nand U47878 (N_47878,N_43868,N_40182);
xnor U47879 (N_47879,N_42871,N_44271);
nor U47880 (N_47880,N_42661,N_40872);
nor U47881 (N_47881,N_42337,N_42252);
nor U47882 (N_47882,N_42142,N_42704);
xor U47883 (N_47883,N_41241,N_44472);
nand U47884 (N_47884,N_40620,N_44030);
xor U47885 (N_47885,N_42284,N_43626);
or U47886 (N_47886,N_43331,N_42377);
nor U47887 (N_47887,N_43312,N_42321);
nor U47888 (N_47888,N_40866,N_40753);
or U47889 (N_47889,N_43714,N_42962);
and U47890 (N_47890,N_41230,N_44439);
or U47891 (N_47891,N_44094,N_40108);
or U47892 (N_47892,N_42763,N_43027);
nand U47893 (N_47893,N_41200,N_41117);
nor U47894 (N_47894,N_43351,N_44379);
xor U47895 (N_47895,N_40726,N_43428);
nand U47896 (N_47896,N_40690,N_41820);
and U47897 (N_47897,N_43406,N_43776);
nor U47898 (N_47898,N_41930,N_41190);
or U47899 (N_47899,N_43438,N_42032);
nor U47900 (N_47900,N_44196,N_43401);
and U47901 (N_47901,N_42348,N_41960);
nor U47902 (N_47902,N_42605,N_44730);
and U47903 (N_47903,N_44140,N_40281);
nand U47904 (N_47904,N_41313,N_43473);
or U47905 (N_47905,N_44331,N_41782);
and U47906 (N_47906,N_41146,N_42959);
or U47907 (N_47907,N_41905,N_40531);
or U47908 (N_47908,N_44920,N_42234);
nand U47909 (N_47909,N_43823,N_41169);
nand U47910 (N_47910,N_44101,N_40601);
nand U47911 (N_47911,N_42947,N_42786);
and U47912 (N_47912,N_41980,N_42870);
and U47913 (N_47913,N_40296,N_44076);
nand U47914 (N_47914,N_42189,N_44303);
nand U47915 (N_47915,N_44753,N_42407);
nor U47916 (N_47916,N_41484,N_40980);
xnor U47917 (N_47917,N_42412,N_40552);
nand U47918 (N_47918,N_44338,N_41743);
xnor U47919 (N_47919,N_40395,N_43278);
or U47920 (N_47920,N_41857,N_41586);
nor U47921 (N_47921,N_43318,N_44881);
nor U47922 (N_47922,N_41548,N_41617);
and U47923 (N_47923,N_44099,N_40256);
and U47924 (N_47924,N_40398,N_41266);
and U47925 (N_47925,N_42000,N_44869);
nor U47926 (N_47926,N_40046,N_40597);
or U47927 (N_47927,N_42730,N_42668);
xnor U47928 (N_47928,N_42169,N_44124);
or U47929 (N_47929,N_40412,N_40238);
nand U47930 (N_47930,N_41094,N_40505);
or U47931 (N_47931,N_43226,N_44216);
xnor U47932 (N_47932,N_44398,N_41755);
and U47933 (N_47933,N_44611,N_44614);
nand U47934 (N_47934,N_42414,N_42591);
and U47935 (N_47935,N_43929,N_41056);
nor U47936 (N_47936,N_41735,N_42569);
and U47937 (N_47937,N_42786,N_40567);
xor U47938 (N_47938,N_43033,N_41453);
nor U47939 (N_47939,N_43107,N_41416);
and U47940 (N_47940,N_42824,N_41308);
nand U47941 (N_47941,N_43044,N_42879);
xor U47942 (N_47942,N_40075,N_40812);
nor U47943 (N_47943,N_40683,N_42610);
nand U47944 (N_47944,N_43105,N_41319);
and U47945 (N_47945,N_41589,N_43620);
xor U47946 (N_47946,N_44869,N_40901);
nor U47947 (N_47947,N_42599,N_41037);
nand U47948 (N_47948,N_40141,N_44360);
nor U47949 (N_47949,N_43895,N_40562);
or U47950 (N_47950,N_44896,N_43567);
nor U47951 (N_47951,N_43529,N_43261);
nand U47952 (N_47952,N_41271,N_44261);
xor U47953 (N_47953,N_40547,N_40123);
nand U47954 (N_47954,N_41864,N_41354);
and U47955 (N_47955,N_43392,N_40784);
nor U47956 (N_47956,N_42588,N_41997);
or U47957 (N_47957,N_40401,N_44758);
xor U47958 (N_47958,N_41383,N_41231);
nor U47959 (N_47959,N_41968,N_42621);
and U47960 (N_47960,N_43619,N_44015);
and U47961 (N_47961,N_44077,N_43146);
or U47962 (N_47962,N_41152,N_40594);
and U47963 (N_47963,N_44741,N_44115);
or U47964 (N_47964,N_43389,N_42650);
xor U47965 (N_47965,N_40259,N_42803);
or U47966 (N_47966,N_41468,N_42616);
nand U47967 (N_47967,N_42606,N_40504);
xor U47968 (N_47968,N_40069,N_44262);
or U47969 (N_47969,N_40650,N_44967);
nor U47970 (N_47970,N_43714,N_42508);
nor U47971 (N_47971,N_44185,N_42139);
nor U47972 (N_47972,N_42758,N_44511);
or U47973 (N_47973,N_42804,N_40065);
and U47974 (N_47974,N_41795,N_42420);
and U47975 (N_47975,N_41086,N_44630);
nand U47976 (N_47976,N_44125,N_41380);
nor U47977 (N_47977,N_41388,N_41400);
xor U47978 (N_47978,N_42056,N_41252);
nand U47979 (N_47979,N_40902,N_43185);
or U47980 (N_47980,N_41398,N_40000);
and U47981 (N_47981,N_43773,N_42381);
nand U47982 (N_47982,N_40579,N_44899);
xnor U47983 (N_47983,N_41067,N_44040);
nand U47984 (N_47984,N_40705,N_40354);
xnor U47985 (N_47985,N_41242,N_41522);
nor U47986 (N_47986,N_44184,N_42622);
nand U47987 (N_47987,N_44251,N_44690);
nand U47988 (N_47988,N_43457,N_44495);
xnor U47989 (N_47989,N_43938,N_43362);
nand U47990 (N_47990,N_43183,N_41778);
and U47991 (N_47991,N_44837,N_41952);
or U47992 (N_47992,N_41682,N_42657);
or U47993 (N_47993,N_40432,N_41381);
xnor U47994 (N_47994,N_42092,N_41972);
nand U47995 (N_47995,N_44779,N_43118);
or U47996 (N_47996,N_43510,N_43836);
and U47997 (N_47997,N_42982,N_44569);
or U47998 (N_47998,N_41153,N_43282);
nor U47999 (N_47999,N_41457,N_44855);
nand U48000 (N_48000,N_40606,N_41920);
nand U48001 (N_48001,N_42662,N_41257);
and U48002 (N_48002,N_40547,N_41887);
nand U48003 (N_48003,N_40860,N_43080);
xor U48004 (N_48004,N_42792,N_43454);
nor U48005 (N_48005,N_44381,N_40469);
nor U48006 (N_48006,N_44990,N_43195);
nor U48007 (N_48007,N_43909,N_43762);
nor U48008 (N_48008,N_40525,N_44249);
xnor U48009 (N_48009,N_41171,N_43926);
or U48010 (N_48010,N_43315,N_41942);
or U48011 (N_48011,N_43612,N_40153);
or U48012 (N_48012,N_41787,N_43544);
and U48013 (N_48013,N_43460,N_40033);
nor U48014 (N_48014,N_40611,N_40349);
nand U48015 (N_48015,N_41947,N_42527);
and U48016 (N_48016,N_42784,N_43979);
and U48017 (N_48017,N_40810,N_44426);
and U48018 (N_48018,N_41101,N_43439);
or U48019 (N_48019,N_41682,N_43149);
nor U48020 (N_48020,N_44007,N_43362);
or U48021 (N_48021,N_42687,N_44924);
or U48022 (N_48022,N_41800,N_44170);
and U48023 (N_48023,N_41375,N_41270);
or U48024 (N_48024,N_43642,N_42097);
nor U48025 (N_48025,N_40657,N_41203);
nor U48026 (N_48026,N_41461,N_40825);
xor U48027 (N_48027,N_42503,N_43517);
nand U48028 (N_48028,N_42044,N_43224);
nand U48029 (N_48029,N_42546,N_43783);
nor U48030 (N_48030,N_42265,N_44010);
xnor U48031 (N_48031,N_42037,N_41057);
nor U48032 (N_48032,N_43174,N_43954);
and U48033 (N_48033,N_43924,N_42490);
nor U48034 (N_48034,N_41852,N_42224);
nand U48035 (N_48035,N_43867,N_40981);
nor U48036 (N_48036,N_44638,N_43320);
nand U48037 (N_48037,N_43971,N_40338);
nand U48038 (N_48038,N_42245,N_43315);
nor U48039 (N_48039,N_41186,N_42835);
nor U48040 (N_48040,N_41996,N_41381);
and U48041 (N_48041,N_44777,N_42053);
nor U48042 (N_48042,N_43965,N_43011);
xnor U48043 (N_48043,N_42923,N_44366);
or U48044 (N_48044,N_42757,N_40886);
or U48045 (N_48045,N_43718,N_41120);
or U48046 (N_48046,N_41652,N_43816);
or U48047 (N_48047,N_43783,N_41459);
nor U48048 (N_48048,N_40976,N_40812);
xor U48049 (N_48049,N_41468,N_42449);
xor U48050 (N_48050,N_40757,N_44185);
xor U48051 (N_48051,N_44661,N_43014);
or U48052 (N_48052,N_42899,N_42405);
and U48053 (N_48053,N_40745,N_44328);
nand U48054 (N_48054,N_43225,N_41549);
nand U48055 (N_48055,N_42238,N_40496);
and U48056 (N_48056,N_43554,N_42452);
xnor U48057 (N_48057,N_42829,N_44387);
or U48058 (N_48058,N_40205,N_40975);
nand U48059 (N_48059,N_41750,N_41968);
or U48060 (N_48060,N_42702,N_42551);
xor U48061 (N_48061,N_40758,N_43564);
or U48062 (N_48062,N_44553,N_40831);
xor U48063 (N_48063,N_43645,N_42665);
nor U48064 (N_48064,N_44464,N_42405);
nor U48065 (N_48065,N_44907,N_42908);
nand U48066 (N_48066,N_41034,N_41285);
xnor U48067 (N_48067,N_40114,N_42257);
nor U48068 (N_48068,N_40418,N_40653);
and U48069 (N_48069,N_40269,N_40676);
or U48070 (N_48070,N_42103,N_41470);
and U48071 (N_48071,N_44100,N_44760);
or U48072 (N_48072,N_40592,N_42357);
nand U48073 (N_48073,N_42408,N_43675);
nand U48074 (N_48074,N_42109,N_43812);
or U48075 (N_48075,N_44419,N_41192);
nor U48076 (N_48076,N_42190,N_41616);
and U48077 (N_48077,N_41369,N_44904);
nand U48078 (N_48078,N_42430,N_44772);
and U48079 (N_48079,N_42185,N_42481);
and U48080 (N_48080,N_41781,N_41686);
or U48081 (N_48081,N_40974,N_40412);
nand U48082 (N_48082,N_44737,N_41597);
xnor U48083 (N_48083,N_40810,N_44854);
nor U48084 (N_48084,N_43002,N_41735);
nor U48085 (N_48085,N_40588,N_40885);
or U48086 (N_48086,N_42919,N_43622);
nand U48087 (N_48087,N_44997,N_43774);
and U48088 (N_48088,N_42529,N_40939);
nand U48089 (N_48089,N_44639,N_43553);
nor U48090 (N_48090,N_44867,N_44579);
and U48091 (N_48091,N_40015,N_40699);
nor U48092 (N_48092,N_41637,N_43168);
nand U48093 (N_48093,N_43452,N_40843);
and U48094 (N_48094,N_44529,N_41974);
or U48095 (N_48095,N_43512,N_44630);
xor U48096 (N_48096,N_40153,N_42790);
and U48097 (N_48097,N_44870,N_42503);
nor U48098 (N_48098,N_42266,N_42957);
nand U48099 (N_48099,N_42772,N_41493);
or U48100 (N_48100,N_41705,N_42481);
nor U48101 (N_48101,N_42960,N_42794);
and U48102 (N_48102,N_43517,N_42764);
or U48103 (N_48103,N_41458,N_40920);
xnor U48104 (N_48104,N_43947,N_40829);
or U48105 (N_48105,N_44716,N_43069);
nand U48106 (N_48106,N_43722,N_44669);
xor U48107 (N_48107,N_42050,N_43179);
xor U48108 (N_48108,N_41735,N_43719);
and U48109 (N_48109,N_42213,N_43072);
xnor U48110 (N_48110,N_41035,N_40402);
and U48111 (N_48111,N_42041,N_43269);
and U48112 (N_48112,N_42119,N_42629);
nor U48113 (N_48113,N_43378,N_44788);
or U48114 (N_48114,N_42773,N_41625);
and U48115 (N_48115,N_40202,N_43517);
or U48116 (N_48116,N_43276,N_44151);
nor U48117 (N_48117,N_43256,N_40626);
xor U48118 (N_48118,N_42960,N_43525);
nand U48119 (N_48119,N_44705,N_40004);
nand U48120 (N_48120,N_40518,N_40968);
xnor U48121 (N_48121,N_43052,N_40669);
and U48122 (N_48122,N_43230,N_41162);
nor U48123 (N_48123,N_44299,N_44638);
nor U48124 (N_48124,N_43082,N_44994);
nand U48125 (N_48125,N_43276,N_40588);
or U48126 (N_48126,N_42488,N_43681);
nor U48127 (N_48127,N_44911,N_44212);
or U48128 (N_48128,N_40959,N_43555);
nand U48129 (N_48129,N_41275,N_44059);
nand U48130 (N_48130,N_41937,N_43724);
and U48131 (N_48131,N_41592,N_44021);
and U48132 (N_48132,N_43496,N_40897);
and U48133 (N_48133,N_40048,N_40920);
xnor U48134 (N_48134,N_41030,N_40756);
nor U48135 (N_48135,N_41816,N_41880);
xor U48136 (N_48136,N_43615,N_44370);
nor U48137 (N_48137,N_42926,N_40840);
nand U48138 (N_48138,N_44398,N_42955);
or U48139 (N_48139,N_40929,N_41892);
or U48140 (N_48140,N_41732,N_43272);
nor U48141 (N_48141,N_43170,N_44402);
nand U48142 (N_48142,N_42073,N_40946);
and U48143 (N_48143,N_44685,N_44416);
nor U48144 (N_48144,N_40156,N_40726);
xnor U48145 (N_48145,N_40778,N_40511);
or U48146 (N_48146,N_40154,N_42326);
nand U48147 (N_48147,N_43658,N_43301);
nand U48148 (N_48148,N_42435,N_44393);
nand U48149 (N_48149,N_43304,N_40681);
nand U48150 (N_48150,N_40509,N_41952);
or U48151 (N_48151,N_40083,N_44430);
and U48152 (N_48152,N_43154,N_43978);
nand U48153 (N_48153,N_41563,N_44293);
and U48154 (N_48154,N_44793,N_44371);
or U48155 (N_48155,N_44003,N_44464);
xor U48156 (N_48156,N_42969,N_43430);
nand U48157 (N_48157,N_41294,N_41184);
or U48158 (N_48158,N_43594,N_40866);
and U48159 (N_48159,N_43010,N_42658);
nor U48160 (N_48160,N_42248,N_42403);
or U48161 (N_48161,N_42595,N_44576);
nor U48162 (N_48162,N_40656,N_40438);
or U48163 (N_48163,N_44398,N_41702);
and U48164 (N_48164,N_40437,N_40498);
nor U48165 (N_48165,N_40089,N_43718);
or U48166 (N_48166,N_41281,N_44576);
nand U48167 (N_48167,N_44783,N_42334);
nor U48168 (N_48168,N_42427,N_41166);
xor U48169 (N_48169,N_44533,N_40506);
nand U48170 (N_48170,N_43521,N_40420);
nor U48171 (N_48171,N_42937,N_42931);
nor U48172 (N_48172,N_42537,N_41573);
or U48173 (N_48173,N_42423,N_41929);
nor U48174 (N_48174,N_43187,N_42704);
or U48175 (N_48175,N_44958,N_40682);
or U48176 (N_48176,N_43355,N_44899);
and U48177 (N_48177,N_41958,N_43199);
or U48178 (N_48178,N_40998,N_40440);
xnor U48179 (N_48179,N_42002,N_44396);
nand U48180 (N_48180,N_41560,N_43866);
xor U48181 (N_48181,N_42867,N_41832);
or U48182 (N_48182,N_42004,N_42357);
nand U48183 (N_48183,N_40317,N_41288);
nand U48184 (N_48184,N_41352,N_41756);
nor U48185 (N_48185,N_42735,N_44240);
and U48186 (N_48186,N_40012,N_43910);
and U48187 (N_48187,N_41773,N_44307);
or U48188 (N_48188,N_40657,N_42548);
nand U48189 (N_48189,N_43088,N_43563);
nand U48190 (N_48190,N_40647,N_41900);
xnor U48191 (N_48191,N_44561,N_42253);
nor U48192 (N_48192,N_41949,N_42195);
nand U48193 (N_48193,N_41621,N_43625);
nand U48194 (N_48194,N_40550,N_41305);
xor U48195 (N_48195,N_42784,N_42245);
and U48196 (N_48196,N_43836,N_41753);
nor U48197 (N_48197,N_44831,N_42547);
and U48198 (N_48198,N_42671,N_41792);
and U48199 (N_48199,N_44409,N_44875);
and U48200 (N_48200,N_41506,N_41984);
and U48201 (N_48201,N_44914,N_43115);
xnor U48202 (N_48202,N_42804,N_42857);
xnor U48203 (N_48203,N_40581,N_40005);
or U48204 (N_48204,N_43333,N_42910);
or U48205 (N_48205,N_43468,N_42398);
xor U48206 (N_48206,N_44061,N_41354);
xnor U48207 (N_48207,N_41065,N_44329);
and U48208 (N_48208,N_44379,N_42709);
or U48209 (N_48209,N_42489,N_44446);
or U48210 (N_48210,N_44596,N_40531);
and U48211 (N_48211,N_44709,N_41874);
nor U48212 (N_48212,N_40011,N_43381);
nand U48213 (N_48213,N_42594,N_41185);
nand U48214 (N_48214,N_44669,N_43214);
and U48215 (N_48215,N_43142,N_42553);
xor U48216 (N_48216,N_44126,N_42899);
xor U48217 (N_48217,N_42683,N_40054);
xor U48218 (N_48218,N_44933,N_43867);
xnor U48219 (N_48219,N_40840,N_42521);
nand U48220 (N_48220,N_41528,N_40800);
nor U48221 (N_48221,N_43313,N_40514);
nor U48222 (N_48222,N_43309,N_42125);
or U48223 (N_48223,N_44306,N_44071);
nand U48224 (N_48224,N_40436,N_40386);
or U48225 (N_48225,N_42515,N_43004);
xor U48226 (N_48226,N_40960,N_44254);
xor U48227 (N_48227,N_43800,N_41319);
or U48228 (N_48228,N_42198,N_43314);
or U48229 (N_48229,N_44328,N_43158);
or U48230 (N_48230,N_40856,N_41825);
nand U48231 (N_48231,N_41794,N_42185);
nand U48232 (N_48232,N_41532,N_42831);
xor U48233 (N_48233,N_42399,N_42262);
xor U48234 (N_48234,N_41833,N_44518);
xor U48235 (N_48235,N_41060,N_41445);
xnor U48236 (N_48236,N_41923,N_42162);
and U48237 (N_48237,N_40061,N_40551);
or U48238 (N_48238,N_44298,N_41263);
nand U48239 (N_48239,N_41711,N_41367);
or U48240 (N_48240,N_44812,N_42177);
and U48241 (N_48241,N_40136,N_42464);
nand U48242 (N_48242,N_43249,N_43291);
nor U48243 (N_48243,N_40777,N_40648);
xnor U48244 (N_48244,N_41075,N_41463);
xnor U48245 (N_48245,N_40454,N_42277);
or U48246 (N_48246,N_40821,N_43229);
and U48247 (N_48247,N_42217,N_42570);
or U48248 (N_48248,N_41591,N_42497);
or U48249 (N_48249,N_42980,N_41519);
nor U48250 (N_48250,N_44151,N_43226);
nand U48251 (N_48251,N_41044,N_42497);
nor U48252 (N_48252,N_42646,N_40551);
and U48253 (N_48253,N_44030,N_42184);
or U48254 (N_48254,N_41095,N_43742);
and U48255 (N_48255,N_41503,N_43625);
nor U48256 (N_48256,N_44435,N_42398);
or U48257 (N_48257,N_44718,N_42258);
xor U48258 (N_48258,N_40248,N_42816);
xnor U48259 (N_48259,N_41414,N_44131);
or U48260 (N_48260,N_41412,N_40641);
nor U48261 (N_48261,N_41480,N_41582);
nand U48262 (N_48262,N_42325,N_44715);
and U48263 (N_48263,N_41360,N_41507);
nor U48264 (N_48264,N_44708,N_41549);
nand U48265 (N_48265,N_42538,N_43712);
or U48266 (N_48266,N_40907,N_42755);
nor U48267 (N_48267,N_42000,N_41454);
xnor U48268 (N_48268,N_42323,N_43625);
or U48269 (N_48269,N_40767,N_44587);
or U48270 (N_48270,N_43021,N_44333);
xor U48271 (N_48271,N_43139,N_42632);
and U48272 (N_48272,N_44190,N_44594);
or U48273 (N_48273,N_40867,N_41578);
nor U48274 (N_48274,N_43110,N_41818);
xnor U48275 (N_48275,N_42203,N_40306);
nor U48276 (N_48276,N_44230,N_41073);
or U48277 (N_48277,N_40087,N_41612);
nor U48278 (N_48278,N_43418,N_43860);
xnor U48279 (N_48279,N_43726,N_42541);
nand U48280 (N_48280,N_41479,N_44547);
and U48281 (N_48281,N_41228,N_44831);
nor U48282 (N_48282,N_42079,N_40436);
xor U48283 (N_48283,N_40519,N_44399);
or U48284 (N_48284,N_44437,N_40909);
nand U48285 (N_48285,N_44004,N_43637);
nor U48286 (N_48286,N_40704,N_44399);
or U48287 (N_48287,N_43619,N_43578);
and U48288 (N_48288,N_42285,N_40393);
xor U48289 (N_48289,N_44724,N_43932);
nor U48290 (N_48290,N_43998,N_44676);
and U48291 (N_48291,N_42764,N_40552);
nor U48292 (N_48292,N_44681,N_43669);
nand U48293 (N_48293,N_43816,N_40303);
xor U48294 (N_48294,N_40364,N_43906);
or U48295 (N_48295,N_44881,N_43634);
nor U48296 (N_48296,N_41100,N_44111);
nor U48297 (N_48297,N_43463,N_40824);
and U48298 (N_48298,N_40400,N_41304);
nor U48299 (N_48299,N_42149,N_44845);
or U48300 (N_48300,N_43556,N_42655);
xor U48301 (N_48301,N_44946,N_40599);
xor U48302 (N_48302,N_41881,N_41539);
and U48303 (N_48303,N_40329,N_42407);
xor U48304 (N_48304,N_40286,N_40913);
xor U48305 (N_48305,N_40174,N_40520);
nand U48306 (N_48306,N_44064,N_42969);
xnor U48307 (N_48307,N_44694,N_43363);
xnor U48308 (N_48308,N_43320,N_43302);
or U48309 (N_48309,N_41752,N_40355);
nand U48310 (N_48310,N_44879,N_43532);
xnor U48311 (N_48311,N_41522,N_42299);
nor U48312 (N_48312,N_43144,N_44598);
and U48313 (N_48313,N_42566,N_44952);
or U48314 (N_48314,N_41376,N_42784);
and U48315 (N_48315,N_43337,N_42654);
and U48316 (N_48316,N_40296,N_42488);
or U48317 (N_48317,N_41338,N_41176);
xor U48318 (N_48318,N_44215,N_42313);
nor U48319 (N_48319,N_41909,N_44323);
nand U48320 (N_48320,N_42257,N_42196);
nor U48321 (N_48321,N_41056,N_40597);
and U48322 (N_48322,N_41823,N_44740);
and U48323 (N_48323,N_44569,N_44817);
nor U48324 (N_48324,N_43160,N_41588);
xnor U48325 (N_48325,N_40063,N_42369);
or U48326 (N_48326,N_42439,N_42785);
and U48327 (N_48327,N_40629,N_42355);
nand U48328 (N_48328,N_42790,N_42807);
nor U48329 (N_48329,N_43065,N_41027);
nor U48330 (N_48330,N_41155,N_41523);
nor U48331 (N_48331,N_44162,N_44303);
nor U48332 (N_48332,N_42058,N_44370);
and U48333 (N_48333,N_40676,N_43810);
or U48334 (N_48334,N_40807,N_44103);
nand U48335 (N_48335,N_41365,N_44144);
and U48336 (N_48336,N_41850,N_40323);
or U48337 (N_48337,N_41413,N_40804);
nand U48338 (N_48338,N_44939,N_44570);
xor U48339 (N_48339,N_40839,N_42515);
nand U48340 (N_48340,N_42479,N_43357);
xor U48341 (N_48341,N_40040,N_40835);
nand U48342 (N_48342,N_40914,N_41545);
nand U48343 (N_48343,N_40783,N_44939);
and U48344 (N_48344,N_40313,N_43170);
xnor U48345 (N_48345,N_41699,N_41827);
nand U48346 (N_48346,N_44685,N_41672);
nor U48347 (N_48347,N_40644,N_40700);
or U48348 (N_48348,N_44991,N_41200);
xor U48349 (N_48349,N_40367,N_44889);
xor U48350 (N_48350,N_44546,N_40058);
or U48351 (N_48351,N_43991,N_41071);
nor U48352 (N_48352,N_42687,N_42795);
xnor U48353 (N_48353,N_43783,N_44443);
nand U48354 (N_48354,N_43641,N_40313);
xnor U48355 (N_48355,N_42838,N_43051);
nor U48356 (N_48356,N_40477,N_44890);
xor U48357 (N_48357,N_43142,N_41662);
xnor U48358 (N_48358,N_43253,N_40120);
nor U48359 (N_48359,N_41391,N_43259);
and U48360 (N_48360,N_42192,N_40361);
nor U48361 (N_48361,N_43278,N_43366);
nor U48362 (N_48362,N_43831,N_41199);
nand U48363 (N_48363,N_43048,N_41270);
and U48364 (N_48364,N_44795,N_42915);
nand U48365 (N_48365,N_40589,N_42064);
nor U48366 (N_48366,N_44140,N_44748);
nand U48367 (N_48367,N_42005,N_43773);
nor U48368 (N_48368,N_41047,N_43346);
nand U48369 (N_48369,N_44446,N_41574);
nor U48370 (N_48370,N_44591,N_41736);
nor U48371 (N_48371,N_41591,N_40170);
or U48372 (N_48372,N_41531,N_40767);
or U48373 (N_48373,N_44818,N_44135);
and U48374 (N_48374,N_44185,N_42542);
and U48375 (N_48375,N_40972,N_42042);
nand U48376 (N_48376,N_43086,N_41876);
nor U48377 (N_48377,N_44443,N_41917);
nand U48378 (N_48378,N_40172,N_44536);
xor U48379 (N_48379,N_44848,N_43432);
or U48380 (N_48380,N_43948,N_44585);
nand U48381 (N_48381,N_40271,N_44428);
or U48382 (N_48382,N_42813,N_41692);
xnor U48383 (N_48383,N_41502,N_40192);
nand U48384 (N_48384,N_42263,N_41439);
and U48385 (N_48385,N_43706,N_44103);
nand U48386 (N_48386,N_42702,N_43848);
nand U48387 (N_48387,N_40976,N_44192);
nand U48388 (N_48388,N_42302,N_42033);
xnor U48389 (N_48389,N_43721,N_44789);
xnor U48390 (N_48390,N_42966,N_40611);
xor U48391 (N_48391,N_44551,N_43788);
nor U48392 (N_48392,N_41237,N_43339);
xor U48393 (N_48393,N_44045,N_43050);
nor U48394 (N_48394,N_43377,N_42807);
nand U48395 (N_48395,N_43000,N_42660);
xnor U48396 (N_48396,N_44566,N_41815);
nor U48397 (N_48397,N_40038,N_42865);
and U48398 (N_48398,N_44358,N_42951);
or U48399 (N_48399,N_44272,N_43101);
xnor U48400 (N_48400,N_43049,N_43760);
xor U48401 (N_48401,N_44732,N_41629);
and U48402 (N_48402,N_42196,N_44138);
nand U48403 (N_48403,N_42139,N_43440);
xor U48404 (N_48404,N_40006,N_44344);
xor U48405 (N_48405,N_41165,N_41517);
nor U48406 (N_48406,N_43699,N_43645);
nor U48407 (N_48407,N_43792,N_43102);
xor U48408 (N_48408,N_43350,N_40255);
nand U48409 (N_48409,N_41936,N_42606);
xor U48410 (N_48410,N_40215,N_42168);
nand U48411 (N_48411,N_42477,N_44054);
and U48412 (N_48412,N_40321,N_41216);
nand U48413 (N_48413,N_41973,N_44764);
nor U48414 (N_48414,N_42868,N_42370);
or U48415 (N_48415,N_41153,N_44356);
nor U48416 (N_48416,N_40363,N_43740);
or U48417 (N_48417,N_41711,N_44018);
xor U48418 (N_48418,N_41819,N_41733);
nor U48419 (N_48419,N_43312,N_43641);
nand U48420 (N_48420,N_41920,N_42618);
or U48421 (N_48421,N_44247,N_41333);
xnor U48422 (N_48422,N_42802,N_44617);
or U48423 (N_48423,N_42182,N_40422);
xor U48424 (N_48424,N_43137,N_44675);
nor U48425 (N_48425,N_41546,N_41495);
xor U48426 (N_48426,N_42275,N_44920);
and U48427 (N_48427,N_41129,N_44062);
or U48428 (N_48428,N_43325,N_42421);
and U48429 (N_48429,N_44682,N_43611);
xnor U48430 (N_48430,N_40110,N_42146);
xor U48431 (N_48431,N_43435,N_44542);
and U48432 (N_48432,N_41154,N_44335);
nor U48433 (N_48433,N_40087,N_40278);
or U48434 (N_48434,N_43198,N_40055);
and U48435 (N_48435,N_42951,N_44731);
xnor U48436 (N_48436,N_41267,N_41920);
nor U48437 (N_48437,N_43046,N_40233);
and U48438 (N_48438,N_42347,N_43775);
or U48439 (N_48439,N_41898,N_42502);
xor U48440 (N_48440,N_43072,N_42978);
xnor U48441 (N_48441,N_40231,N_44355);
nand U48442 (N_48442,N_40070,N_43620);
nor U48443 (N_48443,N_43473,N_40943);
or U48444 (N_48444,N_43099,N_43830);
nand U48445 (N_48445,N_43512,N_44611);
and U48446 (N_48446,N_40294,N_41084);
nand U48447 (N_48447,N_43189,N_41371);
or U48448 (N_48448,N_40419,N_43714);
nand U48449 (N_48449,N_41977,N_43247);
nor U48450 (N_48450,N_43192,N_44383);
xnor U48451 (N_48451,N_43511,N_43716);
nor U48452 (N_48452,N_41339,N_43651);
or U48453 (N_48453,N_41525,N_41708);
nand U48454 (N_48454,N_44245,N_42682);
nand U48455 (N_48455,N_42840,N_40824);
xnor U48456 (N_48456,N_44190,N_44366);
or U48457 (N_48457,N_41794,N_44984);
nand U48458 (N_48458,N_44577,N_40862);
or U48459 (N_48459,N_42727,N_40200);
nor U48460 (N_48460,N_42299,N_42080);
nor U48461 (N_48461,N_44624,N_43022);
nor U48462 (N_48462,N_44653,N_40669);
nand U48463 (N_48463,N_40087,N_43278);
xor U48464 (N_48464,N_40930,N_44296);
xnor U48465 (N_48465,N_41017,N_41225);
or U48466 (N_48466,N_41062,N_43745);
nand U48467 (N_48467,N_44489,N_44655);
nand U48468 (N_48468,N_42251,N_43248);
nand U48469 (N_48469,N_42735,N_40530);
xor U48470 (N_48470,N_40064,N_41852);
xor U48471 (N_48471,N_41696,N_43491);
nand U48472 (N_48472,N_42593,N_41691);
nand U48473 (N_48473,N_41561,N_41281);
or U48474 (N_48474,N_44770,N_43693);
nor U48475 (N_48475,N_40172,N_40471);
or U48476 (N_48476,N_42134,N_44397);
nor U48477 (N_48477,N_42512,N_43619);
and U48478 (N_48478,N_41146,N_43690);
nand U48479 (N_48479,N_40616,N_43771);
xor U48480 (N_48480,N_40609,N_40838);
nor U48481 (N_48481,N_43920,N_44686);
or U48482 (N_48482,N_42184,N_41788);
nor U48483 (N_48483,N_41812,N_43894);
nor U48484 (N_48484,N_42817,N_41842);
or U48485 (N_48485,N_44493,N_41060);
nand U48486 (N_48486,N_42947,N_43526);
nand U48487 (N_48487,N_42348,N_41765);
xor U48488 (N_48488,N_43369,N_42567);
xnor U48489 (N_48489,N_40905,N_44296);
nand U48490 (N_48490,N_43704,N_44162);
nand U48491 (N_48491,N_44826,N_41132);
nand U48492 (N_48492,N_42330,N_41645);
and U48493 (N_48493,N_44387,N_40764);
and U48494 (N_48494,N_40442,N_41620);
xnor U48495 (N_48495,N_41434,N_44244);
or U48496 (N_48496,N_40467,N_43140);
or U48497 (N_48497,N_44670,N_43986);
xor U48498 (N_48498,N_42368,N_42173);
and U48499 (N_48499,N_40906,N_44101);
nand U48500 (N_48500,N_41169,N_41079);
and U48501 (N_48501,N_41043,N_43709);
and U48502 (N_48502,N_43931,N_41640);
or U48503 (N_48503,N_44729,N_43148);
nor U48504 (N_48504,N_43440,N_41736);
and U48505 (N_48505,N_44175,N_41026);
and U48506 (N_48506,N_41633,N_43646);
nand U48507 (N_48507,N_43246,N_44947);
xnor U48508 (N_48508,N_44485,N_42198);
xor U48509 (N_48509,N_41430,N_44440);
xnor U48510 (N_48510,N_44972,N_41617);
and U48511 (N_48511,N_44414,N_44835);
and U48512 (N_48512,N_42669,N_44474);
nor U48513 (N_48513,N_42532,N_43016);
or U48514 (N_48514,N_43511,N_44901);
nand U48515 (N_48515,N_40237,N_40514);
or U48516 (N_48516,N_44296,N_44812);
nand U48517 (N_48517,N_42802,N_42033);
xnor U48518 (N_48518,N_40057,N_42730);
nand U48519 (N_48519,N_43219,N_43986);
nand U48520 (N_48520,N_40910,N_44319);
xnor U48521 (N_48521,N_40237,N_42283);
xor U48522 (N_48522,N_43348,N_43362);
xor U48523 (N_48523,N_43736,N_43103);
xor U48524 (N_48524,N_42300,N_43119);
and U48525 (N_48525,N_44263,N_41415);
or U48526 (N_48526,N_44052,N_43035);
nor U48527 (N_48527,N_42847,N_43396);
nor U48528 (N_48528,N_41428,N_43165);
nand U48529 (N_48529,N_42202,N_42603);
nor U48530 (N_48530,N_41466,N_40572);
nor U48531 (N_48531,N_41552,N_44477);
nand U48532 (N_48532,N_41054,N_44074);
xnor U48533 (N_48533,N_43384,N_44582);
nand U48534 (N_48534,N_43631,N_44679);
and U48535 (N_48535,N_42866,N_40621);
nor U48536 (N_48536,N_43248,N_44352);
nand U48537 (N_48537,N_42376,N_43807);
xnor U48538 (N_48538,N_40008,N_40599);
or U48539 (N_48539,N_44134,N_44158);
and U48540 (N_48540,N_41726,N_40342);
or U48541 (N_48541,N_43963,N_44090);
or U48542 (N_48542,N_44549,N_41290);
xnor U48543 (N_48543,N_41063,N_43975);
nor U48544 (N_48544,N_41661,N_44547);
and U48545 (N_48545,N_44420,N_42462);
nor U48546 (N_48546,N_44718,N_40325);
and U48547 (N_48547,N_40049,N_43170);
nor U48548 (N_48548,N_41519,N_43735);
nor U48549 (N_48549,N_40262,N_43087);
and U48550 (N_48550,N_40859,N_41800);
nor U48551 (N_48551,N_44842,N_43402);
nor U48552 (N_48552,N_42908,N_41025);
xnor U48553 (N_48553,N_41681,N_43859);
xor U48554 (N_48554,N_43038,N_42744);
nand U48555 (N_48555,N_43839,N_44096);
and U48556 (N_48556,N_43729,N_42568);
nor U48557 (N_48557,N_40557,N_41578);
nand U48558 (N_48558,N_43811,N_44746);
and U48559 (N_48559,N_41105,N_40797);
and U48560 (N_48560,N_43862,N_41198);
nor U48561 (N_48561,N_43657,N_42585);
or U48562 (N_48562,N_44890,N_44573);
xnor U48563 (N_48563,N_43948,N_40972);
nor U48564 (N_48564,N_41213,N_43121);
or U48565 (N_48565,N_40251,N_44383);
or U48566 (N_48566,N_41750,N_44769);
and U48567 (N_48567,N_40478,N_40813);
nand U48568 (N_48568,N_40285,N_43369);
nor U48569 (N_48569,N_43451,N_41000);
or U48570 (N_48570,N_44256,N_41196);
nor U48571 (N_48571,N_40350,N_43390);
nor U48572 (N_48572,N_44152,N_40533);
and U48573 (N_48573,N_44079,N_43904);
xor U48574 (N_48574,N_44965,N_42944);
or U48575 (N_48575,N_42682,N_42479);
nor U48576 (N_48576,N_43228,N_40488);
and U48577 (N_48577,N_44196,N_42386);
and U48578 (N_48578,N_42756,N_43562);
nand U48579 (N_48579,N_42899,N_44971);
or U48580 (N_48580,N_42425,N_44529);
and U48581 (N_48581,N_40904,N_40959);
xor U48582 (N_48582,N_41743,N_42440);
xnor U48583 (N_48583,N_42887,N_41612);
nand U48584 (N_48584,N_40195,N_43144);
nor U48585 (N_48585,N_42804,N_41083);
and U48586 (N_48586,N_43258,N_42426);
and U48587 (N_48587,N_42810,N_40418);
nor U48588 (N_48588,N_40866,N_43114);
nor U48589 (N_48589,N_43731,N_40499);
nor U48590 (N_48590,N_43070,N_41987);
and U48591 (N_48591,N_43996,N_40016);
and U48592 (N_48592,N_43684,N_40141);
and U48593 (N_48593,N_40583,N_44181);
or U48594 (N_48594,N_41440,N_44255);
and U48595 (N_48595,N_42863,N_40496);
nor U48596 (N_48596,N_44038,N_41983);
xor U48597 (N_48597,N_42904,N_41656);
xor U48598 (N_48598,N_40561,N_42990);
xor U48599 (N_48599,N_43466,N_43118);
and U48600 (N_48600,N_43899,N_40431);
nor U48601 (N_48601,N_42688,N_43311);
nand U48602 (N_48602,N_42064,N_43550);
or U48603 (N_48603,N_40047,N_43683);
nor U48604 (N_48604,N_42945,N_43158);
nand U48605 (N_48605,N_43434,N_43754);
nand U48606 (N_48606,N_40217,N_43633);
nand U48607 (N_48607,N_43380,N_43212);
and U48608 (N_48608,N_40369,N_44122);
xnor U48609 (N_48609,N_44934,N_41997);
and U48610 (N_48610,N_42229,N_43428);
xnor U48611 (N_48611,N_44605,N_41158);
or U48612 (N_48612,N_41922,N_41331);
nor U48613 (N_48613,N_44647,N_44246);
nor U48614 (N_48614,N_43227,N_40884);
nor U48615 (N_48615,N_42537,N_40419);
and U48616 (N_48616,N_41708,N_42586);
or U48617 (N_48617,N_41952,N_40562);
nand U48618 (N_48618,N_43770,N_41291);
and U48619 (N_48619,N_41801,N_41593);
nand U48620 (N_48620,N_41491,N_42797);
or U48621 (N_48621,N_40239,N_41601);
nand U48622 (N_48622,N_42381,N_43447);
and U48623 (N_48623,N_44146,N_44171);
nand U48624 (N_48624,N_40879,N_44077);
and U48625 (N_48625,N_43218,N_41213);
or U48626 (N_48626,N_41870,N_42668);
nor U48627 (N_48627,N_41225,N_42775);
xor U48628 (N_48628,N_44324,N_42387);
nand U48629 (N_48629,N_41092,N_44684);
or U48630 (N_48630,N_42294,N_43414);
nor U48631 (N_48631,N_41557,N_42188);
and U48632 (N_48632,N_41026,N_44399);
and U48633 (N_48633,N_40240,N_43689);
xnor U48634 (N_48634,N_40480,N_40211);
nand U48635 (N_48635,N_44314,N_43545);
or U48636 (N_48636,N_42270,N_40766);
nand U48637 (N_48637,N_44047,N_42331);
or U48638 (N_48638,N_41264,N_44766);
nor U48639 (N_48639,N_43251,N_44909);
or U48640 (N_48640,N_44575,N_44194);
and U48641 (N_48641,N_42401,N_42036);
or U48642 (N_48642,N_40612,N_44573);
nand U48643 (N_48643,N_41594,N_42732);
nor U48644 (N_48644,N_43837,N_40823);
nor U48645 (N_48645,N_44661,N_42560);
nand U48646 (N_48646,N_42735,N_43908);
nor U48647 (N_48647,N_42398,N_42039);
xor U48648 (N_48648,N_42622,N_41995);
nor U48649 (N_48649,N_43984,N_40957);
xnor U48650 (N_48650,N_42795,N_44655);
xnor U48651 (N_48651,N_40358,N_44079);
and U48652 (N_48652,N_42641,N_44015);
xor U48653 (N_48653,N_44226,N_43971);
nor U48654 (N_48654,N_40085,N_40614);
or U48655 (N_48655,N_43187,N_43179);
nand U48656 (N_48656,N_42760,N_43998);
nand U48657 (N_48657,N_43474,N_42716);
nand U48658 (N_48658,N_43859,N_43140);
xnor U48659 (N_48659,N_41514,N_44872);
nand U48660 (N_48660,N_40161,N_41425);
or U48661 (N_48661,N_41943,N_40096);
and U48662 (N_48662,N_40855,N_40476);
nor U48663 (N_48663,N_40365,N_40997);
nand U48664 (N_48664,N_40352,N_42574);
nor U48665 (N_48665,N_41827,N_41544);
or U48666 (N_48666,N_43088,N_40116);
nor U48667 (N_48667,N_41525,N_42155);
and U48668 (N_48668,N_42711,N_41110);
nand U48669 (N_48669,N_40812,N_44064);
nand U48670 (N_48670,N_42213,N_42480);
or U48671 (N_48671,N_40170,N_42376);
and U48672 (N_48672,N_44225,N_42608);
xnor U48673 (N_48673,N_42371,N_43458);
and U48674 (N_48674,N_42267,N_42471);
nor U48675 (N_48675,N_42725,N_43431);
or U48676 (N_48676,N_40680,N_41196);
nor U48677 (N_48677,N_40518,N_41550);
xor U48678 (N_48678,N_41967,N_40397);
nand U48679 (N_48679,N_43845,N_44989);
or U48680 (N_48680,N_43360,N_41271);
or U48681 (N_48681,N_42619,N_44083);
nor U48682 (N_48682,N_42315,N_42631);
nor U48683 (N_48683,N_42696,N_41962);
nand U48684 (N_48684,N_42966,N_42456);
or U48685 (N_48685,N_40686,N_40239);
nor U48686 (N_48686,N_40978,N_43218);
and U48687 (N_48687,N_41728,N_42481);
xnor U48688 (N_48688,N_40134,N_40874);
xor U48689 (N_48689,N_42866,N_41876);
nand U48690 (N_48690,N_43913,N_40609);
nand U48691 (N_48691,N_41735,N_44630);
and U48692 (N_48692,N_43685,N_42599);
nand U48693 (N_48693,N_40483,N_40642);
or U48694 (N_48694,N_44509,N_41817);
or U48695 (N_48695,N_41176,N_41360);
nand U48696 (N_48696,N_42414,N_41761);
xnor U48697 (N_48697,N_42399,N_44975);
nand U48698 (N_48698,N_43785,N_43587);
or U48699 (N_48699,N_44285,N_43833);
nand U48700 (N_48700,N_43355,N_43922);
and U48701 (N_48701,N_41202,N_44322);
xnor U48702 (N_48702,N_42145,N_42413);
xor U48703 (N_48703,N_43777,N_40259);
and U48704 (N_48704,N_44007,N_42310);
or U48705 (N_48705,N_44823,N_43986);
nor U48706 (N_48706,N_43358,N_42110);
nand U48707 (N_48707,N_41828,N_42689);
nor U48708 (N_48708,N_41962,N_43105);
xnor U48709 (N_48709,N_43396,N_42922);
and U48710 (N_48710,N_43769,N_42444);
and U48711 (N_48711,N_41299,N_42865);
or U48712 (N_48712,N_43211,N_41892);
or U48713 (N_48713,N_41216,N_40341);
nor U48714 (N_48714,N_40816,N_41262);
or U48715 (N_48715,N_44456,N_44465);
nor U48716 (N_48716,N_42721,N_42863);
xor U48717 (N_48717,N_41828,N_43556);
xor U48718 (N_48718,N_40593,N_44129);
xor U48719 (N_48719,N_44934,N_40509);
nor U48720 (N_48720,N_41375,N_41306);
nor U48721 (N_48721,N_44085,N_42318);
or U48722 (N_48722,N_41530,N_42534);
nand U48723 (N_48723,N_41126,N_43937);
nand U48724 (N_48724,N_41813,N_43250);
nor U48725 (N_48725,N_43488,N_41610);
xnor U48726 (N_48726,N_43308,N_40155);
and U48727 (N_48727,N_40198,N_44657);
or U48728 (N_48728,N_43196,N_43521);
nand U48729 (N_48729,N_40494,N_43060);
or U48730 (N_48730,N_40300,N_41805);
xor U48731 (N_48731,N_42538,N_43969);
or U48732 (N_48732,N_43081,N_42390);
xnor U48733 (N_48733,N_40796,N_42576);
or U48734 (N_48734,N_44817,N_40187);
xnor U48735 (N_48735,N_43753,N_44832);
nand U48736 (N_48736,N_40414,N_44170);
or U48737 (N_48737,N_40959,N_42570);
nor U48738 (N_48738,N_42066,N_40136);
and U48739 (N_48739,N_43054,N_43389);
nand U48740 (N_48740,N_40019,N_40336);
nand U48741 (N_48741,N_44464,N_40217);
nand U48742 (N_48742,N_41577,N_42487);
and U48743 (N_48743,N_42727,N_41289);
and U48744 (N_48744,N_44209,N_43053);
nor U48745 (N_48745,N_44880,N_42725);
and U48746 (N_48746,N_41547,N_40526);
nor U48747 (N_48747,N_44454,N_43688);
xor U48748 (N_48748,N_41240,N_44260);
or U48749 (N_48749,N_44679,N_42997);
and U48750 (N_48750,N_42042,N_44401);
and U48751 (N_48751,N_40215,N_40487);
xnor U48752 (N_48752,N_43533,N_44302);
nand U48753 (N_48753,N_44645,N_42333);
xor U48754 (N_48754,N_44907,N_43459);
nor U48755 (N_48755,N_44266,N_40226);
nand U48756 (N_48756,N_44464,N_44023);
and U48757 (N_48757,N_44230,N_41194);
xor U48758 (N_48758,N_41648,N_40747);
nand U48759 (N_48759,N_44917,N_44361);
and U48760 (N_48760,N_43644,N_42975);
or U48761 (N_48761,N_44783,N_42159);
xnor U48762 (N_48762,N_40958,N_44284);
nor U48763 (N_48763,N_43478,N_41177);
nand U48764 (N_48764,N_42637,N_42789);
xor U48765 (N_48765,N_43106,N_43616);
nor U48766 (N_48766,N_41224,N_42666);
or U48767 (N_48767,N_44898,N_40124);
nand U48768 (N_48768,N_41154,N_42643);
or U48769 (N_48769,N_44745,N_43630);
nand U48770 (N_48770,N_42531,N_43282);
xor U48771 (N_48771,N_42458,N_43333);
or U48772 (N_48772,N_41017,N_43892);
and U48773 (N_48773,N_40454,N_44006);
or U48774 (N_48774,N_42001,N_42942);
xor U48775 (N_48775,N_43438,N_42138);
or U48776 (N_48776,N_44162,N_40701);
nor U48777 (N_48777,N_42571,N_44324);
nor U48778 (N_48778,N_41828,N_41152);
or U48779 (N_48779,N_40699,N_41490);
nand U48780 (N_48780,N_42938,N_40459);
xor U48781 (N_48781,N_41640,N_44781);
nor U48782 (N_48782,N_40314,N_41272);
or U48783 (N_48783,N_42935,N_40421);
xor U48784 (N_48784,N_41376,N_42229);
nor U48785 (N_48785,N_44338,N_40490);
xnor U48786 (N_48786,N_42636,N_43905);
xnor U48787 (N_48787,N_43347,N_43434);
nor U48788 (N_48788,N_43082,N_41984);
nand U48789 (N_48789,N_42555,N_42236);
nand U48790 (N_48790,N_42326,N_44469);
nor U48791 (N_48791,N_43079,N_44172);
and U48792 (N_48792,N_41672,N_40349);
nor U48793 (N_48793,N_41620,N_44081);
xor U48794 (N_48794,N_43442,N_41705);
nor U48795 (N_48795,N_41434,N_42333);
or U48796 (N_48796,N_40006,N_40689);
and U48797 (N_48797,N_44357,N_44126);
and U48798 (N_48798,N_41382,N_42974);
and U48799 (N_48799,N_43387,N_42886);
nand U48800 (N_48800,N_41087,N_40494);
nand U48801 (N_48801,N_40556,N_43581);
nand U48802 (N_48802,N_42946,N_42285);
xnor U48803 (N_48803,N_41785,N_40171);
xnor U48804 (N_48804,N_43838,N_42813);
xnor U48805 (N_48805,N_40180,N_40911);
nor U48806 (N_48806,N_44771,N_44251);
nor U48807 (N_48807,N_41178,N_43164);
xnor U48808 (N_48808,N_41053,N_42553);
and U48809 (N_48809,N_44545,N_41124);
or U48810 (N_48810,N_42400,N_43871);
and U48811 (N_48811,N_41556,N_44664);
or U48812 (N_48812,N_44687,N_44662);
xnor U48813 (N_48813,N_44046,N_40806);
nor U48814 (N_48814,N_40748,N_43705);
xnor U48815 (N_48815,N_40861,N_40724);
nand U48816 (N_48816,N_44834,N_43964);
xnor U48817 (N_48817,N_42261,N_43006);
xnor U48818 (N_48818,N_44625,N_42883);
nand U48819 (N_48819,N_43411,N_44757);
or U48820 (N_48820,N_40136,N_44764);
or U48821 (N_48821,N_42958,N_40589);
nand U48822 (N_48822,N_41922,N_43474);
and U48823 (N_48823,N_41169,N_42821);
xnor U48824 (N_48824,N_43398,N_40841);
or U48825 (N_48825,N_40596,N_41911);
nand U48826 (N_48826,N_43081,N_43672);
and U48827 (N_48827,N_41999,N_40043);
nor U48828 (N_48828,N_42315,N_40932);
or U48829 (N_48829,N_41886,N_44945);
xnor U48830 (N_48830,N_40348,N_43743);
nand U48831 (N_48831,N_42981,N_40483);
xor U48832 (N_48832,N_42891,N_43516);
nand U48833 (N_48833,N_44762,N_43100);
or U48834 (N_48834,N_43197,N_40976);
or U48835 (N_48835,N_41620,N_44941);
nand U48836 (N_48836,N_40710,N_43040);
xor U48837 (N_48837,N_43248,N_42370);
nand U48838 (N_48838,N_44744,N_40078);
or U48839 (N_48839,N_43206,N_43416);
nor U48840 (N_48840,N_42045,N_44312);
xnor U48841 (N_48841,N_40537,N_41604);
or U48842 (N_48842,N_42546,N_41521);
or U48843 (N_48843,N_42124,N_42679);
xnor U48844 (N_48844,N_43897,N_44200);
or U48845 (N_48845,N_40090,N_41624);
nor U48846 (N_48846,N_44620,N_43165);
xor U48847 (N_48847,N_44724,N_42134);
and U48848 (N_48848,N_44986,N_41204);
nand U48849 (N_48849,N_40832,N_40486);
and U48850 (N_48850,N_41456,N_43459);
xor U48851 (N_48851,N_41071,N_43299);
xnor U48852 (N_48852,N_41947,N_43608);
or U48853 (N_48853,N_41399,N_42407);
and U48854 (N_48854,N_42767,N_44737);
and U48855 (N_48855,N_44314,N_40462);
xor U48856 (N_48856,N_44720,N_42549);
or U48857 (N_48857,N_41950,N_44474);
or U48858 (N_48858,N_43503,N_44588);
and U48859 (N_48859,N_41806,N_41280);
or U48860 (N_48860,N_40942,N_44737);
and U48861 (N_48861,N_44684,N_42529);
and U48862 (N_48862,N_44861,N_43851);
nor U48863 (N_48863,N_41269,N_41635);
nand U48864 (N_48864,N_41701,N_44265);
or U48865 (N_48865,N_43746,N_44052);
and U48866 (N_48866,N_40889,N_40485);
and U48867 (N_48867,N_43387,N_40767);
and U48868 (N_48868,N_41763,N_41852);
or U48869 (N_48869,N_44642,N_40035);
and U48870 (N_48870,N_40967,N_44255);
nor U48871 (N_48871,N_43358,N_41590);
or U48872 (N_48872,N_41019,N_43983);
xor U48873 (N_48873,N_43391,N_40414);
xnor U48874 (N_48874,N_40481,N_42350);
and U48875 (N_48875,N_44244,N_44291);
xor U48876 (N_48876,N_43235,N_43328);
nor U48877 (N_48877,N_43792,N_40288);
nand U48878 (N_48878,N_43036,N_40810);
or U48879 (N_48879,N_42731,N_44512);
nand U48880 (N_48880,N_42172,N_40595);
nor U48881 (N_48881,N_44696,N_43935);
or U48882 (N_48882,N_40263,N_40474);
xnor U48883 (N_48883,N_43397,N_44254);
and U48884 (N_48884,N_44133,N_41943);
nor U48885 (N_48885,N_40534,N_40851);
xor U48886 (N_48886,N_40434,N_42637);
xor U48887 (N_48887,N_42117,N_43642);
nor U48888 (N_48888,N_41434,N_43559);
or U48889 (N_48889,N_43081,N_42093);
or U48890 (N_48890,N_42681,N_41031);
or U48891 (N_48891,N_42147,N_44155);
xor U48892 (N_48892,N_42985,N_43771);
nor U48893 (N_48893,N_40698,N_41309);
xor U48894 (N_48894,N_44918,N_44542);
nor U48895 (N_48895,N_44560,N_40455);
and U48896 (N_48896,N_42545,N_44483);
xor U48897 (N_48897,N_41619,N_44129);
xnor U48898 (N_48898,N_41743,N_40328);
nor U48899 (N_48899,N_41763,N_41373);
xnor U48900 (N_48900,N_40731,N_40002);
nand U48901 (N_48901,N_41457,N_44787);
nand U48902 (N_48902,N_40800,N_42473);
nor U48903 (N_48903,N_41220,N_40766);
nand U48904 (N_48904,N_44624,N_44980);
or U48905 (N_48905,N_43509,N_40735);
or U48906 (N_48906,N_41161,N_43778);
xnor U48907 (N_48907,N_44110,N_41760);
and U48908 (N_48908,N_42061,N_44940);
nand U48909 (N_48909,N_43957,N_40791);
nor U48910 (N_48910,N_44311,N_42806);
and U48911 (N_48911,N_42111,N_43848);
or U48912 (N_48912,N_42725,N_44504);
or U48913 (N_48913,N_40765,N_42115);
nor U48914 (N_48914,N_41947,N_41159);
nor U48915 (N_48915,N_40992,N_42075);
xnor U48916 (N_48916,N_43960,N_40797);
nor U48917 (N_48917,N_44741,N_43276);
xor U48918 (N_48918,N_41779,N_40752);
or U48919 (N_48919,N_44987,N_41070);
or U48920 (N_48920,N_42611,N_43423);
nand U48921 (N_48921,N_42596,N_43430);
nor U48922 (N_48922,N_40592,N_42274);
nand U48923 (N_48923,N_43350,N_40470);
nand U48924 (N_48924,N_40380,N_40824);
xnor U48925 (N_48925,N_44578,N_43527);
nand U48926 (N_48926,N_44995,N_44840);
nor U48927 (N_48927,N_40289,N_44138);
xnor U48928 (N_48928,N_44293,N_40043);
or U48929 (N_48929,N_40576,N_42789);
nand U48930 (N_48930,N_44705,N_44849);
nand U48931 (N_48931,N_40133,N_42705);
and U48932 (N_48932,N_42486,N_41664);
xor U48933 (N_48933,N_41707,N_40488);
or U48934 (N_48934,N_42295,N_42385);
xor U48935 (N_48935,N_44955,N_44373);
nor U48936 (N_48936,N_44436,N_40530);
nor U48937 (N_48937,N_42182,N_42840);
and U48938 (N_48938,N_40744,N_41938);
and U48939 (N_48939,N_43005,N_40465);
nand U48940 (N_48940,N_43080,N_40377);
or U48941 (N_48941,N_43315,N_40902);
and U48942 (N_48942,N_41576,N_43275);
xnor U48943 (N_48943,N_44849,N_44797);
nand U48944 (N_48944,N_43484,N_41497);
nor U48945 (N_48945,N_41769,N_42470);
or U48946 (N_48946,N_40246,N_42516);
nand U48947 (N_48947,N_40828,N_41982);
nor U48948 (N_48948,N_42156,N_40050);
nand U48949 (N_48949,N_44572,N_44901);
or U48950 (N_48950,N_41053,N_41058);
nor U48951 (N_48951,N_44400,N_44226);
and U48952 (N_48952,N_43249,N_42570);
nor U48953 (N_48953,N_40260,N_42426);
nand U48954 (N_48954,N_41259,N_44310);
nor U48955 (N_48955,N_40570,N_44409);
xnor U48956 (N_48956,N_41324,N_42432);
xnor U48957 (N_48957,N_42208,N_42697);
xor U48958 (N_48958,N_42530,N_40257);
or U48959 (N_48959,N_41131,N_43186);
nand U48960 (N_48960,N_43946,N_41501);
xor U48961 (N_48961,N_43978,N_44121);
xor U48962 (N_48962,N_41221,N_43617);
xor U48963 (N_48963,N_42994,N_44281);
xnor U48964 (N_48964,N_40773,N_41110);
nor U48965 (N_48965,N_40220,N_40241);
nand U48966 (N_48966,N_41512,N_42956);
or U48967 (N_48967,N_41520,N_44880);
nor U48968 (N_48968,N_42812,N_41333);
or U48969 (N_48969,N_41515,N_44897);
nor U48970 (N_48970,N_42835,N_40716);
nor U48971 (N_48971,N_44136,N_41742);
xor U48972 (N_48972,N_44981,N_42911);
and U48973 (N_48973,N_41704,N_40771);
or U48974 (N_48974,N_40944,N_43005);
nand U48975 (N_48975,N_44626,N_42289);
or U48976 (N_48976,N_40552,N_43669);
and U48977 (N_48977,N_44629,N_42522);
nand U48978 (N_48978,N_44353,N_41168);
nand U48979 (N_48979,N_41649,N_44597);
and U48980 (N_48980,N_42030,N_44756);
xnor U48981 (N_48981,N_44179,N_41791);
or U48982 (N_48982,N_43454,N_42114);
nor U48983 (N_48983,N_40597,N_43759);
nor U48984 (N_48984,N_44390,N_43028);
or U48985 (N_48985,N_43190,N_42573);
or U48986 (N_48986,N_44629,N_40579);
and U48987 (N_48987,N_40822,N_43691);
xor U48988 (N_48988,N_40683,N_42886);
nor U48989 (N_48989,N_44247,N_41962);
xnor U48990 (N_48990,N_41026,N_40519);
and U48991 (N_48991,N_41244,N_41524);
and U48992 (N_48992,N_44884,N_41810);
and U48993 (N_48993,N_42519,N_43482);
and U48994 (N_48994,N_41369,N_44757);
nand U48995 (N_48995,N_42506,N_43559);
or U48996 (N_48996,N_42207,N_41125);
nor U48997 (N_48997,N_41969,N_40523);
and U48998 (N_48998,N_42364,N_41734);
or U48999 (N_48999,N_43487,N_40302);
xor U49000 (N_49000,N_42602,N_42545);
nand U49001 (N_49001,N_42798,N_40969);
nand U49002 (N_49002,N_41540,N_41400);
and U49003 (N_49003,N_41210,N_43768);
and U49004 (N_49004,N_40413,N_43242);
nand U49005 (N_49005,N_44981,N_44523);
nand U49006 (N_49006,N_42398,N_44592);
nand U49007 (N_49007,N_40863,N_40821);
or U49008 (N_49008,N_41331,N_42437);
and U49009 (N_49009,N_44821,N_44280);
and U49010 (N_49010,N_40705,N_40927);
xor U49011 (N_49011,N_40235,N_44417);
nor U49012 (N_49012,N_42400,N_41705);
and U49013 (N_49013,N_42543,N_44170);
nand U49014 (N_49014,N_44066,N_43387);
xor U49015 (N_49015,N_43741,N_43024);
xor U49016 (N_49016,N_43976,N_41750);
and U49017 (N_49017,N_43539,N_41450);
or U49018 (N_49018,N_41314,N_43609);
or U49019 (N_49019,N_41439,N_43837);
and U49020 (N_49020,N_43619,N_44427);
nand U49021 (N_49021,N_40724,N_44710);
or U49022 (N_49022,N_44056,N_43859);
nand U49023 (N_49023,N_41947,N_40130);
and U49024 (N_49024,N_40864,N_44221);
nor U49025 (N_49025,N_41820,N_42268);
and U49026 (N_49026,N_44390,N_41589);
xnor U49027 (N_49027,N_41714,N_41341);
nand U49028 (N_49028,N_43186,N_41560);
and U49029 (N_49029,N_42057,N_42139);
or U49030 (N_49030,N_42246,N_41052);
xnor U49031 (N_49031,N_42618,N_43623);
or U49032 (N_49032,N_44476,N_42964);
nor U49033 (N_49033,N_43147,N_44805);
nor U49034 (N_49034,N_41347,N_40197);
and U49035 (N_49035,N_41935,N_40501);
nor U49036 (N_49036,N_42989,N_40465);
nor U49037 (N_49037,N_43648,N_44303);
or U49038 (N_49038,N_41468,N_40591);
xnor U49039 (N_49039,N_42288,N_44481);
nor U49040 (N_49040,N_42320,N_42552);
nor U49041 (N_49041,N_42317,N_43388);
nor U49042 (N_49042,N_41467,N_40755);
and U49043 (N_49043,N_44458,N_40246);
and U49044 (N_49044,N_44831,N_41795);
xnor U49045 (N_49045,N_44804,N_42245);
xor U49046 (N_49046,N_41223,N_43064);
and U49047 (N_49047,N_42742,N_44816);
or U49048 (N_49048,N_43871,N_41342);
nor U49049 (N_49049,N_43629,N_41206);
xnor U49050 (N_49050,N_42531,N_40425);
nor U49051 (N_49051,N_43817,N_40529);
nand U49052 (N_49052,N_43450,N_44395);
nor U49053 (N_49053,N_41033,N_40895);
xnor U49054 (N_49054,N_42917,N_41730);
or U49055 (N_49055,N_42029,N_44494);
xor U49056 (N_49056,N_40641,N_41082);
or U49057 (N_49057,N_40934,N_44758);
nand U49058 (N_49058,N_44621,N_40358);
and U49059 (N_49059,N_44861,N_42234);
nand U49060 (N_49060,N_44534,N_40625);
and U49061 (N_49061,N_44003,N_42835);
and U49062 (N_49062,N_44145,N_42458);
or U49063 (N_49063,N_40654,N_40317);
nand U49064 (N_49064,N_41196,N_44409);
nand U49065 (N_49065,N_44593,N_40168);
nor U49066 (N_49066,N_44059,N_42522);
and U49067 (N_49067,N_42871,N_43409);
nand U49068 (N_49068,N_41341,N_43958);
or U49069 (N_49069,N_42124,N_41040);
and U49070 (N_49070,N_40607,N_43474);
nand U49071 (N_49071,N_44778,N_44332);
nand U49072 (N_49072,N_41502,N_41997);
or U49073 (N_49073,N_42536,N_44667);
nand U49074 (N_49074,N_43076,N_44464);
nor U49075 (N_49075,N_42304,N_44980);
or U49076 (N_49076,N_41229,N_40426);
or U49077 (N_49077,N_43217,N_41555);
or U49078 (N_49078,N_41035,N_41481);
xor U49079 (N_49079,N_41066,N_41665);
nor U49080 (N_49080,N_41832,N_43177);
nand U49081 (N_49081,N_42812,N_40374);
xor U49082 (N_49082,N_43138,N_44345);
and U49083 (N_49083,N_41978,N_43440);
and U49084 (N_49084,N_41717,N_43951);
or U49085 (N_49085,N_43494,N_43479);
and U49086 (N_49086,N_42912,N_41795);
nand U49087 (N_49087,N_40930,N_42197);
nand U49088 (N_49088,N_44481,N_42725);
xor U49089 (N_49089,N_40021,N_42761);
nand U49090 (N_49090,N_41958,N_43959);
nor U49091 (N_49091,N_41430,N_42299);
xor U49092 (N_49092,N_41323,N_44536);
or U49093 (N_49093,N_43555,N_40291);
and U49094 (N_49094,N_42891,N_40228);
or U49095 (N_49095,N_42529,N_43062);
and U49096 (N_49096,N_44496,N_40650);
nor U49097 (N_49097,N_40175,N_42663);
and U49098 (N_49098,N_42511,N_43102);
xor U49099 (N_49099,N_43369,N_42167);
nand U49100 (N_49100,N_43801,N_42738);
nand U49101 (N_49101,N_43549,N_43598);
xor U49102 (N_49102,N_42446,N_42962);
nor U49103 (N_49103,N_40608,N_43728);
nand U49104 (N_49104,N_42552,N_40025);
nor U49105 (N_49105,N_42928,N_41574);
and U49106 (N_49106,N_40628,N_40541);
nand U49107 (N_49107,N_43782,N_43995);
xnor U49108 (N_49108,N_44029,N_43684);
and U49109 (N_49109,N_40323,N_42835);
and U49110 (N_49110,N_41369,N_43704);
xor U49111 (N_49111,N_41353,N_42406);
nor U49112 (N_49112,N_41300,N_42361);
nor U49113 (N_49113,N_40639,N_43773);
nor U49114 (N_49114,N_40255,N_44301);
or U49115 (N_49115,N_44589,N_40725);
or U49116 (N_49116,N_41908,N_44824);
or U49117 (N_49117,N_40094,N_44203);
or U49118 (N_49118,N_42547,N_43151);
xor U49119 (N_49119,N_41276,N_44852);
nand U49120 (N_49120,N_40015,N_42921);
nand U49121 (N_49121,N_43563,N_41378);
and U49122 (N_49122,N_40046,N_41487);
nand U49123 (N_49123,N_43355,N_40057);
or U49124 (N_49124,N_40494,N_44879);
xnor U49125 (N_49125,N_40845,N_40967);
nand U49126 (N_49126,N_41320,N_41403);
and U49127 (N_49127,N_40751,N_41857);
nand U49128 (N_49128,N_41282,N_40584);
nor U49129 (N_49129,N_41565,N_42119);
nand U49130 (N_49130,N_41956,N_41875);
nor U49131 (N_49131,N_42457,N_44649);
and U49132 (N_49132,N_43189,N_41936);
and U49133 (N_49133,N_44081,N_43685);
nand U49134 (N_49134,N_40469,N_44429);
and U49135 (N_49135,N_43462,N_41299);
and U49136 (N_49136,N_42592,N_41770);
nor U49137 (N_49137,N_40034,N_41064);
nor U49138 (N_49138,N_40434,N_41346);
or U49139 (N_49139,N_43026,N_40156);
nand U49140 (N_49140,N_44406,N_40852);
nor U49141 (N_49141,N_42990,N_44492);
or U49142 (N_49142,N_43104,N_42399);
or U49143 (N_49143,N_42129,N_41451);
nor U49144 (N_49144,N_44265,N_43466);
xnor U49145 (N_49145,N_43332,N_43581);
or U49146 (N_49146,N_44550,N_42694);
xor U49147 (N_49147,N_40093,N_44643);
xor U49148 (N_49148,N_41816,N_43568);
or U49149 (N_49149,N_44007,N_43630);
nor U49150 (N_49150,N_42776,N_44506);
nor U49151 (N_49151,N_41635,N_42074);
nor U49152 (N_49152,N_40420,N_41491);
nor U49153 (N_49153,N_41052,N_44258);
xor U49154 (N_49154,N_41956,N_40396);
xor U49155 (N_49155,N_40476,N_41218);
and U49156 (N_49156,N_43722,N_42404);
nand U49157 (N_49157,N_43557,N_41730);
nand U49158 (N_49158,N_42339,N_44532);
xor U49159 (N_49159,N_44166,N_40838);
and U49160 (N_49160,N_44600,N_42000);
and U49161 (N_49161,N_41606,N_43413);
nand U49162 (N_49162,N_40964,N_43132);
xor U49163 (N_49163,N_44711,N_40050);
and U49164 (N_49164,N_44267,N_40071);
xnor U49165 (N_49165,N_42380,N_40123);
and U49166 (N_49166,N_43107,N_40294);
or U49167 (N_49167,N_42814,N_44649);
nor U49168 (N_49168,N_44136,N_42817);
nor U49169 (N_49169,N_40926,N_41358);
nand U49170 (N_49170,N_41820,N_43789);
nand U49171 (N_49171,N_43959,N_44162);
nand U49172 (N_49172,N_44229,N_41941);
and U49173 (N_49173,N_41961,N_42702);
nor U49174 (N_49174,N_44677,N_40341);
nor U49175 (N_49175,N_41614,N_43428);
or U49176 (N_49176,N_40449,N_40037);
xor U49177 (N_49177,N_42889,N_44486);
or U49178 (N_49178,N_42588,N_40592);
and U49179 (N_49179,N_44987,N_42053);
nand U49180 (N_49180,N_44286,N_44378);
xnor U49181 (N_49181,N_41959,N_41988);
and U49182 (N_49182,N_42602,N_42209);
or U49183 (N_49183,N_43899,N_42916);
xnor U49184 (N_49184,N_43653,N_44040);
xor U49185 (N_49185,N_43141,N_40241);
xnor U49186 (N_49186,N_40692,N_41608);
nand U49187 (N_49187,N_42170,N_42650);
or U49188 (N_49188,N_42548,N_43092);
nand U49189 (N_49189,N_41851,N_42616);
or U49190 (N_49190,N_42048,N_41635);
and U49191 (N_49191,N_41207,N_43380);
nand U49192 (N_49192,N_42115,N_44012);
xor U49193 (N_49193,N_40522,N_43050);
nand U49194 (N_49194,N_43184,N_41224);
nand U49195 (N_49195,N_41501,N_42660);
and U49196 (N_49196,N_40271,N_40421);
and U49197 (N_49197,N_41249,N_42166);
and U49198 (N_49198,N_41615,N_40646);
nor U49199 (N_49199,N_42755,N_43369);
and U49200 (N_49200,N_41746,N_41807);
nand U49201 (N_49201,N_40005,N_43635);
nand U49202 (N_49202,N_44169,N_44168);
xor U49203 (N_49203,N_41291,N_40928);
and U49204 (N_49204,N_43008,N_41201);
or U49205 (N_49205,N_40929,N_44098);
nor U49206 (N_49206,N_44755,N_44494);
nor U49207 (N_49207,N_41441,N_43297);
nand U49208 (N_49208,N_42432,N_41939);
nand U49209 (N_49209,N_41823,N_40154);
nand U49210 (N_49210,N_40925,N_40183);
and U49211 (N_49211,N_42750,N_42904);
and U49212 (N_49212,N_40229,N_40966);
and U49213 (N_49213,N_43952,N_41313);
nand U49214 (N_49214,N_43590,N_44252);
nand U49215 (N_49215,N_42343,N_42332);
and U49216 (N_49216,N_43249,N_41802);
or U49217 (N_49217,N_42345,N_42602);
or U49218 (N_49218,N_42563,N_44676);
xor U49219 (N_49219,N_40099,N_42633);
and U49220 (N_49220,N_42436,N_43681);
xnor U49221 (N_49221,N_43980,N_40114);
and U49222 (N_49222,N_40041,N_42387);
or U49223 (N_49223,N_44691,N_42911);
and U49224 (N_49224,N_44949,N_41605);
or U49225 (N_49225,N_41408,N_40583);
or U49226 (N_49226,N_40158,N_41005);
and U49227 (N_49227,N_40630,N_44250);
or U49228 (N_49228,N_42128,N_41106);
and U49229 (N_49229,N_42923,N_41524);
nor U49230 (N_49230,N_43124,N_42975);
and U49231 (N_49231,N_43541,N_40523);
and U49232 (N_49232,N_43175,N_40034);
xnor U49233 (N_49233,N_42713,N_43450);
nand U49234 (N_49234,N_41078,N_42948);
or U49235 (N_49235,N_43990,N_44309);
nor U49236 (N_49236,N_41957,N_42192);
and U49237 (N_49237,N_42874,N_41957);
nand U49238 (N_49238,N_42913,N_40884);
and U49239 (N_49239,N_44829,N_42662);
nand U49240 (N_49240,N_43613,N_44038);
nor U49241 (N_49241,N_40466,N_44734);
xor U49242 (N_49242,N_44260,N_44537);
or U49243 (N_49243,N_42632,N_42553);
nor U49244 (N_49244,N_42362,N_41221);
nand U49245 (N_49245,N_42945,N_43260);
nand U49246 (N_49246,N_42632,N_41757);
xnor U49247 (N_49247,N_42012,N_41713);
nand U49248 (N_49248,N_44407,N_42885);
xor U49249 (N_49249,N_40757,N_42293);
nand U49250 (N_49250,N_40521,N_40694);
and U49251 (N_49251,N_41809,N_41630);
or U49252 (N_49252,N_41616,N_42082);
xnor U49253 (N_49253,N_41885,N_43631);
and U49254 (N_49254,N_44149,N_41378);
and U49255 (N_49255,N_40093,N_41836);
nor U49256 (N_49256,N_43010,N_43428);
xor U49257 (N_49257,N_40380,N_42507);
xor U49258 (N_49258,N_42615,N_44327);
xnor U49259 (N_49259,N_44242,N_41513);
nand U49260 (N_49260,N_42963,N_40589);
xnor U49261 (N_49261,N_44147,N_40078);
nand U49262 (N_49262,N_44788,N_44598);
or U49263 (N_49263,N_41324,N_43736);
xnor U49264 (N_49264,N_40110,N_44776);
xnor U49265 (N_49265,N_41840,N_40790);
xor U49266 (N_49266,N_42700,N_41421);
nand U49267 (N_49267,N_42049,N_43891);
xor U49268 (N_49268,N_42134,N_44665);
nand U49269 (N_49269,N_43545,N_44759);
nor U49270 (N_49270,N_41344,N_40309);
xor U49271 (N_49271,N_40379,N_41003);
nand U49272 (N_49272,N_40826,N_41861);
xnor U49273 (N_49273,N_40333,N_44790);
xor U49274 (N_49274,N_41332,N_41824);
nor U49275 (N_49275,N_43077,N_44809);
xnor U49276 (N_49276,N_40430,N_42320);
and U49277 (N_49277,N_43173,N_40338);
nand U49278 (N_49278,N_43144,N_40941);
xnor U49279 (N_49279,N_42769,N_41745);
nand U49280 (N_49280,N_43703,N_42668);
nand U49281 (N_49281,N_40047,N_41057);
nor U49282 (N_49282,N_41423,N_44017);
and U49283 (N_49283,N_42552,N_41360);
and U49284 (N_49284,N_41163,N_42523);
xnor U49285 (N_49285,N_40008,N_43061);
and U49286 (N_49286,N_44147,N_43292);
and U49287 (N_49287,N_44891,N_41012);
and U49288 (N_49288,N_43322,N_41971);
nand U49289 (N_49289,N_42930,N_40172);
and U49290 (N_49290,N_40247,N_42233);
and U49291 (N_49291,N_42202,N_44313);
and U49292 (N_49292,N_42222,N_44799);
xor U49293 (N_49293,N_44443,N_40568);
nor U49294 (N_49294,N_42508,N_43330);
nor U49295 (N_49295,N_42401,N_44408);
xnor U49296 (N_49296,N_41452,N_40084);
nor U49297 (N_49297,N_40249,N_42559);
and U49298 (N_49298,N_44940,N_42128);
nor U49299 (N_49299,N_41397,N_44590);
or U49300 (N_49300,N_40533,N_42608);
xnor U49301 (N_49301,N_43578,N_41704);
xor U49302 (N_49302,N_43027,N_40065);
nor U49303 (N_49303,N_41445,N_41758);
nand U49304 (N_49304,N_41147,N_44793);
or U49305 (N_49305,N_42203,N_40302);
and U49306 (N_49306,N_40152,N_43951);
or U49307 (N_49307,N_40738,N_41068);
xnor U49308 (N_49308,N_43645,N_40959);
or U49309 (N_49309,N_40617,N_41171);
xor U49310 (N_49310,N_42194,N_44227);
xnor U49311 (N_49311,N_43430,N_44363);
nor U49312 (N_49312,N_44032,N_43200);
or U49313 (N_49313,N_40688,N_40669);
nor U49314 (N_49314,N_40823,N_40309);
nor U49315 (N_49315,N_42591,N_42813);
or U49316 (N_49316,N_43403,N_43284);
xor U49317 (N_49317,N_40522,N_44669);
xnor U49318 (N_49318,N_44313,N_40158);
or U49319 (N_49319,N_41742,N_40919);
nand U49320 (N_49320,N_44544,N_41003);
nand U49321 (N_49321,N_42976,N_41344);
and U49322 (N_49322,N_42978,N_44533);
nor U49323 (N_49323,N_42575,N_40608);
and U49324 (N_49324,N_43695,N_41355);
nor U49325 (N_49325,N_42234,N_44457);
xor U49326 (N_49326,N_41337,N_44183);
or U49327 (N_49327,N_40165,N_43469);
and U49328 (N_49328,N_44454,N_40830);
nand U49329 (N_49329,N_42904,N_44131);
nor U49330 (N_49330,N_40026,N_42269);
and U49331 (N_49331,N_42312,N_43459);
nor U49332 (N_49332,N_42138,N_40411);
or U49333 (N_49333,N_41205,N_41190);
and U49334 (N_49334,N_41294,N_43681);
or U49335 (N_49335,N_42431,N_41820);
nand U49336 (N_49336,N_44675,N_42251);
nand U49337 (N_49337,N_44887,N_44759);
or U49338 (N_49338,N_40487,N_40966);
or U49339 (N_49339,N_42394,N_40532);
or U49340 (N_49340,N_41143,N_42872);
xor U49341 (N_49341,N_43442,N_40448);
or U49342 (N_49342,N_40079,N_40167);
xor U49343 (N_49343,N_44335,N_43145);
nand U49344 (N_49344,N_41118,N_41475);
or U49345 (N_49345,N_44695,N_41862);
and U49346 (N_49346,N_41347,N_41827);
nand U49347 (N_49347,N_44264,N_44173);
xnor U49348 (N_49348,N_43223,N_40989);
nand U49349 (N_49349,N_42795,N_42210);
and U49350 (N_49350,N_43246,N_43925);
or U49351 (N_49351,N_40168,N_41923);
nand U49352 (N_49352,N_44781,N_44842);
or U49353 (N_49353,N_42053,N_40286);
or U49354 (N_49354,N_42003,N_43276);
xnor U49355 (N_49355,N_43242,N_41072);
nand U49356 (N_49356,N_41332,N_41908);
nand U49357 (N_49357,N_40126,N_43149);
or U49358 (N_49358,N_43227,N_44942);
or U49359 (N_49359,N_44787,N_42453);
nand U49360 (N_49360,N_42349,N_42884);
nor U49361 (N_49361,N_44508,N_42125);
or U49362 (N_49362,N_42112,N_44031);
or U49363 (N_49363,N_41530,N_44339);
xor U49364 (N_49364,N_40040,N_43473);
and U49365 (N_49365,N_40128,N_44149);
or U49366 (N_49366,N_43927,N_43215);
nor U49367 (N_49367,N_42077,N_40556);
and U49368 (N_49368,N_44837,N_41330);
and U49369 (N_49369,N_43593,N_44359);
and U49370 (N_49370,N_40735,N_40000);
or U49371 (N_49371,N_40268,N_40142);
or U49372 (N_49372,N_44709,N_41902);
and U49373 (N_49373,N_41598,N_43307);
or U49374 (N_49374,N_42762,N_41818);
nor U49375 (N_49375,N_41886,N_43599);
and U49376 (N_49376,N_44259,N_43327);
or U49377 (N_49377,N_40062,N_41259);
nor U49378 (N_49378,N_43540,N_41331);
and U49379 (N_49379,N_44725,N_44156);
nor U49380 (N_49380,N_40531,N_40017);
or U49381 (N_49381,N_40296,N_44254);
nand U49382 (N_49382,N_41940,N_41314);
or U49383 (N_49383,N_41697,N_42666);
nand U49384 (N_49384,N_44191,N_40938);
and U49385 (N_49385,N_44207,N_41581);
or U49386 (N_49386,N_44970,N_42188);
nor U49387 (N_49387,N_42200,N_43929);
nand U49388 (N_49388,N_40218,N_41202);
xnor U49389 (N_49389,N_42487,N_41746);
nor U49390 (N_49390,N_40574,N_43866);
xnor U49391 (N_49391,N_44051,N_40598);
nor U49392 (N_49392,N_43170,N_42389);
nor U49393 (N_49393,N_41805,N_42012);
nor U49394 (N_49394,N_41325,N_41437);
xor U49395 (N_49395,N_44343,N_43066);
nor U49396 (N_49396,N_44789,N_41727);
nor U49397 (N_49397,N_43867,N_41508);
xor U49398 (N_49398,N_40103,N_40828);
or U49399 (N_49399,N_44798,N_43282);
nor U49400 (N_49400,N_42187,N_44584);
nand U49401 (N_49401,N_43420,N_44085);
nand U49402 (N_49402,N_43625,N_40602);
and U49403 (N_49403,N_44678,N_44851);
or U49404 (N_49404,N_44302,N_43784);
or U49405 (N_49405,N_41210,N_44195);
and U49406 (N_49406,N_42849,N_42958);
or U49407 (N_49407,N_41109,N_44626);
nor U49408 (N_49408,N_44546,N_41954);
xnor U49409 (N_49409,N_41201,N_40063);
and U49410 (N_49410,N_42060,N_40087);
xnor U49411 (N_49411,N_43769,N_40470);
nor U49412 (N_49412,N_43965,N_41018);
xor U49413 (N_49413,N_41400,N_42190);
nor U49414 (N_49414,N_42472,N_40258);
or U49415 (N_49415,N_41181,N_42273);
and U49416 (N_49416,N_42734,N_40515);
nor U49417 (N_49417,N_40939,N_41360);
nand U49418 (N_49418,N_44087,N_40191);
nand U49419 (N_49419,N_44464,N_40718);
and U49420 (N_49420,N_42734,N_44586);
nand U49421 (N_49421,N_42147,N_43654);
nand U49422 (N_49422,N_40760,N_44829);
or U49423 (N_49423,N_43352,N_42731);
xor U49424 (N_49424,N_42685,N_41605);
xor U49425 (N_49425,N_41688,N_43214);
nor U49426 (N_49426,N_44548,N_41948);
or U49427 (N_49427,N_41824,N_43536);
xnor U49428 (N_49428,N_41072,N_40266);
nor U49429 (N_49429,N_43303,N_44423);
nand U49430 (N_49430,N_43558,N_42377);
nand U49431 (N_49431,N_40617,N_44947);
or U49432 (N_49432,N_41145,N_41749);
nor U49433 (N_49433,N_40976,N_43761);
nor U49434 (N_49434,N_43137,N_43521);
or U49435 (N_49435,N_42479,N_41201);
nand U49436 (N_49436,N_42229,N_40684);
nor U49437 (N_49437,N_44130,N_40314);
nor U49438 (N_49438,N_43996,N_42805);
xor U49439 (N_49439,N_40789,N_43146);
xnor U49440 (N_49440,N_42660,N_41118);
and U49441 (N_49441,N_42761,N_44457);
and U49442 (N_49442,N_42770,N_41173);
nor U49443 (N_49443,N_42479,N_44946);
xnor U49444 (N_49444,N_41510,N_40683);
nand U49445 (N_49445,N_44484,N_43839);
xnor U49446 (N_49446,N_43709,N_44729);
xor U49447 (N_49447,N_40361,N_44116);
xor U49448 (N_49448,N_44883,N_42531);
xor U49449 (N_49449,N_41390,N_42967);
or U49450 (N_49450,N_41035,N_43786);
nand U49451 (N_49451,N_43680,N_43314);
nor U49452 (N_49452,N_43011,N_44032);
nand U49453 (N_49453,N_42021,N_44994);
nor U49454 (N_49454,N_44274,N_44884);
xnor U49455 (N_49455,N_42828,N_42041);
nand U49456 (N_49456,N_40512,N_41300);
or U49457 (N_49457,N_40613,N_44994);
xor U49458 (N_49458,N_44942,N_43649);
or U49459 (N_49459,N_42838,N_43737);
or U49460 (N_49460,N_44661,N_43971);
and U49461 (N_49461,N_43996,N_41420);
xnor U49462 (N_49462,N_41403,N_40141);
xor U49463 (N_49463,N_43249,N_40567);
and U49464 (N_49464,N_44471,N_41210);
and U49465 (N_49465,N_43677,N_42696);
or U49466 (N_49466,N_41907,N_41852);
or U49467 (N_49467,N_40450,N_43720);
or U49468 (N_49468,N_43760,N_41679);
nand U49469 (N_49469,N_40638,N_40919);
and U49470 (N_49470,N_44670,N_43133);
and U49471 (N_49471,N_40675,N_43170);
nor U49472 (N_49472,N_41723,N_44642);
or U49473 (N_49473,N_44643,N_42050);
xnor U49474 (N_49474,N_41486,N_44560);
or U49475 (N_49475,N_41864,N_44689);
and U49476 (N_49476,N_42304,N_44724);
nor U49477 (N_49477,N_41920,N_44162);
nor U49478 (N_49478,N_41004,N_40744);
nand U49479 (N_49479,N_41966,N_40548);
and U49480 (N_49480,N_42498,N_42715);
nand U49481 (N_49481,N_42578,N_41173);
and U49482 (N_49482,N_40610,N_42540);
and U49483 (N_49483,N_43755,N_41823);
nand U49484 (N_49484,N_40183,N_40097);
nor U49485 (N_49485,N_40473,N_43219);
and U49486 (N_49486,N_42313,N_43094);
or U49487 (N_49487,N_41746,N_41925);
nand U49488 (N_49488,N_44509,N_40446);
nand U49489 (N_49489,N_40905,N_44562);
nor U49490 (N_49490,N_40537,N_44259);
and U49491 (N_49491,N_44725,N_42321);
nor U49492 (N_49492,N_44210,N_44533);
nor U49493 (N_49493,N_42921,N_43688);
xor U49494 (N_49494,N_42421,N_43720);
or U49495 (N_49495,N_42726,N_41212);
nand U49496 (N_49496,N_41786,N_44120);
nor U49497 (N_49497,N_42148,N_40897);
xnor U49498 (N_49498,N_44202,N_40769);
and U49499 (N_49499,N_42774,N_44214);
or U49500 (N_49500,N_41166,N_43187);
nand U49501 (N_49501,N_40391,N_42988);
nor U49502 (N_49502,N_41384,N_42386);
and U49503 (N_49503,N_40895,N_44019);
xnor U49504 (N_49504,N_40906,N_41225);
nor U49505 (N_49505,N_42318,N_41277);
nor U49506 (N_49506,N_43184,N_41154);
xnor U49507 (N_49507,N_44545,N_44681);
xnor U49508 (N_49508,N_41040,N_44677);
nor U49509 (N_49509,N_42663,N_44806);
or U49510 (N_49510,N_44948,N_40374);
nand U49511 (N_49511,N_40416,N_43973);
nand U49512 (N_49512,N_41736,N_43311);
xnor U49513 (N_49513,N_42911,N_42697);
or U49514 (N_49514,N_40073,N_43428);
nor U49515 (N_49515,N_43055,N_41310);
or U49516 (N_49516,N_41778,N_42531);
nand U49517 (N_49517,N_40277,N_44722);
and U49518 (N_49518,N_42487,N_41665);
nand U49519 (N_49519,N_41254,N_44584);
or U49520 (N_49520,N_44261,N_41418);
xor U49521 (N_49521,N_42211,N_40868);
nand U49522 (N_49522,N_44035,N_40130);
nand U49523 (N_49523,N_40917,N_40850);
nand U49524 (N_49524,N_43242,N_41609);
nand U49525 (N_49525,N_41445,N_42327);
nand U49526 (N_49526,N_42531,N_42398);
nor U49527 (N_49527,N_41663,N_40072);
nor U49528 (N_49528,N_44949,N_44094);
nand U49529 (N_49529,N_43988,N_40075);
and U49530 (N_49530,N_42633,N_42197);
nor U49531 (N_49531,N_43361,N_41639);
nand U49532 (N_49532,N_42568,N_40469);
or U49533 (N_49533,N_42702,N_41563);
nand U49534 (N_49534,N_42951,N_43306);
xor U49535 (N_49535,N_44435,N_43122);
nand U49536 (N_49536,N_41365,N_44710);
or U49537 (N_49537,N_44342,N_44788);
or U49538 (N_49538,N_42082,N_40645);
nor U49539 (N_49539,N_44627,N_41335);
and U49540 (N_49540,N_44530,N_44752);
nand U49541 (N_49541,N_42143,N_42396);
and U49542 (N_49542,N_40946,N_43910);
nor U49543 (N_49543,N_43025,N_44398);
and U49544 (N_49544,N_40413,N_41115);
or U49545 (N_49545,N_41843,N_40308);
xor U49546 (N_49546,N_41542,N_40045);
nand U49547 (N_49547,N_41086,N_44171);
xor U49548 (N_49548,N_41436,N_44485);
nor U49549 (N_49549,N_42175,N_42896);
or U49550 (N_49550,N_41361,N_44485);
and U49551 (N_49551,N_42853,N_44056);
or U49552 (N_49552,N_40233,N_42867);
nor U49553 (N_49553,N_41077,N_42475);
nor U49554 (N_49554,N_40137,N_43804);
xor U49555 (N_49555,N_44743,N_40468);
nor U49556 (N_49556,N_40319,N_42922);
or U49557 (N_49557,N_42895,N_44652);
xor U49558 (N_49558,N_41653,N_44948);
nor U49559 (N_49559,N_44178,N_44786);
xor U49560 (N_49560,N_42423,N_42146);
or U49561 (N_49561,N_42279,N_41824);
or U49562 (N_49562,N_43178,N_42054);
and U49563 (N_49563,N_44862,N_40929);
nand U49564 (N_49564,N_43610,N_40271);
xor U49565 (N_49565,N_41228,N_43936);
nand U49566 (N_49566,N_42190,N_42613);
xnor U49567 (N_49567,N_44040,N_44016);
nor U49568 (N_49568,N_42335,N_41877);
and U49569 (N_49569,N_42471,N_44715);
or U49570 (N_49570,N_40891,N_42154);
nand U49571 (N_49571,N_43290,N_43805);
nand U49572 (N_49572,N_43130,N_42543);
or U49573 (N_49573,N_44578,N_44362);
xnor U49574 (N_49574,N_44341,N_41371);
nand U49575 (N_49575,N_44899,N_44676);
nor U49576 (N_49576,N_44916,N_41605);
and U49577 (N_49577,N_42455,N_42898);
and U49578 (N_49578,N_44068,N_42167);
nand U49579 (N_49579,N_43360,N_41829);
and U49580 (N_49580,N_43049,N_43604);
nor U49581 (N_49581,N_43878,N_40679);
nor U49582 (N_49582,N_41560,N_44054);
nor U49583 (N_49583,N_40331,N_44685);
nand U49584 (N_49584,N_41521,N_41937);
xor U49585 (N_49585,N_41894,N_42987);
or U49586 (N_49586,N_43597,N_44431);
nand U49587 (N_49587,N_41603,N_40675);
and U49588 (N_49588,N_40079,N_42304);
and U49589 (N_49589,N_43728,N_41203);
and U49590 (N_49590,N_41066,N_43599);
or U49591 (N_49591,N_42080,N_43724);
nand U49592 (N_49592,N_44292,N_40730);
nand U49593 (N_49593,N_44066,N_40428);
nand U49594 (N_49594,N_43183,N_44291);
nand U49595 (N_49595,N_43907,N_42027);
nand U49596 (N_49596,N_43885,N_40829);
xor U49597 (N_49597,N_40364,N_44907);
nor U49598 (N_49598,N_43432,N_40690);
and U49599 (N_49599,N_43607,N_41056);
xnor U49600 (N_49600,N_44022,N_42762);
nor U49601 (N_49601,N_41661,N_43424);
xor U49602 (N_49602,N_43750,N_42204);
nand U49603 (N_49603,N_42787,N_44874);
nor U49604 (N_49604,N_41878,N_40359);
or U49605 (N_49605,N_44688,N_43532);
and U49606 (N_49606,N_44254,N_44773);
nor U49607 (N_49607,N_44723,N_43635);
nand U49608 (N_49608,N_43094,N_43665);
xor U49609 (N_49609,N_40526,N_41545);
nor U49610 (N_49610,N_41575,N_41099);
or U49611 (N_49611,N_43970,N_42932);
and U49612 (N_49612,N_40541,N_44410);
and U49613 (N_49613,N_40238,N_42842);
or U49614 (N_49614,N_40652,N_42846);
or U49615 (N_49615,N_42215,N_44296);
xor U49616 (N_49616,N_42038,N_40601);
nand U49617 (N_49617,N_42436,N_43398);
nand U49618 (N_49618,N_41702,N_44359);
nand U49619 (N_49619,N_44098,N_42675);
or U49620 (N_49620,N_41088,N_43908);
nand U49621 (N_49621,N_41507,N_40591);
xor U49622 (N_49622,N_41175,N_44326);
and U49623 (N_49623,N_44718,N_42958);
nor U49624 (N_49624,N_42866,N_41186);
nand U49625 (N_49625,N_43149,N_40332);
nor U49626 (N_49626,N_40879,N_40617);
xnor U49627 (N_49627,N_43620,N_40326);
or U49628 (N_49628,N_42186,N_43105);
nand U49629 (N_49629,N_42962,N_41639);
or U49630 (N_49630,N_41645,N_40214);
nor U49631 (N_49631,N_41708,N_41328);
and U49632 (N_49632,N_42858,N_40810);
or U49633 (N_49633,N_43670,N_42746);
or U49634 (N_49634,N_43762,N_42306);
nand U49635 (N_49635,N_40255,N_42242);
nand U49636 (N_49636,N_44079,N_41566);
xnor U49637 (N_49637,N_42502,N_44290);
nor U49638 (N_49638,N_40538,N_44834);
nor U49639 (N_49639,N_42659,N_44723);
or U49640 (N_49640,N_42897,N_43867);
nand U49641 (N_49641,N_41014,N_40306);
and U49642 (N_49642,N_41412,N_44878);
nor U49643 (N_49643,N_43875,N_40447);
and U49644 (N_49644,N_42115,N_41271);
nand U49645 (N_49645,N_41931,N_42222);
xor U49646 (N_49646,N_44574,N_44130);
nor U49647 (N_49647,N_41137,N_41722);
and U49648 (N_49648,N_40413,N_42035);
nor U49649 (N_49649,N_41259,N_44025);
nor U49650 (N_49650,N_43538,N_41710);
xor U49651 (N_49651,N_42596,N_44134);
nor U49652 (N_49652,N_43988,N_43602);
or U49653 (N_49653,N_44867,N_41154);
nor U49654 (N_49654,N_43578,N_43982);
and U49655 (N_49655,N_44472,N_44576);
xnor U49656 (N_49656,N_44414,N_43208);
and U49657 (N_49657,N_41470,N_41113);
xor U49658 (N_49658,N_40878,N_44994);
xor U49659 (N_49659,N_42386,N_43559);
nor U49660 (N_49660,N_41576,N_43426);
nor U49661 (N_49661,N_42230,N_40024);
nand U49662 (N_49662,N_44296,N_44374);
nor U49663 (N_49663,N_41910,N_40826);
nand U49664 (N_49664,N_43137,N_41168);
xnor U49665 (N_49665,N_43895,N_42265);
or U49666 (N_49666,N_42126,N_44565);
and U49667 (N_49667,N_42929,N_44131);
nor U49668 (N_49668,N_43016,N_40429);
nor U49669 (N_49669,N_40292,N_43259);
or U49670 (N_49670,N_42724,N_42008);
and U49671 (N_49671,N_40949,N_43466);
and U49672 (N_49672,N_43564,N_44352);
nor U49673 (N_49673,N_43672,N_44425);
nand U49674 (N_49674,N_44236,N_44125);
nand U49675 (N_49675,N_42821,N_42784);
nor U49676 (N_49676,N_43428,N_40693);
and U49677 (N_49677,N_41902,N_42251);
and U49678 (N_49678,N_41033,N_44837);
or U49679 (N_49679,N_40533,N_44442);
nand U49680 (N_49680,N_43697,N_40615);
or U49681 (N_49681,N_43857,N_43437);
and U49682 (N_49682,N_42398,N_41441);
and U49683 (N_49683,N_40215,N_42438);
nor U49684 (N_49684,N_43298,N_43235);
and U49685 (N_49685,N_44442,N_42438);
or U49686 (N_49686,N_42037,N_42294);
or U49687 (N_49687,N_41715,N_44647);
xor U49688 (N_49688,N_41666,N_40274);
nand U49689 (N_49689,N_42614,N_42655);
nor U49690 (N_49690,N_42403,N_43492);
xor U49691 (N_49691,N_41577,N_43661);
xnor U49692 (N_49692,N_40652,N_43449);
xor U49693 (N_49693,N_43001,N_40124);
or U49694 (N_49694,N_42080,N_41623);
and U49695 (N_49695,N_41972,N_43936);
nand U49696 (N_49696,N_40986,N_41746);
or U49697 (N_49697,N_40539,N_43043);
nor U49698 (N_49698,N_42412,N_43428);
or U49699 (N_49699,N_40757,N_43341);
nor U49700 (N_49700,N_44193,N_41554);
nand U49701 (N_49701,N_40467,N_40048);
xnor U49702 (N_49702,N_42405,N_43898);
nand U49703 (N_49703,N_44935,N_43894);
or U49704 (N_49704,N_43966,N_41848);
nor U49705 (N_49705,N_40379,N_44518);
xor U49706 (N_49706,N_42145,N_40255);
or U49707 (N_49707,N_42168,N_42837);
and U49708 (N_49708,N_42593,N_42251);
nand U49709 (N_49709,N_42188,N_40055);
nor U49710 (N_49710,N_43261,N_40153);
nor U49711 (N_49711,N_43072,N_44160);
xnor U49712 (N_49712,N_41767,N_42392);
and U49713 (N_49713,N_42105,N_44089);
and U49714 (N_49714,N_42400,N_44722);
and U49715 (N_49715,N_42533,N_43117);
and U49716 (N_49716,N_44023,N_41780);
nand U49717 (N_49717,N_44084,N_43455);
xor U49718 (N_49718,N_42918,N_40458);
nand U49719 (N_49719,N_43668,N_43960);
or U49720 (N_49720,N_42301,N_44677);
nor U49721 (N_49721,N_42536,N_43428);
or U49722 (N_49722,N_44020,N_43586);
and U49723 (N_49723,N_43406,N_44454);
nand U49724 (N_49724,N_40885,N_40052);
and U49725 (N_49725,N_41121,N_43960);
nor U49726 (N_49726,N_42660,N_40724);
nor U49727 (N_49727,N_44504,N_43264);
or U49728 (N_49728,N_41302,N_41597);
or U49729 (N_49729,N_40827,N_41527);
and U49730 (N_49730,N_40959,N_44820);
nor U49731 (N_49731,N_41227,N_42815);
xor U49732 (N_49732,N_44838,N_40101);
and U49733 (N_49733,N_44980,N_41993);
xnor U49734 (N_49734,N_40535,N_43580);
nor U49735 (N_49735,N_41989,N_43020);
xnor U49736 (N_49736,N_40637,N_44716);
nor U49737 (N_49737,N_41677,N_41037);
and U49738 (N_49738,N_41309,N_40823);
nor U49739 (N_49739,N_42567,N_43498);
and U49740 (N_49740,N_40199,N_40121);
or U49741 (N_49741,N_41432,N_42243);
nand U49742 (N_49742,N_44160,N_44377);
and U49743 (N_49743,N_42873,N_42154);
nand U49744 (N_49744,N_40299,N_44436);
xnor U49745 (N_49745,N_43528,N_40093);
and U49746 (N_49746,N_44143,N_43480);
nor U49747 (N_49747,N_41041,N_44152);
nor U49748 (N_49748,N_43368,N_41336);
or U49749 (N_49749,N_42530,N_40153);
and U49750 (N_49750,N_43977,N_43720);
nand U49751 (N_49751,N_40225,N_43023);
or U49752 (N_49752,N_41024,N_40193);
nand U49753 (N_49753,N_40073,N_40559);
and U49754 (N_49754,N_40180,N_44645);
xor U49755 (N_49755,N_41077,N_41513);
nand U49756 (N_49756,N_40098,N_41713);
nand U49757 (N_49757,N_40767,N_42100);
nor U49758 (N_49758,N_42007,N_44535);
nand U49759 (N_49759,N_44645,N_44556);
xnor U49760 (N_49760,N_42863,N_44691);
and U49761 (N_49761,N_40779,N_44922);
nand U49762 (N_49762,N_43586,N_41073);
nand U49763 (N_49763,N_44159,N_41171);
xnor U49764 (N_49764,N_44413,N_40759);
nor U49765 (N_49765,N_43774,N_42054);
nand U49766 (N_49766,N_43626,N_43562);
nand U49767 (N_49767,N_40165,N_42830);
nand U49768 (N_49768,N_41142,N_44172);
and U49769 (N_49769,N_44826,N_44853);
nand U49770 (N_49770,N_42016,N_41925);
nor U49771 (N_49771,N_44002,N_44223);
and U49772 (N_49772,N_41230,N_40176);
and U49773 (N_49773,N_43315,N_44979);
nor U49774 (N_49774,N_40599,N_40474);
or U49775 (N_49775,N_42485,N_41106);
nor U49776 (N_49776,N_44103,N_43923);
nand U49777 (N_49777,N_40284,N_43784);
nand U49778 (N_49778,N_43132,N_42236);
or U49779 (N_49779,N_42247,N_41278);
nand U49780 (N_49780,N_40621,N_42271);
nand U49781 (N_49781,N_40416,N_43987);
nor U49782 (N_49782,N_42535,N_43570);
and U49783 (N_49783,N_43278,N_40602);
xnor U49784 (N_49784,N_42903,N_40954);
or U49785 (N_49785,N_42325,N_40521);
or U49786 (N_49786,N_41357,N_40400);
or U49787 (N_49787,N_44105,N_40979);
and U49788 (N_49788,N_40132,N_44933);
xnor U49789 (N_49789,N_44632,N_43734);
nor U49790 (N_49790,N_44265,N_40488);
xor U49791 (N_49791,N_41345,N_44343);
nand U49792 (N_49792,N_44475,N_42348);
nor U49793 (N_49793,N_42148,N_44080);
and U49794 (N_49794,N_42597,N_42814);
xnor U49795 (N_49795,N_42292,N_44034);
nand U49796 (N_49796,N_44593,N_42479);
or U49797 (N_49797,N_42468,N_41175);
xor U49798 (N_49798,N_43274,N_41473);
or U49799 (N_49799,N_40360,N_43614);
nand U49800 (N_49800,N_40683,N_42416);
and U49801 (N_49801,N_41003,N_40723);
xnor U49802 (N_49802,N_40114,N_40258);
or U49803 (N_49803,N_42367,N_43962);
nand U49804 (N_49804,N_40209,N_41724);
or U49805 (N_49805,N_43369,N_40776);
nor U49806 (N_49806,N_43984,N_40021);
and U49807 (N_49807,N_42793,N_44825);
xnor U49808 (N_49808,N_40402,N_44196);
and U49809 (N_49809,N_41934,N_40276);
nand U49810 (N_49810,N_44487,N_42582);
or U49811 (N_49811,N_40376,N_42299);
xor U49812 (N_49812,N_41246,N_40870);
nor U49813 (N_49813,N_41434,N_40001);
nor U49814 (N_49814,N_43728,N_42790);
nand U49815 (N_49815,N_44927,N_42522);
or U49816 (N_49816,N_42782,N_40428);
nand U49817 (N_49817,N_41712,N_41470);
xnor U49818 (N_49818,N_41940,N_43467);
nand U49819 (N_49819,N_43993,N_40035);
or U49820 (N_49820,N_44245,N_41546);
and U49821 (N_49821,N_44006,N_41528);
and U49822 (N_49822,N_43959,N_42043);
or U49823 (N_49823,N_42904,N_41945);
or U49824 (N_49824,N_41365,N_42423);
xor U49825 (N_49825,N_41204,N_44404);
nor U49826 (N_49826,N_42149,N_42845);
nand U49827 (N_49827,N_43284,N_40891);
xor U49828 (N_49828,N_40674,N_42107);
nor U49829 (N_49829,N_44173,N_40178);
xor U49830 (N_49830,N_42260,N_43536);
or U49831 (N_49831,N_42367,N_41869);
or U49832 (N_49832,N_41557,N_40595);
nor U49833 (N_49833,N_41872,N_44698);
xnor U49834 (N_49834,N_41345,N_42997);
or U49835 (N_49835,N_41501,N_41566);
nand U49836 (N_49836,N_43932,N_42614);
or U49837 (N_49837,N_40222,N_42394);
or U49838 (N_49838,N_41887,N_42346);
xor U49839 (N_49839,N_41738,N_44365);
xnor U49840 (N_49840,N_42022,N_44289);
nor U49841 (N_49841,N_44613,N_42491);
and U49842 (N_49842,N_40299,N_42264);
or U49843 (N_49843,N_43289,N_43454);
xnor U49844 (N_49844,N_40166,N_44364);
nor U49845 (N_49845,N_41954,N_40314);
and U49846 (N_49846,N_44775,N_41079);
nand U49847 (N_49847,N_43496,N_40250);
or U49848 (N_49848,N_40673,N_43667);
xor U49849 (N_49849,N_44470,N_41609);
or U49850 (N_49850,N_40868,N_42392);
and U49851 (N_49851,N_42357,N_44453);
xor U49852 (N_49852,N_42807,N_43537);
or U49853 (N_49853,N_41596,N_43076);
and U49854 (N_49854,N_44656,N_44622);
nand U49855 (N_49855,N_43882,N_42955);
and U49856 (N_49856,N_44096,N_44327);
xnor U49857 (N_49857,N_44831,N_43038);
xor U49858 (N_49858,N_41796,N_41261);
nor U49859 (N_49859,N_44822,N_40535);
or U49860 (N_49860,N_41532,N_42437);
nor U49861 (N_49861,N_42308,N_42791);
nand U49862 (N_49862,N_41663,N_41504);
nor U49863 (N_49863,N_42230,N_41913);
and U49864 (N_49864,N_44199,N_40898);
nand U49865 (N_49865,N_40717,N_40283);
nand U49866 (N_49866,N_40067,N_43679);
or U49867 (N_49867,N_43674,N_42553);
and U49868 (N_49868,N_42719,N_44059);
and U49869 (N_49869,N_41285,N_42878);
nand U49870 (N_49870,N_40393,N_44136);
xnor U49871 (N_49871,N_43979,N_40326);
or U49872 (N_49872,N_44448,N_40479);
or U49873 (N_49873,N_44522,N_40624);
xnor U49874 (N_49874,N_43519,N_44396);
nor U49875 (N_49875,N_42280,N_43773);
xnor U49876 (N_49876,N_41140,N_44046);
and U49877 (N_49877,N_42091,N_42980);
nand U49878 (N_49878,N_43003,N_40354);
nor U49879 (N_49879,N_43080,N_41038);
xnor U49880 (N_49880,N_41175,N_44754);
or U49881 (N_49881,N_40914,N_44875);
nand U49882 (N_49882,N_43511,N_41892);
nor U49883 (N_49883,N_40534,N_44503);
or U49884 (N_49884,N_43416,N_42750);
or U49885 (N_49885,N_42216,N_42292);
nand U49886 (N_49886,N_42896,N_42176);
xnor U49887 (N_49887,N_40160,N_42164);
xor U49888 (N_49888,N_44387,N_42172);
or U49889 (N_49889,N_40640,N_44096);
nor U49890 (N_49890,N_43318,N_41893);
or U49891 (N_49891,N_43220,N_42485);
xnor U49892 (N_49892,N_44342,N_40425);
nand U49893 (N_49893,N_40456,N_43224);
xor U49894 (N_49894,N_40130,N_40791);
and U49895 (N_49895,N_42925,N_43877);
or U49896 (N_49896,N_43299,N_44010);
nor U49897 (N_49897,N_44465,N_41325);
nand U49898 (N_49898,N_44801,N_42172);
nor U49899 (N_49899,N_41140,N_40377);
and U49900 (N_49900,N_41535,N_44024);
nand U49901 (N_49901,N_42449,N_40284);
nand U49902 (N_49902,N_43493,N_44969);
nand U49903 (N_49903,N_41799,N_43250);
nor U49904 (N_49904,N_40389,N_42021);
nor U49905 (N_49905,N_40600,N_44917);
nor U49906 (N_49906,N_43410,N_42714);
nor U49907 (N_49907,N_43037,N_41511);
xnor U49908 (N_49908,N_44865,N_43875);
and U49909 (N_49909,N_44393,N_44194);
or U49910 (N_49910,N_44073,N_40769);
or U49911 (N_49911,N_42270,N_41214);
or U49912 (N_49912,N_43453,N_40835);
or U49913 (N_49913,N_42543,N_40052);
nand U49914 (N_49914,N_41583,N_43649);
nand U49915 (N_49915,N_40426,N_43549);
and U49916 (N_49916,N_42212,N_43771);
or U49917 (N_49917,N_42812,N_41247);
or U49918 (N_49918,N_40245,N_40439);
nand U49919 (N_49919,N_43390,N_40790);
xnor U49920 (N_49920,N_42445,N_41913);
or U49921 (N_49921,N_44449,N_41937);
nor U49922 (N_49922,N_43988,N_40858);
or U49923 (N_49923,N_41101,N_44892);
nand U49924 (N_49924,N_40445,N_40462);
nor U49925 (N_49925,N_43751,N_41733);
xnor U49926 (N_49926,N_40439,N_40894);
or U49927 (N_49927,N_40029,N_44250);
xor U49928 (N_49928,N_41737,N_43154);
and U49929 (N_49929,N_43841,N_43542);
and U49930 (N_49930,N_43810,N_40527);
xor U49931 (N_49931,N_42097,N_42889);
and U49932 (N_49932,N_41142,N_42098);
and U49933 (N_49933,N_44035,N_42976);
nor U49934 (N_49934,N_42969,N_40224);
nor U49935 (N_49935,N_43423,N_41234);
nor U49936 (N_49936,N_44879,N_43722);
or U49937 (N_49937,N_44386,N_44671);
nand U49938 (N_49938,N_40764,N_41596);
nor U49939 (N_49939,N_40209,N_42044);
or U49940 (N_49940,N_42316,N_42027);
or U49941 (N_49941,N_40065,N_42026);
nand U49942 (N_49942,N_41438,N_40184);
nand U49943 (N_49943,N_42020,N_42958);
or U49944 (N_49944,N_43941,N_42058);
nor U49945 (N_49945,N_41063,N_42894);
and U49946 (N_49946,N_40531,N_44393);
xnor U49947 (N_49947,N_44456,N_42740);
nand U49948 (N_49948,N_43799,N_41936);
nand U49949 (N_49949,N_44213,N_41884);
nor U49950 (N_49950,N_44308,N_42498);
xor U49951 (N_49951,N_42693,N_43791);
or U49952 (N_49952,N_41672,N_43654);
or U49953 (N_49953,N_42354,N_43967);
xnor U49954 (N_49954,N_41670,N_42537);
xor U49955 (N_49955,N_40313,N_43077);
or U49956 (N_49956,N_40660,N_41169);
or U49957 (N_49957,N_43961,N_42954);
xnor U49958 (N_49958,N_44349,N_43167);
nor U49959 (N_49959,N_42082,N_44215);
xnor U49960 (N_49960,N_41721,N_41114);
nor U49961 (N_49961,N_41099,N_40099);
nor U49962 (N_49962,N_44814,N_42149);
xnor U49963 (N_49963,N_43956,N_44003);
xnor U49964 (N_49964,N_44774,N_44430);
nor U49965 (N_49965,N_40431,N_43451);
and U49966 (N_49966,N_43582,N_41181);
xor U49967 (N_49967,N_44030,N_42490);
nor U49968 (N_49968,N_42786,N_41282);
nand U49969 (N_49969,N_43839,N_40960);
and U49970 (N_49970,N_44466,N_42510);
and U49971 (N_49971,N_40416,N_40337);
nor U49972 (N_49972,N_44848,N_43301);
xor U49973 (N_49973,N_43720,N_41384);
nand U49974 (N_49974,N_44364,N_44177);
and U49975 (N_49975,N_40104,N_44994);
nand U49976 (N_49976,N_41299,N_40466);
nor U49977 (N_49977,N_42965,N_44937);
nand U49978 (N_49978,N_44164,N_42961);
or U49979 (N_49979,N_44895,N_44794);
and U49980 (N_49980,N_40736,N_43468);
xnor U49981 (N_49981,N_42137,N_44927);
nand U49982 (N_49982,N_42004,N_41156);
nor U49983 (N_49983,N_42211,N_41155);
xnor U49984 (N_49984,N_42167,N_40207);
xnor U49985 (N_49985,N_42115,N_41421);
nor U49986 (N_49986,N_41930,N_44503);
nor U49987 (N_49987,N_40071,N_41362);
xnor U49988 (N_49988,N_43000,N_42114);
nand U49989 (N_49989,N_44672,N_44967);
xor U49990 (N_49990,N_40043,N_41806);
nand U49991 (N_49991,N_43933,N_44450);
xor U49992 (N_49992,N_42489,N_41997);
or U49993 (N_49993,N_44685,N_43422);
xor U49994 (N_49994,N_44101,N_40800);
nor U49995 (N_49995,N_42498,N_41573);
xnor U49996 (N_49996,N_44358,N_42312);
xnor U49997 (N_49997,N_41891,N_41415);
xnor U49998 (N_49998,N_44804,N_44762);
or U49999 (N_49999,N_41027,N_42897);
and UO_0 (O_0,N_46218,N_47542);
and UO_1 (O_1,N_46236,N_47972);
and UO_2 (O_2,N_47883,N_45378);
or UO_3 (O_3,N_46292,N_49823);
nor UO_4 (O_4,N_48518,N_47073);
or UO_5 (O_5,N_46221,N_49048);
nor UO_6 (O_6,N_49039,N_48822);
xor UO_7 (O_7,N_45922,N_45894);
or UO_8 (O_8,N_47392,N_49782);
nor UO_9 (O_9,N_46954,N_49362);
xor UO_10 (O_10,N_46510,N_46732);
and UO_11 (O_11,N_46868,N_46648);
or UO_12 (O_12,N_45110,N_47534);
xor UO_13 (O_13,N_45301,N_48167);
or UO_14 (O_14,N_49311,N_45565);
xnor UO_15 (O_15,N_49399,N_45929);
nand UO_16 (O_16,N_48444,N_45082);
and UO_17 (O_17,N_46775,N_45850);
and UO_18 (O_18,N_49634,N_46205);
or UO_19 (O_19,N_45830,N_49401);
nor UO_20 (O_20,N_45447,N_45789);
or UO_21 (O_21,N_48891,N_49101);
and UO_22 (O_22,N_49808,N_46386);
nand UO_23 (O_23,N_46610,N_45375);
nand UO_24 (O_24,N_49678,N_45485);
or UO_25 (O_25,N_49174,N_46631);
and UO_26 (O_26,N_46969,N_47094);
and UO_27 (O_27,N_49290,N_49935);
and UO_28 (O_28,N_46837,N_47588);
nand UO_29 (O_29,N_48412,N_49995);
and UO_30 (O_30,N_47430,N_47614);
nor UO_31 (O_31,N_48787,N_46201);
or UO_32 (O_32,N_46663,N_47292);
or UO_33 (O_33,N_46655,N_49377);
nand UO_34 (O_34,N_45801,N_46077);
nor UO_35 (O_35,N_47772,N_45455);
nor UO_36 (O_36,N_45585,N_48343);
or UO_37 (O_37,N_46107,N_45359);
xor UO_38 (O_38,N_45518,N_48575);
and UO_39 (O_39,N_47721,N_49503);
nor UO_40 (O_40,N_47291,N_45824);
xnor UO_41 (O_41,N_46257,N_47113);
nand UO_42 (O_42,N_45078,N_46829);
nor UO_43 (O_43,N_45890,N_45113);
xor UO_44 (O_44,N_49276,N_46030);
nor UO_45 (O_45,N_47598,N_48374);
or UO_46 (O_46,N_45318,N_48869);
nand UO_47 (O_47,N_49599,N_47572);
or UO_48 (O_48,N_49971,N_48665);
nand UO_49 (O_49,N_47606,N_46770);
nor UO_50 (O_50,N_48257,N_45664);
or UO_51 (O_51,N_48661,N_49024);
xor UO_52 (O_52,N_46358,N_46237);
nand UO_53 (O_53,N_49735,N_47499);
xor UO_54 (O_54,N_47160,N_45472);
and UO_55 (O_55,N_47016,N_46822);
xnor UO_56 (O_56,N_49996,N_46842);
and UO_57 (O_57,N_46855,N_45554);
xor UO_58 (O_58,N_46135,N_46017);
nand UO_59 (O_59,N_45845,N_45062);
nor UO_60 (O_60,N_45169,N_46513);
or UO_61 (O_61,N_45813,N_46883);
xnor UO_62 (O_62,N_46724,N_47685);
xnor UO_63 (O_63,N_48692,N_45193);
nand UO_64 (O_64,N_48625,N_47311);
nor UO_65 (O_65,N_46181,N_45796);
or UO_66 (O_66,N_48218,N_46376);
nor UO_67 (O_67,N_45874,N_47293);
nor UO_68 (O_68,N_48835,N_45288);
nor UO_69 (O_69,N_48560,N_48874);
nor UO_70 (O_70,N_45241,N_49451);
or UO_71 (O_71,N_45178,N_46499);
nand UO_72 (O_72,N_47237,N_46688);
xnor UO_73 (O_73,N_46457,N_49711);
xor UO_74 (O_74,N_49908,N_49686);
and UO_75 (O_75,N_46823,N_45903);
nand UO_76 (O_76,N_45885,N_48678);
nand UO_77 (O_77,N_46667,N_47530);
nor UO_78 (O_78,N_46794,N_45423);
nor UO_79 (O_79,N_47624,N_49523);
nor UO_80 (O_80,N_45938,N_48384);
nand UO_81 (O_81,N_45559,N_48759);
or UO_82 (O_82,N_45299,N_45376);
nor UO_83 (O_83,N_49153,N_48839);
xnor UO_84 (O_84,N_48233,N_45791);
nand UO_85 (O_85,N_46032,N_47363);
nand UO_86 (O_86,N_48350,N_45363);
or UO_87 (O_87,N_48573,N_47154);
xnor UO_88 (O_88,N_48349,N_47521);
nor UO_89 (O_89,N_48019,N_47429);
xor UO_90 (O_90,N_48214,N_49616);
xnor UO_91 (O_91,N_47699,N_47440);
nand UO_92 (O_92,N_46361,N_49904);
nand UO_93 (O_93,N_49856,N_48760);
and UO_94 (O_94,N_45228,N_46149);
nand UO_95 (O_95,N_49674,N_48655);
nor UO_96 (O_96,N_49287,N_49506);
and UO_97 (O_97,N_47503,N_49977);
and UO_98 (O_98,N_46113,N_49932);
nor UO_99 (O_99,N_48305,N_46561);
xnor UO_100 (O_100,N_47462,N_49939);
and UO_101 (O_101,N_47826,N_49387);
and UO_102 (O_102,N_47129,N_48878);
nand UO_103 (O_103,N_49901,N_47824);
nand UO_104 (O_104,N_45064,N_46546);
nand UO_105 (O_105,N_45456,N_46338);
nor UO_106 (O_106,N_46023,N_46910);
nor UO_107 (O_107,N_45340,N_46197);
and UO_108 (O_108,N_46179,N_47677);
xor UO_109 (O_109,N_49976,N_49407);
nor UO_110 (O_110,N_47528,N_47726);
nand UO_111 (O_111,N_49345,N_48932);
nor UO_112 (O_112,N_46932,N_46227);
and UO_113 (O_113,N_47642,N_49254);
or UO_114 (O_114,N_47495,N_47807);
nor UO_115 (O_115,N_49860,N_45045);
xnor UO_116 (O_116,N_47885,N_47581);
and UO_117 (O_117,N_47197,N_46702);
and UO_118 (O_118,N_48544,N_49396);
or UO_119 (O_119,N_46613,N_47181);
xnor UO_120 (O_120,N_47746,N_46831);
and UO_121 (O_121,N_49398,N_45943);
nor UO_122 (O_122,N_49405,N_49463);
nand UO_123 (O_123,N_48771,N_45323);
xnor UO_124 (O_124,N_46101,N_46843);
xor UO_125 (O_125,N_46184,N_46176);
xnor UO_126 (O_126,N_49811,N_49741);
and UO_127 (O_127,N_49117,N_47298);
xor UO_128 (O_128,N_46255,N_45616);
or UO_129 (O_129,N_48387,N_49059);
xor UO_130 (O_130,N_48959,N_49304);
nand UO_131 (O_131,N_47285,N_47817);
nand UO_132 (O_132,N_48428,N_45581);
and UO_133 (O_133,N_49491,N_47355);
nor UO_134 (O_134,N_49371,N_46712);
nor UO_135 (O_135,N_49431,N_49184);
or UO_136 (O_136,N_49704,N_46646);
and UO_137 (O_137,N_47156,N_47271);
nand UO_138 (O_138,N_46050,N_47706);
xor UO_139 (O_139,N_49617,N_47587);
or UO_140 (O_140,N_48543,N_46084);
nand UO_141 (O_141,N_46432,N_45727);
and UO_142 (O_142,N_49216,N_46196);
nand UO_143 (O_143,N_47803,N_47133);
or UO_144 (O_144,N_48506,N_46565);
xnor UO_145 (O_145,N_46366,N_48422);
or UO_146 (O_146,N_45511,N_49084);
or UO_147 (O_147,N_48075,N_47489);
or UO_148 (O_148,N_46899,N_48056);
nor UO_149 (O_149,N_46295,N_49979);
and UO_150 (O_150,N_49981,N_47123);
xnor UO_151 (O_151,N_49150,N_48016);
nor UO_152 (O_152,N_45441,N_49676);
nand UO_153 (O_153,N_46389,N_45770);
xor UO_154 (O_154,N_49601,N_48918);
and UO_155 (O_155,N_47928,N_48974);
xnor UO_156 (O_156,N_49945,N_46920);
and UO_157 (O_157,N_45736,N_45923);
or UO_158 (O_158,N_47947,N_47047);
nand UO_159 (O_159,N_49326,N_47012);
nand UO_160 (O_160,N_47681,N_45059);
nor UO_161 (O_161,N_48884,N_45973);
xnor UO_162 (O_162,N_47715,N_49192);
nor UO_163 (O_163,N_49687,N_45865);
xnor UO_164 (O_164,N_48315,N_45075);
nand UO_165 (O_165,N_45729,N_48391);
nand UO_166 (O_166,N_47185,N_47391);
nand UO_167 (O_167,N_47433,N_48729);
nand UO_168 (O_168,N_45704,N_49364);
nand UO_169 (O_169,N_47964,N_49056);
xor UO_170 (O_170,N_45209,N_45802);
xor UO_171 (O_171,N_45927,N_45848);
or UO_172 (O_172,N_49814,N_47860);
and UO_173 (O_173,N_45568,N_48215);
nand UO_174 (O_174,N_46870,N_45852);
and UO_175 (O_175,N_49115,N_46750);
xnor UO_176 (O_176,N_46998,N_48670);
and UO_177 (O_177,N_46460,N_46244);
xnor UO_178 (O_178,N_47060,N_48746);
nand UO_179 (O_179,N_45195,N_48105);
xnor UO_180 (O_180,N_48934,N_49966);
or UO_181 (O_181,N_48631,N_45017);
nor UO_182 (O_182,N_48613,N_47981);
nor UO_183 (O_183,N_45302,N_47401);
or UO_184 (O_184,N_47035,N_49365);
or UO_185 (O_185,N_46015,N_49854);
and UO_186 (O_186,N_49521,N_47805);
nor UO_187 (O_187,N_45250,N_46298);
and UO_188 (O_188,N_45767,N_47457);
and UO_189 (O_189,N_46154,N_46745);
or UO_190 (O_190,N_48364,N_48042);
and UO_191 (O_191,N_49881,N_45679);
and UO_192 (O_192,N_48750,N_45379);
nand UO_193 (O_193,N_45374,N_46497);
xnor UO_194 (O_194,N_45305,N_48170);
nand UO_195 (O_195,N_48534,N_46103);
or UO_196 (O_196,N_47134,N_47646);
nand UO_197 (O_197,N_47762,N_48495);
nand UO_198 (O_198,N_48357,N_46812);
nand UO_199 (O_199,N_49736,N_46375);
or UO_200 (O_200,N_48967,N_46583);
or UO_201 (O_201,N_48273,N_45694);
nor UO_202 (O_202,N_49133,N_48209);
and UO_203 (O_203,N_46264,N_47211);
nand UO_204 (O_204,N_49423,N_45899);
or UO_205 (O_205,N_48720,N_48321);
or UO_206 (O_206,N_45742,N_49961);
or UO_207 (O_207,N_49828,N_47932);
or UO_208 (O_208,N_45454,N_48377);
nor UO_209 (O_209,N_48805,N_48652);
and UO_210 (O_210,N_48980,N_49352);
nor UO_211 (O_211,N_45372,N_48265);
or UO_212 (O_212,N_46765,N_48324);
xnor UO_213 (O_213,N_49170,N_49843);
xor UO_214 (O_214,N_49189,N_48603);
or UO_215 (O_215,N_45598,N_49335);
xor UO_216 (O_216,N_45353,N_49508);
nor UO_217 (O_217,N_47628,N_49889);
and UO_218 (O_218,N_48496,N_47791);
nand UO_219 (O_219,N_46132,N_48614);
nor UO_220 (O_220,N_47985,N_45660);
xnor UO_221 (O_221,N_49812,N_48332);
nand UO_222 (O_222,N_46002,N_48636);
and UO_223 (O_223,N_48401,N_49750);
or UO_224 (O_224,N_45344,N_48731);
and UO_225 (O_225,N_49307,N_47438);
xnor UO_226 (O_226,N_46437,N_47436);
or UO_227 (O_227,N_47225,N_46085);
and UO_228 (O_228,N_48303,N_46469);
nand UO_229 (O_229,N_45438,N_46683);
or UO_230 (O_230,N_45107,N_47763);
xor UO_231 (O_231,N_48820,N_45643);
xor UO_232 (O_232,N_49195,N_46144);
nor UO_233 (O_233,N_48504,N_46817);
xor UO_234 (O_234,N_49716,N_45474);
nand UO_235 (O_235,N_48448,N_48572);
nor UO_236 (O_236,N_46130,N_49459);
nand UO_237 (O_237,N_49847,N_49085);
xnor UO_238 (O_238,N_49303,N_45457);
and UO_239 (O_239,N_46632,N_48256);
or UO_240 (O_240,N_46861,N_49638);
xnor UO_241 (O_241,N_47830,N_47340);
nor UO_242 (O_242,N_45762,N_47477);
nand UO_243 (O_243,N_45158,N_47583);
xor UO_244 (O_244,N_48668,N_46708);
or UO_245 (O_245,N_47557,N_49688);
or UO_246 (O_246,N_48298,N_49761);
xor UO_247 (O_247,N_46167,N_47552);
xor UO_248 (O_248,N_48398,N_48053);
xnor UO_249 (O_249,N_45297,N_46027);
and UO_250 (O_250,N_45776,N_45129);
nor UO_251 (O_251,N_48378,N_45071);
nand UO_252 (O_252,N_47039,N_45837);
or UO_253 (O_253,N_49342,N_48576);
or UO_254 (O_254,N_48538,N_46518);
or UO_255 (O_255,N_48453,N_49283);
nor UO_256 (O_256,N_49705,N_45192);
xor UO_257 (O_257,N_49298,N_47270);
xor UO_258 (O_258,N_46636,N_49253);
nand UO_259 (O_259,N_46479,N_49288);
xnor UO_260 (O_260,N_48045,N_48996);
nor UO_261 (O_261,N_46100,N_49827);
or UO_262 (O_262,N_46297,N_47901);
nand UO_263 (O_263,N_47309,N_46448);
nand UO_264 (O_264,N_48671,N_47616);
xnor UO_265 (O_265,N_46270,N_49809);
nor UO_266 (O_266,N_48411,N_49744);
xor UO_267 (O_267,N_47629,N_47818);
nor UO_268 (O_268,N_48467,N_45902);
nor UO_269 (O_269,N_48443,N_49568);
and UO_270 (O_270,N_49989,N_47075);
nor UO_271 (O_271,N_46607,N_49820);
xnor UO_272 (O_272,N_49635,N_45503);
or UO_273 (O_273,N_47924,N_48730);
and UO_274 (O_274,N_46947,N_45146);
and UO_275 (O_275,N_48870,N_47651);
or UO_276 (O_276,N_47087,N_46277);
nand UO_277 (O_277,N_45752,N_46730);
xnor UO_278 (O_278,N_47705,N_49985);
or UO_279 (O_279,N_45798,N_47464);
or UO_280 (O_280,N_46080,N_49957);
or UO_281 (O_281,N_45834,N_47356);
nand UO_282 (O_282,N_45974,N_48049);
and UO_283 (O_283,N_45861,N_48188);
nor UO_284 (O_284,N_45406,N_45948);
nand UO_285 (O_285,N_48246,N_46756);
and UO_286 (O_286,N_45965,N_49111);
nor UO_287 (O_287,N_48072,N_48922);
and UO_288 (O_288,N_46529,N_48253);
nand UO_289 (O_289,N_45815,N_49504);
xnor UO_290 (O_290,N_45829,N_48068);
nand UO_291 (O_291,N_47623,N_48946);
and UO_292 (O_292,N_47832,N_45433);
nor UO_293 (O_293,N_46145,N_48108);
xor UO_294 (O_294,N_47479,N_47383);
nor UO_295 (O_295,N_48834,N_47447);
nand UO_296 (O_296,N_48341,N_45040);
xor UO_297 (O_297,N_47954,N_48030);
nor UO_298 (O_298,N_45575,N_49998);
or UO_299 (O_299,N_48548,N_46355);
or UO_300 (O_300,N_45847,N_46128);
nor UO_301 (O_301,N_46230,N_48077);
or UO_302 (O_302,N_48125,N_49746);
and UO_303 (O_303,N_49437,N_46302);
and UO_304 (O_304,N_49268,N_46054);
or UO_305 (O_305,N_47332,N_47516);
or UO_306 (O_306,N_47114,N_49592);
and UO_307 (O_307,N_45892,N_47455);
xnor UO_308 (O_308,N_48048,N_49718);
and UO_309 (O_309,N_47441,N_48131);
xnor UO_310 (O_310,N_46423,N_46836);
xnor UO_311 (O_311,N_47835,N_48565);
and UO_312 (O_312,N_46401,N_48858);
nand UO_313 (O_313,N_49202,N_46534);
nor UO_314 (O_314,N_46795,N_49186);
and UO_315 (O_315,N_49509,N_49021);
and UO_316 (O_316,N_48450,N_45719);
and UO_317 (O_317,N_47314,N_46716);
or UO_318 (O_318,N_47235,N_48015);
xor UO_319 (O_319,N_46304,N_49751);
nor UO_320 (O_320,N_48340,N_47158);
xor UO_321 (O_321,N_47619,N_46946);
nand UO_322 (O_322,N_49682,N_47543);
xnor UO_323 (O_323,N_46525,N_45147);
xor UO_324 (O_324,N_49691,N_49074);
xor UO_325 (O_325,N_48442,N_45536);
nor UO_326 (O_326,N_49830,N_45296);
and UO_327 (O_327,N_49323,N_46447);
and UO_328 (O_328,N_48469,N_49714);
nor UO_329 (O_329,N_46059,N_49850);
and UO_330 (O_330,N_49378,N_46504);
or UO_331 (O_331,N_45324,N_46788);
nor UO_332 (O_332,N_48087,N_47893);
nor UO_333 (O_333,N_49694,N_47115);
xnor UO_334 (O_334,N_45135,N_45317);
or UO_335 (O_335,N_48112,N_48252);
nand UO_336 (O_336,N_46413,N_47770);
nor UO_337 (O_337,N_45783,N_45538);
and UO_338 (O_338,N_45428,N_49524);
nor UO_339 (O_339,N_46689,N_47944);
or UO_340 (O_340,N_47412,N_46974);
nand UO_341 (O_341,N_48675,N_46291);
nand UO_342 (O_342,N_48796,N_49888);
xnor UO_343 (O_343,N_49089,N_47913);
or UO_344 (O_344,N_48404,N_45876);
xor UO_345 (O_345,N_45049,N_49123);
xor UO_346 (O_346,N_49144,N_47609);
or UO_347 (O_347,N_48235,N_49962);
xnor UO_348 (O_348,N_47978,N_49087);
or UO_349 (O_349,N_45465,N_48331);
and UO_350 (O_350,N_45415,N_45649);
or UO_351 (O_351,N_48707,N_45398);
nor UO_352 (O_352,N_47338,N_46827);
or UO_353 (O_353,N_49650,N_47009);
and UO_354 (O_354,N_47408,N_48530);
nand UO_355 (O_355,N_49080,N_47361);
nand UO_356 (O_356,N_46368,N_46599);
and UO_357 (O_357,N_48510,N_46495);
and UO_358 (O_358,N_48200,N_47130);
nand UO_359 (O_359,N_45699,N_48903);
and UO_360 (O_360,N_49797,N_45364);
xor UO_361 (O_361,N_46266,N_47904);
nor UO_362 (O_362,N_46464,N_47630);
xnor UO_363 (O_363,N_47252,N_49376);
or UO_364 (O_364,N_46679,N_49062);
nor UO_365 (O_365,N_48395,N_46962);
nand UO_366 (O_366,N_49222,N_45571);
nand UO_367 (O_367,N_45619,N_49492);
nor UO_368 (O_368,N_48308,N_46186);
or UO_369 (O_369,N_49269,N_49008);
nand UO_370 (O_370,N_45496,N_47352);
or UO_371 (O_371,N_48521,N_45484);
xor UO_372 (O_372,N_45832,N_45137);
and UO_373 (O_373,N_46143,N_48230);
or UO_374 (O_374,N_46593,N_49855);
and UO_375 (O_375,N_45726,N_46581);
and UO_376 (O_376,N_45006,N_48290);
nor UO_377 (O_377,N_49968,N_46347);
or UO_378 (O_378,N_45276,N_48983);
xnor UO_379 (O_379,N_46336,N_46909);
and UO_380 (O_380,N_48727,N_46582);
nor UO_381 (O_381,N_46308,N_47882);
or UO_382 (O_382,N_46246,N_45185);
and UO_383 (O_383,N_49050,N_45483);
and UO_384 (O_384,N_47790,N_45096);
and UO_385 (O_385,N_45267,N_45092);
or UO_386 (O_386,N_49005,N_45004);
xnor UO_387 (O_387,N_47905,N_46570);
or UO_388 (O_388,N_49563,N_49514);
nor UO_389 (O_389,N_48351,N_46299);
nand UO_390 (O_390,N_47753,N_45222);
and UO_391 (O_391,N_49777,N_45684);
xnor UO_392 (O_392,N_49815,N_48054);
nand UO_393 (O_393,N_46047,N_46844);
xor UO_394 (O_394,N_49498,N_47859);
nor UO_395 (O_395,N_46833,N_47544);
and UO_396 (O_396,N_48580,N_48992);
nand UO_397 (O_397,N_46229,N_48687);
and UO_398 (O_398,N_49236,N_48611);
nor UO_399 (O_399,N_46485,N_45275);
nor UO_400 (O_400,N_45255,N_49707);
nor UO_401 (O_401,N_47398,N_48910);
or UO_402 (O_402,N_47132,N_48234);
and UO_403 (O_403,N_47232,N_45358);
xor UO_404 (O_404,N_45860,N_45001);
nand UO_405 (O_405,N_47149,N_48683);
nand UO_406 (O_406,N_45515,N_45785);
xor UO_407 (O_407,N_46832,N_47312);
or UO_408 (O_408,N_46860,N_48837);
nor UO_409 (O_409,N_48078,N_49934);
and UO_410 (O_410,N_47059,N_46288);
xor UO_411 (O_411,N_49064,N_47618);
or UO_412 (O_412,N_48713,N_47217);
or UO_413 (O_413,N_47632,N_47890);
and UO_414 (O_414,N_45201,N_48699);
and UO_415 (O_415,N_46383,N_45126);
nand UO_416 (O_416,N_47707,N_47316);
and UO_417 (O_417,N_48312,N_47145);
xnor UO_418 (O_418,N_49511,N_45733);
or UO_419 (O_419,N_45630,N_48899);
xnor UO_420 (O_420,N_47005,N_47604);
and UO_421 (O_421,N_46643,N_49265);
xnor UO_422 (O_422,N_48923,N_48930);
xnor UO_423 (O_423,N_45805,N_47966);
or UO_424 (O_424,N_46532,N_46315);
xnor UO_425 (O_425,N_46791,N_46300);
nand UO_426 (O_426,N_45673,N_45426);
xor UO_427 (O_427,N_49149,N_48579);
and UO_428 (O_428,N_45794,N_45077);
nor UO_429 (O_429,N_49629,N_47099);
xnor UO_430 (O_430,N_45003,N_45909);
nand UO_431 (O_431,N_49267,N_47262);
or UO_432 (O_432,N_48266,N_45361);
nand UO_433 (O_433,N_48302,N_47128);
or UO_434 (O_434,N_48705,N_48104);
xor UO_435 (O_435,N_48174,N_46664);
and UO_436 (O_436,N_47950,N_46848);
xor UO_437 (O_437,N_48915,N_47750);
nor UO_438 (O_438,N_45542,N_49826);
nand UO_439 (O_439,N_46478,N_49938);
or UO_440 (O_440,N_49091,N_45934);
nand UO_441 (O_441,N_47065,N_48427);
nand UO_442 (O_442,N_49570,N_49068);
nand UO_443 (O_443,N_47601,N_48409);
or UO_444 (O_444,N_45970,N_49250);
nor UO_445 (O_445,N_46170,N_46125);
xor UO_446 (O_446,N_49067,N_45044);
nor UO_447 (O_447,N_48978,N_49347);
nand UO_448 (O_448,N_48163,N_49569);
nor UO_449 (O_449,N_49086,N_49280);
nor UO_450 (O_450,N_45856,N_48180);
xor UO_451 (O_451,N_48561,N_49781);
nor UO_452 (O_452,N_48637,N_46815);
nor UO_453 (O_453,N_49737,N_45658);
xnor UO_454 (O_454,N_47472,N_47336);
and UO_455 (O_455,N_46373,N_49622);
xor UO_456 (O_456,N_47296,N_48571);
xnor UO_457 (O_457,N_48733,N_46010);
nor UO_458 (O_458,N_46487,N_46159);
and UO_459 (O_459,N_46904,N_47082);
nor UO_460 (O_460,N_49789,N_46012);
nor UO_461 (O_461,N_48976,N_48301);
and UO_462 (O_462,N_49432,N_46605);
xnor UO_463 (O_463,N_49426,N_48639);
nor UO_464 (O_464,N_48310,N_46552);
nand UO_465 (O_465,N_47712,N_46150);
or UO_466 (O_466,N_47370,N_49546);
nor UO_467 (O_467,N_46314,N_48187);
nor UO_468 (O_468,N_45763,N_45429);
and UO_469 (O_469,N_45661,N_45208);
xnor UO_470 (O_470,N_48314,N_46577);
nor UO_471 (O_471,N_49251,N_48982);
nand UO_472 (O_472,N_47416,N_47254);
xnor UO_473 (O_473,N_47852,N_49413);
xor UO_474 (O_474,N_49681,N_48232);
nand UO_475 (O_475,N_45879,N_47036);
nand UO_476 (O_476,N_47969,N_49978);
and UO_477 (O_477,N_47939,N_47856);
nor UO_478 (O_478,N_47213,N_47376);
nand UO_479 (O_479,N_48224,N_47205);
nor UO_480 (O_480,N_49651,N_47845);
nor UO_481 (O_481,N_46147,N_49762);
nor UO_482 (O_482,N_48833,N_45809);
or UO_483 (O_483,N_47349,N_46062);
and UO_484 (O_484,N_49659,N_47157);
or UO_485 (O_485,N_45610,N_46615);
nor UO_486 (O_486,N_45857,N_45439);
or UO_487 (O_487,N_49548,N_48319);
or UO_488 (O_488,N_45866,N_47582);
nand UO_489 (O_489,N_48160,N_48279);
and UO_490 (O_490,N_45101,N_47889);
nand UO_491 (O_491,N_48009,N_46097);
xnor UO_492 (O_492,N_48993,N_49906);
nand UO_493 (O_493,N_48508,N_49515);
or UO_494 (O_494,N_46141,N_46792);
or UO_495 (O_495,N_49642,N_47175);
nand UO_496 (O_496,N_46949,N_47864);
or UO_497 (O_497,N_45248,N_46879);
or UO_498 (O_498,N_45983,N_48662);
and UO_499 (O_499,N_45099,N_45862);
nor UO_500 (O_500,N_48219,N_45817);
nand UO_501 (O_501,N_45336,N_45806);
nand UO_502 (O_502,N_45460,N_48278);
and UO_503 (O_503,N_45298,N_48255);
xnor UO_504 (O_504,N_47341,N_45534);
and UO_505 (O_505,N_49792,N_48231);
nor UO_506 (O_506,N_46285,N_47857);
nor UO_507 (O_507,N_46545,N_45797);
or UO_508 (O_508,N_46618,N_45367);
nand UO_509 (O_509,N_48058,N_48654);
nand UO_510 (O_510,N_48540,N_49355);
or UO_511 (O_511,N_49620,N_46785);
and UO_512 (O_512,N_49281,N_49669);
xnor UO_513 (O_513,N_48457,N_46682);
nand UO_514 (O_514,N_49199,N_49057);
nand UO_515 (O_515,N_46950,N_46105);
nand UO_516 (O_516,N_48120,N_46456);
nand UO_517 (O_517,N_48901,N_47473);
nor UO_518 (O_518,N_45034,N_45997);
and UO_519 (O_519,N_47929,N_49055);
xor UO_520 (O_520,N_48095,N_47594);
nor UO_521 (O_521,N_47709,N_46108);
or UO_522 (O_522,N_48994,N_47781);
nand UO_523 (O_523,N_48083,N_46074);
xnor UO_524 (O_524,N_49698,N_49393);
or UO_525 (O_525,N_48449,N_45968);
or UO_526 (O_526,N_49794,N_49770);
or UO_527 (O_527,N_45310,N_47297);
and UO_528 (O_528,N_49956,N_45284);
nor UO_529 (O_529,N_47765,N_46160);
xor UO_530 (O_530,N_49337,N_49520);
and UO_531 (O_531,N_45124,N_47403);
and UO_532 (O_532,N_45123,N_47574);
nor UO_533 (O_533,N_48882,N_45102);
nor UO_534 (O_534,N_48509,N_45921);
and UO_535 (O_535,N_47320,N_48626);
nand UO_536 (O_536,N_49921,N_46551);
xor UO_537 (O_537,N_45705,N_46262);
or UO_538 (O_538,N_45108,N_46758);
or UO_539 (O_539,N_46119,N_45512);
or UO_540 (O_540,N_46796,N_46737);
or UO_541 (O_541,N_49851,N_48052);
nor UO_542 (O_542,N_48533,N_47573);
or UO_543 (O_543,N_46365,N_45950);
and UO_544 (O_544,N_45795,N_45068);
and UO_545 (O_545,N_46451,N_48781);
nor UO_546 (O_546,N_47808,N_45606);
and UO_547 (O_547,N_46041,N_45530);
xor UO_548 (O_548,N_49029,N_47989);
nor UO_549 (O_549,N_46690,N_49613);
or UO_550 (O_550,N_48810,N_46671);
xor UO_551 (O_551,N_47048,N_45166);
nor UO_552 (O_552,N_49963,N_47131);
or UO_553 (O_553,N_47084,N_46514);
and UO_554 (O_554,N_45939,N_45569);
or UO_555 (O_555,N_48515,N_49301);
xnor UO_556 (O_556,N_48949,N_46657);
and UO_557 (O_557,N_45319,N_47888);
nand UO_558 (O_558,N_48386,N_46574);
nor UO_559 (O_559,N_48205,N_49270);
nor UO_560 (O_560,N_48069,N_48900);
nand UO_561 (O_561,N_46214,N_49473);
or UO_562 (O_562,N_47446,N_49249);
or UO_563 (O_563,N_48451,N_48818);
xnor UO_564 (O_564,N_47096,N_47325);
or UO_565 (O_565,N_47188,N_46903);
nand UO_566 (O_566,N_49313,N_47454);
nand UO_567 (O_567,N_49041,N_46849);
nor UO_568 (O_568,N_47633,N_48537);
nand UO_569 (O_569,N_47773,N_49666);
or UO_570 (O_570,N_47467,N_45893);
xnor UO_571 (O_571,N_47110,N_47164);
or UO_572 (O_572,N_47529,N_45143);
nand UO_573 (O_573,N_48865,N_46706);
nand UO_574 (O_574,N_49558,N_45490);
or UO_575 (O_575,N_48886,N_49724);
or UO_576 (O_576,N_45434,N_46568);
and UO_577 (O_577,N_47431,N_46418);
or UO_578 (O_578,N_46979,N_47346);
or UO_579 (O_579,N_47218,N_48583);
and UO_580 (O_580,N_48926,N_45867);
and UO_581 (O_581,N_49094,N_49880);
or UO_582 (O_582,N_49185,N_47641);
nand UO_583 (O_583,N_45468,N_49673);
or UO_584 (O_584,N_49832,N_48271);
or UO_585 (O_585,N_49447,N_47081);
nor UO_586 (O_586,N_47117,N_48455);
or UO_587 (O_587,N_48610,N_48744);
nand UO_588 (O_588,N_49722,N_49930);
xnor UO_589 (O_589,N_45510,N_48981);
or UO_590 (O_590,N_46869,N_46713);
and UO_591 (O_591,N_47470,N_47760);
xor UO_592 (O_592,N_48955,N_47116);
nor UO_593 (O_593,N_48648,N_46665);
or UO_594 (O_594,N_45846,N_46908);
xnor UO_595 (O_595,N_49760,N_46595);
nor UO_596 (O_596,N_45682,N_45355);
or UO_597 (O_597,N_46675,N_48149);
xnor UO_598 (O_598,N_49867,N_49799);
nand UO_599 (O_599,N_49286,N_47567);
xnor UO_600 (O_600,N_45432,N_45521);
or UO_601 (O_601,N_46654,N_49776);
or UO_602 (O_602,N_45171,N_46064);
xnor UO_603 (O_603,N_48329,N_46994);
nand UO_604 (O_604,N_47359,N_47491);
nand UO_605 (O_605,N_47877,N_48578);
nand UO_606 (O_606,N_47537,N_48739);
or UO_607 (O_607,N_48897,N_49507);
or UO_608 (O_608,N_46472,N_46492);
nor UO_609 (O_609,N_46405,N_47226);
and UO_610 (O_610,N_45118,N_49767);
xnor UO_611 (O_611,N_48309,N_45401);
nand UO_612 (O_612,N_49118,N_46740);
and UO_613 (O_613,N_48827,N_48094);
and UO_614 (O_614,N_47821,N_46764);
and UO_615 (O_615,N_45932,N_48086);
and UO_616 (O_616,N_46473,N_46428);
xor UO_617 (O_617,N_46118,N_48186);
nand UO_618 (O_618,N_46575,N_46452);
xnor UO_619 (O_619,N_46850,N_45427);
and UO_620 (O_620,N_49227,N_45295);
and UO_621 (O_621,N_48140,N_45253);
nand UO_622 (O_622,N_48494,N_47306);
nor UO_623 (O_623,N_49984,N_49800);
nand UO_624 (O_624,N_48766,N_47339);
and UO_625 (O_625,N_48222,N_46163);
and UO_626 (O_626,N_48216,N_47741);
and UO_627 (O_627,N_47796,N_47909);
xor UO_628 (O_628,N_47827,N_45421);
xor UO_629 (O_629,N_48653,N_48944);
nor UO_630 (O_630,N_46281,N_47621);
nand UO_631 (O_631,N_47187,N_47379);
nand UO_632 (O_632,N_46362,N_47050);
and UO_633 (O_633,N_45424,N_46987);
and UO_634 (O_634,N_46232,N_47690);
and UO_635 (O_635,N_48318,N_49302);
xnor UO_636 (O_636,N_49804,N_47069);
nand UO_637 (O_637,N_45187,N_48354);
xor UO_638 (O_638,N_46474,N_46173);
or UO_639 (O_639,N_46798,N_46226);
xor UO_640 (O_640,N_46517,N_47103);
xnor UO_641 (O_641,N_49436,N_48189);
or UO_642 (O_642,N_48500,N_47754);
nand UO_643 (O_643,N_46274,N_49656);
or UO_644 (O_644,N_48371,N_45089);
and UO_645 (O_645,N_49176,N_49660);
nor UO_646 (O_646,N_46660,N_46396);
nand UO_647 (O_647,N_46042,N_49483);
nand UO_648 (O_648,N_45587,N_46136);
nor UO_649 (O_649,N_46426,N_45414);
nor UO_650 (O_650,N_45008,N_46283);
and UO_651 (O_651,N_45548,N_46455);
and UO_652 (O_652,N_46559,N_48997);
nor UO_653 (O_653,N_49545,N_47063);
or UO_654 (O_654,N_47163,N_49566);
nand UO_655 (O_655,N_45712,N_47993);
or UO_656 (O_656,N_46476,N_46963);
nor UO_657 (O_657,N_48931,N_46013);
nor UO_658 (O_658,N_48970,N_48817);
or UO_659 (O_659,N_45469,N_48587);
nand UO_660 (O_660,N_46537,N_47483);
xor UO_661 (O_661,N_48914,N_45487);
nor UO_662 (O_662,N_49237,N_48498);
or UO_663 (O_663,N_49912,N_48070);
xor UO_664 (O_664,N_48987,N_46929);
nor UO_665 (O_665,N_48300,N_45900);
xor UO_666 (O_666,N_49322,N_45625);
or UO_667 (O_667,N_45692,N_47421);
xnor UO_668 (O_668,N_49664,N_49852);
nor UO_669 (O_669,N_49456,N_46656);
nand UO_670 (O_670,N_45686,N_47198);
nand UO_671 (O_671,N_46056,N_46960);
nand UO_672 (O_672,N_47662,N_46584);
or UO_673 (O_673,N_45588,N_47871);
or UO_674 (O_674,N_47720,N_49403);
xnor UO_675 (O_675,N_45261,N_45714);
nor UO_676 (O_676,N_48889,N_45517);
nor UO_677 (O_677,N_49255,N_47659);
and UO_678 (O_678,N_49485,N_46993);
and UO_679 (O_679,N_46854,N_48697);
xnor UO_680 (O_680,N_47926,N_47032);
and UO_681 (O_681,N_45029,N_49279);
and UO_682 (O_682,N_45940,N_49312);
xor UO_683 (O_683,N_46001,N_46727);
and UO_684 (O_684,N_49412,N_45448);
nand UO_685 (O_685,N_49708,N_47916);
or UO_686 (O_686,N_48961,N_49607);
and UO_687 (O_687,N_47461,N_48452);
or UO_688 (O_688,N_45999,N_48280);
nor UO_689 (O_689,N_48547,N_45563);
and UO_690 (O_690,N_45329,N_45012);
and UO_691 (O_691,N_48020,N_46482);
and UO_692 (O_692,N_48634,N_49765);
nand UO_693 (O_693,N_46335,N_47850);
or UO_694 (O_694,N_48562,N_47540);
nor UO_695 (O_695,N_48563,N_46185);
xor UO_696 (O_696,N_49655,N_48181);
and UO_697 (O_697,N_46206,N_49206);
nor UO_698 (O_698,N_48645,N_47020);
and UO_699 (O_699,N_47549,N_45737);
and UO_700 (O_700,N_45803,N_47927);
and UO_701 (O_701,N_49877,N_47884);
nand UO_702 (O_702,N_48063,N_48768);
nor UO_703 (O_703,N_46953,N_48542);
nand UO_704 (O_704,N_45786,N_45949);
nor UO_705 (O_705,N_45654,N_45031);
nand UO_706 (O_706,N_49452,N_49061);
xnor UO_707 (O_707,N_46549,N_49165);
and UO_708 (O_708,N_46076,N_47930);
nor UO_709 (O_709,N_49536,N_49294);
xor UO_710 (O_710,N_48883,N_47591);
nor UO_711 (O_711,N_47697,N_47109);
and UO_712 (O_712,N_46771,N_45311);
nand UO_713 (O_713,N_47234,N_45853);
xnor UO_714 (O_714,N_45604,N_46014);
and UO_715 (O_715,N_45603,N_48345);
or UO_716 (O_716,N_48067,N_45662);
nor UO_717 (O_717,N_48433,N_45870);
nor UO_718 (O_718,N_46948,N_48753);
xor UO_719 (O_719,N_46981,N_45133);
nor UO_720 (O_720,N_46364,N_48285);
and UO_721 (O_721,N_48114,N_48826);
xnor UO_722 (O_722,N_48383,N_46721);
nand UO_723 (O_723,N_45992,N_46816);
nor UO_724 (O_724,N_48908,N_46808);
and UO_725 (O_725,N_45629,N_48193);
and UO_726 (O_726,N_49103,N_46621);
or UO_727 (O_727,N_45327,N_48038);
or UO_728 (O_728,N_49495,N_46111);
xnor UO_729 (O_729,N_46757,N_45345);
and UO_730 (O_730,N_49226,N_45037);
xnor UO_731 (O_731,N_48825,N_47874);
nor UO_732 (O_732,N_45828,N_48440);
xnor UO_733 (O_733,N_49769,N_45480);
nor UO_734 (O_734,N_46462,N_46328);
nand UO_735 (O_735,N_49168,N_47735);
or UO_736 (O_736,N_47143,N_47224);
nand UO_737 (O_737,N_48079,N_47167);
or UO_738 (O_738,N_45611,N_49745);
xnor UO_739 (O_739,N_48468,N_46332);
nor UO_740 (O_740,N_46500,N_48811);
xor UO_741 (O_741,N_45657,N_45823);
or UO_742 (O_742,N_49344,N_45254);
or UO_743 (O_743,N_47976,N_46259);
nor UO_744 (O_744,N_47313,N_45269);
and UO_745 (O_745,N_45523,N_47192);
or UO_746 (O_746,N_46467,N_49053);
nor UO_747 (O_747,N_48373,N_45417);
nor UO_748 (O_748,N_49825,N_47334);
or UO_749 (O_749,N_48523,N_48485);
nand UO_750 (O_750,N_48711,N_49210);
and UO_751 (O_751,N_49639,N_46697);
nor UO_752 (O_752,N_48765,N_46542);
and UO_753 (O_753,N_46784,N_48097);
xor UO_754 (O_754,N_45309,N_46446);
and UO_755 (O_755,N_49713,N_45841);
nor UO_756 (O_756,N_45346,N_47369);
nor UO_757 (O_757,N_47273,N_47259);
nor UO_758 (O_758,N_47797,N_47778);
or UO_759 (O_759,N_49680,N_48370);
nand UO_760 (O_760,N_46983,N_48328);
nor UO_761 (O_761,N_47236,N_49873);
and UO_762 (O_762,N_46563,N_47010);
nand UO_763 (O_763,N_49129,N_46975);
and UO_764 (O_764,N_48938,N_49649);
nand UO_765 (O_765,N_45788,N_48943);
xnor UO_766 (O_766,N_48559,N_46131);
or UO_767 (O_767,N_48132,N_47843);
nand UO_768 (O_768,N_46494,N_45493);
nand UO_769 (O_769,N_47736,N_47631);
xor UO_770 (O_770,N_47739,N_46165);
xnor UO_771 (O_771,N_45482,N_47200);
nand UO_772 (O_772,N_48935,N_47894);
xor UO_773 (O_773,N_48158,N_47732);
nand UO_774 (O_774,N_45168,N_48389);
xnor UO_775 (O_775,N_45875,N_45648);
nand UO_776 (O_776,N_46940,N_45953);
and UO_777 (O_777,N_46433,N_45858);
or UO_778 (O_778,N_45908,N_45519);
or UO_779 (O_779,N_46235,N_47660);
and UO_780 (O_780,N_45030,N_49444);
or UO_781 (O_781,N_49875,N_46161);
xnor UO_782 (O_782,N_48867,N_49586);
nand UO_783 (O_783,N_46294,N_46895);
and UO_784 (O_784,N_46880,N_47716);
and UO_785 (O_785,N_49581,N_47404);
nand UO_786 (O_786,N_46239,N_48348);
nor UO_787 (O_787,N_48465,N_46127);
nand UO_788 (O_788,N_47196,N_45646);
xor UO_789 (O_789,N_45645,N_45540);
nand UO_790 (O_790,N_45182,N_45498);
or UO_791 (O_791,N_46095,N_47360);
and UO_792 (O_792,N_47183,N_47899);
nand UO_793 (O_793,N_46318,N_46484);
nand UO_794 (O_794,N_46866,N_47364);
nand UO_795 (O_795,N_48135,N_49731);
nand UO_796 (O_796,N_49058,N_45735);
and UO_797 (O_797,N_48358,N_48414);
nor UO_798 (O_798,N_49550,N_48717);
xnor UO_799 (O_799,N_46334,N_45307);
and UO_800 (O_800,N_48526,N_47411);
xnor UO_801 (O_801,N_49119,N_47568);
nor UO_802 (O_802,N_46172,N_45151);
and UO_803 (O_803,N_46079,N_46630);
xor UO_804 (O_804,N_45980,N_49246);
or UO_805 (O_805,N_49846,N_47144);
or UO_806 (O_806,N_49677,N_47553);
and UO_807 (O_807,N_46496,N_46260);
and UO_808 (O_808,N_47925,N_46965);
and UO_809 (O_809,N_48282,N_49623);
and UO_810 (O_810,N_45039,N_46692);
or UO_811 (O_811,N_47056,N_48407);
and UO_812 (O_812,N_48689,N_47578);
nor UO_813 (O_813,N_46444,N_46628);
and UO_814 (O_814,N_46761,N_45579);
nand UO_815 (O_815,N_45525,N_47903);
xor UO_816 (O_816,N_49663,N_45680);
xnor UO_817 (O_817,N_46427,N_48551);
or UO_818 (O_818,N_45747,N_47900);
nand UO_819 (O_819,N_48748,N_49951);
nor UO_820 (O_820,N_47704,N_45996);
and UO_821 (O_821,N_47592,N_47724);
or UO_822 (O_822,N_46888,N_46865);
nand UO_823 (O_823,N_45766,N_48134);
xnor UO_824 (O_824,N_45759,N_45459);
or UO_825 (O_825,N_45373,N_48263);
nand UO_826 (O_826,N_48871,N_46591);
and UO_827 (O_827,N_46070,N_48029);
and UO_828 (O_828,N_49252,N_48724);
and UO_829 (O_829,N_47854,N_46280);
or UO_830 (O_830,N_46068,N_47776);
or UO_831 (O_831,N_49598,N_47393);
and UO_832 (O_832,N_47727,N_45047);
nor UO_833 (O_833,N_48264,N_45500);
nand UO_834 (O_834,N_48210,N_46731);
xor UO_835 (O_835,N_48691,N_48862);
or UO_836 (O_836,N_47960,N_46527);
and UO_837 (O_837,N_46234,N_46356);
and UO_838 (O_838,N_49049,N_47151);
or UO_839 (O_839,N_45928,N_47918);
or UO_840 (O_840,N_45206,N_47804);
and UO_841 (O_841,N_48921,N_49142);
nor UO_842 (O_842,N_47600,N_48172);
xor UO_843 (O_843,N_48487,N_49339);
nand UO_844 (O_844,N_47170,N_45811);
xor UO_845 (O_845,N_47751,N_47661);
and UO_846 (O_846,N_45816,N_46480);
xnor UO_847 (O_847,N_45989,N_45057);
or UO_848 (O_848,N_49203,N_46544);
xor UO_849 (O_849,N_46768,N_48435);
nand UO_850 (O_850,N_48202,N_47420);
or UO_851 (O_851,N_48192,N_47866);
nand UO_852 (O_852,N_48213,N_48642);
or UO_853 (O_853,N_49665,N_49348);
nand UO_854 (O_854,N_47282,N_49727);
xor UO_855 (O_855,N_45226,N_49299);
or UO_856 (O_856,N_49416,N_47558);
or UO_857 (O_857,N_46290,N_49844);
and UO_858 (O_858,N_47239,N_47626);
or UO_859 (O_859,N_49484,N_49872);
nor UO_860 (O_860,N_49155,N_45971);
or UO_861 (O_861,N_47488,N_49449);
xnor UO_862 (O_862,N_49940,N_45435);
nor UO_863 (O_863,N_49571,N_49685);
xor UO_864 (O_864,N_48165,N_49990);
and UO_865 (O_865,N_46020,N_45628);
and UO_866 (O_866,N_48399,N_47299);
and UO_867 (O_867,N_48879,N_45917);
and UO_868 (O_868,N_48306,N_45396);
and UO_869 (O_869,N_46434,N_49600);
xnor UO_870 (O_870,N_48139,N_48299);
nand UO_871 (O_871,N_45933,N_49964);
nand UO_872 (O_872,N_48906,N_48338);
and UO_873 (O_873,N_45189,N_47524);
nand UO_874 (O_874,N_49461,N_45190);
and UO_875 (O_875,N_47414,N_49740);
and UO_876 (O_876,N_46714,N_45995);
xor UO_877 (O_877,N_49167,N_49319);
nand UO_878 (O_878,N_45728,N_45778);
nor UO_879 (O_879,N_45873,N_47322);
nand UO_880 (O_880,N_47450,N_48732);
xor UO_881 (O_881,N_46573,N_47173);
nor UO_882 (O_882,N_46242,N_47645);
nand UO_883 (O_883,N_49207,N_46440);
xor UO_884 (O_884,N_45066,N_48403);
and UO_885 (O_885,N_45403,N_47290);
nor UO_886 (O_886,N_45094,N_45352);
or UO_887 (O_887,N_47471,N_47547);
nor UO_888 (O_888,N_48641,N_48549);
and UO_889 (O_889,N_48718,N_47640);
nor UO_890 (O_890,N_48317,N_47153);
nand UO_891 (O_891,N_48966,N_46344);
and UO_892 (O_892,N_47280,N_45966);
nor UO_893 (O_893,N_46579,N_45156);
nor UO_894 (O_894,N_48606,N_47896);
nand UO_895 (O_895,N_47711,N_49217);
nor UO_896 (O_896,N_48894,N_49679);
nand UO_897 (O_897,N_46729,N_49469);
nor UO_898 (O_898,N_45958,N_49965);
nand UO_899 (O_899,N_48898,N_48885);
nor UO_900 (O_900,N_49723,N_47608);
nand UO_901 (O_901,N_46847,N_47119);
nor UO_902 (O_902,N_49516,N_45272);
xnor UO_903 (O_903,N_48482,N_48893);
and UO_904 (O_904,N_48335,N_45602);
nor UO_905 (O_905,N_47172,N_49063);
xor UO_906 (O_906,N_49555,N_48741);
and UO_907 (O_907,N_47545,N_49857);
nand UO_908 (O_908,N_48473,N_46701);
or UO_909 (O_909,N_45333,N_45868);
nor UO_910 (O_910,N_45279,N_45961);
xnor UO_911 (O_911,N_46258,N_49513);
nor UO_912 (O_912,N_46354,N_47342);
nor UO_913 (O_913,N_48761,N_45240);
nor UO_914 (O_914,N_49243,N_46924);
nor UO_915 (O_915,N_45777,N_47008);
and UO_916 (O_916,N_48507,N_49228);
nand UO_917 (O_917,N_45659,N_47043);
nand UO_918 (O_918,N_46845,N_46746);
nand UO_919 (O_919,N_45286,N_49899);
and UO_920 (O_920,N_48659,N_47987);
nand UO_921 (O_921,N_46109,N_48754);
xnor UO_922 (O_922,N_46420,N_46498);
nand UO_923 (O_923,N_46182,N_47559);
nand UO_924 (O_924,N_46322,N_49160);
nor UO_925 (O_925,N_49009,N_45964);
or UO_926 (O_926,N_47879,N_47920);
xnor UO_927 (O_927,N_46382,N_46011);
or UO_928 (O_928,N_47399,N_48410);
nand UO_929 (O_929,N_49122,N_49277);
nor UO_930 (O_930,N_49445,N_47142);
nand UO_931 (O_931,N_45271,N_49466);
nand UO_932 (O_932,N_47089,N_49726);
nand UO_933 (O_933,N_46254,N_46191);
nor UO_934 (O_934,N_49178,N_47137);
nand UO_935 (O_935,N_48111,N_48632);
nor UO_936 (O_936,N_47015,N_47936);
or UO_937 (O_937,N_47955,N_45993);
xnor UO_938 (O_938,N_49824,N_45334);
xnor UO_939 (O_939,N_46151,N_45050);
xnor UO_940 (O_940,N_49927,N_46178);
nand UO_941 (O_941,N_45476,N_46918);
nor UO_942 (O_942,N_49897,N_48339);
xor UO_943 (O_943,N_45609,N_46093);
or UO_944 (O_944,N_46286,N_46379);
nand UO_945 (O_945,N_45061,N_45626);
nor UO_946 (O_946,N_46877,N_45239);
or UO_947 (O_947,N_46249,N_45772);
xnor UO_948 (O_948,N_47620,N_45138);
or UO_949 (O_949,N_47657,N_49743);
xor UO_950 (O_950,N_46466,N_48846);
xnor UO_951 (O_951,N_45405,N_46642);
and UO_952 (O_952,N_49774,N_48850);
nor UO_953 (O_953,N_46459,N_46021);
nand UO_954 (O_954,N_47875,N_46668);
or UO_955 (O_955,N_46233,N_45963);
xor UO_956 (O_956,N_47809,N_45706);
nor UO_957 (O_957,N_45635,N_47782);
or UO_958 (O_958,N_47813,N_46148);
nor UO_959 (O_959,N_48183,N_48896);
and UO_960 (O_960,N_46878,N_49803);
and UO_961 (O_961,N_45180,N_47738);
xor UO_962 (O_962,N_47426,N_46611);
nor UO_963 (O_963,N_47556,N_46958);
xnor UO_964 (O_964,N_49356,N_45698);
nor UO_965 (O_965,N_46576,N_48682);
nand UO_966 (O_966,N_46330,N_47490);
nand UO_967 (O_967,N_47041,N_46051);
or UO_968 (O_968,N_49734,N_46099);
or UO_969 (O_969,N_47643,N_45577);
nor UO_970 (O_970,N_48505,N_49983);
and UO_971 (O_971,N_45316,N_46863);
nor UO_972 (O_972,N_46773,N_49876);
nand UO_973 (O_973,N_45227,N_45173);
xnor UO_974 (O_974,N_49821,N_49081);
or UO_975 (O_975,N_49611,N_46454);
xor UO_976 (O_976,N_47748,N_47025);
and UO_977 (O_977,N_47256,N_46104);
and UO_978 (O_978,N_48740,N_49429);
nor UO_979 (O_979,N_47590,N_45172);
nor UO_980 (O_980,N_49950,N_48463);
nand UO_981 (O_981,N_45773,N_45463);
nor UO_982 (O_982,N_49942,N_48736);
or UO_983 (O_983,N_46776,N_46156);
nor UO_984 (O_984,N_45882,N_49354);
nand UO_985 (O_985,N_47742,N_45915);
xnor UO_986 (O_986,N_48025,N_46580);
nand UO_987 (O_987,N_49408,N_48342);
xnor UO_988 (O_988,N_46194,N_48801);
or UO_989 (O_989,N_49937,N_47500);
nand UO_990 (O_990,N_47512,N_48940);
nor UO_991 (O_991,N_47931,N_45289);
and UO_992 (O_992,N_48831,N_45621);
or UO_993 (O_993,N_45093,N_47676);
nor UO_994 (O_994,N_49919,N_49019);
and UO_995 (O_995,N_46633,N_46370);
and UO_996 (O_996,N_47825,N_47374);
nand UO_997 (O_997,N_49567,N_46766);
nor UO_998 (O_998,N_47554,N_49434);
xor UO_999 (O_999,N_46133,N_49054);
or UO_1000 (O_1000,N_48799,N_49858);
or UO_1001 (O_1001,N_47539,N_47329);
and UO_1002 (O_1002,N_47502,N_48567);
nor UO_1003 (O_1003,N_48553,N_49419);
nand UO_1004 (O_1004,N_49154,N_46902);
xor UO_1005 (O_1005,N_48635,N_45251);
or UO_1006 (O_1006,N_45838,N_47417);
xnor UO_1007 (O_1007,N_48947,N_45256);
nor UO_1008 (O_1008,N_48081,N_45038);
nand UO_1009 (O_1009,N_46753,N_48700);
nand UO_1010 (O_1010,N_45990,N_47092);
nor UO_1011 (O_1011,N_48330,N_45265);
and UO_1012 (O_1012,N_46984,N_46083);
nand UO_1013 (O_1013,N_45451,N_49528);
nor UO_1014 (O_1014,N_48382,N_46889);
or UO_1015 (O_1015,N_49095,N_47186);
and UO_1016 (O_1016,N_49869,N_47510);
or UO_1017 (O_1017,N_45765,N_45945);
nor UO_1018 (O_1018,N_48161,N_49013);
and UO_1019 (O_1019,N_45905,N_48933);
nor UO_1020 (O_1020,N_47046,N_45339);
or UO_1021 (O_1021,N_48145,N_48715);
or UO_1022 (O_1022,N_45709,N_47566);
xnor UO_1023 (O_1023,N_45849,N_49868);
or UO_1024 (O_1024,N_48026,N_45268);
and UO_1025 (O_1025,N_45067,N_46431);
nand UO_1026 (O_1026,N_49542,N_46876);
xnor UO_1027 (O_1027,N_47841,N_45262);
or UO_1028 (O_1028,N_45052,N_48249);
xor UO_1029 (O_1029,N_45871,N_49433);
xor UO_1030 (O_1030,N_47400,N_49296);
nor UO_1031 (O_1031,N_46912,N_46110);
or UO_1032 (O_1032,N_47886,N_47422);
nor UO_1033 (O_1033,N_48963,N_49532);
and UO_1034 (O_1034,N_47833,N_49430);
or UO_1035 (O_1035,N_46471,N_45109);
nor UO_1036 (O_1036,N_45872,N_47596);
nor UO_1037 (O_1037,N_46463,N_45131);
nor UO_1038 (O_1038,N_46112,N_45825);
or UO_1039 (O_1039,N_49619,N_48393);
nand UO_1040 (O_1040,N_45700,N_45021);
or UO_1041 (O_1041,N_46790,N_46009);
or UO_1042 (O_1042,N_45112,N_45343);
or UO_1043 (O_1043,N_47694,N_45574);
or UO_1044 (O_1044,N_48912,N_46968);
and UO_1045 (O_1045,N_47203,N_49274);
nor UO_1046 (O_1046,N_48710,N_48782);
xnor UO_1047 (O_1047,N_47249,N_49148);
nand UO_1048 (O_1048,N_45330,N_45740);
nor UO_1049 (O_1049,N_46162,N_46703);
nand UO_1050 (O_1050,N_48681,N_47992);
or UO_1051 (O_1051,N_45243,N_47849);
and UO_1052 (O_1052,N_45717,N_49813);
xnor UO_1053 (O_1053,N_45931,N_45325);
nand UO_1054 (O_1054,N_46438,N_49675);
xnor UO_1055 (O_1055,N_49092,N_45084);
nand UO_1056 (O_1056,N_45020,N_45756);
or UO_1057 (O_1057,N_48074,N_47669);
nor UO_1058 (O_1058,N_49197,N_45000);
or UO_1059 (O_1059,N_48064,N_46026);
xnor UO_1060 (O_1060,N_45217,N_47756);
or UO_1061 (O_1061,N_48554,N_48059);
nand UO_1062 (O_1062,N_49147,N_47674);
nor UO_1063 (O_1063,N_46157,N_48043);
or UO_1064 (O_1064,N_46594,N_46006);
and UO_1065 (O_1065,N_49141,N_47475);
and UO_1066 (O_1066,N_46210,N_49556);
xnor UO_1067 (O_1067,N_49332,N_45710);
nor UO_1068 (O_1068,N_49164,N_49810);
nor UO_1069 (O_1069,N_45165,N_49683);
xnor UO_1070 (O_1070,N_49501,N_46759);
nand UO_1071 (O_1071,N_45622,N_49128);
and UO_1072 (O_1072,N_49840,N_46116);
nor UO_1073 (O_1073,N_47982,N_46989);
xnor UO_1074 (O_1074,N_49952,N_48243);
or UO_1075 (O_1075,N_45722,N_47190);
nor UO_1076 (O_1076,N_46970,N_48242);
or UO_1077 (O_1077,N_45026,N_46123);
nand UO_1078 (O_1078,N_48238,N_49047);
nor UO_1079 (O_1079,N_45183,N_48786);
or UO_1080 (O_1080,N_46986,N_49032);
and UO_1081 (O_1081,N_47090,N_46967);
or UO_1082 (O_1082,N_49747,N_46043);
xnor UO_1083 (O_1083,N_49551,N_46398);
and UO_1084 (O_1084,N_46972,N_45792);
or UO_1085 (O_1085,N_47951,N_47083);
xnor UO_1086 (O_1086,N_49420,N_47284);
and UO_1087 (O_1087,N_47569,N_48294);
and UO_1088 (O_1088,N_46282,N_46789);
or UO_1089 (O_1089,N_47308,N_47548);
and UO_1090 (O_1090,N_48646,N_47654);
or UO_1091 (O_1091,N_49953,N_49670);
and UO_1092 (O_1092,N_45014,N_49822);
or UO_1093 (O_1093,N_47362,N_47579);
and UO_1094 (O_1094,N_46617,N_48669);
or UO_1095 (O_1095,N_47152,N_48968);
nor UO_1096 (O_1096,N_47286,N_45174);
xor UO_1097 (O_1097,N_48199,N_46907);
and UO_1098 (O_1098,N_49181,N_46048);
nand UO_1099 (O_1099,N_47589,N_48347);
xnor UO_1100 (O_1100,N_48795,N_46780);
or UO_1101 (O_1101,N_47159,N_47448);
nor UO_1102 (O_1102,N_49380,N_49224);
or UO_1103 (O_1103,N_46520,N_46890);
xor UO_1104 (O_1104,N_46208,N_48679);
nor UO_1105 (O_1105,N_48153,N_48133);
or UO_1106 (O_1106,N_49894,N_49766);
and UO_1107 (O_1107,N_47141,N_49076);
nand UO_1108 (O_1108,N_48948,N_49402);
nor UO_1109 (O_1109,N_49275,N_47725);
or UO_1110 (O_1110,N_49025,N_48162);
nand UO_1111 (O_1111,N_48829,N_47767);
and UO_1112 (O_1112,N_46681,N_45445);
nor UO_1113 (O_1113,N_46220,N_46388);
xnor UO_1114 (O_1114,N_48368,N_45273);
xor UO_1115 (O_1115,N_47678,N_45111);
or UO_1116 (O_1116,N_45672,N_47611);
or UO_1117 (O_1117,N_49272,N_46639);
xor UO_1118 (O_1118,N_45884,N_45597);
xor UO_1119 (O_1119,N_45002,N_48489);
nor UO_1120 (O_1120,N_45810,N_46211);
xor UO_1121 (O_1121,N_48593,N_49890);
or UO_1122 (O_1122,N_46169,N_49069);
and UO_1123 (O_1123,N_49244,N_49152);
nand UO_1124 (O_1124,N_47305,N_49648);
or UO_1125 (O_1125,N_46619,N_45669);
xor UO_1126 (O_1126,N_46190,N_48035);
nor UO_1127 (O_1127,N_49549,N_47057);
and UO_1128 (O_1128,N_45844,N_45936);
nor UO_1129 (O_1129,N_49835,N_48320);
and UO_1130 (O_1130,N_46409,N_45155);
or UO_1131 (O_1131,N_45342,N_47793);
nor UO_1132 (O_1132,N_49177,N_45869);
xor UO_1133 (O_1133,N_49106,N_49787);
nand UO_1134 (O_1134,N_49194,N_49564);
nand UO_1135 (O_1135,N_47688,N_45925);
xor UO_1136 (O_1136,N_47402,N_48143);
nand UO_1137 (O_1137,N_47378,N_48240);
nand UO_1138 (O_1138,N_47675,N_49414);
and UO_1139 (O_1139,N_46039,N_49261);
and UO_1140 (O_1140,N_46060,N_47425);
or UO_1141 (O_1141,N_45573,N_48385);
and UO_1142 (O_1142,N_45153,N_49082);
and UO_1143 (O_1143,N_47243,N_48437);
and UO_1144 (O_1144,N_46256,N_46985);
nand UO_1145 (O_1145,N_46867,N_46503);
and UO_1146 (O_1146,N_48260,N_47783);
nand UO_1147 (O_1147,N_48424,N_46864);
nand UO_1148 (O_1148,N_45612,N_49654);
xnor UO_1149 (O_1149,N_45547,N_48259);
and UO_1150 (O_1150,N_47774,N_49717);
xnor UO_1151 (O_1151,N_49489,N_47068);
nand UO_1152 (O_1152,N_48488,N_49831);
xor UO_1153 (O_1153,N_49327,N_48841);
and UO_1154 (O_1154,N_47029,N_49201);
nor UO_1155 (O_1155,N_47868,N_46894);
nor UO_1156 (O_1156,N_47494,N_46022);
nor UO_1157 (O_1157,N_46421,N_46523);
nor UO_1158 (O_1158,N_47603,N_46526);
nor UO_1159 (O_1159,N_49480,N_47018);
nor UO_1160 (O_1160,N_48904,N_48311);
and UO_1161 (O_1161,N_48085,N_46066);
xor UO_1162 (O_1162,N_47289,N_48090);
or UO_1163 (O_1163,N_48267,N_47769);
or UO_1164 (O_1164,N_45238,N_45701);
nor UO_1165 (O_1165,N_48446,N_48021);
xnor UO_1166 (O_1166,N_48481,N_48036);
nand UO_1167 (O_1167,N_45826,N_49657);
nor UO_1168 (O_1168,N_45492,N_47505);
xnor UO_1169 (O_1169,N_46566,N_48060);
nor UO_1170 (O_1170,N_46016,N_46276);
and UO_1171 (O_1171,N_47733,N_45413);
nor UO_1172 (O_1172,N_46088,N_45144);
xor UO_1173 (O_1173,N_45891,N_48148);
and UO_1174 (O_1174,N_49671,N_48466);
and UO_1175 (O_1175,N_46937,N_46071);
nor UO_1176 (O_1176,N_47288,N_48622);
or UO_1177 (O_1177,N_48176,N_47527);
xor UO_1178 (O_1178,N_49709,N_46616);
nor UO_1179 (O_1179,N_47638,N_45063);
nand UO_1180 (O_1180,N_46142,N_45707);
and UO_1181 (O_1181,N_49496,N_47333);
and UO_1182 (O_1182,N_45119,N_47463);
xor UO_1183 (O_1183,N_48703,N_49404);
and UO_1184 (O_1184,N_48274,N_49752);
or UO_1185 (O_1185,N_49749,N_49093);
nand UO_1186 (O_1186,N_49796,N_49046);
xor UO_1187 (O_1187,N_45854,N_45696);
nor UO_1188 (O_1188,N_45141,N_49490);
and UO_1189 (O_1189,N_47702,N_48142);
nor UO_1190 (O_1190,N_45978,N_45058);
xnor UO_1191 (O_1191,N_46999,N_48492);
nand UO_1192 (O_1192,N_47671,N_46782);
nor UO_1193 (O_1193,N_48336,N_49034);
and UO_1194 (O_1194,N_47062,N_45175);
and UO_1195 (O_1195,N_48917,N_48843);
xor UO_1196 (O_1196,N_49725,N_48514);
and UO_1197 (O_1197,N_48092,N_46363);
xor UO_1198 (O_1198,N_45516,N_45446);
and UO_1199 (O_1199,N_46956,N_45148);
xnor UO_1200 (O_1200,N_49779,N_45437);
and UO_1201 (O_1201,N_46892,N_45467);
and UO_1202 (O_1202,N_48129,N_47961);
xor UO_1203 (O_1203,N_45695,N_49702);
or UO_1204 (O_1204,N_48103,N_47967);
or UO_1205 (O_1205,N_49472,N_46412);
and UO_1206 (O_1206,N_45292,N_49096);
nor UO_1207 (O_1207,N_48124,N_49668);
or UO_1208 (O_1208,N_49505,N_45976);
and UO_1209 (O_1209,N_47906,N_48803);
or UO_1210 (O_1210,N_46996,N_45145);
and UO_1211 (O_1211,N_47207,N_48617);
or UO_1212 (O_1212,N_46061,N_48585);
nor UO_1213 (O_1213,N_48663,N_45181);
or UO_1214 (O_1214,N_48615,N_47405);
or UO_1215 (O_1215,N_47923,N_47202);
and UO_1216 (O_1216,N_46742,N_46666);
nor UO_1217 (O_1217,N_47229,N_47088);
nor UO_1218 (O_1218,N_46578,N_45937);
or UO_1219 (O_1219,N_48777,N_49866);
and UO_1220 (O_1220,N_47872,N_49162);
and UO_1221 (O_1221,N_49297,N_46857);
nand UO_1222 (O_1222,N_48096,N_49343);
nand UO_1223 (O_1223,N_45836,N_49474);
and UO_1224 (O_1224,N_48362,N_46158);
or UO_1225 (O_1225,N_46606,N_48763);
or UO_1226 (O_1226,N_45697,N_45494);
nor UO_1227 (O_1227,N_46604,N_45366);
or UO_1228 (O_1228,N_48144,N_49346);
xnor UO_1229 (O_1229,N_46536,N_47184);
and UO_1230 (O_1230,N_45808,N_45599);
xnor UO_1231 (O_1231,N_45687,N_46340);
or UO_1232 (O_1232,N_48952,N_49608);
and UO_1233 (O_1233,N_45191,N_47080);
nand UO_1234 (O_1234,N_47942,N_49305);
nand UO_1235 (O_1235,N_46458,N_45464);
xnor UO_1236 (O_1236,N_49214,N_46873);
nand UO_1237 (O_1237,N_45987,N_49470);
nand UO_1238 (O_1238,N_48269,N_46627);
xnor UO_1239 (O_1239,N_47223,N_48775);
nor UO_1240 (O_1240,N_49465,N_49690);
xor UO_1241 (O_1241,N_45278,N_45225);
xnor UO_1242 (O_1242,N_45157,N_46905);
xor UO_1243 (O_1243,N_45461,N_45486);
or UO_1244 (O_1244,N_47834,N_49079);
nand UO_1245 (O_1245,N_45098,N_45557);
xor UO_1246 (O_1246,N_46777,N_47343);
xnor UO_1247 (O_1247,N_48284,N_49918);
and UO_1248 (O_1248,N_47994,N_48528);
or UO_1249 (O_1249,N_45984,N_45105);
or UO_1250 (O_1250,N_49336,N_46045);
nor UO_1251 (O_1251,N_48012,N_47261);
or UO_1252 (O_1252,N_48629,N_46676);
or UO_1253 (O_1253,N_49088,N_47258);
xnor UO_1254 (O_1254,N_48643,N_48397);
and UO_1255 (O_1255,N_45443,N_45244);
nand UO_1256 (O_1256,N_45663,N_48304);
nor UO_1257 (O_1257,N_49325,N_46767);
xnor UO_1258 (O_1258,N_48792,N_47111);
nor UO_1259 (O_1259,N_48464,N_47541);
or UO_1260 (O_1260,N_45023,N_49486);
xnor UO_1261 (O_1261,N_48254,N_46810);
or UO_1262 (O_1262,N_47348,N_46893);
nand UO_1263 (O_1263,N_49375,N_46935);
nor UO_1264 (O_1264,N_48001,N_45357);
and UO_1265 (O_1265,N_45215,N_47344);
xor UO_1266 (O_1266,N_47551,N_46289);
nand UO_1267 (O_1267,N_49488,N_46783);
nand UO_1268 (O_1268,N_49028,N_46367);
or UO_1269 (O_1269,N_45618,N_47365);
xor UO_1270 (O_1270,N_45920,N_46253);
or UO_1271 (O_1271,N_49394,N_45580);
or UO_1272 (O_1272,N_48630,N_46973);
xnor UO_1273 (O_1273,N_46339,N_47386);
and UO_1274 (O_1274,N_45914,N_46231);
xor UO_1275 (O_1275,N_48844,N_49525);
or UO_1276 (O_1276,N_46252,N_45314);
nor UO_1277 (O_1277,N_48037,N_47949);
and UO_1278 (O_1278,N_46859,N_48247);
nor UO_1279 (O_1279,N_49788,N_47914);
nand UO_1280 (O_1280,N_48130,N_47064);
or UO_1281 (O_1281,N_49728,N_46976);
or UO_1282 (O_1282,N_48873,N_47098);
xor UO_1283 (O_1283,N_45771,N_48476);
nand UO_1284 (O_1284,N_49931,N_46483);
nand UO_1285 (O_1285,N_47347,N_45210);
and UO_1286 (O_1286,N_49510,N_45586);
xnor UO_1287 (O_1287,N_49967,N_48477);
xor UO_1288 (O_1288,N_45723,N_46505);
nor UO_1289 (O_1289,N_45954,N_46738);
and UO_1290 (O_1290,N_45739,N_48714);
or UO_1291 (O_1291,N_45550,N_47324);
nor UO_1292 (O_1292,N_45822,N_49755);
xnor UO_1293 (O_1293,N_47970,N_48337);
xor UO_1294 (O_1294,N_45321,N_48574);
xnor UO_1295 (O_1295,N_45216,N_47209);
or UO_1296 (O_1296,N_48876,N_49754);
or UO_1297 (O_1297,N_45590,N_45159);
and UO_1298 (O_1298,N_46219,N_47912);
nor UO_1299 (O_1299,N_45104,N_46337);
or UO_1300 (O_1300,N_49529,N_46557);
and UO_1301 (O_1301,N_45904,N_45653);
and UO_1302 (O_1302,N_48023,N_48905);
nand UO_1303 (O_1303,N_45473,N_47995);
or UO_1304 (O_1304,N_47124,N_45768);
xnor UO_1305 (O_1305,N_49886,N_45514);
xor UO_1306 (O_1306,N_47493,N_48516);
nor UO_1307 (O_1307,N_45743,N_49158);
or UO_1308 (O_1308,N_47051,N_49271);
nor UO_1309 (O_1309,N_46623,N_47752);
nor UO_1310 (O_1310,N_47161,N_48566);
nor UO_1311 (O_1311,N_49870,N_45385);
nand UO_1312 (O_1312,N_45362,N_45079);
nor UO_1313 (O_1313,N_49892,N_48586);
nand UO_1314 (O_1314,N_47278,N_47301);
xnor UO_1315 (O_1315,N_47876,N_49878);
nand UO_1316 (O_1316,N_49605,N_46089);
xnor UO_1317 (O_1317,N_47508,N_48456);
nand UO_1318 (O_1318,N_47267,N_47555);
xnor UO_1319 (O_1319,N_47136,N_45152);
or UO_1320 (O_1320,N_47779,N_45009);
or UO_1321 (O_1321,N_48024,N_47245);
nand UO_1322 (O_1322,N_47310,N_48644);
or UO_1323 (O_1323,N_46058,N_45507);
and UO_1324 (O_1324,N_49729,N_47919);
or UO_1325 (O_1325,N_47780,N_46124);
or UO_1326 (O_1326,N_47497,N_46592);
nor UO_1327 (O_1327,N_49701,N_49987);
or UO_1328 (O_1328,N_48821,N_46092);
nand UO_1329 (O_1329,N_45115,N_46126);
nor UO_1330 (O_1330,N_48107,N_49494);
or UO_1331 (O_1331,N_49471,N_45539);
or UO_1332 (O_1332,N_49612,N_49384);
nand UO_1333 (O_1333,N_46153,N_47272);
nand UO_1334 (O_1334,N_46620,N_47873);
nand UO_1335 (O_1335,N_49487,N_46122);
or UO_1336 (O_1336,N_46138,N_47387);
nor UO_1337 (O_1337,N_45689,N_47496);
or UO_1338 (O_1338,N_45091,N_46587);
xnor UO_1339 (O_1339,N_49333,N_46046);
xnor UO_1340 (O_1340,N_46033,N_45229);
and UO_1341 (O_1341,N_48577,N_49802);
nor UO_1342 (O_1342,N_47350,N_49898);
or UO_1343 (O_1343,N_45186,N_48756);
and UO_1344 (O_1344,N_49836,N_45634);
and UO_1345 (O_1345,N_48721,N_45194);
nor UO_1346 (O_1346,N_46830,N_48552);
xnor UO_1347 (O_1347,N_49368,N_49242);
and UO_1348 (O_1348,N_46449,N_45247);
xnor UO_1349 (O_1349,N_49606,N_45994);
nor UO_1350 (O_1350,N_49022,N_48664);
or UO_1351 (O_1351,N_49644,N_46661);
nand UO_1352 (O_1352,N_48845,N_47672);
or UO_1353 (O_1353,N_46090,N_48849);
nand UO_1354 (O_1354,N_48367,N_47613);
and UO_1355 (O_1355,N_48198,N_48033);
xnor UO_1356 (O_1356,N_46658,N_49282);
and UO_1357 (O_1357,N_46645,N_48484);
nor UO_1358 (O_1358,N_48220,N_45650);
and UO_1359 (O_1359,N_49574,N_48696);
and UO_1360 (O_1360,N_47853,N_48783);
and UO_1361 (O_1361,N_47381,N_47996);
nand UO_1362 (O_1362,N_46670,N_45212);
xnor UO_1363 (O_1363,N_47911,N_45390);
nor UO_1364 (O_1364,N_48431,N_47498);
nand UO_1365 (O_1365,N_47575,N_47990);
xnor UO_1366 (O_1366,N_49330,N_49051);
nor UO_1367 (O_1367,N_48546,N_47428);
and UO_1368 (O_1368,N_46598,N_47097);
or UO_1369 (O_1369,N_48379,N_47647);
xor UO_1370 (O_1370,N_45688,N_49994);
and UO_1371 (O_1371,N_46684,N_48602);
or UO_1372 (O_1372,N_46700,N_46377);
nor UO_1373 (O_1373,N_49134,N_48223);
nor UO_1374 (O_1374,N_49338,N_49324);
nor UO_1375 (O_1375,N_47610,N_46224);
nor UO_1376 (O_1376,N_46760,N_49604);
nand UO_1377 (O_1377,N_47570,N_46710);
and UO_1378 (O_1378,N_46279,N_46650);
or UO_1379 (O_1379,N_49848,N_48044);
nor UO_1380 (O_1380,N_47520,N_48184);
nand UO_1381 (O_1381,N_46402,N_48539);
and UO_1382 (O_1382,N_48429,N_45751);
and UO_1383 (O_1383,N_47585,N_49014);
nand UO_1384 (O_1384,N_49329,N_47250);
or UO_1385 (O_1385,N_49273,N_48600);
xor UO_1386 (O_1386,N_47880,N_45907);
nor UO_1387 (O_1387,N_49692,N_48770);
nor UO_1388 (O_1388,N_45985,N_48283);
and UO_1389 (O_1389,N_45683,N_45125);
xor UO_1390 (O_1390,N_47898,N_45053);
nor UO_1391 (O_1391,N_46073,N_47511);
xnor UO_1392 (O_1392,N_48953,N_48995);
or UO_1393 (O_1393,N_46374,N_46804);
xnor UO_1394 (O_1394,N_49381,N_48047);
nor UO_1395 (O_1395,N_46393,N_49043);
nor UO_1396 (O_1396,N_45051,N_45270);
xnor UO_1397 (O_1397,N_45955,N_47268);
nand UO_1398 (O_1398,N_48420,N_47908);
and UO_1399 (O_1399,N_46524,N_48334);
xor UO_1400 (O_1400,N_49955,N_47231);
nor UO_1401 (O_1401,N_46614,N_49944);
xnor UO_1402 (O_1402,N_48604,N_49602);
and UO_1403 (O_1403,N_46562,N_49030);
xnor UO_1404 (O_1404,N_49991,N_45088);
and UO_1405 (O_1405,N_48239,N_45818);
and UO_1406 (O_1406,N_47432,N_48702);
nand UO_1407 (O_1407,N_45851,N_45734);
nor UO_1408 (O_1408,N_49883,N_45032);
or UO_1409 (O_1409,N_46251,N_48211);
nand UO_1410 (O_1410,N_47714,N_49842);
and UO_1411 (O_1411,N_45926,N_48960);
nor UO_1412 (O_1412,N_46203,N_47670);
xor UO_1413 (O_1413,N_49215,N_49706);
nor UO_1414 (O_1414,N_48002,N_45322);
nor UO_1415 (O_1415,N_47100,N_45556);
nand UO_1416 (O_1416,N_49589,N_45749);
or UO_1417 (O_1417,N_47484,N_48390);
nand UO_1418 (O_1418,N_47279,N_47689);
or UO_1419 (O_1419,N_48830,N_49263);
nand UO_1420 (O_1420,N_49475,N_45898);
xnor UO_1421 (O_1421,N_45205,N_46443);
or UO_1422 (O_1422,N_45300,N_49035);
nor UO_1423 (O_1423,N_48788,N_46590);
and UO_1424 (O_1424,N_45956,N_49801);
xnor UO_1425 (O_1425,N_47775,N_49070);
nand UO_1426 (O_1426,N_48226,N_48418);
xor UO_1427 (O_1427,N_45693,N_45479);
nor UO_1428 (O_1428,N_48098,N_48784);
nor UO_1429 (O_1429,N_46352,N_48359);
nor UO_1430 (O_1430,N_49090,N_49947);
nor UO_1431 (O_1431,N_48939,N_48875);
nand UO_1432 (O_1432,N_49590,N_47679);
xnor UO_1433 (O_1433,N_49913,N_47650);
and UO_1434 (O_1434,N_49328,N_46008);
and UO_1435 (O_1435,N_45676,N_49481);
nand UO_1436 (O_1436,N_48031,N_47943);
nand UO_1437 (O_1437,N_45395,N_49882);
nand UO_1438 (O_1438,N_45821,N_47837);
nand UO_1439 (O_1439,N_49107,N_46415);
nand UO_1440 (O_1440,N_48942,N_47743);
xor UO_1441 (O_1441,N_49137,N_45043);
and UO_1442 (O_1442,N_48066,N_46063);
and UO_1443 (O_1443,N_47792,N_45282);
xnor UO_1444 (O_1444,N_47139,N_48757);
and UO_1445 (O_1445,N_48101,N_45315);
nor UO_1446 (O_1446,N_48880,N_45170);
or UO_1447 (O_1447,N_46069,N_49798);
xor UO_1448 (O_1448,N_48073,N_48680);
or UO_1449 (O_1449,N_48478,N_47074);
nand UO_1450 (O_1450,N_48854,N_45506);
or UO_1451 (O_1451,N_48595,N_46342);
and UO_1452 (O_1452,N_48535,N_46649);
nor UO_1453 (O_1453,N_46034,N_47812);
and UO_1454 (O_1454,N_48887,N_46424);
nand UO_1455 (O_1455,N_47165,N_48356);
nor UO_1456 (O_1456,N_48458,N_49715);
nor UO_1457 (O_1457,N_45354,N_45690);
nand UO_1458 (O_1458,N_49895,N_45436);
xnor UO_1459 (O_1459,N_45337,N_45025);
xor UO_1460 (O_1460,N_48084,N_46647);
xor UO_1461 (O_1461,N_49223,N_45775);
nor UO_1462 (O_1462,N_48028,N_48737);
xor UO_1463 (O_1463,N_46982,N_45675);
nand UO_1464 (O_1464,N_46404,N_46075);
xnor UO_1465 (O_1465,N_48519,N_45895);
xor UO_1466 (O_1466,N_48480,N_46558);
xor UO_1467 (O_1467,N_45242,N_47974);
nand UO_1468 (O_1468,N_47550,N_48623);
or UO_1469 (O_1469,N_45280,N_47731);
and UO_1470 (O_1470,N_45562,N_46839);
nand UO_1471 (O_1471,N_45246,N_48911);
xnor UO_1472 (O_1472,N_45260,N_46625);
or UO_1473 (O_1473,N_47851,N_49518);
nor UO_1474 (O_1474,N_48150,N_46997);
and UO_1475 (O_1475,N_47396,N_48055);
or UO_1476 (O_1476,N_48773,N_49618);
nand UO_1477 (O_1477,N_48128,N_48276);
or UO_1478 (O_1478,N_45757,N_48779);
and UO_1479 (O_1479,N_45495,N_47532);
nor UO_1480 (O_1480,N_46436,N_47634);
nand UO_1481 (O_1481,N_45132,N_46884);
xor UO_1482 (O_1482,N_48182,N_45274);
xnor UO_1483 (O_1483,N_47247,N_49759);
and UO_1484 (O_1484,N_47126,N_47358);
or UO_1485 (O_1485,N_48270,N_45748);
nand UO_1486 (O_1486,N_46507,N_45600);
or UO_1487 (O_1487,N_48154,N_49585);
or UO_1488 (O_1488,N_46307,N_48046);
xor UO_1489 (O_1489,N_45410,N_49603);
or UO_1490 (O_1490,N_48268,N_48501);
xor UO_1491 (O_1491,N_45787,N_47842);
nand UO_1492 (O_1492,N_47118,N_47999);
and UO_1493 (O_1493,N_49784,N_49502);
nor UO_1494 (O_1494,N_48752,N_48704);
nand UO_1495 (O_1495,N_49667,N_47244);
xor UO_1496 (O_1496,N_49171,N_49538);
or UO_1497 (O_1497,N_45203,N_47963);
or UO_1498 (O_1498,N_48228,N_46055);
or UO_1499 (O_1499,N_45666,N_47395);
and UO_1500 (O_1500,N_47373,N_47330);
and UO_1501 (O_1501,N_49732,N_49131);
and UO_1502 (O_1502,N_47971,N_47802);
nand UO_1503 (O_1503,N_47740,N_49315);
nor UO_1504 (O_1504,N_47150,N_45380);
and UO_1505 (O_1505,N_47241,N_48250);
and UO_1506 (O_1506,N_47337,N_45780);
xnor UO_1507 (O_1507,N_48316,N_46739);
nor UO_1508 (O_1508,N_47692,N_47935);
or UO_1509 (O_1509,N_48780,N_45369);
xnor UO_1510 (O_1510,N_46896,N_46793);
xnor UO_1511 (O_1511,N_48751,N_47327);
nand UO_1512 (O_1512,N_49756,N_49169);
nand UO_1513 (O_1513,N_48861,N_47013);
or UO_1514 (O_1514,N_47561,N_47007);
and UO_1515 (O_1515,N_45998,N_45420);
and UO_1516 (O_1516,N_49758,N_47565);
nand UO_1517 (O_1517,N_45404,N_45399);
xnor UO_1518 (O_1518,N_47839,N_46086);
xor UO_1519 (O_1519,N_47240,N_48541);
or UO_1520 (O_1520,N_49493,N_45715);
nand UO_1521 (O_1521,N_49543,N_48666);
nor UO_1522 (O_1522,N_47580,N_49007);
or UO_1523 (O_1523,N_45790,N_46445);
and UO_1524 (O_1524,N_46391,N_47861);
nand UO_1525 (O_1525,N_48774,N_47878);
nor UO_1526 (O_1526,N_46400,N_48327);
nor UO_1527 (O_1527,N_49580,N_48262);
xnor UO_1528 (O_1528,N_47212,N_47011);
nand UO_1529 (O_1529,N_45744,N_47915);
nor UO_1530 (O_1530,N_45442,N_49986);
and UO_1531 (O_1531,N_48179,N_46966);
xnor UO_1532 (O_1532,N_47560,N_47576);
or UO_1533 (O_1533,N_49188,N_45591);
or UO_1534 (O_1534,N_46556,N_46728);
or UO_1535 (O_1535,N_46934,N_47787);
xor UO_1536 (O_1536,N_47998,N_49248);
nand UO_1537 (O_1537,N_49775,N_49075);
nor UO_1538 (O_1538,N_48864,N_47353);
nor UO_1539 (O_1539,N_47658,N_47372);
xor UO_1540 (O_1540,N_48532,N_48415);
or UO_1541 (O_1541,N_47179,N_45200);
and UO_1542 (O_1542,N_48989,N_45582);
or UO_1543 (O_1543,N_47956,N_46769);
and UO_1544 (O_1544,N_45595,N_45620);
and UO_1545 (O_1545,N_46774,N_49026);
or UO_1546 (O_1546,N_46977,N_46925);
xor UO_1547 (O_1547,N_46856,N_46263);
and UO_1548 (O_1548,N_47458,N_47266);
or UO_1549 (O_1549,N_48388,N_48360);
xor UO_1550 (O_1550,N_46705,N_46603);
xnor UO_1551 (O_1551,N_49512,N_48421);
xor UO_1552 (O_1552,N_46271,N_45754);
nand UO_1553 (O_1553,N_48376,N_48755);
nand UO_1554 (O_1554,N_49163,N_48517);
xnor UO_1555 (O_1555,N_46875,N_46501);
and UO_1556 (O_1556,N_47127,N_45452);
or UO_1557 (O_1557,N_47246,N_45281);
xor UO_1558 (O_1558,N_49643,N_46781);
or UO_1559 (O_1559,N_45074,N_46209);
or UO_1560 (O_1560,N_45450,N_45497);
xor UO_1561 (O_1561,N_47979,N_49662);
and UO_1562 (O_1562,N_48159,N_47482);
nor UO_1563 (O_1563,N_48863,N_48769);
or UO_1564 (O_1564,N_47125,N_45886);
or UO_1565 (O_1565,N_45522,N_46923);
or UO_1566 (O_1566,N_47938,N_48091);
nor UO_1567 (O_1567,N_45085,N_48840);
or UO_1568 (O_1568,N_46442,N_45839);
or UO_1569 (O_1569,N_46541,N_45444);
nand UO_1570 (O_1570,N_46586,N_46351);
xnor UO_1571 (O_1571,N_45665,N_47120);
and UO_1572 (O_1572,N_45287,N_46539);
or UO_1573 (O_1573,N_48258,N_48291);
nor UO_1574 (O_1574,N_47452,N_47354);
nand UO_1575 (O_1575,N_45277,N_45703);
or UO_1576 (O_1576,N_47786,N_48520);
or UO_1577 (O_1577,N_48207,N_49104);
and UO_1578 (O_1578,N_45069,N_47933);
nand UO_1579 (O_1579,N_45086,N_45402);
xor UO_1580 (O_1580,N_48620,N_46754);
nor UO_1581 (O_1581,N_46762,N_46662);
nand UO_1582 (O_1582,N_45543,N_47593);
and UO_1583 (O_1583,N_48674,N_49763);
nand UO_1584 (O_1584,N_48372,N_46403);
nand UO_1585 (O_1585,N_47106,N_46215);
or UO_1586 (O_1586,N_45537,N_46468);
nor UO_1587 (O_1587,N_46543,N_48089);
or UO_1588 (O_1588,N_49441,N_49138);
nand UO_1589 (O_1589,N_47054,N_45623);
and UO_1590 (O_1590,N_47535,N_45449);
xor UO_1591 (O_1591,N_45758,N_45015);
and UO_1592 (O_1592,N_48709,N_45639);
or UO_1593 (O_1593,N_49266,N_46477);
and UO_1594 (O_1594,N_47443,N_46200);
and UO_1595 (O_1595,N_49905,N_48459);
and UO_1596 (O_1596,N_49166,N_46038);
or UO_1597 (O_1597,N_45527,N_49559);
xor UO_1598 (O_1598,N_45431,N_49438);
nor UO_1599 (O_1599,N_47171,N_49849);
nand UO_1600 (O_1600,N_45383,N_46936);
xor UO_1601 (O_1601,N_49926,N_49862);
xor UO_1602 (O_1602,N_45982,N_45655);
and UO_1603 (O_1603,N_46394,N_49386);
nor UO_1604 (O_1604,N_46564,N_45501);
xor UO_1605 (O_1605,N_45368,N_49948);
and UO_1606 (O_1606,N_46959,N_47424);
or UO_1607 (O_1607,N_45685,N_46371);
or UO_1608 (O_1608,N_45235,N_47599);
xnor UO_1609 (O_1609,N_46018,N_48402);
nand UO_1610 (O_1610,N_46851,N_47531);
or UO_1611 (O_1611,N_47434,N_49015);
nor UO_1612 (O_1612,N_47836,N_45010);
nand UO_1613 (O_1613,N_49406,N_47973);
and UO_1614 (O_1614,N_48598,N_45221);
nor UO_1615 (O_1615,N_48597,N_49229);
nor UO_1616 (O_1616,N_48619,N_45013);
nor UO_1617 (O_1617,N_48531,N_48608);
and UO_1618 (O_1618,N_48138,N_45725);
and UO_1619 (O_1619,N_48237,N_45048);
and UO_1620 (O_1620,N_49245,N_45090);
or UO_1621 (O_1621,N_49230,N_49719);
or UO_1622 (O_1622,N_49703,N_45952);
nor UO_1623 (O_1623,N_49859,N_47233);
nor UO_1624 (O_1624,N_45644,N_45231);
nand UO_1625 (O_1625,N_46800,N_49151);
nor UO_1626 (O_1626,N_49553,N_46846);
xor UO_1627 (O_1627,N_48017,N_48812);
and UO_1628 (O_1628,N_45140,N_46067);
nor UO_1629 (O_1629,N_48344,N_49218);
nand UO_1630 (O_1630,N_49969,N_48838);
or UO_1631 (O_1631,N_46554,N_46301);
nand UO_1632 (O_1632,N_46943,N_47958);
xor UO_1633 (O_1633,N_47806,N_48088);
nor UO_1634 (O_1634,N_45508,N_47091);
xnor UO_1635 (O_1635,N_46193,N_49016);
and UO_1636 (O_1636,N_46486,N_49625);
and UO_1637 (O_1637,N_47519,N_49478);
and UO_1638 (O_1638,N_49036,N_47525);
nand UO_1639 (O_1639,N_48694,N_49175);
or UO_1640 (O_1640,N_46540,N_47959);
and UO_1641 (O_1641,N_49145,N_48375);
nand UO_1642 (O_1642,N_46516,N_48536);
xnor UO_1643 (O_1643,N_47789,N_47265);
nor UO_1644 (O_1644,N_45677,N_47617);
nand UO_1645 (O_1645,N_46450,N_48973);
or UO_1646 (O_1646,N_46241,N_45652);
nand UO_1647 (O_1647,N_46261,N_45991);
nand UO_1648 (O_1648,N_49360,N_45080);
nand UO_1649 (O_1649,N_48909,N_45481);
nand UO_1650 (O_1650,N_46535,N_45167);
xnor UO_1651 (O_1651,N_45959,N_48808);
xor UO_1652 (O_1652,N_49120,N_46312);
nand UO_1653 (O_1653,N_48164,N_45389);
or UO_1654 (O_1654,N_48325,N_48988);
nor UO_1655 (O_1655,N_46811,N_45668);
nand UO_1656 (O_1656,N_49293,N_46821);
and UO_1657 (O_1657,N_49837,N_48022);
nor UO_1658 (O_1658,N_48950,N_49027);
and UO_1659 (O_1659,N_45418,N_46803);
nor UO_1660 (O_1660,N_47121,N_45746);
or UO_1661 (O_1661,N_49519,N_48117);
nand UO_1662 (O_1662,N_46406,N_49640);
xnor UO_1663 (O_1663,N_46509,N_47385);
nand UO_1664 (O_1664,N_49409,N_45878);
nor UO_1665 (O_1665,N_46882,N_46612);
nand UO_1666 (O_1666,N_48483,N_46694);
nand UO_1667 (O_1667,N_48816,N_49232);
or UO_1668 (O_1668,N_46183,N_49805);
and UO_1669 (O_1669,N_46028,N_48847);
xnor UO_1670 (O_1670,N_49289,N_49373);
nand UO_1671 (O_1671,N_47140,N_48426);
xor UO_1672 (O_1672,N_49829,N_49841);
and UO_1673 (O_1673,N_48512,N_49833);
nor UO_1674 (O_1674,N_46115,N_47946);
or UO_1675 (O_1675,N_47228,N_47302);
or UO_1676 (O_1676,N_49997,N_46707);
nor UO_1677 (O_1677,N_46858,N_47323);
or UO_1678 (O_1678,N_48685,N_45223);
nor UO_1679 (O_1679,N_49367,N_48472);
and UO_1680 (O_1680,N_45162,N_48447);
and UO_1681 (O_1681,N_49078,N_45294);
nor UO_1682 (O_1682,N_48065,N_45230);
or UO_1683 (O_1683,N_48722,N_49125);
or UO_1684 (O_1684,N_48082,N_49388);
and UO_1685 (O_1685,N_47138,N_48958);
and UO_1686 (O_1686,N_46392,N_47515);
nand UO_1687 (O_1687,N_48605,N_45219);
or UO_1688 (O_1688,N_45526,N_46331);
and UO_1689 (O_1689,N_47028,N_47155);
nor UO_1690 (O_1690,N_46978,N_47838);
nand UO_1691 (O_1691,N_47953,N_46481);
and UO_1692 (O_1692,N_46192,N_46360);
nand UO_1693 (O_1693,N_48640,N_45793);
xor UO_1694 (O_1694,N_47319,N_47991);
or UO_1695 (O_1695,N_47815,N_46465);
and UO_1696 (O_1696,N_49928,N_48990);
or UO_1697 (O_1697,N_48557,N_48706);
nand UO_1698 (O_1698,N_48853,N_47283);
nand UO_1699 (O_1699,N_49198,N_46321);
nor UO_1700 (O_1700,N_46673,N_47439);
nor UO_1701 (O_1701,N_48601,N_49349);
nand UO_1702 (O_1702,N_47734,N_46470);
or UO_1703 (O_1703,N_48004,N_48027);
or UO_1704 (O_1704,N_45750,N_46417);
xor UO_1705 (O_1705,N_49499,N_48439);
nor UO_1706 (O_1706,N_48986,N_45624);
nor UO_1707 (O_1707,N_45804,N_45617);
nor UO_1708 (O_1708,N_47941,N_46324);
nand UO_1709 (O_1709,N_49190,N_48400);
or UO_1710 (O_1710,N_45935,N_47221);
and UO_1711 (O_1711,N_48570,N_49023);
or UO_1712 (O_1712,N_49000,N_45918);
nand UO_1713 (O_1713,N_47384,N_48813);
nor UO_1714 (O_1714,N_48425,N_45627);
and UO_1715 (O_1715,N_46874,N_45564);
or UO_1716 (O_1716,N_45916,N_49424);
nor UO_1717 (O_1717,N_47615,N_49410);
nor UO_1718 (O_1718,N_48099,N_48018);
nor UO_1719 (O_1719,N_45055,N_47465);
nand UO_1720 (O_1720,N_46384,N_46961);
xnor UO_1721 (O_1721,N_46350,N_47148);
and UO_1722 (O_1722,N_48493,N_45513);
xnor UO_1723 (O_1723,N_46425,N_49077);
xnor UO_1724 (O_1724,N_47388,N_48147);
nand UO_1725 (O_1725,N_46199,N_46349);
nand UO_1726 (O_1726,N_49807,N_45642);
nor UO_1727 (O_1727,N_47107,N_49697);
or UO_1728 (O_1728,N_46841,N_45671);
nand UO_1729 (O_1729,N_46772,N_46715);
or UO_1730 (O_1730,N_48000,N_49941);
nand UO_1731 (O_1731,N_49200,N_46506);
nand UO_1732 (O_1732,N_46359,N_47112);
nand UO_1733 (O_1733,N_47485,N_45799);
xor UO_1734 (O_1734,N_46898,N_49382);
nor UO_1735 (O_1735,N_47945,N_46065);
or UO_1736 (O_1736,N_48584,N_46007);
and UO_1737 (O_1737,N_48627,N_45549);
nand UO_1738 (O_1738,N_45453,N_47345);
nand UO_1739 (O_1739,N_49331,N_48366);
or UO_1740 (O_1740,N_45720,N_48261);
nand UO_1741 (O_1741,N_46000,N_48353);
nor UO_1742 (O_1742,N_46735,N_45572);
nor UO_1743 (O_1743,N_49464,N_47419);
nand UO_1744 (O_1744,N_45924,N_48191);
nand UO_1745 (O_1745,N_49936,N_48954);
or UO_1746 (O_1746,N_49780,N_47357);
and UO_1747 (O_1747,N_47607,N_46044);
nor UO_1748 (O_1748,N_45656,N_49909);
and UO_1749 (O_1749,N_49597,N_49786);
xor UO_1750 (O_1750,N_45054,N_46930);
nand UO_1751 (O_1751,N_48695,N_49066);
or UO_1752 (O_1752,N_45350,N_46164);
nand UO_1753 (O_1753,N_46686,N_45388);
xnor UO_1754 (O_1754,N_45812,N_48307);
xor UO_1755 (O_1755,N_49462,N_49350);
xnor UO_1756 (O_1756,N_46955,N_45041);
or UO_1757 (O_1757,N_47215,N_47189);
xor UO_1758 (O_1758,N_45083,N_45060);
nor UO_1759 (O_1759,N_46799,N_49960);
xnor UO_1760 (O_1760,N_45941,N_46624);
or UO_1761 (O_1761,N_49083,N_46813);
xor UO_1762 (O_1762,N_45912,N_46040);
xor UO_1763 (O_1763,N_49044,N_46601);
nor UO_1764 (O_1764,N_49560,N_49925);
nor UO_1765 (O_1765,N_48365,N_46493);
and UO_1766 (O_1766,N_48051,N_48723);
nand UO_1767 (O_1767,N_49970,N_46840);
nor UO_1768 (O_1768,N_49143,N_47653);
nor UO_1769 (O_1769,N_49187,N_48434);
nand UO_1770 (O_1770,N_49533,N_49221);
nor UO_1771 (O_1771,N_49891,N_49785);
nor UO_1772 (O_1772,N_46137,N_46838);
or UO_1773 (O_1773,N_46004,N_46003);
nor UO_1774 (O_1774,N_47174,N_46303);
or UO_1775 (O_1775,N_47784,N_47828);
or UO_1776 (O_1776,N_46571,N_48892);
xor UO_1777 (O_1777,N_46862,N_49900);
nor UO_1778 (O_1778,N_48208,N_49795);
and UO_1779 (O_1779,N_46019,N_48888);
xnor UO_1780 (O_1780,N_49993,N_49259);
xnor UO_1781 (O_1781,N_45117,N_46310);
xnor UO_1782 (O_1782,N_48568,N_48588);
nand UO_1783 (O_1783,N_48924,N_47562);
and UO_1784 (O_1784,N_47768,N_49591);
and UO_1785 (O_1785,N_46528,N_45199);
and UO_1786 (O_1786,N_49211,N_46699);
or UO_1787 (O_1787,N_45691,N_46390);
nand UO_1788 (O_1788,N_46519,N_46267);
nor UO_1789 (O_1789,N_48212,N_45880);
nand UO_1790 (O_1790,N_48928,N_49341);
nor UO_1791 (O_1791,N_47635,N_45328);
and UO_1792 (O_1792,N_45142,N_46072);
or UO_1793 (O_1793,N_46140,N_47022);
nor UO_1794 (O_1794,N_48363,N_49853);
xor UO_1795 (O_1795,N_46939,N_49204);
nor UO_1796 (O_1796,N_48591,N_46669);
xnor UO_1797 (O_1797,N_45724,N_49127);
nand UO_1798 (O_1798,N_48907,N_49973);
nor UO_1799 (O_1799,N_49102,N_48941);
and UO_1800 (O_1800,N_45913,N_49863);
and UO_1801 (O_1801,N_45258,N_49440);
or UO_1802 (O_1802,N_46704,N_46596);
and UO_1803 (O_1803,N_45263,N_48392);
or UO_1804 (O_1804,N_45596,N_47683);
and UO_1805 (O_1805,N_47193,N_49109);
nor UO_1806 (O_1806,N_48638,N_46278);
and UO_1807 (O_1807,N_49108,N_49773);
and UO_1808 (O_1808,N_49699,N_45024);
or UO_1809 (O_1809,N_47049,N_48836);
or UO_1810 (O_1810,N_46828,N_46602);
nand UO_1811 (O_1811,N_49072,N_45237);
xor UO_1812 (O_1812,N_45946,N_45532);
nor UO_1813 (O_1813,N_49240,N_49012);
and UO_1814 (O_1814,N_49385,N_48807);
xnor UO_1815 (O_1815,N_45641,N_48738);
nor UO_1816 (O_1816,N_45613,N_45708);
nand UO_1817 (O_1817,N_47177,N_45774);
nor UO_1818 (O_1818,N_46343,N_45103);
nand UO_1819 (O_1819,N_46659,N_45056);
and UO_1820 (O_1820,N_48014,N_48432);
nor UO_1821 (O_1821,N_45188,N_45988);
nand UO_1822 (O_1822,N_46906,N_46951);
xnor UO_1823 (O_1823,N_48152,N_47242);
nand UO_1824 (O_1824,N_48798,N_47269);
and UO_1825 (O_1825,N_47655,N_46547);
nor UO_1826 (O_1826,N_49578,N_48628);
xnor UO_1827 (O_1827,N_48522,N_49383);
and UO_1828 (O_1828,N_46644,N_46944);
or UO_1829 (O_1829,N_45732,N_49098);
and UO_1830 (O_1830,N_48503,N_49100);
or UO_1831 (O_1831,N_48445,N_49427);
and UO_1832 (O_1832,N_46187,N_47644);
or UO_1833 (O_1833,N_46461,N_46805);
nand UO_1834 (O_1834,N_45888,N_49116);
and UO_1835 (O_1835,N_46177,N_47648);
nand UO_1836 (O_1836,N_49689,N_49225);
nand UO_1837 (O_1837,N_46488,N_45570);
or UO_1838 (O_1838,N_48003,N_49911);
xnor UO_1839 (O_1839,N_45419,N_45160);
or UO_1840 (O_1840,N_47442,N_48851);
xor UO_1841 (O_1841,N_45883,N_47563);
and UO_1842 (O_1842,N_49442,N_48688);
nor UO_1843 (O_1843,N_45245,N_47002);
and UO_1844 (O_1844,N_49366,N_49306);
nand UO_1845 (O_1845,N_48470,N_47691);
and UO_1846 (O_1846,N_45667,N_46341);
xor UO_1847 (O_1847,N_46453,N_46637);
xor UO_1848 (O_1848,N_49661,N_48406);
nor UO_1849 (O_1849,N_47001,N_48157);
nor UO_1850 (O_1850,N_47253,N_49136);
nor UO_1851 (O_1851,N_49819,N_48815);
nor UO_1852 (O_1852,N_48206,N_48295);
nand UO_1853 (O_1853,N_45745,N_49693);
nor UO_1854 (O_1854,N_47892,N_47816);
nor UO_1855 (O_1855,N_47636,N_47030);
nor UO_1856 (O_1856,N_48916,N_45551);
and UO_1857 (O_1857,N_47317,N_45901);
nor UO_1858 (O_1858,N_45906,N_49417);
nand UO_1859 (O_1859,N_49949,N_46035);
xor UO_1860 (O_1860,N_47178,N_47371);
nor UO_1861 (O_1861,N_49065,N_47093);
xnor UO_1862 (O_1862,N_47078,N_47449);
nand UO_1863 (O_1863,N_48034,N_49180);
and UO_1864 (O_1864,N_47693,N_49879);
xor UO_1865 (O_1865,N_46414,N_48745);
xor UO_1866 (O_1866,N_48126,N_49038);
and UO_1867 (O_1867,N_47819,N_45640);
nor UO_1868 (O_1868,N_47605,N_46988);
or UO_1869 (O_1869,N_48762,N_48229);
and UO_1870 (O_1870,N_47326,N_45594);
nand UO_1871 (O_1871,N_49778,N_49317);
xor UO_1872 (O_1872,N_49684,N_49389);
or UO_1873 (O_1873,N_47040,N_46508);
and UO_1874 (O_1874,N_47867,N_48592);
and UO_1875 (O_1875,N_47021,N_45097);
or UO_1876 (O_1876,N_48185,N_49838);
or UO_1877 (O_1877,N_48333,N_45070);
xnor UO_1878 (O_1878,N_45560,N_48123);
nor UO_1879 (O_1879,N_47038,N_49615);
nor UO_1880 (O_1880,N_48475,N_47665);
and UO_1881 (O_1881,N_45341,N_48007);
xnor UO_1882 (O_1882,N_47199,N_47460);
and UO_1883 (O_1883,N_48913,N_46327);
nand UO_1884 (O_1884,N_46372,N_48110);
and UO_1885 (O_1885,N_49183,N_49002);
or UO_1886 (O_1886,N_47000,N_47988);
and UO_1887 (O_1887,N_45184,N_45633);
xnor UO_1888 (O_1888,N_47034,N_45306);
nand UO_1889 (O_1889,N_46685,N_47410);
and UO_1890 (O_1890,N_48197,N_49353);
nor UO_1891 (O_1891,N_48832,N_47526);
xnor UO_1892 (O_1892,N_47722,N_48109);
xor UO_1893 (O_1893,N_45567,N_47977);
nor UO_1894 (O_1894,N_49121,N_48594);
nor UO_1895 (O_1895,N_48136,N_48728);
or UO_1896 (O_1896,N_46082,N_46695);
nor UO_1897 (O_1897,N_47451,N_48972);
or UO_1898 (O_1898,N_46991,N_49610);
nor UO_1899 (O_1899,N_46957,N_47287);
or UO_1900 (O_1900,N_45897,N_48767);
nor UO_1901 (O_1901,N_47086,N_48607);
or UO_1902 (O_1902,N_45042,N_45730);
or UO_1903 (O_1903,N_46223,N_46885);
xnor UO_1904 (O_1904,N_49903,N_48991);
nor UO_1905 (O_1905,N_49114,N_47501);
and UO_1906 (O_1906,N_47147,N_47848);
nor UO_1907 (O_1907,N_48173,N_47146);
xnor UO_1908 (O_1908,N_46629,N_49146);
nor UO_1909 (O_1909,N_47729,N_47844);
nand UO_1910 (O_1910,N_45647,N_46567);
xnor UO_1911 (O_1911,N_49738,N_45605);
xnor UO_1912 (O_1912,N_48115,N_46348);
nor UO_1913 (O_1913,N_47006,N_48742);
or UO_1914 (O_1914,N_45150,N_48062);
or UO_1915 (O_1915,N_49173,N_48790);
xnor UO_1916 (O_1916,N_46653,N_49479);
nand UO_1917 (O_1917,N_46726,N_47627);
and UO_1918 (O_1918,N_49621,N_47663);
nor UO_1919 (O_1919,N_49712,N_48119);
or UO_1920 (O_1920,N_47847,N_48734);
xnor UO_1921 (O_1921,N_49700,N_45889);
xnor UO_1922 (O_1922,N_47522,N_45741);
nand UO_1923 (O_1923,N_49818,N_47602);
nand UO_1924 (O_1924,N_46553,N_48322);
or UO_1925 (O_1925,N_48747,N_46419);
and UO_1926 (O_1926,N_46919,N_45338);
and UO_1927 (O_1927,N_46502,N_48155);
xor UO_1928 (O_1928,N_48999,N_47708);
and UO_1929 (O_1929,N_46802,N_46687);
xnor UO_1930 (O_1930,N_48956,N_49887);
or UO_1931 (O_1931,N_46711,N_48667);
and UO_1932 (O_1932,N_48758,N_48596);
xnor UO_1933 (O_1933,N_49562,N_48647);
and UO_1934 (O_1934,N_47194,N_45458);
and UO_1935 (O_1935,N_47747,N_49645);
or UO_1936 (O_1936,N_49316,N_49839);
nor UO_1937 (O_1937,N_45397,N_45409);
nor UO_1938 (O_1938,N_48277,N_45944);
xor UO_1939 (O_1939,N_48890,N_49369);
xnor UO_1940 (O_1940,N_49902,N_48471);
xnor UO_1941 (O_1941,N_47456,N_49003);
and UO_1942 (O_1942,N_48190,N_45264);
nor UO_1943 (O_1943,N_48361,N_47004);
or UO_1944 (O_1944,N_49710,N_46914);
nor UO_1945 (O_1945,N_49658,N_46835);
nor UO_1946 (O_1946,N_45979,N_46512);
nand UO_1947 (O_1947,N_47737,N_46725);
nand UO_1948 (O_1948,N_48296,N_49739);
nand UO_1949 (O_1949,N_49552,N_48743);
and UO_1950 (O_1950,N_46248,N_45392);
and UO_1951 (O_1951,N_46677,N_48486);
nand UO_1952 (O_1952,N_46672,N_46265);
xnor UO_1953 (O_1953,N_48979,N_45711);
nor UO_1954 (O_1954,N_47869,N_45681);
nand UO_1955 (O_1955,N_47294,N_45555);
and UO_1956 (O_1956,N_45387,N_49933);
or UO_1957 (O_1957,N_45019,N_48558);
or UO_1958 (O_1958,N_47468,N_48175);
nand UO_1959 (O_1959,N_45291,N_47375);
nand UO_1960 (O_1960,N_47206,N_48589);
xnor UO_1961 (O_1961,N_46763,N_45632);
nor UO_1962 (O_1962,N_49579,N_46399);
nor UO_1963 (O_1963,N_45520,N_49045);
nand UO_1964 (O_1964,N_45121,N_47230);
xnor UO_1965 (O_1965,N_49628,N_49573);
and UO_1966 (O_1966,N_48925,N_45566);
xnor UO_1967 (O_1967,N_47577,N_47263);
and UO_1968 (O_1968,N_46718,N_49422);
xor UO_1969 (O_1969,N_47684,N_46600);
and UO_1970 (O_1970,N_47668,N_46005);
or UO_1971 (O_1971,N_46901,N_46533);
xor UO_1972 (O_1972,N_45351,N_48881);
xnor UO_1973 (O_1973,N_48196,N_46198);
and UO_1974 (O_1974,N_47758,N_47486);
nor UO_1975 (O_1975,N_45303,N_49572);
nor UO_1976 (O_1976,N_47377,N_49544);
or UO_1977 (O_1977,N_45394,N_47664);
xor UO_1978 (O_1978,N_49179,N_49626);
nor UO_1979 (O_1979,N_47814,N_47085);
nor UO_1980 (O_1980,N_47264,N_47169);
nor UO_1981 (O_1981,N_48355,N_45349);
or UO_1982 (O_1982,N_49541,N_46225);
or UO_1983 (O_1983,N_47182,N_45381);
xnor UO_1984 (O_1984,N_46818,N_46155);
and UO_1985 (O_1985,N_49113,N_49310);
or UO_1986 (O_1986,N_47639,N_49446);
and UO_1987 (O_1987,N_48116,N_46240);
and UO_1988 (O_1988,N_48281,N_49453);
nor UO_1989 (O_1989,N_45760,N_45960);
or UO_1990 (O_1990,N_46515,N_45266);
and UO_1991 (O_1991,N_46134,N_46926);
or UO_1992 (O_1992,N_46826,N_49374);
and UO_1993 (O_1993,N_45638,N_48369);
and UO_1994 (O_1994,N_46852,N_47027);
nand UO_1995 (O_1995,N_45755,N_49247);
nor UO_1996 (O_1996,N_45784,N_46698);
or UO_1997 (O_1997,N_47586,N_48032);
nor UO_1998 (O_1998,N_46204,N_49219);
and UO_1999 (O_1999,N_45163,N_45347);
xnor UO_2000 (O_2000,N_49764,N_48957);
and UO_2001 (O_2001,N_47696,N_47487);
and UO_2002 (O_2002,N_45835,N_49917);
nor UO_2003 (O_2003,N_46585,N_48100);
nor UO_2004 (O_2004,N_48848,N_49999);
xnor UO_2005 (O_2005,N_47968,N_47135);
and UO_2006 (O_2006,N_45440,N_45781);
nor UO_2007 (O_2007,N_47759,N_48937);
xor UO_2008 (O_2008,N_47986,N_48203);
and UO_2009 (O_2009,N_49653,N_47940);
nand UO_2010 (O_2010,N_48177,N_46094);
nor UO_2011 (O_2011,N_47757,N_48423);
nand UO_2012 (O_2012,N_49467,N_47444);
and UO_2013 (O_2013,N_45553,N_49596);
and UO_2014 (O_2014,N_48474,N_46741);
xnor UO_2015 (O_2015,N_45257,N_47831);
xor UO_2016 (O_2016,N_49517,N_48394);
and UO_2017 (O_2017,N_46696,N_45576);
or UO_2018 (O_2018,N_48236,N_49696);
xor UO_2019 (O_2019,N_45313,N_46180);
nand UO_2020 (O_2020,N_48039,N_48971);
or UO_2021 (O_2021,N_48686,N_48919);
or UO_2022 (O_2022,N_45637,N_47536);
and UO_2023 (O_2023,N_45713,N_48618);
nor UO_2024 (O_2024,N_49526,N_48460);
nand UO_2025 (O_2025,N_47037,N_45593);
xor UO_2026 (O_2026,N_45533,N_47667);
and UO_2027 (O_2027,N_46381,N_48288);
nand UO_2028 (O_2028,N_47480,N_47984);
or UO_2029 (O_2029,N_46572,N_46825);
or UO_2030 (O_2030,N_46931,N_46212);
and UO_2031 (O_2031,N_47303,N_45670);
and UO_2032 (O_2032,N_45154,N_46243);
and UO_2033 (O_2033,N_48609,N_47794);
nor UO_2034 (O_2034,N_48726,N_47017);
nor UO_2035 (O_2035,N_49291,N_49577);
nand UO_2036 (O_2036,N_48430,N_48040);
and UO_2037 (O_2037,N_49587,N_46635);
nor UO_2038 (O_2038,N_49748,N_46087);
or UO_2039 (O_2039,N_48201,N_47168);
xnor UO_2040 (O_2040,N_45541,N_47934);
xnor UO_2041 (O_2041,N_45535,N_46511);
and UO_2042 (O_2042,N_46293,N_48204);
xnor UO_2043 (O_2043,N_48346,N_46037);
nand UO_2044 (O_2044,N_45116,N_45769);
or UO_2045 (O_2045,N_46588,N_46640);
nand UO_2046 (O_2046,N_48800,N_46269);
or UO_2047 (O_2047,N_49418,N_49235);
nor UO_2048 (O_2048,N_49314,N_49627);
and UO_2049 (O_2049,N_48856,N_47509);
or UO_2050 (O_2050,N_46806,N_49018);
nor UO_2051 (O_2051,N_47870,N_47070);
or UO_2052 (O_2052,N_49010,N_47666);
xnor UO_2053 (O_2053,N_46755,N_46608);
nor UO_2054 (O_2054,N_46891,N_45877);
nand UO_2055 (O_2055,N_47571,N_46778);
xnor UO_2056 (O_2056,N_49468,N_46309);
or UO_2057 (O_2057,N_49370,N_47260);
xnor UO_2058 (O_2058,N_49482,N_48776);
nor UO_2059 (O_2059,N_47481,N_45283);
and UO_2060 (O_2060,N_46900,N_48396);
and UO_2061 (O_2061,N_46316,N_49561);
or UO_2062 (O_2062,N_45087,N_45214);
nor UO_2063 (O_2063,N_45546,N_49161);
and UO_2064 (O_2064,N_49205,N_48660);
xnor UO_2065 (O_2065,N_49448,N_46207);
or UO_2066 (O_2066,N_47730,N_46024);
nor UO_2067 (O_2067,N_49321,N_47948);
nand UO_2068 (O_2068,N_49308,N_47937);
or UO_2069 (O_2069,N_45488,N_46385);
or UO_2070 (O_2070,N_45509,N_47251);
nor UO_2071 (O_2071,N_45545,N_48122);
xor UO_2072 (O_2072,N_49861,N_47514);
nor UO_2073 (O_2073,N_48649,N_46117);
or UO_2074 (O_2074,N_45384,N_46139);
xor UO_2075 (O_2075,N_47504,N_47492);
xor UO_2076 (O_2076,N_48868,N_49972);
and UO_2077 (O_2077,N_48555,N_47917);
and UO_2078 (O_2078,N_47076,N_46397);
nor UO_2079 (O_2079,N_45072,N_46995);
nand UO_2080 (O_2080,N_46922,N_45106);
xnor UO_2081 (O_2081,N_46634,N_46435);
and UO_2082 (O_2082,N_48194,N_49213);
nor UO_2083 (O_2083,N_48802,N_46439);
nand UO_2084 (O_2084,N_49239,N_45528);
nor UO_2085 (O_2085,N_49455,N_45678);
xnor UO_2086 (O_2086,N_47024,N_48041);
and UO_2087 (O_2087,N_45176,N_46326);
nand UO_2088 (O_2088,N_49320,N_45864);
nand UO_2089 (O_2089,N_45471,N_48293);
or UO_2090 (O_2090,N_46317,N_47788);
and UO_2091 (O_2091,N_49260,N_45855);
nand UO_2092 (O_2092,N_47975,N_48590);
nand UO_2093 (O_2093,N_49636,N_48113);
and UO_2094 (O_2094,N_47390,N_49457);
or UO_2095 (O_2095,N_47597,N_49397);
or UO_2096 (O_2096,N_46416,N_46928);
nor UO_2097 (O_2097,N_46216,N_48479);
and UO_2098 (O_2098,N_48633,N_49450);
and UO_2099 (O_2099,N_46430,N_45065);
or UO_2100 (O_2100,N_48616,N_47335);
xnor UO_2101 (O_2101,N_46609,N_49907);
nor UO_2102 (O_2102,N_46319,N_49637);
and UO_2103 (O_2103,N_45128,N_47766);
xor UO_2104 (O_2104,N_45782,N_49893);
nor UO_2105 (O_2105,N_48076,N_46078);
and UO_2106 (O_2106,N_47952,N_47238);
and UO_2107 (O_2107,N_47728,N_45400);
and UO_2108 (O_2108,N_46651,N_47785);
and UO_2109 (O_2109,N_45840,N_49262);
or UO_2110 (O_2110,N_48061,N_46275);
nand UO_2111 (O_2111,N_45631,N_47810);
and UO_2112 (O_2112,N_45356,N_45827);
nand UO_2113 (O_2113,N_49295,N_49126);
or UO_2114 (O_2114,N_47276,N_47469);
nor UO_2115 (O_2115,N_48405,N_47052);
or UO_2116 (O_2116,N_49783,N_48676);
nand UO_2117 (O_2117,N_45100,N_47703);
xor UO_2118 (O_2118,N_45470,N_46175);
nand UO_2119 (O_2119,N_49351,N_45544);
xnor UO_2120 (O_2120,N_45177,N_46323);
nand UO_2121 (O_2121,N_47507,N_46387);
xnor UO_2122 (O_2122,N_48872,N_46031);
or UO_2123 (O_2123,N_49139,N_48436);
nand UO_2124 (O_2124,N_45370,N_48093);
nand UO_2125 (O_2125,N_47095,N_46369);
xnor UO_2126 (O_2126,N_46921,N_47195);
and UO_2127 (O_2127,N_45887,N_47744);
nand UO_2128 (O_2128,N_48624,N_47506);
and UO_2129 (O_2129,N_48672,N_48951);
and UO_2130 (O_2130,N_47105,N_49040);
nor UO_2131 (O_2131,N_46719,N_49234);
nand UO_2132 (O_2132,N_45149,N_47584);
and UO_2133 (O_2133,N_45425,N_47673);
and UO_2134 (O_2134,N_47902,N_46245);
nand UO_2135 (O_2135,N_49130,N_45430);
nand UO_2136 (O_2136,N_45290,N_45552);
nand UO_2137 (O_2137,N_45331,N_49864);
and UO_2138 (O_2138,N_45018,N_46152);
xnor UO_2139 (O_2139,N_48227,N_46407);
nor UO_2140 (O_2140,N_46872,N_49695);
nor UO_2141 (O_2141,N_49071,N_47208);
nor UO_2142 (O_2142,N_45365,N_46311);
nand UO_2143 (O_2143,N_49334,N_45320);
nand UO_2144 (O_2144,N_45164,N_45114);
or UO_2145 (O_2145,N_45947,N_48529);
nand UO_2146 (O_2146,N_48764,N_49284);
nor UO_2147 (O_2147,N_48245,N_49614);
nand UO_2148 (O_2148,N_45911,N_46174);
and UO_2149 (O_2149,N_49915,N_48582);
and UO_2150 (O_2150,N_47406,N_49033);
xor UO_2151 (O_2151,N_49042,N_48166);
and UO_2152 (O_2152,N_46053,N_48417);
xor UO_2153 (O_2153,N_48380,N_48651);
and UO_2154 (O_2154,N_47367,N_45233);
xnor UO_2155 (O_2155,N_49258,N_49193);
nor UO_2156 (O_2156,N_49594,N_46548);
or UO_2157 (O_2157,N_46121,N_45393);
xor UO_2158 (O_2158,N_45412,N_48438);
nand UO_2159 (O_2159,N_48823,N_45377);
xor UO_2160 (O_2160,N_45814,N_45218);
xor UO_2161 (O_2161,N_45005,N_48701);
and UO_2162 (O_2162,N_47055,N_46809);
nand UO_2163 (O_2163,N_49943,N_49806);
or UO_2164 (O_2164,N_47014,N_49954);
nand UO_2165 (O_2165,N_49753,N_48793);
nor UO_2166 (O_2166,N_48556,N_45615);
or UO_2167 (O_2167,N_48860,N_48502);
or UO_2168 (O_2168,N_47637,N_46530);
nor UO_2169 (O_2169,N_46353,N_48684);
nor UO_2170 (O_2170,N_47474,N_49771);
and UO_2171 (O_2171,N_47304,N_47518);
nand UO_2172 (O_2172,N_47227,N_47427);
nand UO_2173 (O_2173,N_46195,N_46098);
and UO_2174 (O_2174,N_48178,N_47680);
nor UO_2175 (O_2175,N_45224,N_46752);
xor UO_2176 (O_2176,N_46980,N_45011);
or UO_2177 (O_2177,N_46313,N_47071);
nand UO_2178 (O_2178,N_48050,N_49742);
or UO_2179 (O_2179,N_45738,N_49031);
xor UO_2180 (O_2180,N_45607,N_46202);
nor UO_2181 (O_2181,N_45407,N_49988);
or UO_2182 (O_2182,N_49390,N_46797);
xnor UO_2183 (O_2183,N_45285,N_49209);
xor UO_2184 (O_2184,N_48524,N_47546);
or UO_2185 (O_2185,N_46626,N_48581);
nor UO_2186 (O_2186,N_49458,N_49757);
or UO_2187 (O_2187,N_49400,N_46272);
nor UO_2188 (O_2188,N_45007,N_49132);
xor UO_2189 (O_2189,N_49547,N_45332);
nand UO_2190 (O_2190,N_45035,N_47983);
nand UO_2191 (O_2191,N_49428,N_49140);
nand UO_2192 (O_2192,N_49011,N_47717);
nor UO_2193 (O_2193,N_45136,N_45232);
and UO_2194 (O_2194,N_49834,N_46120);
nor UO_2195 (O_2195,N_46952,N_48824);
and UO_2196 (O_2196,N_47023,N_46641);
xor UO_2197 (O_2197,N_47382,N_49097);
or UO_2198 (O_2198,N_46284,N_48809);
or UO_2199 (O_2199,N_46678,N_47437);
nor UO_2200 (O_2200,N_49884,N_48772);
nand UO_2201 (O_2201,N_47980,N_46897);
or UO_2202 (O_2202,N_48381,N_48171);
nor UO_2203 (O_2203,N_49531,N_48698);
or UO_2204 (O_2204,N_48118,N_48785);
and UO_2205 (O_2205,N_49300,N_45202);
nor UO_2206 (O_2206,N_47513,N_47058);
or UO_2207 (O_2207,N_46992,N_46102);
nor UO_2208 (O_2208,N_49358,N_45731);
nand UO_2209 (O_2209,N_45601,N_47415);
and UO_2210 (O_2210,N_48156,N_47331);
xor UO_2211 (O_2211,N_49646,N_49871);
and UO_2212 (O_2212,N_49191,N_49537);
or UO_2213 (O_2213,N_46622,N_47687);
nor UO_2214 (O_2214,N_47079,N_45211);
or UO_2215 (O_2215,N_46166,N_45578);
or UO_2216 (O_2216,N_48102,N_46189);
nor UO_2217 (O_2217,N_45130,N_49630);
nand UO_2218 (O_2218,N_47962,N_46680);
nand UO_2219 (O_2219,N_49721,N_49231);
xnor UO_2220 (O_2220,N_49159,N_48221);
nor UO_2221 (O_2221,N_46305,N_48289);
and UO_2222 (O_2222,N_48569,N_47564);
or UO_2223 (O_2223,N_48441,N_48287);
and UO_2224 (O_2224,N_46550,N_49557);
xor UO_2225 (O_2225,N_49379,N_47122);
nor UO_2226 (O_2226,N_47277,N_49439);
or UO_2227 (O_2227,N_47656,N_47101);
nand UO_2228 (O_2228,N_45981,N_48936);
or UO_2229 (O_2229,N_48121,N_47019);
and UO_2230 (O_2230,N_49730,N_49425);
nand UO_2231 (O_2231,N_46380,N_48454);
or UO_2232 (O_2232,N_49522,N_47822);
nand UO_2233 (O_2233,N_47723,N_46814);
nand UO_2234 (O_2234,N_48499,N_47380);
or UO_2235 (O_2235,N_48828,N_47413);
nor UO_2236 (O_2236,N_49652,N_49575);
xnor UO_2237 (O_2237,N_49340,N_49052);
nand UO_2238 (O_2238,N_45831,N_45326);
nor UO_2239 (O_2239,N_45529,N_49196);
nor UO_2240 (O_2240,N_45896,N_47318);
or UO_2241 (O_2241,N_46674,N_48735);
nor UO_2242 (O_2242,N_45252,N_49530);
and UO_2243 (O_2243,N_46938,N_47368);
nor UO_2244 (O_2244,N_45859,N_45957);
nor UO_2245 (O_2245,N_48127,N_47476);
or UO_2246 (O_2246,N_45134,N_45807);
or UO_2247 (O_2247,N_45819,N_46422);
and UO_2248 (O_2248,N_48146,N_49135);
and UO_2249 (O_2249,N_49910,N_49595);
and UO_2250 (O_2250,N_48225,N_47701);
nor UO_2251 (O_2251,N_47219,N_48855);
nor UO_2252 (O_2252,N_48013,N_45220);
or UO_2253 (O_2253,N_45608,N_45592);
and UO_2254 (O_2254,N_45462,N_46036);
nand UO_2255 (O_2255,N_45411,N_45161);
xor UO_2256 (O_2256,N_49992,N_46887);
and UO_2257 (O_2257,N_46081,N_49257);
nor UO_2258 (O_2258,N_49583,N_46213);
or UO_2259 (O_2259,N_48461,N_48169);
or UO_2260 (O_2260,N_45196,N_46429);
nand UO_2261 (O_2261,N_48969,N_47622);
nor UO_2262 (O_2262,N_49001,N_45204);
and UO_2263 (O_2263,N_45122,N_48292);
or UO_2264 (O_2264,N_48945,N_45967);
or UO_2265 (O_2265,N_46306,N_46569);
xnor UO_2266 (O_2266,N_47718,N_46787);
xnor UO_2267 (O_2267,N_45962,N_49975);
nand UO_2268 (O_2268,N_46871,N_47749);
nand UO_2269 (O_2269,N_47466,N_49264);
nor UO_2270 (O_2270,N_49790,N_45197);
xnor UO_2271 (O_2271,N_47321,N_47533);
and UO_2272 (O_2272,N_48977,N_48326);
nand UO_2273 (O_2273,N_49361,N_46325);
nor UO_2274 (O_2274,N_49584,N_49037);
nand UO_2275 (O_2275,N_45820,N_49017);
xor UO_2276 (O_2276,N_48929,N_48998);
nor UO_2277 (O_2277,N_49793,N_46807);
nand UO_2278 (O_2278,N_49411,N_47061);
xnor UO_2279 (O_2279,N_49633,N_49443);
xnor UO_2280 (O_2280,N_48902,N_48564);
or UO_2281 (O_2281,N_47771,N_45127);
xnor UO_2282 (O_2282,N_46329,N_46057);
and UO_2283 (O_2283,N_49212,N_45081);
or UO_2284 (O_2284,N_48005,N_46217);
nor UO_2285 (O_2285,N_46250,N_49182);
or UO_2286 (O_2286,N_49220,N_47800);
nand UO_2287 (O_2287,N_49476,N_49534);
nand UO_2288 (O_2288,N_46779,N_47077);
nand UO_2289 (O_2289,N_45478,N_49421);
and UO_2290 (O_2290,N_47698,N_45335);
and UO_2291 (O_2291,N_47423,N_47255);
nor UO_2292 (O_2292,N_47858,N_47862);
xnor UO_2293 (O_2293,N_46717,N_47652);
or UO_2294 (O_2294,N_47881,N_48241);
xnor UO_2295 (O_2295,N_49539,N_47965);
xor UO_2296 (O_2296,N_45721,N_46129);
nand UO_2297 (O_2297,N_45761,N_48071);
nor UO_2298 (O_2298,N_47351,N_48080);
nor UO_2299 (O_2299,N_47713,N_46238);
or UO_2300 (O_2300,N_49415,N_48010);
and UO_2301 (O_2301,N_46834,N_46345);
and UO_2302 (O_2302,N_46942,N_49554);
nand UO_2303 (O_2303,N_46638,N_47166);
nor UO_2304 (O_2304,N_46748,N_45753);
or UO_2305 (O_2305,N_49241,N_46106);
or UO_2306 (O_2306,N_47066,N_49060);
and UO_2307 (O_2307,N_46025,N_48525);
and UO_2308 (O_2308,N_48272,N_49609);
nor UO_2309 (O_2309,N_45408,N_47275);
xor UO_2310 (O_2310,N_46560,N_49593);
or UO_2311 (O_2311,N_47295,N_46886);
and UO_2312 (O_2312,N_48195,N_46247);
or UO_2313 (O_2313,N_46709,N_48789);
xor UO_2314 (O_2314,N_48491,N_46747);
nor UO_2315 (O_2315,N_45583,N_46693);
nand UO_2316 (O_2316,N_49647,N_49500);
nand UO_2317 (O_2317,N_48964,N_49073);
xor UO_2318 (O_2318,N_47445,N_46222);
or UO_2319 (O_2319,N_45951,N_45022);
xnor UO_2320 (O_2320,N_46819,N_48297);
nor UO_2321 (O_2321,N_47846,N_48650);
and UO_2322 (O_2322,N_47695,N_46049);
or UO_2323 (O_2323,N_49733,N_49392);
nor UO_2324 (O_2324,N_46052,N_49923);
nor UO_2325 (O_2325,N_48599,N_47795);
and UO_2326 (O_2326,N_45491,N_47300);
nor UO_2327 (O_2327,N_46378,N_46188);
and UO_2328 (O_2328,N_48621,N_46171);
and UO_2329 (O_2329,N_48965,N_47823);
xor UO_2330 (O_2330,N_46916,N_47719);
xnor UO_2331 (O_2331,N_45502,N_47397);
xor UO_2332 (O_2332,N_47216,N_46531);
nand UO_2333 (O_2333,N_48011,N_49285);
or UO_2334 (O_2334,N_49914,N_46538);
nand UO_2335 (O_2335,N_49916,N_45614);
or UO_2336 (O_2336,N_45308,N_45561);
xnor UO_2337 (O_2337,N_45382,N_46801);
or UO_2338 (O_2338,N_47108,N_47394);
nor UO_2339 (O_2339,N_49292,N_46114);
nor UO_2340 (O_2340,N_45702,N_46652);
xnor UO_2341 (O_2341,N_47026,N_46091);
xor UO_2342 (O_2342,N_47595,N_48275);
and UO_2343 (O_2343,N_47517,N_48927);
nor UO_2344 (O_2344,N_45881,N_45589);
and UO_2345 (O_2345,N_49582,N_47907);
and UO_2346 (O_2346,N_48920,N_49540);
or UO_2347 (O_2347,N_48984,N_49435);
nor UO_2348 (O_2348,N_46490,N_46820);
and UO_2349 (O_2349,N_46744,N_49817);
nor UO_2350 (O_2350,N_47686,N_47997);
xor UO_2351 (O_2351,N_47274,N_49641);
or UO_2352 (O_2352,N_48545,N_46268);
and UO_2353 (O_2353,N_46786,N_45179);
nand UO_2354 (O_2354,N_49772,N_48511);
and UO_2355 (O_2355,N_45046,N_47710);
nand UO_2356 (O_2356,N_48859,N_45466);
nor UO_2357 (O_2357,N_47201,N_48413);
nor UO_2358 (O_2358,N_47478,N_46913);
or UO_2359 (O_2359,N_48217,N_48814);
and UO_2360 (O_2360,N_49974,N_48612);
or UO_2361 (O_2361,N_49497,N_47044);
or UO_2362 (O_2362,N_47538,N_47210);
and UO_2363 (O_2363,N_48248,N_46911);
or UO_2364 (O_2364,N_49006,N_45779);
or UO_2365 (O_2365,N_46964,N_48550);
nor UO_2366 (O_2366,N_49099,N_46522);
or UO_2367 (O_2367,N_45636,N_48057);
nand UO_2368 (O_2368,N_49278,N_49624);
nor UO_2369 (O_2369,N_49233,N_47407);
nor UO_2370 (O_2370,N_47453,N_46917);
xor UO_2371 (O_2371,N_47315,N_46296);
nor UO_2372 (O_2372,N_46441,N_49309);
or UO_2373 (O_2373,N_45391,N_48877);
xor UO_2374 (O_2374,N_47855,N_47801);
or UO_2375 (O_2375,N_46146,N_45505);
nand UO_2376 (O_2376,N_45207,N_47891);
nand UO_2377 (O_2377,N_47820,N_49958);
nand UO_2378 (O_2378,N_46410,N_48490);
or UO_2379 (O_2379,N_47612,N_45833);
nor UO_2380 (O_2380,N_47191,N_47204);
and UO_2381 (O_2381,N_48673,N_48656);
nor UO_2382 (O_2382,N_47811,N_45234);
nand UO_2383 (O_2383,N_45198,N_47031);
or UO_2384 (O_2384,N_46357,N_45718);
or UO_2385 (O_2385,N_45422,N_47435);
xnor UO_2386 (O_2386,N_49454,N_45386);
nor UO_2387 (O_2387,N_49110,N_46320);
nand UO_2388 (O_2388,N_49946,N_46489);
xnor UO_2389 (O_2389,N_46927,N_47067);
or UO_2390 (O_2390,N_45972,N_45716);
and UO_2391 (O_2391,N_48725,N_45800);
and UO_2392 (O_2392,N_46168,N_47214);
xnor UO_2393 (O_2393,N_48806,N_48819);
and UO_2394 (O_2394,N_48985,N_47761);
nand UO_2395 (O_2395,N_46723,N_49020);
or UO_2396 (O_2396,N_46941,N_45524);
xor UO_2397 (O_2397,N_49395,N_48716);
nor UO_2398 (O_2398,N_46597,N_45842);
nand UO_2399 (O_2399,N_45416,N_45076);
or UO_2400 (O_2400,N_49720,N_46720);
and UO_2401 (O_2401,N_47222,N_47176);
nand UO_2402 (O_2402,N_49816,N_45843);
nor UO_2403 (O_2403,N_46990,N_46734);
nand UO_2404 (O_2404,N_45027,N_49124);
and UO_2405 (O_2405,N_45977,N_49156);
xor UO_2406 (O_2406,N_45036,N_47248);
nand UO_2407 (O_2407,N_48719,N_48513);
nor UO_2408 (O_2408,N_48657,N_48708);
nor UO_2409 (O_2409,N_48323,N_46945);
and UO_2410 (O_2410,N_46333,N_45475);
or UO_2411 (O_2411,N_49105,N_47957);
and UO_2412 (O_2412,N_47777,N_48462);
or UO_2413 (O_2413,N_49112,N_46971);
and UO_2414 (O_2414,N_48352,N_46743);
nor UO_2415 (O_2415,N_46751,N_47102);
xor UO_2416 (O_2416,N_45651,N_45095);
and UO_2417 (O_2417,N_47418,N_47162);
or UO_2418 (O_2418,N_47895,N_47307);
or UO_2419 (O_2419,N_47003,N_49924);
nand UO_2420 (O_2420,N_45863,N_45969);
nand UO_2421 (O_2421,N_46853,N_47829);
nand UO_2422 (O_2422,N_45371,N_46824);
and UO_2423 (O_2423,N_46029,N_49372);
nor UO_2424 (O_2424,N_46736,N_46521);
nor UO_2425 (O_2425,N_49631,N_47281);
or UO_2426 (O_2426,N_49980,N_49922);
and UO_2427 (O_2427,N_45304,N_45975);
and UO_2428 (O_2428,N_45139,N_45028);
or UO_2429 (O_2429,N_46228,N_45033);
nand UO_2430 (O_2430,N_49768,N_49527);
and UO_2431 (O_2431,N_49357,N_49672);
and UO_2432 (O_2432,N_45919,N_45259);
or UO_2433 (O_2433,N_45764,N_46555);
and UO_2434 (O_2434,N_46589,N_45213);
xor UO_2435 (O_2435,N_48137,N_48151);
and UO_2436 (O_2436,N_48006,N_45016);
nand UO_2437 (O_2437,N_46287,N_46395);
nand UO_2438 (O_2438,N_48791,N_48693);
xnor UO_2439 (O_2439,N_49238,N_48251);
and UO_2440 (O_2440,N_49896,N_47897);
nor UO_2441 (O_2441,N_46691,N_47328);
and UO_2442 (O_2442,N_45930,N_49157);
and UO_2443 (O_2443,N_45236,N_47745);
or UO_2444 (O_2444,N_48658,N_48857);
or UO_2445 (O_2445,N_47865,N_47104);
nand UO_2446 (O_2446,N_47799,N_45348);
nand UO_2447 (O_2447,N_49565,N_49632);
nand UO_2448 (O_2448,N_49929,N_45674);
xnor UO_2449 (O_2449,N_45942,N_46733);
nor UO_2450 (O_2450,N_47755,N_48690);
or UO_2451 (O_2451,N_49791,N_47389);
or UO_2452 (O_2452,N_49359,N_48975);
or UO_2453 (O_2453,N_47922,N_46475);
or UO_2454 (O_2454,N_48008,N_49477);
xnor UO_2455 (O_2455,N_48749,N_45584);
nor UO_2456 (O_2456,N_47072,N_48244);
or UO_2457 (O_2457,N_46273,N_45312);
nand UO_2458 (O_2458,N_45360,N_47910);
or UO_2459 (O_2459,N_48168,N_47033);
or UO_2460 (O_2460,N_48962,N_49256);
nand UO_2461 (O_2461,N_47887,N_47523);
nand UO_2462 (O_2462,N_49004,N_48286);
or UO_2463 (O_2463,N_45986,N_46346);
nand UO_2464 (O_2464,N_49172,N_45910);
nor UO_2465 (O_2465,N_48106,N_47459);
or UO_2466 (O_2466,N_48141,N_46915);
nand UO_2467 (O_2467,N_49535,N_48677);
nor UO_2468 (O_2468,N_45489,N_46881);
or UO_2469 (O_2469,N_48842,N_49959);
or UO_2470 (O_2470,N_49588,N_48419);
or UO_2471 (O_2471,N_47921,N_48866);
or UO_2472 (O_2472,N_47257,N_48794);
or UO_2473 (O_2473,N_46722,N_49576);
xor UO_2474 (O_2474,N_47366,N_49208);
or UO_2475 (O_2475,N_45558,N_47045);
and UO_2476 (O_2476,N_47625,N_46096);
and UO_2477 (O_2477,N_46749,N_45477);
or UO_2478 (O_2478,N_47840,N_49363);
xnor UO_2479 (O_2479,N_47180,N_49845);
nor UO_2480 (O_2480,N_48313,N_48778);
and UO_2481 (O_2481,N_47798,N_47700);
and UO_2482 (O_2482,N_48408,N_48895);
nor UO_2483 (O_2483,N_46491,N_47682);
nand UO_2484 (O_2484,N_47863,N_45499);
or UO_2485 (O_2485,N_48852,N_48497);
xor UO_2486 (O_2486,N_45293,N_45249);
xnor UO_2487 (O_2487,N_49318,N_45504);
nor UO_2488 (O_2488,N_49460,N_47042);
xnor UO_2489 (O_2489,N_47220,N_49391);
and UO_2490 (O_2490,N_49982,N_47053);
nor UO_2491 (O_2491,N_48797,N_47649);
and UO_2492 (O_2492,N_49874,N_45531);
nor UO_2493 (O_2493,N_48712,N_46933);
and UO_2494 (O_2494,N_49865,N_49920);
nand UO_2495 (O_2495,N_47764,N_48804);
or UO_2496 (O_2496,N_48527,N_47409);
or UO_2497 (O_2497,N_48416,N_45120);
nor UO_2498 (O_2498,N_46411,N_45073);
xor UO_2499 (O_2499,N_49885,N_46408);
or UO_2500 (O_2500,N_46458,N_48353);
xor UO_2501 (O_2501,N_49019,N_48826);
and UO_2502 (O_2502,N_49817,N_45355);
nand UO_2503 (O_2503,N_49920,N_49074);
nor UO_2504 (O_2504,N_49146,N_48810);
nor UO_2505 (O_2505,N_47049,N_48530);
or UO_2506 (O_2506,N_48588,N_46173);
and UO_2507 (O_2507,N_49809,N_46068);
and UO_2508 (O_2508,N_47592,N_46173);
or UO_2509 (O_2509,N_47771,N_45914);
xnor UO_2510 (O_2510,N_48377,N_45511);
nand UO_2511 (O_2511,N_48462,N_45013);
and UO_2512 (O_2512,N_48664,N_48573);
nor UO_2513 (O_2513,N_49332,N_47792);
nor UO_2514 (O_2514,N_45139,N_49471);
nor UO_2515 (O_2515,N_48796,N_47409);
and UO_2516 (O_2516,N_47140,N_46042);
and UO_2517 (O_2517,N_45505,N_45605);
and UO_2518 (O_2518,N_49601,N_48627);
or UO_2519 (O_2519,N_49000,N_45341);
and UO_2520 (O_2520,N_48386,N_48049);
nor UO_2521 (O_2521,N_49841,N_46531);
or UO_2522 (O_2522,N_45807,N_47914);
or UO_2523 (O_2523,N_45269,N_48925);
and UO_2524 (O_2524,N_46984,N_45630);
and UO_2525 (O_2525,N_45837,N_46612);
and UO_2526 (O_2526,N_47065,N_45704);
or UO_2527 (O_2527,N_47029,N_49717);
and UO_2528 (O_2528,N_45493,N_46756);
nor UO_2529 (O_2529,N_45057,N_46026);
or UO_2530 (O_2530,N_46118,N_48423);
or UO_2531 (O_2531,N_47744,N_48856);
nor UO_2532 (O_2532,N_48804,N_45488);
nand UO_2533 (O_2533,N_46963,N_47316);
or UO_2534 (O_2534,N_46130,N_45716);
xor UO_2535 (O_2535,N_47462,N_47624);
xor UO_2536 (O_2536,N_46002,N_48402);
or UO_2537 (O_2537,N_46565,N_45538);
and UO_2538 (O_2538,N_45201,N_47254);
and UO_2539 (O_2539,N_47813,N_46556);
or UO_2540 (O_2540,N_47252,N_45955);
xnor UO_2541 (O_2541,N_45454,N_47736);
and UO_2542 (O_2542,N_45227,N_45332);
nor UO_2543 (O_2543,N_48758,N_48968);
or UO_2544 (O_2544,N_48436,N_49656);
and UO_2545 (O_2545,N_46687,N_45182);
nand UO_2546 (O_2546,N_48795,N_47272);
xor UO_2547 (O_2547,N_47310,N_46491);
or UO_2548 (O_2548,N_49618,N_46937);
nor UO_2549 (O_2549,N_49121,N_48140);
nand UO_2550 (O_2550,N_48447,N_48302);
nor UO_2551 (O_2551,N_46560,N_49461);
or UO_2552 (O_2552,N_49470,N_49688);
or UO_2553 (O_2553,N_48632,N_48443);
and UO_2554 (O_2554,N_45725,N_45340);
xnor UO_2555 (O_2555,N_46443,N_47529);
or UO_2556 (O_2556,N_45080,N_49336);
nor UO_2557 (O_2557,N_46643,N_47457);
nand UO_2558 (O_2558,N_49839,N_49816);
nor UO_2559 (O_2559,N_45935,N_46318);
xor UO_2560 (O_2560,N_45905,N_45838);
or UO_2561 (O_2561,N_46821,N_46464);
or UO_2562 (O_2562,N_45034,N_45942);
nand UO_2563 (O_2563,N_49013,N_45039);
nor UO_2564 (O_2564,N_46359,N_48214);
xnor UO_2565 (O_2565,N_48933,N_46897);
or UO_2566 (O_2566,N_48360,N_46111);
or UO_2567 (O_2567,N_45031,N_46965);
nor UO_2568 (O_2568,N_45130,N_48816);
nand UO_2569 (O_2569,N_49200,N_45487);
nand UO_2570 (O_2570,N_46763,N_45922);
or UO_2571 (O_2571,N_45222,N_48127);
nand UO_2572 (O_2572,N_48597,N_47789);
nand UO_2573 (O_2573,N_45461,N_45798);
xor UO_2574 (O_2574,N_48278,N_46624);
or UO_2575 (O_2575,N_47075,N_49836);
nor UO_2576 (O_2576,N_48631,N_48260);
xor UO_2577 (O_2577,N_49454,N_47107);
nand UO_2578 (O_2578,N_48181,N_46663);
or UO_2579 (O_2579,N_49042,N_48513);
and UO_2580 (O_2580,N_45582,N_45526);
and UO_2581 (O_2581,N_48456,N_47775);
nor UO_2582 (O_2582,N_46519,N_45824);
and UO_2583 (O_2583,N_47655,N_46090);
nand UO_2584 (O_2584,N_45596,N_49180);
xor UO_2585 (O_2585,N_47283,N_47296);
nor UO_2586 (O_2586,N_46638,N_49900);
xor UO_2587 (O_2587,N_47501,N_46872);
or UO_2588 (O_2588,N_49277,N_49788);
xnor UO_2589 (O_2589,N_47859,N_46980);
or UO_2590 (O_2590,N_47049,N_48692);
or UO_2591 (O_2591,N_47982,N_48988);
nor UO_2592 (O_2592,N_48526,N_46359);
xnor UO_2593 (O_2593,N_48634,N_47584);
xnor UO_2594 (O_2594,N_45164,N_49341);
and UO_2595 (O_2595,N_47215,N_47589);
and UO_2596 (O_2596,N_47407,N_48395);
nand UO_2597 (O_2597,N_45295,N_48600);
and UO_2598 (O_2598,N_46375,N_49759);
xor UO_2599 (O_2599,N_46519,N_46487);
or UO_2600 (O_2600,N_49063,N_47342);
nor UO_2601 (O_2601,N_45549,N_49173);
nor UO_2602 (O_2602,N_48631,N_49568);
nor UO_2603 (O_2603,N_45123,N_46803);
or UO_2604 (O_2604,N_46256,N_47764);
and UO_2605 (O_2605,N_48287,N_48280);
nor UO_2606 (O_2606,N_48329,N_45589);
nor UO_2607 (O_2607,N_48648,N_48896);
xnor UO_2608 (O_2608,N_45496,N_45414);
and UO_2609 (O_2609,N_46649,N_48441);
xor UO_2610 (O_2610,N_46801,N_45403);
xor UO_2611 (O_2611,N_47891,N_48035);
or UO_2612 (O_2612,N_47252,N_47638);
xor UO_2613 (O_2613,N_48526,N_49527);
or UO_2614 (O_2614,N_46358,N_48140);
nor UO_2615 (O_2615,N_49299,N_49865);
nand UO_2616 (O_2616,N_47007,N_49334);
or UO_2617 (O_2617,N_48549,N_45823);
nand UO_2618 (O_2618,N_45608,N_45956);
nor UO_2619 (O_2619,N_47680,N_47521);
xnor UO_2620 (O_2620,N_46110,N_45628);
xor UO_2621 (O_2621,N_47907,N_47733);
nand UO_2622 (O_2622,N_48974,N_47214);
and UO_2623 (O_2623,N_47812,N_45023);
xor UO_2624 (O_2624,N_49593,N_48403);
xnor UO_2625 (O_2625,N_49607,N_45630);
xnor UO_2626 (O_2626,N_49209,N_48309);
and UO_2627 (O_2627,N_46948,N_46021);
xnor UO_2628 (O_2628,N_48137,N_46290);
nand UO_2629 (O_2629,N_45789,N_45889);
xnor UO_2630 (O_2630,N_46252,N_45590);
nor UO_2631 (O_2631,N_46492,N_47823);
and UO_2632 (O_2632,N_45984,N_46181);
nor UO_2633 (O_2633,N_45341,N_48924);
or UO_2634 (O_2634,N_47874,N_48078);
nand UO_2635 (O_2635,N_45387,N_47493);
nor UO_2636 (O_2636,N_47668,N_46891);
nor UO_2637 (O_2637,N_48011,N_49324);
or UO_2638 (O_2638,N_49272,N_46220);
nor UO_2639 (O_2639,N_46965,N_47549);
nor UO_2640 (O_2640,N_48004,N_45257);
or UO_2641 (O_2641,N_49213,N_46630);
or UO_2642 (O_2642,N_45226,N_45989);
nand UO_2643 (O_2643,N_48885,N_49190);
xnor UO_2644 (O_2644,N_45176,N_46103);
or UO_2645 (O_2645,N_49551,N_48190);
xor UO_2646 (O_2646,N_45259,N_47104);
nand UO_2647 (O_2647,N_48411,N_47531);
nand UO_2648 (O_2648,N_45304,N_48763);
or UO_2649 (O_2649,N_48815,N_48735);
xnor UO_2650 (O_2650,N_47690,N_46559);
and UO_2651 (O_2651,N_45961,N_46127);
nand UO_2652 (O_2652,N_49659,N_46335);
and UO_2653 (O_2653,N_47124,N_46044);
nand UO_2654 (O_2654,N_45228,N_48977);
or UO_2655 (O_2655,N_48920,N_49353);
nor UO_2656 (O_2656,N_48636,N_47215);
nor UO_2657 (O_2657,N_47145,N_48822);
nand UO_2658 (O_2658,N_45051,N_47916);
and UO_2659 (O_2659,N_49963,N_49538);
or UO_2660 (O_2660,N_49061,N_49266);
xor UO_2661 (O_2661,N_49943,N_46742);
nor UO_2662 (O_2662,N_48549,N_47626);
xor UO_2663 (O_2663,N_49030,N_48410);
nand UO_2664 (O_2664,N_46605,N_48855);
xnor UO_2665 (O_2665,N_46398,N_46345);
nand UO_2666 (O_2666,N_46687,N_46466);
and UO_2667 (O_2667,N_46721,N_46848);
nor UO_2668 (O_2668,N_45166,N_45886);
nand UO_2669 (O_2669,N_45141,N_48522);
nor UO_2670 (O_2670,N_47759,N_47363);
or UO_2671 (O_2671,N_46996,N_46685);
nor UO_2672 (O_2672,N_48253,N_48827);
nor UO_2673 (O_2673,N_47946,N_46653);
nor UO_2674 (O_2674,N_47388,N_48982);
and UO_2675 (O_2675,N_45198,N_45735);
and UO_2676 (O_2676,N_48267,N_45939);
xor UO_2677 (O_2677,N_46204,N_47716);
nand UO_2678 (O_2678,N_47714,N_45602);
nor UO_2679 (O_2679,N_47880,N_48146);
and UO_2680 (O_2680,N_49810,N_46698);
and UO_2681 (O_2681,N_45906,N_45189);
nand UO_2682 (O_2682,N_47935,N_49618);
nor UO_2683 (O_2683,N_47115,N_48049);
and UO_2684 (O_2684,N_47077,N_48969);
or UO_2685 (O_2685,N_47756,N_46591);
xor UO_2686 (O_2686,N_47351,N_46356);
or UO_2687 (O_2687,N_45299,N_49178);
or UO_2688 (O_2688,N_47111,N_47728);
nor UO_2689 (O_2689,N_46458,N_48951);
and UO_2690 (O_2690,N_46865,N_48397);
and UO_2691 (O_2691,N_48191,N_46503);
xnor UO_2692 (O_2692,N_45146,N_47735);
or UO_2693 (O_2693,N_47881,N_48347);
nand UO_2694 (O_2694,N_45951,N_47544);
and UO_2695 (O_2695,N_46386,N_45614);
and UO_2696 (O_2696,N_47089,N_47503);
nor UO_2697 (O_2697,N_48906,N_48957);
xnor UO_2698 (O_2698,N_49597,N_48534);
xor UO_2699 (O_2699,N_48345,N_45193);
nor UO_2700 (O_2700,N_48489,N_46468);
nor UO_2701 (O_2701,N_47753,N_49620);
nor UO_2702 (O_2702,N_48356,N_48238);
or UO_2703 (O_2703,N_48099,N_47899);
and UO_2704 (O_2704,N_49071,N_45050);
or UO_2705 (O_2705,N_45167,N_46628);
or UO_2706 (O_2706,N_48706,N_45342);
nor UO_2707 (O_2707,N_46770,N_46024);
nor UO_2708 (O_2708,N_49216,N_49365);
nand UO_2709 (O_2709,N_48620,N_49649);
or UO_2710 (O_2710,N_47308,N_46659);
or UO_2711 (O_2711,N_45621,N_47104);
xor UO_2712 (O_2712,N_49730,N_48607);
nand UO_2713 (O_2713,N_45225,N_49240);
nand UO_2714 (O_2714,N_46387,N_49765);
xnor UO_2715 (O_2715,N_47255,N_45512);
or UO_2716 (O_2716,N_45660,N_47503);
and UO_2717 (O_2717,N_48317,N_48085);
or UO_2718 (O_2718,N_45283,N_49034);
nor UO_2719 (O_2719,N_45174,N_49021);
and UO_2720 (O_2720,N_46689,N_46942);
xnor UO_2721 (O_2721,N_49626,N_49092);
and UO_2722 (O_2722,N_45784,N_49688);
or UO_2723 (O_2723,N_45415,N_48131);
xor UO_2724 (O_2724,N_48202,N_49656);
or UO_2725 (O_2725,N_46260,N_49581);
or UO_2726 (O_2726,N_46453,N_48732);
nor UO_2727 (O_2727,N_49933,N_49487);
nand UO_2728 (O_2728,N_49306,N_47117);
or UO_2729 (O_2729,N_49301,N_49661);
nand UO_2730 (O_2730,N_47027,N_47259);
or UO_2731 (O_2731,N_46614,N_48395);
nand UO_2732 (O_2732,N_45910,N_49526);
xnor UO_2733 (O_2733,N_45494,N_47916);
nand UO_2734 (O_2734,N_48722,N_49461);
nand UO_2735 (O_2735,N_47717,N_47619);
nand UO_2736 (O_2736,N_48943,N_47950);
xnor UO_2737 (O_2737,N_46720,N_48640);
xnor UO_2738 (O_2738,N_49175,N_47061);
xor UO_2739 (O_2739,N_45142,N_49977);
and UO_2740 (O_2740,N_46502,N_49785);
or UO_2741 (O_2741,N_45957,N_46492);
xor UO_2742 (O_2742,N_49347,N_48738);
nor UO_2743 (O_2743,N_47281,N_45686);
and UO_2744 (O_2744,N_48772,N_46378);
xnor UO_2745 (O_2745,N_45556,N_46036);
nor UO_2746 (O_2746,N_45741,N_48912);
nor UO_2747 (O_2747,N_49934,N_45654);
or UO_2748 (O_2748,N_47563,N_45689);
nand UO_2749 (O_2749,N_45762,N_46431);
nand UO_2750 (O_2750,N_46961,N_46294);
xor UO_2751 (O_2751,N_48460,N_49823);
or UO_2752 (O_2752,N_47085,N_48784);
nand UO_2753 (O_2753,N_48272,N_45496);
xor UO_2754 (O_2754,N_47328,N_47996);
xor UO_2755 (O_2755,N_49396,N_46585);
nor UO_2756 (O_2756,N_45894,N_48870);
nand UO_2757 (O_2757,N_49031,N_49345);
and UO_2758 (O_2758,N_45610,N_49752);
and UO_2759 (O_2759,N_48849,N_47596);
and UO_2760 (O_2760,N_48845,N_47880);
or UO_2761 (O_2761,N_49158,N_45018);
or UO_2762 (O_2762,N_47254,N_48393);
nor UO_2763 (O_2763,N_46188,N_46269);
nor UO_2764 (O_2764,N_49410,N_49167);
xnor UO_2765 (O_2765,N_45644,N_48130);
nand UO_2766 (O_2766,N_47709,N_48108);
xor UO_2767 (O_2767,N_45061,N_45336);
and UO_2768 (O_2768,N_45891,N_46702);
or UO_2769 (O_2769,N_47240,N_48481);
nor UO_2770 (O_2770,N_47740,N_46014);
or UO_2771 (O_2771,N_48401,N_45157);
and UO_2772 (O_2772,N_48435,N_48222);
nor UO_2773 (O_2773,N_49016,N_48317);
nor UO_2774 (O_2774,N_47124,N_47901);
nor UO_2775 (O_2775,N_46574,N_45187);
xnor UO_2776 (O_2776,N_48133,N_47142);
nor UO_2777 (O_2777,N_48776,N_49582);
xor UO_2778 (O_2778,N_46908,N_47788);
and UO_2779 (O_2779,N_47634,N_49761);
nor UO_2780 (O_2780,N_48105,N_47033);
and UO_2781 (O_2781,N_48185,N_48170);
nor UO_2782 (O_2782,N_48692,N_49136);
nor UO_2783 (O_2783,N_45325,N_45092);
or UO_2784 (O_2784,N_48613,N_48371);
xor UO_2785 (O_2785,N_48073,N_45793);
nand UO_2786 (O_2786,N_45899,N_46602);
nor UO_2787 (O_2787,N_46360,N_45765);
or UO_2788 (O_2788,N_46129,N_48561);
nand UO_2789 (O_2789,N_45428,N_45262);
or UO_2790 (O_2790,N_45738,N_48987);
nand UO_2791 (O_2791,N_46231,N_48721);
or UO_2792 (O_2792,N_46124,N_49102);
nand UO_2793 (O_2793,N_47311,N_46061);
xor UO_2794 (O_2794,N_49110,N_48498);
or UO_2795 (O_2795,N_47412,N_47711);
xor UO_2796 (O_2796,N_49766,N_46118);
nand UO_2797 (O_2797,N_45891,N_47873);
nor UO_2798 (O_2798,N_45546,N_46594);
nand UO_2799 (O_2799,N_45322,N_49098);
nor UO_2800 (O_2800,N_49930,N_49465);
nor UO_2801 (O_2801,N_48671,N_46928);
nor UO_2802 (O_2802,N_45341,N_48200);
and UO_2803 (O_2803,N_46568,N_47966);
nand UO_2804 (O_2804,N_46571,N_49326);
nand UO_2805 (O_2805,N_48074,N_48791);
nor UO_2806 (O_2806,N_49612,N_49773);
and UO_2807 (O_2807,N_45522,N_47792);
or UO_2808 (O_2808,N_47984,N_48001);
nor UO_2809 (O_2809,N_49126,N_49577);
xor UO_2810 (O_2810,N_47093,N_45070);
nand UO_2811 (O_2811,N_47411,N_47194);
and UO_2812 (O_2812,N_48543,N_48338);
nor UO_2813 (O_2813,N_47318,N_48406);
nand UO_2814 (O_2814,N_45279,N_47327);
xor UO_2815 (O_2815,N_47254,N_46715);
or UO_2816 (O_2816,N_48392,N_49107);
and UO_2817 (O_2817,N_47296,N_47494);
nor UO_2818 (O_2818,N_47132,N_48044);
xnor UO_2819 (O_2819,N_47092,N_48724);
and UO_2820 (O_2820,N_47218,N_49445);
and UO_2821 (O_2821,N_47642,N_47420);
nor UO_2822 (O_2822,N_45171,N_47481);
nand UO_2823 (O_2823,N_47330,N_48970);
nand UO_2824 (O_2824,N_48486,N_48234);
nor UO_2825 (O_2825,N_48637,N_47111);
and UO_2826 (O_2826,N_48687,N_46354);
or UO_2827 (O_2827,N_47938,N_46000);
and UO_2828 (O_2828,N_49124,N_47609);
nor UO_2829 (O_2829,N_45817,N_49343);
or UO_2830 (O_2830,N_49779,N_46301);
and UO_2831 (O_2831,N_47353,N_45160);
and UO_2832 (O_2832,N_47040,N_49652);
nand UO_2833 (O_2833,N_49689,N_48408);
or UO_2834 (O_2834,N_49496,N_47958);
nor UO_2835 (O_2835,N_47947,N_49562);
xnor UO_2836 (O_2836,N_45542,N_48062);
xor UO_2837 (O_2837,N_49892,N_46006);
or UO_2838 (O_2838,N_48830,N_46699);
nand UO_2839 (O_2839,N_47932,N_48936);
xor UO_2840 (O_2840,N_47523,N_48475);
nor UO_2841 (O_2841,N_48338,N_48108);
and UO_2842 (O_2842,N_46985,N_45160);
nor UO_2843 (O_2843,N_47144,N_46400);
and UO_2844 (O_2844,N_49255,N_47051);
xor UO_2845 (O_2845,N_48453,N_47071);
and UO_2846 (O_2846,N_47708,N_49248);
or UO_2847 (O_2847,N_45438,N_48315);
nand UO_2848 (O_2848,N_48554,N_47754);
xor UO_2849 (O_2849,N_46784,N_49160);
xnor UO_2850 (O_2850,N_46560,N_45356);
nor UO_2851 (O_2851,N_46000,N_47646);
nor UO_2852 (O_2852,N_47584,N_45953);
nand UO_2853 (O_2853,N_48823,N_45116);
nor UO_2854 (O_2854,N_49195,N_49032);
and UO_2855 (O_2855,N_46526,N_45782);
nand UO_2856 (O_2856,N_45239,N_46676);
nand UO_2857 (O_2857,N_45054,N_47111);
xor UO_2858 (O_2858,N_46820,N_49949);
nor UO_2859 (O_2859,N_46844,N_47011);
or UO_2860 (O_2860,N_47226,N_45837);
nor UO_2861 (O_2861,N_45136,N_45515);
and UO_2862 (O_2862,N_46525,N_49581);
nand UO_2863 (O_2863,N_49122,N_49323);
nor UO_2864 (O_2864,N_46964,N_49407);
and UO_2865 (O_2865,N_49661,N_47641);
or UO_2866 (O_2866,N_48384,N_48554);
or UO_2867 (O_2867,N_45406,N_46223);
nor UO_2868 (O_2868,N_49307,N_48898);
or UO_2869 (O_2869,N_49594,N_47076);
or UO_2870 (O_2870,N_48874,N_48676);
nand UO_2871 (O_2871,N_45270,N_46444);
xnor UO_2872 (O_2872,N_47172,N_45375);
or UO_2873 (O_2873,N_47815,N_47542);
and UO_2874 (O_2874,N_46195,N_46989);
xor UO_2875 (O_2875,N_46263,N_47053);
and UO_2876 (O_2876,N_49041,N_49453);
nand UO_2877 (O_2877,N_45709,N_45272);
xnor UO_2878 (O_2878,N_48142,N_49745);
nor UO_2879 (O_2879,N_45453,N_46874);
xor UO_2880 (O_2880,N_45724,N_46413);
xnor UO_2881 (O_2881,N_47754,N_46867);
nand UO_2882 (O_2882,N_45588,N_49995);
or UO_2883 (O_2883,N_46357,N_45623);
nor UO_2884 (O_2884,N_49956,N_45639);
nand UO_2885 (O_2885,N_47889,N_47559);
xor UO_2886 (O_2886,N_46561,N_49390);
nand UO_2887 (O_2887,N_47792,N_46756);
or UO_2888 (O_2888,N_45483,N_48616);
nand UO_2889 (O_2889,N_47572,N_45594);
nor UO_2890 (O_2890,N_45451,N_45351);
or UO_2891 (O_2891,N_45318,N_49026);
or UO_2892 (O_2892,N_48071,N_49186);
nor UO_2893 (O_2893,N_47812,N_45820);
and UO_2894 (O_2894,N_47103,N_45638);
and UO_2895 (O_2895,N_46784,N_47915);
nor UO_2896 (O_2896,N_49062,N_45845);
or UO_2897 (O_2897,N_46707,N_48989);
and UO_2898 (O_2898,N_46778,N_45565);
or UO_2899 (O_2899,N_49107,N_47206);
nand UO_2900 (O_2900,N_47489,N_48097);
nand UO_2901 (O_2901,N_46073,N_45414);
and UO_2902 (O_2902,N_46990,N_45967);
nor UO_2903 (O_2903,N_46226,N_47708);
or UO_2904 (O_2904,N_45293,N_45115);
nand UO_2905 (O_2905,N_46035,N_48544);
and UO_2906 (O_2906,N_48394,N_46253);
or UO_2907 (O_2907,N_47853,N_49315);
and UO_2908 (O_2908,N_45300,N_49905);
nor UO_2909 (O_2909,N_45159,N_48019);
or UO_2910 (O_2910,N_48043,N_49560);
or UO_2911 (O_2911,N_45919,N_46938);
nor UO_2912 (O_2912,N_48331,N_48970);
nand UO_2913 (O_2913,N_46465,N_46454);
and UO_2914 (O_2914,N_48325,N_48865);
xnor UO_2915 (O_2915,N_46029,N_49048);
xnor UO_2916 (O_2916,N_46762,N_47899);
nand UO_2917 (O_2917,N_49723,N_46745);
or UO_2918 (O_2918,N_45347,N_46767);
nand UO_2919 (O_2919,N_49850,N_49123);
nor UO_2920 (O_2920,N_45920,N_48092);
nor UO_2921 (O_2921,N_46407,N_48369);
nor UO_2922 (O_2922,N_47540,N_47181);
or UO_2923 (O_2923,N_45924,N_47126);
and UO_2924 (O_2924,N_46363,N_49021);
nand UO_2925 (O_2925,N_45952,N_47628);
xnor UO_2926 (O_2926,N_48369,N_45007);
xnor UO_2927 (O_2927,N_46672,N_47227);
and UO_2928 (O_2928,N_47222,N_48556);
and UO_2929 (O_2929,N_46212,N_46415);
and UO_2930 (O_2930,N_49084,N_48904);
and UO_2931 (O_2931,N_48602,N_45773);
and UO_2932 (O_2932,N_47555,N_47688);
nor UO_2933 (O_2933,N_48659,N_45520);
or UO_2934 (O_2934,N_48910,N_45049);
xnor UO_2935 (O_2935,N_49477,N_47859);
xnor UO_2936 (O_2936,N_45189,N_47187);
nor UO_2937 (O_2937,N_47570,N_48002);
and UO_2938 (O_2938,N_49405,N_48342);
and UO_2939 (O_2939,N_45148,N_47222);
or UO_2940 (O_2940,N_47633,N_45703);
nand UO_2941 (O_2941,N_49313,N_48929);
nand UO_2942 (O_2942,N_45823,N_49328);
nand UO_2943 (O_2943,N_47140,N_45260);
or UO_2944 (O_2944,N_46398,N_49790);
xnor UO_2945 (O_2945,N_45875,N_47281);
xor UO_2946 (O_2946,N_48242,N_48359);
nor UO_2947 (O_2947,N_47866,N_49093);
nand UO_2948 (O_2948,N_49512,N_46788);
and UO_2949 (O_2949,N_47766,N_47204);
nand UO_2950 (O_2950,N_45024,N_45841);
nand UO_2951 (O_2951,N_45019,N_49805);
nor UO_2952 (O_2952,N_46644,N_49417);
xor UO_2953 (O_2953,N_47089,N_47170);
xor UO_2954 (O_2954,N_47720,N_49806);
or UO_2955 (O_2955,N_45476,N_48476);
nor UO_2956 (O_2956,N_47005,N_47314);
and UO_2957 (O_2957,N_49039,N_46530);
nand UO_2958 (O_2958,N_47000,N_46131);
nand UO_2959 (O_2959,N_48992,N_45805);
nor UO_2960 (O_2960,N_47485,N_46652);
nand UO_2961 (O_2961,N_47249,N_48727);
xnor UO_2962 (O_2962,N_47550,N_47582);
and UO_2963 (O_2963,N_49146,N_47261);
and UO_2964 (O_2964,N_46483,N_47549);
xnor UO_2965 (O_2965,N_46050,N_48506);
nor UO_2966 (O_2966,N_49364,N_49470);
xor UO_2967 (O_2967,N_47371,N_49799);
xor UO_2968 (O_2968,N_48275,N_46144);
nand UO_2969 (O_2969,N_47065,N_48842);
nor UO_2970 (O_2970,N_46021,N_49217);
nor UO_2971 (O_2971,N_48110,N_45883);
nand UO_2972 (O_2972,N_48267,N_47312);
xnor UO_2973 (O_2973,N_47799,N_48201);
nor UO_2974 (O_2974,N_47177,N_46857);
xor UO_2975 (O_2975,N_47689,N_46742);
or UO_2976 (O_2976,N_47210,N_46658);
or UO_2977 (O_2977,N_46250,N_48553);
nor UO_2978 (O_2978,N_45587,N_46089);
nand UO_2979 (O_2979,N_46917,N_46172);
or UO_2980 (O_2980,N_48181,N_49307);
and UO_2981 (O_2981,N_48922,N_49863);
nand UO_2982 (O_2982,N_46006,N_49654);
nand UO_2983 (O_2983,N_49634,N_49504);
nand UO_2984 (O_2984,N_49986,N_48829);
xnor UO_2985 (O_2985,N_45517,N_47664);
nand UO_2986 (O_2986,N_45639,N_47247);
nor UO_2987 (O_2987,N_46696,N_48003);
xnor UO_2988 (O_2988,N_46068,N_48033);
or UO_2989 (O_2989,N_48115,N_46492);
xor UO_2990 (O_2990,N_46250,N_49920);
nor UO_2991 (O_2991,N_48255,N_45923);
xnor UO_2992 (O_2992,N_46790,N_49475);
or UO_2993 (O_2993,N_49219,N_48900);
nand UO_2994 (O_2994,N_45359,N_46449);
and UO_2995 (O_2995,N_45114,N_47154);
xnor UO_2996 (O_2996,N_49016,N_46664);
or UO_2997 (O_2997,N_45228,N_46849);
nor UO_2998 (O_2998,N_48895,N_49373);
or UO_2999 (O_2999,N_46112,N_46750);
xnor UO_3000 (O_3000,N_48874,N_45890);
nor UO_3001 (O_3001,N_46217,N_49682);
nand UO_3002 (O_3002,N_49921,N_46343);
nand UO_3003 (O_3003,N_48542,N_49999);
nor UO_3004 (O_3004,N_49968,N_47271);
nor UO_3005 (O_3005,N_49228,N_45573);
or UO_3006 (O_3006,N_48284,N_49293);
xnor UO_3007 (O_3007,N_49370,N_46790);
and UO_3008 (O_3008,N_48725,N_47494);
nand UO_3009 (O_3009,N_48112,N_48377);
nor UO_3010 (O_3010,N_45890,N_48421);
nand UO_3011 (O_3011,N_45956,N_49872);
and UO_3012 (O_3012,N_47834,N_45845);
nand UO_3013 (O_3013,N_45693,N_49066);
and UO_3014 (O_3014,N_47158,N_45872);
nand UO_3015 (O_3015,N_45014,N_46933);
nand UO_3016 (O_3016,N_45624,N_46935);
or UO_3017 (O_3017,N_47298,N_48183);
nor UO_3018 (O_3018,N_49032,N_48581);
nand UO_3019 (O_3019,N_45563,N_46366);
nand UO_3020 (O_3020,N_49758,N_46874);
and UO_3021 (O_3021,N_46053,N_46570);
or UO_3022 (O_3022,N_49846,N_45977);
xor UO_3023 (O_3023,N_48082,N_45466);
xor UO_3024 (O_3024,N_45790,N_49683);
nor UO_3025 (O_3025,N_46300,N_45128);
xnor UO_3026 (O_3026,N_49744,N_47994);
nor UO_3027 (O_3027,N_47050,N_46909);
xnor UO_3028 (O_3028,N_46471,N_48130);
xor UO_3029 (O_3029,N_49315,N_46448);
and UO_3030 (O_3030,N_48683,N_48354);
nand UO_3031 (O_3031,N_45010,N_45571);
nor UO_3032 (O_3032,N_48630,N_47224);
nand UO_3033 (O_3033,N_47810,N_49511);
xnor UO_3034 (O_3034,N_46433,N_45721);
nor UO_3035 (O_3035,N_49006,N_47721);
or UO_3036 (O_3036,N_48134,N_45069);
and UO_3037 (O_3037,N_48642,N_46832);
and UO_3038 (O_3038,N_47111,N_47621);
xnor UO_3039 (O_3039,N_48716,N_48765);
or UO_3040 (O_3040,N_49940,N_49594);
xor UO_3041 (O_3041,N_48692,N_46971);
or UO_3042 (O_3042,N_45720,N_48215);
or UO_3043 (O_3043,N_45668,N_48211);
nand UO_3044 (O_3044,N_45368,N_49171);
xor UO_3045 (O_3045,N_47767,N_48320);
or UO_3046 (O_3046,N_47532,N_48691);
and UO_3047 (O_3047,N_45262,N_47697);
or UO_3048 (O_3048,N_49182,N_46449);
nor UO_3049 (O_3049,N_46824,N_46020);
and UO_3050 (O_3050,N_46649,N_47762);
or UO_3051 (O_3051,N_49122,N_45238);
or UO_3052 (O_3052,N_48558,N_48600);
and UO_3053 (O_3053,N_47217,N_49088);
and UO_3054 (O_3054,N_48001,N_49483);
or UO_3055 (O_3055,N_49006,N_49086);
and UO_3056 (O_3056,N_47581,N_46117);
nand UO_3057 (O_3057,N_45724,N_47657);
nor UO_3058 (O_3058,N_49230,N_45736);
nand UO_3059 (O_3059,N_48195,N_47972);
or UO_3060 (O_3060,N_49547,N_49445);
or UO_3061 (O_3061,N_48195,N_45305);
nor UO_3062 (O_3062,N_49177,N_45641);
or UO_3063 (O_3063,N_48191,N_46231);
nand UO_3064 (O_3064,N_45967,N_49833);
nand UO_3065 (O_3065,N_49301,N_49286);
nor UO_3066 (O_3066,N_46173,N_46181);
or UO_3067 (O_3067,N_47107,N_47234);
or UO_3068 (O_3068,N_45816,N_47714);
and UO_3069 (O_3069,N_45965,N_49410);
and UO_3070 (O_3070,N_48006,N_46461);
or UO_3071 (O_3071,N_45241,N_45445);
and UO_3072 (O_3072,N_46050,N_49469);
and UO_3073 (O_3073,N_49587,N_46473);
xnor UO_3074 (O_3074,N_45841,N_46984);
nand UO_3075 (O_3075,N_49980,N_47498);
xnor UO_3076 (O_3076,N_49615,N_46248);
or UO_3077 (O_3077,N_49332,N_46997);
nor UO_3078 (O_3078,N_48460,N_46534);
nand UO_3079 (O_3079,N_47064,N_48554);
and UO_3080 (O_3080,N_49097,N_47569);
nor UO_3081 (O_3081,N_45735,N_48726);
xnor UO_3082 (O_3082,N_47399,N_47314);
or UO_3083 (O_3083,N_49726,N_46787);
and UO_3084 (O_3084,N_48997,N_47039);
nor UO_3085 (O_3085,N_49248,N_46829);
or UO_3086 (O_3086,N_45494,N_47329);
nand UO_3087 (O_3087,N_49230,N_46845);
nand UO_3088 (O_3088,N_47643,N_48101);
and UO_3089 (O_3089,N_49219,N_47707);
nor UO_3090 (O_3090,N_45179,N_46244);
or UO_3091 (O_3091,N_48558,N_46956);
nand UO_3092 (O_3092,N_46583,N_46590);
nand UO_3093 (O_3093,N_49109,N_47897);
xor UO_3094 (O_3094,N_49472,N_47568);
xnor UO_3095 (O_3095,N_49346,N_46374);
xnor UO_3096 (O_3096,N_48372,N_49053);
nor UO_3097 (O_3097,N_48694,N_47887);
and UO_3098 (O_3098,N_45323,N_49247);
nand UO_3099 (O_3099,N_46849,N_45097);
and UO_3100 (O_3100,N_49686,N_45389);
nand UO_3101 (O_3101,N_48681,N_49836);
or UO_3102 (O_3102,N_46286,N_49789);
and UO_3103 (O_3103,N_49094,N_49470);
xor UO_3104 (O_3104,N_47943,N_45885);
and UO_3105 (O_3105,N_49104,N_46042);
and UO_3106 (O_3106,N_47640,N_47838);
nor UO_3107 (O_3107,N_47838,N_48751);
nand UO_3108 (O_3108,N_47154,N_47261);
xor UO_3109 (O_3109,N_49608,N_47563);
nand UO_3110 (O_3110,N_45644,N_45540);
or UO_3111 (O_3111,N_48885,N_47602);
xnor UO_3112 (O_3112,N_46909,N_47349);
nor UO_3113 (O_3113,N_48099,N_48717);
nand UO_3114 (O_3114,N_49297,N_45635);
and UO_3115 (O_3115,N_45608,N_48641);
xnor UO_3116 (O_3116,N_49925,N_49579);
nor UO_3117 (O_3117,N_45396,N_46731);
nor UO_3118 (O_3118,N_47391,N_48742);
nand UO_3119 (O_3119,N_45479,N_46016);
xnor UO_3120 (O_3120,N_46895,N_49767);
or UO_3121 (O_3121,N_46900,N_48317);
or UO_3122 (O_3122,N_45735,N_48824);
nor UO_3123 (O_3123,N_45595,N_47087);
nand UO_3124 (O_3124,N_48121,N_48462);
nor UO_3125 (O_3125,N_49905,N_49992);
and UO_3126 (O_3126,N_48126,N_48069);
and UO_3127 (O_3127,N_45618,N_49227);
nor UO_3128 (O_3128,N_47666,N_46655);
or UO_3129 (O_3129,N_46273,N_45212);
or UO_3130 (O_3130,N_45183,N_45553);
or UO_3131 (O_3131,N_45023,N_47111);
xnor UO_3132 (O_3132,N_46300,N_46705);
nand UO_3133 (O_3133,N_46653,N_49768);
or UO_3134 (O_3134,N_49081,N_46048);
xor UO_3135 (O_3135,N_45117,N_49138);
or UO_3136 (O_3136,N_47864,N_45330);
and UO_3137 (O_3137,N_49723,N_45169);
or UO_3138 (O_3138,N_47308,N_48335);
xor UO_3139 (O_3139,N_46039,N_45585);
nand UO_3140 (O_3140,N_45149,N_45816);
nand UO_3141 (O_3141,N_46262,N_46518);
nor UO_3142 (O_3142,N_49313,N_47508);
nand UO_3143 (O_3143,N_49750,N_45517);
or UO_3144 (O_3144,N_47428,N_46715);
nor UO_3145 (O_3145,N_46307,N_45036);
nand UO_3146 (O_3146,N_48911,N_45295);
nand UO_3147 (O_3147,N_48009,N_47314);
or UO_3148 (O_3148,N_49917,N_46888);
xnor UO_3149 (O_3149,N_47144,N_49629);
and UO_3150 (O_3150,N_49033,N_45359);
and UO_3151 (O_3151,N_47687,N_46956);
nor UO_3152 (O_3152,N_48714,N_45389);
or UO_3153 (O_3153,N_49875,N_49920);
and UO_3154 (O_3154,N_47082,N_49547);
nand UO_3155 (O_3155,N_46216,N_49882);
xnor UO_3156 (O_3156,N_45851,N_47398);
nand UO_3157 (O_3157,N_48941,N_49665);
nand UO_3158 (O_3158,N_45947,N_47114);
xor UO_3159 (O_3159,N_48929,N_46845);
nand UO_3160 (O_3160,N_48581,N_49231);
nand UO_3161 (O_3161,N_46764,N_47924);
nor UO_3162 (O_3162,N_49677,N_47942);
or UO_3163 (O_3163,N_49244,N_49496);
nor UO_3164 (O_3164,N_49485,N_49875);
nand UO_3165 (O_3165,N_46501,N_49802);
or UO_3166 (O_3166,N_45543,N_45849);
and UO_3167 (O_3167,N_46020,N_46535);
nand UO_3168 (O_3168,N_48272,N_46513);
xor UO_3169 (O_3169,N_49902,N_47407);
xor UO_3170 (O_3170,N_45016,N_46416);
xnor UO_3171 (O_3171,N_48898,N_49556);
nand UO_3172 (O_3172,N_48496,N_46143);
nor UO_3173 (O_3173,N_45159,N_47893);
nor UO_3174 (O_3174,N_49490,N_45908);
nand UO_3175 (O_3175,N_47211,N_49076);
nor UO_3176 (O_3176,N_49950,N_45085);
nand UO_3177 (O_3177,N_46389,N_47243);
xnor UO_3178 (O_3178,N_45873,N_46048);
xor UO_3179 (O_3179,N_48650,N_47728);
nand UO_3180 (O_3180,N_49868,N_46682);
xor UO_3181 (O_3181,N_49873,N_49808);
nand UO_3182 (O_3182,N_47556,N_49938);
or UO_3183 (O_3183,N_46174,N_47248);
nand UO_3184 (O_3184,N_47263,N_47622);
nand UO_3185 (O_3185,N_48808,N_45283);
nor UO_3186 (O_3186,N_48736,N_46684);
nand UO_3187 (O_3187,N_49561,N_45623);
xnor UO_3188 (O_3188,N_45917,N_46452);
and UO_3189 (O_3189,N_46466,N_49389);
nand UO_3190 (O_3190,N_49824,N_45278);
xnor UO_3191 (O_3191,N_49645,N_46456);
nor UO_3192 (O_3192,N_47689,N_46751);
nand UO_3193 (O_3193,N_46904,N_45243);
xor UO_3194 (O_3194,N_45001,N_48225);
and UO_3195 (O_3195,N_48718,N_49134);
xor UO_3196 (O_3196,N_49755,N_47072);
xnor UO_3197 (O_3197,N_45742,N_47379);
or UO_3198 (O_3198,N_48299,N_45387);
nand UO_3199 (O_3199,N_47829,N_45535);
and UO_3200 (O_3200,N_49333,N_46028);
nand UO_3201 (O_3201,N_48964,N_46373);
nand UO_3202 (O_3202,N_48808,N_49797);
nand UO_3203 (O_3203,N_47080,N_46941);
xnor UO_3204 (O_3204,N_48014,N_47280);
nand UO_3205 (O_3205,N_46128,N_46427);
nor UO_3206 (O_3206,N_45231,N_48749);
xnor UO_3207 (O_3207,N_49353,N_46034);
nand UO_3208 (O_3208,N_46920,N_48086);
nand UO_3209 (O_3209,N_49804,N_48211);
nand UO_3210 (O_3210,N_49358,N_47638);
and UO_3211 (O_3211,N_46565,N_48330);
xor UO_3212 (O_3212,N_45083,N_47488);
xnor UO_3213 (O_3213,N_47418,N_49707);
nand UO_3214 (O_3214,N_47780,N_48424);
or UO_3215 (O_3215,N_46424,N_48211);
or UO_3216 (O_3216,N_45136,N_48273);
nand UO_3217 (O_3217,N_49158,N_45521);
xnor UO_3218 (O_3218,N_49262,N_45359);
and UO_3219 (O_3219,N_45488,N_46509);
and UO_3220 (O_3220,N_45868,N_48643);
or UO_3221 (O_3221,N_48284,N_46807);
xnor UO_3222 (O_3222,N_47791,N_48856);
and UO_3223 (O_3223,N_48409,N_49318);
nand UO_3224 (O_3224,N_48588,N_48360);
xor UO_3225 (O_3225,N_45573,N_48123);
nor UO_3226 (O_3226,N_48923,N_49633);
nor UO_3227 (O_3227,N_48483,N_49384);
and UO_3228 (O_3228,N_49574,N_47825);
xnor UO_3229 (O_3229,N_47768,N_48452);
nor UO_3230 (O_3230,N_46300,N_45254);
or UO_3231 (O_3231,N_49556,N_45184);
and UO_3232 (O_3232,N_47735,N_48838);
nand UO_3233 (O_3233,N_46089,N_46536);
xor UO_3234 (O_3234,N_45743,N_49198);
and UO_3235 (O_3235,N_45162,N_48434);
nand UO_3236 (O_3236,N_47098,N_46780);
xnor UO_3237 (O_3237,N_49811,N_48541);
or UO_3238 (O_3238,N_45607,N_49096);
and UO_3239 (O_3239,N_46236,N_47961);
xor UO_3240 (O_3240,N_46225,N_45676);
nor UO_3241 (O_3241,N_46978,N_45101);
xnor UO_3242 (O_3242,N_49395,N_48891);
and UO_3243 (O_3243,N_45614,N_46873);
xnor UO_3244 (O_3244,N_45969,N_48868);
nand UO_3245 (O_3245,N_47572,N_49107);
xor UO_3246 (O_3246,N_46364,N_49676);
and UO_3247 (O_3247,N_49717,N_48478);
and UO_3248 (O_3248,N_48946,N_46127);
or UO_3249 (O_3249,N_47505,N_49098);
nor UO_3250 (O_3250,N_49639,N_49014);
nor UO_3251 (O_3251,N_49095,N_45757);
and UO_3252 (O_3252,N_48637,N_47683);
and UO_3253 (O_3253,N_49502,N_48753);
and UO_3254 (O_3254,N_48928,N_46613);
nor UO_3255 (O_3255,N_48733,N_49791);
xor UO_3256 (O_3256,N_46081,N_47591);
xnor UO_3257 (O_3257,N_48176,N_48522);
nand UO_3258 (O_3258,N_46577,N_46059);
or UO_3259 (O_3259,N_46136,N_46815);
and UO_3260 (O_3260,N_46628,N_47426);
and UO_3261 (O_3261,N_48169,N_49590);
nor UO_3262 (O_3262,N_48184,N_47211);
and UO_3263 (O_3263,N_46203,N_46481);
or UO_3264 (O_3264,N_45862,N_48936);
or UO_3265 (O_3265,N_46007,N_49286);
and UO_3266 (O_3266,N_46686,N_46095);
nand UO_3267 (O_3267,N_47479,N_45090);
and UO_3268 (O_3268,N_45860,N_49745);
xnor UO_3269 (O_3269,N_46920,N_46838);
and UO_3270 (O_3270,N_45176,N_49439);
and UO_3271 (O_3271,N_47712,N_46463);
nor UO_3272 (O_3272,N_45941,N_48041);
nor UO_3273 (O_3273,N_47086,N_47712);
or UO_3274 (O_3274,N_45978,N_47147);
nor UO_3275 (O_3275,N_49694,N_49114);
or UO_3276 (O_3276,N_46249,N_45946);
nand UO_3277 (O_3277,N_47362,N_48983);
xnor UO_3278 (O_3278,N_49903,N_45731);
or UO_3279 (O_3279,N_45176,N_48939);
nor UO_3280 (O_3280,N_47618,N_46873);
or UO_3281 (O_3281,N_47269,N_48285);
nand UO_3282 (O_3282,N_47856,N_47299);
nand UO_3283 (O_3283,N_49076,N_49072);
nor UO_3284 (O_3284,N_49162,N_49534);
or UO_3285 (O_3285,N_49005,N_46412);
nand UO_3286 (O_3286,N_49648,N_47468);
xnor UO_3287 (O_3287,N_48894,N_48979);
nor UO_3288 (O_3288,N_46044,N_46061);
or UO_3289 (O_3289,N_48243,N_48911);
and UO_3290 (O_3290,N_45243,N_48388);
nor UO_3291 (O_3291,N_45270,N_49871);
xor UO_3292 (O_3292,N_48613,N_49558);
xor UO_3293 (O_3293,N_46383,N_48698);
and UO_3294 (O_3294,N_45200,N_48715);
and UO_3295 (O_3295,N_49107,N_46976);
nand UO_3296 (O_3296,N_46149,N_48779);
or UO_3297 (O_3297,N_47791,N_47252);
xnor UO_3298 (O_3298,N_48781,N_47050);
nand UO_3299 (O_3299,N_45780,N_45988);
or UO_3300 (O_3300,N_47132,N_48049);
xor UO_3301 (O_3301,N_46052,N_47993);
nor UO_3302 (O_3302,N_45892,N_46475);
or UO_3303 (O_3303,N_49300,N_48894);
nand UO_3304 (O_3304,N_46387,N_45076);
nor UO_3305 (O_3305,N_47199,N_48230);
xnor UO_3306 (O_3306,N_48447,N_46261);
xor UO_3307 (O_3307,N_48538,N_46850);
nand UO_3308 (O_3308,N_49979,N_46007);
or UO_3309 (O_3309,N_46204,N_48761);
nor UO_3310 (O_3310,N_45430,N_49701);
xnor UO_3311 (O_3311,N_47271,N_47305);
and UO_3312 (O_3312,N_48984,N_45454);
nand UO_3313 (O_3313,N_47693,N_45175);
nand UO_3314 (O_3314,N_47985,N_47569);
xnor UO_3315 (O_3315,N_45527,N_46632);
nor UO_3316 (O_3316,N_46156,N_49371);
or UO_3317 (O_3317,N_49112,N_48635);
nand UO_3318 (O_3318,N_49116,N_48943);
xnor UO_3319 (O_3319,N_46415,N_45001);
nand UO_3320 (O_3320,N_49098,N_48992);
xor UO_3321 (O_3321,N_48247,N_48910);
or UO_3322 (O_3322,N_47859,N_49097);
and UO_3323 (O_3323,N_45459,N_47180);
xor UO_3324 (O_3324,N_47457,N_47773);
nand UO_3325 (O_3325,N_48667,N_49624);
xor UO_3326 (O_3326,N_49173,N_48252);
nand UO_3327 (O_3327,N_49604,N_47052);
xor UO_3328 (O_3328,N_49741,N_47031);
or UO_3329 (O_3329,N_49730,N_46061);
nand UO_3330 (O_3330,N_47359,N_48001);
and UO_3331 (O_3331,N_49829,N_48970);
or UO_3332 (O_3332,N_46682,N_46461);
nor UO_3333 (O_3333,N_45639,N_47742);
and UO_3334 (O_3334,N_46557,N_48180);
nor UO_3335 (O_3335,N_49074,N_46282);
nand UO_3336 (O_3336,N_47666,N_45103);
nand UO_3337 (O_3337,N_46960,N_46995);
nand UO_3338 (O_3338,N_49564,N_47191);
xor UO_3339 (O_3339,N_49569,N_48069);
or UO_3340 (O_3340,N_49572,N_48855);
and UO_3341 (O_3341,N_45663,N_48094);
xnor UO_3342 (O_3342,N_45702,N_49400);
nor UO_3343 (O_3343,N_49793,N_47784);
nor UO_3344 (O_3344,N_46256,N_47811);
xor UO_3345 (O_3345,N_48489,N_47327);
nand UO_3346 (O_3346,N_47349,N_46006);
or UO_3347 (O_3347,N_46985,N_49988);
or UO_3348 (O_3348,N_47681,N_49586);
nand UO_3349 (O_3349,N_47746,N_46744);
xnor UO_3350 (O_3350,N_47107,N_46377);
nand UO_3351 (O_3351,N_48841,N_48793);
xor UO_3352 (O_3352,N_45662,N_46971);
nor UO_3353 (O_3353,N_46796,N_47819);
nand UO_3354 (O_3354,N_48275,N_45935);
or UO_3355 (O_3355,N_45495,N_48407);
and UO_3356 (O_3356,N_46502,N_47637);
nand UO_3357 (O_3357,N_48749,N_45152);
nor UO_3358 (O_3358,N_46491,N_47034);
xnor UO_3359 (O_3359,N_45102,N_45565);
nand UO_3360 (O_3360,N_49297,N_49911);
and UO_3361 (O_3361,N_46501,N_47590);
xor UO_3362 (O_3362,N_45617,N_47846);
xnor UO_3363 (O_3363,N_46740,N_49194);
or UO_3364 (O_3364,N_47586,N_48193);
and UO_3365 (O_3365,N_49911,N_47042);
or UO_3366 (O_3366,N_47094,N_47071);
nand UO_3367 (O_3367,N_48074,N_46054);
and UO_3368 (O_3368,N_47247,N_45354);
nor UO_3369 (O_3369,N_49977,N_49425);
nor UO_3370 (O_3370,N_46649,N_45916);
xor UO_3371 (O_3371,N_47414,N_48707);
and UO_3372 (O_3372,N_48933,N_46369);
xnor UO_3373 (O_3373,N_46237,N_46352);
xor UO_3374 (O_3374,N_47776,N_45643);
and UO_3375 (O_3375,N_47157,N_47343);
nand UO_3376 (O_3376,N_45662,N_45366);
nand UO_3377 (O_3377,N_46260,N_49286);
and UO_3378 (O_3378,N_45202,N_46613);
xnor UO_3379 (O_3379,N_47863,N_49328);
or UO_3380 (O_3380,N_45485,N_47621);
nand UO_3381 (O_3381,N_47237,N_45074);
nand UO_3382 (O_3382,N_47260,N_47330);
or UO_3383 (O_3383,N_49680,N_46897);
nand UO_3384 (O_3384,N_45675,N_45687);
nor UO_3385 (O_3385,N_48084,N_46250);
xnor UO_3386 (O_3386,N_46445,N_45782);
nor UO_3387 (O_3387,N_47250,N_45743);
and UO_3388 (O_3388,N_49510,N_46741);
or UO_3389 (O_3389,N_45026,N_45461);
xor UO_3390 (O_3390,N_47459,N_48670);
or UO_3391 (O_3391,N_49411,N_48649);
nand UO_3392 (O_3392,N_48311,N_48429);
and UO_3393 (O_3393,N_48631,N_48242);
and UO_3394 (O_3394,N_49352,N_45081);
nand UO_3395 (O_3395,N_45937,N_48131);
and UO_3396 (O_3396,N_47554,N_45195);
xor UO_3397 (O_3397,N_47440,N_45087);
nand UO_3398 (O_3398,N_47215,N_49664);
xnor UO_3399 (O_3399,N_48694,N_47486);
or UO_3400 (O_3400,N_48777,N_45515);
and UO_3401 (O_3401,N_49930,N_48788);
xnor UO_3402 (O_3402,N_46914,N_46713);
or UO_3403 (O_3403,N_48614,N_45950);
or UO_3404 (O_3404,N_46163,N_48405);
nand UO_3405 (O_3405,N_48238,N_46390);
and UO_3406 (O_3406,N_47818,N_46336);
or UO_3407 (O_3407,N_47745,N_46478);
and UO_3408 (O_3408,N_45170,N_47349);
xnor UO_3409 (O_3409,N_49240,N_46614);
and UO_3410 (O_3410,N_49760,N_49992);
xor UO_3411 (O_3411,N_49425,N_48329);
xor UO_3412 (O_3412,N_47922,N_48636);
and UO_3413 (O_3413,N_47847,N_48340);
and UO_3414 (O_3414,N_48845,N_46175);
nor UO_3415 (O_3415,N_46121,N_45221);
and UO_3416 (O_3416,N_48624,N_46293);
xnor UO_3417 (O_3417,N_45726,N_49942);
or UO_3418 (O_3418,N_47374,N_48999);
xnor UO_3419 (O_3419,N_48603,N_46826);
nand UO_3420 (O_3420,N_48334,N_47394);
nand UO_3421 (O_3421,N_46900,N_45167);
and UO_3422 (O_3422,N_48747,N_46122);
nor UO_3423 (O_3423,N_49544,N_45778);
or UO_3424 (O_3424,N_48622,N_49522);
xnor UO_3425 (O_3425,N_45719,N_46825);
nand UO_3426 (O_3426,N_46032,N_45883);
and UO_3427 (O_3427,N_49309,N_46966);
xnor UO_3428 (O_3428,N_45747,N_45831);
or UO_3429 (O_3429,N_45229,N_46870);
xnor UO_3430 (O_3430,N_49591,N_49727);
nand UO_3431 (O_3431,N_48901,N_48588);
xor UO_3432 (O_3432,N_46636,N_45980);
or UO_3433 (O_3433,N_45753,N_48034);
and UO_3434 (O_3434,N_48470,N_48050);
nor UO_3435 (O_3435,N_46207,N_47281);
or UO_3436 (O_3436,N_48141,N_46947);
xnor UO_3437 (O_3437,N_45231,N_45795);
xnor UO_3438 (O_3438,N_45458,N_49333);
xor UO_3439 (O_3439,N_46588,N_49882);
and UO_3440 (O_3440,N_45853,N_48691);
nand UO_3441 (O_3441,N_47166,N_49078);
or UO_3442 (O_3442,N_49127,N_46988);
xnor UO_3443 (O_3443,N_49405,N_48951);
and UO_3444 (O_3444,N_46965,N_47494);
and UO_3445 (O_3445,N_48157,N_48884);
nand UO_3446 (O_3446,N_46056,N_45431);
and UO_3447 (O_3447,N_46555,N_49616);
and UO_3448 (O_3448,N_48303,N_45711);
nor UO_3449 (O_3449,N_47613,N_48220);
or UO_3450 (O_3450,N_48672,N_45736);
xnor UO_3451 (O_3451,N_48589,N_47088);
and UO_3452 (O_3452,N_48095,N_49889);
xnor UO_3453 (O_3453,N_45970,N_48451);
nor UO_3454 (O_3454,N_47256,N_45708);
nor UO_3455 (O_3455,N_49918,N_48011);
or UO_3456 (O_3456,N_47287,N_45185);
nand UO_3457 (O_3457,N_48926,N_46648);
or UO_3458 (O_3458,N_45843,N_47920);
or UO_3459 (O_3459,N_49282,N_46444);
nor UO_3460 (O_3460,N_48579,N_45650);
xor UO_3461 (O_3461,N_49299,N_49336);
nand UO_3462 (O_3462,N_48302,N_48842);
and UO_3463 (O_3463,N_45180,N_45388);
xnor UO_3464 (O_3464,N_47544,N_49596);
nor UO_3465 (O_3465,N_45625,N_46746);
nor UO_3466 (O_3466,N_47309,N_49028);
xnor UO_3467 (O_3467,N_47522,N_49914);
xnor UO_3468 (O_3468,N_48501,N_45007);
and UO_3469 (O_3469,N_45157,N_45448);
nand UO_3470 (O_3470,N_46119,N_46057);
nand UO_3471 (O_3471,N_49109,N_48981);
nand UO_3472 (O_3472,N_46101,N_48875);
xor UO_3473 (O_3473,N_45355,N_46914);
or UO_3474 (O_3474,N_47010,N_45772);
or UO_3475 (O_3475,N_48124,N_47543);
xnor UO_3476 (O_3476,N_46608,N_45353);
nor UO_3477 (O_3477,N_49392,N_46864);
or UO_3478 (O_3478,N_47595,N_48055);
nor UO_3479 (O_3479,N_46634,N_46195);
and UO_3480 (O_3480,N_49376,N_47792);
nor UO_3481 (O_3481,N_49649,N_46657);
nor UO_3482 (O_3482,N_45598,N_46401);
nand UO_3483 (O_3483,N_46205,N_48312);
nand UO_3484 (O_3484,N_49092,N_46024);
and UO_3485 (O_3485,N_49006,N_49611);
nand UO_3486 (O_3486,N_49635,N_47346);
and UO_3487 (O_3487,N_48800,N_46752);
xor UO_3488 (O_3488,N_49932,N_45248);
and UO_3489 (O_3489,N_46702,N_47998);
nor UO_3490 (O_3490,N_46881,N_46504);
or UO_3491 (O_3491,N_46852,N_49125);
and UO_3492 (O_3492,N_46473,N_47106);
xnor UO_3493 (O_3493,N_48756,N_46771);
and UO_3494 (O_3494,N_48385,N_49073);
xnor UO_3495 (O_3495,N_47840,N_49490);
or UO_3496 (O_3496,N_49763,N_48008);
xor UO_3497 (O_3497,N_46609,N_49027);
xor UO_3498 (O_3498,N_45858,N_47701);
xnor UO_3499 (O_3499,N_48457,N_48612);
or UO_3500 (O_3500,N_45254,N_46819);
and UO_3501 (O_3501,N_48526,N_45604);
and UO_3502 (O_3502,N_47363,N_49550);
xor UO_3503 (O_3503,N_49921,N_47201);
nor UO_3504 (O_3504,N_47993,N_49308);
nor UO_3505 (O_3505,N_46951,N_48703);
nand UO_3506 (O_3506,N_49420,N_46928);
nor UO_3507 (O_3507,N_45733,N_47617);
and UO_3508 (O_3508,N_48890,N_48844);
xnor UO_3509 (O_3509,N_48836,N_48899);
nor UO_3510 (O_3510,N_48160,N_49020);
xnor UO_3511 (O_3511,N_49855,N_48993);
nor UO_3512 (O_3512,N_47095,N_45533);
or UO_3513 (O_3513,N_46403,N_45100);
nor UO_3514 (O_3514,N_49930,N_48092);
nor UO_3515 (O_3515,N_47884,N_45158);
or UO_3516 (O_3516,N_47404,N_46944);
and UO_3517 (O_3517,N_45980,N_49116);
nor UO_3518 (O_3518,N_49021,N_46081);
and UO_3519 (O_3519,N_48466,N_48917);
and UO_3520 (O_3520,N_47199,N_47803);
or UO_3521 (O_3521,N_48544,N_45738);
nor UO_3522 (O_3522,N_48742,N_45837);
nor UO_3523 (O_3523,N_45370,N_45372);
and UO_3524 (O_3524,N_45377,N_46997);
nor UO_3525 (O_3525,N_46649,N_47464);
nand UO_3526 (O_3526,N_47053,N_49716);
nand UO_3527 (O_3527,N_46129,N_49374);
or UO_3528 (O_3528,N_45903,N_47262);
xor UO_3529 (O_3529,N_46588,N_46004);
nand UO_3530 (O_3530,N_45184,N_47705);
xor UO_3531 (O_3531,N_49126,N_47393);
or UO_3532 (O_3532,N_49628,N_47100);
nand UO_3533 (O_3533,N_48536,N_46916);
nor UO_3534 (O_3534,N_46808,N_45279);
nand UO_3535 (O_3535,N_47018,N_47755);
or UO_3536 (O_3536,N_45476,N_46324);
or UO_3537 (O_3537,N_46933,N_46638);
xor UO_3538 (O_3538,N_48648,N_49797);
or UO_3539 (O_3539,N_47640,N_46587);
xor UO_3540 (O_3540,N_45434,N_46020);
or UO_3541 (O_3541,N_46503,N_46456);
or UO_3542 (O_3542,N_47450,N_46859);
and UO_3543 (O_3543,N_49510,N_45180);
nand UO_3544 (O_3544,N_49640,N_46790);
xor UO_3545 (O_3545,N_47628,N_49813);
nand UO_3546 (O_3546,N_49289,N_46171);
nand UO_3547 (O_3547,N_46987,N_46285);
or UO_3548 (O_3548,N_49529,N_47128);
or UO_3549 (O_3549,N_46208,N_49494);
nand UO_3550 (O_3550,N_46211,N_47003);
or UO_3551 (O_3551,N_45269,N_46722);
nand UO_3552 (O_3552,N_46469,N_48538);
nand UO_3553 (O_3553,N_45900,N_47591);
xnor UO_3554 (O_3554,N_49473,N_48464);
nand UO_3555 (O_3555,N_45896,N_45652);
xnor UO_3556 (O_3556,N_46666,N_45250);
xnor UO_3557 (O_3557,N_49800,N_49862);
or UO_3558 (O_3558,N_46765,N_49028);
and UO_3559 (O_3559,N_49348,N_49135);
and UO_3560 (O_3560,N_47193,N_47766);
nand UO_3561 (O_3561,N_45278,N_49798);
nand UO_3562 (O_3562,N_48300,N_46825);
nor UO_3563 (O_3563,N_46619,N_49921);
or UO_3564 (O_3564,N_48056,N_47228);
nand UO_3565 (O_3565,N_45527,N_48506);
and UO_3566 (O_3566,N_45630,N_46961);
xor UO_3567 (O_3567,N_48929,N_45993);
and UO_3568 (O_3568,N_46740,N_45664);
nand UO_3569 (O_3569,N_47034,N_47809);
xnor UO_3570 (O_3570,N_46492,N_49402);
xor UO_3571 (O_3571,N_45439,N_48743);
nand UO_3572 (O_3572,N_48601,N_48564);
nor UO_3573 (O_3573,N_48207,N_48383);
xor UO_3574 (O_3574,N_48527,N_45230);
xor UO_3575 (O_3575,N_49244,N_45001);
or UO_3576 (O_3576,N_47711,N_45429);
nand UO_3577 (O_3577,N_48966,N_46220);
or UO_3578 (O_3578,N_45054,N_46519);
nand UO_3579 (O_3579,N_46251,N_46001);
and UO_3580 (O_3580,N_49266,N_48723);
nand UO_3581 (O_3581,N_49010,N_47231);
or UO_3582 (O_3582,N_47315,N_48948);
and UO_3583 (O_3583,N_49833,N_45398);
or UO_3584 (O_3584,N_45408,N_47235);
nand UO_3585 (O_3585,N_46517,N_48523);
and UO_3586 (O_3586,N_49653,N_49577);
nor UO_3587 (O_3587,N_49492,N_46194);
xnor UO_3588 (O_3588,N_48306,N_45055);
and UO_3589 (O_3589,N_47981,N_48289);
xnor UO_3590 (O_3590,N_45359,N_46635);
and UO_3591 (O_3591,N_45462,N_46112);
nand UO_3592 (O_3592,N_46925,N_45571);
or UO_3593 (O_3593,N_46200,N_46170);
xor UO_3594 (O_3594,N_48076,N_48575);
xor UO_3595 (O_3595,N_49095,N_45570);
nand UO_3596 (O_3596,N_48670,N_48722);
or UO_3597 (O_3597,N_46427,N_46135);
or UO_3598 (O_3598,N_49724,N_48771);
nor UO_3599 (O_3599,N_45916,N_47686);
nor UO_3600 (O_3600,N_45192,N_47195);
or UO_3601 (O_3601,N_48777,N_48094);
nand UO_3602 (O_3602,N_49368,N_47465);
nor UO_3603 (O_3603,N_47537,N_49898);
and UO_3604 (O_3604,N_46394,N_49686);
or UO_3605 (O_3605,N_47972,N_49877);
xnor UO_3606 (O_3606,N_49258,N_47781);
and UO_3607 (O_3607,N_48435,N_45958);
and UO_3608 (O_3608,N_46819,N_45499);
nor UO_3609 (O_3609,N_49748,N_46432);
or UO_3610 (O_3610,N_45526,N_49455);
nand UO_3611 (O_3611,N_49391,N_48895);
xnor UO_3612 (O_3612,N_49267,N_49653);
and UO_3613 (O_3613,N_46353,N_49965);
and UO_3614 (O_3614,N_45547,N_49174);
or UO_3615 (O_3615,N_46730,N_49353);
and UO_3616 (O_3616,N_49306,N_49490);
nand UO_3617 (O_3617,N_49013,N_49773);
or UO_3618 (O_3618,N_47718,N_48123);
and UO_3619 (O_3619,N_48348,N_46396);
xor UO_3620 (O_3620,N_47094,N_46991);
nor UO_3621 (O_3621,N_47161,N_48665);
nor UO_3622 (O_3622,N_45522,N_47913);
and UO_3623 (O_3623,N_48675,N_46713);
nor UO_3624 (O_3624,N_49271,N_49441);
nor UO_3625 (O_3625,N_49996,N_48146);
xor UO_3626 (O_3626,N_48837,N_46163);
nor UO_3627 (O_3627,N_45024,N_48920);
xor UO_3628 (O_3628,N_49906,N_46730);
nor UO_3629 (O_3629,N_48832,N_47556);
nor UO_3630 (O_3630,N_45735,N_47782);
xnor UO_3631 (O_3631,N_47911,N_47529);
and UO_3632 (O_3632,N_48064,N_47572);
nand UO_3633 (O_3633,N_47266,N_45574);
nand UO_3634 (O_3634,N_47351,N_45436);
and UO_3635 (O_3635,N_47471,N_46888);
nand UO_3636 (O_3636,N_46526,N_47339);
or UO_3637 (O_3637,N_49640,N_46672);
xnor UO_3638 (O_3638,N_47023,N_46276);
xnor UO_3639 (O_3639,N_45210,N_49461);
xnor UO_3640 (O_3640,N_47265,N_48676);
xnor UO_3641 (O_3641,N_48277,N_49375);
and UO_3642 (O_3642,N_47771,N_47621);
xor UO_3643 (O_3643,N_45256,N_47289);
nor UO_3644 (O_3644,N_46632,N_49373);
or UO_3645 (O_3645,N_49708,N_45064);
or UO_3646 (O_3646,N_48659,N_47286);
and UO_3647 (O_3647,N_49136,N_45352);
xnor UO_3648 (O_3648,N_49266,N_45733);
and UO_3649 (O_3649,N_46354,N_47642);
xnor UO_3650 (O_3650,N_45221,N_48167);
or UO_3651 (O_3651,N_48269,N_47598);
and UO_3652 (O_3652,N_47973,N_45937);
nor UO_3653 (O_3653,N_45894,N_46762);
xor UO_3654 (O_3654,N_49281,N_45358);
or UO_3655 (O_3655,N_48986,N_48122);
nor UO_3656 (O_3656,N_45563,N_47232);
and UO_3657 (O_3657,N_48885,N_45011);
or UO_3658 (O_3658,N_45003,N_48014);
xor UO_3659 (O_3659,N_46047,N_46755);
and UO_3660 (O_3660,N_48684,N_45166);
nand UO_3661 (O_3661,N_48036,N_48423);
nand UO_3662 (O_3662,N_48415,N_48268);
and UO_3663 (O_3663,N_47129,N_48712);
and UO_3664 (O_3664,N_47055,N_49069);
xnor UO_3665 (O_3665,N_45381,N_47176);
nand UO_3666 (O_3666,N_48069,N_46275);
nor UO_3667 (O_3667,N_46712,N_48592);
or UO_3668 (O_3668,N_45378,N_49535);
or UO_3669 (O_3669,N_48390,N_45122);
xnor UO_3670 (O_3670,N_47478,N_48504);
nor UO_3671 (O_3671,N_47419,N_46458);
nand UO_3672 (O_3672,N_47170,N_45600);
or UO_3673 (O_3673,N_47032,N_46909);
xor UO_3674 (O_3674,N_48593,N_46953);
nand UO_3675 (O_3675,N_49141,N_47384);
nor UO_3676 (O_3676,N_48224,N_45767);
or UO_3677 (O_3677,N_48512,N_46338);
nand UO_3678 (O_3678,N_49702,N_45870);
nor UO_3679 (O_3679,N_48650,N_46176);
nor UO_3680 (O_3680,N_49989,N_48936);
or UO_3681 (O_3681,N_48085,N_46633);
and UO_3682 (O_3682,N_47137,N_46272);
and UO_3683 (O_3683,N_47459,N_47269);
nand UO_3684 (O_3684,N_48831,N_45503);
nor UO_3685 (O_3685,N_48588,N_47269);
xnor UO_3686 (O_3686,N_49034,N_49024);
nand UO_3687 (O_3687,N_45620,N_45518);
nor UO_3688 (O_3688,N_47430,N_45615);
and UO_3689 (O_3689,N_47205,N_46021);
xor UO_3690 (O_3690,N_48503,N_48068);
nor UO_3691 (O_3691,N_47535,N_46019);
and UO_3692 (O_3692,N_46572,N_45139);
nand UO_3693 (O_3693,N_49865,N_46180);
nand UO_3694 (O_3694,N_45201,N_49624);
and UO_3695 (O_3695,N_45232,N_46944);
and UO_3696 (O_3696,N_48487,N_49430);
or UO_3697 (O_3697,N_47753,N_49020);
xor UO_3698 (O_3698,N_47800,N_46371);
xor UO_3699 (O_3699,N_46681,N_49583);
nand UO_3700 (O_3700,N_45453,N_46365);
xnor UO_3701 (O_3701,N_45867,N_47702);
or UO_3702 (O_3702,N_46716,N_46744);
xnor UO_3703 (O_3703,N_48003,N_46275);
or UO_3704 (O_3704,N_45194,N_47146);
or UO_3705 (O_3705,N_45114,N_45094);
xnor UO_3706 (O_3706,N_49703,N_49689);
and UO_3707 (O_3707,N_46635,N_47700);
nor UO_3708 (O_3708,N_48087,N_48857);
or UO_3709 (O_3709,N_45953,N_46660);
or UO_3710 (O_3710,N_46959,N_46785);
or UO_3711 (O_3711,N_48321,N_46833);
nor UO_3712 (O_3712,N_46118,N_47831);
xnor UO_3713 (O_3713,N_45175,N_46548);
xnor UO_3714 (O_3714,N_48929,N_46036);
and UO_3715 (O_3715,N_49175,N_45900);
xnor UO_3716 (O_3716,N_48133,N_46293);
and UO_3717 (O_3717,N_48688,N_45914);
or UO_3718 (O_3718,N_48622,N_45870);
and UO_3719 (O_3719,N_47123,N_45520);
and UO_3720 (O_3720,N_46568,N_47188);
xor UO_3721 (O_3721,N_49454,N_47619);
nor UO_3722 (O_3722,N_46863,N_47011);
and UO_3723 (O_3723,N_48355,N_46475);
or UO_3724 (O_3724,N_48917,N_45857);
nor UO_3725 (O_3725,N_49152,N_46127);
nand UO_3726 (O_3726,N_46744,N_49963);
xor UO_3727 (O_3727,N_46432,N_48998);
and UO_3728 (O_3728,N_48260,N_49081);
or UO_3729 (O_3729,N_46844,N_45840);
and UO_3730 (O_3730,N_49512,N_45672);
xor UO_3731 (O_3731,N_49948,N_49100);
nor UO_3732 (O_3732,N_46356,N_45367);
and UO_3733 (O_3733,N_45204,N_46877);
nor UO_3734 (O_3734,N_48082,N_45799);
nand UO_3735 (O_3735,N_45848,N_48331);
or UO_3736 (O_3736,N_47907,N_46091);
or UO_3737 (O_3737,N_46141,N_46452);
nand UO_3738 (O_3738,N_46715,N_48227);
and UO_3739 (O_3739,N_48024,N_47917);
xor UO_3740 (O_3740,N_47535,N_49461);
nand UO_3741 (O_3741,N_47005,N_45161);
nand UO_3742 (O_3742,N_48331,N_47906);
nand UO_3743 (O_3743,N_49803,N_46854);
xor UO_3744 (O_3744,N_45136,N_47531);
nor UO_3745 (O_3745,N_46816,N_47654);
or UO_3746 (O_3746,N_46266,N_49167);
nand UO_3747 (O_3747,N_48302,N_49395);
xor UO_3748 (O_3748,N_49960,N_46017);
xor UO_3749 (O_3749,N_48571,N_46686);
nor UO_3750 (O_3750,N_49700,N_45627);
or UO_3751 (O_3751,N_48899,N_49970);
nand UO_3752 (O_3752,N_48510,N_47610);
nand UO_3753 (O_3753,N_47682,N_47674);
xor UO_3754 (O_3754,N_49010,N_45733);
nand UO_3755 (O_3755,N_45959,N_46983);
or UO_3756 (O_3756,N_47332,N_49069);
xor UO_3757 (O_3757,N_48488,N_48840);
and UO_3758 (O_3758,N_45013,N_47560);
and UO_3759 (O_3759,N_49934,N_47988);
xnor UO_3760 (O_3760,N_48501,N_47426);
or UO_3761 (O_3761,N_45963,N_48106);
or UO_3762 (O_3762,N_45323,N_46230);
nor UO_3763 (O_3763,N_49329,N_46389);
xor UO_3764 (O_3764,N_48699,N_46583);
and UO_3765 (O_3765,N_49900,N_47877);
or UO_3766 (O_3766,N_47659,N_45965);
nor UO_3767 (O_3767,N_46362,N_48323);
nand UO_3768 (O_3768,N_49422,N_49686);
or UO_3769 (O_3769,N_47747,N_47513);
nor UO_3770 (O_3770,N_46067,N_46928);
xnor UO_3771 (O_3771,N_45013,N_49583);
xnor UO_3772 (O_3772,N_49263,N_49127);
nor UO_3773 (O_3773,N_49353,N_47264);
nor UO_3774 (O_3774,N_48852,N_45560);
and UO_3775 (O_3775,N_49939,N_48399);
nand UO_3776 (O_3776,N_48918,N_47766);
nor UO_3777 (O_3777,N_49205,N_45363);
and UO_3778 (O_3778,N_47739,N_45002);
nor UO_3779 (O_3779,N_46670,N_49655);
or UO_3780 (O_3780,N_49565,N_48833);
nor UO_3781 (O_3781,N_49156,N_45726);
nand UO_3782 (O_3782,N_48526,N_49943);
and UO_3783 (O_3783,N_46695,N_47005);
nand UO_3784 (O_3784,N_46772,N_46188);
xnor UO_3785 (O_3785,N_48159,N_45026);
nor UO_3786 (O_3786,N_49168,N_46428);
nand UO_3787 (O_3787,N_46267,N_46235);
xnor UO_3788 (O_3788,N_46849,N_47890);
or UO_3789 (O_3789,N_49068,N_48361);
xor UO_3790 (O_3790,N_46670,N_49464);
and UO_3791 (O_3791,N_49638,N_45818);
nor UO_3792 (O_3792,N_47317,N_45605);
nand UO_3793 (O_3793,N_46518,N_45844);
or UO_3794 (O_3794,N_47051,N_45706);
nor UO_3795 (O_3795,N_46530,N_46785);
or UO_3796 (O_3796,N_47353,N_45023);
xor UO_3797 (O_3797,N_47187,N_48696);
xnor UO_3798 (O_3798,N_46129,N_46977);
nor UO_3799 (O_3799,N_49788,N_49040);
nor UO_3800 (O_3800,N_47035,N_49205);
nor UO_3801 (O_3801,N_49128,N_48422);
xnor UO_3802 (O_3802,N_46031,N_49843);
xnor UO_3803 (O_3803,N_48011,N_49416);
or UO_3804 (O_3804,N_46309,N_49975);
nor UO_3805 (O_3805,N_45321,N_49483);
xnor UO_3806 (O_3806,N_49977,N_48100);
nand UO_3807 (O_3807,N_48789,N_48504);
nor UO_3808 (O_3808,N_47390,N_49018);
and UO_3809 (O_3809,N_45858,N_46269);
nand UO_3810 (O_3810,N_46701,N_46816);
xor UO_3811 (O_3811,N_45190,N_48137);
and UO_3812 (O_3812,N_48985,N_45442);
nand UO_3813 (O_3813,N_47998,N_48630);
and UO_3814 (O_3814,N_45387,N_48424);
and UO_3815 (O_3815,N_46121,N_48472);
nor UO_3816 (O_3816,N_46627,N_49375);
xnor UO_3817 (O_3817,N_46646,N_47198);
nand UO_3818 (O_3818,N_47864,N_48139);
nand UO_3819 (O_3819,N_47604,N_48854);
xnor UO_3820 (O_3820,N_49752,N_45973);
nor UO_3821 (O_3821,N_45681,N_47826);
nor UO_3822 (O_3822,N_45402,N_46268);
or UO_3823 (O_3823,N_47807,N_46122);
or UO_3824 (O_3824,N_46192,N_45461);
nor UO_3825 (O_3825,N_45445,N_48359);
nand UO_3826 (O_3826,N_48441,N_45191);
or UO_3827 (O_3827,N_49467,N_47551);
or UO_3828 (O_3828,N_46459,N_47508);
xor UO_3829 (O_3829,N_45730,N_45629);
xnor UO_3830 (O_3830,N_46207,N_49820);
and UO_3831 (O_3831,N_49980,N_48527);
and UO_3832 (O_3832,N_47157,N_49413);
nor UO_3833 (O_3833,N_48462,N_46896);
or UO_3834 (O_3834,N_46210,N_49568);
and UO_3835 (O_3835,N_45942,N_49120);
nor UO_3836 (O_3836,N_45537,N_45508);
xnor UO_3837 (O_3837,N_49329,N_48260);
nand UO_3838 (O_3838,N_46260,N_48070);
or UO_3839 (O_3839,N_47016,N_49324);
or UO_3840 (O_3840,N_45499,N_45885);
or UO_3841 (O_3841,N_45426,N_45390);
or UO_3842 (O_3842,N_46635,N_45217);
nor UO_3843 (O_3843,N_47891,N_45036);
nand UO_3844 (O_3844,N_48068,N_48439);
nand UO_3845 (O_3845,N_49028,N_45868);
nor UO_3846 (O_3846,N_46680,N_46806);
and UO_3847 (O_3847,N_49130,N_46503);
or UO_3848 (O_3848,N_45299,N_47717);
nand UO_3849 (O_3849,N_47611,N_48623);
or UO_3850 (O_3850,N_46903,N_45948);
nor UO_3851 (O_3851,N_46386,N_46647);
nand UO_3852 (O_3852,N_46891,N_49304);
xor UO_3853 (O_3853,N_45445,N_48451);
nor UO_3854 (O_3854,N_46710,N_45227);
nor UO_3855 (O_3855,N_49101,N_48415);
xnor UO_3856 (O_3856,N_45770,N_48593);
or UO_3857 (O_3857,N_49794,N_45970);
nand UO_3858 (O_3858,N_45012,N_46524);
or UO_3859 (O_3859,N_46212,N_45282);
nand UO_3860 (O_3860,N_47772,N_46905);
xor UO_3861 (O_3861,N_46870,N_46288);
nand UO_3862 (O_3862,N_49628,N_48355);
xnor UO_3863 (O_3863,N_49048,N_45194);
nor UO_3864 (O_3864,N_47981,N_48011);
nor UO_3865 (O_3865,N_47719,N_46110);
nor UO_3866 (O_3866,N_45380,N_46131);
xnor UO_3867 (O_3867,N_45061,N_46203);
nand UO_3868 (O_3868,N_45551,N_48035);
xnor UO_3869 (O_3869,N_47319,N_46579);
nor UO_3870 (O_3870,N_48741,N_46855);
and UO_3871 (O_3871,N_46750,N_48152);
or UO_3872 (O_3872,N_49176,N_48481);
and UO_3873 (O_3873,N_49625,N_46775);
nand UO_3874 (O_3874,N_48261,N_48521);
or UO_3875 (O_3875,N_48949,N_48081);
xor UO_3876 (O_3876,N_47370,N_46777);
nand UO_3877 (O_3877,N_47361,N_49230);
or UO_3878 (O_3878,N_47278,N_45330);
xnor UO_3879 (O_3879,N_47016,N_49322);
and UO_3880 (O_3880,N_48971,N_49080);
and UO_3881 (O_3881,N_47129,N_46639);
or UO_3882 (O_3882,N_47737,N_45794);
xnor UO_3883 (O_3883,N_47806,N_45999);
nor UO_3884 (O_3884,N_47770,N_46815);
xor UO_3885 (O_3885,N_49970,N_48054);
xor UO_3886 (O_3886,N_46170,N_49961);
nand UO_3887 (O_3887,N_48405,N_46495);
nand UO_3888 (O_3888,N_49679,N_49103);
or UO_3889 (O_3889,N_46775,N_47132);
nor UO_3890 (O_3890,N_46442,N_46702);
or UO_3891 (O_3891,N_48971,N_47575);
nor UO_3892 (O_3892,N_47223,N_47954);
and UO_3893 (O_3893,N_45185,N_49002);
nor UO_3894 (O_3894,N_46527,N_46917);
or UO_3895 (O_3895,N_47125,N_46121);
and UO_3896 (O_3896,N_45882,N_46719);
nand UO_3897 (O_3897,N_47398,N_45184);
xor UO_3898 (O_3898,N_49319,N_47466);
xor UO_3899 (O_3899,N_45972,N_47848);
nor UO_3900 (O_3900,N_49307,N_47586);
and UO_3901 (O_3901,N_47389,N_48460);
and UO_3902 (O_3902,N_45522,N_48257);
or UO_3903 (O_3903,N_48138,N_47986);
and UO_3904 (O_3904,N_48609,N_47406);
nand UO_3905 (O_3905,N_45202,N_46569);
nor UO_3906 (O_3906,N_45514,N_47057);
xnor UO_3907 (O_3907,N_45580,N_49831);
nand UO_3908 (O_3908,N_49114,N_45673);
and UO_3909 (O_3909,N_46688,N_45164);
nand UO_3910 (O_3910,N_48751,N_47782);
nand UO_3911 (O_3911,N_48770,N_47664);
or UO_3912 (O_3912,N_49732,N_46304);
nor UO_3913 (O_3913,N_45361,N_48840);
and UO_3914 (O_3914,N_48640,N_48601);
xnor UO_3915 (O_3915,N_47246,N_49616);
nand UO_3916 (O_3916,N_45303,N_46369);
or UO_3917 (O_3917,N_48467,N_46389);
or UO_3918 (O_3918,N_49431,N_49958);
and UO_3919 (O_3919,N_45068,N_48284);
xor UO_3920 (O_3920,N_46416,N_48266);
xor UO_3921 (O_3921,N_47086,N_48652);
or UO_3922 (O_3922,N_46385,N_48659);
nor UO_3923 (O_3923,N_47697,N_49168);
xnor UO_3924 (O_3924,N_48483,N_48167);
and UO_3925 (O_3925,N_49369,N_49147);
nor UO_3926 (O_3926,N_48692,N_46438);
nand UO_3927 (O_3927,N_48873,N_47228);
xor UO_3928 (O_3928,N_45419,N_48215);
nand UO_3929 (O_3929,N_48726,N_48185);
or UO_3930 (O_3930,N_48485,N_48699);
nor UO_3931 (O_3931,N_49193,N_46441);
nor UO_3932 (O_3932,N_47977,N_46931);
or UO_3933 (O_3933,N_47296,N_47442);
nor UO_3934 (O_3934,N_46509,N_47026);
and UO_3935 (O_3935,N_47066,N_46780);
nor UO_3936 (O_3936,N_45484,N_46327);
and UO_3937 (O_3937,N_45574,N_47920);
or UO_3938 (O_3938,N_47123,N_47312);
or UO_3939 (O_3939,N_48066,N_45156);
xor UO_3940 (O_3940,N_45598,N_47962);
nand UO_3941 (O_3941,N_47875,N_47482);
xor UO_3942 (O_3942,N_46954,N_47595);
xnor UO_3943 (O_3943,N_49501,N_45463);
nor UO_3944 (O_3944,N_46588,N_47863);
xnor UO_3945 (O_3945,N_47451,N_45518);
or UO_3946 (O_3946,N_45447,N_49793);
nand UO_3947 (O_3947,N_49290,N_48146);
nand UO_3948 (O_3948,N_47287,N_48860);
and UO_3949 (O_3949,N_49583,N_45835);
nor UO_3950 (O_3950,N_46541,N_49699);
and UO_3951 (O_3951,N_47376,N_48037);
nand UO_3952 (O_3952,N_46229,N_48969);
nor UO_3953 (O_3953,N_48448,N_48888);
or UO_3954 (O_3954,N_49529,N_49444);
and UO_3955 (O_3955,N_46541,N_45775);
nand UO_3956 (O_3956,N_49151,N_46152);
or UO_3957 (O_3957,N_45047,N_49659);
nand UO_3958 (O_3958,N_45088,N_46446);
nand UO_3959 (O_3959,N_46695,N_45247);
xnor UO_3960 (O_3960,N_49173,N_47590);
nand UO_3961 (O_3961,N_45575,N_45868);
or UO_3962 (O_3962,N_45314,N_47255);
xor UO_3963 (O_3963,N_47487,N_48939);
xnor UO_3964 (O_3964,N_48413,N_46896);
nand UO_3965 (O_3965,N_47933,N_46215);
nand UO_3966 (O_3966,N_47781,N_45839);
nand UO_3967 (O_3967,N_46169,N_46922);
nand UO_3968 (O_3968,N_45885,N_49903);
nand UO_3969 (O_3969,N_49048,N_49187);
nor UO_3970 (O_3970,N_46824,N_48578);
or UO_3971 (O_3971,N_47205,N_49598);
and UO_3972 (O_3972,N_47751,N_48035);
xnor UO_3973 (O_3973,N_46316,N_46621);
and UO_3974 (O_3974,N_48872,N_48295);
or UO_3975 (O_3975,N_47218,N_47196);
xnor UO_3976 (O_3976,N_45210,N_48807);
nand UO_3977 (O_3977,N_48098,N_47100);
xor UO_3978 (O_3978,N_48793,N_45185);
nor UO_3979 (O_3979,N_48872,N_48088);
and UO_3980 (O_3980,N_46035,N_45808);
or UO_3981 (O_3981,N_47425,N_48879);
nor UO_3982 (O_3982,N_47409,N_49560);
or UO_3983 (O_3983,N_49956,N_49663);
nand UO_3984 (O_3984,N_47208,N_49565);
or UO_3985 (O_3985,N_47234,N_45814);
and UO_3986 (O_3986,N_45544,N_47560);
nor UO_3987 (O_3987,N_47392,N_47215);
or UO_3988 (O_3988,N_47068,N_48314);
or UO_3989 (O_3989,N_48644,N_45464);
and UO_3990 (O_3990,N_46371,N_47693);
and UO_3991 (O_3991,N_47437,N_47721);
nor UO_3992 (O_3992,N_47197,N_45909);
xnor UO_3993 (O_3993,N_46723,N_49249);
xnor UO_3994 (O_3994,N_46313,N_45274);
nor UO_3995 (O_3995,N_47820,N_46292);
nand UO_3996 (O_3996,N_49679,N_48135);
and UO_3997 (O_3997,N_48535,N_45814);
xor UO_3998 (O_3998,N_48717,N_46025);
xnor UO_3999 (O_3999,N_45118,N_45441);
nor UO_4000 (O_4000,N_45602,N_45007);
and UO_4001 (O_4001,N_48578,N_47194);
nand UO_4002 (O_4002,N_49004,N_46712);
xor UO_4003 (O_4003,N_48634,N_49345);
or UO_4004 (O_4004,N_48431,N_49186);
nand UO_4005 (O_4005,N_47201,N_49382);
and UO_4006 (O_4006,N_48904,N_45500);
nor UO_4007 (O_4007,N_47439,N_46359);
or UO_4008 (O_4008,N_46419,N_48728);
xor UO_4009 (O_4009,N_46954,N_46081);
nor UO_4010 (O_4010,N_45623,N_45981);
nand UO_4011 (O_4011,N_49046,N_45813);
xnor UO_4012 (O_4012,N_48946,N_45033);
or UO_4013 (O_4013,N_47259,N_47029);
or UO_4014 (O_4014,N_49428,N_45724);
or UO_4015 (O_4015,N_47623,N_49463);
and UO_4016 (O_4016,N_46724,N_48848);
or UO_4017 (O_4017,N_47193,N_47286);
or UO_4018 (O_4018,N_45614,N_46810);
xnor UO_4019 (O_4019,N_49056,N_46336);
nor UO_4020 (O_4020,N_46112,N_46297);
or UO_4021 (O_4021,N_46428,N_47506);
nor UO_4022 (O_4022,N_48595,N_48104);
nand UO_4023 (O_4023,N_45141,N_47739);
or UO_4024 (O_4024,N_47315,N_45129);
nor UO_4025 (O_4025,N_47145,N_48863);
or UO_4026 (O_4026,N_47944,N_46610);
xnor UO_4027 (O_4027,N_49083,N_45858);
and UO_4028 (O_4028,N_49143,N_49572);
or UO_4029 (O_4029,N_45966,N_48095);
or UO_4030 (O_4030,N_49830,N_49094);
or UO_4031 (O_4031,N_45214,N_48951);
nand UO_4032 (O_4032,N_47685,N_47450);
xor UO_4033 (O_4033,N_46716,N_46578);
and UO_4034 (O_4034,N_49115,N_47866);
nor UO_4035 (O_4035,N_47202,N_48163);
nor UO_4036 (O_4036,N_46570,N_45760);
and UO_4037 (O_4037,N_45277,N_47349);
or UO_4038 (O_4038,N_47299,N_48578);
xnor UO_4039 (O_4039,N_47550,N_48206);
nand UO_4040 (O_4040,N_45907,N_49712);
nor UO_4041 (O_4041,N_46457,N_45703);
xnor UO_4042 (O_4042,N_47253,N_48760);
and UO_4043 (O_4043,N_48800,N_49024);
xnor UO_4044 (O_4044,N_49383,N_47313);
nor UO_4045 (O_4045,N_47826,N_46215);
or UO_4046 (O_4046,N_46168,N_47907);
or UO_4047 (O_4047,N_46895,N_49034);
nor UO_4048 (O_4048,N_46206,N_46636);
nand UO_4049 (O_4049,N_48540,N_45084);
xor UO_4050 (O_4050,N_48832,N_45877);
nand UO_4051 (O_4051,N_46945,N_48228);
and UO_4052 (O_4052,N_47820,N_49682);
nor UO_4053 (O_4053,N_45489,N_48851);
and UO_4054 (O_4054,N_46475,N_48933);
nand UO_4055 (O_4055,N_46823,N_49449);
nand UO_4056 (O_4056,N_48894,N_49139);
or UO_4057 (O_4057,N_48343,N_46488);
nor UO_4058 (O_4058,N_46282,N_46638);
or UO_4059 (O_4059,N_48642,N_45777);
xor UO_4060 (O_4060,N_46839,N_47759);
nor UO_4061 (O_4061,N_47503,N_49525);
and UO_4062 (O_4062,N_48446,N_46202);
and UO_4063 (O_4063,N_45746,N_47944);
nand UO_4064 (O_4064,N_49363,N_45545);
nand UO_4065 (O_4065,N_46408,N_49481);
or UO_4066 (O_4066,N_49730,N_49360);
nand UO_4067 (O_4067,N_49445,N_45658);
or UO_4068 (O_4068,N_46331,N_47347);
nand UO_4069 (O_4069,N_49840,N_47925);
xor UO_4070 (O_4070,N_45213,N_49946);
nand UO_4071 (O_4071,N_49447,N_45159);
xor UO_4072 (O_4072,N_48054,N_49213);
or UO_4073 (O_4073,N_47214,N_48226);
and UO_4074 (O_4074,N_48194,N_48011);
or UO_4075 (O_4075,N_46769,N_48400);
nand UO_4076 (O_4076,N_45813,N_45495);
xor UO_4077 (O_4077,N_49544,N_46172);
or UO_4078 (O_4078,N_49967,N_48955);
and UO_4079 (O_4079,N_47316,N_49162);
or UO_4080 (O_4080,N_45679,N_46264);
nand UO_4081 (O_4081,N_49765,N_45705);
nand UO_4082 (O_4082,N_48267,N_49235);
or UO_4083 (O_4083,N_47179,N_49575);
or UO_4084 (O_4084,N_49771,N_48194);
or UO_4085 (O_4085,N_49799,N_48210);
nor UO_4086 (O_4086,N_46527,N_48208);
xnor UO_4087 (O_4087,N_45580,N_47035);
nand UO_4088 (O_4088,N_45603,N_49871);
or UO_4089 (O_4089,N_46385,N_48192);
nor UO_4090 (O_4090,N_48062,N_48557);
or UO_4091 (O_4091,N_46139,N_47828);
xnor UO_4092 (O_4092,N_47845,N_46855);
and UO_4093 (O_4093,N_46079,N_45757);
nor UO_4094 (O_4094,N_46149,N_49702);
nor UO_4095 (O_4095,N_46770,N_46583);
nand UO_4096 (O_4096,N_47380,N_45338);
and UO_4097 (O_4097,N_45498,N_48449);
or UO_4098 (O_4098,N_47781,N_45693);
and UO_4099 (O_4099,N_46152,N_46622);
or UO_4100 (O_4100,N_49686,N_49112);
nor UO_4101 (O_4101,N_45812,N_45689);
nor UO_4102 (O_4102,N_46888,N_47122);
nand UO_4103 (O_4103,N_47433,N_49019);
nand UO_4104 (O_4104,N_49672,N_47096);
and UO_4105 (O_4105,N_49637,N_45035);
nand UO_4106 (O_4106,N_49813,N_48321);
nor UO_4107 (O_4107,N_48988,N_48601);
xnor UO_4108 (O_4108,N_49020,N_49489);
and UO_4109 (O_4109,N_46129,N_47833);
nor UO_4110 (O_4110,N_48531,N_45583);
xnor UO_4111 (O_4111,N_48528,N_49653);
xor UO_4112 (O_4112,N_46742,N_45888);
or UO_4113 (O_4113,N_48941,N_46817);
nand UO_4114 (O_4114,N_47558,N_45552);
nand UO_4115 (O_4115,N_49980,N_49907);
or UO_4116 (O_4116,N_49232,N_49971);
and UO_4117 (O_4117,N_49179,N_49920);
nand UO_4118 (O_4118,N_45158,N_47268);
nor UO_4119 (O_4119,N_46997,N_49762);
nor UO_4120 (O_4120,N_47488,N_49467);
nor UO_4121 (O_4121,N_47452,N_46896);
and UO_4122 (O_4122,N_48632,N_48659);
or UO_4123 (O_4123,N_48286,N_45507);
or UO_4124 (O_4124,N_49664,N_47115);
and UO_4125 (O_4125,N_46112,N_46474);
or UO_4126 (O_4126,N_48801,N_45745);
xnor UO_4127 (O_4127,N_46719,N_45393);
nand UO_4128 (O_4128,N_49918,N_46701);
xnor UO_4129 (O_4129,N_47958,N_49710);
nor UO_4130 (O_4130,N_47687,N_49378);
nor UO_4131 (O_4131,N_47063,N_47741);
or UO_4132 (O_4132,N_49725,N_45513);
xnor UO_4133 (O_4133,N_45899,N_45318);
or UO_4134 (O_4134,N_49051,N_45447);
and UO_4135 (O_4135,N_46359,N_47586);
nand UO_4136 (O_4136,N_47243,N_45759);
nand UO_4137 (O_4137,N_48488,N_46635);
nor UO_4138 (O_4138,N_47138,N_48666);
xor UO_4139 (O_4139,N_45317,N_49782);
xnor UO_4140 (O_4140,N_49741,N_47510);
and UO_4141 (O_4141,N_45232,N_49094);
nand UO_4142 (O_4142,N_47891,N_49087);
and UO_4143 (O_4143,N_45060,N_47874);
and UO_4144 (O_4144,N_46930,N_46570);
and UO_4145 (O_4145,N_45171,N_46342);
or UO_4146 (O_4146,N_47519,N_49596);
or UO_4147 (O_4147,N_49337,N_49212);
or UO_4148 (O_4148,N_48962,N_49211);
nand UO_4149 (O_4149,N_45542,N_48857);
xnor UO_4150 (O_4150,N_47251,N_47610);
nor UO_4151 (O_4151,N_46673,N_47756);
xor UO_4152 (O_4152,N_45695,N_49915);
or UO_4153 (O_4153,N_48016,N_45488);
and UO_4154 (O_4154,N_49264,N_48799);
nand UO_4155 (O_4155,N_46356,N_45318);
nor UO_4156 (O_4156,N_48979,N_45641);
or UO_4157 (O_4157,N_46961,N_47188);
xor UO_4158 (O_4158,N_49447,N_49770);
nand UO_4159 (O_4159,N_49205,N_49416);
nand UO_4160 (O_4160,N_47322,N_45044);
and UO_4161 (O_4161,N_47191,N_47771);
nor UO_4162 (O_4162,N_49097,N_46354);
nand UO_4163 (O_4163,N_49833,N_45762);
and UO_4164 (O_4164,N_48647,N_48460);
nand UO_4165 (O_4165,N_47378,N_46468);
xnor UO_4166 (O_4166,N_45867,N_47849);
xor UO_4167 (O_4167,N_48067,N_49025);
or UO_4168 (O_4168,N_46098,N_45688);
and UO_4169 (O_4169,N_49004,N_45968);
xnor UO_4170 (O_4170,N_49624,N_46264);
nor UO_4171 (O_4171,N_46894,N_48440);
nand UO_4172 (O_4172,N_48840,N_49336);
xor UO_4173 (O_4173,N_45382,N_45904);
xor UO_4174 (O_4174,N_45840,N_49687);
xor UO_4175 (O_4175,N_45504,N_49987);
and UO_4176 (O_4176,N_48714,N_45011);
and UO_4177 (O_4177,N_48200,N_49715);
nand UO_4178 (O_4178,N_49284,N_47939);
nand UO_4179 (O_4179,N_48510,N_47326);
xor UO_4180 (O_4180,N_45367,N_45357);
or UO_4181 (O_4181,N_45439,N_46310);
and UO_4182 (O_4182,N_45298,N_46504);
nor UO_4183 (O_4183,N_47931,N_48737);
nor UO_4184 (O_4184,N_46004,N_46103);
xnor UO_4185 (O_4185,N_49274,N_49935);
and UO_4186 (O_4186,N_48950,N_47051);
and UO_4187 (O_4187,N_45083,N_46275);
nor UO_4188 (O_4188,N_45138,N_45089);
nand UO_4189 (O_4189,N_45970,N_47246);
nand UO_4190 (O_4190,N_46264,N_47542);
or UO_4191 (O_4191,N_46569,N_45109);
nand UO_4192 (O_4192,N_47659,N_46208);
nand UO_4193 (O_4193,N_47908,N_47047);
xnor UO_4194 (O_4194,N_48105,N_45406);
and UO_4195 (O_4195,N_46173,N_48818);
or UO_4196 (O_4196,N_49137,N_45274);
xnor UO_4197 (O_4197,N_49371,N_48139);
xnor UO_4198 (O_4198,N_49996,N_48780);
nand UO_4199 (O_4199,N_45418,N_48568);
or UO_4200 (O_4200,N_48224,N_46663);
nor UO_4201 (O_4201,N_45433,N_46903);
nand UO_4202 (O_4202,N_49520,N_45484);
nand UO_4203 (O_4203,N_49626,N_45527);
xor UO_4204 (O_4204,N_46568,N_46917);
nor UO_4205 (O_4205,N_46098,N_45310);
xnor UO_4206 (O_4206,N_48789,N_45607);
xor UO_4207 (O_4207,N_45224,N_46494);
and UO_4208 (O_4208,N_47172,N_48638);
and UO_4209 (O_4209,N_48376,N_48266);
nor UO_4210 (O_4210,N_45407,N_47272);
and UO_4211 (O_4211,N_49076,N_47701);
xor UO_4212 (O_4212,N_46158,N_47811);
xor UO_4213 (O_4213,N_47768,N_49777);
or UO_4214 (O_4214,N_45369,N_47649);
xor UO_4215 (O_4215,N_49795,N_48868);
and UO_4216 (O_4216,N_47493,N_45541);
nand UO_4217 (O_4217,N_47291,N_49294);
nor UO_4218 (O_4218,N_49644,N_47250);
nand UO_4219 (O_4219,N_45699,N_46819);
xnor UO_4220 (O_4220,N_49740,N_49783);
nand UO_4221 (O_4221,N_48177,N_48250);
nor UO_4222 (O_4222,N_47585,N_46284);
nor UO_4223 (O_4223,N_49838,N_47977);
xnor UO_4224 (O_4224,N_49504,N_47305);
or UO_4225 (O_4225,N_45031,N_49029);
xnor UO_4226 (O_4226,N_48887,N_46915);
nor UO_4227 (O_4227,N_49038,N_45172);
xnor UO_4228 (O_4228,N_46815,N_48246);
nor UO_4229 (O_4229,N_45476,N_49572);
nand UO_4230 (O_4230,N_46410,N_45797);
or UO_4231 (O_4231,N_48658,N_49056);
nand UO_4232 (O_4232,N_46419,N_49354);
nor UO_4233 (O_4233,N_45684,N_48573);
xor UO_4234 (O_4234,N_47617,N_49920);
or UO_4235 (O_4235,N_48025,N_49908);
xor UO_4236 (O_4236,N_47445,N_49747);
and UO_4237 (O_4237,N_46008,N_47897);
nand UO_4238 (O_4238,N_45234,N_45655);
or UO_4239 (O_4239,N_45147,N_48516);
nand UO_4240 (O_4240,N_48553,N_45423);
xor UO_4241 (O_4241,N_45646,N_48308);
and UO_4242 (O_4242,N_45235,N_45298);
nor UO_4243 (O_4243,N_47824,N_49606);
nor UO_4244 (O_4244,N_46850,N_47091);
and UO_4245 (O_4245,N_48774,N_45262);
nand UO_4246 (O_4246,N_47615,N_46874);
and UO_4247 (O_4247,N_48894,N_48050);
or UO_4248 (O_4248,N_49266,N_46895);
nor UO_4249 (O_4249,N_49232,N_46602);
or UO_4250 (O_4250,N_46843,N_46669);
xnor UO_4251 (O_4251,N_47528,N_47615);
or UO_4252 (O_4252,N_46345,N_48363);
or UO_4253 (O_4253,N_45450,N_48507);
xor UO_4254 (O_4254,N_45860,N_48722);
and UO_4255 (O_4255,N_48374,N_49921);
xnor UO_4256 (O_4256,N_46348,N_47576);
nor UO_4257 (O_4257,N_49780,N_47449);
or UO_4258 (O_4258,N_48771,N_49905);
nand UO_4259 (O_4259,N_45952,N_49493);
nor UO_4260 (O_4260,N_45218,N_47873);
nor UO_4261 (O_4261,N_49325,N_48657);
or UO_4262 (O_4262,N_46512,N_48662);
and UO_4263 (O_4263,N_47703,N_47631);
xor UO_4264 (O_4264,N_48659,N_46485);
nand UO_4265 (O_4265,N_45156,N_45863);
and UO_4266 (O_4266,N_47002,N_48330);
xor UO_4267 (O_4267,N_47502,N_49887);
nand UO_4268 (O_4268,N_48611,N_48791);
xor UO_4269 (O_4269,N_49982,N_48541);
or UO_4270 (O_4270,N_49575,N_45733);
nand UO_4271 (O_4271,N_46095,N_46974);
nor UO_4272 (O_4272,N_46573,N_48549);
or UO_4273 (O_4273,N_49151,N_49192);
xor UO_4274 (O_4274,N_48227,N_49087);
and UO_4275 (O_4275,N_45728,N_48522);
nand UO_4276 (O_4276,N_46953,N_47514);
xor UO_4277 (O_4277,N_46117,N_46754);
or UO_4278 (O_4278,N_47790,N_47667);
and UO_4279 (O_4279,N_47483,N_49104);
xor UO_4280 (O_4280,N_49713,N_46118);
nand UO_4281 (O_4281,N_46828,N_45291);
and UO_4282 (O_4282,N_47292,N_47457);
nor UO_4283 (O_4283,N_48686,N_48082);
or UO_4284 (O_4284,N_48780,N_49764);
and UO_4285 (O_4285,N_48499,N_48602);
or UO_4286 (O_4286,N_45357,N_48040);
or UO_4287 (O_4287,N_45773,N_49239);
nand UO_4288 (O_4288,N_49194,N_49861);
and UO_4289 (O_4289,N_49042,N_49488);
nor UO_4290 (O_4290,N_48544,N_49093);
nor UO_4291 (O_4291,N_47042,N_48330);
nor UO_4292 (O_4292,N_49706,N_46513);
nor UO_4293 (O_4293,N_45624,N_49190);
nand UO_4294 (O_4294,N_46858,N_48959);
or UO_4295 (O_4295,N_48925,N_48536);
nand UO_4296 (O_4296,N_48109,N_47727);
xnor UO_4297 (O_4297,N_48564,N_45724);
or UO_4298 (O_4298,N_45393,N_45513);
xor UO_4299 (O_4299,N_49178,N_49963);
and UO_4300 (O_4300,N_49797,N_46894);
or UO_4301 (O_4301,N_45318,N_47823);
or UO_4302 (O_4302,N_46620,N_46934);
and UO_4303 (O_4303,N_48470,N_49757);
and UO_4304 (O_4304,N_49959,N_47904);
nor UO_4305 (O_4305,N_45426,N_48593);
or UO_4306 (O_4306,N_47388,N_46033);
xor UO_4307 (O_4307,N_46783,N_46044);
and UO_4308 (O_4308,N_48711,N_45122);
nand UO_4309 (O_4309,N_46503,N_48833);
and UO_4310 (O_4310,N_47689,N_47646);
or UO_4311 (O_4311,N_45484,N_47883);
nor UO_4312 (O_4312,N_49140,N_48305);
or UO_4313 (O_4313,N_45835,N_49442);
or UO_4314 (O_4314,N_45556,N_46376);
and UO_4315 (O_4315,N_45477,N_47522);
nand UO_4316 (O_4316,N_46781,N_45812);
nor UO_4317 (O_4317,N_45205,N_45034);
and UO_4318 (O_4318,N_46018,N_49890);
or UO_4319 (O_4319,N_48725,N_46495);
xnor UO_4320 (O_4320,N_48105,N_48468);
and UO_4321 (O_4321,N_47645,N_49202);
or UO_4322 (O_4322,N_46510,N_49841);
nand UO_4323 (O_4323,N_49245,N_45515);
nand UO_4324 (O_4324,N_45198,N_49104);
nand UO_4325 (O_4325,N_45928,N_46139);
and UO_4326 (O_4326,N_45680,N_48040);
xor UO_4327 (O_4327,N_46960,N_48835);
and UO_4328 (O_4328,N_45684,N_45031);
xnor UO_4329 (O_4329,N_46517,N_46496);
and UO_4330 (O_4330,N_46235,N_48190);
nor UO_4331 (O_4331,N_49855,N_46668);
or UO_4332 (O_4332,N_45975,N_48360);
xor UO_4333 (O_4333,N_47097,N_47399);
or UO_4334 (O_4334,N_48968,N_46214);
nand UO_4335 (O_4335,N_49766,N_49456);
nand UO_4336 (O_4336,N_46485,N_49007);
or UO_4337 (O_4337,N_46802,N_48847);
xor UO_4338 (O_4338,N_49659,N_45832);
nand UO_4339 (O_4339,N_49755,N_47862);
xor UO_4340 (O_4340,N_47780,N_48092);
xor UO_4341 (O_4341,N_48176,N_48189);
nand UO_4342 (O_4342,N_47175,N_48256);
xor UO_4343 (O_4343,N_46852,N_47399);
xnor UO_4344 (O_4344,N_47992,N_46233);
xnor UO_4345 (O_4345,N_48452,N_47003);
or UO_4346 (O_4346,N_46730,N_48234);
nand UO_4347 (O_4347,N_48973,N_49691);
or UO_4348 (O_4348,N_46467,N_45198);
or UO_4349 (O_4349,N_47374,N_48805);
nand UO_4350 (O_4350,N_48739,N_49244);
nor UO_4351 (O_4351,N_49768,N_45659);
and UO_4352 (O_4352,N_48578,N_47333);
nor UO_4353 (O_4353,N_48404,N_46060);
or UO_4354 (O_4354,N_48595,N_46773);
and UO_4355 (O_4355,N_47700,N_45183);
nand UO_4356 (O_4356,N_49015,N_45365);
xor UO_4357 (O_4357,N_49331,N_49355);
and UO_4358 (O_4358,N_45701,N_45751);
xor UO_4359 (O_4359,N_47429,N_47707);
nand UO_4360 (O_4360,N_46204,N_47129);
nor UO_4361 (O_4361,N_49529,N_46263);
nor UO_4362 (O_4362,N_48334,N_48430);
nand UO_4363 (O_4363,N_48859,N_49885);
or UO_4364 (O_4364,N_45718,N_45135);
xnor UO_4365 (O_4365,N_47096,N_48124);
or UO_4366 (O_4366,N_48566,N_48542);
and UO_4367 (O_4367,N_47470,N_48814);
or UO_4368 (O_4368,N_45647,N_46367);
nor UO_4369 (O_4369,N_47232,N_49936);
xnor UO_4370 (O_4370,N_49101,N_49801);
and UO_4371 (O_4371,N_47430,N_49803);
nand UO_4372 (O_4372,N_47139,N_45546);
nor UO_4373 (O_4373,N_47731,N_47049);
xor UO_4374 (O_4374,N_46131,N_45227);
nand UO_4375 (O_4375,N_45465,N_47998);
xnor UO_4376 (O_4376,N_45054,N_47979);
nor UO_4377 (O_4377,N_49742,N_45028);
and UO_4378 (O_4378,N_47582,N_48259);
and UO_4379 (O_4379,N_48645,N_48223);
xor UO_4380 (O_4380,N_45288,N_48519);
or UO_4381 (O_4381,N_47782,N_47008);
xnor UO_4382 (O_4382,N_48589,N_49084);
nor UO_4383 (O_4383,N_49501,N_45030);
xor UO_4384 (O_4384,N_45598,N_48846);
xnor UO_4385 (O_4385,N_45098,N_46899);
or UO_4386 (O_4386,N_48756,N_47434);
or UO_4387 (O_4387,N_47338,N_48342);
xor UO_4388 (O_4388,N_49170,N_48913);
xnor UO_4389 (O_4389,N_48460,N_45273);
nor UO_4390 (O_4390,N_45672,N_46065);
nor UO_4391 (O_4391,N_48392,N_47235);
nand UO_4392 (O_4392,N_46961,N_49109);
nor UO_4393 (O_4393,N_48010,N_49920);
nor UO_4394 (O_4394,N_47191,N_47708);
xnor UO_4395 (O_4395,N_46858,N_45079);
xnor UO_4396 (O_4396,N_47531,N_45296);
nor UO_4397 (O_4397,N_47341,N_47267);
xor UO_4398 (O_4398,N_48755,N_46815);
nand UO_4399 (O_4399,N_48495,N_46806);
or UO_4400 (O_4400,N_48828,N_47572);
nand UO_4401 (O_4401,N_47401,N_47694);
nand UO_4402 (O_4402,N_47780,N_46133);
nor UO_4403 (O_4403,N_49221,N_49086);
nand UO_4404 (O_4404,N_48311,N_45327);
nand UO_4405 (O_4405,N_48564,N_47067);
and UO_4406 (O_4406,N_48558,N_48210);
nor UO_4407 (O_4407,N_46752,N_48867);
nor UO_4408 (O_4408,N_48836,N_45022);
nand UO_4409 (O_4409,N_49188,N_45054);
or UO_4410 (O_4410,N_46120,N_48735);
and UO_4411 (O_4411,N_45264,N_46376);
xnor UO_4412 (O_4412,N_45530,N_49196);
or UO_4413 (O_4413,N_48586,N_49728);
or UO_4414 (O_4414,N_49495,N_46119);
and UO_4415 (O_4415,N_47163,N_46885);
xnor UO_4416 (O_4416,N_49941,N_47383);
nand UO_4417 (O_4417,N_47001,N_47178);
and UO_4418 (O_4418,N_49264,N_46450);
nor UO_4419 (O_4419,N_48019,N_46393);
or UO_4420 (O_4420,N_48342,N_49805);
xor UO_4421 (O_4421,N_46984,N_49352);
xor UO_4422 (O_4422,N_47621,N_47958);
nand UO_4423 (O_4423,N_47258,N_46680);
and UO_4424 (O_4424,N_46288,N_46701);
nor UO_4425 (O_4425,N_48527,N_46266);
and UO_4426 (O_4426,N_47356,N_48751);
and UO_4427 (O_4427,N_45931,N_48213);
nand UO_4428 (O_4428,N_45815,N_45479);
xor UO_4429 (O_4429,N_45295,N_48858);
or UO_4430 (O_4430,N_49533,N_46530);
or UO_4431 (O_4431,N_47396,N_49644);
nand UO_4432 (O_4432,N_48460,N_49724);
nor UO_4433 (O_4433,N_47749,N_45583);
and UO_4434 (O_4434,N_45337,N_45476);
xnor UO_4435 (O_4435,N_49047,N_47437);
xor UO_4436 (O_4436,N_47656,N_47068);
nor UO_4437 (O_4437,N_45982,N_49479);
nand UO_4438 (O_4438,N_47083,N_48871);
or UO_4439 (O_4439,N_48658,N_45191);
nor UO_4440 (O_4440,N_47180,N_48683);
nor UO_4441 (O_4441,N_46450,N_49535);
or UO_4442 (O_4442,N_49139,N_49841);
nand UO_4443 (O_4443,N_47135,N_46441);
nor UO_4444 (O_4444,N_49206,N_46782);
xnor UO_4445 (O_4445,N_45224,N_46152);
or UO_4446 (O_4446,N_46092,N_46175);
or UO_4447 (O_4447,N_46168,N_45343);
and UO_4448 (O_4448,N_45659,N_45711);
nand UO_4449 (O_4449,N_47486,N_49510);
and UO_4450 (O_4450,N_46772,N_48449);
and UO_4451 (O_4451,N_49054,N_47897);
or UO_4452 (O_4452,N_47369,N_45296);
nand UO_4453 (O_4453,N_48318,N_49338);
or UO_4454 (O_4454,N_47646,N_47433);
or UO_4455 (O_4455,N_46503,N_49392);
and UO_4456 (O_4456,N_49983,N_45526);
xnor UO_4457 (O_4457,N_46585,N_49200);
or UO_4458 (O_4458,N_47640,N_46452);
and UO_4459 (O_4459,N_47093,N_48397);
or UO_4460 (O_4460,N_45780,N_46929);
xor UO_4461 (O_4461,N_49028,N_49538);
xor UO_4462 (O_4462,N_49484,N_45521);
nand UO_4463 (O_4463,N_48277,N_47412);
and UO_4464 (O_4464,N_48771,N_45322);
nor UO_4465 (O_4465,N_49121,N_46386);
or UO_4466 (O_4466,N_49188,N_49777);
or UO_4467 (O_4467,N_46660,N_46451);
nand UO_4468 (O_4468,N_47664,N_46335);
and UO_4469 (O_4469,N_47443,N_45766);
nand UO_4470 (O_4470,N_49984,N_46297);
xnor UO_4471 (O_4471,N_46375,N_45023);
nor UO_4472 (O_4472,N_47078,N_48465);
xor UO_4473 (O_4473,N_48268,N_48155);
or UO_4474 (O_4474,N_46955,N_45222);
nor UO_4475 (O_4475,N_45951,N_46103);
xnor UO_4476 (O_4476,N_45118,N_45335);
xnor UO_4477 (O_4477,N_45764,N_48035);
xor UO_4478 (O_4478,N_49939,N_48238);
nor UO_4479 (O_4479,N_46885,N_48933);
or UO_4480 (O_4480,N_49068,N_48760);
and UO_4481 (O_4481,N_48214,N_46142);
or UO_4482 (O_4482,N_49325,N_45286);
nor UO_4483 (O_4483,N_45286,N_47684);
and UO_4484 (O_4484,N_46041,N_48464);
or UO_4485 (O_4485,N_46498,N_46781);
nor UO_4486 (O_4486,N_48608,N_49781);
xor UO_4487 (O_4487,N_49875,N_48037);
xnor UO_4488 (O_4488,N_46652,N_45228);
nor UO_4489 (O_4489,N_46523,N_49702);
or UO_4490 (O_4490,N_49593,N_48909);
xor UO_4491 (O_4491,N_49533,N_47198);
nor UO_4492 (O_4492,N_45594,N_48238);
nor UO_4493 (O_4493,N_47602,N_46645);
xnor UO_4494 (O_4494,N_47057,N_47687);
nor UO_4495 (O_4495,N_49544,N_47088);
and UO_4496 (O_4496,N_48419,N_46715);
or UO_4497 (O_4497,N_48097,N_48815);
xnor UO_4498 (O_4498,N_49950,N_45965);
nor UO_4499 (O_4499,N_48821,N_46536);
nor UO_4500 (O_4500,N_45773,N_47532);
nor UO_4501 (O_4501,N_47125,N_49185);
xnor UO_4502 (O_4502,N_45424,N_46095);
or UO_4503 (O_4503,N_45167,N_47097);
nand UO_4504 (O_4504,N_45250,N_49557);
xor UO_4505 (O_4505,N_48564,N_47850);
and UO_4506 (O_4506,N_45157,N_46343);
or UO_4507 (O_4507,N_48988,N_49520);
or UO_4508 (O_4508,N_48189,N_45566);
nand UO_4509 (O_4509,N_45906,N_48595);
or UO_4510 (O_4510,N_46078,N_49178);
or UO_4511 (O_4511,N_48697,N_45276);
nor UO_4512 (O_4512,N_49862,N_49637);
nor UO_4513 (O_4513,N_45460,N_47370);
nand UO_4514 (O_4514,N_45377,N_49776);
nor UO_4515 (O_4515,N_48031,N_46222);
xnor UO_4516 (O_4516,N_49850,N_45967);
or UO_4517 (O_4517,N_47225,N_47356);
nor UO_4518 (O_4518,N_46326,N_48191);
and UO_4519 (O_4519,N_48380,N_45020);
nor UO_4520 (O_4520,N_48539,N_47396);
or UO_4521 (O_4521,N_47343,N_47175);
or UO_4522 (O_4522,N_49321,N_48570);
or UO_4523 (O_4523,N_47564,N_46527);
and UO_4524 (O_4524,N_49012,N_45003);
and UO_4525 (O_4525,N_47636,N_49772);
or UO_4526 (O_4526,N_48680,N_49162);
nand UO_4527 (O_4527,N_45867,N_46832);
or UO_4528 (O_4528,N_49841,N_48780);
and UO_4529 (O_4529,N_45954,N_47661);
or UO_4530 (O_4530,N_46110,N_47283);
and UO_4531 (O_4531,N_47767,N_49589);
or UO_4532 (O_4532,N_47964,N_45468);
nand UO_4533 (O_4533,N_46486,N_46406);
or UO_4534 (O_4534,N_48466,N_49259);
or UO_4535 (O_4535,N_45199,N_46657);
or UO_4536 (O_4536,N_45032,N_49856);
xnor UO_4537 (O_4537,N_47477,N_45436);
and UO_4538 (O_4538,N_47605,N_47869);
nor UO_4539 (O_4539,N_49036,N_47988);
nand UO_4540 (O_4540,N_45791,N_45553);
and UO_4541 (O_4541,N_46833,N_45312);
xnor UO_4542 (O_4542,N_49168,N_46847);
and UO_4543 (O_4543,N_45046,N_47540);
xor UO_4544 (O_4544,N_49987,N_47982);
nand UO_4545 (O_4545,N_47927,N_45427);
and UO_4546 (O_4546,N_46012,N_46593);
xor UO_4547 (O_4547,N_49109,N_49391);
nor UO_4548 (O_4548,N_47200,N_49073);
and UO_4549 (O_4549,N_49176,N_49337);
nand UO_4550 (O_4550,N_45252,N_49568);
or UO_4551 (O_4551,N_47832,N_48598);
nor UO_4552 (O_4552,N_47027,N_48554);
and UO_4553 (O_4553,N_49377,N_49351);
nand UO_4554 (O_4554,N_48107,N_49580);
nor UO_4555 (O_4555,N_48448,N_49116);
and UO_4556 (O_4556,N_46336,N_46769);
or UO_4557 (O_4557,N_45043,N_49412);
xor UO_4558 (O_4558,N_47242,N_46265);
xnor UO_4559 (O_4559,N_45151,N_48443);
and UO_4560 (O_4560,N_48981,N_49072);
and UO_4561 (O_4561,N_45488,N_47544);
nor UO_4562 (O_4562,N_46046,N_45654);
or UO_4563 (O_4563,N_48175,N_45622);
xor UO_4564 (O_4564,N_49362,N_49352);
xnor UO_4565 (O_4565,N_49780,N_46841);
or UO_4566 (O_4566,N_45008,N_48527);
xor UO_4567 (O_4567,N_47056,N_46195);
nand UO_4568 (O_4568,N_48920,N_45879);
or UO_4569 (O_4569,N_46806,N_46261);
or UO_4570 (O_4570,N_47724,N_45935);
or UO_4571 (O_4571,N_48454,N_45235);
nand UO_4572 (O_4572,N_45204,N_49849);
and UO_4573 (O_4573,N_45545,N_49217);
and UO_4574 (O_4574,N_47288,N_46672);
xnor UO_4575 (O_4575,N_46964,N_47222);
or UO_4576 (O_4576,N_49981,N_49093);
xnor UO_4577 (O_4577,N_45042,N_49288);
and UO_4578 (O_4578,N_47375,N_46910);
or UO_4579 (O_4579,N_45546,N_46850);
nor UO_4580 (O_4580,N_46815,N_47073);
nand UO_4581 (O_4581,N_47540,N_46583);
xor UO_4582 (O_4582,N_48476,N_49135);
xor UO_4583 (O_4583,N_48300,N_49592);
nand UO_4584 (O_4584,N_49056,N_45925);
and UO_4585 (O_4585,N_46657,N_47042);
or UO_4586 (O_4586,N_45821,N_49994);
or UO_4587 (O_4587,N_48185,N_47692);
nand UO_4588 (O_4588,N_49355,N_46006);
xor UO_4589 (O_4589,N_47896,N_48358);
nor UO_4590 (O_4590,N_46084,N_45154);
nor UO_4591 (O_4591,N_47900,N_46345);
nand UO_4592 (O_4592,N_49757,N_48363);
nor UO_4593 (O_4593,N_45751,N_48992);
and UO_4594 (O_4594,N_45050,N_48860);
nand UO_4595 (O_4595,N_48175,N_45960);
and UO_4596 (O_4596,N_47591,N_46732);
nand UO_4597 (O_4597,N_47136,N_47713);
xnor UO_4598 (O_4598,N_48213,N_46693);
and UO_4599 (O_4599,N_48267,N_46116);
nor UO_4600 (O_4600,N_49228,N_47249);
xnor UO_4601 (O_4601,N_46350,N_49037);
nand UO_4602 (O_4602,N_46779,N_49996);
nand UO_4603 (O_4603,N_48116,N_49572);
xor UO_4604 (O_4604,N_48160,N_47029);
and UO_4605 (O_4605,N_46110,N_49620);
nand UO_4606 (O_4606,N_46758,N_46587);
nand UO_4607 (O_4607,N_45770,N_49768);
or UO_4608 (O_4608,N_49261,N_48023);
and UO_4609 (O_4609,N_46670,N_49816);
and UO_4610 (O_4610,N_46499,N_48240);
nand UO_4611 (O_4611,N_47348,N_49241);
nor UO_4612 (O_4612,N_47446,N_46982);
and UO_4613 (O_4613,N_46718,N_46223);
and UO_4614 (O_4614,N_48180,N_48368);
or UO_4615 (O_4615,N_46506,N_46860);
and UO_4616 (O_4616,N_49583,N_47223);
nand UO_4617 (O_4617,N_49507,N_48054);
nor UO_4618 (O_4618,N_47892,N_47640);
or UO_4619 (O_4619,N_46211,N_47213);
xnor UO_4620 (O_4620,N_46333,N_48371);
nor UO_4621 (O_4621,N_48311,N_49189);
nor UO_4622 (O_4622,N_45591,N_47727);
nand UO_4623 (O_4623,N_48121,N_49120);
xnor UO_4624 (O_4624,N_46734,N_49341);
xnor UO_4625 (O_4625,N_45691,N_48843);
xor UO_4626 (O_4626,N_49659,N_46777);
xor UO_4627 (O_4627,N_48965,N_49646);
xor UO_4628 (O_4628,N_48654,N_48186);
and UO_4629 (O_4629,N_47017,N_48293);
nand UO_4630 (O_4630,N_45776,N_46382);
and UO_4631 (O_4631,N_45603,N_47484);
nand UO_4632 (O_4632,N_48641,N_47426);
nand UO_4633 (O_4633,N_46221,N_47266);
and UO_4634 (O_4634,N_49283,N_46896);
nor UO_4635 (O_4635,N_45042,N_49464);
nand UO_4636 (O_4636,N_46657,N_49619);
nand UO_4637 (O_4637,N_48355,N_48759);
nand UO_4638 (O_4638,N_48366,N_45335);
or UO_4639 (O_4639,N_48687,N_48561);
xor UO_4640 (O_4640,N_48691,N_48903);
nor UO_4641 (O_4641,N_46204,N_46441);
xnor UO_4642 (O_4642,N_49367,N_49479);
xnor UO_4643 (O_4643,N_47821,N_47725);
nand UO_4644 (O_4644,N_48591,N_45241);
nor UO_4645 (O_4645,N_47785,N_47246);
and UO_4646 (O_4646,N_49147,N_48808);
or UO_4647 (O_4647,N_45376,N_46831);
nand UO_4648 (O_4648,N_45865,N_47411);
and UO_4649 (O_4649,N_46219,N_49871);
and UO_4650 (O_4650,N_47462,N_47186);
nand UO_4651 (O_4651,N_48415,N_49376);
and UO_4652 (O_4652,N_48846,N_46607);
nand UO_4653 (O_4653,N_47635,N_48112);
xnor UO_4654 (O_4654,N_49887,N_45692);
and UO_4655 (O_4655,N_47722,N_47261);
xnor UO_4656 (O_4656,N_49745,N_46940);
xnor UO_4657 (O_4657,N_46788,N_49131);
and UO_4658 (O_4658,N_48764,N_46112);
nand UO_4659 (O_4659,N_45535,N_49622);
or UO_4660 (O_4660,N_49720,N_47948);
or UO_4661 (O_4661,N_46829,N_45256);
and UO_4662 (O_4662,N_49193,N_46258);
or UO_4663 (O_4663,N_48407,N_48609);
nor UO_4664 (O_4664,N_48688,N_48704);
xor UO_4665 (O_4665,N_48771,N_48762);
or UO_4666 (O_4666,N_46516,N_48219);
xnor UO_4667 (O_4667,N_47301,N_46331);
nor UO_4668 (O_4668,N_47398,N_45603);
and UO_4669 (O_4669,N_49892,N_47736);
or UO_4670 (O_4670,N_47447,N_49999);
and UO_4671 (O_4671,N_48718,N_46146);
nor UO_4672 (O_4672,N_47210,N_45364);
nand UO_4673 (O_4673,N_47012,N_48068);
xnor UO_4674 (O_4674,N_47233,N_46964);
and UO_4675 (O_4675,N_48393,N_47143);
nand UO_4676 (O_4676,N_46682,N_46496);
nor UO_4677 (O_4677,N_46996,N_49302);
or UO_4678 (O_4678,N_49701,N_48059);
xnor UO_4679 (O_4679,N_48469,N_49712);
nand UO_4680 (O_4680,N_45718,N_45750);
xnor UO_4681 (O_4681,N_46718,N_49640);
or UO_4682 (O_4682,N_49793,N_48215);
nand UO_4683 (O_4683,N_48334,N_48346);
xnor UO_4684 (O_4684,N_45714,N_48288);
nor UO_4685 (O_4685,N_46813,N_45366);
or UO_4686 (O_4686,N_49651,N_48286);
or UO_4687 (O_4687,N_45513,N_49258);
and UO_4688 (O_4688,N_48462,N_49502);
and UO_4689 (O_4689,N_45120,N_45396);
nor UO_4690 (O_4690,N_49980,N_48491);
nand UO_4691 (O_4691,N_48940,N_45663);
xor UO_4692 (O_4692,N_46078,N_48851);
xnor UO_4693 (O_4693,N_45131,N_49621);
or UO_4694 (O_4694,N_46819,N_49146);
xnor UO_4695 (O_4695,N_46111,N_48965);
nor UO_4696 (O_4696,N_49339,N_48385);
xnor UO_4697 (O_4697,N_46130,N_48099);
nand UO_4698 (O_4698,N_47711,N_47135);
xnor UO_4699 (O_4699,N_48065,N_45536);
nand UO_4700 (O_4700,N_47959,N_48228);
nor UO_4701 (O_4701,N_48142,N_49997);
nand UO_4702 (O_4702,N_49776,N_49672);
nand UO_4703 (O_4703,N_49074,N_49051);
or UO_4704 (O_4704,N_49032,N_46268);
xnor UO_4705 (O_4705,N_48973,N_46609);
nor UO_4706 (O_4706,N_47436,N_48778);
nand UO_4707 (O_4707,N_46039,N_47214);
nor UO_4708 (O_4708,N_46740,N_46687);
nand UO_4709 (O_4709,N_46635,N_47910);
nand UO_4710 (O_4710,N_49399,N_46242);
nor UO_4711 (O_4711,N_49696,N_45983);
nand UO_4712 (O_4712,N_46676,N_49139);
nor UO_4713 (O_4713,N_49147,N_45094);
nand UO_4714 (O_4714,N_48210,N_48437);
xnor UO_4715 (O_4715,N_47928,N_49709);
and UO_4716 (O_4716,N_45869,N_45179);
nand UO_4717 (O_4717,N_47684,N_47585);
and UO_4718 (O_4718,N_48047,N_49219);
and UO_4719 (O_4719,N_48494,N_49195);
nor UO_4720 (O_4720,N_47226,N_49837);
or UO_4721 (O_4721,N_47492,N_49593);
xnor UO_4722 (O_4722,N_47959,N_49766);
or UO_4723 (O_4723,N_45245,N_46932);
xor UO_4724 (O_4724,N_47239,N_49624);
or UO_4725 (O_4725,N_49793,N_45720);
and UO_4726 (O_4726,N_49078,N_46265);
nand UO_4727 (O_4727,N_46404,N_46549);
nand UO_4728 (O_4728,N_47778,N_45292);
or UO_4729 (O_4729,N_48130,N_49722);
nor UO_4730 (O_4730,N_46881,N_46485);
and UO_4731 (O_4731,N_49735,N_47847);
nand UO_4732 (O_4732,N_49988,N_45381);
or UO_4733 (O_4733,N_45845,N_45313);
xor UO_4734 (O_4734,N_46882,N_48744);
xor UO_4735 (O_4735,N_47230,N_47092);
xor UO_4736 (O_4736,N_47469,N_49426);
xnor UO_4737 (O_4737,N_49814,N_45679);
or UO_4738 (O_4738,N_47185,N_48992);
nand UO_4739 (O_4739,N_47483,N_48796);
or UO_4740 (O_4740,N_49698,N_49568);
nor UO_4741 (O_4741,N_46462,N_48667);
nor UO_4742 (O_4742,N_46165,N_47870);
and UO_4743 (O_4743,N_49695,N_45647);
xor UO_4744 (O_4744,N_49324,N_46802);
nor UO_4745 (O_4745,N_48121,N_47622);
xnor UO_4746 (O_4746,N_48919,N_48920);
xor UO_4747 (O_4747,N_48503,N_46975);
xor UO_4748 (O_4748,N_47719,N_45180);
nand UO_4749 (O_4749,N_46968,N_48572);
and UO_4750 (O_4750,N_49265,N_47815);
nor UO_4751 (O_4751,N_48517,N_46811);
and UO_4752 (O_4752,N_48269,N_48853);
nand UO_4753 (O_4753,N_47455,N_49447);
nor UO_4754 (O_4754,N_46188,N_49002);
nor UO_4755 (O_4755,N_49418,N_46092);
nor UO_4756 (O_4756,N_48756,N_47698);
nor UO_4757 (O_4757,N_47155,N_47064);
xor UO_4758 (O_4758,N_45793,N_49971);
nor UO_4759 (O_4759,N_48993,N_49442);
nor UO_4760 (O_4760,N_49205,N_48070);
xor UO_4761 (O_4761,N_46955,N_47549);
or UO_4762 (O_4762,N_49725,N_46985);
nand UO_4763 (O_4763,N_47154,N_48542);
nand UO_4764 (O_4764,N_48100,N_45170);
or UO_4765 (O_4765,N_49943,N_45250);
nand UO_4766 (O_4766,N_48377,N_47066);
or UO_4767 (O_4767,N_47806,N_46047);
and UO_4768 (O_4768,N_48108,N_49319);
nor UO_4769 (O_4769,N_49404,N_49162);
nor UO_4770 (O_4770,N_48025,N_48685);
nor UO_4771 (O_4771,N_49164,N_45435);
and UO_4772 (O_4772,N_49698,N_49091);
nand UO_4773 (O_4773,N_47527,N_45218);
nor UO_4774 (O_4774,N_45321,N_46267);
or UO_4775 (O_4775,N_47794,N_45610);
xor UO_4776 (O_4776,N_46234,N_45294);
and UO_4777 (O_4777,N_49986,N_49502);
nor UO_4778 (O_4778,N_45022,N_45559);
nor UO_4779 (O_4779,N_49330,N_49055);
xnor UO_4780 (O_4780,N_49595,N_46087);
or UO_4781 (O_4781,N_45901,N_47997);
nand UO_4782 (O_4782,N_48267,N_47613);
or UO_4783 (O_4783,N_46755,N_47350);
and UO_4784 (O_4784,N_46630,N_49441);
nor UO_4785 (O_4785,N_47436,N_49974);
xor UO_4786 (O_4786,N_49202,N_49973);
nor UO_4787 (O_4787,N_49216,N_47366);
and UO_4788 (O_4788,N_45035,N_47612);
or UO_4789 (O_4789,N_45735,N_47633);
or UO_4790 (O_4790,N_48611,N_45207);
or UO_4791 (O_4791,N_45215,N_45383);
xor UO_4792 (O_4792,N_46236,N_47292);
or UO_4793 (O_4793,N_46925,N_46994);
nand UO_4794 (O_4794,N_46934,N_46713);
and UO_4795 (O_4795,N_45505,N_45163);
and UO_4796 (O_4796,N_47425,N_46633);
and UO_4797 (O_4797,N_46501,N_49884);
xor UO_4798 (O_4798,N_47513,N_49725);
xor UO_4799 (O_4799,N_48832,N_47275);
xnor UO_4800 (O_4800,N_45048,N_46071);
nand UO_4801 (O_4801,N_46917,N_47892);
xnor UO_4802 (O_4802,N_48831,N_49920);
xor UO_4803 (O_4803,N_45026,N_49682);
xor UO_4804 (O_4804,N_47763,N_46357);
nand UO_4805 (O_4805,N_47270,N_45561);
and UO_4806 (O_4806,N_48574,N_47271);
and UO_4807 (O_4807,N_48955,N_48978);
or UO_4808 (O_4808,N_46867,N_45522);
or UO_4809 (O_4809,N_48985,N_49156);
and UO_4810 (O_4810,N_48120,N_47712);
nor UO_4811 (O_4811,N_49074,N_47519);
nor UO_4812 (O_4812,N_45563,N_45937);
xnor UO_4813 (O_4813,N_49591,N_49199);
and UO_4814 (O_4814,N_49078,N_48550);
and UO_4815 (O_4815,N_45876,N_46192);
nor UO_4816 (O_4816,N_48138,N_48932);
xnor UO_4817 (O_4817,N_49226,N_47436);
xnor UO_4818 (O_4818,N_47316,N_47948);
xnor UO_4819 (O_4819,N_45763,N_48593);
or UO_4820 (O_4820,N_47545,N_47684);
and UO_4821 (O_4821,N_46488,N_47848);
and UO_4822 (O_4822,N_48870,N_46239);
nand UO_4823 (O_4823,N_45337,N_48962);
nor UO_4824 (O_4824,N_49479,N_47824);
or UO_4825 (O_4825,N_49919,N_49701);
xnor UO_4826 (O_4826,N_48167,N_49234);
or UO_4827 (O_4827,N_47996,N_46737);
or UO_4828 (O_4828,N_49808,N_45213);
and UO_4829 (O_4829,N_49529,N_49914);
nor UO_4830 (O_4830,N_45402,N_45199);
or UO_4831 (O_4831,N_45916,N_45383);
nor UO_4832 (O_4832,N_49361,N_46017);
nor UO_4833 (O_4833,N_46845,N_49848);
nor UO_4834 (O_4834,N_49371,N_47320);
xor UO_4835 (O_4835,N_49616,N_47642);
nand UO_4836 (O_4836,N_48288,N_48185);
and UO_4837 (O_4837,N_46210,N_47766);
and UO_4838 (O_4838,N_49777,N_47075);
nand UO_4839 (O_4839,N_46975,N_48961);
nand UO_4840 (O_4840,N_46157,N_49484);
or UO_4841 (O_4841,N_48297,N_47637);
xor UO_4842 (O_4842,N_46366,N_45870);
nand UO_4843 (O_4843,N_49331,N_48104);
xor UO_4844 (O_4844,N_48996,N_48253);
or UO_4845 (O_4845,N_47627,N_47679);
or UO_4846 (O_4846,N_47930,N_47368);
or UO_4847 (O_4847,N_47457,N_47637);
nand UO_4848 (O_4848,N_47373,N_45611);
or UO_4849 (O_4849,N_47165,N_45564);
nor UO_4850 (O_4850,N_46910,N_46163);
nor UO_4851 (O_4851,N_47426,N_45950);
xor UO_4852 (O_4852,N_49573,N_45033);
and UO_4853 (O_4853,N_46672,N_45717);
xor UO_4854 (O_4854,N_46785,N_47808);
and UO_4855 (O_4855,N_46369,N_48556);
xnor UO_4856 (O_4856,N_47289,N_49596);
nor UO_4857 (O_4857,N_46173,N_48290);
xnor UO_4858 (O_4858,N_47213,N_49296);
or UO_4859 (O_4859,N_49472,N_49528);
and UO_4860 (O_4860,N_47069,N_47157);
and UO_4861 (O_4861,N_46958,N_45957);
nand UO_4862 (O_4862,N_46255,N_46244);
xor UO_4863 (O_4863,N_48170,N_45054);
or UO_4864 (O_4864,N_48071,N_46616);
and UO_4865 (O_4865,N_48353,N_47539);
nor UO_4866 (O_4866,N_49011,N_47358);
or UO_4867 (O_4867,N_49518,N_45732);
xnor UO_4868 (O_4868,N_47447,N_48129);
and UO_4869 (O_4869,N_47079,N_46801);
or UO_4870 (O_4870,N_48180,N_48135);
xor UO_4871 (O_4871,N_48885,N_46741);
xor UO_4872 (O_4872,N_49638,N_47491);
xnor UO_4873 (O_4873,N_45198,N_45087);
nand UO_4874 (O_4874,N_46404,N_48246);
and UO_4875 (O_4875,N_46537,N_49851);
or UO_4876 (O_4876,N_45286,N_46554);
and UO_4877 (O_4877,N_47369,N_48756);
and UO_4878 (O_4878,N_49206,N_49942);
and UO_4879 (O_4879,N_45339,N_49976);
xnor UO_4880 (O_4880,N_45203,N_46071);
nand UO_4881 (O_4881,N_48619,N_47161);
nor UO_4882 (O_4882,N_45739,N_49180);
or UO_4883 (O_4883,N_48441,N_48284);
and UO_4884 (O_4884,N_49096,N_49277);
or UO_4885 (O_4885,N_46721,N_47390);
and UO_4886 (O_4886,N_45453,N_49677);
xnor UO_4887 (O_4887,N_49643,N_49628);
nand UO_4888 (O_4888,N_48234,N_47557);
xor UO_4889 (O_4889,N_48158,N_49043);
nor UO_4890 (O_4890,N_47663,N_46442);
and UO_4891 (O_4891,N_45640,N_47484);
and UO_4892 (O_4892,N_49493,N_45272);
nor UO_4893 (O_4893,N_49091,N_48801);
nand UO_4894 (O_4894,N_46664,N_49496);
nand UO_4895 (O_4895,N_45080,N_45529);
nand UO_4896 (O_4896,N_48779,N_49225);
or UO_4897 (O_4897,N_49166,N_49999);
nand UO_4898 (O_4898,N_45039,N_47420);
and UO_4899 (O_4899,N_46274,N_45792);
and UO_4900 (O_4900,N_49267,N_47603);
nand UO_4901 (O_4901,N_45381,N_45240);
nand UO_4902 (O_4902,N_48686,N_48957);
nor UO_4903 (O_4903,N_46705,N_48862);
nor UO_4904 (O_4904,N_46596,N_48725);
or UO_4905 (O_4905,N_49443,N_46390);
nand UO_4906 (O_4906,N_47082,N_46144);
xnor UO_4907 (O_4907,N_45087,N_48069);
or UO_4908 (O_4908,N_46475,N_49824);
and UO_4909 (O_4909,N_49738,N_48188);
nand UO_4910 (O_4910,N_49719,N_49477);
nor UO_4911 (O_4911,N_48992,N_48576);
or UO_4912 (O_4912,N_47805,N_46979);
xor UO_4913 (O_4913,N_49225,N_48368);
nand UO_4914 (O_4914,N_48262,N_48765);
xor UO_4915 (O_4915,N_49611,N_46909);
nand UO_4916 (O_4916,N_48139,N_48381);
nor UO_4917 (O_4917,N_46421,N_48884);
nor UO_4918 (O_4918,N_46753,N_47890);
or UO_4919 (O_4919,N_46188,N_47163);
nor UO_4920 (O_4920,N_48349,N_46707);
nor UO_4921 (O_4921,N_47925,N_47680);
nor UO_4922 (O_4922,N_46697,N_49670);
nand UO_4923 (O_4923,N_49923,N_49439);
nor UO_4924 (O_4924,N_45627,N_48194);
xor UO_4925 (O_4925,N_47826,N_49109);
nand UO_4926 (O_4926,N_48041,N_48293);
nor UO_4927 (O_4927,N_49326,N_49620);
and UO_4928 (O_4928,N_47621,N_48228);
or UO_4929 (O_4929,N_45541,N_45401);
and UO_4930 (O_4930,N_45622,N_45183);
nand UO_4931 (O_4931,N_48600,N_45184);
nand UO_4932 (O_4932,N_45591,N_46414);
xor UO_4933 (O_4933,N_47815,N_47569);
nand UO_4934 (O_4934,N_45130,N_46692);
nor UO_4935 (O_4935,N_45304,N_45904);
and UO_4936 (O_4936,N_45465,N_49800);
or UO_4937 (O_4937,N_47321,N_47906);
nand UO_4938 (O_4938,N_49075,N_49602);
and UO_4939 (O_4939,N_47975,N_47917);
and UO_4940 (O_4940,N_47756,N_48421);
nor UO_4941 (O_4941,N_47211,N_48528);
xor UO_4942 (O_4942,N_45539,N_46667);
nor UO_4943 (O_4943,N_47533,N_47968);
and UO_4944 (O_4944,N_47601,N_48710);
or UO_4945 (O_4945,N_45607,N_49987);
xnor UO_4946 (O_4946,N_49491,N_45006);
nand UO_4947 (O_4947,N_46632,N_46607);
or UO_4948 (O_4948,N_47898,N_46602);
nor UO_4949 (O_4949,N_46177,N_48209);
nand UO_4950 (O_4950,N_46722,N_46582);
and UO_4951 (O_4951,N_45687,N_46281);
nor UO_4952 (O_4952,N_47426,N_49338);
xor UO_4953 (O_4953,N_46890,N_48779);
or UO_4954 (O_4954,N_48646,N_45873);
nor UO_4955 (O_4955,N_46028,N_46867);
and UO_4956 (O_4956,N_47842,N_45064);
and UO_4957 (O_4957,N_47803,N_49619);
or UO_4958 (O_4958,N_45160,N_47528);
nand UO_4959 (O_4959,N_45378,N_49556);
nand UO_4960 (O_4960,N_48263,N_47558);
and UO_4961 (O_4961,N_47853,N_49333);
nor UO_4962 (O_4962,N_49073,N_46381);
xor UO_4963 (O_4963,N_48985,N_47580);
and UO_4964 (O_4964,N_49089,N_45837);
or UO_4965 (O_4965,N_47084,N_45307);
and UO_4966 (O_4966,N_46892,N_47273);
nand UO_4967 (O_4967,N_48232,N_47008);
nand UO_4968 (O_4968,N_47683,N_48786);
and UO_4969 (O_4969,N_46637,N_45701);
nand UO_4970 (O_4970,N_47474,N_46370);
nand UO_4971 (O_4971,N_48315,N_47644);
xor UO_4972 (O_4972,N_45441,N_48715);
and UO_4973 (O_4973,N_47883,N_45781);
nand UO_4974 (O_4974,N_45321,N_45751);
or UO_4975 (O_4975,N_49321,N_46988);
and UO_4976 (O_4976,N_49790,N_45077);
or UO_4977 (O_4977,N_49496,N_45731);
xor UO_4978 (O_4978,N_49451,N_49344);
nand UO_4979 (O_4979,N_49105,N_45076);
and UO_4980 (O_4980,N_46188,N_47577);
nor UO_4981 (O_4981,N_48112,N_47415);
or UO_4982 (O_4982,N_47231,N_47436);
nor UO_4983 (O_4983,N_47581,N_47389);
and UO_4984 (O_4984,N_49576,N_46345);
nor UO_4985 (O_4985,N_48885,N_49337);
nand UO_4986 (O_4986,N_46437,N_49928);
nand UO_4987 (O_4987,N_48878,N_49181);
nand UO_4988 (O_4988,N_49086,N_48824);
nand UO_4989 (O_4989,N_45665,N_49230);
or UO_4990 (O_4990,N_45652,N_48177);
nor UO_4991 (O_4991,N_45915,N_47509);
nor UO_4992 (O_4992,N_46522,N_47236);
nand UO_4993 (O_4993,N_45536,N_45234);
or UO_4994 (O_4994,N_48356,N_47022);
or UO_4995 (O_4995,N_47481,N_47385);
xnor UO_4996 (O_4996,N_46230,N_45155);
and UO_4997 (O_4997,N_47684,N_48939);
xnor UO_4998 (O_4998,N_49245,N_48322);
xor UO_4999 (O_4999,N_48082,N_48105);
endmodule